

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4289, n4290, n4291, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374;

  AND2_X1 U4792 ( .A1(n8543), .A2(n8542), .ZN(n8755) );
  INV_X1 U4793 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10066) );
  NAND2_X1 U4794 ( .A1(n5369), .A2(n5368), .ZN(n9950) );
  NAND2_X1 U4795 ( .A1(n5694), .A2(n5693), .ZN(n9459) );
  INV_X1 U4796 ( .A(n7772), .ZN(n7809) );
  NAND2_X1 U4797 ( .A1(n9322), .A2(n9416), .ZN(n9240) );
  INV_X1 U4798 ( .A(n7767), .ZN(n7770) );
  NAND2_X1 U4799 ( .A1(n5159), .A2(n5158), .ZN(n9857) );
  BUF_X1 U4800 ( .A(n8948), .Z(n4293) );
  INV_X2 U4801 ( .A(n4294), .ZN(n7040) );
  NAND2_X1 U4802 ( .A1(n6209), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5817) );
  AND2_X1 U4803 ( .A1(n6685), .A2(n9267), .ZN(n6491) );
  BUF_X1 U4804 ( .A(n5890), .Z(n6007) );
  NAND2_X1 U4805 ( .A1(n5434), .A2(n5435), .ZN(n5458) );
  INV_X1 U4808 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X2 U4809 ( .B1(n6194), .B2(n8212), .A(n6183), .ZN(n8512) );
  NAND2_X1 U4810 ( .A1(n6687), .A2(n6686), .ZN(n6688) );
  NAND2_X1 U4812 ( .A1(n9950), .A2(n9219), .ZN(n9361) );
  NAND2_X1 U4813 ( .A1(n7770), .A2(n7882), .ZN(n8143) );
  OR2_X1 U4814 ( .A1(n5705), .A2(n5704), .ZN(n5715) );
  INV_X2 U4816 ( .A(n5241), .ZN(n6449) );
  AND2_X1 U4817 ( .A1(n7286), .A2(n9395), .ZN(n9384) );
  INV_X1 U4818 ( .A(n8270), .ZN(n7882) );
  AND2_X2 U4819 ( .A1(n6259), .A2(n8242), .ZN(n8245) );
  NAND2_X1 U4820 ( .A1(n6093), .A2(n6092), .ZN(n8636) );
  NAND2_X1 U4821 ( .A1(n8215), .A2(n8216), .ZN(n8212) );
  NAND2_X1 U4822 ( .A1(n6489), .A2(n4560), .ZN(n4446) );
  INV_X1 U4823 ( .A(n8273), .ZN(n7423) );
  INV_X1 U4824 ( .A(n8122), .ZN(n10151) );
  NAND2_X1 U4825 ( .A1(n6097), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  AND2_X1 U4826 ( .A1(n5491), .A2(n5472), .ZN(n5465) );
  NAND2_X1 U4828 ( .A1(n9348), .A2(n9257), .ZN(n9680) );
  AND2_X1 U4829 ( .A1(n9789), .A2(n4317), .ZN(n9723) );
  NAND2_X1 U4830 ( .A1(n9304), .A2(n9326), .ZN(n9804) );
  AND4_X1 U4831 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n7884)
         );
  XNOR2_X1 U4832 ( .A(n5817), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6213) );
  INV_X1 U4833 ( .A(n9965), .ZN(n9683) );
  AND4_X1 U4834 ( .A1(n5576), .A2(n5575), .A3(n5574), .A4(n5573), .ZN(n8828)
         );
  NAND2_X1 U4835 ( .A1(n6172), .A2(n6171), .ZN(n8520) );
  INV_X1 U4836 ( .A(n7452), .ZN(n7349) );
  INV_X1 U4837 ( .A(n6736), .ZN(n9470) );
  NAND2_X1 U4838 ( .A1(n5436), .A2(n5458), .ZN(n9267) );
  OR2_X2 U4840 ( .A1(n8157), .A2(n8267), .ZN(n8160) );
  NAND2_X2 U4841 ( .A1(n4446), .A2(n6024), .ZN(n8157) );
  NAND2_X2 U4842 ( .A1(n6781), .A2(n6780), .ZN(n9555) );
  NAND2_X1 U4843 ( .A1(n6585), .A2(n5859), .ZN(n5888) );
  OR2_X2 U4844 ( .A1(n9816), .A2(n5616), .ZN(n9817) );
  AOI21_X2 U4845 ( .B1(n5789), .B2(n9846), .A(n5788), .ZN(n6382) );
  NAND3_X2 U4846 ( .A1(n7482), .A2(n4578), .A3(n4577), .ZN(n4905) );
  INV_X1 U4847 ( .A(n5452), .ZN(n5030) );
  NAND2_X2 U4848 ( .A1(n7897), .A2(n7898), .ZN(n7896) );
  NAND2_X2 U4849 ( .A1(n7927), .A2(n7808), .ZN(n7897) );
  XNOR2_X2 U4850 ( .A(n5033), .B(n5032), .ZN(n7708) );
  NAND2_X2 U4851 ( .A1(n7994), .A2(n4404), .ZN(n4852) );
  NAND2_X2 U4852 ( .A1(n7896), .A2(n7812), .ZN(n7994) );
  AND2_X4 U4853 ( .A1(n4496), .A2(n4495), .ZN(n6585) );
  NAND2_X2 U4854 ( .A1(n5078), .A2(n5077), .ZN(n5122) );
  NAND3_X2 U4855 ( .A1(n5073), .A2(n5072), .A3(n5071), .ZN(n5078) );
  AOI211_X2 U4856 ( .C1(n9007), .C2(n9011), .A(n9010), .B(n8842), .ZN(n8843)
         );
  NAND2_X2 U4857 ( .A1(n5219), .A2(n5218), .ZN(n5226) );
  NAND2_X2 U4858 ( .A1(n4681), .A2(n5871), .ZN(n6851) );
  NAND2_X2 U4859 ( .A1(n5815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6096) );
  XNOR2_X2 U4860 ( .A(n6732), .B(n6731), .ZN(n6734) );
  BUF_X1 U4861 ( .A(n6685), .Z(n4300) );
  XNOR2_X1 U4862 ( .A(n5433), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6685) );
  XNOR2_X2 U4863 ( .A(n5846), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5852) );
  OAI22_X2 U4864 ( .A1(n8385), .A2(n8384), .B1(n8383), .B2(n8391), .ZN(n8404)
         );
  AOI22_X2 U4865 ( .A1(n8357), .A2(n8356), .B1(n8355), .B2(n8354), .ZN(n8385)
         );
  NAND2_X4 U4866 ( .A1(n6214), .A2(n6578), .ZN(n5858) );
  XNOR2_X2 U4867 ( .A(n5837), .B(n5842), .ZN(n6578) );
  OAI21_X2 U4868 ( .B1(n5220), .B2(SI_13_), .A(n5227), .ZN(n5224) );
  XNOR2_X1 U4869 ( .A(n8153), .B(n8268), .ZN(n8150) );
  NAND2_X2 U4870 ( .A1(n6011), .A2(n6010), .ZN(n8153) );
  OAI22_X2 U4871 ( .A1(n8332), .A2(n8331), .B1(n8330), .B2(n8329), .ZN(n8357)
         );
  AOI22_X2 U4872 ( .A1(n8307), .A2(n8306), .B1(n8305), .B2(n8304), .ZN(n8332)
         );
  NOR2_X4 U4873 ( .A1(n6714), .A2(n6713), .ZN(n6733) );
  INV_X1 U4874 ( .A(n8922), .ZN(n4289) );
  INV_X1 U4875 ( .A(n8922), .ZN(n4290) );
  OAI22_X2 U4876 ( .A1(n6733), .A2(n6734), .B1(n6732), .B2(n6731), .ZN(n7039)
         );
  OAI22_X2 U4877 ( .A1(n7145), .A2(n4653), .B1(n4655), .B2(n4652), .ZN(n8282)
         );
  NAND2_X1 U4878 ( .A1(n7723), .A2(n8177), .ZN(n8651) );
  NAND2_X1 U4879 ( .A1(n8160), .A2(n8161), .ZN(n8059) );
  NAND2_X1 U4880 ( .A1(n5767), .A2(n7233), .ZN(n7232) );
  NAND2_X1 U4881 ( .A1(n7532), .A2(n9467), .ZN(n5767) );
  INV_X2 U4882 ( .A(n7221), .ZN(n7532) );
  NAND2_X1 U4883 ( .A1(n5760), .A2(n9401), .ZN(n7251) );
  INV_X1 U4884 ( .A(n7542), .ZN(n7054) );
  NAND2_X2 U4885 ( .A1(n8080), .A2(n8088), .ZN(n7135) );
  NAND2_X2 U4886 ( .A1(n7330), .A2(n9470), .ZN(n9403) );
  INV_X1 U4887 ( .A(n9384), .ZN(n9382) );
  AND4_X1 U4888 ( .A1(n5523), .A2(n5522), .A3(n5521), .A4(n5520), .ZN(n6956)
         );
  INV_X1 U4889 ( .A(n8222), .ZN(n8235) );
  INV_X1 U4890 ( .A(n9474), .ZN(n4291) );
  CLKBUF_X2 U4891 ( .A(n5986), .Z(n6202) );
  BUF_X2 U4892 ( .A(n5511), .Z(n5782) );
  BUF_X1 U4893 ( .A(n5753), .Z(n4301) );
  XNOR2_X1 U4894 ( .A(n5467), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5753) );
  CLKBUF_X2 U4895 ( .A(n6218), .Z(n4297) );
  NAND2_X1 U4896 ( .A1(n5432), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U4897 ( .A1(n5849), .A2(n5848), .ZN(n5882) );
  NAND2_X2 U4898 ( .A1(n5056), .A2(n7708), .ZN(n5067) );
  CLKBUF_X2 U4899 ( .A(n5056), .Z(n7763) );
  AND3_X1 U4900 ( .A1(n5016), .A2(n5015), .A3(n5190), .ZN(n5022) );
  AND4_X1 U4901 ( .A1(n5828), .A2(n5827), .A3(n6095), .A4(n6242), .ZN(n5830)
         );
  NOR2_X1 U4902 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5808) );
  MUX2_X1 U4903 ( .A(n9868), .B(n9867), .S(n10117), .Z(n9869) );
  OAI21_X1 U4904 ( .B1(n6407), .B2(n6406), .A(n6405), .ZN(n6411) );
  AOI21_X1 U4905 ( .B1(n4372), .B2(n8345), .A(n4472), .ZN(n4447) );
  NAND2_X1 U4906 ( .A1(n9078), .A2(n8957), .ZN(n9195) );
  AND2_X1 U4907 ( .A1(n4731), .A2(n4730), .ZN(n8468) );
  AND2_X1 U4908 ( .A1(n4732), .A2(n8466), .ZN(n4730) );
  OR2_X1 U4909 ( .A1(n8446), .A2(n8445), .ZN(n4732) );
  NAND2_X1 U4910 ( .A1(n6142), .A2(n6141), .ZN(n8569) );
  AOI21_X1 U4911 ( .B1(n4769), .B2(n4768), .A(n4414), .ZN(n4767) );
  NAND2_X1 U4912 ( .A1(n8031), .A2(n8030), .ZN(n8742) );
  NAND2_X1 U4913 ( .A1(n8233), .A2(n8032), .ZN(n8227) );
  NAND2_X1 U4914 ( .A1(n8902), .A2(n9183), .ZN(n9026) );
  NAND2_X1 U4915 ( .A1(n8647), .A2(n8173), .ZN(n8626) );
  NAND2_X2 U4916 ( .A1(n9803), .A2(n5617), .ZN(n9788) );
  NAND2_X1 U4917 ( .A1(n8651), .A2(n8062), .ZN(n4705) );
  XNOR2_X1 U4918 ( .A(n5406), .B(SI_29_), .ZN(n8815) );
  NAND2_X2 U4919 ( .A1(n7435), .A2(n5593), .ZN(n7493) );
  NAND2_X1 U4920 ( .A1(n9064), .A2(n8860), .ZN(n9153) );
  INV_X1 U4921 ( .A(n9923), .ZN(n9307) );
  NAND2_X1 U4922 ( .A1(n4592), .A2(n4593), .ZN(n5371) );
  NAND2_X1 U4923 ( .A1(n6067), .A2(n6066), .ZN(n8737) );
  NAND2_X1 U4924 ( .A1(n5341), .A2(n5340), .ZN(n9667) );
  OR2_X1 U4925 ( .A1(n8287), .A2(n8298), .ZN(n8288) );
  NAND2_X1 U4926 ( .A1(n4468), .A2(n4467), .ZN(n5009) );
  AND2_X1 U4927 ( .A1(n5332), .A2(n5331), .ZN(n9965) );
  NAND2_X2 U4928 ( .A1(n7197), .A2(n5561), .ZN(n7228) );
  NAND2_X1 U4929 ( .A1(n5345), .A2(n5344), .ZN(n5353) );
  NOR2_X1 U4930 ( .A1(n4307), .A2(n4350), .ZN(n4854) );
  NAND2_X1 U4931 ( .A1(n6182), .A2(n6181), .ZN(n8572) );
  NAND2_X2 U4932 ( .A1(n5244), .A2(n5243), .ZN(n9929) );
  NAND2_X1 U4933 ( .A1(n4588), .A2(n4586), .ZN(n5326) );
  NAND2_X1 U4934 ( .A1(n7157), .A2(n7156), .ZN(n4723) );
  NAND2_X1 U4935 ( .A1(n5627), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5645) );
  OR2_X1 U4936 ( .A1(n7971), .A2(n7884), .ZN(n8147) );
  NAND2_X1 U4937 ( .A1(n5217), .A2(n5216), .ZN(n8856) );
  AND2_X1 U4938 ( .A1(n4343), .A2(n7150), .ZN(n7093) );
  OAI21_X1 U4939 ( .B1(n5253), .B2(SI_14_), .A(n5255), .ZN(n5236) );
  NAND2_X1 U4940 ( .A1(n5194), .A2(n5193), .ZN(n9019) );
  OR2_X1 U4941 ( .A1(n6764), .A2(n6765), .ZN(n4448) );
  NAND2_X1 U4942 ( .A1(n4445), .A2(n5206), .ZN(n5219) );
  NAND2_X2 U4943 ( .A1(n9280), .A2(n9403), .ZN(n5763) );
  NAND2_X1 U4944 ( .A1(n10151), .A2(n8274), .ZN(n8106) );
  NAND2_X1 U4945 ( .A1(n9471), .A2(n10111), .ZN(n9402) );
  CLKBUF_X2 U4946 ( .A(n6684), .Z(n10101) );
  AND2_X1 U4947 ( .A1(n5115), .A2(n5114), .ZN(n7542) );
  CLKBUF_X1 U4948 ( .A(n6851), .Z(n8277) );
  BUF_X2 U4949 ( .A(n6709), .Z(n8947) );
  NAND2_X1 U4950 ( .A1(n6448), .A2(n6674), .ZN(n10099) );
  XNOR2_X1 U4951 ( .A(n5171), .B(n5178), .ZN(n6453) );
  AND2_X1 U4952 ( .A1(n5147), .A2(n5140), .ZN(n6441) );
  AND4_X1 U4953 ( .A1(n5568), .A2(n5567), .A3(n5566), .A4(n5565), .ZN(n9137)
         );
  NAND4_X1 U4954 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n8270)
         );
  NAND2_X1 U4955 ( .A1(n4770), .A2(n6748), .ZN(n6874) );
  NAND2_X1 U4956 ( .A1(n5050), .A2(n4567), .ZN(n10073) );
  NAND2_X1 U4957 ( .A1(n4329), .A2(n5930), .ZN(n8274) );
  NAND2_X2 U4958 ( .A1(n6213), .A2(n8255), .ZN(n8222) );
  INV_X1 U4959 ( .A(n6014), .ZN(n6013) );
  NAND4_X2 U4960 ( .A1(n5508), .A2(n5507), .A3(n5506), .A4(n5505), .ZN(n9474)
         );
  CLKBUF_X3 U4961 ( .A(n5528), .Z(n5738) );
  AOI21_X1 U4962 ( .B1(n4921), .B2(n4923), .A(n4920), .ZN(n4919) );
  NAND2_X1 U4963 ( .A1(n6233), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U4964 ( .A1(n6209), .A2(n6208), .ZN(n8242) );
  CLKBUF_X1 U4965 ( .A(n8029), .Z(n4474) );
  BUF_X2 U4966 ( .A(n6218), .Z(n4298) );
  CLKBUF_X3 U4967 ( .A(n5882), .Z(n5971) );
  CLKBUF_X3 U4968 ( .A(n5141), .Z(n5422) );
  AOI21_X1 U4969 ( .B1(n5062), .B2(n6530), .A(n4568), .ZN(n4567) );
  OR2_X1 U4970 ( .A1(n5525), .A2(n5497), .ZN(n5501) );
  AND2_X1 U4971 ( .A1(n5504), .A2(n5445), .ZN(n5512) );
  INV_X1 U4972 ( .A(n4931), .ZN(n4928) );
  NAND2_X4 U4973 ( .A1(n7827), .A2(n5848), .ZN(n5957) );
  INV_X4 U4974 ( .A(n8477), .ZN(n8405) );
  INV_X1 U4975 ( .A(n6214), .ZN(n8477) );
  INV_X1 U4976 ( .A(n5445), .ZN(n9991) );
  OAI211_X1 U4977 ( .C1(n5301), .C2(n5300), .A(n5299), .B(n5298), .ZN(n5485)
         );
  AND2_X1 U4978 ( .A1(n5461), .A2(n4321), .ZN(n5472) );
  NOR2_X1 U4979 ( .A1(n5105), .A2(n5104), .ZN(n5123) );
  OR2_X1 U4980 ( .A1(n5571), .A2(n5570), .ZN(n5579) );
  MUX2_X1 U4981 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5440), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5441) );
  OR2_X1 U4982 ( .A1(n5442), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n9986) );
  XNOR2_X1 U4983 ( .A(n5031), .B(n5439), .ZN(n5056) );
  NOR2_X1 U4984 ( .A1(n4544), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9990) );
  NOR2_X2 U4985 ( .A1(n6047), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U4986 ( .A1(n6237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U4987 ( .A1(n4461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5031) );
  NAND2_X1 U4988 ( .A1(n5150), .A2(n4545), .ZN(n5168) );
  NAND2_X1 U4989 ( .A1(n5098), .A2(SI_5_), .ZN(n5125) );
  NAND2_X1 U4990 ( .A1(n5463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5033) );
  NOR2_X2 U4991 ( .A1(n5084), .A2(n5083), .ZN(n9488) );
  OR2_X1 U4992 ( .A1(n5925), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5942) );
  AND2_X1 U4993 ( .A1(n5029), .A2(n4423), .ZN(n4422) );
  NAND2_X1 U4994 ( .A1(n5030), .A2(n5029), .ZN(n5463) );
  AND2_X1 U4995 ( .A1(n5029), .A2(n4957), .ZN(n4424) );
  BUF_X2 U4996 ( .A(n5149), .Z(n4543) );
  INV_X1 U4997 ( .A(n5931), .ZN(n4438) );
  NAND4_X2 U4998 ( .A1(n5080), .A2(n5022), .A3(n5021), .A4(n5153), .ZN(n5452)
         );
  NAND2_X1 U4999 ( .A1(n5537), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5556) );
  AND2_X1 U5000 ( .A1(n5018), .A2(n5017), .ZN(n5021) );
  NOR2_X1 U5001 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5020) );
  NOR2_X1 U5002 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5015) );
  NOR2_X1 U5003 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5018) );
  NOR2_X1 U5004 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5019) );
  NOR2_X1 U5005 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5016) );
  NOR2_X1 U5006 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5017) );
  INV_X1 U5007 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7482) );
  INV_X1 U5008 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5190) );
  INV_X1 U5009 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5952) );
  INV_X4 U5010 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5011 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5435) );
  INV_X1 U5012 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6095) );
  INV_X1 U5013 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5820) );
  INV_X1 U5014 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5814) );
  INV_X1 U5015 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4904) );
  INV_X1 U5016 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4577) );
  INV_X1 U5017 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4578) );
  INV_X1 U5018 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5827) );
  INV_X1 U5019 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6242) );
  NOR2_X2 U5020 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5034) );
  INV_X1 U5021 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7130) );
  OR2_X1 U5022 ( .A1(n6232), .A2(n6231), .ZN(n6234) );
  AND2_X1 U5023 ( .A1(n6852), .A2(n6928), .ZN(n6853) );
  OAI22_X2 U5024 ( .A1(n8282), .A2(n8281), .B1(n8280), .B2(n8279), .ZN(n8307)
         );
  INV_X4 U5025 ( .A(n8964), .ZN(n9034) );
  BUF_X4 U5026 ( .A(n8948), .Z(n4294) );
  OAI22_X2 U5028 ( .A1(n9153), .A2(n4819), .B1(n4368), .B2(n8872), .ZN(n9087)
         );
  AOI21_X2 U5029 ( .B1(n7696), .B2(n6046), .A(n6045), .ZN(n7730) );
  INV_X1 U5030 ( .A(n5960), .ZN(n4295) );
  CLKBUF_X1 U5031 ( .A(n6218), .Z(n4296) );
  INV_X1 U5032 ( .A(n5939), .ZN(n6218) );
  INV_X1 U5033 ( .A(n4862), .ZN(n7760) );
  OAI21_X1 U5034 ( .B1(n7752), .B2(n7648), .A(n4863), .ZN(n4862) );
  OR2_X1 U5035 ( .A1(n7827), .A2(n5852), .ZN(n5939) );
  AOI21_X1 U5036 ( .B1(n4626), .B2(n9360), .A(n4625), .ZN(n4624) );
  INV_X1 U5037 ( .A(n9357), .ZN(n4625) );
  INV_X1 U5038 ( .A(n5218), .ZN(n4923) );
  NAND2_X1 U5039 ( .A1(n5381), .A2(n5380), .ZN(n5396) );
  INV_X1 U5040 ( .A(n4597), .ZN(n4596) );
  OAI21_X1 U5041 ( .B1(n5352), .B2(n4598), .A(n5361), .ZN(n4597) );
  INV_X1 U5042 ( .A(n6491), .ZN(n4431) );
  AND2_X1 U5043 ( .A1(n9237), .A2(n9443), .ZN(n6676) );
  AOI21_X1 U5044 ( .B1(n9635), .B2(n9354), .A(n4628), .ZN(n4514) );
  OR2_X1 U5045 ( .A1(n5746), .A2(n7022), .ZN(n9378) );
  NAND2_X1 U5046 ( .A1(n4299), .A2(n5790), .ZN(n9394) );
  INV_X1 U5047 ( .A(n5971), .ZN(n6216) );
  INV_X1 U5048 ( .A(n4688), .ZN(n4687) );
  AOI21_X1 U5049 ( .B1(n4688), .B2(n4686), .A(n4371), .ZN(n4685) );
  AND2_X1 U5050 ( .A1(n4689), .A2(n8223), .ZN(n4688) );
  OR2_X1 U5051 ( .A1(n8751), .A2(n8533), .ZN(n8223) );
  AND2_X1 U5052 ( .A1(n4301), .A2(n4300), .ZN(n9237) );
  INV_X1 U5053 ( .A(n5546), .ZN(n5781) );
  AND2_X1 U5054 ( .A1(n5471), .A2(n6678), .ZN(n6448) );
  AND2_X1 U5055 ( .A1(n6677), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5471) );
  NAND2_X1 U5056 ( .A1(n8149), .A2(n8150), .ZN(n4674) );
  NOR2_X1 U5057 ( .A1(n9414), .A2(n4638), .ZN(n4637) );
  NAND2_X1 U5058 ( .A1(n9416), .A2(n9302), .ZN(n4638) );
  AOI21_X1 U5059 ( .B1(n4914), .B2(n4915), .A(n4910), .ZN(n4420) );
  NAND2_X1 U5060 ( .A1(n4539), .A2(n8217), .ZN(n4536) );
  NOR2_X1 U5061 ( .A1(n8226), .A2(n8227), .ZN(n4667) );
  INV_X1 U5062 ( .A(n6152), .ZN(n4892) );
  OAI21_X1 U5063 ( .B1(n4623), .B2(n4626), .A(n4364), .ZN(n4622) );
  AOI21_X1 U5064 ( .B1(n9356), .B2(n5778), .A(n9355), .ZN(n9365) );
  INV_X1 U5065 ( .A(n5011), .ZN(n4840) );
  NOR2_X1 U5066 ( .A1(n5005), .A2(n5452), .ZN(n4430) );
  OAI21_X1 U5067 ( .B1(n4919), .B2(n4304), .A(n5267), .ZN(n4602) );
  NAND2_X1 U5068 ( .A1(n5269), .A2(n5268), .ZN(n5274) );
  NOR2_X1 U5069 ( .A1(n8230), .A2(n8231), .ZN(n4678) );
  NAND2_X1 U5070 ( .A1(n8297), .A2(n8296), .ZN(n4773) );
  NAND2_X1 U5071 ( .A1(n4767), .A2(n8451), .ZN(n4760) );
  NAND2_X1 U5072 ( .A1(n6184), .A2(n10249), .ZN(n6197) );
  OR2_X1 U5073 ( .A1(n8726), .A2(n8659), .ZN(n8173) );
  AND2_X1 U5074 ( .A1(n7767), .A2(n8270), .ZN(n8132) );
  AND2_X1 U5075 ( .A1(n6295), .A2(n8553), .ZN(n8206) );
  OR2_X1 U5076 ( .A1(n7854), .A2(n8638), .ZN(n8594) );
  AND2_X1 U5077 ( .A1(n8594), .A2(n8188), .ZN(n8625) );
  OR2_X1 U5078 ( .A1(n8800), .A2(n8637), .ZN(n8062) );
  NOR2_X1 U5079 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5831) );
  AOI21_X1 U5080 ( .B1(n8993), .B2(n9164), .A(n8995), .ZN(n8932) );
  NOR2_X1 U5081 ( .A1(n4344), .A2(n4824), .ZN(n4823) );
  AOI21_X1 U5082 ( .B1(n9437), .B2(n9232), .A(n9435), .ZN(n9234) );
  NAND2_X1 U5083 ( .A1(n9997), .A2(n9991), .ZN(n5525) );
  NAND2_X1 U5084 ( .A1(n4436), .A2(n4435), .ZN(n5429) );
  INV_X1 U5085 ( .A(n5452), .ZN(n4436) );
  OR2_X1 U5086 ( .A1(n8981), .A2(n9199), .ZN(n9358) );
  AOI21_X1 U5087 ( .B1(n4564), .B2(n4975), .A(n4359), .ZN(n4563) );
  OR2_X1 U5088 ( .A1(n9929), .A2(n9811), .ZN(n9306) );
  AND2_X1 U5089 ( .A1(n5769), .A2(n9284), .ZN(n9412) );
  AOI21_X1 U5090 ( .B1(n9298), .B2(n9293), .A(n9296), .ZN(n5769) );
  NAND2_X1 U5091 ( .A1(n4524), .A2(n4523), .ZN(n9249) );
  INV_X1 U5092 ( .A(n9292), .ZN(n4523) );
  NOR2_X1 U5093 ( .A1(n5768), .A2(n9278), .ZN(n4524) );
  NAND2_X1 U5094 ( .A1(n4967), .A2(n4966), .ZN(n9802) );
  AOI21_X1 U5095 ( .B1(n4968), .B2(n4970), .A(n4362), .ZN(n4966) );
  NAND2_X1 U5096 ( .A1(n7493), .A2(n4968), .ZN(n4967) );
  AOI21_X1 U5097 ( .B1(n10099), .B2(n5486), .A(n6676), .ZN(n5749) );
  OAI21_X1 U5098 ( .B1(n5407), .B2(n5406), .A(n5405), .ZN(n5417) );
  AND2_X1 U5099 ( .A1(n5363), .A2(n5358), .ZN(n5361) );
  OAI21_X1 U5100 ( .B1(n5326), .B2(n5325), .A(n5324), .ZN(n5335) );
  INV_X1 U5101 ( .A(n5316), .ZN(n5322) );
  NAND2_X1 U5102 ( .A1(n4603), .A2(n4919), .ZN(n5253) );
  AND2_X1 U5103 ( .A1(n4908), .A2(n4909), .ZN(n5179) );
  INV_X2 U5104 ( .A(n5116), .ZN(n5149) );
  AND2_X1 U5105 ( .A1(n6304), .A2(n6266), .ZN(n6819) );
  NAND2_X1 U5106 ( .A1(n4751), .A2(n4748), .ZN(n4747) );
  OR2_X1 U5107 ( .A1(n7292), .A2(n7300), .ZN(n7293) );
  OAI22_X1 U5108 ( .A1(n4767), .A2(n8451), .B1(n8418), .B2(n4764), .ZN(n8459)
         );
  NAND2_X1 U5109 ( .A1(n4765), .A2(n4768), .ZN(n4764) );
  NAND2_X1 U5110 ( .A1(n4761), .A2(n8462), .ZN(n8463) );
  INV_X1 U5111 ( .A(n4762), .ZN(n4761) );
  OAI21_X1 U5112 ( .B1(n4760), .B2(n4759), .A(n4757), .ZN(n4762) );
  AOI21_X1 U5113 ( .B1(n4767), .B2(n4411), .A(n4758), .ZN(n4757) );
  NAND2_X1 U5114 ( .A1(n6240), .A2(n6239), .ZN(n6813) );
  AOI21_X1 U5115 ( .B1(n4879), .B2(n4878), .A(n4361), .ZN(n4877) );
  INV_X1 U5116 ( .A(n6124), .ZN(n4878) );
  NAND3_X1 U5117 ( .A1(n5861), .A2(n5860), .A3(n4333), .ZN(n5862) );
  OR2_X1 U5118 ( .A1(n6404), .A2(n6403), .ZN(n6842) );
  AND2_X1 U5119 ( .A1(n10144), .A2(n8245), .ZN(n6399) );
  NAND2_X1 U5120 ( .A1(n8223), .A2(n8224), .ZN(n8516) );
  NAND2_X1 U5121 ( .A1(n6193), .A2(n6192), .ZN(n8751) );
  NAND2_X1 U5122 ( .A1(n8519), .A2(n8571), .ZN(n8522) );
  NAND2_X1 U5123 ( .A1(n6297), .A2(n8199), .ZN(n6408) );
  OR2_X1 U5124 ( .A1(n8222), .A2(n6824), .ZN(n8658) );
  OR2_X1 U5125 ( .A1(n8222), .A2(n6855), .ZN(n8656) );
  INV_X1 U5126 ( .A(n8658), .ZN(n8571) );
  INV_X1 U5127 ( .A(n8656), .ZN(n8573) );
  AND2_X1 U5128 ( .A1(n6847), .A2(n7288), .ZN(n10144) );
  OR2_X1 U5129 ( .A1(n8222), .A2(n6299), .ZN(n6856) );
  AND2_X1 U5130 ( .A1(n6819), .A2(n6820), .ZN(n6858) );
  AND2_X1 U5131 ( .A1(n6813), .A2(n6486), .ZN(n6820) );
  NOR2_X1 U5132 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4900) );
  NAND2_X1 U5133 ( .A1(n6096), .A2(n4858), .ZN(n6209) );
  AND2_X1 U5134 ( .A1(n5816), .A2(n4859), .ZN(n4858) );
  INV_X1 U5135 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4859) );
  INV_X1 U5136 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4495) );
  INV_X1 U5137 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4496) );
  AOI21_X1 U5138 ( .B1(n9110), .B2(n4817), .A(n4816), .ZN(n4815) );
  INV_X1 U5139 ( .A(n9111), .ZN(n4817) );
  INV_X1 U5140 ( .A(n8943), .ZN(n4816) );
  INV_X1 U5141 ( .A(n9457), .ZN(n9198) );
  NAND2_X1 U5142 ( .A1(n9267), .A2(n9765), .ZN(n9443) );
  AOI21_X2 U5143 ( .B1(n9685), .B2(n5738), .A(n5683), .ZN(n9055) );
  INV_X1 U5144 ( .A(n5782), .ZN(n5736) );
  INV_X1 U5145 ( .A(n5738), .ZN(n5725) );
  INV_X1 U5146 ( .A(n5525), .ZN(n5511) );
  AND2_X1 U5147 ( .A1(n9991), .A2(n5504), .ZN(n5528) );
  OR2_X1 U5148 ( .A1(n5723), .A2(n8978), .ZN(n5793) );
  NOR2_X1 U5149 ( .A1(n4508), .A2(n9620), .ZN(n4506) );
  INV_X1 U5150 ( .A(n4514), .ZN(n4508) );
  AND2_X1 U5151 ( .A1(n4341), .A2(n5695), .ZN(n4971) );
  NAND2_X1 U5152 ( .A1(n5774), .A2(n4351), .ZN(n9738) );
  INV_X1 U5153 ( .A(n9740), .ZN(n5775) );
  AOI21_X1 U5154 ( .B1(n9807), .B2(n4942), .A(n4941), .ZN(n4940) );
  INV_X1 U5155 ( .A(n9326), .ZN(n4941) );
  NAND2_X1 U5156 ( .A1(n7493), .A2(n9240), .ZN(n7494) );
  XNOR2_X1 U5157 ( .A(n5444), .B(n5443), .ZN(n5445) );
  INV_X1 U5158 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5443) );
  NAND2_X1 U5159 ( .A1(n4421), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5444) );
  NAND2_X1 U5160 ( .A1(n5030), .A2(n4422), .ZN(n4421) );
  NAND2_X1 U5161 ( .A1(n5458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5433) );
  NAND2_X1 U5162 ( .A1(n5840), .A2(n5839), .ZN(n8505) );
  NAND2_X1 U5163 ( .A1(n8545), .A2(n6216), .ZN(n6172) );
  XNOR2_X1 U5164 ( .A(n5470), .B(n5469), .ZN(n6678) );
  NAND2_X1 U5165 ( .A1(n6702), .A2(n9852), .ZN(n9215) );
  NAND2_X1 U5166 ( .A1(n8108), .A2(n8222), .ZN(n8119) );
  NAND2_X1 U5167 ( .A1(n8114), .A2(n8113), .ZN(n8117) );
  INV_X1 U5168 ( .A(n8142), .ZN(n4675) );
  INV_X1 U5169 ( .A(n4674), .ZN(n4672) );
  OR2_X1 U5170 ( .A1(n4673), .A2(n4674), .ZN(n4669) );
  INV_X1 U5171 ( .A(n8151), .ZN(n4673) );
  NOR2_X1 U5172 ( .A1(n9804), .A2(n4942), .ZN(n4925) );
  INV_X1 U5173 ( .A(n4634), .ZN(n4633) );
  INV_X1 U5174 ( .A(n9314), .ZN(n4643) );
  AOI21_X1 U5175 ( .B1(n8654), .B2(n4347), .A(n4311), .ZN(n4548) );
  NOR2_X1 U5176 ( .A1(n4345), .A2(n9384), .ZN(n4505) );
  NOR2_X1 U5177 ( .A1(n4520), .A2(n4521), .ZN(n4912) );
  NOR2_X1 U5178 ( .A1(n4614), .A2(n4613), .ZN(n4610) );
  NAND2_X1 U5179 ( .A1(n4918), .A2(n4312), .ZN(n4614) );
  OAI21_X1 U5180 ( .B1(n4615), .B2(n4613), .A(n4617), .ZN(n4612) );
  INV_X1 U5181 ( .A(n9350), .ZN(n4617) );
  AOI21_X1 U5182 ( .B1(n4918), .B2(n4616), .A(n4917), .ZN(n4615) );
  NAND2_X1 U5183 ( .A1(n4684), .A2(n8193), .ZN(n8202) );
  OAI21_X1 U5184 ( .B1(n8187), .B2(n8186), .A(n8191), .ZN(n4684) );
  NOR2_X1 U5185 ( .A1(n4536), .A2(n4356), .ZN(n4535) );
  NAND2_X1 U5186 ( .A1(n8202), .A2(n8598), .ZN(n8197) );
  AND2_X1 U5187 ( .A1(n4667), .A2(n4538), .ZN(n4537) );
  AND2_X1 U5188 ( .A1(n7362), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4744) );
  NOR2_X1 U5189 ( .A1(n8512), .A2(n4892), .ZN(n4891) );
  INV_X1 U5190 ( .A(n6141), .ZN(n4884) );
  NAND2_X1 U5191 ( .A1(n4890), .A2(n4888), .ZN(n4887) );
  NOR2_X1 U5192 ( .A1(n4889), .A2(n4892), .ZN(n4888) );
  OR2_X1 U5193 ( .A1(n9154), .A2(n4821), .ZN(n4820) );
  AND2_X1 U5194 ( .A1(n9378), .A2(n9366), .ZN(n4607) );
  NAND2_X1 U5195 ( .A1(n4607), .A2(n4606), .ZN(n9230) );
  INV_X1 U5196 ( .A(n9363), .ZN(n4606) );
  AOI21_X1 U5197 ( .B1(n4621), .B2(n4623), .A(n4620), .ZN(n4619) );
  INV_X1 U5198 ( .A(n9359), .ZN(n4620) );
  NAND2_X1 U5199 ( .A1(n4808), .A2(n9870), .ZN(n4807) );
  INV_X1 U5200 ( .A(n5354), .ZN(n4598) );
  OAI21_X1 U5201 ( .B1(n6430), .B2(P1_DATAO_REG_7__SCAN_IN), .A(n5134), .ZN(
        n5136) );
  OR2_X1 U5202 ( .A1(n5149), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n5134) );
  OAI211_X1 U5203 ( .C1(n5116), .C2(P1_DATAO_REG_0__SCAN_IN), .A(n4516), .B(
        SI_0_), .ZN(n5041) );
  NOR2_X1 U5204 ( .A1(n4839), .A2(n4366), .ZN(n4838) );
  NOR2_X1 U5205 ( .A1(n4841), .A2(n4840), .ZN(n4839) );
  NAND2_X1 U5206 ( .A1(n4838), .A2(n4840), .ZN(n4836) );
  AND2_X1 U5207 ( .A1(n7796), .A2(n7870), .ZN(n7797) );
  AND2_X1 U5208 ( .A1(n7775), .A2(n7886), .ZN(n7776) );
  OR2_X1 U5209 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  NOR2_X1 U5210 ( .A1(n8516), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U5211 ( .A1(n8540), .A2(n4719), .ZN(n4718) );
  OR2_X1 U5212 ( .A1(n8342), .A2(n8341), .ZN(n8343) );
  AND2_X1 U5213 ( .A1(n8393), .A2(n8392), .ZN(n8394) );
  OR2_X1 U5214 ( .A1(n8380), .A2(n8388), .ZN(n8381) );
  NAND2_X1 U5215 ( .A1(n8422), .A2(n4494), .ZN(n8425) );
  OR2_X1 U5216 ( .A1(n8424), .A2(n8423), .ZN(n4494) );
  NAND2_X1 U5217 ( .A1(n8239), .A2(n8519), .ZN(n4689) );
  OR2_X1 U5218 ( .A1(n6197), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7753) );
  INV_X1 U5219 ( .A(n6269), .ZN(n5910) );
  OR2_X1 U5220 ( .A1(n6261), .A2(n6258), .ZN(n6303) );
  OR2_X1 U5221 ( .A1(n8769), .A2(n7850), .ZN(n8199) );
  OR2_X1 U5222 ( .A1(n8706), .A2(n8608), .ZN(n8201) );
  OR2_X1 U5223 ( .A1(n8002), .A2(n7838), .ZN(n8169) );
  NAND2_X1 U5224 ( .A1(n6034), .A2(n4871), .ZN(n4869) );
  NAND2_X1 U5225 ( .A1(n6006), .A2(n4872), .ZN(n4871) );
  AND2_X1 U5226 ( .A1(n7622), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U5227 ( .A1(n6033), .A2(n6006), .ZN(n4870) );
  NAND2_X1 U5228 ( .A1(n7644), .A2(n5993), .ZN(n7597) );
  NOR2_X1 U5229 ( .A1(n8132), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5230 ( .A1(n8147), .A2(n8148), .ZN(n7768) );
  NAND2_X1 U5231 ( .A1(n9117), .A2(n7047), .ZN(n7050) );
  AOI21_X1 U5232 ( .B1(n7321), .B2(n4305), .A(n4831), .ZN(n4830) );
  NOR2_X1 U5233 ( .A1(n7579), .A2(n7580), .ZN(n4831) );
  OR2_X1 U5234 ( .A1(n4291), .A2(n4294), .ZN(n6493) );
  OR2_X1 U5235 ( .A1(n9374), .A2(n9376), .ZN(n4934) );
  INV_X1 U5236 ( .A(n9997), .ZN(n5504) );
  NOR2_X1 U5237 ( .A1(n10005), .A2(n4458), .ZN(n9567) );
  AND2_X1 U5238 ( .A1(n10006), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n4458) );
  NOR2_X1 U5239 ( .A1(n5746), .A2(n4807), .ZN(n4806) );
  NAND2_X1 U5240 ( .A1(n4331), .A2(n5722), .ZN(n4987) );
  NOR2_X1 U5241 ( .A1(n9259), .A2(n4989), .ZN(n4988) );
  INV_X1 U5242 ( .A(n5722), .ZN(n4989) );
  OR2_X1 U5243 ( .A1(n9045), .A2(n9031), .ZN(n9366) );
  NOR2_X1 U5244 ( .A1(n9667), .A2(n4800), .ZN(n4799) );
  INV_X1 U5245 ( .A(n4801), .ZN(n4800) );
  NAND2_X1 U5246 ( .A1(n4517), .A2(n4346), .ZN(n9223) );
  NAND2_X1 U5247 ( .A1(n4519), .A2(n4522), .ZN(n4518) );
  INV_X1 U5248 ( .A(n5636), .ZN(n4976) );
  NOR2_X1 U5249 ( .A1(n8845), .A2(n4795), .ZN(n4794) );
  INV_X1 U5250 ( .A(n4796), .ZN(n4795) );
  NAND2_X1 U5251 ( .A1(n4499), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5603) );
  INV_X1 U5252 ( .A(n5595), .ZN(n4499) );
  NAND2_X1 U5253 ( .A1(n5577), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5587) );
  INV_X1 U5254 ( .A(n5579), .ZN(n5577) );
  OR2_X1 U5255 ( .A1(n8830), .A2(n8828), .ZN(n9316) );
  OAI211_X1 U5256 ( .C1(n5396), .C2(n5395), .A(n5394), .B(n4585), .ZN(n5406)
         );
  NAND2_X1 U5257 ( .A1(n5396), .A2(n4399), .ZN(n4585) );
  NAND2_X1 U5258 ( .A1(n5373), .A2(n5372), .ZN(n5381) );
  INV_X1 U5259 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5454) );
  NOR2_X2 U5260 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5453) );
  AND2_X1 U5261 ( .A1(n5354), .A2(n5349), .ZN(n5352) );
  NOR2_X2 U5262 ( .A1(n5429), .A2(n5428), .ZN(n5434) );
  AOI21_X1 U5263 ( .B1(n4589), .B2(n4591), .A(n4587), .ZN(n4586) );
  INV_X1 U5264 ( .A(n5306), .ZN(n4587) );
  INV_X1 U5265 ( .A(n5287), .ZN(n4591) );
  INV_X1 U5266 ( .A(n4602), .ZN(n4601) );
  NOR2_X1 U5267 ( .A1(n4922), .A2(n4304), .ZN(n4600) );
  OAI21_X1 U5268 ( .B1(n6430), .B2(P1_DATAO_REG_9__SCAN_IN), .A(n4486), .ZN(
        n5181) );
  NAND2_X1 U5269 ( .A1(n6430), .A2(n6454), .ZN(n4486) );
  INV_X1 U5270 ( .A(n5186), .ZN(n5185) );
  NAND2_X1 U5271 ( .A1(n7685), .A2(n8271), .ZN(n4484) );
  INV_X1 U5272 ( .A(n4855), .ZN(n7456) );
  NOR2_X1 U5273 ( .A1(n4326), .A2(n4861), .ZN(n4860) );
  NAND2_X1 U5274 ( .A1(n5896), .A2(n7130), .ZN(n5913) );
  NAND2_X1 U5275 ( .A1(n7421), .A2(n4856), .ZN(n4855) );
  NOR2_X1 U5276 ( .A1(n7458), .A2(n4857), .ZN(n4856) );
  INV_X1 U5277 ( .A(n7420), .ZN(n4857) );
  AND3_X1 U5278 ( .A1(n7860), .A2(n7861), .A3(n7859), .ZN(n7869) );
  NAND2_X1 U5279 ( .A1(n6104), .A2(n4715), .ZN(n6128) );
  NAND2_X1 U5280 ( .A1(n7959), .A2(n7960), .ZN(n7958) );
  INV_X1 U5281 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n4714) );
  XNOR2_X1 U5282 ( .A(n6854), .B(n10126), .ZN(n6895) );
  NAND2_X1 U5283 ( .A1(n7023), .A2(n7009), .ZN(n4482) );
  NAND2_X1 U5284 ( .A1(n4552), .A2(n4551), .ZN(n8246) );
  NAND2_X1 U5285 ( .A1(n4676), .A2(n4330), .ZN(n4551) );
  AOI21_X1 U5286 ( .B1(n8238), .B2(n8239), .A(n8237), .ZN(n4676) );
  BUF_X1 U5287 ( .A(n5939), .Z(n8022) );
  NAND2_X1 U5288 ( .A1(n6057), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5883) );
  OR2_X1 U5289 ( .A1(n5939), .A2(n5847), .ZN(n5857) );
  OR2_X1 U5290 ( .A1(n5957), .A2(n10157), .ZN(n5871) );
  OAI22_X1 U5291 ( .A1(n5939), .A2(n7137), .B1(n5870), .B2(n5882), .ZN(n4682)
         );
  OAI21_X1 U5292 ( .B1(n6606), .B2(n6586), .A(n6618), .ZN(n6587) );
  NOR2_X1 U5293 ( .A1(n6587), .A2(n7137), .ZN(n6620) );
  AOI21_X1 U5294 ( .B1(n6581), .B2(n6580), .A(n6611), .ZN(n6582) );
  XNOR2_X1 U5295 ( .A(n6607), .B(n6606), .ZN(n6575) );
  NAND3_X1 U5296 ( .A1(n6663), .A2(n6747), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n6750) );
  OR2_X1 U5297 ( .A1(n6875), .A2(n6966), .ZN(n5001) );
  NOR2_X1 U5298 ( .A1(n4755), .A2(n4749), .ZN(n6979) );
  NAND2_X1 U5299 ( .A1(n4753), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4749) );
  NAND2_X1 U5300 ( .A1(n7099), .A2(n7098), .ZN(n7155) );
  NAND2_X1 U5301 ( .A1(n4725), .A2(n7143), .ZN(n4724) );
  AND3_X1 U5302 ( .A1(n4724), .A2(n7155), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n7158) );
  NAND2_X1 U5303 ( .A1(n7299), .A2(n4306), .ZN(n4785) );
  NAND2_X1 U5304 ( .A1(n7299), .A2(n7298), .ZN(n4777) );
  INV_X1 U5305 ( .A(n7308), .ZN(n4660) );
  NOR2_X1 U5306 ( .A1(n7300), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4782) );
  AND2_X1 U5307 ( .A1(n4781), .A2(n4779), .ZN(n4778) );
  CLKBUF_X1 U5308 ( .A(n5818), .Z(n5819) );
  NAND2_X1 U5309 ( .A1(n4736), .A2(n4740), .ZN(n8365) );
  INV_X1 U5310 ( .A(n4760), .ZN(n4756) );
  NAND2_X1 U5311 ( .A1(n8425), .A2(n4765), .ZN(n8446) );
  NAND2_X1 U5312 ( .A1(n6102), .A2(n6101), .ZN(n7854) );
  AND2_X1 U5313 ( .A1(n6112), .A2(n6094), .ZN(n4901) );
  INV_X1 U5314 ( .A(n8625), .ZN(n6112) );
  NAND2_X1 U5315 ( .A1(n6104), .A2(n6103), .ZN(n6116) );
  AOI21_X1 U5316 ( .B1(n4875), .B2(n8171), .A(n4357), .ZN(n4874) );
  NAND2_X1 U5317 ( .A1(n7718), .A2(n4338), .ZN(n4873) );
  NAND2_X1 U5318 ( .A1(n6052), .A2(n4711), .ZN(n6085) );
  AND2_X1 U5319 ( .A1(n4318), .A2(n4712), .ZN(n4711) );
  INV_X1 U5320 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n4712) );
  NAND2_X1 U5321 ( .A1(n7718), .A2(n6290), .ZN(n7721) );
  NAND2_X1 U5322 ( .A1(n6052), .A2(n6051), .ZN(n6068) );
  NAND2_X1 U5323 ( .A1(n5973), .A2(n5972), .ZN(n5987) );
  INV_X1 U5324 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5972) );
  INV_X1 U5325 ( .A(n5974), .ZN(n5973) );
  NAND2_X1 U5326 ( .A1(n7189), .A2(n5949), .ZN(n4898) );
  NAND2_X1 U5327 ( .A1(n5941), .A2(n5940), .ZN(n5958) );
  INV_X1 U5328 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5940) );
  INV_X1 U5329 ( .A(n5942), .ZN(n5941) );
  AND2_X1 U5330 ( .A1(n6296), .A2(n8198), .ZN(n4702) );
  AND2_X1 U5331 ( .A1(n8769), .A2(n8572), .ZN(n8551) );
  NAND2_X1 U5332 ( .A1(n8579), .A2(n8203), .ZN(n4703) );
  OR2_X1 U5333 ( .A1(n8703), .A2(n8591), .ZN(n8198) );
  OR2_X1 U5334 ( .A1(n8711), .A2(n8621), .ZN(n8595) );
  NAND2_X1 U5335 ( .A1(n7721), .A2(n6073), .ZN(n8652) );
  AND2_X1 U5336 ( .A1(n6091), .A2(n6090), .ZN(n8659) );
  AND3_X1 U5337 ( .A1(n6072), .A2(n6071), .A3(n6070), .ZN(n8657) );
  NOR2_X1 U5338 ( .A1(n6284), .A2(n4696), .ZN(n4695) );
  INV_X1 U5339 ( .A(n7768), .ZN(n8058) );
  AND2_X1 U5340 ( .A1(n6238), .A2(n6237), .ZN(n6246) );
  NAND2_X1 U5341 ( .A1(n5834), .A2(n5833), .ZN(n6235) );
  NOR2_X1 U5342 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), .ZN(
        n4849) );
  NAND2_X1 U5343 ( .A1(n6063), .A2(n5814), .ZN(n6074) );
  NAND2_X1 U5344 ( .A1(n4476), .A2(n4475), .ZN(n4832) );
  INV_X1 U5345 ( .A(n7215), .ZN(n4475) );
  INV_X1 U5346 ( .A(n7216), .ZN(n4476) );
  AND2_X1 U5347 ( .A1(n8968), .A2(n8967), .ZN(n9046) );
  AOI21_X1 U5348 ( .B1(n7040), .B2(n10090), .A(n4466), .ZN(n6496) );
  AND2_X1 U5349 ( .A1(n6495), .A2(n4469), .ZN(n4466) );
  NAND2_X1 U5350 ( .A1(n9051), .A2(n8921), .ZN(n8992) );
  NAND2_X1 U5351 ( .A1(n8891), .A2(n8893), .ZN(n8894) );
  INV_X1 U5352 ( .A(n5539), .ZN(n5537) );
  NAND2_X1 U5353 ( .A1(n8999), .A2(n4815), .ZN(n4813) );
  INV_X1 U5354 ( .A(n9080), .ZN(n4812) );
  AND3_X1 U5355 ( .A1(n5533), .A2(n5532), .A3(n5531), .ZN(n6736) );
  AND2_X1 U5356 ( .A1(n5530), .A2(n5529), .ZN(n5531) );
  AND2_X1 U5357 ( .A1(n9259), .A2(n9361), .ZN(n4953) );
  NAND2_X1 U5358 ( .A1(n5714), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U5359 ( .A1(n9647), .A2(n9351), .ZN(n9631) );
  NAND2_X1 U5360 ( .A1(n9631), .A2(n9635), .ZN(n9630) );
  NAND2_X1 U5361 ( .A1(n9349), .A2(n9257), .ZN(n4947) );
  OR2_X1 U5362 ( .A1(n4949), .A2(n5776), .ZN(n4946) );
  AND2_X1 U5363 ( .A1(n9664), .A2(n4950), .ZN(n4949) );
  NAND2_X1 U5364 ( .A1(n4951), .A2(n9257), .ZN(n4950) );
  INV_X1 U5365 ( .A(n9348), .ZN(n4951) );
  NAND2_X1 U5366 ( .A1(n9679), .A2(n9348), .ZN(n4948) );
  AOI21_X1 U5367 ( .B1(n4980), .B2(n4979), .A(n4370), .ZN(n4978) );
  AND2_X1 U5368 ( .A1(n9340), .A2(n9428), .ZN(n9729) );
  NAND2_X1 U5369 ( .A1(n9757), .A2(n4342), .ZN(n5774) );
  NAND2_X1 U5370 ( .A1(n4939), .A2(n4352), .ZN(n9794) );
  NAND2_X1 U5371 ( .A1(n9838), .A2(n4940), .ZN(n4939) );
  NAND2_X1 U5372 ( .A1(n4940), .A2(n9804), .ZN(n4938) );
  AND2_X1 U5373 ( .A1(n9306), .A2(n9327), .ZN(n9796) );
  NAND2_X1 U5374 ( .A1(n7495), .A2(n9416), .ZN(n9839) );
  INV_X1 U5375 ( .A(n4969), .ZN(n4968) );
  OAI21_X1 U5376 ( .B1(n9240), .B2(n4970), .A(n9827), .ZN(n4969) );
  INV_X1 U5377 ( .A(n5601), .ZN(n4970) );
  NAND2_X1 U5378 ( .A1(n5772), .A2(n4956), .ZN(n7495) );
  AND2_X1 U5379 ( .A1(n5773), .A2(n9318), .ZN(n4956) );
  NAND2_X1 U5380 ( .A1(n7436), .A2(n9241), .ZN(n7435) );
  INV_X1 U5381 ( .A(n9250), .ZN(n5770) );
  NAND2_X1 U5382 ( .A1(n9412), .A2(n7065), .ZN(n4952) );
  NAND2_X1 U5383 ( .A1(n5769), .A2(n9249), .ZN(n9410) );
  NAND2_X1 U5384 ( .A1(n4569), .A2(n4962), .ZN(n7276) );
  AOI21_X1 U5385 ( .B1(n4963), .B2(n4965), .A(n4360), .ZN(n4962) );
  NAND2_X1 U5386 ( .A1(n7228), .A2(n4963), .ZN(n4569) );
  INV_X1 U5387 ( .A(n9841), .ZN(n9808) );
  INV_X1 U5388 ( .A(n5569), .ZN(n4965) );
  INV_X1 U5389 ( .A(n4964), .ZN(n4963) );
  OAI21_X1 U5390 ( .B1(n7236), .B2(n4965), .A(n7384), .ZN(n4964) );
  NAND2_X1 U5391 ( .A1(n7228), .A2(n7236), .ZN(n7229) );
  NAND2_X1 U5392 ( .A1(n4958), .A2(n4570), .ZN(n7197) );
  INV_X1 U5393 ( .A(n4571), .ZN(n4570) );
  OAI21_X1 U5394 ( .B1(n7199), .B2(n4961), .A(n7232), .ZN(n4571) );
  NAND2_X1 U5395 ( .A1(n4937), .A2(n4935), .ZN(n9275) );
  NOR2_X1 U5396 ( .A1(n5762), .A2(n4936), .ZN(n4935) );
  INV_X1 U5397 ( .A(n9279), .ZN(n4936) );
  AND2_X1 U5398 ( .A1(n6801), .A2(n7263), .ZN(n7177) );
  AND2_X1 U5399 ( .A1(n9237), .A2(n6517), .ZN(n9841) );
  AND2_X1 U5400 ( .A1(n9237), .A2(n7763), .ZN(n9843) );
  INV_X1 U5401 ( .A(n9846), .ZN(n9761) );
  INV_X1 U5402 ( .A(n9843), .ZN(n9810) );
  INV_X1 U5403 ( .A(n5067), .ZN(n5062) );
  CLKBUF_X1 U5404 ( .A(n5067), .Z(n5241) );
  AND2_X1 U5405 ( .A1(n5492), .A2(n9985), .ZN(n6672) );
  NAND2_X1 U5406 ( .A1(n5360), .A2(n5359), .ZN(n9637) );
  INV_X1 U5407 ( .A(n5423), .ZN(n5397) );
  AND2_X1 U5408 ( .A1(n5749), .A2(n5488), .ZN(n5804) );
  AND2_X1 U5409 ( .A1(n5463), .A2(n5464), .ZN(n5487) );
  MUX2_X1 U5410 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5462), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5464) );
  AND2_X1 U5411 ( .A1(n5344), .A2(n5339), .ZN(n5342) );
  XNOR2_X1 U5412 ( .A(n5245), .B(n5237), .ZN(n6727) );
  XNOR2_X1 U5413 ( .A(n5253), .B(n5228), .ZN(n6593) );
  OR2_X1 U5414 ( .A1(n5214), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5229) );
  NOR2_X1 U5415 ( .A1(n5173), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5212) );
  OR2_X1 U5416 ( .A1(n5156), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5173) );
  BUF_X1 U5417 ( .A(n5080), .Z(n5154) );
  NAND2_X1 U5418 ( .A1(n5055), .A2(n4902), .ZN(n5049) );
  INV_X1 U5419 ( .A(n8751), .ZN(n7834) );
  INV_X1 U5420 ( .A(n7833), .ZN(n4464) );
  NOR2_X1 U5421 ( .A1(n7828), .A2(n4851), .ZN(n4850) );
  INV_X1 U5422 ( .A(n4853), .ZN(n4851) );
  NAND2_X1 U5423 ( .A1(n6827), .A2(n8643), .ZN(n7998) );
  INV_X1 U5424 ( .A(n7998), .ZN(n8015) );
  NAND4_X2 U5425 ( .A1(n5866), .A2(n5865), .A3(n5864), .A4(n5863), .ZN(n8278)
         );
  NOR2_X1 U5426 ( .A1(n4651), .A2(n4650), .ZN(n4649) );
  INV_X1 U5427 ( .A(n6659), .ZN(n4650) );
  INV_X1 U5428 ( .A(n6648), .ZN(n4651) );
  AND2_X1 U5429 ( .A1(n4319), .A2(n7293), .ZN(n7364) );
  XNOR2_X1 U5430 ( .A(n5984), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8295) );
  XNOR2_X1 U5431 ( .A(n6009), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8338) );
  OR2_X2 U5432 ( .A1(n6813), .A2(n6426), .ZN(n8457) );
  AOI21_X1 U5433 ( .B1(n8484), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8458), .ZN(
        n4663) );
  NAND2_X1 U5434 ( .A1(n4320), .A2(n4664), .ZN(n4473) );
  AOI21_X1 U5435 ( .B1(n6344), .B2(n8640), .A(n4864), .ZN(n4863) );
  INV_X1 U5436 ( .A(n6351), .ZN(n4864) );
  NOR2_X1 U5437 ( .A1(n6224), .A2(n6223), .ZN(n6225) );
  NOR2_X1 U5438 ( .A1(n8533), .A2(n8656), .ZN(n6224) );
  AND2_X1 U5439 ( .A1(n8634), .A2(n8042), .ZN(n4704) );
  AND2_X1 U5440 ( .A1(n8663), .A2(n6409), .ZN(n8678) );
  NAND2_X1 U5441 ( .A1(n6399), .A2(n6820), .ZN(n8643) );
  AND2_X1 U5442 ( .A1(n10168), .A2(n10144), .ZN(n8733) );
  NAND2_X1 U5443 ( .A1(n4690), .A2(n8223), .ZN(n6329) );
  NAND2_X1 U5444 ( .A1(n8522), .A2(n8521), .ZN(n8523) );
  OR2_X1 U5445 ( .A1(n6826), .A2(n6311), .ZN(n6312) );
  AND2_X1 U5446 ( .A1(n4900), .A2(n4390), .ZN(n4679) );
  INV_X1 U5447 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4680) );
  INV_X1 U5448 ( .A(n7181), .ZN(n10111) );
  AND4_X1 U5449 ( .A1(n5592), .A2(n5591), .A3(n5590), .A4(n5589), .ZN(n9072)
         );
  NAND2_X1 U5450 ( .A1(n4814), .A2(n9110), .ZN(n9114) );
  NAND2_X1 U5451 ( .A1(n9112), .A2(n9111), .ZN(n4814) );
  INV_X1 U5452 ( .A(n9210), .ZN(n9165) );
  AND2_X1 U5453 ( .A1(n6698), .A2(n6696), .ZN(n9196) );
  AND3_X1 U5454 ( .A1(n5633), .A2(n5632), .A3(n5631), .ZN(n9764) );
  NOR2_X1 U5455 ( .A1(n4335), .A2(n9395), .ZN(n4584) );
  INV_X1 U5456 ( .A(n9452), .ZN(n4581) );
  NAND2_X1 U5457 ( .A1(n5700), .A2(n5699), .ZN(n9458) );
  OR2_X1 U5458 ( .A1(n9669), .A2(n5725), .ZN(n5694) );
  OAI21_X1 U5459 ( .B1(n10070), .B2(n9595), .A(n9594), .ZN(n4490) );
  NOR2_X1 U5460 ( .A1(n5437), .A2(n9832), .ZN(n9596) );
  NAND2_X1 U5461 ( .A1(n9635), .A2(n9620), .ZN(n4513) );
  NAND2_X1 U5462 ( .A1(n5751), .A2(n6448), .ZN(n9852) );
  NAND2_X1 U5463 ( .A1(n9267), .A2(n9395), .ZN(n10088) );
  NAND2_X1 U5464 ( .A1(n9950), .A2(n9899), .ZN(n4576) );
  AOI21_X1 U5465 ( .B1(n6381), .B2(n6380), .A(n4997), .ZN(n6383) );
  OR2_X1 U5466 ( .A1(n6381), .A2(n6374), .ZN(n6384) );
  NOR2_X1 U5467 ( .A1(n6413), .A2(n9981), .ZN(n6415) );
  OAI21_X1 U5468 ( .B1(n7751), .B2(n9943), .A(n6364), .ZN(n6368) );
  NAND2_X1 U5469 ( .A1(n6326), .A2(n9950), .ZN(n4527) );
  NAND2_X1 U5470 ( .A1(n9872), .A2(n4528), .ZN(n9949) );
  INV_X1 U5471 ( .A(n4529), .ZN(n4528) );
  OAI21_X1 U5472 ( .B1(n9873), .B2(n9943), .A(n9871), .ZN(n4529) );
  INV_X1 U5473 ( .A(n9409), .ZN(n4641) );
  OAI21_X1 U5474 ( .B1(n4639), .B2(n4636), .A(n9419), .ZN(n4634) );
  INV_X1 U5475 ( .A(n9416), .ZN(n4636) );
  AND2_X1 U5476 ( .A1(n4401), .A2(n4640), .ZN(n4639) );
  NAND2_X1 U5477 ( .A1(n4642), .A2(n4641), .ZN(n4640) );
  OAI21_X1 U5478 ( .B1(n9301), .B2(n9300), .A(n9299), .ZN(n9317) );
  OAI21_X1 U5479 ( .B1(n4670), .B2(n4367), .A(n4671), .ZN(n4558) );
  NAND2_X1 U5480 ( .A1(n8118), .A2(n8119), .ZN(n4670) );
  NAND2_X1 U5481 ( .A1(n8159), .A2(n8160), .ZN(n4554) );
  AND2_X1 U5482 ( .A1(n4669), .A2(n8156), .ZN(n4668) );
  INV_X1 U5483 ( .A(n8163), .ZN(n4557) );
  NAND2_X1 U5484 ( .A1(n8168), .A2(n8167), .ZN(n8178) );
  NAND2_X1 U5485 ( .A1(n4556), .A2(n4555), .ZN(n8168) );
  INV_X1 U5486 ( .A(n8166), .ZN(n4555) );
  OAI21_X1 U5487 ( .B1(n4553), .B2(n4558), .A(n4369), .ZN(n4556) );
  INV_X1 U5488 ( .A(n4924), .ZN(n9309) );
  OR2_X1 U5489 ( .A1(n4916), .A2(n9313), .ZN(n4915) );
  AOI21_X1 U5490 ( .B1(n4924), .B2(n4348), .A(n4643), .ZN(n4916) );
  INV_X1 U5491 ( .A(n9760), .ZN(n4910) );
  INV_X1 U5492 ( .A(n9680), .ZN(n4918) );
  AND2_X1 U5493 ( .A1(n9347), .A2(n9382), .ZN(n4917) );
  INV_X1 U5494 ( .A(n9346), .ZN(n4616) );
  AOI21_X1 U5495 ( .B1(n4548), .B2(n8171), .A(n4373), .ZN(n4547) );
  INV_X1 U5496 ( .A(n8221), .ZN(n4539) );
  NAND2_X1 U5497 ( .A1(n4376), .A2(n8217), .ZN(n4531) );
  NAND2_X1 U5498 ( .A1(n4379), .A2(n8217), .ZN(n4530) );
  INV_X1 U5499 ( .A(n4363), .ZN(n4627) );
  INV_X1 U5500 ( .A(n4612), .ZN(n4611) );
  OAI21_X1 U5501 ( .B1(n9343), .B2(n9342), .A(n4365), .ZN(n4504) );
  INV_X1 U5502 ( .A(SI_16_), .ZN(n5257) );
  INV_X1 U5503 ( .A(n6153), .ZN(n4889) );
  INV_X1 U5504 ( .A(n8512), .ZN(n4890) );
  AOI22_X1 U5505 ( .A1(n10300), .A2(n5258), .B1(n5259), .B2(n5257), .ZN(n5254)
         );
  OAI211_X1 U5506 ( .C1(n4542), .C2(n4532), .A(n4302), .B(n4534), .ZN(n8229)
         );
  NAND2_X1 U5507 ( .A1(n8213), .A2(n4535), .ZN(n4534) );
  INV_X1 U5508 ( .A(n8073), .ZN(n4719) );
  OR2_X1 U5509 ( .A1(n8212), .A2(n8563), .ZN(n4721) );
  OR2_X1 U5510 ( .A1(n8737), .A2(n8657), .ZN(n8179) );
  INV_X1 U5511 ( .A(n5993), .ZN(n4872) );
  INV_X1 U5512 ( .A(n8921), .ZN(n4824) );
  AOI211_X1 U5513 ( .C1(n9365), .C2(n4629), .A(n9364), .B(n9363), .ZN(n9368)
         );
  OR2_X1 U5514 ( .A1(n9968), .A2(n8917), .ZN(n9344) );
  NOR2_X1 U5515 ( .A1(n9019), .A2(n8830), .ZN(n4796) );
  INV_X1 U5516 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5025) );
  NOR2_X1 U5517 ( .A1(n5305), .A2(n4590), .ZN(n4589) );
  INV_X1 U5518 ( .A(n5290), .ZN(n4590) );
  INV_X1 U5519 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5426) );
  INV_X1 U5520 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5277) );
  INV_X1 U5521 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5278) );
  INV_X1 U5522 ( .A(n5256), .ZN(n5258) );
  INV_X1 U5523 ( .A(n5227), .ZN(n4920) );
  NAND2_X1 U5524 ( .A1(n5220), .A2(SI_13_), .ZN(n5227) );
  NAND2_X1 U5525 ( .A1(n5149), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n4545) );
  OR2_X1 U5526 ( .A1(n5149), .A2(n5148), .ZN(n5150) );
  INV_X1 U5527 ( .A(n7804), .ZN(n4861) );
  AND2_X1 U5528 ( .A1(n6103), .A2(n4716), .ZN(n4715) );
  INV_X1 U5529 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n4716) );
  INV_X1 U5530 ( .A(n6303), .ZN(n6307) );
  NAND2_X1 U5531 ( .A1(n5853), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5854) );
  NOR2_X1 U5532 ( .A1(n6887), .A2(n4750), .ZN(n4748) );
  INV_X1 U5533 ( .A(n6977), .ZN(n4750) );
  OR2_X1 U5534 ( .A1(n4306), .A2(n7569), .ZN(n4781) );
  NAND2_X1 U5535 ( .A1(n4780), .A2(n7300), .ZN(n4779) );
  INV_X1 U5536 ( .A(n7298), .ZN(n4780) );
  OAI211_X1 U5537 ( .C1(n4743), .C2(n4742), .A(n4745), .B(n4741), .ZN(n8287)
         );
  NAND2_X1 U5538 ( .A1(n7361), .A2(n4744), .ZN(n4743) );
  INV_X1 U5539 ( .A(n7293), .ZN(n4742) );
  INV_X1 U5540 ( .A(n8418), .ZN(n4759) );
  INV_X1 U5541 ( .A(n8224), .ZN(n4686) );
  INV_X1 U5542 ( .A(n4891), .ZN(n4885) );
  AND2_X1 U5543 ( .A1(n4886), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U5544 ( .A1(n4891), .A2(n4884), .ZN(n4883) );
  NAND2_X1 U5545 ( .A1(n8611), .A2(n6124), .ZN(n4881) );
  INV_X1 U5546 ( .A(n6105), .ZN(n6104) );
  INV_X1 U5547 ( .A(n6073), .ZN(n4875) );
  INV_X1 U5548 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n4713) );
  INV_X1 U5549 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6051) );
  INV_X1 U5550 ( .A(n6053), .ZN(n6052) );
  NOR2_X1 U5551 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_12__SCAN_IN), 
        .ZN(n4710) );
  NAND2_X1 U5552 ( .A1(n6851), .A2(n10122), .ZN(n8080) );
  OR2_X1 U5553 ( .A1(n8756), .A2(n7991), .ZN(n8067) );
  AND2_X1 U5554 ( .A1(n8756), .A2(n7991), .ZN(n8219) );
  INV_X1 U5555 ( .A(n8147), .ZN(n4694) );
  INV_X1 U5556 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5821) );
  INV_X1 U5557 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4899) );
  NOR2_X1 U5558 ( .A1(n5645), .A2(n5644), .ZN(n4501) );
  NAND2_X1 U5559 ( .A1(n4830), .A2(n4828), .ZN(n4827) );
  INV_X1 U5560 ( .A(n9008), .ZN(n4828) );
  NAND2_X1 U5561 ( .A1(n8867), .A2(n4822), .ZN(n4819) );
  OAI211_X1 U5562 ( .C1(n9230), .C2(n9231), .A(n4605), .B(n4604), .ZN(n9435)
         );
  NAND2_X1 U5563 ( .A1(n4607), .A2(n9367), .ZN(n4604) );
  NOR2_X1 U5564 ( .A1(n9229), .A2(n4327), .ZN(n4605) );
  NOR2_X1 U5565 ( .A1(n9683), .A2(n9968), .ZN(n4801) );
  INV_X1 U5566 ( .A(n4324), .ZN(n4979) );
  AND2_X1 U5567 ( .A1(n9344), .A2(n9345), .ZN(n9239) );
  INV_X1 U5568 ( .A(n9729), .ZN(n4522) );
  AOI21_X1 U5569 ( .B1(n9729), .B2(n4521), .A(n4520), .ZN(n4519) );
  NAND2_X1 U5570 ( .A1(n9771), .A2(n9778), .ZN(n9757) );
  NAND2_X1 U5571 ( .A1(n4456), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5620) );
  INV_X1 U5572 ( .A(n5610), .ZN(n4456) );
  NAND2_X1 U5573 ( .A1(n4457), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5610) );
  INV_X1 U5574 ( .A(n5603), .ZN(n4457) );
  NAND2_X1 U5575 ( .A1(n4500), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5595) );
  INV_X1 U5576 ( .A(n5587), .ZN(n4500) );
  NAND2_X1 U5577 ( .A1(n5562), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5571) );
  INV_X1 U5578 ( .A(n5563), .ZN(n5562) );
  INV_X1 U5579 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U5580 ( .A1(n5553), .A2(n5552), .ZN(n5563) );
  AND2_X1 U5581 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n5552) );
  INV_X1 U5582 ( .A(n5556), .ZN(n5553) );
  INV_X1 U5583 ( .A(n5551), .ZN(n4961) );
  NOR2_X1 U5584 ( .A1(n4961), .A2(n4960), .ZN(n4959) );
  INV_X1 U5585 ( .A(n5545), .ZN(n4960) );
  NAND2_X1 U5586 ( .A1(n4492), .A2(n4493), .ZN(n7252) );
  INV_X1 U5587 ( .A(n7254), .ZN(n4492) );
  INV_X1 U5588 ( .A(n7251), .ZN(n4493) );
  INV_X1 U5589 ( .A(n4807), .ZN(n4805) );
  NAND2_X1 U5590 ( .A1(n9695), .A2(n9697), .ZN(n9696) );
  NAND2_X1 U5591 ( .A1(n7379), .A2(n4794), .ZN(n7499) );
  NAND2_X1 U5592 ( .A1(n7379), .A2(n9142), .ZN(n7378) );
  AND2_X1 U5593 ( .A1(n4957), .A2(n4632), .ZN(n4423) );
  INV_X1 U5594 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4632) );
  NOR2_X1 U5595 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n4957) );
  NAND2_X1 U5596 ( .A1(n5396), .A2(n5393), .ZN(n5401) );
  AND2_X1 U5597 ( .A1(n5393), .A2(n5377), .ZN(n5380) );
  AOI21_X1 U5598 ( .B1(n4596), .B2(n4598), .A(n4594), .ZN(n4593) );
  INV_X1 U5599 ( .A(n5363), .ZN(n4594) );
  INV_X1 U5600 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5427) );
  NAND2_X1 U5601 ( .A1(n4932), .A2(n5195), .ZN(n4931) );
  NAND2_X1 U5602 ( .A1(n5137), .A2(SI_7_), .ZN(n5162) );
  NAND2_X1 U5603 ( .A1(n5122), .A2(n5121), .ZN(n5128) );
  INV_X1 U5604 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5014) );
  INV_X1 U5605 ( .A(n5042), .ZN(n5040) );
  INV_X1 U5606 ( .A(n5068), .ZN(n4902) );
  NAND2_X1 U5607 ( .A1(n7958), .A2(n7804), .ZN(n7846) );
  NAND2_X1 U5608 ( .A1(n7991), .A2(n7992), .ZN(n4853) );
  AND2_X1 U5609 ( .A1(n4836), .A2(n7797), .ZN(n4835) );
  AOI21_X1 U5610 ( .B1(n7776), .B2(n4354), .A(n4313), .ZN(n4847) );
  INV_X1 U5611 ( .A(n7776), .ZN(n4848) );
  INV_X1 U5612 ( .A(n4846), .ZN(n7883) );
  NAND2_X1 U5613 ( .A1(n4837), .A2(n5011), .ZN(n7856) );
  NAND2_X1 U5614 ( .A1(n8004), .A2(n4841), .ZN(n4837) );
  NAND2_X1 U5615 ( .A1(n5912), .A2(n5911), .ZN(n5925) );
  INV_X1 U5616 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5911) );
  INV_X1 U5617 ( .A(n5913), .ZN(n5912) );
  OR2_X1 U5618 ( .A1(n6305), .A2(n10144), .ZN(n6807) );
  AOI21_X1 U5619 ( .B1(n8071), .B2(n6847), .A(n8070), .ZN(n8243) );
  AND2_X1 U5620 ( .A1(n8234), .A2(n8069), .ZN(n4717) );
  AND2_X1 U5621 ( .A1(n8027), .A2(n8026), .ZN(n8076) );
  OR2_X1 U5622 ( .A1(n5986), .A2(n5924), .ZN(n5929) );
  NAND2_X1 U5623 ( .A1(n5853), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5863) );
  OAI21_X1 U5624 ( .B1(n8477), .B2(n10157), .A(n4450), .ZN(n6607) );
  NAND2_X1 U5625 ( .A1(n8477), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4450) );
  NOR2_X1 U5626 ( .A1(n6752), .A2(n6656), .ZN(n6657) );
  AND2_X1 U5627 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  NAND2_X1 U5628 ( .A1(n6750), .A2(n6747), .ZN(n4770) );
  INV_X1 U5629 ( .A(n4755), .ZN(n4752) );
  NAND2_X1 U5630 ( .A1(n4448), .A2(n4314), .ZN(n4647) );
  INV_X1 U5631 ( .A(n6882), .ZN(n4648) );
  AOI21_X1 U5632 ( .B1(n6971), .B2(n4776), .A(n4417), .ZN(n4774) );
  NAND2_X1 U5633 ( .A1(n4413), .A2(n5001), .ZN(n6972) );
  NOR2_X1 U5634 ( .A1(n6965), .A2(n4644), .ZN(n6969) );
  NOR2_X1 U5635 ( .A1(n4645), .A2(n6887), .ZN(n4644) );
  INV_X1 U5636 ( .A(n6967), .ZN(n4645) );
  NAND2_X1 U5637 ( .A1(n4481), .A2(n6585), .ZN(n5931) );
  AND2_X1 U5638 ( .A1(n5813), .A2(n5812), .ZN(n4481) );
  NOR2_X1 U5639 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5812) );
  NOR2_X1 U5640 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5813) );
  INV_X1 U5641 ( .A(n7155), .ZN(n7157) );
  OR2_X1 U5642 ( .A1(n5983), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5994) );
  INV_X1 U5643 ( .A(n7358), .ZN(n4656) );
  NAND2_X1 U5644 ( .A1(n4785), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4784) );
  NAND2_X1 U5645 ( .A1(n4772), .A2(n8305), .ZN(n4771) );
  AOI21_X1 U5646 ( .B1(n8358), .B2(n4789), .A(n4418), .ZN(n4788) );
  NAND2_X1 U5647 ( .A1(n4395), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n8359) );
  NOR2_X1 U5648 ( .A1(n8394), .A2(n8402), .ZN(n8414) );
  NAND2_X1 U5649 ( .A1(n4471), .A2(n4727), .ZN(n8422) );
  AOI21_X1 U5650 ( .B1(n8408), .B2(n4728), .A(n4419), .ZN(n4727) );
  NAND2_X1 U5651 ( .A1(n4332), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n8409) );
  OAI22_X1 U5652 ( .A1(n8432), .A2(n8431), .B1(n8430), .B2(n8438), .ZN(n8453)
         );
  NOR2_X1 U5653 ( .A1(n8482), .A2(n8475), .ZN(n4664) );
  OAI21_X1 U5654 ( .B1(n8476), .B2(n8475), .A(n8474), .ZN(n8481) );
  AND2_X1 U5655 ( .A1(n6579), .A2(n8819), .ZN(n6596) );
  NOR2_X1 U5656 ( .A1(n7818), .A2(n8658), .ZN(n6223) );
  AND2_X1 U5657 ( .A1(n6156), .A2(n4707), .ZN(n4706) );
  INV_X1 U5658 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n4707) );
  AOI21_X1 U5659 ( .B1(n8583), .B2(n6216), .A(n6140), .ZN(n8591) );
  AOI21_X1 U5660 ( .B1(n8600), .B2(n6216), .A(n6133), .ZN(n8608) );
  OR2_X1 U5661 ( .A1(n8605), .A2(n8611), .ZN(n8607) );
  NAND2_X1 U5662 ( .A1(n8636), .A2(n6094), .ZN(n8619) );
  OR2_X2 U5663 ( .A1(n6085), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6105) );
  AND2_X1 U5664 ( .A1(n6111), .A2(n6110), .ZN(n8638) );
  NAND2_X1 U5665 ( .A1(n6052), .A2(n4318), .ZN(n6078) );
  INV_X1 U5666 ( .A(n6290), .ZN(n8065) );
  NAND2_X1 U5667 ( .A1(n6013), .A2(n4708), .ZN(n6053) );
  AND2_X1 U5668 ( .A1(n4710), .A2(n4709), .ZN(n4708) );
  INV_X1 U5669 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4709) );
  NAND2_X1 U5670 ( .A1(n6013), .A2(n4710), .ZN(n6039) );
  NAND2_X1 U5671 ( .A1(n6013), .A2(n6012), .ZN(n6025) );
  INV_X1 U5672 ( .A(n8267), .ZN(n7888) );
  CLKBUF_X1 U5673 ( .A(n7643), .Z(n7644) );
  INV_X1 U5674 ( .A(n7455), .ZN(n7557) );
  NAND2_X1 U5675 ( .A1(n8139), .A2(n8129), .ZN(n8043) );
  AND2_X1 U5676 ( .A1(n8127), .A2(n8134), .ZN(n8125) );
  INV_X1 U5677 ( .A(n4895), .ZN(n4894) );
  OAI21_X1 U5678 ( .B1(n7008), .B2(n4896), .A(n7163), .ZN(n4895) );
  INV_X1 U5679 ( .A(n7008), .ZN(n8049) );
  NAND2_X1 U5680 ( .A1(n7123), .A2(n8093), .ZN(n7111) );
  NAND2_X1 U5681 ( .A1(n6272), .A2(n5879), .ZN(n6929) );
  OAI21_X1 U5682 ( .B1(n6926), .B2(n6928), .A(n10122), .ZN(n5878) );
  OAI211_X1 U5683 ( .C1(n6300), .C2(n8241), .A(n10150), .B(n6856), .ZN(n7648)
         );
  AND2_X1 U5684 ( .A1(n8498), .A2(n8497), .ZN(n8743) );
  INV_X1 U5685 ( .A(n8516), .ZN(n8517) );
  INV_X1 U5686 ( .A(n8215), .ZN(n4701) );
  OR2_X1 U5687 ( .A1(n8206), .A2(n8041), .ZN(n8570) );
  AND2_X1 U5688 ( .A1(n8595), .A2(n8596), .ZN(n8611) );
  INV_X1 U5689 ( .A(n8266), .ZN(n7950) );
  INV_X1 U5690 ( .A(n8160), .ZN(n4866) );
  INV_X1 U5691 ( .A(n10144), .ZN(n10150) );
  NAND2_X1 U5692 ( .A1(n6228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6232) );
  INV_X1 U5693 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6231) );
  XNOR2_X1 U5694 ( .A(n6241), .B(n6242), .ZN(n7392) );
  OR2_X1 U5695 ( .A1(n5888), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5903) );
  INV_X1 U5696 ( .A(n4501), .ZN(n5655) );
  NAND2_X1 U5697 ( .A1(n6690), .A2(n8964), .ZN(n4428) );
  NAND2_X1 U5698 ( .A1(n9143), .A2(n8913), .ZN(n9052) );
  NAND2_X1 U5699 ( .A1(n7050), .A2(n7049), .ZN(n7210) );
  INV_X1 U5700 ( .A(n7049), .ZN(n4467) );
  INV_X1 U5701 ( .A(n7050), .ZN(n4468) );
  NAND2_X1 U5702 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5539) );
  NAND2_X1 U5703 ( .A1(n9119), .A2(n9118), .ZN(n9117) );
  NAND2_X1 U5704 ( .A1(n7322), .A2(n4305), .ZN(n4829) );
  NAND2_X1 U5705 ( .A1(n9153), .A2(n9154), .ZN(n9152) );
  OAI22_X1 U5706 ( .A1(n5509), .A2(n4294), .B1(n6684), .B2(n8922), .ZN(n6689)
         );
  CLKBUF_X1 U5707 ( .A(n9099), .Z(n4479) );
  CLKBUF_X1 U5708 ( .A(n7320), .Z(n7322) );
  AND2_X1 U5709 ( .A1(n9600), .A2(n9376), .ZN(n9438) );
  AOI21_X1 U5710 ( .B1(n4608), .B2(n9389), .A(n9388), .ZN(n9390) );
  AOI21_X1 U5711 ( .B1(n9041), .B2(n5738), .A(n5737), .ZN(n9031) );
  AND2_X1 U5712 ( .A1(n5730), .A2(n5729), .ZN(n9199) );
  OR2_X1 U5713 ( .A1(n9609), .A2(n5725), .ZN(n5730) );
  AND3_X1 U5714 ( .A1(n4392), .A2(n4630), .A3(n5558), .ZN(n7218) );
  NAND2_X1 U5715 ( .A1(n5732), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n4630) );
  OR2_X1 U5716 ( .A1(n6560), .A2(n6559), .ZN(n6631) );
  OR2_X1 U5717 ( .A1(n6640), .A2(n6641), .ZN(n6781) );
  OR2_X1 U5718 ( .A1(n6633), .A2(n6634), .ZN(n6771) );
  INV_X1 U5719 ( .A(n6783), .ZN(n4487) );
  INV_X1 U5720 ( .A(n6784), .ZN(n4488) );
  OR2_X1 U5721 ( .A1(n6995), .A2(n6996), .ZN(n9564) );
  OR2_X1 U5722 ( .A1(n6988), .A2(n6989), .ZN(n9578) );
  AND2_X1 U5723 ( .A1(n10003), .A2(n10002), .ZN(n10005) );
  OR2_X1 U5724 ( .A1(n10056), .A2(n10057), .ZN(n10053) );
  NAND2_X1 U5725 ( .A1(n4455), .A2(n4454), .ZN(n10058) );
  INV_X1 U5726 ( .A(n10062), .ZN(n4454) );
  INV_X1 U5727 ( .A(n10061), .ZN(n4455) );
  AND2_X1 U5728 ( .A1(n6318), .A2(n4386), .ZN(n9601) );
  INV_X1 U5729 ( .A(n4986), .ZN(n4985) );
  OAI21_X1 U5730 ( .B1(n9259), .B2(n4987), .A(n5731), .ZN(n4986) );
  AND2_X1 U5731 ( .A1(n9366), .A2(n9359), .ZN(n9262) );
  NAND2_X1 U5732 ( .A1(n4512), .A2(n9260), .ZN(n4511) );
  NAND2_X1 U5733 ( .A1(n4514), .A2(n4515), .ZN(n4512) );
  AND2_X1 U5734 ( .A1(n4799), .A2(n4798), .ZN(n4797) );
  AND2_X1 U5735 ( .A1(n5686), .A2(n5010), .ZN(n4572) );
  AND2_X1 U5736 ( .A1(n4944), .A2(n5778), .ZN(n4943) );
  NAND2_X1 U5737 ( .A1(n4946), .A2(n4947), .ZN(n4944) );
  NAND2_X1 U5738 ( .A1(n9695), .A2(n4799), .ZN(n9665) );
  OR2_X1 U5739 ( .A1(n5663), .A2(n9148), .ZN(n5670) );
  OAI21_X1 U5740 ( .B1(n9738), .B2(n4522), .A(n4519), .ZN(n9709) );
  INV_X1 U5741 ( .A(n5662), .ZN(n4981) );
  NAND2_X1 U5742 ( .A1(n4983), .A2(n4324), .ZN(n4982) );
  NAND2_X1 U5743 ( .A1(n9789), .A2(n4303), .ZN(n9745) );
  AND2_X1 U5744 ( .A1(n4973), .A2(n4565), .ZN(n4564) );
  INV_X1 U5745 ( .A(n5626), .ZN(n4566) );
  AND2_X1 U5746 ( .A1(n9331), .A2(n9337), .ZN(n9760) );
  NAND2_X1 U5747 ( .A1(n4470), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5629) );
  INV_X1 U5748 ( .A(n5620), .ZN(n4470) );
  AND2_X1 U5749 ( .A1(n5634), .A2(n9776), .ZN(n5635) );
  NAND2_X1 U5750 ( .A1(n9788), .A2(n5626), .ZN(n9777) );
  INV_X1 U5751 ( .A(n5634), .ZN(n9778) );
  NAND2_X1 U5752 ( .A1(n9838), .A2(n9417), .ZN(n9806) );
  AND2_X1 U5753 ( .A1(n4794), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U5754 ( .A1(n7277), .A2(n5585), .ZN(n7436) );
  NAND2_X1 U5755 ( .A1(n5133), .A2(n7339), .ZN(n7198) );
  NAND2_X1 U5756 ( .A1(n7061), .A2(n7199), .ZN(n7062) );
  NAND2_X1 U5757 ( .A1(n6908), .A2(n5766), .ZN(n6907) );
  INV_X1 U5758 ( .A(n9782), .ZN(n9832) );
  AND2_X1 U5759 ( .A1(n4937), .A2(n5761), .ZN(n9282) );
  NAND2_X1 U5760 ( .A1(n7252), .A2(n5760), .ZN(n6795) );
  NAND2_X1 U5761 ( .A1(n7251), .A2(n7256), .ZN(n7255) );
  AND2_X1 U5762 ( .A1(n5449), .A2(n9376), .ZN(n9864) );
  OR2_X1 U5763 ( .A1(n6356), .A2(n9262), .ZN(n6381) );
  NAND2_X1 U5764 ( .A1(n5309), .A2(n5308), .ZN(n9903) );
  NAND2_X1 U5765 ( .A1(n5223), .A2(n5222), .ZN(n9939) );
  XNOR2_X1 U5766 ( .A(n5421), .B(n5420), .ZN(n8809) );
  XNOR2_X1 U5767 ( .A(n5401), .B(n5400), .ZN(n7761) );
  XNOR2_X1 U5768 ( .A(n5381), .B(n5380), .ZN(n7707) );
  NAND2_X1 U5769 ( .A1(n4595), .A2(n5354), .ZN(n5362) );
  NAND2_X1 U5770 ( .A1(n5353), .A2(n5352), .ZN(n4595) );
  OAI21_X2 U5771 ( .B1(n5458), .B2(n5457), .A(n5456), .ZN(n5491) );
  OAI21_X1 U5772 ( .B1(n5291), .B2(n4591), .A(n5290), .ZN(n5304) );
  XNOR2_X1 U5773 ( .A(n5203), .B(n5204), .ZN(n6474) );
  CLKBUF_X1 U5774 ( .A(n5179), .Z(n5171) );
  OR2_X1 U5775 ( .A1(n5108), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5110) );
  AND2_X1 U5776 ( .A1(n4902), .A2(n5070), .ZN(n5051) );
  INV_X1 U5777 ( .A(n4543), .ZN(n4544) );
  NAND2_X1 U5778 ( .A1(n7421), .A2(n7420), .ZN(n7457) );
  AND3_X1 U5779 ( .A1(n6060), .A2(n6059), .A3(n6058), .ZN(n7838) );
  AOI21_X1 U5780 ( .B1(n4846), .B2(n4845), .A(n4843), .ZN(n7836) );
  NOR2_X1 U5781 ( .A1(n4848), .A2(n4410), .ZN(n4845) );
  OAI21_X1 U5782 ( .B1(n4847), .B2(n4410), .A(n4844), .ZN(n4843) );
  INV_X1 U5783 ( .A(n7947), .ZN(n4844) );
  INV_X1 U5784 ( .A(n8572), .ZN(n7850) );
  OAI22_X1 U5785 ( .A1(n6898), .A2(n6897), .B1(n6476), .B2(n6896), .ZN(n6899)
         );
  AND2_X1 U5786 ( .A1(n6123), .A2(n6122), .ZN(n8621) );
  AND4_X1 U5787 ( .A1(n5980), .A2(n5979), .A3(n5978), .A4(n5977), .ZN(n7560)
         );
  OAI21_X1 U5788 ( .B1(n7883), .B2(n4848), .A(n4847), .ZN(n7949) );
  NAND2_X1 U5789 ( .A1(n7079), .A2(n7078), .ZN(n7421) );
  AND2_X1 U5790 ( .A1(n6191), .A2(n6190), .ZN(n8533) );
  NAND2_X1 U5791 ( .A1(n6858), .A2(n6825), .ZN(n8009) );
  NAND2_X1 U5792 ( .A1(n6823), .A2(n6822), .ZN(n8011) );
  XNOR2_X1 U5793 ( .A(n5825), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8255) );
  INV_X1 U5794 ( .A(n8076), .ZN(n8498) );
  NAND2_X1 U5795 ( .A1(n6205), .A2(n6204), .ZN(n8519) );
  INV_X1 U5796 ( .A(n8533), .ZN(n8259) );
  NAND2_X1 U5797 ( .A1(n6151), .A2(n6150), .ZN(n8553) );
  INV_X1 U5798 ( .A(n8591), .ZN(n8574) );
  INV_X1 U5799 ( .A(n8659), .ZN(n8263) );
  AND3_X1 U5800 ( .A1(n6082), .A2(n6081), .A3(n6080), .ZN(n8637) );
  INV_X1 U5801 ( .A(n8657), .ZN(n8264) );
  NAND4_X2 U5802 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n8273)
         );
  OR2_X1 U5803 ( .A1(n5971), .A2(n7117), .ZN(n5899) );
  OAI21_X1 U5804 ( .B1(n8405), .B2(n6584), .A(n6574), .ZN(n6598) );
  INV_X1 U5805 ( .A(n8371), .ZN(n8484) );
  INV_X1 U5806 ( .A(n4448), .ZN(n6880) );
  AND2_X1 U5807 ( .A1(n4647), .A2(n4646), .ZN(n6965) );
  INV_X1 U5808 ( .A(n6883), .ZN(n4646) );
  INV_X1 U5809 ( .A(n4647), .ZN(n6884) );
  INV_X1 U5810 ( .A(n4753), .ZN(n6978) );
  NAND2_X1 U5811 ( .A1(n4724), .A2(n7155), .ZN(n7100) );
  AOI21_X1 U5812 ( .B1(n7145), .B2(n7144), .A(n4662), .ZN(n7309) );
  NAND2_X1 U5813 ( .A1(n4654), .A2(n4657), .ZN(n7359) );
  NAND2_X1 U5814 ( .A1(n7145), .A2(n4658), .ZN(n4654) );
  OAI21_X1 U5815 ( .B1(n7364), .B2(n7363), .A(n7362), .ZN(n8285) );
  INV_X1 U5816 ( .A(n4661), .ZN(n4652) );
  NAND2_X1 U5817 ( .A1(n4657), .A2(n4661), .ZN(n4653) );
  AOI21_X1 U5818 ( .B1(n4659), .B2(n4657), .A(n4656), .ZN(n4655) );
  INV_X1 U5819 ( .A(n4735), .ZN(n4738) );
  NAND2_X1 U5820 ( .A1(n8427), .A2(n8446), .ZN(n8429) );
  AND2_X1 U5821 ( .A1(n8462), .A2(n4763), .ZN(n8439) );
  NAND2_X1 U5822 ( .A1(n4756), .A2(n4310), .ZN(n4763) );
  AND2_X1 U5823 ( .A1(n4733), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4729) );
  INV_X1 U5824 ( .A(n8445), .ZN(n4733) );
  AND2_X1 U5825 ( .A1(n6596), .A2(n8405), .ZN(n8492) );
  XNOR2_X1 U5826 ( .A(n8017), .B(n8227), .ZN(n7752) );
  NAND2_X1 U5827 ( .A1(n6135), .A2(n6134), .ZN(n8703) );
  NAND2_X1 U5828 ( .A1(n6127), .A2(n6126), .ZN(n8706) );
  NAND2_X1 U5829 ( .A1(n6115), .A2(n6114), .ZN(n8711) );
  NAND2_X1 U5830 ( .A1(n6084), .A2(n6083), .ZN(n8726) );
  INV_X1 U5831 ( .A(n10132), .ZN(n4700) );
  NAND2_X1 U5832 ( .A1(n10144), .A2(n6306), .ZN(n8671) );
  INV_X1 U5833 ( .A(n8643), .ZN(n8677) );
  INV_X1 U5834 ( .A(n8666), .ZN(n8630) );
  AND3_X2 U5835 ( .A1(n6267), .A2(n6404), .A3(n6308), .ZN(n10168) );
  INV_X1 U5836 ( .A(n10168), .ZN(n10165) );
  NAND2_X1 U5837 ( .A1(n6396), .A2(n6395), .ZN(n6397) );
  NAND2_X1 U5838 ( .A1(n8572), .A2(n8573), .ZN(n6395) );
  NAND2_X1 U5839 ( .A1(n6174), .A2(n6173), .ZN(n8769) );
  CLKBUF_X1 U5840 ( .A(n8560), .Z(n8561) );
  NAND2_X1 U5841 ( .A1(n6144), .A2(n6143), .ZN(n8775) );
  NAND2_X1 U5842 ( .A1(n6077), .A2(n6076), .ZN(n8800) );
  NAND2_X1 U5843 ( .A1(n8652), .A2(n8171), .ZN(n8661) );
  NAND2_X1 U5844 ( .A1(n6050), .A2(n6049), .ZN(n8002) );
  NAND2_X1 U5845 ( .A1(n6038), .A2(n6037), .ZN(n7839) );
  CLKBUF_X1 U5846 ( .A(n7700), .Z(n7701) );
  NAND2_X1 U5847 ( .A1(n4692), .A2(n8147), .ZN(n7656) );
  NAND2_X1 U5848 ( .A1(n4697), .A2(n4695), .ZN(n4692) );
  AND2_X1 U5849 ( .A1(n7601), .A2(n7600), .ZN(n7610) );
  NAND2_X1 U5850 ( .A1(n4697), .A2(n8143), .ZN(n7603) );
  NAND2_X1 U5851 ( .A1(n4561), .A2(n4560), .ZN(n4559) );
  INV_X1 U5852 ( .A(n6465), .ZN(n4561) );
  AND2_X1 U5853 ( .A1(n6263), .A2(n6262), .ZN(n8808) );
  AND2_X1 U5854 ( .A1(n7392), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6486) );
  INV_X1 U5855 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n5843) );
  INV_X1 U5856 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7669) );
  INV_X1 U5857 ( .A(n6246), .ZN(n7671) );
  INV_X1 U5858 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7638) );
  INV_X1 U5859 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7654) );
  INV_X1 U5860 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7394) );
  INV_X1 U5861 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7290) );
  INV_X1 U5862 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7250) );
  INV_X1 U5863 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7110) );
  NAND2_X1 U5864 ( .A1(n6096), .A2(n5816), .ZN(n6207) );
  INV_X1 U5865 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7006) );
  INV_X1 U5866 ( .A(n6259), .ZN(n8487) );
  NOR2_X1 U5867 ( .A1(n4543), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8820) );
  INV_X1 U5868 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6724) );
  INV_X1 U5869 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6830) );
  INV_X1 U5870 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5871 ( .A1(n5859), .A2(n8811), .ZN(n4790) );
  NAND2_X1 U5872 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4791) );
  INV_X1 U5873 ( .A(n6585), .ZN(n5873) );
  OAI21_X1 U5874 ( .B1(n7322), .B2(n7321), .A(n4832), .ZN(n7581) );
  NAND2_X1 U5875 ( .A1(n9152), .A2(n8867), .ZN(n8987) );
  NOR3_X1 U5876 ( .A1(n9162), .A2(n8998), .A3(n8997), .ZN(n9001) );
  AND2_X1 U5877 ( .A1(n4402), .A2(n8894), .ZN(n4833) );
  OAI21_X1 U5878 ( .B1(n9112), .B2(n4818), .A(n4815), .ZN(n9079) );
  AND4_X1 U5879 ( .A1(n5600), .A2(n5599), .A3(n5598), .A4(n5597), .ZN(n9157)
         );
  AND4_X1 U5880 ( .A1(n5584), .A2(n5583), .A3(n5582), .A4(n5581), .ZN(n9178)
         );
  NAND2_X1 U5881 ( .A1(n4479), .A2(n8894), .ZN(n9185) );
  AND2_X1 U5882 ( .A1(n6683), .A2(n6682), .ZN(n9210) );
  INV_X1 U5883 ( .A(n9215), .ZN(n9205) );
  INV_X1 U5884 ( .A(n9196), .ZN(n9217) );
  AND2_X1 U5885 ( .A1(n5745), .A2(n5744), .ZN(n7022) );
  OR2_X1 U5886 ( .A1(n9622), .A2(n5725), .ZN(n5721) );
  NAND2_X1 U5887 ( .A1(n5711), .A2(n5710), .ZN(n9457) );
  OR2_X1 U5888 ( .A1(n9639), .A2(n5725), .ZN(n5711) );
  INV_X1 U5889 ( .A(n9178), .ZN(n9464) );
  INV_X1 U5890 ( .A(n7218), .ZN(n9467) );
  NAND4_X1 U5891 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n9469)
         );
  NAND4_X1 U5892 ( .A1(n5517), .A2(n5516), .A3(n5515), .A4(n5514), .ZN(n9472)
         );
  NAND2_X1 U5893 ( .A1(n5511), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5517) );
  CLKBUF_X1 U5894 ( .A(n5502), .Z(n6715) );
  NAND2_X1 U5895 ( .A1(n5511), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5506) );
  OR2_X1 U5896 ( .A1(n6545), .A2(n6546), .ZN(n6638) );
  OR2_X1 U5897 ( .A1(n6775), .A2(n6776), .ZN(n6986) );
  AND2_X1 U5898 ( .A1(n5215), .A2(n5229), .ZN(n6788) );
  AND2_X1 U5899 ( .A1(n10001), .A2(n10000), .ZN(n10009) );
  AOI211_X1 U5900 ( .C1(n9603), .C2(n9602), .A(n9832), .B(n9601), .ZN(n9865)
         );
  AND2_X1 U5901 ( .A1(n4954), .A2(n9361), .ZN(n6321) );
  XNOR2_X1 U5902 ( .A(n9619), .B(n9260), .ZN(n9873) );
  NAND2_X1 U5903 ( .A1(n4948), .A2(n9257), .ZN(n9659) );
  NAND2_X1 U5904 ( .A1(n4573), .A2(n5686), .ZN(n9663) );
  NAND2_X1 U5905 ( .A1(n9728), .A2(n9729), .ZN(n9727) );
  NAND2_X1 U5906 ( .A1(n9738), .A2(n9338), .ZN(n9728) );
  NAND2_X1 U5907 ( .A1(n5273), .A2(n5272), .ZN(n9919) );
  OAI21_X1 U5908 ( .B1(n9838), .B2(n9804), .A(n4940), .ZN(n9795) );
  OAI21_X1 U5909 ( .B1(n7493), .B2(n4970), .A(n4968), .ZN(n9826) );
  NAND2_X1 U5910 ( .A1(n7494), .A2(n5601), .ZN(n9828) );
  NAND2_X1 U5911 ( .A1(n5772), .A2(n9318), .ZN(n7497) );
  NAND2_X1 U5912 ( .A1(n4952), .A2(n9410), .ZN(n7280) );
  OAI21_X1 U5913 ( .B1(n7228), .B2(n4965), .A(n4963), .ZN(n7377) );
  NAND2_X1 U5914 ( .A1(n7229), .A2(n5569), .ZN(n7376) );
  OR2_X1 U5915 ( .A1(n5796), .A2(n5795), .ZN(n9783) );
  NAND2_X1 U5916 ( .A1(n5423), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4809) );
  AND2_X1 U5917 ( .A1(n9855), .A2(n6699), .ZN(n10074) );
  AND2_X1 U5918 ( .A1(n9855), .A2(n5758), .ZN(n10071) );
  INV_X1 U5919 ( .A(n10074), .ZN(n9836) );
  AND2_X1 U5920 ( .A1(n7286), .A2(n6686), .ZN(n10089) );
  OR2_X1 U5921 ( .A1(n5796), .A2(n6672), .ZN(n5752) );
  NAND2_X1 U5922 ( .A1(n4631), .A2(n5146), .ZN(n7221) );
  NAND2_X1 U5923 ( .A1(n6441), .A2(n5422), .ZN(n4631) );
  AND2_X1 U5924 ( .A1(n5241), .A2(n4387), .ZN(n4568) );
  INV_X1 U5925 ( .A(n9637), .ZN(n9955) );
  INV_X1 U5926 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7672) );
  INV_X1 U5927 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7639) );
  INV_X1 U5928 ( .A(n5472), .ZN(n7641) );
  INV_X1 U5929 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10231) );
  INV_X1 U5930 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7287) );
  INV_X1 U5931 ( .A(n4301), .ZN(n7286) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7248) );
  NAND2_X1 U5933 ( .A1(n4433), .A2(n4432), .ZN(n5436) );
  NAND2_X1 U5934 ( .A1(n5435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4432) );
  INV_X1 U5935 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7108) );
  AND2_X1 U5936 ( .A1(n5284), .A2(n5283), .ZN(n10065) );
  INV_X1 U5937 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6726) );
  INV_X1 U5938 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6832) );
  AND2_X1 U5939 ( .A1(n5238), .A2(n5232), .ZN(n10006) );
  AND2_X1 U5940 ( .A1(n5157), .A2(n5173), .ZN(n9540) );
  CLKBUF_X2 U5941 ( .A(P1_IR_REG_0__SCAN_IN), .Z(n4469) );
  NOR2_X1 U5942 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  NOR2_X1 U5943 ( .A1(n7834), .A2(n8015), .ZN(n4463) );
  NAND2_X1 U5944 ( .A1(n4666), .A2(n8475), .ZN(n4665) );
  OAI21_X1 U5945 ( .B1(n4320), .B2(n8457), .A(n8488), .ZN(n4666) );
  NAND2_X1 U5946 ( .A1(n4478), .A2(n4477), .ZN(P2_U3205) );
  NAND2_X1 U5947 ( .A1(n8510), .A2(n8663), .ZN(n4477) );
  INV_X1 U5948 ( .A(n8509), .ZN(n4478) );
  NAND2_X1 U5949 ( .A1(n8528), .A2(n4441), .ZN(P2_U3206) );
  INV_X1 U5950 ( .A(n4442), .ZN(n4441) );
  OAI21_X1 U5951 ( .B1(n8754), .B2(n8669), .A(n8527), .ZN(n4442) );
  OR2_X1 U5952 ( .A1(n8508), .A2(n8716), .ZN(n6301) );
  NAND2_X1 U5953 ( .A1(n8689), .A2(n4443), .ZN(P2_U3486) );
  INV_X1 U5954 ( .A(n4444), .ZN(n4443) );
  OAI21_X1 U5955 ( .B1(n8754), .B2(n8716), .A(n8688), .ZN(n4444) );
  NOR2_X1 U5956 ( .A1(n6353), .A2(n4994), .ZN(n6354) );
  NAND2_X1 U5957 ( .A1(n8753), .A2(n4439), .ZN(P2_U3454) );
  INV_X1 U5958 ( .A(n4440), .ZN(n4439) );
  OAI21_X1 U5959 ( .B1(n8754), .B2(n8790), .A(n8752), .ZN(n4440) );
  NAND2_X1 U5960 ( .A1(n9048), .A2(n9049), .ZN(n4426) );
  NAND2_X1 U5961 ( .A1(n4453), .A2(n4451), .ZN(P1_U3229) );
  NOR2_X1 U5962 ( .A1(n9116), .A2(n4452), .ZN(n4451) );
  AND2_X1 U5963 ( .A1(n9652), .A2(n9215), .ZN(n4452) );
  OR2_X1 U5964 ( .A1(n9451), .A2(n9450), .ZN(n4579) );
  NAND2_X1 U5965 ( .A1(n4491), .A2(n4489), .ZN(P1_U3262) );
  AOI21_X1 U5966 ( .B1(n9592), .B2(n9765), .A(n4490), .ZN(n4489) );
  AOI21_X1 U5967 ( .B1(n9391), .B2(n9899), .A(n5494), .ZN(n5495) );
  NAND2_X1 U5968 ( .A1(n5746), .A2(n9899), .ZN(n6387) );
  OAI21_X1 U5969 ( .B1(n4808), .B2(n6370), .A(n6369), .ZN(n6371) );
  AOI21_X1 U5970 ( .B1(n9949), .B2(n10117), .A(n4574), .ZN(n9874) );
  NAND2_X1 U5971 ( .A1(n4576), .A2(n4575), .ZN(n4574) );
  NAND2_X1 U5972 ( .A1(n10118), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n4575) );
  NOR2_X1 U5973 ( .A1(n6415), .A2(n6414), .ZN(n6416) );
  AOI21_X1 U5974 ( .B1(n9949), .B2(n10348), .A(n4525), .ZN(n9951) );
  NAND2_X1 U5975 ( .A1(n4527), .A2(n4526), .ZN(n4525) );
  NAND2_X1 U5976 ( .A1(n10346), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n4526) );
  AND3_X1 U5977 ( .A1(n4537), .A2(n4393), .A3(n4316), .ZN(n4302) );
  AND2_X1 U5978 ( .A1(n4308), .A2(n4803), .ZN(n4303) );
  BUF_X1 U5979 ( .A(n5960), .Z(n5986) );
  INV_X2 U5980 ( .A(n5960), .ZN(n6057) );
  NAND2_X1 U5981 ( .A1(n5254), .A2(n5013), .ZN(n4304) );
  AND2_X1 U5982 ( .A1(n4353), .A2(n4832), .ZN(n4305) );
  INV_X1 U5983 ( .A(n7339), .ZN(n7317) );
  AND2_X1 U5984 ( .A1(n5132), .A2(n5131), .ZN(n7339) );
  INV_X1 U5985 ( .A(n9804), .ZN(n9807) );
  INV_X1 U5986 ( .A(n5207), .ZN(n5206) );
  INV_X1 U5987 ( .A(n9338), .ZN(n4521) );
  AND2_X1 U5988 ( .A1(n7298), .A2(n7357), .ZN(n4306) );
  INV_X1 U5989 ( .A(n9417), .ZN(n4942) );
  AND2_X1 U5990 ( .A1(n7424), .A2(n7423), .ZN(n4307) );
  AND2_X1 U5991 ( .A1(n9307), .A2(n9108), .ZN(n4308) );
  AND4_X1 U5992 ( .A1(n8068), .A2(n4720), .A3(n4718), .A4(n4334), .ZN(n4309)
         );
  OR2_X1 U5993 ( .A1(n8418), .A2(n8417), .ZN(n4310) );
  AND2_X1 U5994 ( .A1(n8172), .A2(n8235), .ZN(n4311) );
  AND2_X1 U5995 ( .A1(n9335), .A2(n9384), .ZN(n4312) );
  AND2_X1 U5996 ( .A1(n7777), .A2(n8268), .ZN(n4313) );
  INV_X1 U5997 ( .A(n8416), .ZN(n4769) );
  OR2_X1 U5998 ( .A1(n4648), .A2(n6768), .ZN(n4314) );
  OR2_X1 U5999 ( .A1(n9637), .A2(n9198), .ZN(n9362) );
  INV_X1 U6000 ( .A(n9362), .ZN(n4628) );
  AOI21_X1 U6001 ( .B1(n4658), .B2(n4662), .A(n4375), .ZN(n4657) );
  INV_X1 U6002 ( .A(n8872), .ZN(n4822) );
  AND2_X1 U6003 ( .A1(n7156), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4315) );
  OR2_X1 U6004 ( .A1(n8221), .A2(n4531), .ZN(n4316) );
  AND2_X1 U6005 ( .A1(n4303), .A2(n4802), .ZN(n4317) );
  AOI21_X1 U6006 ( .B1(n8418), .B2(n8416), .A(n8417), .ZN(n4766) );
  AND2_X1 U6007 ( .A1(n6051), .A2(n4713), .ZN(n4318) );
  AND2_X1 U6008 ( .A1(n7361), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4319) );
  NAND2_X1 U6009 ( .A1(n4751), .A2(n6966), .ZN(n4753) );
  OR2_X1 U6010 ( .A1(n5616), .A2(n9211), .ZN(n9304) );
  OR2_X1 U6011 ( .A1(n8476), .A2(n8456), .ZN(n4320) );
  NAND2_X1 U6012 ( .A1(n7597), .A2(n6006), .ZN(n7595) );
  NAND2_X1 U6013 ( .A1(n4982), .A2(n4980), .ZN(n9675) );
  INV_X1 U6014 ( .A(n7813), .ZN(n7772) );
  NAND2_X1 U6015 ( .A1(n9789), .A2(n4308), .ZN(n9744) );
  NAND2_X1 U6016 ( .A1(n4829), .A2(n4830), .ZN(n8844) );
  AND2_X1 U6017 ( .A1(n9723), .A2(n9717), .ZN(n9695) );
  INV_X1 U6018 ( .A(n5512), .ZN(n5546) );
  NAND2_X1 U6019 ( .A1(n4430), .A2(n5024), .ZN(n4321) );
  OR2_X1 U6020 ( .A1(n9667), .A2(n9220), .ZN(n4322) );
  NAND2_X1 U6021 ( .A1(n9789), .A2(n9307), .ZN(n4323) );
  NAND2_X1 U6022 ( .A1(n9777), .A2(n5635), .ZN(n9775) );
  INV_X1 U6023 ( .A(n9472), .ZN(n5518) );
  NAND2_X1 U6024 ( .A1(n9908), .A2(n9462), .ZN(n4324) );
  AND2_X1 U6025 ( .A1(n6849), .A2(n8039), .ZN(n4325) );
  NOR2_X1 U6026 ( .A1(n7844), .A2(n8553), .ZN(n4326) );
  AND2_X1 U6027 ( .A1(n9602), .A2(n9383), .ZN(n4327) );
  NAND2_X1 U6028 ( .A1(n5067), .A2(n6430), .ZN(n5210) );
  AND2_X1 U6029 ( .A1(n9701), .A2(n9700), .ZN(n9713) );
  AND3_X1 U6030 ( .A1(n5917), .A2(n5916), .A3(n5915), .ZN(n4328) );
  AND3_X1 U6031 ( .A1(n5929), .A2(n5928), .A3(n5927), .ZN(n4329) );
  NAND2_X1 U6032 ( .A1(n4927), .A2(n4929), .ZN(n5208) );
  NAND2_X1 U6033 ( .A1(n9402), .A2(n9279), .ZN(n6950) );
  OR2_X1 U6034 ( .A1(n8229), .A2(n8228), .ZN(n4330) );
  NAND2_X1 U6035 ( .A1(n8607), .A2(n6124), .ZN(n8589) );
  NAND2_X1 U6036 ( .A1(n4972), .A2(n5695), .ZN(n9645) );
  NAND2_X1 U6037 ( .A1(n9775), .A2(n5636), .ZN(n9754) );
  NAND2_X1 U6038 ( .A1(n4703), .A2(n8198), .ZN(n8568) );
  INV_X1 U6039 ( .A(n9240), .ZN(n5773) );
  INV_X1 U6040 ( .A(n9428), .ZN(n4520) );
  NOR2_X1 U6041 ( .A1(n9950), .A2(n9456), .ZN(n4331) );
  INV_X1 U6042 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5842) );
  AND2_X1 U6043 ( .A1(n8381), .A2(n8408), .ZN(n4332) );
  OR2_X1 U6044 ( .A1(n5858), .A2(n6659), .ZN(n4333) );
  NAND2_X1 U6045 ( .A1(n5315), .A2(n5314), .ZN(n9968) );
  NAND2_X1 U6046 ( .A1(n5774), .A2(n9331), .ZN(n9737) );
  NAND2_X1 U6047 ( .A1(n5414), .A2(n5413), .ZN(n9602) );
  INV_X1 U6048 ( .A(n9602), .ZN(n4804) );
  NOR4_X1 U6049 ( .A1(n8570), .A2(n8066), .A3(n8200), .A4(n8590), .ZN(n4334)
         );
  NOR3_X1 U6050 ( .A1(n9265), .A2(n9438), .A3(n9440), .ZN(n4335) );
  NAND2_X1 U6051 ( .A1(n4873), .A2(n4874), .ZN(n8633) );
  OR2_X1 U6052 ( .A1(n5858), .A2(n6762), .ZN(n4336) );
  AND2_X1 U6053 ( .A1(n8505), .A2(n8078), .ZN(n4337) );
  AND2_X1 U6054 ( .A1(n8171), .A2(n6290), .ZN(n4338) );
  AND2_X1 U6055 ( .A1(n9304), .A2(n9382), .ZN(n4339) );
  AND2_X1 U6056 ( .A1(n5891), .A2(n4336), .ZN(n4340) );
  OR2_X1 U6057 ( .A1(n9652), .A2(n9458), .ZN(n4341) );
  AND2_X1 U6058 ( .A1(n9758), .A2(n9760), .ZN(n4342) );
  NAND2_X1 U6059 ( .A1(n4705), .A2(n8042), .ZN(n8648) );
  OR2_X1 U6060 ( .A1(n7092), .A2(n7098), .ZN(n4343) );
  NAND2_X1 U6061 ( .A1(n4982), .A2(n5662), .ZN(n9712) );
  NOR2_X1 U6062 ( .A1(n8993), .A2(n9164), .ZN(n4344) );
  OR2_X1 U6063 ( .A1(n9680), .A2(n4613), .ZN(n4345) );
  INV_X1 U6064 ( .A(n9360), .ZN(n4629) );
  NAND2_X1 U6065 ( .A1(n5200), .A2(n5199), .ZN(n8845) );
  INV_X1 U6066 ( .A(n9361), .ZN(n4955) );
  AND2_X1 U6067 ( .A1(n9432), .A2(n4518), .ZN(n4346) );
  NAND2_X1 U6068 ( .A1(n8177), .A2(n8235), .ZN(n4347) );
  AND2_X1 U6069 ( .A1(n9306), .A2(n4339), .ZN(n4348) );
  OR2_X1 U6070 ( .A1(n8250), .A2(n8249), .ZN(n4349) );
  NOR2_X1 U6071 ( .A1(n7556), .A2(n7557), .ZN(n4350) );
  NAND2_X1 U6072 ( .A1(n5399), .A2(n5398), .ZN(n5746) );
  AND2_X1 U6073 ( .A1(n5775), .A2(n9331), .ZN(n4351) );
  AND2_X1 U6074 ( .A1(n8173), .A2(n8079), .ZN(n8634) );
  INV_X1 U6075 ( .A(n8200), .ZN(n4541) );
  AND2_X1 U6076 ( .A1(n9796), .A2(n4938), .ZN(n4352) );
  OR2_X1 U6077 ( .A1(n7578), .A2(n7577), .ZN(n4353) );
  INV_X1 U6078 ( .A(n4922), .ZN(n4921) );
  OAI21_X1 U6079 ( .B1(n5206), .B2(n4923), .A(n5225), .ZN(n4922) );
  NAND2_X1 U6080 ( .A1(n7968), .A2(n7766), .ZN(n4354) );
  INV_X1 U6081 ( .A(n9414), .ZN(n4642) );
  OR2_X1 U6082 ( .A1(n8159), .A2(n8162), .ZN(n4355) );
  INV_X1 U6083 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8811) );
  NAND4_X1 U6084 ( .A1(n8204), .A2(n8203), .A3(n8222), .A4(n8562), .ZN(n4356)
         );
  AND2_X1 U6085 ( .A1(n8800), .A2(n7783), .ZN(n4357) );
  OR2_X1 U6086 ( .A1(n5245), .A2(SI_15_), .ZN(n4358) );
  NOR2_X1 U6087 ( .A1(n9747), .A2(n9730), .ZN(n4359) );
  NOR2_X1 U6088 ( .A1(n8830), .A2(n9465), .ZN(n4360) );
  NOR2_X1 U6089 ( .A1(n8706), .A2(n8260), .ZN(n4361) );
  NOR2_X1 U6090 ( .A1(n9939), .A2(n9075), .ZN(n4362) );
  INV_X1 U6091 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5586) );
  INV_X1 U6092 ( .A(n8214), .ZN(n4540) );
  INV_X1 U6093 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5439) );
  OR2_X1 U6094 ( .A1(n9950), .A2(n9219), .ZN(n4363) );
  AND2_X1 U6095 ( .A1(n9366), .A2(n9358), .ZN(n4364) );
  AND2_X1 U6096 ( .A1(n4505), .A2(n9432), .ZN(n4365) );
  OR2_X1 U6097 ( .A1(n7790), .A2(n7789), .ZN(n4366) );
  INV_X1 U6098 ( .A(n4659), .ZN(n4658) );
  OAI21_X1 U6099 ( .B1(n7144), .B2(n4662), .A(n4660), .ZN(n4659) );
  INV_X1 U6100 ( .A(n4322), .ZN(n4613) );
  OR2_X1 U6101 ( .A1(n8142), .A2(n4674), .ZN(n4367) );
  INV_X1 U6102 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5822) );
  AND2_X1 U6103 ( .A1(n4820), .A2(n8873), .ZN(n4368) );
  INV_X1 U6104 ( .A(n9391), .ZN(n9600) );
  NAND2_X1 U6105 ( .A1(n5425), .A2(n5424), .ZN(n9391) );
  AND2_X1 U6106 ( .A1(n4557), .A2(n4355), .ZN(n4369) );
  NAND2_X1 U6107 ( .A1(n9677), .A2(n9676), .ZN(n4370) );
  INV_X1 U6108 ( .A(n9635), .ZN(n4515) );
  AND2_X1 U6109 ( .A1(n9362), .A2(n9226), .ZN(n9635) );
  AND2_X1 U6110 ( .A1(n4689), .A2(n4337), .ZN(n4371) );
  OR2_X1 U6111 ( .A1(n8467), .A2(n8448), .ZN(n4372) );
  NAND2_X1 U6112 ( .A1(n8594), .A2(n8173), .ZN(n4373) );
  INV_X1 U6113 ( .A(n8867), .ZN(n4821) );
  NAND2_X1 U6114 ( .A1(n6318), .A2(n4805), .ZN(n4374) );
  NOR2_X1 U6115 ( .A1(n7307), .A2(n7306), .ZN(n4375) );
  AND2_X1 U6116 ( .A1(n4540), .A2(n8200), .ZN(n4376) );
  AND2_X1 U6117 ( .A1(n8843), .A2(n4305), .ZN(n4377) );
  INV_X1 U6118 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U6119 ( .A1(n9695), .A2(n4801), .ZN(n4378) );
  OR2_X1 U6120 ( .A1(n8212), .A2(n8211), .ZN(n4379) );
  NAND2_X1 U6121 ( .A1(n9378), .A2(n9377), .ZN(n9370) );
  INV_X1 U6122 ( .A(n9370), .ZN(n4502) );
  AND3_X1 U6123 ( .A1(n9288), .A2(n9287), .A3(n9286), .ZN(n4380) );
  OR2_X1 U6124 ( .A1(n9349), .A2(n9382), .ZN(n4381) );
  OR2_X1 U6125 ( .A1(n6763), .A2(n6762), .ZN(n4382) );
  OR2_X1 U6126 ( .A1(n8131), .A2(n8126), .ZN(n4383) );
  AND2_X1 U6127 ( .A1(n9919), .A2(n9772), .ZN(n4384) );
  AND2_X1 U6128 ( .A1(n4698), .A2(n8147), .ZN(n4385) );
  AND2_X1 U6129 ( .A1(n4806), .A2(n4804), .ZN(n4386) );
  NOR2_X1 U6130 ( .A1(n9713), .A2(n4981), .ZN(n4980) );
  AND2_X1 U6131 ( .A1(n5149), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4387) );
  NAND2_X1 U6132 ( .A1(n4700), .A2(n6894), .ZN(n8093) );
  AND2_X1 U6133 ( .A1(n9260), .A2(n9362), .ZN(n4388) );
  AND2_X1 U6134 ( .A1(n5012), .A2(n5950), .ZN(n4389) );
  INV_X1 U6135 ( .A(n7166), .ZN(n4896) );
  AND2_X1 U6136 ( .A1(n5842), .A2(n4680), .ZN(n4390) );
  OR2_X1 U6137 ( .A1(n8029), .A2(n5039), .ZN(n4391) );
  AND2_X1 U6138 ( .A1(n5559), .A2(n5560), .ZN(n4392) );
  INV_X1 U6139 ( .A(n4880), .ZN(n4879) );
  NAND2_X1 U6140 ( .A1(n8590), .A2(n4881), .ZN(n4880) );
  OR2_X1 U6141 ( .A1(n8221), .A2(n4530), .ZN(n4393) );
  OR2_X1 U6142 ( .A1(n4750), .A2(n4754), .ZN(n4394) );
  OR2_X1 U6143 ( .A1(n8218), .A2(n8219), .ZN(n8540) );
  INV_X1 U6144 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5032) );
  INV_X1 U6145 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n4435) );
  INV_X1 U6146 ( .A(n5890), .ZN(n5907) );
  INV_X1 U6147 ( .A(n6007), .ZN(n4560) );
  NAND2_X1 U6148 ( .A1(n6842), .A2(n8643), .ZN(n8663) );
  NAND2_X1 U6149 ( .A1(n5383), .A2(n5382), .ZN(n9045) );
  INV_X1 U6150 ( .A(n9045), .ZN(n4808) );
  NAND2_X1 U6151 ( .A1(n7408), .A2(n4698), .ZN(n4697) );
  NAND2_X1 U6152 ( .A1(n5351), .A2(n5350), .ZN(n9652) );
  INV_X1 U6153 ( .A(n9652), .ZN(n4798) );
  AND2_X1 U6154 ( .A1(n8343), .A2(n8358), .ZN(n4395) );
  NAND2_X1 U6155 ( .A1(n6809), .A2(n6808), .ZN(n8003) );
  NAND2_X1 U6156 ( .A1(n4437), .A2(n8103), .ZN(n7007) );
  NOR2_X1 U6157 ( .A1(n4784), .A2(n4783), .ZN(n4396) );
  NAND2_X1 U6158 ( .A1(n4897), .A2(n7008), .ZN(n7010) );
  NOR2_X1 U6159 ( .A1(n8487), .A2(n8242), .ZN(n4397) );
  AND2_X1 U6160 ( .A1(n7379), .A2(n4796), .ZN(n4398) );
  INV_X2 U6161 ( .A(n10156), .ZN(n10155) );
  INV_X1 U6162 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n4776) );
  NAND2_X1 U6163 ( .A1(n4898), .A2(n5950), .ZN(n7273) );
  INV_X1 U6164 ( .A(n9110), .ZN(n4818) );
  NAND2_X1 U6165 ( .A1(n5906), .A2(n5920), .ZN(n6881) );
  NAND2_X1 U6166 ( .A1(n7062), .A2(n5551), .ZN(n7196) );
  AND3_X1 U6167 ( .A1(n5402), .A2(n5393), .A3(n5403), .ZN(n4399) );
  AND2_X1 U6168 ( .A1(n9339), .A2(n9331), .ZN(n4400) );
  AND2_X1 U6169 ( .A1(n9322), .A2(n9318), .ZN(n4401) );
  NAND2_X1 U6170 ( .A1(n4773), .A2(n8298), .ZN(n8320) );
  INV_X1 U6171 ( .A(n7143), .ZN(n7098) );
  OR2_X1 U6172 ( .A1(n8901), .A2(n8900), .ZN(n4402) );
  AND2_X1 U6173 ( .A1(n4738), .A2(n4740), .ZN(n4403) );
  INV_X1 U6174 ( .A(n8981), .ZN(n9870) );
  NAND2_X1 U6175 ( .A1(n5379), .A2(n5378), .ZN(n8981) );
  INV_X1 U6176 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5609) );
  INV_X1 U6177 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5602) );
  INV_X1 U6178 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6012) );
  OR2_X1 U6179 ( .A1(n7991), .A2(n7992), .ZN(n4404) );
  AND2_X1 U6180 ( .A1(n8334), .A2(n8355), .ZN(n4405) );
  OR2_X1 U6181 ( .A1(n9961), .A2(n9205), .ZN(n4406) );
  AND2_X1 U6182 ( .A1(n4715), .A2(n4714), .ZN(n4407) );
  AND2_X1 U6183 ( .A1(n4771), .A2(n8320), .ZN(n4408) );
  NOR2_X2 U6184 ( .A1(n6518), .A2(n6517), .ZN(n4409) );
  AND2_X1 U6185 ( .A1(n6871), .A2(n6887), .ZN(n4755) );
  NAND2_X1 U6186 ( .A1(n5286), .A2(n5285), .ZN(n9747) );
  INV_X1 U6187 ( .A(n9747), .ZN(n4803) );
  INV_X1 U6188 ( .A(n8856), .ZN(n4793) );
  AND2_X1 U6189 ( .A1(n8039), .A2(n6211), .ZN(n8653) );
  INV_X1 U6190 ( .A(n8653), .ZN(n8640) );
  AND2_X2 U6191 ( .A1(n5804), .A2(n6672), .ZN(n10117) );
  NAND2_X1 U6192 ( .A1(n5303), .A2(n5302), .ZN(n9908) );
  INV_X1 U6193 ( .A(n9908), .ZN(n4802) );
  AND2_X1 U6194 ( .A1(n7778), .A2(n7888), .ZN(n4410) );
  NAND2_X1 U6195 ( .A1(n6905), .A2(n5545), .ZN(n7061) );
  NAND2_X1 U6196 ( .A1(n4777), .A2(n7300), .ZN(n7368) );
  INV_X1 U6197 ( .A(n7368), .ZN(n4783) );
  AND2_X1 U6198 ( .A1(n8451), .A2(n8417), .ZN(n4411) );
  INV_X1 U6199 ( .A(n8417), .ZN(n4768) );
  NAND2_X1 U6200 ( .A1(n4723), .A2(n4722), .ZN(n4412) );
  INV_X1 U6201 ( .A(n7123), .ZN(n8048) );
  NAND2_X1 U6202 ( .A1(n8102), .A2(n8093), .ZN(n7123) );
  AND2_X1 U6203 ( .A1(n6971), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4413) );
  AND2_X1 U6204 ( .A1(n8438), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n4414) );
  AND2_X1 U6205 ( .A1(n4752), .A2(n4753), .ZN(n4415) );
  AND2_X1 U6206 ( .A1(n5001), .A2(n6971), .ZN(n4416) );
  XOR2_X1 U6207 ( .A(n7095), .B(P2_REG1_REG_6__SCAN_IN), .Z(n4417) );
  XOR2_X1 U6208 ( .A(n8378), .B(P2_REG1_REG_14__SCAN_IN), .Z(n4418) );
  XOR2_X1 U6209 ( .A(n8424), .B(P2_REG2_REG_16__SCAN_IN), .Z(n4419) );
  BUF_X1 U6210 ( .A(n5485), .Z(n9765) );
  AND2_X1 U6211 ( .A1(n8487), .A2(n8242), .ZN(n8241) );
  INV_X1 U6212 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4754) );
  INV_X1 U6213 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n4728) );
  INV_X1 U6214 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n4758) );
  INV_X1 U6215 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n4789) );
  INV_X1 U6216 ( .A(n8451), .ZN(n4765) );
  XNOR2_X1 U6217 ( .A(n6075), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8451) );
  NAND2_X1 U6218 ( .A1(n4438), .A2(n5810), .ZN(n5951) );
  NAND2_X1 U6219 ( .A1(n7559), .A2(n7558), .ZN(n7687) );
  NAND2_X1 U6220 ( .A1(n7807), .A2(n7806), .ZN(n7927) );
  NAND2_X1 U6221 ( .A1(n6940), .A2(n6941), .ZN(n7024) );
  XNOR2_X2 U6222 ( .A(n6099), .B(P2_IR_REG_19__SCAN_IN), .ZN(n6259) );
  NAND2_X1 U6223 ( .A1(n7873), .A2(n7802), .ZN(n7959) );
  NAND2_X2 U6224 ( .A1(n6848), .A2(n4325), .ZN(n6854) );
  OAI21_X2 U6225 ( .B1(n9026), .B2(n9024), .A(n9022), .ZN(n9144) );
  OAI21_X1 U6226 ( .B1(n9392), .B2(n9391), .A(n9390), .ZN(n9398) );
  NOR4_X1 U6227 ( .A1(n9329), .A2(n9328), .A3(n9382), .A4(n9422), .ZN(n9330)
         );
  NAND2_X1 U6228 ( .A1(n5030), .A2(n4424), .ZN(n5442) );
  NAND2_X1 U6229 ( .A1(n4913), .A2(n4912), .ZN(n9333) );
  NAND2_X1 U6230 ( .A1(n9336), .A2(n4610), .ZN(n4609) );
  NAND2_X1 U6231 ( .A1(n4911), .A2(n4420), .ZN(n9341) );
  NAND2_X1 U6232 ( .A1(n9144), .A2(n9145), .ZN(n9143) );
  OAI21_X1 U6233 ( .B1(n9065), .B2(n9067), .A(n9066), .ZN(n9064) );
  INV_X4 U6234 ( .A(n5149), .ZN(n6430) );
  NAND2_X1 U6235 ( .A1(n6690), .A2(n6494), .ZN(n6692) );
  AND2_X1 U6236 ( .A1(n6492), .A2(n6493), .ZN(n6690) );
  AOI21_X1 U6237 ( .B1(n7320), .B2(n4377), .A(n4825), .ZN(n9065) );
  NOR2_X1 U6238 ( .A1(n4427), .A2(n4426), .ZN(n4425) );
  INV_X1 U6239 ( .A(n5503), .ZN(n6684) );
  OAI211_X1 U6240 ( .C1(n9282), .C2(n9281), .A(n9280), .B(n9279), .ZN(n9283)
         );
  NOR2_X1 U6241 ( .A1(n9040), .A2(n4810), .ZN(n4427) );
  NAND2_X1 U6242 ( .A1(n6692), .A2(n6691), .ZN(n4429) );
  NAND2_X1 U6243 ( .A1(n9093), .A2(n8887), .ZN(n9100) );
  NAND2_X1 U6244 ( .A1(n9050), .A2(n4425), .ZN(P1_U3220) );
  AND2_X2 U6245 ( .A1(n6693), .A2(n6694), .ZN(n6714) );
  AND2_X1 U6246 ( .A1(n4429), .A2(n4428), .ZN(n6693) );
  INV_X1 U6247 ( .A(n4430), .ZN(n5460) );
  NAND2_X1 U6248 ( .A1(n4434), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4433) );
  OR2_X1 U6249 ( .A1(n5434), .A2(n5035), .ZN(n4434) );
  INV_X1 U6250 ( .A(n9115), .ZN(n4453) );
  AND2_X2 U6251 ( .A1(n9195), .A2(n8975), .ZN(n9040) );
  NAND2_X1 U6252 ( .A1(n7112), .A2(n6275), .ZN(n4437) );
  NAND2_X2 U6253 ( .A1(n4705), .A2(n4704), .ZN(n8647) );
  NAND2_X2 U6254 ( .A1(n6928), .A2(n7138), .ZN(n8088) );
  NOR2_X1 U6255 ( .A1(n4683), .A2(n4682), .ZN(n4681) );
  OAI22_X1 U6256 ( .A1(n4931), .A2(n5185), .B1(n5202), .B2(SI_11_), .ZN(n4930)
         );
  NAND2_X1 U6257 ( .A1(n4539), .A2(n8540), .ZN(n4538) );
  NAND2_X1 U6258 ( .A1(n4601), .A2(n4599), .ZN(n5276) );
  OAI211_X1 U6259 ( .C1(n8232), .C2(n8519), .A(n4330), .B(n4678), .ZN(n4677)
         );
  NAND2_X1 U6260 ( .A1(n4677), .A2(n8240), .ZN(n4552) );
  NAND2_X2 U6261 ( .A1(n6234), .A2(n6233), .ZN(n6243) );
  NOR2_X1 U6262 ( .A1(n6899), .A2(n6900), .ZN(n6938) );
  NAND2_X2 U6263 ( .A1(n7733), .A2(n6061), .ZN(n7718) );
  INV_X1 U6264 ( .A(n5208), .ZN(n4445) );
  NAND2_X1 U6265 ( .A1(n7007), .A2(n6276), .ZN(n6283) );
  NAND2_X1 U6266 ( .A1(n4447), .A2(n4665), .ZN(P2_U3200) );
  NOR2_X2 U6267 ( .A1(n6647), .A2(n4649), .ZN(n6650) );
  NOR2_X1 U6268 ( .A1(n6597), .A2(n6575), .ZN(n6608) );
  AND2_X4 U6269 ( .A1(n4449), .A2(n4438), .ZN(n5834) );
  NOR2_X2 U6270 ( .A1(n5818), .A2(n5811), .ZN(n4449) );
  NOR2_X1 U6271 ( .A1(n8455), .A2(n8454), .ZN(n8476) );
  NAND2_X1 U6272 ( .A1(n6761), .A2(n4382), .ZN(n6764) );
  OAI21_X1 U6273 ( .B1(n8483), .B2(n8482), .A(n8490), .ZN(n8491) );
  NOR2_X1 U6274 ( .A1(n6608), .A2(n5004), .ZN(n6610) );
  NAND2_X1 U6275 ( .A1(n6969), .A2(n6968), .ZN(n7087) );
  NAND2_X1 U6276 ( .A1(n6650), .A2(n6649), .ZN(n6761) );
  NOR2_X1 U6277 ( .A1(n6610), .A2(n6609), .ZN(n6647) );
  NAND3_X1 U6278 ( .A1(n8248), .A2(n8247), .A3(n4349), .ZN(n8257) );
  NAND2_X1 U6279 ( .A1(n6287), .A2(n6286), .ZN(n7700) );
  NAND2_X1 U6280 ( .A1(n4488), .A2(n4487), .ZN(n6993) );
  XNOR2_X2 U6281 ( .A(n5036), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6530) );
  NAND2_X1 U6282 ( .A1(n5669), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U6283 ( .A1(n9553), .A2(n6782), .ZN(n6784) );
  AOI21_X1 U6284 ( .B1(n9266), .B2(n4584), .A(n4583), .ZN(n4582) );
  NAND2_X1 U6285 ( .A1(n9593), .A2(n9395), .ZN(n4491) );
  AOI21_X1 U6286 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10037), .A(n10028), .ZN(
        n10042) );
  NOR2_X1 U6287 ( .A1(n9568), .A2(n10019), .ZN(n10030) );
  NAND2_X1 U6288 ( .A1(n5685), .A2(n5684), .ZN(n4573) );
  NAND2_X1 U6289 ( .A1(n4974), .A2(n4566), .ZN(n4565) );
  AOI21_X1 U6290 ( .B1(n4974), .B2(n4976), .A(n4384), .ZN(n4973) );
  OAI21_X2 U6291 ( .B1(n9634), .B2(n5712), .A(n5713), .ZN(n9619) );
  NAND2_X2 U6292 ( .A1(n9223), .A2(n9224), .ZN(n9679) );
  NAND3_X1 U6293 ( .A1(n6382), .A2(n6384), .A3(n6383), .ZN(n6412) );
  INV_X1 U6294 ( .A(n5041), .ZN(n5043) );
  NAND2_X1 U6295 ( .A1(n4954), .A2(n4953), .ZN(n6320) );
  NAND2_X1 U6296 ( .A1(n4459), .A2(n4381), .ZN(n9356) );
  NAND3_X1 U6297 ( .A1(n4504), .A2(n4611), .A3(n4609), .ZN(n4459) );
  OAI211_X1 U6298 ( .C1(n9399), .C2(n9291), .A(n4460), .B(n9290), .ZN(n9301)
         );
  NAND2_X1 U6299 ( .A1(n9289), .A2(n4380), .ZN(n4460) );
  OAI21_X1 U6300 ( .B1(n4582), .B2(n9446), .A(n4581), .ZN(n4580) );
  NAND3_X1 U6301 ( .A1(n5030), .A2(n5032), .A3(n5029), .ZN(n4461) );
  AOI21_X2 U6302 ( .B1(n7039), .B2(n7038), .A(n4998), .ZN(n9119) );
  XNOR2_X2 U6303 ( .A(n6854), .B(n10122), .ZN(n6852) );
  NAND2_X1 U6304 ( .A1(n4465), .A2(n4462), .ZN(P2_U3154) );
  NAND3_X1 U6305 ( .A1(n4483), .A2(n8003), .A3(n7830), .ZN(n4465) );
  NAND2_X1 U6306 ( .A1(n8006), .A2(n8005), .ZN(n8004) );
  NAND2_X1 U6307 ( .A1(n7024), .A2(n4482), .ZN(n7077) );
  NAND2_X2 U6308 ( .A1(n4813), .A2(n4811), .ZN(n9078) );
  NAND2_X1 U6309 ( .A1(n8933), .A2(n8932), .ZN(n8999) );
  NAND2_X2 U6310 ( .A1(n5465), .A2(n5487), .ZN(n6677) );
  NAND2_X1 U6311 ( .A1(n4485), .A2(n4484), .ZN(n4846) );
  NAND2_X1 U6312 ( .A1(n9421), .A2(n9758), .ZN(n5634) );
  OAI21_X1 U6313 ( .B1(n9619), .B2(n4331), .A(n5722), .ZN(n6317) );
  INV_X1 U6314 ( .A(n4975), .ZN(n4974) );
  NAND2_X1 U6315 ( .A1(n5689), .A2(n5705), .ZN(n9669) );
  NOR2_X2 U6316 ( .A1(n5678), .A2(n5677), .ZN(n4498) );
  NAND2_X1 U6317 ( .A1(n4501), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5663) );
  NAND2_X2 U6318 ( .A1(n8618), .A2(n6113), .ZN(n8605) );
  AOI21_X1 U6319 ( .B1(n6389), .B2(n8513), .A(n8512), .ZN(n8515) );
  NAND2_X1 U6320 ( .A1(n5179), .A2(n5178), .ZN(n5183) );
  NAND3_X1 U6321 ( .A1(n5069), .A2(n5070), .A3(SI_1_), .ZN(n5072) );
  NAND2_X1 U6322 ( .A1(n4933), .A2(n5185), .ZN(n5196) );
  XNOR2_X2 U6323 ( .A(n5226), .B(n5224), .ZN(n6489) );
  OAI21_X1 U6324 ( .B1(n8246), .B2(n6299), .A(n4550), .ZN(n4549) );
  NAND2_X1 U6325 ( .A1(n4726), .A2(n8408), .ZN(n4471) );
  NAND2_X1 U6326 ( .A1(n4731), .A2(n4732), .ZN(n8467) );
  INV_X1 U6327 ( .A(n4746), .ZN(n7097) );
  NAND3_X1 U6328 ( .A1(n4473), .A2(n8465), .A3(n4663), .ZN(n4472) );
  AOI21_X1 U6329 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6881), .A(n6870), .ZN(
        n6871) );
  NAND2_X2 U6330 ( .A1(n5858), .A2(n6430), .ZN(n8029) );
  OAI21_X2 U6331 ( .B1(n7114), .B2(n5910), .A(n6270), .ZN(n7011) );
  OR2_X2 U6332 ( .A1(n8605), .A2(n4880), .ZN(n4876) );
  NAND2_X2 U6333 ( .A1(n8092), .A2(n8094), .ZN(n6272) );
  NAND2_X1 U6334 ( .A1(n7687), .A2(n7686), .ZN(n4485) );
  NAND2_X1 U6335 ( .A1(n7411), .A2(n5981), .ZN(n7412) );
  NAND2_X1 U6336 ( .A1(n9100), .A2(n9101), .ZN(n9099) );
  OAI21_X2 U6337 ( .B1(n5335), .B2(n5334), .A(n5333), .ZN(n5343) );
  INV_X1 U6338 ( .A(n4533), .ZN(n4532) );
  OR2_X2 U6339 ( .A1(n8516), .A2(n8220), .ZN(n8221) );
  AOI21_X1 U6340 ( .B1(n4815), .B2(n4818), .A(n4812), .ZN(n4811) );
  INV_X1 U6341 ( .A(n4930), .ZN(n4929) );
  INV_X1 U6342 ( .A(n5203), .ZN(n4932) );
  NAND2_X1 U6343 ( .A1(n4445), .A2(n4921), .ZN(n4603) );
  BUF_X1 U6344 ( .A(n7040), .Z(n4480) );
  OAI21_X1 U6345 ( .B1(n5635), .B2(n4976), .A(n5642), .ZN(n4975) );
  NAND2_X1 U6346 ( .A1(n4358), .A2(n5247), .ZN(n5249) );
  XNOR2_X1 U6347 ( .A(n5249), .B(n5248), .ZN(n6062) );
  BUF_X2 U6348 ( .A(n5852), .Z(n5848) );
  INV_X1 U6349 ( .A(n4549), .ZN(n8248) );
  AND2_X1 U6350 ( .A1(n4295), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4683) );
  NAND2_X1 U6351 ( .A1(n8250), .A2(n8487), .ZN(n4550) );
  AOI21_X1 U6352 ( .B1(n8038), .B2(n8037), .A(n8036), .ZN(n8040) );
  NAND2_X1 U6353 ( .A1(n7829), .A2(n7828), .ZN(n4483) );
  NAND2_X1 U6354 ( .A1(n4867), .A2(n4865), .ZN(n7696) );
  NAND2_X1 U6355 ( .A1(n5196), .A2(n5195), .ZN(n5204) );
  INV_X1 U6356 ( .A(n5187), .ZN(n4933) );
  NAND2_X2 U6357 ( .A1(n5999), .A2(n5998), .ZN(n7971) );
  NAND2_X1 U6358 ( .A1(n4926), .A2(n4925), .ZN(n4924) );
  OAI21_X1 U6359 ( .B1(n4755), .B2(n4394), .A(n4747), .ZN(n4746) );
  NAND2_X1 U6360 ( .A1(n9369), .A2(n9384), .ZN(n4503) );
  NAND2_X1 U6361 ( .A1(n9341), .A2(n4400), .ZN(n4913) );
  OAI21_X1 U6362 ( .B1(n9308), .B2(n9309), .A(n9307), .ZN(n9310) );
  NAND3_X1 U6363 ( .A1(n8427), .A2(P2_REG2_REG_17__SCAN_IN), .A3(n8446), .ZN(
        n8447) );
  NAND2_X1 U6364 ( .A1(n4497), .A2(n9382), .ZN(n9371) );
  NAND2_X1 U6365 ( .A1(n4619), .A2(n4618), .ZN(n4497) );
  INV_X1 U6366 ( .A(n4624), .ZN(n4623) );
  INV_X1 U6367 ( .A(n4498), .ZN(n5688) );
  NAND2_X1 U6368 ( .A1(n4498), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5705) );
  INV_X1 U6369 ( .A(n4622), .ZN(n4621) );
  NAND3_X1 U6370 ( .A1(n9006), .A2(n9005), .A3(n4406), .ZN(P1_U3216) );
  NAND2_X2 U6371 ( .A1(n9052), .A2(n9053), .ZN(n9051) );
  NAND3_X1 U6372 ( .A1(n4503), .A2(n9371), .A3(n4502), .ZN(n4608) );
  NAND2_X1 U6373 ( .A1(n4580), .A2(n4579), .ZN(P1_U3242) );
  NAND2_X2 U6374 ( .A1(n9839), .A2(n9840), .ZN(n9838) );
  NAND2_X1 U6375 ( .A1(n9647), .A2(n4506), .ZN(n4509) );
  NAND2_X1 U6376 ( .A1(n4511), .A2(n4507), .ZN(n4510) );
  NAND2_X1 U6377 ( .A1(n4514), .A2(n9620), .ZN(n4507) );
  OAI211_X1 U6378 ( .C1(n9647), .C2(n4513), .A(n4510), .B(n4509), .ZN(n9618)
         );
  NAND2_X1 U6379 ( .A1(n5116), .A2(n5037), .ZN(n4516) );
  NAND2_X4 U6380 ( .A1(n4905), .A2(n4903), .ZN(n5116) );
  NAND2_X1 U6381 ( .A1(n9738), .A2(n4519), .ZN(n4517) );
  NAND3_X1 U6382 ( .A1(n4952), .A2(n5770), .A3(n9410), .ZN(n7278) );
  NOR2_X1 U6383 ( .A1(n4536), .A2(n8214), .ZN(n4533) );
  NAND2_X1 U6384 ( .A1(n8197), .A2(n8196), .ZN(n4542) );
  NAND2_X2 U6385 ( .A1(P1_U3086), .A2(n4544), .ZN(n9993) );
  MUX2_X1 U6386 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n5149), .Z(n5205) );
  MUX2_X1 U6387 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n5149), .Z(n5256) );
  MUX2_X1 U6388 ( .A(n6832), .B(n6830), .S(n4543), .Z(n5259) );
  MUX2_X1 U6389 ( .A(n5277), .B(n5278), .S(n4543), .Z(n5288) );
  MUX2_X1 U6390 ( .A(n6726), .B(n6724), .S(n4543), .Z(n5269) );
  MUX2_X1 U6391 ( .A(n7108), .B(n7110), .S(n4543), .Z(n5319) );
  MUX2_X1 U6392 ( .A(n7248), .B(n7250), .S(n4543), .Z(n5316) );
  MUX2_X1 U6393 ( .A(n7287), .B(n7290), .S(n4543), .Z(n5328) );
  MUX2_X1 U6394 ( .A(n7573), .B(n7654), .S(n4543), .Z(n5347) );
  MUX2_X1 U6395 ( .A(n7639), .B(n7638), .S(n4543), .Z(n5356) );
  MUX2_X1 U6396 ( .A(n7709), .B(n7717), .S(n4543), .Z(n5375) );
  MUX2_X1 U6397 ( .A(n7762), .B(n5838), .S(n4543), .Z(n5392) );
  MUX2_X1 U6398 ( .A(n5418), .B(n8028), .S(n4543), .Z(n5419) );
  NAND2_X1 U6399 ( .A1(n8170), .A2(n4548), .ZN(n4546) );
  NAND2_X1 U6400 ( .A1(n4546), .A2(n4547), .ZN(n8174) );
  OAI21_X1 U6401 ( .B1(n8170), .B2(n8171), .A(n4548), .ZN(n8183) );
  NAND2_X1 U6402 ( .A1(n4668), .A2(n4554), .ZN(n4553) );
  AND2_X2 U6403 ( .A1(n4559), .A2(n5985), .ZN(n7767) );
  OAI21_X1 U6404 ( .B1(n9788), .B2(n4975), .A(n4564), .ZN(n9736) );
  NAND2_X1 U6405 ( .A1(n4563), .A2(n4562), .ZN(n5654) );
  NAND2_X1 U6406 ( .A1(n9788), .A2(n4564), .ZN(n4562) );
  AND2_X2 U6407 ( .A1(n5067), .A2(n5149), .ZN(n5423) );
  NAND2_X1 U6408 ( .A1(n4573), .A2(n4572), .ZN(n4972) );
  AND3_X2 U6409 ( .A1(n5027), .A2(n5028), .A3(n5026), .ZN(n5029) );
  NAND3_X1 U6410 ( .A1(n9447), .A2(n9269), .A3(n9268), .ZN(n4583) );
  NAND2_X1 U6411 ( .A1(n5291), .A2(n4589), .ZN(n4588) );
  NAND2_X1 U6412 ( .A1(n5353), .A2(n4596), .ZN(n4592) );
  NAND2_X1 U6413 ( .A1(n4445), .A2(n4600), .ZN(n4599) );
  AOI21_X1 U6414 ( .B1(n4608), .B2(n9375), .A(n4934), .ZN(n9392) );
  NAND2_X1 U6415 ( .A1(n9365), .A2(n4621), .ZN(n4618) );
  AOI21_X1 U6416 ( .B1(n4629), .B2(n4628), .A(n4627), .ZN(n4626) );
  NAND2_X1 U6417 ( .A1(n7218), .A2(n7221), .ZN(n7233) );
  NAND2_X1 U6418 ( .A1(n9317), .A2(n4637), .ZN(n4635) );
  NAND2_X1 U6419 ( .A1(n4635), .A2(n4633), .ZN(n4926) );
  NAND2_X1 U6420 ( .A1(n7356), .A2(n7357), .ZN(n4661) );
  AND2_X1 U6421 ( .A1(n7142), .A2(n7143), .ZN(n4662) );
  NAND3_X1 U6422 ( .A1(n4672), .A2(n4675), .A3(n4383), .ZN(n4671) );
  NAND4_X1 U6423 ( .A1(n5834), .A2(n5833), .A3(n4900), .A4(n5842), .ZN(n5845)
         );
  AND3_X2 U6424 ( .A1(n5834), .A2(n5833), .A3(n4679), .ZN(n8810) );
  NAND3_X1 U6425 ( .A1(n5834), .A2(n5833), .A3(n4900), .ZN(n5841) );
  INV_X2 U6426 ( .A(n6851), .ZN(n6928) );
  NAND2_X1 U6427 ( .A1(n8511), .A2(n8224), .ZN(n4690) );
  OAI21_X2 U6428 ( .B1(n8511), .B2(n4687), .A(n4685), .ZN(n8017) );
  NAND2_X1 U6429 ( .A1(n7407), .A2(n4385), .ZN(n4691) );
  NAND3_X1 U6430 ( .A1(n4693), .A2(n8150), .A3(n4691), .ZN(n7658) );
  INV_X1 U6431 ( .A(n8143), .ZN(n4696) );
  OR2_X1 U6432 ( .A1(n4695), .A2(n4694), .ZN(n4693) );
  NAND2_X1 U6433 ( .A1(n7408), .A2(n8139), .ZN(n7642) );
  INV_X1 U6434 ( .A(n8139), .ZN(n4699) );
  NAND2_X1 U6435 ( .A1(n6271), .A2(n4700), .ZN(n5893) );
  NAND2_X1 U6436 ( .A1(n7998), .A2(n4700), .ZN(n6891) );
  AOI22_X1 U6437 ( .A1(n8666), .A2(n4700), .B1(n7130), .B2(n8677), .ZN(n7131)
         );
  AND2_X2 U6438 ( .A1(n5892), .A2(n4340), .ZN(n10132) );
  OAI21_X2 U6439 ( .B1(n6408), .B2(n4701), .A(n8216), .ZN(n8547) );
  OAI21_X2 U6440 ( .B1(n7700), .B2(n8165), .A(n7697), .ZN(n7729) );
  INV_X2 U6441 ( .A(n7138), .ZN(n10122) );
  NAND3_X1 U6442 ( .A1(n5875), .A2(n5876), .A3(n4391), .ZN(n7138) );
  NAND2_X1 U6443 ( .A1(n4703), .A2(n4702), .ZN(n8560) );
  NAND3_X1 U6444 ( .A1(n5834), .A2(n4899), .A3(n5833), .ZN(n6237) );
  NAND2_X1 U6445 ( .A1(n6167), .A2(n6185), .ZN(n8545) );
  NAND2_X1 U6446 ( .A1(n6157), .A2(n4706), .ZN(n6185) );
  NAND2_X1 U6447 ( .A1(n6157), .A2(n6156), .ZN(n6166) );
  NAND2_X1 U6448 ( .A1(n6104), .A2(n4407), .ZN(n6136) );
  NAND3_X1 U6449 ( .A1(n6334), .A2(n4309), .A3(n4717), .ZN(n8071) );
  NAND3_X1 U6450 ( .A1(n4723), .A2(n4990), .A3(n4722), .ZN(n7292) );
  NAND3_X1 U6451 ( .A1(n4724), .A2(n7155), .A3(n4315), .ZN(n4722) );
  INV_X1 U6452 ( .A(n7099), .ZN(n4725) );
  INV_X1 U6453 ( .A(n8381), .ZN(n4726) );
  NAND3_X1 U6454 ( .A1(n8427), .A2(n8446), .A3(n4729), .ZN(n4731) );
  INV_X1 U6455 ( .A(n8335), .ZN(n4734) );
  AOI21_X1 U6456 ( .B1(n4734), .B2(n8341), .A(n4737), .ZN(n4736) );
  AOI21_X1 U6457 ( .B1(n8335), .B2(n8334), .A(n8355), .ZN(n4735) );
  NAND2_X1 U6458 ( .A1(n8335), .A2(n4405), .ZN(n4740) );
  OAI21_X1 U6459 ( .B1(n8334), .B2(n8355), .A(P2_REG2_REG_13__SCAN_IN), .ZN(
        n4737) );
  NAND2_X1 U6460 ( .A1(n4739), .A2(n8341), .ZN(n8363) );
  NAND2_X1 U6461 ( .A1(n8335), .A2(n8334), .ZN(n4739) );
  NAND2_X1 U6462 ( .A1(n7363), .A2(n7362), .ZN(n4741) );
  NAND2_X1 U6463 ( .A1(n7293), .A2(n7361), .ZN(n7294) );
  OR2_X1 U6464 ( .A1(n8295), .A2(n8286), .ZN(n4745) );
  INV_X1 U6465 ( .A(n6871), .ZN(n4751) );
  NOR2_X1 U6466 ( .A1(n8289), .A2(n8290), .ZN(n8313) );
  NAND2_X1 U6467 ( .A1(n8310), .A2(n8288), .ZN(n8289) );
  NAND2_X1 U6468 ( .A1(n8379), .A2(n5008), .ZN(n8380) );
  AND2_X1 U6469 ( .A1(n6196), .A2(n4887), .ZN(n4886) );
  OAI21_X2 U6470 ( .B1(n8313), .B2(n8312), .A(n8311), .ZN(n8335) );
  NAND2_X2 U6471 ( .A1(n5874), .A2(n5873), .ZN(n6606) );
  OAI21_X2 U6472 ( .B1(n7089), .B2(n7088), .A(n7087), .ZN(n7145) );
  OR2_X4 U6473 ( .A1(n6145), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6175) );
  AND2_X1 U6474 ( .A1(n6663), .A2(n6747), .ZN(n6664) );
  NAND3_X1 U6475 ( .A1(n4771), .A2(P2_REG1_REG_11__SCAN_IN), .A3(n8320), .ZN(
        n8321) );
  INV_X1 U6476 ( .A(n4773), .ZN(n4772) );
  OAI21_X2 U6477 ( .B1(n4775), .B2(n5001), .A(n4774), .ZN(n7091) );
  INV_X1 U6478 ( .A(n6971), .ZN(n4775) );
  OAI21_X1 U6479 ( .B1(n7299), .B2(n4782), .A(n4778), .ZN(n7370) );
  NAND2_X1 U6480 ( .A1(n7368), .A2(n4785), .ZN(n7301) );
  INV_X1 U6481 ( .A(n8343), .ZN(n4786) );
  NAND2_X1 U6482 ( .A1(n4786), .A2(n8358), .ZN(n4787) );
  NAND2_X1 U6483 ( .A1(n4787), .A2(n4788), .ZN(n8393) );
  OAI211_X2 U6484 ( .C1(n6585), .C2(n4791), .A(n5888), .B(n4790), .ZN(n6659)
         );
  AND2_X2 U6485 ( .A1(n7379), .A2(n4792), .ZN(n9830) );
  AND2_X2 U6486 ( .A1(n9695), .A2(n4797), .ZN(n9651) );
  NAND2_X1 U6487 ( .A1(n6318), .A2(n4806), .ZN(n9603) );
  NAND2_X1 U6488 ( .A1(n6318), .A2(n9870), .ZN(n6362) );
  NAND3_X1 U6489 ( .A1(n5085), .A2(n5086), .A3(n4809), .ZN(n7181) );
  NAND3_X1 U6490 ( .A1(n9038), .A2(n9196), .A3(n9039), .ZN(n4810) );
  NAND2_X1 U6491 ( .A1(n9087), .A2(n8879), .ZN(n8885) );
  NAND2_X1 U6492 ( .A1(n9051), .A2(n4823), .ZN(n8933) );
  NAND2_X1 U6493 ( .A1(n4826), .A2(n5007), .ZN(n4825) );
  NAND2_X1 U6494 ( .A1(n8843), .A2(n4827), .ZN(n4826) );
  NAND2_X1 U6495 ( .A1(n9099), .A2(n4833), .ZN(n8902) );
  NAND2_X1 U6496 ( .A1(n8004), .A2(n4838), .ZN(n4834) );
  NAND2_X1 U6497 ( .A1(n4834), .A2(n4835), .ZN(n7801) );
  NAND2_X1 U6498 ( .A1(n8004), .A2(n5000), .ZN(n7906) );
  NOR2_X1 U6499 ( .A1(n7787), .A2(n4842), .ZN(n4841) );
  INV_X1 U6500 ( .A(n5000), .ZN(n4842) );
  NAND2_X1 U6501 ( .A1(n6063), .A2(n4849), .ZN(n5815) );
  NAND2_X1 U6502 ( .A1(n4852), .A2(n4853), .ZN(n7829) );
  NAND2_X2 U6503 ( .A1(n4852), .A2(n4850), .ZN(n7830) );
  NAND2_X1 U6504 ( .A1(n4855), .A2(n4854), .ZN(n7559) );
  NOR2_X1 U6505 ( .A1(n7456), .A2(n4307), .ZN(n7555) );
  NAND2_X1 U6506 ( .A1(n7958), .A2(n4860), .ZN(n7807) );
  NAND2_X2 U6507 ( .A1(n5834), .A2(n5827), .ZN(n6047) );
  OAI21_X1 U6508 ( .B1(n7643), .B2(n4870), .A(n4868), .ZN(n7627) );
  AOI21_X2 U6509 ( .B1(n4868), .B2(n4870), .A(n4866), .ZN(n4865) );
  NAND2_X1 U6510 ( .A1(n7643), .A2(n4868), .ZN(n4867) );
  NAND2_X2 U6511 ( .A1(n4869), .A2(n6033), .ZN(n4868) );
  NAND2_X1 U6512 ( .A1(n4876), .A2(n4877), .ZN(n8580) );
  OAI21_X1 U6513 ( .B1(n6142), .B2(n4885), .A(n4882), .ZN(n6332) );
  INV_X1 U6514 ( .A(n6332), .ZN(n6343) );
  OAI21_X2 U6515 ( .B1(n8569), .B2(n6153), .A(n6152), .ZN(n6389) );
  INV_X1 U6516 ( .A(n7011), .ZN(n4897) );
  NAND2_X1 U6517 ( .A1(n4893), .A2(n4894), .ZN(n7165) );
  NAND2_X1 U6518 ( .A1(n7011), .A2(n7166), .ZN(n4893) );
  NAND2_X1 U6519 ( .A1(n4898), .A2(n4389), .ZN(n7411) );
  NAND2_X1 U6520 ( .A1(n8636), .A2(n4901), .ZN(n8618) );
  AND2_X1 U6521 ( .A1(n5043), .A2(n5042), .ZN(n5068) );
  NAND3_X1 U6522 ( .A1(n4904), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4903) );
  NAND3_X1 U6523 ( .A1(n5128), .A2(n5127), .A3(n4906), .ZN(n4908) );
  NOR2_X1 U6524 ( .A1(n5166), .A2(n4907), .ZN(n4906) );
  INV_X1 U6525 ( .A(n5170), .ZN(n4907) );
  NAND2_X1 U6526 ( .A1(n5165), .A2(n5170), .ZN(n4909) );
  NAND2_X1 U6527 ( .A1(n5128), .A2(n5127), .ZN(n5167) );
  NAND2_X1 U6528 ( .A1(n9312), .A2(n4914), .ZN(n4911) );
  INV_X1 U6529 ( .A(n9330), .ZN(n4914) );
  NAND2_X1 U6530 ( .A1(n5187), .A2(n4928), .ZN(n4927) );
  NAND2_X1 U6531 ( .A1(n6795), .A2(n9404), .ZN(n4937) );
  NAND2_X1 U6532 ( .A1(n9275), .A2(n5764), .ZN(n6908) );
  AND2_X2 U6533 ( .A1(n5034), .A2(n5014), .ZN(n5080) );
  NAND2_X1 U6534 ( .A1(n9806), .A2(n9807), .ZN(n9805) );
  NAND2_X1 U6535 ( .A1(n9679), .A2(n4946), .ZN(n4945) );
  OAI21_X1 U6536 ( .B1(n9679), .B2(n4947), .A(n4946), .ZN(n9648) );
  NAND2_X2 U6537 ( .A1(n4945), .A2(n4943), .ZN(n9647) );
  NAND2_X1 U6538 ( .A1(n9630), .A2(n4388), .ZN(n4954) );
  NAND2_X1 U6539 ( .A1(n6905), .A2(n4959), .ZN(n4958) );
  NAND2_X1 U6540 ( .A1(n4972), .A2(n4971), .ZN(n5702) );
  INV_X1 U6541 ( .A(n9722), .ZN(n4983) );
  NAND2_X1 U6542 ( .A1(n4977), .A2(n4978), .ZN(n5685) );
  NAND2_X1 U6543 ( .A1(n9722), .A2(n4980), .ZN(n4977) );
  NAND2_X1 U6544 ( .A1(n9619), .A2(n4988), .ZN(n4984) );
  NAND2_X1 U6545 ( .A1(n4984), .A2(n4985), .ZN(n6356) );
  INV_X1 U6546 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9595) );
  XOR2_X1 U6547 ( .A(n8511), .B(n8516), .Z(n8754) );
  AOI21_X1 U6548 ( .B1(n6398), .B2(n8640), .A(n6397), .ZN(n8760) );
  OAI21_X1 U6549 ( .B1(n6394), .B2(n8212), .A(n8539), .ZN(n6398) );
  NAND2_X1 U6550 ( .A1(n8520), .A2(n8573), .ZN(n8521) );
  NAND2_X1 U6551 ( .A1(n8520), .A2(n8571), .ZN(n6396) );
  NAND2_X1 U6552 ( .A1(n8017), .A2(n8233), .ZN(n8038) );
  NAND2_X2 U6553 ( .A1(n5046), .A2(n5045), .ZN(n5069) );
  INV_X1 U6554 ( .A(n5502), .ZN(n5509) );
  MUX2_X2 U6555 ( .A(n8690), .B(n8755), .S(n10168), .Z(n8692) );
  MUX2_X2 U6556 ( .A(n10301), .B(n8755), .S(n10155), .Z(n8759) );
  CLKBUF_X1 U6557 ( .A(n8321), .Z(n8317) );
  MUX2_X2 U6558 ( .A(n8544), .B(n8755), .S(n8663), .Z(n8550) );
  NAND2_X1 U6559 ( .A1(n8342), .A2(n8341), .ZN(n8358) );
  INV_X1 U6560 ( .A(n6213), .ZN(n6847) );
  NAND2_X1 U6561 ( .A1(n7093), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7147) );
  CLKBUF_X1 U6562 ( .A(n9757), .Z(n9770) );
  NAND2_X1 U6563 ( .A1(n5236), .A2(n5235), .ZN(n5245) );
  AND2_X1 U6564 ( .A1(n9234), .A2(n9376), .ZN(n9235) );
  AND2_X1 U6565 ( .A1(n6659), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6652) );
  CLKBUF_X1 U6566 ( .A(n9065), .Z(n9175) );
  OAI21_X1 U6567 ( .B1(n5417), .B2(n5416), .A(n5415), .ZN(n5421) );
  AOI21_X2 U6568 ( .B1(n6864), .B2(n6863), .A(n6853), .ZN(n6898) );
  XNOR2_X2 U6569 ( .A(n6852), .B(n8277), .ZN(n6864) );
  AND2_X1 U6570 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  INV_X1 U6571 ( .A(n4300), .ZN(n6686) );
  INV_X1 U6572 ( .A(n5487), .ZN(n7674) );
  NAND2_X1 U6573 ( .A1(n5474), .A2(n5487), .ZN(n6674) );
  OAI21_X1 U6574 ( .B1(n5116), .B2(n5097), .A(n5096), .ZN(n5098) );
  NAND2_X1 U6575 ( .A1(n5116), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5096) );
  OAI21_X1 U6576 ( .B1(n5116), .B2(n5039), .A(n5038), .ZN(n5042) );
  NAND2_X1 U6577 ( .A1(n5116), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5038) );
  OAI21_X2 U6578 ( .B1(n8547), .B2(n8219), .A(n8067), .ZN(n8511) );
  INV_X1 U6579 ( .A(n6956), .ZN(n9471) );
  NAND2_X1 U6580 ( .A1(n5880), .A2(n5862), .ZN(n8094) );
  CLKBUF_X3 U6581 ( .A(n5513), .Z(n5732) );
  INV_X1 U6582 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U6583 ( .A1(n7827), .A2(n8818), .ZN(n5960) );
  INV_X1 U6584 ( .A(n7827), .ZN(n5849) );
  OR2_X1 U6585 ( .A1(n7297), .A2(n7291), .ZN(n4990) );
  INV_X1 U6586 ( .A(n5513), .ZN(n5742) );
  AND2_X1 U6587 ( .A1(n8204), .A2(n8562), .ZN(n4991) );
  NOR4_X1 U6588 ( .A1(n9646), .A2(n9703), .A3(n9258), .A4(n9680), .ZN(n4992)
         );
  AND2_X1 U6589 ( .A1(n6820), .A2(n6261), .ZN(n6484) );
  NAND2_X2 U6590 ( .A1(n5752), .A2(n9852), .ZN(n9855) );
  AND2_X1 U6591 ( .A1(n10117), .A2(n9940), .ZN(n9899) );
  INV_X1 U6592 ( .A(n9981), .ZN(n6326) );
  OR2_X1 U6593 ( .A1(n9600), .A2(n9981), .ZN(n4993) );
  AND2_X1 U6594 ( .A1(n10156), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n4994) );
  AND2_X1 U6595 ( .A1(n7900), .A2(n8677), .ZN(n4995) );
  OR2_X1 U6596 ( .A1(n9385), .A2(n9383), .ZN(n4996) );
  INV_X1 U6597 ( .A(n8206), .ZN(n6296) );
  AND2_X1 U6598 ( .A1(n6419), .A2(n8801), .ZN(n6353) );
  NAND2_X1 U6599 ( .A1(n6379), .A2(n6378), .ZN(n4997) );
  AND2_X1 U6600 ( .A1(n7037), .A2(n7036), .ZN(n4998) );
  AND2_X1 U6601 ( .A1(n7780), .A2(n7950), .ZN(n4999) );
  OR2_X1 U6602 ( .A1(n7782), .A2(n7838), .ZN(n5000) );
  XOR2_X1 U6603 ( .A(n7767), .B(n7813), .Z(n5002) );
  AND2_X1 U6604 ( .A1(n9092), .A2(n8884), .ZN(n5003) );
  INV_X1 U6605 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5039) );
  INV_X1 U6606 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5151) );
  NOR2_X1 U6607 ( .A1(n4808), .A2(n9981), .ZN(n6365) );
  AND2_X1 U6608 ( .A1(n6607), .A2(n6606), .ZN(n5004) );
  OR2_X1 U6609 ( .A1(n5451), .A2(n5450), .ZN(n5005) );
  INV_X1 U6610 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6098) );
  INV_X1 U6611 ( .A(n6509), .ZN(n5061) );
  AND2_X1 U6612 ( .A1(n7814), .A2(n8003), .ZN(n5006) );
  AND2_X1 U6613 ( .A1(n9173), .A2(n8851), .ZN(n5007) );
  OR2_X1 U6614 ( .A1(n8378), .A2(n8377), .ZN(n5008) );
  INV_X1 U6615 ( .A(n10113), .ZN(n9943) );
  NAND2_X1 U6616 ( .A1(n9667), .A2(n9459), .ZN(n5010) );
  INV_X1 U6617 ( .A(n9349), .ZN(n5776) );
  AND2_X1 U6618 ( .A1(n7786), .A2(n7978), .ZN(n5011) );
  XNOR2_X1 U6619 ( .A(n5313), .B(n5312), .ZN(n6125) );
  OR2_X1 U6620 ( .A1(n7429), .A2(n7557), .ZN(n5012) );
  OR2_X1 U6621 ( .A1(n5255), .A2(SI_14_), .ZN(n5013) );
  AND2_X1 U6622 ( .A1(n8082), .A2(n8255), .ZN(n8083) );
  MUX2_X1 U6623 ( .A(n8222), .B(n8089), .S(n8088), .Z(n8091) );
  NOR2_X1 U6624 ( .A1(n8115), .A2(n8222), .ZN(n8116) );
  NAND2_X1 U6625 ( .A1(n8117), .A2(n8116), .ZN(n8118) );
  AND2_X1 U6626 ( .A1(n9701), .A2(n9340), .ZN(n9332) );
  INV_X1 U6627 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5810) );
  INV_X1 U6628 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5828) );
  NAND2_X1 U6629 ( .A1(n7938), .A2(n7788), .ZN(n7789) );
  AND2_X1 U6630 ( .A1(n8100), .A2(n7111), .ZN(n6275) );
  AND2_X1 U6631 ( .A1(n8114), .A2(n8127), .ZN(n7401) );
  INV_X1 U6632 ( .A(n9007), .ZN(n8849) );
  INV_X1 U6633 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5024) );
  OR2_X1 U6634 ( .A1(n8338), .A2(n8333), .ZN(n8334) );
  INV_X1 U6635 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U6636 ( .A1(n8850), .A2(n8849), .ZN(n8851) );
  AND2_X1 U6637 ( .A1(n5025), .A2(n5024), .ZN(n5026) );
  OR2_X1 U6638 ( .A1(n7419), .A2(n8123), .ZN(n7420) );
  NAND2_X1 U6639 ( .A1(n6214), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U6640 ( .A1(n8278), .A2(n6850), .ZN(n6926) );
  INV_X1 U6641 ( .A(n9646), .ZN(n5778) );
  INV_X1 U6642 ( .A(SI_15_), .ZN(n10300) );
  NAND2_X1 U6643 ( .A1(n5509), .A2(n5503), .ZN(n5760) );
  NAND2_X1 U6644 ( .A1(n5431), .A2(n5430), .ZN(n5432) );
  INV_X1 U6645 ( .A(SI_19_), .ZN(n5292) );
  INV_X1 U6646 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10223) );
  OR2_X1 U6647 ( .A1(n7803), .A2(n8574), .ZN(n7804) );
  AND2_X1 U6648 ( .A1(n8072), .A2(n8742), .ZN(n8036) );
  INV_X1 U6649 ( .A(n8865), .ZN(n8866) );
  AND2_X1 U6650 ( .A1(n8943), .A2(n8942), .ZN(n9110) );
  NAND2_X1 U6651 ( .A1(n5062), .A2(n5061), .ZN(n5063) );
  INV_X1 U6652 ( .A(n5210), .ZN(n5141) );
  INV_X1 U6653 ( .A(n8845), .ZN(n5201) );
  NAND2_X1 U6654 ( .A1(n6736), .A2(n9123), .ZN(n9280) );
  INV_X1 U6655 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n10206) );
  AND2_X1 U6656 ( .A1(n10101), .A2(n7265), .ZN(n7263) );
  NAND2_X1 U6657 ( .A1(n5293), .A2(n5292), .ZN(n5306) );
  NAND2_X1 U6658 ( .A1(n5205), .A2(SI_12_), .ZN(n5218) );
  INV_X1 U6659 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5896) );
  OR2_X1 U6660 ( .A1(P2_U3150), .A2(n6573), .ZN(n8371) );
  INV_X1 U6661 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6420) );
  OR2_X1 U6662 ( .A1(n8165), .A2(n8164), .ZN(n8163) );
  INV_X1 U6663 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6229) );
  AOI22_X1 U6664 ( .A1(n5423), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6449), .B2(
        n6548), .ZN(n5095) );
  INV_X1 U6665 ( .A(n5746), .ZN(n6413) );
  AND2_X1 U6666 ( .A1(n10089), .A2(n9267), .ZN(n9782) );
  AND4_X1 U6667 ( .A1(n5608), .A2(n5607), .A3(n5606), .A4(n5605), .ZN(n9809)
         );
  NOR2_X2 U6668 ( .A1(n7198), .A2(n7221), .ZN(n7230) );
  AND2_X1 U6669 ( .A1(n5372), .A2(n5367), .ZN(n5370) );
  XNOR2_X1 U6670 ( .A(n5288), .B(SI_18_), .ZN(n5287) );
  XNOR2_X1 U6671 ( .A(n5168), .B(SI_8_), .ZN(n5161) );
  INV_X1 U6672 ( .A(n8009), .ZN(n7984) );
  AOI22_X1 U6673 ( .A1(n7077), .A2(n7076), .B1(n7075), .B2(n7074), .ZN(n7079)
         );
  AOI21_X1 U6674 ( .B1(n7836), .B2(n7835), .A(n4999), .ZN(n8006) );
  INV_X1 U6675 ( .A(n8488), .ZN(n8373) );
  INV_X1 U6676 ( .A(n8681), .ZN(n6405) );
  NOR2_X1 U6677 ( .A1(n7755), .A2(n8696), .ZN(n6422) );
  INV_X1 U6678 ( .A(n8716), .ZN(n8734) );
  INV_X1 U6679 ( .A(n8790), .ZN(n8802) );
  NAND2_X1 U6680 ( .A1(n7648), .A2(n10127), .ZN(n10153) );
  INV_X1 U6681 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5469) );
  INV_X1 U6682 ( .A(n9167), .ZN(n9202) );
  AND4_X1 U6683 ( .A1(n5615), .A2(n5614), .A3(n5613), .A4(n5612), .ZN(n9211)
         );
  INV_X1 U6684 ( .A(n10055), .ZN(n10047) );
  INV_X1 U6685 ( .A(n9239), .ZN(n9703) );
  INV_X1 U6686 ( .A(n9783), .ZN(n10076) );
  NAND2_X1 U6687 ( .A1(n5780), .A2(n9394), .ZN(n9846) );
  NOR2_X1 U6688 ( .A1(n10117), .A2(n5493), .ZN(n5494) );
  AND2_X1 U6689 ( .A1(n10089), .A2(n9443), .ZN(n9940) );
  NAND2_X1 U6690 ( .A1(n9815), .A2(n7547), .ZN(n10113) );
  INV_X1 U6691 ( .A(n6672), .ZN(n5803) );
  AND2_X1 U6692 ( .A1(n5192), .A2(n5197), .ZN(n6779) );
  INV_X1 U6693 ( .A(n8011), .ZN(n7953) );
  INV_X1 U6694 ( .A(n8003), .ZN(n8000) );
  AND2_X1 U6695 ( .A1(n8027), .A2(n6222), .ZN(n7818) );
  INV_X1 U6696 ( .A(n8638), .ZN(n8262) );
  OR2_X1 U6697 ( .A1(n6571), .A2(n6570), .ZN(n8488) );
  OR2_X1 U6698 ( .A1(n8457), .A2(n8251), .ZN(n8482) );
  OR2_X1 U6699 ( .A1(n6583), .A2(n8405), .ZN(n8495) );
  INV_X1 U6700 ( .A(n8663), .ZN(n8681) );
  INV_X1 U6701 ( .A(n8678), .ZN(n8669) );
  NOR2_X1 U6702 ( .A1(n6422), .A2(n6421), .ZN(n6423) );
  INV_X1 U6703 ( .A(n8733), .ZN(n8696) );
  OR2_X1 U6704 ( .A1(n8508), .A2(n8790), .ZN(n6315) );
  OR2_X1 U6705 ( .A1(n10156), .A2(n10133), .ZN(n8790) );
  AND2_X1 U6706 ( .A1(n6313), .A2(n6312), .ZN(n10156) );
  INV_X1 U6707 ( .A(n6484), .ZN(n6478) );
  INV_X1 U6708 ( .A(n5852), .ZN(n8818) );
  INV_X1 U6709 ( .A(n8255), .ZN(n7288) );
  INV_X1 U6710 ( .A(n7357), .ZN(n7300) );
  INV_X1 U6711 ( .A(n9968), .ZN(n9697) );
  INV_X1 U6712 ( .A(n9903), .ZN(n9717) );
  INV_X1 U6713 ( .A(n9939), .ZN(n9837) );
  INV_X1 U6714 ( .A(n9950), .ZN(n9625) );
  INV_X1 U6715 ( .A(n9199), .ZN(n9455) );
  OR2_X1 U6716 ( .A1(n6518), .A2(n9448), .ZN(n10060) );
  OR2_X1 U6717 ( .A1(n6518), .A2(n6514), .ZN(n10055) );
  INV_X1 U6718 ( .A(n10033), .ZN(n10070) );
  NAND2_X1 U6719 ( .A1(n6381), .A2(n6357), .ZN(n7751) );
  INV_X1 U6720 ( .A(n10071), .ZN(n9850) );
  INV_X2 U6721 ( .A(n10117), .ZN(n10118) );
  NAND2_X1 U6722 ( .A1(n10348), .A2(n9940), .ZN(n9981) );
  INV_X1 U6723 ( .A(n10348), .ZN(n10346) );
  AND2_X2 U6724 ( .A1(n5804), .A2(n5803), .ZN(n10348) );
  INV_X1 U6725 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7573) );
  INV_X1 U6726 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7004) );
  INV_X1 U6727 ( .A(n8457), .ZN(P2_U3893) );
  NAND2_X1 U6728 ( .A1(n6411), .A2(n6410), .ZN(P2_U3208) );
  AND2_X1 U6729 ( .A1(n6425), .A2(n6678), .ZN(P1_U3973) );
  AND2_X2 U6730 ( .A1(n5020), .A2(n5019), .ZN(n5153) );
  NOR2_X1 U6731 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5023) );
  NAND3_X1 U6732 ( .A1(n5453), .A2(n5023), .A3(n5426), .ZN(n5451) );
  INV_X1 U6733 ( .A(n5451), .ZN(n5028) );
  INV_X2 U6734 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5281) );
  NAND4_X1 U6735 ( .A1(n5435), .A2(n4435), .A3(n5281), .A4(n5454), .ZN(n5450)
         );
  INV_X1 U6736 ( .A(n5450), .ZN(n5027) );
  INV_X1 U6737 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5035) );
  OR2_X1 U6738 ( .A1(n5034), .A2(n5035), .ZN(n5036) );
  INV_X1 U6739 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5868) );
  INV_X1 U6740 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5037) );
  INV_X1 U6741 ( .A(SI_0_), .ZN(n5867) );
  NAND2_X1 U6742 ( .A1(n5041), .A2(n5040), .ZN(n5070) );
  NAND2_X1 U6743 ( .A1(n5051), .A2(SI_1_), .ZN(n5055) );
  INV_X1 U6744 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6438) );
  INV_X1 U6745 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5044) );
  MUX2_X1 U6746 ( .A(n6438), .B(n5044), .S(n5116), .Z(n5046) );
  INV_X1 U6747 ( .A(SI_2_), .ZN(n5045) );
  INV_X1 U6748 ( .A(n5046), .ZN(n5047) );
  NAND2_X1 U6749 ( .A1(n5047), .A2(SI_2_), .ZN(n5071) );
  NAND2_X1 U6750 ( .A1(n5069), .A2(n5071), .ZN(n5048) );
  XNOR2_X1 U6751 ( .A(n5049), .B(n5048), .ZN(n6437) );
  NAND2_X1 U6752 ( .A1(n6437), .A2(n5141), .ZN(n5050) );
  INV_X2 U6753 ( .A(n10073), .ZN(n6801) );
  INV_X1 U6754 ( .A(n5051), .ZN(n5053) );
  INV_X1 U6755 ( .A(SI_1_), .ZN(n5052) );
  NAND2_X1 U6756 ( .A1(n5053), .A2(n5052), .ZN(n5054) );
  NAND2_X1 U6757 ( .A1(n5055), .A2(n5054), .ZN(n6461) );
  OR2_X1 U6758 ( .A1(n6461), .A2(n5210), .ZN(n5065) );
  INV_X1 U6759 ( .A(n7763), .ZN(n6517) );
  INV_X1 U6760 ( .A(n7708), .ZN(n6514) );
  AND2_X1 U6761 ( .A1(n5149), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5057) );
  OAI21_X1 U6762 ( .B1(n6517), .B2(n6514), .A(n5057), .ZN(n5064) );
  NAND2_X1 U6763 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4469), .ZN(n5058) );
  MUX2_X1 U6764 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5058), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5060) );
  INV_X1 U6765 ( .A(n5034), .ZN(n5059) );
  NAND2_X1 U6766 ( .A1(n5060), .A2(n5059), .ZN(n6509) );
  NAND3_X1 U6767 ( .A1(n5065), .A2(n5064), .A3(n5063), .ZN(n5503) );
  NAND2_X1 U6768 ( .A1(n6430), .A2(SI_0_), .ZN(n5066) );
  XNOR2_X1 U6769 ( .A(n5066), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9999) );
  MUX2_X1 U6770 ( .A(n4469), .B(n9999), .S(n5067), .Z(n10090) );
  INV_X1 U6771 ( .A(n10090), .ZN(n7265) );
  INV_X1 U6772 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U6773 ( .A1(n5068), .A2(n5069), .ZN(n5073) );
  INV_X1 U6774 ( .A(n5078), .ZN(n5075) );
  MUX2_X1 U6775 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5116), .Z(n5074) );
  NAND2_X1 U6776 ( .A1(n5074), .A2(SI_3_), .ZN(n5101) );
  OAI21_X1 U6777 ( .B1(n5074), .B2(SI_3_), .A(n5101), .ZN(n5076) );
  NAND2_X1 U6778 ( .A1(n5075), .A2(n5076), .ZN(n5079) );
  INV_X1 U6779 ( .A(n5076), .ZN(n5077) );
  NAND2_X1 U6780 ( .A1(n5079), .A2(n5122), .ZN(n6458) );
  OR2_X1 U6781 ( .A1(n6458), .A2(n5210), .ZN(n5086) );
  NOR2_X1 U6782 ( .A1(n5154), .A2(n5035), .ZN(n5081) );
  MUX2_X1 U6783 ( .A(n5035), .B(n5081), .S(P1_IR_REG_3__SCAN_IN), .Z(n5084) );
  INV_X1 U6784 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U6785 ( .A1(n5154), .A2(n5082), .ZN(n5108) );
  INV_X1 U6786 ( .A(n5108), .ZN(n5083) );
  NAND2_X1 U6787 ( .A1(n6449), .A2(n9488), .ZN(n5085) );
  NAND2_X1 U6788 ( .A1(n7177), .A2(n10111), .ZN(n7176) );
  NAND2_X1 U6789 ( .A1(n5108), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U6790 ( .A(n5087), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6548) );
  NAND2_X1 U6791 ( .A1(n5122), .A2(n5101), .ZN(n5092) );
  MUX2_X1 U6792 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n5116), .Z(n5088) );
  NAND2_X1 U6793 ( .A1(n5088), .A2(SI_4_), .ZN(n5100) );
  INV_X1 U6794 ( .A(n5088), .ZN(n5090) );
  INV_X1 U6795 ( .A(SI_4_), .ZN(n5089) );
  NAND2_X1 U6796 ( .A1(n5090), .A2(n5089), .ZN(n5103) );
  AND2_X1 U6797 ( .A1(n5100), .A2(n5103), .ZN(n5091) );
  OR2_X1 U6798 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  NAND2_X1 U6799 ( .A1(n5092), .A2(n5091), .ZN(n5099) );
  AND2_X1 U6800 ( .A1(n5093), .A2(n5099), .ZN(n6429) );
  NAND2_X1 U6801 ( .A1(n6429), .A2(n5141), .ZN(n5094) );
  NAND2_X2 U6802 ( .A1(n5095), .A2(n5094), .ZN(n9123) );
  NOR2_X2 U6803 ( .A1(n7176), .A2(n9123), .ZN(n6953) );
  OAI21_X1 U6804 ( .B1(n5098), .B2(SI_5_), .A(n5125), .ZN(n5105) );
  NAND3_X1 U6805 ( .A1(n5099), .A2(n5100), .A3(n5105), .ZN(n5107) );
  NAND2_X1 U6806 ( .A1(n5101), .A2(n5100), .ZN(n5120) );
  INV_X1 U6807 ( .A(n5120), .ZN(n5102) );
  NAND2_X1 U6808 ( .A1(n5122), .A2(n5102), .ZN(n5106) );
  INV_X1 U6809 ( .A(n5103), .ZN(n5104) );
  NAND2_X1 U6810 ( .A1(n5106), .A2(n5123), .ZN(n5118) );
  NAND2_X1 U6811 ( .A1(n5107), .A2(n5118), .ZN(n6455) );
  OR2_X1 U6812 ( .A1(n6455), .A2(n5210), .ZN(n5115) );
  NAND2_X1 U6813 ( .A1(n5110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5109) );
  MUX2_X1 U6814 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5109), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5113) );
  INV_X1 U6815 ( .A(n5110), .ZN(n5112) );
  INV_X1 U6816 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6817 ( .A1(n5112), .A2(n5111), .ZN(n5130) );
  NAND2_X1 U6818 ( .A1(n5113), .A2(n5130), .ZN(n6551) );
  INV_X1 U6819 ( .A(n6551), .ZN(n9501) );
  AOI22_X1 U6820 ( .A1(n5423), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6449), .B2(
        n9501), .ZN(n5114) );
  NAND2_X1 U6821 ( .A1(n6953), .A2(n7542), .ZN(n7064) );
  INV_X1 U6822 ( .A(n7064), .ZN(n5133) );
  MUX2_X1 U6823 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5116), .Z(n5117) );
  NAND2_X1 U6824 ( .A1(n5117), .A2(SI_6_), .ZN(n5164) );
  OAI21_X1 U6825 ( .B1(n5117), .B2(SI_6_), .A(n5164), .ZN(n5124) );
  NAND3_X1 U6826 ( .A1(n5118), .A2(n5125), .A3(n5124), .ZN(n5129) );
  INV_X1 U6827 ( .A(n5125), .ZN(n5119) );
  NOR2_X1 U6828 ( .A1(n5120), .A2(n5119), .ZN(n5121) );
  INV_X1 U6829 ( .A(n5123), .ZN(n5126) );
  AOI21_X1 U6830 ( .B1(n5126), .B2(n5125), .A(n5124), .ZN(n5127) );
  NAND2_X1 U6831 ( .A1(n5129), .A2(n5167), .ZN(n6436) );
  OR2_X1 U6832 ( .A1(n6436), .A2(n5210), .ZN(n5132) );
  NAND2_X1 U6833 ( .A1(n5130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5143) );
  XNOR2_X1 U6834 ( .A(n5143), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9514) );
  AOI22_X1 U6835 ( .A1(n5423), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6449), .B2(
        n9514), .ZN(n5131) );
  NAND2_X1 U6836 ( .A1(n5167), .A2(n5164), .ZN(n5139) );
  INV_X1 U6837 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10205) );
  INV_X1 U6838 ( .A(SI_7_), .ZN(n5135) );
  NAND2_X1 U6839 ( .A1(n5136), .A2(n5135), .ZN(n5160) );
  INV_X1 U6840 ( .A(n5136), .ZN(n5137) );
  AND2_X1 U6841 ( .A1(n5160), .A2(n5162), .ZN(n5138) );
  NAND2_X1 U6842 ( .A1(n5139), .A2(n5138), .ZN(n5147) );
  OR2_X1 U6843 ( .A1(n5139), .A2(n5138), .ZN(n5140) );
  INV_X1 U6844 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U6845 ( .A1(n5143), .A2(n5142), .ZN(n5144) );
  NAND2_X1 U6846 ( .A1(n5144), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5145) );
  XNOR2_X1 U6847 ( .A(n5145), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U6848 ( .A1(n5423), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6449), .B2(
        n9527), .ZN(n5146) );
  NAND2_X1 U6849 ( .A1(n5147), .A2(n5162), .ZN(n5152) );
  INV_X1 U6850 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5148) );
  XNOR2_X1 U6851 ( .A(n5152), .B(n5161), .ZN(n6442) );
  NAND2_X1 U6852 ( .A1(n6442), .A2(n5422), .ZN(n5159) );
  NAND3_X1 U6853 ( .A1(n5154), .A2(n5153), .A3(n10223), .ZN(n5156) );
  NAND2_X1 U6854 ( .A1(n5156), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5155) );
  MUX2_X1 U6855 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5155), .S(
        P1_IR_REG_8__SCAN_IN), .Z(n5157) );
  AOI22_X1 U6856 ( .A1(n5423), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6449), .B2(
        n9540), .ZN(n5158) );
  INV_X1 U6857 ( .A(n9857), .ZN(n7244) );
  AND2_X2 U6858 ( .A1(n7230), .A2(n7244), .ZN(n7379) );
  INV_X1 U6859 ( .A(n5160), .ZN(n5166) );
  INV_X1 U6860 ( .A(n5161), .ZN(n5163) );
  OAI211_X1 U6861 ( .C1(n5166), .C2(n5164), .A(n5163), .B(n5162), .ZN(n5165)
         );
  INV_X1 U6862 ( .A(n5168), .ZN(n5169) );
  INV_X1 U6863 ( .A(SI_8_), .ZN(n10204) );
  NAND2_X1 U6864 ( .A1(n5169), .A2(n10204), .ZN(n5170) );
  INV_X1 U6865 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6462) );
  INV_X1 U6866 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6454) );
  XNOR2_X1 U6867 ( .A(n5181), .B(SI_9_), .ZN(n5178) );
  NAND2_X1 U6868 ( .A1(n6453), .A2(n5422), .ZN(n5177) );
  NAND2_X1 U6869 ( .A1(n5173), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5172) );
  MUX2_X1 U6870 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5172), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n5175) );
  INV_X1 U6871 ( .A(n5212), .ZN(n5174) );
  NAND2_X1 U6872 ( .A1(n5175), .A2(n5174), .ZN(n6636) );
  INV_X1 U6873 ( .A(n6636), .ZN(n6564) );
  AOI22_X1 U6874 ( .A1(n5423), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6449), .B2(
        n6564), .ZN(n5176) );
  NAND2_X1 U6875 ( .A1(n5177), .A2(n5176), .ZN(n8830) );
  INV_X1 U6876 ( .A(n8830), .ZN(n9142) );
  INV_X1 U6877 ( .A(SI_9_), .ZN(n5180) );
  NAND2_X1 U6878 ( .A1(n5181), .A2(n5180), .ZN(n5182) );
  NAND2_X1 U6879 ( .A1(n5183), .A2(n5182), .ZN(n5187) );
  MUX2_X1 U6880 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6430), .Z(n5184) );
  NAND2_X1 U6881 ( .A1(n5184), .A2(SI_10_), .ZN(n5195) );
  OAI21_X1 U6882 ( .B1(n5184), .B2(SI_10_), .A(n5195), .ZN(n5186) );
  NAND2_X1 U6883 ( .A1(n5187), .A2(n5186), .ZN(n5188) );
  NAND2_X1 U6884 ( .A1(n5196), .A2(n5188), .ZN(n6465) );
  OR2_X1 U6885 ( .A1(n6465), .A2(n5210), .ZN(n5194) );
  NOR2_X1 U6886 ( .A1(n5212), .A2(n5035), .ZN(n5189) );
  NAND2_X1 U6887 ( .A1(n5189), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5192) );
  INV_X1 U6888 ( .A(n5189), .ZN(n5191) );
  NAND2_X1 U6889 ( .A1(n5191), .A2(n5190), .ZN(n5197) );
  AOI22_X1 U6890 ( .A1(n5423), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6449), .B2(
        n6779), .ZN(n5193) );
  MUX2_X1 U6891 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6430), .Z(n5202) );
  XNOR2_X1 U6892 ( .A(n5202), .B(SI_11_), .ZN(n5203) );
  NAND2_X1 U6893 ( .A1(n6474), .A2(n5422), .ZN(n5200) );
  NAND2_X1 U6894 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  XNOR2_X1 U6895 ( .A(n5198), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9559) );
  AOI22_X1 U6896 ( .A1(n5423), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9559), .B2(
        n6449), .ZN(n5199) );
  OAI21_X1 U6897 ( .B1(n5205), .B2(SI_12_), .A(n5218), .ZN(n5207) );
  NAND2_X1 U6898 ( .A1(n5208), .A2(n5207), .ZN(n5209) );
  NAND2_X1 U6899 ( .A1(n5219), .A2(n5209), .ZN(n6482) );
  OR2_X1 U6900 ( .A1(n6482), .A2(n5210), .ZN(n5217) );
  NOR2_X1 U6901 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5211) );
  NAND2_X1 U6902 ( .A1(n5212), .A2(n5211), .ZN(n5214) );
  NAND2_X1 U6903 ( .A1(n5214), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5213) );
  MUX2_X1 U6904 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5213), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5215) );
  AOI22_X1 U6905 ( .A1(n5423), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6449), .B2(
        n6788), .ZN(n5216) );
  MUX2_X1 U6906 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6430), .Z(n5220) );
  NAND2_X1 U6907 ( .A1(n6489), .A2(n5422), .ZN(n5223) );
  NAND2_X1 U6908 ( .A1(n5229), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6909 ( .A(n5221), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9576) );
  AOI22_X1 U6910 ( .A1(n5423), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n9576), .B2(
        n6449), .ZN(n5222) );
  NAND2_X1 U6911 ( .A1(n9830), .A2(n9837), .ZN(n9816) );
  INV_X1 U6912 ( .A(n5224), .ZN(n5225) );
  MUX2_X1 U6913 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6430), .Z(n5255) );
  XNOR2_X1 U6914 ( .A(n5255), .B(SI_14_), .ZN(n5228) );
  NAND2_X1 U6915 ( .A1(n6593), .A2(n5422), .ZN(n5234) );
  OAI21_X1 U6916 ( .B1(n5229), .B2(P1_IR_REG_13__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5231) );
  INV_X1 U6917 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6918 ( .A1(n5231), .A2(n5230), .ZN(n5238) );
  OR2_X1 U6919 ( .A1(n5231), .A2(n5230), .ZN(n5232) );
  AOI22_X1 U6920 ( .A1(n10006), .A2(n6449), .B1(n5423), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5233) );
  NAND2_X2 U6921 ( .A1(n5234), .A2(n5233), .ZN(n5616) );
  NAND2_X1 U6922 ( .A1(n5253), .A2(SI_14_), .ZN(n5235) );
  XNOR2_X1 U6923 ( .A(n5256), .B(SI_15_), .ZN(n5237) );
  NAND2_X1 U6924 ( .A1(n6727), .A2(n5422), .ZN(n5244) );
  NAND2_X1 U6925 ( .A1(n5238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5240) );
  INV_X1 U6926 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5239) );
  XNOR2_X1 U6927 ( .A(n5240), .B(n5239), .ZN(n10015) );
  INV_X1 U6928 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6730) );
  OAI22_X1 U6929 ( .A1(n10015), .A2(n5241), .B1(n5397), .B2(n6730), .ZN(n5242)
         );
  INV_X1 U6930 ( .A(n5242), .ZN(n5243) );
  NOR2_X4 U6931 ( .A1(n9817), .A2(n9929), .ZN(n9789) );
  NAND2_X1 U6932 ( .A1(n5245), .A2(SI_15_), .ZN(n5246) );
  NAND2_X1 U6933 ( .A1(n5246), .A2(n5258), .ZN(n5247) );
  XNOR2_X1 U6934 ( .A(n5259), .B(SI_16_), .ZN(n5248) );
  NAND2_X1 U6935 ( .A1(n6062), .A2(n5422), .ZN(n5252) );
  NAND2_X1 U6936 ( .A1(n5452), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6937 ( .A(n5250), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10037) );
  AOI22_X1 U6938 ( .A1(n5423), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6449), .B2(
        n10037), .ZN(n5251) );
  NAND2_X2 U6939 ( .A1(n5252), .A2(n5251), .ZN(n9923) );
  INV_X1 U6940 ( .A(n5254), .ZN(n5265) );
  NAND2_X1 U6941 ( .A1(n5255), .A2(SI_14_), .ZN(n5264) );
  NAND3_X1 U6942 ( .A1(n5256), .A2(SI_16_), .A3(SI_15_), .ZN(n5263) );
  OAI21_X1 U6943 ( .B1(n5258), .B2(n10300), .A(n5257), .ZN(n5261) );
  INV_X1 U6944 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U6945 ( .A1(n5261), .A2(n5260), .ZN(n5262) );
  OAI211_X1 U6946 ( .C1(n5265), .C2(n5264), .A(n5263), .B(n5262), .ZN(n5266)
         );
  INV_X1 U6947 ( .A(n5266), .ZN(n5267) );
  INV_X1 U6948 ( .A(SI_17_), .ZN(n5268) );
  INV_X1 U6949 ( .A(n5269), .ZN(n5270) );
  NAND2_X1 U6950 ( .A1(n5270), .A2(SI_17_), .ZN(n5271) );
  NAND2_X1 U6951 ( .A1(n5274), .A2(n5271), .ZN(n5275) );
  XNOR2_X1 U6952 ( .A(n5276), .B(n5275), .ZN(n6723) );
  NAND2_X1 U6953 ( .A1(n6723), .A2(n5422), .ZN(n5273) );
  NAND2_X1 U6954 ( .A1(n5429), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5279) );
  XNOR2_X1 U6955 ( .A(n5279), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10045) );
  AOI22_X1 U6956 ( .A1(n5423), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6449), .B2(
        n10045), .ZN(n5272) );
  INV_X1 U6957 ( .A(n9919), .ZN(n9108) );
  OAI21_X2 U6958 ( .B1(n5276), .B2(n5275), .A(n5274), .ZN(n5291) );
  XNOR2_X1 U6959 ( .A(n5291), .B(n5287), .ZN(n6742) );
  NAND2_X1 U6960 ( .A1(n6742), .A2(n5422), .ZN(n5286) );
  NAND2_X1 U6961 ( .A1(n5279), .A2(n5426), .ZN(n5301) );
  AND2_X1 U6962 ( .A1(n5301), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U6963 ( .A1(n5280), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n5284) );
  INV_X1 U6964 ( .A(n5280), .ZN(n5282) );
  NAND2_X1 U6965 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  AOI22_X1 U6966 ( .A1(n5423), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6449), .B2(
        n10065), .ZN(n5285) );
  INV_X1 U6967 ( .A(n5288), .ZN(n5289) );
  NAND2_X1 U6968 ( .A1(n5289), .A2(SI_18_), .ZN(n5290) );
  MUX2_X1 U6969 ( .A(n7006), .B(n7004), .S(n6430), .Z(n5293) );
  INV_X1 U6970 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U6971 ( .A1(n5294), .A2(SI_19_), .ZN(n5295) );
  NAND2_X1 U6972 ( .A1(n5306), .A2(n5295), .ZN(n5305) );
  XNOR2_X1 U6973 ( .A(n5304), .B(n5305), .ZN(n7003) );
  NAND2_X1 U6974 ( .A1(n7003), .A2(n5422), .ZN(n5303) );
  NAND2_X1 U6975 ( .A1(n5281), .A2(n5427), .ZN(n5300) );
  NAND3_X1 U6976 ( .A1(n5301), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_IR_REG_19__SCAN_IN), .ZN(n5299) );
  NAND2_X1 U6977 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n5296) );
  NAND2_X1 U6978 ( .A1(n5296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5297) );
  OAI21_X1 U6979 ( .B1(n5427), .B2(P1_IR_REG_31__SCAN_IN), .A(n5297), .ZN(
        n5298) );
  INV_X2 U6980 ( .A(n5485), .ZN(n9395) );
  AOI22_X1 U6981 ( .A1(n5423), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9395), .B2(
        n6449), .ZN(n5302) );
  XNOR2_X1 U6982 ( .A(n5319), .B(SI_20_), .ZN(n5307) );
  XNOR2_X1 U6983 ( .A(n5326), .B(n5307), .ZN(n7107) );
  NAND2_X1 U6984 ( .A1(n7107), .A2(n5422), .ZN(n5309) );
  OR2_X1 U6985 ( .A1(n5397), .A2(n7108), .ZN(n5308) );
  INV_X1 U6986 ( .A(SI_20_), .ZN(n5318) );
  OAI21_X1 U6987 ( .B1(n5326), .B2(n5318), .A(n5319), .ZN(n5311) );
  NAND2_X1 U6988 ( .A1(n5326), .A2(n5318), .ZN(n5310) );
  NAND2_X1 U6989 ( .A1(n5311), .A2(n5310), .ZN(n5313) );
  XNOR2_X1 U6990 ( .A(n5316), .B(SI_21_), .ZN(n5312) );
  NAND2_X1 U6991 ( .A1(n6125), .A2(n5422), .ZN(n5315) );
  OR2_X1 U6992 ( .A1(n5397), .A2(n7248), .ZN(n5314) );
  INV_X1 U6993 ( .A(n5319), .ZN(n5321) );
  OAI22_X1 U6994 ( .A1(n5321), .A2(SI_20_), .B1(n5322), .B2(SI_21_), .ZN(n5325) );
  INV_X1 U6995 ( .A(SI_21_), .ZN(n5317) );
  OAI21_X1 U6996 ( .B1(n5319), .B2(n5318), .A(n5317), .ZN(n5323) );
  AND2_X1 U6997 ( .A1(SI_21_), .A2(SI_20_), .ZN(n5320) );
  AOI22_X1 U6998 ( .A1(n5323), .A2(n5322), .B1(n5321), .B2(n5320), .ZN(n5324)
         );
  INV_X1 U6999 ( .A(SI_22_), .ZN(n5327) );
  NAND2_X1 U7000 ( .A1(n5328), .A2(n5327), .ZN(n5333) );
  INV_X1 U7001 ( .A(n5328), .ZN(n5329) );
  NAND2_X1 U7002 ( .A1(n5329), .A2(SI_22_), .ZN(n5330) );
  NAND2_X1 U7003 ( .A1(n5333), .A2(n5330), .ZN(n5334) );
  XNOR2_X1 U7004 ( .A(n5335), .B(n5334), .ZN(n7285) );
  NAND2_X1 U7005 ( .A1(n7285), .A2(n5422), .ZN(n5332) );
  OR2_X1 U7006 ( .A1(n5397), .A2(n7287), .ZN(n5331) );
  MUX2_X1 U7007 ( .A(n7394), .B(n10231), .S(n6430), .Z(n5337) );
  INV_X1 U7008 ( .A(SI_23_), .ZN(n5336) );
  NAND2_X1 U7009 ( .A1(n5337), .A2(n5336), .ZN(n5344) );
  INV_X1 U7010 ( .A(n5337), .ZN(n5338) );
  NAND2_X1 U7011 ( .A1(n5338), .A2(SI_23_), .ZN(n5339) );
  XNOR2_X1 U7012 ( .A(n5343), .B(n5342), .ZN(n7396) );
  NAND2_X1 U7013 ( .A1(n7396), .A2(n5422), .ZN(n5341) );
  OR2_X1 U7014 ( .A1(n5397), .A2(n10231), .ZN(n5340) );
  NAND2_X1 U7015 ( .A1(n5343), .A2(n5342), .ZN(n5345) );
  INV_X1 U7016 ( .A(SI_24_), .ZN(n5346) );
  NAND2_X1 U7017 ( .A1(n5347), .A2(n5346), .ZN(n5354) );
  INV_X1 U7018 ( .A(n5347), .ZN(n5348) );
  NAND2_X1 U7019 ( .A1(n5348), .A2(SI_24_), .ZN(n5349) );
  XNOR2_X1 U7020 ( .A(n5353), .B(n5352), .ZN(n7571) );
  NAND2_X1 U7021 ( .A1(n7571), .A2(n5422), .ZN(n5351) );
  OR2_X1 U7022 ( .A1(n5397), .A2(n7573), .ZN(n5350) );
  INV_X1 U7023 ( .A(SI_25_), .ZN(n5355) );
  NAND2_X1 U7024 ( .A1(n5356), .A2(n5355), .ZN(n5363) );
  INV_X1 U7025 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U7026 ( .A1(n5357), .A2(SI_25_), .ZN(n5358) );
  XNOR2_X1 U7027 ( .A(n5362), .B(n5361), .ZN(n7637) );
  NAND2_X1 U7028 ( .A1(n7637), .A2(n5422), .ZN(n5360) );
  OR2_X1 U7029 ( .A1(n5397), .A2(n7639), .ZN(n5359) );
  AND2_X2 U7030 ( .A1(n9651), .A2(n9955), .ZN(n9623) );
  MUX2_X1 U7031 ( .A(n7669), .B(n7672), .S(n6430), .Z(n5365) );
  INV_X1 U7032 ( .A(SI_26_), .ZN(n5364) );
  NAND2_X1 U7033 ( .A1(n5365), .A2(n5364), .ZN(n5372) );
  INV_X1 U7034 ( .A(n5365), .ZN(n5366) );
  NAND2_X1 U7035 ( .A1(n5366), .A2(SI_26_), .ZN(n5367) );
  XNOR2_X1 U7036 ( .A(n5371), .B(n5370), .ZN(n7668) );
  NAND2_X1 U7037 ( .A1(n7668), .A2(n5422), .ZN(n5369) );
  OR2_X1 U7038 ( .A1(n5397), .A2(n7672), .ZN(n5368) );
  AND2_X2 U7039 ( .A1(n9623), .A2(n9625), .ZN(n6318) );
  NAND2_X1 U7040 ( .A1(n5371), .A2(n5370), .ZN(n5373) );
  INV_X1 U7041 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7717) );
  INV_X1 U7042 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7709) );
  INV_X1 U7043 ( .A(SI_27_), .ZN(n5374) );
  NAND2_X1 U7044 ( .A1(n5375), .A2(n5374), .ZN(n5393) );
  INV_X1 U7045 ( .A(n5375), .ZN(n5376) );
  NAND2_X1 U7046 ( .A1(n5376), .A2(SI_27_), .ZN(n5377) );
  NAND2_X1 U7047 ( .A1(n7707), .A2(n5422), .ZN(n5379) );
  OR2_X1 U7048 ( .A1(n5397), .A2(n7709), .ZN(n5378) );
  INV_X1 U7049 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5838) );
  INV_X1 U7050 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7762) );
  XNOR2_X1 U7051 ( .A(n5392), .B(SI_28_), .ZN(n5400) );
  NAND2_X1 U7052 ( .A1(n7761), .A2(n5422), .ZN(n5383) );
  OR2_X1 U7053 ( .A1(n5397), .A2(n7762), .ZN(n5382) );
  INV_X1 U7054 ( .A(n5392), .ZN(n5385) );
  NAND2_X1 U7055 ( .A1(n5385), .A2(SI_28_), .ZN(n5384) );
  MUX2_X1 U7056 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6430), .Z(n5403) );
  INV_X1 U7057 ( .A(n5403), .ZN(n5386) );
  NAND2_X1 U7058 ( .A1(n5384), .A2(n5386), .ZN(n5395) );
  INV_X1 U7059 ( .A(n5395), .ZN(n5390) );
  INV_X1 U7060 ( .A(n5393), .ZN(n5389) );
  INV_X1 U7061 ( .A(SI_28_), .ZN(n5391) );
  OAI21_X1 U7062 ( .B1(n5386), .B2(n5391), .A(n5385), .ZN(n5388) );
  OAI21_X1 U7063 ( .B1(n5403), .B2(SI_28_), .A(n5392), .ZN(n5387) );
  AOI22_X1 U7064 ( .A1(n5390), .A2(n5389), .B1(n5388), .B2(n5387), .ZN(n5394)
         );
  NAND2_X1 U7065 ( .A1(n5392), .A2(n5391), .ZN(n5402) );
  NAND2_X1 U7066 ( .A1(n8815), .A2(n5422), .ZN(n5399) );
  INV_X1 U7067 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9996) );
  OR2_X1 U7068 ( .A1(n5397), .A2(n9996), .ZN(n5398) );
  INV_X1 U7069 ( .A(SI_29_), .ZN(n5407) );
  NAND2_X1 U7070 ( .A1(n5401), .A2(n5400), .ZN(n5404) );
  NAND3_X1 U7071 ( .A1(n5404), .A2(n5403), .A3(n5402), .ZN(n5405) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8019) );
  INV_X1 U7073 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n5408) );
  MUX2_X1 U7074 ( .A(n8019), .B(n5408), .S(n6430), .Z(n5410) );
  INV_X1 U7075 ( .A(SI_30_), .ZN(n5409) );
  NAND2_X1 U7076 ( .A1(n5410), .A2(n5409), .ZN(n5415) );
  INV_X1 U7077 ( .A(n5410), .ZN(n5411) );
  NAND2_X1 U7078 ( .A1(n5411), .A2(SI_30_), .ZN(n5412) );
  NAND2_X1 U7079 ( .A1(n5415), .A2(n5412), .ZN(n5416) );
  XNOR2_X1 U7080 ( .A(n5417), .B(n5416), .ZN(n8018) );
  NAND2_X1 U7081 ( .A1(n8018), .A2(n5422), .ZN(n5414) );
  NAND2_X1 U7082 ( .A1(n5423), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5413) );
  INV_X1 U7083 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8028) );
  INV_X1 U7084 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5418) );
  XNOR2_X1 U7085 ( .A(n5419), .B(SI_31_), .ZN(n5420) );
  NAND2_X1 U7086 ( .A1(n8809), .A2(n5422), .ZN(n5425) );
  NAND2_X1 U7087 ( .A1(n5423), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5424) );
  XNOR2_X1 U7088 ( .A(n9601), .B(n9600), .ZN(n5437) );
  NAND3_X1 U7089 ( .A1(n5281), .A2(n5427), .A3(n5426), .ZN(n5428) );
  INV_X1 U7090 ( .A(n5458), .ZN(n5431) );
  INV_X1 U7091 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U7092 ( .A1(n6514), .A2(P1_B_REG_SCAN_IN), .ZN(n5438) );
  NAND2_X1 U7093 ( .A1(n9843), .A2(n5438), .ZN(n5787) );
  INV_X1 U7094 ( .A(n5787), .ZN(n5449) );
  NAND2_X1 U7095 ( .A1(n5442), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5440) );
  NAND2_X2 U7096 ( .A1(n5441), .A2(n9986), .ZN(n9997) );
  NAND2_X1 U7097 ( .A1(n5781), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U7098 ( .A1(n5782), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n5447) );
  AND2_X2 U7099 ( .A1(n5445), .A2(n9997), .ZN(n5513) );
  NAND2_X1 U7100 ( .A1(n5732), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5446) );
  NAND3_X1 U7101 ( .A1(n5448), .A2(n5447), .A3(n5446), .ZN(n9376) );
  NOR2_X1 U7102 ( .A1(n9596), .A2(n9864), .ZN(n5805) );
  NAND3_X1 U7103 ( .A1(n5460), .A2(n5453), .A3(n5469), .ZN(n5457) );
  XNOR2_X1 U7104 ( .A(n5454), .B(P1_IR_REG_31__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U7105 ( .A1(n5460), .A2(n5455), .ZN(n5456) );
  NAND2_X1 U7106 ( .A1(n5460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5459) );
  MUX2_X1 U7107 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5459), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5461) );
  NAND2_X1 U7108 ( .A1(n4321), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5462) );
  INV_X1 U7109 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7110 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  NAND2_X1 U7111 ( .A1(n5468), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7112 ( .A1(n7641), .A2(P1_B_REG_SCAN_IN), .ZN(n5473) );
  MUX2_X1 U7113 ( .A(n5473), .B(P1_B_REG_SCAN_IN), .S(n5491), .Z(n5474) );
  NOR2_X1 U7114 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n5478) );
  NOR4_X1 U7115 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5477) );
  NOR4_X1 U7116 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5476) );
  NOR4_X1 U7117 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5475) );
  NAND4_X1 U7118 ( .A1(n5478), .A2(n5477), .A3(n5476), .A4(n5475), .ZN(n5484)
         );
  NOR4_X1 U7119 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5482) );
  NOR4_X1 U7120 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5481) );
  NOR4_X1 U7121 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5480) );
  NOR4_X1 U7122 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5479) );
  NAND4_X1 U7123 ( .A1(n5482), .A2(n5481), .A3(n5480), .A4(n5479), .ZN(n5483)
         );
  NOR2_X1 U7124 ( .A1(n5484), .A2(n5483), .ZN(n6675) );
  NAND2_X1 U7125 ( .A1(n6448), .A2(n6675), .ZN(n5486) );
  NAND2_X1 U7126 ( .A1(n9782), .A2(n9395), .ZN(n5750) );
  NAND2_X1 U7127 ( .A1(n7674), .A2(n7641), .ZN(n9984) );
  OAI21_X1 U7128 ( .B1(n6674), .B2(P1_D_REG_1__SCAN_IN), .A(n9984), .ZN(n5748)
         );
  AND2_X1 U7129 ( .A1(n5750), .A2(n5748), .ZN(n5488) );
  INV_X1 U7130 ( .A(n6674), .ZN(n5490) );
  INV_X1 U7131 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5489) );
  NAND2_X1 U7132 ( .A1(n5490), .A2(n5489), .ZN(n5492) );
  INV_X1 U7133 ( .A(n5491), .ZN(n7572) );
  NAND2_X1 U7134 ( .A1(n7674), .A2(n7572), .ZN(n9985) );
  OR2_X1 U7135 ( .A1(n5805), .A2(n10118), .ZN(n5496) );
  INV_X1 U7136 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U7137 ( .A1(n5496), .A2(n5495), .ZN(P1_U3553) );
  INV_X1 U7138 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7139 ( .A1(n5512), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5500) );
  NAND2_X1 U7140 ( .A1(n5513), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5499) );
  NAND3_X1 U7141 ( .A1(n5504), .A2(n9991), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n5498) );
  NAND4_X1 U7142 ( .A1(n5500), .A2(n5501), .A3(n5499), .A4(n5498), .ZN(n5502)
         );
  NAND2_X1 U7143 ( .A1(n5502), .A2(n6684), .ZN(n9401) );
  NAND2_X1 U7144 ( .A1(n5528), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7145 ( .A1(n5512), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U7146 ( .A1(n5513), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U7147 ( .A1(n9474), .A2(n10090), .ZN(n7256) );
  NAND2_X1 U7148 ( .A1(n5509), .A2(n10101), .ZN(n5510) );
  NAND2_X1 U7149 ( .A1(n7255), .A2(n5510), .ZN(n6791) );
  NAND2_X1 U7150 ( .A1(n5528), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7151 ( .A1(n5512), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5515) );
  NAND2_X1 U7152 ( .A1(n5513), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5514) );
  NAND2_X1 U7153 ( .A1(n6801), .A2(n9472), .ZN(n9404) );
  NAND2_X1 U7154 ( .A1(n5518), .A2(n10073), .ZN(n5761) );
  NAND2_X1 U7155 ( .A1(n9404), .A2(n5761), .ZN(n9242) );
  NAND2_X1 U7156 ( .A1(n6791), .A2(n9242), .ZN(n6793) );
  NAND2_X1 U7157 ( .A1(n5518), .A2(n6801), .ZN(n5519) );
  NAND2_X1 U7158 ( .A1(n6793), .A2(n5519), .ZN(n6949) );
  NAND2_X1 U7159 ( .A1(n5782), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5523) );
  INV_X1 U7160 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6739) );
  NAND2_X1 U7161 ( .A1(n5738), .A2(n6739), .ZN(n5522) );
  NAND2_X1 U7162 ( .A1(n5618), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7163 ( .A1(n5732), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7164 ( .A1(n6956), .A2(n7181), .ZN(n9279) );
  NAND2_X1 U7165 ( .A1(n5618), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5533) );
  NAND2_X1 U7166 ( .A1(n5732), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5532) );
  INV_X1 U7167 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n5524) );
  OR2_X1 U7168 ( .A1(n5525), .A2(n5524), .ZN(n5530) );
  INV_X1 U7169 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5526) );
  NAND2_X1 U7170 ( .A1(n6739), .A2(n5526), .ZN(n5527) );
  AND2_X1 U7171 ( .A1(n5527), .A2(n5539), .ZN(n9122) );
  NAND2_X1 U7172 ( .A1(n5528), .A2(n9122), .ZN(n5529) );
  INV_X1 U7173 ( .A(n9123), .ZN(n7330) );
  NAND3_X1 U7174 ( .A1(n6949), .A2(n6950), .A3(n5763), .ZN(n5536) );
  NOR2_X1 U7175 ( .A1(n9471), .A2(n7181), .ZN(n6951) );
  NOR2_X1 U7176 ( .A1(n9123), .A2(n9470), .ZN(n5534) );
  AOI21_X1 U7177 ( .B1(n6951), .B2(n5763), .A(n5534), .ZN(n5535) );
  NAND2_X1 U7178 ( .A1(n5536), .A2(n5535), .ZN(n6904) );
  NAND2_X1 U7179 ( .A1(n5513), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7180 ( .A1(n5618), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5543) );
  INV_X1 U7181 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7182 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AND2_X1 U7183 ( .A1(n5556), .A2(n5540), .ZN(n7539) );
  NAND2_X1 U7184 ( .A1(n5738), .A2(n7539), .ZN(n5542) );
  NAND2_X1 U7185 ( .A1(n5782), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7186 ( .A1(n7542), .A2(n9469), .ZN(n9406) );
  INV_X1 U7187 ( .A(n9469), .ZN(n7051) );
  NAND2_X1 U7188 ( .A1(n7054), .A2(n7051), .ZN(n9286) );
  NAND2_X1 U7189 ( .A1(n9406), .A2(n9286), .ZN(n9243) );
  NAND2_X1 U7190 ( .A1(n6904), .A2(n9243), .ZN(n6905) );
  NAND2_X1 U7191 ( .A1(n7542), .A2(n7051), .ZN(n5545) );
  NAND2_X1 U7192 ( .A1(n5782), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5550) );
  XNOR2_X1 U7193 ( .A(n5556), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n7340) );
  NAND2_X1 U7194 ( .A1(n5738), .A2(n7340), .ZN(n5549) );
  INV_X2 U7195 ( .A(n5546), .ZN(n5618) );
  NAND2_X1 U7196 ( .A1(n5618), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U7197 ( .A1(n5732), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5547) );
  NAND4_X1 U7198 ( .A1(n5550), .A2(n5549), .A3(n5548), .A4(n5547), .ZN(n9468)
         );
  NAND2_X1 U7199 ( .A1(n7339), .A2(n9468), .ZN(n9276) );
  INV_X1 U7200 ( .A(n9468), .ZN(n7212) );
  NAND2_X1 U7201 ( .A1(n7212), .A2(n7317), .ZN(n9284) );
  NAND2_X1 U7202 ( .A1(n9276), .A2(n9284), .ZN(n7199) );
  NAND2_X1 U7203 ( .A1(n7339), .A2(n7212), .ZN(n5551) );
  INV_X1 U7204 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5555) );
  INV_X1 U7205 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5554) );
  OAI21_X1 U7206 ( .B1(n5556), .B2(n5555), .A(n5554), .ZN(n5557) );
  AND2_X1 U7207 ( .A1(n5563), .A2(n5557), .ZN(n7529) );
  NAND2_X1 U7208 ( .A1(n5738), .A2(n7529), .ZN(n5560) );
  NAND2_X1 U7209 ( .A1(n5618), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7210 ( .A1(n5782), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U7211 ( .A1(n7532), .A2(n7218), .ZN(n5561) );
  NAND2_X1 U7212 ( .A1(n5782), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7213 ( .A1(n5732), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5567) );
  INV_X1 U7214 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10273) );
  NAND2_X1 U7215 ( .A1(n5563), .A2(n10273), .ZN(n5564) );
  AND2_X1 U7216 ( .A1(n5571), .A2(n5564), .ZN(n7587) );
  NAND2_X1 U7217 ( .A1(n5738), .A2(n7587), .ZN(n5566) );
  NAND2_X1 U7218 ( .A1(n5618), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5565) );
  OR2_X1 U7219 ( .A1(n9857), .A2(n9137), .ZN(n7381) );
  NAND2_X1 U7220 ( .A1(n9857), .A2(n9137), .ZN(n9294) );
  NAND2_X1 U7221 ( .A1(n7381), .A2(n9294), .ZN(n7236) );
  INV_X1 U7222 ( .A(n9137), .ZN(n9466) );
  OR2_X1 U7223 ( .A1(n9857), .A2(n9466), .ZN(n5569) );
  NAND2_X1 U7224 ( .A1(n5782), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5576) );
  NAND2_X1 U7225 ( .A1(n5732), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U7226 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  AND2_X1 U7227 ( .A1(n5579), .A2(n5572), .ZN(n9135) );
  NAND2_X1 U7228 ( .A1(n5738), .A2(n9135), .ZN(n5574) );
  NAND2_X1 U7229 ( .A1(n5618), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7230 ( .A1(n8830), .A2(n8828), .ZN(n9302) );
  NAND2_X1 U7231 ( .A1(n9316), .A2(n9302), .ZN(n7384) );
  INV_X1 U7232 ( .A(n8828), .ZN(n9465) );
  NAND2_X1 U7233 ( .A1(n5782), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7234 ( .A1(n5732), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5583) );
  INV_X1 U7235 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U7236 ( .A1(n5579), .A2(n5578), .ZN(n5580) );
  AND2_X1 U7237 ( .A1(n5587), .A2(n5580), .ZN(n9014) );
  NAND2_X1 U7238 ( .A1(n5738), .A2(n9014), .ZN(n5582) );
  NAND2_X1 U7239 ( .A1(n5618), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5581) );
  OR2_X1 U7240 ( .A1(n9019), .A2(n9178), .ZN(n9409) );
  NAND2_X1 U7241 ( .A1(n9019), .A2(n9178), .ZN(n9303) );
  NAND2_X1 U7242 ( .A1(n9409), .A2(n9303), .ZN(n9250) );
  NAND2_X1 U7243 ( .A1(n7276), .A2(n9250), .ZN(n7277) );
  OR2_X1 U7244 ( .A1(n9019), .A2(n9464), .ZN(n5585) );
  NAND2_X1 U7245 ( .A1(n5732), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7246 ( .A1(n5782), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5591) );
  NAND2_X1 U7247 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  AND2_X1 U7248 ( .A1(n5595), .A2(n5588), .ZN(n7442) );
  NAND2_X1 U7249 ( .A1(n5738), .A2(n7442), .ZN(n5590) );
  NAND2_X1 U7250 ( .A1(n5618), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5589) );
  OR2_X1 U7251 ( .A1(n8845), .A2(n9072), .ZN(n9318) );
  NAND2_X1 U7252 ( .A1(n8845), .A2(n9072), .ZN(n9319) );
  NAND2_X1 U7253 ( .A1(n9318), .A2(n9319), .ZN(n9241) );
  INV_X1 U7254 ( .A(n9072), .ZN(n9463) );
  OR2_X1 U7255 ( .A1(n8845), .A2(n9463), .ZN(n5593) );
  NAND2_X1 U7256 ( .A1(n5732), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7257 ( .A1(n5618), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5599) );
  INV_X1 U7258 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7259 ( .A1(n5595), .A2(n5594), .ZN(n5596) );
  AND2_X1 U7260 ( .A1(n5603), .A2(n5596), .ZN(n9070) );
  NAND2_X1 U7261 ( .A1(n5738), .A2(n9070), .ZN(n5598) );
  NAND2_X1 U7262 ( .A1(n5782), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5597) );
  OR2_X1 U7263 ( .A1(n8856), .A2(n9157), .ZN(n9322) );
  NAND2_X1 U7264 ( .A1(n8856), .A2(n9157), .ZN(n9416) );
  INV_X1 U7265 ( .A(n9157), .ZN(n9842) );
  OR2_X1 U7266 ( .A1(n8856), .A2(n9842), .ZN(n5601) );
  NAND2_X1 U7267 ( .A1(n5513), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7268 ( .A1(n5782), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5607) );
  NAND2_X1 U7269 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  AND2_X1 U7270 ( .A1(n5610), .A2(n5604), .ZN(n9834) );
  NAND2_X1 U7271 ( .A1(n5738), .A2(n9834), .ZN(n5606) );
  NAND2_X1 U7272 ( .A1(n5618), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5605) );
  OR2_X1 U7273 ( .A1(n9939), .A2(n9809), .ZN(n9419) );
  NAND2_X1 U7274 ( .A1(n9939), .A2(n9809), .ZN(n9417) );
  NAND2_X1 U7275 ( .A1(n9419), .A2(n9417), .ZN(n9827) );
  INV_X1 U7276 ( .A(n9809), .ZN(n9075) );
  NAND2_X1 U7277 ( .A1(n5610), .A2(n5609), .ZN(n5611) );
  AND2_X1 U7278 ( .A1(n5620), .A2(n5611), .ZN(n9819) );
  NAND2_X1 U7279 ( .A1(n9819), .A2(n5738), .ZN(n5615) );
  NAND2_X1 U7280 ( .A1(n5732), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7281 ( .A1(n5781), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7282 ( .A1(n5782), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7283 ( .A1(n5616), .A2(n9211), .ZN(n9326) );
  NAND2_X1 U7284 ( .A1(n9802), .A2(n9804), .ZN(n9803) );
  INV_X1 U7285 ( .A(n9211), .ZN(n9844) );
  OR2_X1 U7286 ( .A1(n5616), .A2(n9844), .ZN(n5617) );
  INV_X1 U7287 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10017) );
  INV_X1 U7288 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U7289 ( .A1(n5620), .A2(n5619), .ZN(n5621) );
  NAND2_X1 U7290 ( .A1(n5629), .A2(n5621), .ZN(n9790) );
  OR2_X1 U7291 ( .A1(n9790), .A2(n5725), .ZN(n5625) );
  NAND2_X1 U7292 ( .A1(n5782), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U7293 ( .A1(n5513), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5622) );
  AND2_X1 U7294 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  OAI211_X1 U7295 ( .C1(n5546), .C2(n10017), .A(n5625), .B(n5624), .ZN(n9773)
         );
  NAND2_X1 U7296 ( .A1(n9929), .A2(n9773), .ZN(n5626) );
  INV_X1 U7297 ( .A(n5629), .ZN(n5627) );
  INV_X1 U7298 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7299 ( .A1(n5629), .A2(n5628), .ZN(n5630) );
  NAND2_X1 U7300 ( .A1(n5645), .A2(n5630), .ZN(n9780) );
  OR2_X1 U7301 ( .A1(n9780), .A2(n5725), .ZN(n5633) );
  AOI22_X1 U7302 ( .A1(n5782), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n5513), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U7303 ( .A1(n5781), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5631) );
  OR2_X1 U7304 ( .A1(n9923), .A2(n9764), .ZN(n9421) );
  NAND2_X1 U7305 ( .A1(n9923), .A2(n9764), .ZN(n9758) );
  OR2_X1 U7306 ( .A1(n9929), .A2(n9773), .ZN(n9776) );
  INV_X1 U7307 ( .A(n9764), .ZN(n9797) );
  NAND2_X1 U7308 ( .A1(n9923), .A2(n9797), .ZN(n5636) );
  XNOR2_X1 U7309 ( .A(n5645), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9103) );
  NAND2_X1 U7310 ( .A1(n9103), .A2(n5738), .ZN(n5641) );
  INV_X1 U7311 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10312) );
  NAND2_X1 U7312 ( .A1(n5513), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7313 ( .A1(n5781), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U7314 ( .C1(n5736), .C2(n10312), .A(n5638), .B(n5637), .ZN(n5639)
         );
  INV_X1 U7315 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7316 ( .A1(n5641), .A2(n5640), .ZN(n9772) );
  OR2_X1 U7317 ( .A1(n9919), .A2(n9772), .ZN(n5642) );
  INV_X1 U7318 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5643) );
  INV_X1 U7319 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9186) );
  OAI21_X1 U7320 ( .B1(n5645), .B2(n5643), .A(n9186), .ZN(n5646) );
  NAND2_X1 U7321 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_REG3_REG_18__SCAN_IN), 
        .ZN(n5644) );
  AND2_X1 U7322 ( .A1(n5646), .A2(n5655), .ZN(n9748) );
  NAND2_X1 U7323 ( .A1(n9748), .A2(n5738), .ZN(n5652) );
  INV_X1 U7324 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7325 ( .A1(n5732), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7326 ( .A1(n5781), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5647) );
  OAI211_X1 U7327 ( .C1(n5736), .C2(n5649), .A(n5648), .B(n5647), .ZN(n5650)
         );
  INV_X1 U7328 ( .A(n5650), .ZN(n5651) );
  NAND2_X1 U7329 ( .A1(n5652), .A2(n5651), .ZN(n9730) );
  NAND2_X1 U7330 ( .A1(n9747), .A2(n9730), .ZN(n5653) );
  NAND2_X1 U7331 ( .A1(n5654), .A2(n5653), .ZN(n9722) );
  INV_X1 U7332 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U7333 ( .A1(n5655), .A2(n10261), .ZN(n5656) );
  NAND2_X1 U7334 ( .A1(n5663), .A2(n5656), .ZN(n9724) );
  OR2_X1 U7335 ( .A1(n9724), .A2(n5725), .ZN(n5661) );
  INV_X1 U7336 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U7337 ( .A1(n5782), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5658) );
  NAND2_X1 U7338 ( .A1(n5781), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5657) );
  OAI211_X1 U7339 ( .C1(n5742), .C2(n10315), .A(n5658), .B(n5657), .ZN(n5659)
         );
  INV_X1 U7340 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7341 ( .A1(n5661), .A2(n5660), .ZN(n9462) );
  OR2_X1 U7342 ( .A1(n9908), .A2(n9462), .ZN(n5662) );
  INV_X1 U7343 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9148) );
  NAND2_X1 U7344 ( .A1(n5663), .A2(n9148), .ZN(n5664) );
  AND2_X1 U7345 ( .A1(n5670), .A2(n5664), .ZN(n9715) );
  INV_X1 U7346 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n5667) );
  NAND2_X1 U7347 ( .A1(n5781), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U7348 ( .A1(n5732), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5665) );
  OAI211_X1 U7349 ( .C1(n5736), .C2(n5667), .A(n5666), .B(n5665), .ZN(n5668)
         );
  AOI21_X1 U7350 ( .B1(n9715), .B2(n5738), .A(n5668), .ZN(n9056) );
  OR2_X1 U7351 ( .A1(n9903), .A2(n9056), .ZN(n9701) );
  NAND2_X1 U7352 ( .A1(n9903), .A2(n9056), .ZN(n9700) );
  INV_X1 U7353 ( .A(n5670), .ZN(n5669) );
  INV_X1 U7354 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U7355 ( .A1(n5670), .A2(n10233), .ZN(n5671) );
  NAND2_X1 U7356 ( .A1(n5678), .A2(n5671), .ZN(n9694) );
  OR2_X1 U7357 ( .A1(n9694), .A2(n5725), .ZN(n5676) );
  INV_X1 U7358 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U7359 ( .A1(n5781), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7360 ( .A1(n5732), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5672) );
  OAI211_X1 U7361 ( .C1(n5736), .C2(n9693), .A(n5673), .B(n5672), .ZN(n5674)
         );
  INV_X1 U7362 ( .A(n5674), .ZN(n5675) );
  NAND2_X1 U7363 ( .A1(n5676), .A2(n5675), .ZN(n9461) );
  NAND2_X1 U7364 ( .A1(n9968), .A2(n9461), .ZN(n9677) );
  INV_X1 U7365 ( .A(n9056), .ZN(n9731) );
  NAND2_X1 U7366 ( .A1(n9903), .A2(n9731), .ZN(n9676) );
  INV_X1 U7367 ( .A(n9461), .ZN(n8917) );
  NAND2_X1 U7368 ( .A1(n9968), .A2(n8917), .ZN(n9345) );
  INV_X1 U7369 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7370 ( .A1(n5678), .A2(n5677), .ZN(n5679) );
  AND2_X1 U7371 ( .A1(n5688), .A2(n5679), .ZN(n9685) );
  INV_X1 U7372 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7373 ( .A1(n5732), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U7374 ( .A1(n5781), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5680) );
  OAI211_X1 U7375 ( .C1(n5682), .C2(n5736), .A(n5681), .B(n5680), .ZN(n5683)
         );
  AOI22_X1 U7376 ( .A1(n9239), .A2(n9677), .B1(n9965), .B2(n9055), .ZN(n5684)
         );
  INV_X1 U7377 ( .A(n9055), .ZN(n9460) );
  NAND2_X1 U7378 ( .A1(n9683), .A2(n9460), .ZN(n5686) );
  INV_X1 U7379 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5687) );
  NAND2_X1 U7380 ( .A1(n5688), .A2(n5687), .ZN(n5689) );
  INV_X1 U7381 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U7382 ( .A1(n5781), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n5691) );
  NAND2_X1 U7383 ( .A1(n5732), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5690) );
  OAI211_X1 U7384 ( .C1(n5736), .C2(n9668), .A(n5691), .B(n5690), .ZN(n5692)
         );
  INV_X1 U7385 ( .A(n5692), .ZN(n5693) );
  OR2_X1 U7386 ( .A1(n9667), .A2(n9459), .ZN(n5695) );
  XNOR2_X1 U7387 ( .A(n5705), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9653) );
  NAND2_X1 U7388 ( .A1(n9653), .A2(n5738), .ZN(n5700) );
  INV_X1 U7389 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10317) );
  NAND2_X1 U7390 ( .A1(n5781), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5697) );
  NAND2_X1 U7391 ( .A1(n5782), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U7392 ( .C1(n5742), .C2(n10317), .A(n5697), .B(n5696), .ZN(n5698)
         );
  INV_X1 U7393 ( .A(n5698), .ZN(n5699) );
  NAND2_X1 U7394 ( .A1(n9652), .A2(n9458), .ZN(n5701) );
  NAND2_X1 U7395 ( .A1(n5702), .A2(n5701), .ZN(n9634) );
  INV_X1 U7396 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5703) );
  INV_X1 U7397 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9082) );
  OAI21_X1 U7398 ( .B1(n5705), .B2(n5703), .A(n9082), .ZN(n5706) );
  NAND2_X1 U7399 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5704) );
  NAND2_X1 U7400 ( .A1(n5706), .A2(n5715), .ZN(n9639) );
  INV_X1 U7401 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U7402 ( .A1(n5781), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U7403 ( .A1(n5732), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5707) );
  OAI211_X1 U7404 ( .C1(n5736), .C2(n9638), .A(n5708), .B(n5707), .ZN(n5709)
         );
  INV_X1 U7405 ( .A(n5709), .ZN(n5710) );
  AND2_X1 U7406 ( .A1(n9637), .A2(n9457), .ZN(n5712) );
  OR2_X1 U7407 ( .A1(n9637), .A2(n9457), .ZN(n5713) );
  INV_X1 U7408 ( .A(n5715), .ZN(n5714) );
  INV_X1 U7409 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9200) );
  NAND2_X1 U7410 ( .A1(n5715), .A2(n9200), .ZN(n5716) );
  NAND2_X1 U7411 ( .A1(n5723), .A2(n5716), .ZN(n9622) );
  INV_X1 U7412 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9621) );
  NAND2_X1 U7413 ( .A1(n5732), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5718) );
  NAND2_X1 U7414 ( .A1(n5781), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5717) );
  OAI211_X1 U7415 ( .C1(n9621), .C2(n5736), .A(n5718), .B(n5717), .ZN(n5719)
         );
  INV_X1 U7416 ( .A(n5719), .ZN(n5720) );
  NAND2_X2 U7417 ( .A1(n5721), .A2(n5720), .ZN(n9456) );
  NAND2_X1 U7418 ( .A1(n9950), .A2(n9456), .ZN(n5722) );
  INV_X1 U7419 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U7420 ( .A1(n5723), .A2(n8978), .ZN(n5724) );
  NAND2_X1 U7421 ( .A1(n5793), .A2(n5724), .ZN(n9609) );
  INV_X1 U7422 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U7423 ( .A1(n5732), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7424 ( .A1(n5782), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5726) );
  OAI211_X1 U7425 ( .C1(n9868), .C2(n5546), .A(n5727), .B(n5726), .ZN(n5728)
         );
  INV_X1 U7426 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U7427 ( .A1(n8981), .A2(n9199), .ZN(n9357) );
  AND2_X2 U7428 ( .A1(n9358), .A2(n9357), .ZN(n9259) );
  OR2_X1 U7429 ( .A1(n8981), .A2(n9455), .ZN(n5731) );
  XNOR2_X1 U7430 ( .A(n5793), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9041) );
  INV_X1 U7431 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7432 ( .A1(n5781), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5734) );
  NAND2_X1 U7433 ( .A1(n5732), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5733) );
  OAI211_X1 U7434 ( .C1(n5736), .C2(n5735), .A(n5734), .B(n5733), .ZN(n5737)
         );
  NAND2_X1 U7435 ( .A1(n9045), .A2(n9031), .ZN(n9359) );
  INV_X1 U7436 ( .A(n9031), .ZN(n9454) );
  NAND2_X1 U7437 ( .A1(n9045), .A2(n9454), .ZN(n6377) );
  NAND2_X1 U7438 ( .A1(n6381), .A2(n6377), .ZN(n5747) );
  NAND2_X1 U7439 ( .A1(n5738), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5739) );
  OR2_X1 U7440 ( .A1(n5793), .A2(n5739), .ZN(n5745) );
  INV_X1 U7441 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10311) );
  NAND2_X1 U7442 ( .A1(n5782), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5741) );
  NAND2_X1 U7443 ( .A1(n5781), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5740) );
  OAI211_X1 U7444 ( .C1(n5742), .C2(n10311), .A(n5741), .B(n5740), .ZN(n5743)
         );
  INV_X1 U7445 ( .A(n5743), .ZN(n5744) );
  NAND2_X1 U7446 ( .A1(n5746), .A2(n7022), .ZN(n9377) );
  XNOR2_X1 U7447 ( .A(n5747), .B(n4502), .ZN(n5759) );
  INV_X1 U7448 ( .A(n5748), .ZN(n6673) );
  NAND2_X1 U7449 ( .A1(n5749), .A2(n6673), .ZN(n5796) );
  INV_X1 U7450 ( .A(n5750), .ZN(n5751) );
  NAND2_X1 U7451 ( .A1(n5753), .A2(n9765), .ZN(n6687) );
  NAND2_X1 U7452 ( .A1(n6687), .A2(n9443), .ZN(n5754) );
  INV_X1 U7453 ( .A(n10089), .ZN(n10085) );
  AND2_X1 U7454 ( .A1(n5754), .A2(n10085), .ZN(n5756) );
  INV_X1 U7455 ( .A(n6687), .ZN(n5755) );
  NAND2_X1 U7456 ( .A1(n5755), .A2(n6491), .ZN(n10086) );
  NAND2_X1 U7457 ( .A1(n5756), .A2(n10086), .ZN(n9815) );
  INV_X1 U7458 ( .A(n10088), .ZN(n5757) );
  NAND2_X1 U7459 ( .A1(n5757), .A2(n4300), .ZN(n7260) );
  NAND2_X1 U7460 ( .A1(n9815), .A2(n7260), .ZN(n5758) );
  NAND2_X1 U7461 ( .A1(n5759), .A2(n10071), .ZN(n5802) );
  NAND2_X1 U7462 ( .A1(n4291), .A2(n10090), .ZN(n7254) );
  INV_X1 U7463 ( .A(n5761), .ZN(n5762) );
  INV_X1 U7464 ( .A(n9402), .ZN(n9281) );
  NOR2_X1 U7465 ( .A1(n5763), .A2(n9281), .ZN(n5764) );
  INV_X1 U7466 ( .A(n9280), .ZN(n5765) );
  NOR2_X1 U7467 ( .A1(n9243), .A2(n5765), .ZN(n5766) );
  NAND2_X1 U7468 ( .A1(n6907), .A2(n9406), .ZN(n7065) );
  AND2_X1 U7469 ( .A1(n9316), .A2(n7381), .ZN(n9298) );
  NAND2_X1 U7470 ( .A1(n9294), .A2(n7233), .ZN(n9293) );
  INV_X1 U7471 ( .A(n9302), .ZN(n9296) );
  NAND2_X1 U7472 ( .A1(n7381), .A2(n5767), .ZN(n9292) );
  INV_X1 U7473 ( .A(n9316), .ZN(n5768) );
  INV_X1 U7474 ( .A(n9276), .ZN(n9278) );
  INV_X1 U7475 ( .A(n9303), .ZN(n9315) );
  NOR2_X1 U7476 ( .A1(n9241), .A2(n9315), .ZN(n5771) );
  NAND2_X1 U7477 ( .A1(n7278), .A2(n5771), .ZN(n5772) );
  INV_X1 U7478 ( .A(n9827), .ZN(n9840) );
  INV_X1 U7479 ( .A(n9773), .ZN(n9811) );
  NAND2_X1 U7480 ( .A1(n9929), .A2(n9811), .ZN(n9327) );
  NAND2_X1 U7481 ( .A1(n9794), .A2(n9327), .ZN(n9771) );
  INV_X1 U7482 ( .A(n9772), .ZN(n9742) );
  OR2_X1 U7483 ( .A1(n9919), .A2(n9742), .ZN(n9331) );
  NAND2_X1 U7484 ( .A1(n9919), .A2(n9742), .ZN(n9337) );
  INV_X1 U7485 ( .A(n9730), .ZN(n9763) );
  OR2_X1 U7486 ( .A1(n9747), .A2(n9763), .ZN(n9339) );
  NAND2_X1 U7487 ( .A1(n9747), .A2(n9763), .ZN(n9338) );
  NAND2_X1 U7488 ( .A1(n9339), .A2(n9338), .ZN(n9740) );
  INV_X1 U7489 ( .A(n9462), .ZN(n9743) );
  OR2_X1 U7490 ( .A1(n9908), .A2(n9743), .ZN(n9340) );
  NAND2_X1 U7491 ( .A1(n9908), .A2(n9743), .ZN(n9428) );
  AND2_X1 U7492 ( .A1(n9344), .A2(n9701), .ZN(n9432) );
  NAND2_X1 U7493 ( .A1(n9345), .A2(n9700), .ZN(n9334) );
  NAND2_X1 U7494 ( .A1(n9334), .A2(n9344), .ZN(n9224) );
  OR2_X1 U7495 ( .A1(n9683), .A2(n9055), .ZN(n9348) );
  NAND2_X1 U7496 ( .A1(n9683), .A2(n9055), .ZN(n9257) );
  XNOR2_X1 U7497 ( .A(n9667), .B(n9459), .ZN(n9664) );
  INV_X1 U7498 ( .A(n9459), .ZN(n9220) );
  NAND2_X1 U7499 ( .A1(n9667), .A2(n9220), .ZN(n9349) );
  INV_X1 U7500 ( .A(n9458), .ZN(n5777) );
  OR2_X1 U7501 ( .A1(n9652), .A2(n5777), .ZN(n9351) );
  NAND2_X1 U7502 ( .A1(n9652), .A2(n5777), .ZN(n9352) );
  NAND2_X1 U7503 ( .A1(n9351), .A2(n9352), .ZN(n9646) );
  NAND2_X1 U7504 ( .A1(n9637), .A2(n9198), .ZN(n9226) );
  INV_X1 U7505 ( .A(n9456), .ZN(n9219) );
  XNOR2_X1 U7506 ( .A(n9950), .B(n9219), .ZN(n9620) );
  NAND2_X1 U7507 ( .A1(n6320), .A2(n9358), .ZN(n6359) );
  NAND2_X1 U7508 ( .A1(n6359), .A2(n9262), .ZN(n6358) );
  NAND2_X1 U7509 ( .A1(n6358), .A2(n9366), .ZN(n5779) );
  XNOR2_X1 U7510 ( .A(n5779), .B(n9370), .ZN(n5789) );
  NAND2_X1 U7511 ( .A1(n4301), .A2(n9395), .ZN(n5780) );
  INV_X1 U7512 ( .A(n9267), .ZN(n5790) );
  NAND2_X1 U7513 ( .A1(n5781), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5785) );
  NAND2_X1 U7514 ( .A1(n5782), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7515 ( .A1(n5513), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5783) );
  AND3_X1 U7516 ( .A1(n5785), .A2(n5784), .A3(n5783), .ZN(n9383) );
  NAND2_X1 U7517 ( .A1(n9454), .A2(n9841), .ZN(n5786) );
  OAI21_X1 U7518 ( .B1(n9383), .B2(n5787), .A(n5786), .ZN(n5788) );
  INV_X2 U7519 ( .A(n9855), .ZN(n10084) );
  AND2_X1 U7520 ( .A1(n10089), .A2(n5790), .ZN(n6699) );
  INV_X1 U7521 ( .A(n9852), .ZN(n10094) );
  NAND2_X1 U7522 ( .A1(n10094), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5792) );
  INV_X1 U7523 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5791) );
  OAI22_X1 U7524 ( .A1(n5793), .A2(n5792), .B1(n5791), .B2(n9855), .ZN(n5798)
         );
  AOI21_X1 U7525 ( .B1(n4374), .B2(n5746), .A(n9832), .ZN(n5794) );
  NAND2_X1 U7526 ( .A1(n5794), .A2(n9603), .ZN(n6379) );
  NAND2_X1 U7527 ( .A1(n5803), .A2(n9765), .ZN(n5795) );
  NOR2_X1 U7528 ( .A1(n6379), .A2(n9783), .ZN(n5797) );
  AOI211_X1 U7529 ( .C1(n10074), .C2(n5746), .A(n5798), .B(n5797), .ZN(n5799)
         );
  OAI21_X1 U7530 ( .B1(n6382), .B2(n10084), .A(n5799), .ZN(n5800) );
  NAND2_X1 U7531 ( .A1(n5802), .A2(n5801), .ZN(P1_U3356) );
  INV_X1 U7532 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5806) );
  MUX2_X1 U7533 ( .A(n5806), .B(n5805), .S(n10348), .Z(n5807) );
  NAND2_X1 U7534 ( .A1(n5807), .A2(n4993), .ZN(P1_U3521) );
  INV_X1 U7535 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6268) );
  NOR2_X1 U7536 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5809) );
  NAND4_X1 U7537 ( .A1(n5809), .A2(n5808), .A3(n5952), .A4(n10206), .ZN(n5818)
         );
  NAND2_X1 U7538 ( .A1(n5820), .A2(n5810), .ZN(n5811) );
  OAI21_X1 U7539 ( .B1(P2_IR_REG_19__SCAN_IN), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  NOR2_X2 U7540 ( .A1(n5951), .A2(n5819), .ZN(n6021) );
  NAND4_X1 U7541 ( .A1(n5831), .A2(n5820), .A3(n5827), .A4(n6095), .ZN(n5823)
         );
  NAND4_X1 U7542 ( .A1(n5814), .A2(n5822), .A3(n6098), .A4(n5821), .ZN(n5826)
         );
  NOR2_X1 U7543 ( .A1(n5823), .A2(n5826), .ZN(n5824) );
  NAND2_X1 U7544 ( .A1(n6021), .A2(n5824), .ZN(n6227) );
  NAND2_X1 U7545 ( .A1(n6227), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5825) );
  INV_X1 U7546 ( .A(n5826), .ZN(n5832) );
  NOR2_X1 U7547 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n5829) );
  AND4_X2 U7548 ( .A1(n5832), .A2(n5831), .A3(n5830), .A4(n5829), .ZN(n5833)
         );
  XNOR2_X2 U7549 ( .A(n5835), .B(n5836), .ZN(n6214) );
  NAND2_X1 U7550 ( .A1(n5841), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5837) );
  NAND2_X1 U7551 ( .A1(n5858), .A2(n4543), .ZN(n5890) );
  NAND2_X1 U7552 ( .A1(n7761), .A2(n4560), .ZN(n5840) );
  OR2_X1 U7553 ( .A1(n4474), .A2(n5838), .ZN(n5839) );
  OR2_X2 U7554 ( .A1(n8810), .A2(n8811), .ZN(n5844) );
  XNOR2_X2 U7555 ( .A(n5844), .B(n5843), .ZN(n7827) );
  NAND2_X1 U7556 ( .A1(n5845), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  INV_X1 U7557 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5847) );
  INV_X1 U7558 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5850) );
  OR2_X1 U7559 ( .A1(n5882), .A2(n5850), .ZN(n5856) );
  INV_X1 U7560 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5851) );
  OR2_X1 U7561 ( .A1(n5960), .A2(n5851), .ZN(n5855) );
  INV_X1 U7562 ( .A(n5957), .ZN(n5853) );
  AND4_X2 U7563 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n5880)
         );
  INV_X2 U7564 ( .A(n5880), .ZN(n6476) );
  NAND2_X1 U7565 ( .A1(n6437), .A2(n5907), .ZN(n5861) );
  OR2_X1 U7566 ( .A1(n8029), .A2(n6438), .ZN(n5860) );
  INV_X2 U7567 ( .A(n5862), .ZN(n10126) );
  NAND2_X1 U7568 ( .A1(n6476), .A2(n10126), .ZN(n8092) );
  NAND2_X1 U7569 ( .A1(n6057), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5866) );
  INV_X1 U7570 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6843) );
  OR2_X1 U7571 ( .A1(n5882), .A2(n6843), .ZN(n5865) );
  INV_X1 U7572 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6584) );
  OR2_X1 U7573 ( .A1(n5939), .A2(n6584), .ZN(n5864) );
  NOR2_X1 U7574 ( .A1(n6430), .A2(n5867), .ZN(n5869) );
  XNOR2_X1 U7575 ( .A(n5869), .B(n5868), .ZN(n8824) );
  MUX2_X1 U7576 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8824), .S(n5858), .Z(n6850) );
  INV_X1 U7577 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10157) );
  INV_X1 U7578 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7579 ( .A1(n5890), .A2(n6461), .ZN(n5876) );
  NAND2_X1 U7580 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5872) );
  MUX2_X1 U7581 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5872), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5874) );
  OR2_X1 U7582 ( .A1(n5858), .A2(n6606), .ZN(n5875) );
  NAND2_X1 U7583 ( .A1(n6926), .A2(n6928), .ZN(n5877) );
  NAND2_X1 U7584 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  NAND2_X1 U7585 ( .A1(n5880), .A2(n10126), .ZN(n5881) );
  NAND2_X1 U7586 ( .A1(n6929), .A2(n5881), .ZN(n7127) );
  OR2_X1 U7587 ( .A1(n5971), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5886) );
  INV_X1 U7588 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10160) );
  OR2_X1 U7589 ( .A1(n5957), .A2(n10160), .ZN(n5885) );
  NAND2_X1 U7590 ( .A1(n4296), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5884) );
  AND4_X2 U7591 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n6894)
         );
  INV_X2 U7592 ( .A(n6894), .ZN(n6271) );
  NAND2_X1 U7593 ( .A1(n5888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5887) );
  MUX2_X1 U7594 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5887), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5889) );
  NAND2_X1 U7595 ( .A1(n5889), .A2(n5903), .ZN(n6762) );
  OR2_X1 U7596 ( .A1(n6007), .A2(n6458), .ZN(n5892) );
  INV_X1 U7597 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6434) );
  OR2_X1 U7598 ( .A1(n8029), .A2(n6434), .ZN(n5891) );
  NAND2_X1 U7599 ( .A1(n7127), .A2(n5893), .ZN(n5895) );
  NAND2_X1 U7600 ( .A1(n6894), .A2(n10132), .ZN(n5894) );
  NAND2_X1 U7601 ( .A1(n5895), .A2(n5894), .ZN(n7114) );
  NAND2_X1 U7602 ( .A1(n4298), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5901) );
  INV_X1 U7603 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10162) );
  OR2_X1 U7604 ( .A1(n5957), .A2(n10162), .ZN(n5900) );
  NAND2_X1 U7605 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5897) );
  AND2_X1 U7606 ( .A1(n5913), .A2(n5897), .ZN(n7117) );
  OR2_X1 U7607 ( .A1(n5986), .A2(n10142), .ZN(n5898) );
  NAND4_X2 U7608 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(n8276)
         );
  INV_X2 U7609 ( .A(n8029), .ZN(n6100) );
  INV_X2 U7610 ( .A(n5858), .ZN(n6570) );
  NAND2_X1 U7611 ( .A1(n5903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5902) );
  MUX2_X1 U7612 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5902), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5906) );
  INV_X1 U7613 ( .A(n5903), .ZN(n5905) );
  INV_X1 U7614 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5904) );
  NAND2_X1 U7615 ( .A1(n5905), .A2(n5904), .ZN(n5920) );
  INV_X1 U7616 ( .A(n6881), .ZN(n6768) );
  AOI22_X1 U7617 ( .A1(n6100), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6570), .B2(
        n6768), .ZN(n5909) );
  NAND2_X1 U7618 ( .A1(n6429), .A2(n5907), .ZN(n5908) );
  NAND2_X1 U7619 ( .A1(n5909), .A2(n5908), .ZN(n7119) );
  OR2_X2 U7620 ( .A1(n8276), .A2(n7119), .ZN(n6269) );
  NAND2_X1 U7621 ( .A1(n8276), .A2(n7119), .ZN(n6270) );
  OR2_X1 U7622 ( .A1(n5957), .A2(n4776), .ZN(n5917) );
  NAND2_X1 U7623 ( .A1(n5913), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5914) );
  AND2_X1 U7624 ( .A1(n5925), .A2(n5914), .ZN(n7034) );
  OR2_X1 U7625 ( .A1(n5971), .A2(n7034), .ZN(n5916) );
  NAND2_X1 U7626 ( .A1(n4298), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5915) );
  INV_X1 U7627 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5918) );
  OR2_X1 U7628 ( .A1(n5986), .A2(n5918), .ZN(n5919) );
  NAND2_X2 U7629 ( .A1(n4328), .A2(n5919), .ZN(n8275) );
  INV_X2 U7630 ( .A(n8275), .ZN(n7075) );
  OR2_X1 U7631 ( .A1(n6455), .A2(n6007), .ZN(n5923) );
  NAND2_X1 U7632 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5921) );
  XNOR2_X1 U7633 ( .A(n5921), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6887) );
  AOI22_X1 U7634 ( .A1(n6100), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6570), .B2(
        n6887), .ZN(n5922) );
  NAND2_X1 U7635 ( .A1(n5923), .A2(n5922), .ZN(n10143) );
  NAND2_X1 U7636 ( .A1(n7075), .A2(n10143), .ZN(n8104) );
  INV_X1 U7637 ( .A(n10143), .ZN(n7025) );
  NAND2_X1 U7638 ( .A1(n7025), .A2(n8275), .ZN(n8110) );
  NAND2_X1 U7639 ( .A1(n8104), .A2(n8110), .ZN(n7008) );
  NAND2_X1 U7640 ( .A1(n7075), .A2(n7025), .ZN(n7166) );
  INV_X1 U7641 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5924) );
  NAND2_X1 U7642 ( .A1(n5925), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5926) );
  AND2_X1 U7643 ( .A1(n5942), .A2(n5926), .ZN(n7170) );
  OR2_X1 U7644 ( .A1(n5971), .A2(n7170), .ZN(n5928) );
  OR2_X1 U7645 ( .A1(n5957), .A2(n10166), .ZN(n5927) );
  NAND2_X1 U7646 ( .A1(n4297), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5930) );
  INV_X2 U7647 ( .A(n8274), .ZN(n8123) );
  OR2_X1 U7648 ( .A1(n6436), .A2(n6007), .ZN(n5934) );
  NAND2_X1 U7649 ( .A1(n5931), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5932) );
  XNOR2_X1 U7650 ( .A(n5932), .B(P2_IR_REG_6__SCAN_IN), .ZN(n7095) );
  AOI22_X1 U7651 ( .A1(n6100), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6570), .B2(
        n7095), .ZN(n5933) );
  NAND2_X1 U7652 ( .A1(n5934), .A2(n5933), .ZN(n8122) );
  NAND2_X1 U7653 ( .A1(n8123), .A2(n8122), .ZN(n6277) );
  NAND2_X1 U7654 ( .A1(n6277), .A2(n8106), .ZN(n7163) );
  NAND2_X1 U7655 ( .A1(n8123), .A2(n10151), .ZN(n5935) );
  NAND2_X1 U7656 ( .A1(n7165), .A2(n5935), .ZN(n7189) );
  NAND2_X1 U7657 ( .A1(n6441), .A2(n5907), .ZN(n5938) );
  NAND2_X1 U7658 ( .A1(n5951), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7659 ( .A(n5936), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7143) );
  AOI22_X1 U7660 ( .A1(n6100), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6570), .B2(
        n7143), .ZN(n5937) );
  NAND2_X1 U7661 ( .A1(n5938), .A2(n5937), .ZN(n7452) );
  INV_X2 U7662 ( .A(n5957), .ZN(n6199) );
  NAND2_X1 U7663 ( .A1(n6199), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5948) );
  INV_X1 U7664 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10245) );
  OR2_X1 U7665 ( .A1(n8022), .A2(n10245), .ZN(n5947) );
  NAND2_X1 U7666 ( .A1(n5942), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5943) );
  AND2_X1 U7667 ( .A1(n5958), .A2(n5943), .ZN(n7449) );
  OR2_X1 U7668 ( .A1(n5971), .A2(n7449), .ZN(n5946) );
  INV_X1 U7669 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7670 ( .A1(n5986), .A2(n5944), .ZN(n5945) );
  NAND2_X1 U7671 ( .A1(n7452), .A2(n8273), .ZN(n5949) );
  NAND2_X1 U7672 ( .A1(n7349), .A2(n7423), .ZN(n5950) );
  NAND2_X1 U7673 ( .A1(n6442), .A2(n5907), .ZN(n5956) );
  INV_X1 U7674 ( .A(n5951), .ZN(n5953) );
  NAND2_X1 U7675 ( .A1(n5953), .A2(n5952), .ZN(n5965) );
  NAND2_X1 U7676 ( .A1(n5965), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5954) );
  XNOR2_X1 U7677 ( .A(n5954), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7297) );
  AOI22_X1 U7678 ( .A1(n6100), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6570), .B2(
        n7297), .ZN(n5955) );
  NAND2_X2 U7679 ( .A1(n5956), .A2(n5955), .ZN(n7429) );
  NAND2_X1 U7680 ( .A1(n4298), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5964) );
  INV_X1 U7681 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7399) );
  OR2_X1 U7682 ( .A1(n5957), .A2(n7399), .ZN(n5963) );
  OR2_X2 U7683 ( .A1(n5958), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5974) );
  NAND2_X1 U7684 ( .A1(n5958), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5959) );
  AND2_X1 U7685 ( .A1(n5974), .A2(n5959), .ZN(n7520) );
  OR2_X1 U7686 ( .A1(n5971), .A2(n7520), .ZN(n5962) );
  INV_X1 U7687 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10211) );
  OR2_X1 U7688 ( .A1(n5986), .A2(n10211), .ZN(n5961) );
  NAND4_X1 U7689 ( .A1(n5964), .A2(n5963), .A3(n5962), .A4(n5961), .ZN(n8272)
         );
  INV_X1 U7690 ( .A(n8272), .ZN(n7455) );
  NAND2_X1 U7691 ( .A1(n6453), .A2(n5907), .ZN(n5970) );
  INV_X1 U7692 ( .A(n5965), .ZN(n5967) );
  INV_X1 U7693 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7694 ( .A1(n5967), .A2(n5966), .ZN(n5983) );
  NAND2_X1 U7695 ( .A1(n5983), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7696 ( .A(n5968), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7357) );
  AOI22_X1 U7697 ( .A1(n6100), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6570), .B2(
        n7357), .ZN(n5969) );
  NAND2_X1 U7698 ( .A1(n5970), .A2(n5969), .ZN(n7567) );
  NAND2_X1 U7699 ( .A1(n4297), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5980) );
  INV_X1 U7700 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7569) );
  OR2_X1 U7701 ( .A1(n5957), .A2(n7569), .ZN(n5979) );
  NAND2_X1 U7702 ( .A1(n5974), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5975) );
  AND2_X1 U7703 ( .A1(n5987), .A2(n5975), .ZN(n7615) );
  OR2_X1 U7704 ( .A1(n5971), .A2(n7615), .ZN(n5978) );
  INV_X1 U7705 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5976) );
  OR2_X1 U7706 ( .A1(n5986), .A2(n5976), .ZN(n5977) );
  OR2_X1 U7707 ( .A1(n7567), .A2(n7560), .ZN(n8139) );
  NAND2_X1 U7708 ( .A1(n7567), .A2(n7560), .ZN(n8129) );
  NAND2_X1 U7709 ( .A1(n7429), .A2(n7557), .ZN(n7410) );
  AND2_X1 U7710 ( .A1(n8043), .A2(n7410), .ZN(n5981) );
  INV_X1 U7711 ( .A(n7560), .ZN(n8271) );
  OR2_X1 U7712 ( .A1(n7567), .A2(n8271), .ZN(n5982) );
  NAND2_X1 U7713 ( .A1(n7412), .A2(n5982), .ZN(n7643) );
  NAND2_X1 U7714 ( .A1(n5994), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5984) );
  AOI22_X1 U7715 ( .A1(n6100), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6570), .B2(
        n8295), .ZN(n5985) );
  NAND2_X1 U7716 ( .A1(n4297), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5992) );
  INV_X1 U7717 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n7650) );
  OR2_X1 U7718 ( .A1(n5986), .A2(n7650), .ZN(n5991) );
  OR2_X2 U7719 ( .A1(n5987), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6000) );
  NAND2_X1 U7720 ( .A1(n5987), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5988) );
  AND2_X1 U7721 ( .A1(n6000), .A2(n5988), .ZN(n7691) );
  OR2_X1 U7722 ( .A1(n5971), .A2(n7691), .ZN(n5990) );
  INV_X1 U7723 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8294) );
  OR2_X1 U7724 ( .A1(n5957), .A2(n8294), .ZN(n5989) );
  NAND2_X1 U7725 ( .A1(n7770), .A2(n8270), .ZN(n5993) );
  NAND2_X1 U7726 ( .A1(n6474), .A2(n4560), .ZN(n5999) );
  INV_X1 U7727 ( .A(n5994), .ZN(n5996) );
  INV_X1 U7728 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7729 ( .A1(n5996), .A2(n5995), .ZN(n6008) );
  NAND2_X1 U7730 ( .A1(n6008), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5997) );
  XNOR2_X1 U7731 ( .A(n5997), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8305) );
  AOI22_X1 U7732 ( .A1(n6100), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6570), .B2(
        n8305), .ZN(n5998) );
  NAND2_X1 U7733 ( .A1(n4297), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6005) );
  INV_X1 U7734 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7606) );
  OR2_X1 U7735 ( .A1(n6202), .A2(n7606), .ZN(n6004) );
  OR2_X2 U7736 ( .A1(n6000), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7737 ( .A1(n6000), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6001) );
  AND2_X1 U7738 ( .A1(n6014), .A2(n6001), .ZN(n7611) );
  OR2_X1 U7739 ( .A1(n5971), .A2(n7611), .ZN(n6003) );
  INV_X1 U7740 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7602) );
  OR2_X1 U7741 ( .A1(n5957), .A2(n7602), .ZN(n6002) );
  NAND2_X1 U7742 ( .A1(n7971), .A2(n7884), .ZN(n8148) );
  OR2_X1 U7743 ( .A1(n7770), .A2(n8270), .ZN(n7596) );
  AND2_X1 U7744 ( .A1(n7768), .A2(n7596), .ZN(n6006) );
  INV_X1 U7745 ( .A(n7884), .ZN(n8269) );
  NAND2_X1 U7746 ( .A1(n7971), .A2(n8269), .ZN(n7659) );
  OR2_X1 U7747 ( .A1(n6482), .A2(n6007), .ZN(n6011) );
  OAI21_X1 U7748 ( .B1(n6008), .B2(P2_IR_REG_11__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6009) );
  AOI22_X1 U7749 ( .A1(n6100), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8338), .B2(
        n6570), .ZN(n6010) );
  NAND2_X1 U7750 ( .A1(n4298), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6019) );
  INV_X1 U7751 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7711) );
  OR2_X1 U7752 ( .A1(n6202), .A2(n7711), .ZN(n6018) );
  NAND2_X1 U7753 ( .A1(n6014), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6015) );
  AND2_X1 U7754 ( .A1(n6025), .A2(n6015), .ZN(n7892) );
  OR2_X1 U7755 ( .A1(n5971), .A2(n7892), .ZN(n6017) );
  INV_X1 U7756 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8337) );
  OR2_X1 U7757 ( .A1(n5957), .A2(n8337), .ZN(n6016) );
  NAND4_X1 U7758 ( .A1(n6019), .A2(n6018), .A3(n6017), .A4(n6016), .ZN(n8268)
         );
  NAND2_X1 U7759 ( .A1(n8153), .A2(n8268), .ZN(n6020) );
  AND2_X1 U7760 ( .A1(n7659), .A2(n6020), .ZN(n7622) );
  INV_X1 U7761 ( .A(n6021), .ZN(n6022) );
  NAND2_X1 U7762 ( .A1(n6022), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6023) );
  XNOR2_X1 U7763 ( .A(n6023), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8355) );
  AOI22_X1 U7764 ( .A1(n6100), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6570), .B2(
        n8355), .ZN(n6024) );
  NAND2_X1 U7765 ( .A1(n6199), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6031) );
  INV_X1 U7766 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8336) );
  OR2_X1 U7767 ( .A1(n8022), .A2(n8336), .ZN(n6030) );
  NAND2_X1 U7768 ( .A1(n6025), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6026) );
  AND2_X1 U7769 ( .A1(n6039), .A2(n6026), .ZN(n7954) );
  OR2_X1 U7770 ( .A1(n5971), .A2(n7954), .ZN(n6029) );
  INV_X1 U7771 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7772 ( .A1(n6202), .A2(n6027), .ZN(n6028) );
  NAND4_X1 U7773 ( .A1(n6031), .A2(n6030), .A3(n6029), .A4(n6028), .ZN(n8267)
         );
  NAND2_X1 U7774 ( .A1(n8157), .A2(n8267), .ZN(n8161) );
  INV_X1 U7775 ( .A(n8059), .ZN(n6032) );
  OR2_X1 U7776 ( .A1(n8153), .A2(n8268), .ZN(n7623) );
  OR2_X1 U7777 ( .A1(n8059), .A2(n7623), .ZN(n6033) );
  NAND2_X1 U7778 ( .A1(n6593), .A2(n4560), .ZN(n6038) );
  INV_X1 U7779 ( .A(n5834), .ZN(n6035) );
  NAND2_X1 U7780 ( .A1(n6035), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6036) );
  XNOR2_X1 U7781 ( .A(n6036), .B(P2_IR_REG_14__SCAN_IN), .ZN(n8378) );
  AOI22_X1 U7782 ( .A1(n6100), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6570), .B2(
        n8378), .ZN(n6037) );
  NAND2_X1 U7783 ( .A1(n6039), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7784 ( .A1(n6053), .A2(n6040), .ZN(n8676) );
  NAND2_X1 U7785 ( .A1(n6216), .A2(n8676), .ZN(n6044) );
  INV_X1 U7786 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8377) );
  OR2_X1 U7787 ( .A1(n8022), .A2(n8377), .ZN(n6043) );
  INV_X1 U7788 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n7699) );
  OR2_X1 U7789 ( .A1(n6202), .A2(n7699), .ZN(n6042) );
  INV_X1 U7790 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7704) );
  OR2_X1 U7791 ( .A1(n5957), .A2(n7704), .ZN(n6041) );
  NAND4_X1 U7792 ( .A1(n6044), .A2(n6043), .A3(n6042), .A4(n6041), .ZN(n8266)
         );
  NAND2_X1 U7793 ( .A1(n7839), .A2(n8266), .ZN(n6046) );
  NOR2_X1 U7794 ( .A1(n7839), .A2(n8266), .ZN(n6045) );
  NAND2_X1 U7795 ( .A1(n6727), .A2(n4560), .ZN(n6050) );
  NAND2_X1 U7796 ( .A1(n6047), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6048) );
  XNOR2_X1 U7797 ( .A(n6048), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8402) );
  AOI22_X1 U7798 ( .A1(n6100), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6570), .B2(
        n8402), .ZN(n6049) );
  NAND2_X1 U7799 ( .A1(n6053), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U7800 ( .A1(n6068), .A2(n6054), .ZN(n8012) );
  NAND2_X1 U7801 ( .A1(n8012), .A2(n6216), .ZN(n6060) );
  NAND2_X1 U7802 ( .A1(n6199), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U7803 ( .A1(n4298), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6055) );
  AND2_X1 U7804 ( .A1(n6056), .A2(n6055), .ZN(n6059) );
  NAND2_X1 U7805 ( .A1(n6057), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7806 ( .A1(n8002), .A2(n7838), .ZN(n8176) );
  NAND2_X1 U7807 ( .A1(n8169), .A2(n8176), .ZN(n8061) );
  NAND2_X1 U7808 ( .A1(n7730), .A2(n8061), .ZN(n7733) );
  INV_X1 U7809 ( .A(n7838), .ZN(n8265) );
  NAND2_X1 U7810 ( .A1(n8002), .A2(n8265), .ZN(n6061) );
  NAND2_X1 U7811 ( .A1(n6062), .A2(n4560), .ZN(n6067) );
  INV_X1 U7812 ( .A(n6063), .ZN(n6064) );
  NAND2_X1 U7813 ( .A1(n6064), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6065) );
  XNOR2_X1 U7814 ( .A(n6065), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8424) );
  AOI22_X1 U7815 ( .A1(n6100), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6570), .B2(
        n8424), .ZN(n6066) );
  NAND2_X1 U7816 ( .A1(n6068), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7817 ( .A1(n6078), .A2(n6069), .ZN(n7910) );
  NAND2_X1 U7818 ( .A1(n7910), .A2(n6216), .ZN(n6072) );
  AOI22_X1 U7819 ( .A1(n6199), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n4298), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n6071) );
  INV_X1 U7820 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n10243) );
  OR2_X1 U7821 ( .A1(n6202), .A2(n10243), .ZN(n6070) );
  NAND2_X1 U7822 ( .A1(n8737), .A2(n8657), .ZN(n8177) );
  NAND2_X1 U7823 ( .A1(n8179), .A2(n8177), .ZN(n6290) );
  NAND2_X1 U7824 ( .A1(n8737), .A2(n8264), .ZN(n6073) );
  NAND2_X1 U7825 ( .A1(n6723), .A2(n4560), .ZN(n6077) );
  NAND2_X1 U7826 ( .A1(n6074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6075) );
  AOI22_X1 U7827 ( .A1(n6100), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6570), .B2(
        n8451), .ZN(n6076) );
  NAND2_X1 U7828 ( .A1(n6078), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7829 ( .A1(n6085), .A2(n6079), .ZN(n8665) );
  NAND2_X1 U7830 ( .A1(n8665), .A2(n6216), .ZN(n6082) );
  AOI22_X1 U7831 ( .A1(n6199), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n4297), .B2(
        P2_REG2_REG_17__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7832 ( .A1(n6057), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7833 ( .A1(n8800), .A2(n8637), .ZN(n8042) );
  NAND2_X1 U7834 ( .A1(n8062), .A2(n8042), .ZN(n8171) );
  INV_X1 U7835 ( .A(n8637), .ZN(n7783) );
  INV_X1 U7836 ( .A(n8633), .ZN(n6093) );
  NAND2_X1 U7837 ( .A1(n6742), .A2(n5907), .ZN(n6084) );
  XNOR2_X1 U7838 ( .A(n6096), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8475) );
  AOI22_X1 U7839 ( .A1(n6100), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6570), .B2(
        n8475), .ZN(n6083) );
  NAND2_X1 U7840 ( .A1(n6085), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7841 ( .A1(n6105), .A2(n6086), .ZN(n8642) );
  NAND2_X1 U7842 ( .A1(n8642), .A2(n6216), .ZN(n6091) );
  INV_X1 U7843 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8796) );
  NAND2_X1 U7844 ( .A1(n6199), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U7845 ( .A1(n4297), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6087) );
  OAI211_X1 U7846 ( .C1(n8796), .C2(n6202), .A(n6088), .B(n6087), .ZN(n6089)
         );
  INV_X1 U7847 ( .A(n6089), .ZN(n6090) );
  NAND2_X1 U7848 ( .A1(n8726), .A2(n8659), .ZN(n8079) );
  INV_X1 U7849 ( .A(n8634), .ZN(n6092) );
  OR2_X1 U7850 ( .A1(n8726), .A2(n8263), .ZN(n6094) );
  NAND2_X1 U7851 ( .A1(n7003), .A2(n4560), .ZN(n6102) );
  NAND2_X1 U7852 ( .A1(n6096), .A2(n6095), .ZN(n6097) );
  AOI22_X1 U7853 ( .A1(n6100), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6259), .B2(
        n6570), .ZN(n6101) );
  INV_X1 U7854 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7855 ( .A1(n6105), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6106) );
  NAND2_X1 U7856 ( .A1(n6116), .A2(n6106), .ZN(n8627) );
  NAND2_X1 U7857 ( .A1(n8627), .A2(n6216), .ZN(n6111) );
  INV_X1 U7858 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U7859 ( .A1(n4298), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7860 ( .A1(n6057), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6107) );
  OAI211_X1 U7861 ( .C1(n5957), .C2(n8723), .A(n6108), .B(n6107), .ZN(n6109)
         );
  INV_X1 U7862 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7863 ( .A1(n7854), .A2(n8638), .ZN(n8188) );
  NAND2_X1 U7864 ( .A1(n7854), .A2(n8262), .ZN(n6113) );
  NAND2_X1 U7865 ( .A1(n7107), .A2(n5907), .ZN(n6115) );
  OR2_X1 U7866 ( .A1(n4474), .A2(n7110), .ZN(n6114) );
  NAND2_X1 U7867 ( .A1(n6116), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7868 ( .A1(n6128), .A2(n6117), .ZN(n8613) );
  NAND2_X1 U7869 ( .A1(n8613), .A2(n6216), .ZN(n6123) );
  INV_X1 U7870 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7871 ( .A1(n6199), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6119) );
  NAND2_X1 U7872 ( .A1(n4297), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6118) );
  OAI211_X1 U7873 ( .C1(n6120), .C2(n6202), .A(n6119), .B(n6118), .ZN(n6121)
         );
  INV_X1 U7874 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7875 ( .A1(n8711), .A2(n8621), .ZN(n8596) );
  INV_X1 U7876 ( .A(n8621), .ZN(n8261) );
  OR2_X1 U7877 ( .A1(n8711), .A2(n8261), .ZN(n6124) );
  NAND2_X1 U7878 ( .A1(n6125), .A2(n4560), .ZN(n6127) );
  OR2_X1 U7879 ( .A1(n4474), .A2(n7250), .ZN(n6126) );
  NAND2_X1 U7880 ( .A1(n6128), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7881 ( .A1(n6136), .A2(n6129), .ZN(n8600) );
  INV_X1 U7882 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7883 ( .A1(n6199), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7884 ( .A1(n4298), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6130) );
  OAI211_X1 U7885 ( .C1(n6132), .C2(n6202), .A(n6131), .B(n6130), .ZN(n6133)
         );
  NAND2_X1 U7886 ( .A1(n8706), .A2(n8608), .ZN(n8194) );
  NAND2_X1 U7887 ( .A1(n8201), .A2(n8194), .ZN(n8590) );
  INV_X1 U7888 ( .A(n8608), .ZN(n8260) );
  NAND2_X1 U7889 ( .A1(n7285), .A2(n4560), .ZN(n6135) );
  OR2_X1 U7890 ( .A1(n4474), .A2(n7290), .ZN(n6134) );
  OR2_X2 U7891 ( .A1(n6136), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6145) );
  NAND2_X1 U7892 ( .A1(n6136), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7893 ( .A1(n6145), .A2(n6137), .ZN(n8583) );
  INV_X1 U7894 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U7895 ( .A1(n6199), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6139) );
  NAND2_X1 U7896 ( .A1(n4297), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6138) );
  OAI211_X1 U7897 ( .C1(n8780), .C2(n6202), .A(n6139), .B(n6138), .ZN(n6140)
         );
  NAND2_X1 U7898 ( .A1(n8703), .A2(n8591), .ZN(n8203) );
  NAND2_X1 U7899 ( .A1(n8198), .A2(n8203), .ZN(n8200) );
  NAND2_X1 U7900 ( .A1(n8580), .A2(n8200), .ZN(n6142) );
  OR2_X1 U7901 ( .A1(n8703), .A2(n8574), .ZN(n6141) );
  NAND2_X1 U7902 ( .A1(n7396), .A2(n4560), .ZN(n6144) );
  OR2_X1 U7903 ( .A1(n4474), .A2(n7394), .ZN(n6143) );
  NAND2_X1 U7904 ( .A1(n6145), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7905 ( .A1(n6175), .A2(n6146), .ZN(n8576) );
  NAND2_X1 U7906 ( .A1(n8576), .A2(n6216), .ZN(n6151) );
  INV_X1 U7907 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10330) );
  NAND2_X1 U7908 ( .A1(n4297), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7909 ( .A1(n6057), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U7910 ( .C1(n5957), .C2(n10330), .A(n6148), .B(n6147), .ZN(n6149)
         );
  INV_X1 U7911 ( .A(n6149), .ZN(n6150) );
  NOR2_X1 U7912 ( .A1(n8775), .A2(n8553), .ZN(n6153) );
  NAND2_X1 U7913 ( .A1(n8775), .A2(n8553), .ZN(n6152) );
  NAND2_X1 U7914 ( .A1(n7637), .A2(n4560), .ZN(n6155) );
  OR2_X1 U7915 ( .A1(n4474), .A2(n7638), .ZN(n6154) );
  NAND2_X2 U7916 ( .A1(n6155), .A2(n6154), .ZN(n8762) );
  NOR2_X4 U7917 ( .A1(n6175), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6157) );
  INV_X1 U7918 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6156) );
  INV_X1 U7919 ( .A(n6157), .ZN(n6177) );
  NAND2_X1 U7920 ( .A1(n6177), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7921 ( .A1(n6166), .A2(n6158), .ZN(n7900) );
  NAND2_X1 U7922 ( .A1(n7900), .A2(n6216), .ZN(n6163) );
  INV_X1 U7923 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n10216) );
  NAND2_X1 U7924 ( .A1(n6057), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6160) );
  NAND2_X1 U7925 ( .A1(n6199), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6159) );
  OAI211_X1 U7926 ( .C1(n8022), .C2(n10216), .A(n6160), .B(n6159), .ZN(n6161)
         );
  INV_X1 U7927 ( .A(n6161), .ZN(n6162) );
  NAND2_X2 U7928 ( .A1(n6163), .A2(n6162), .ZN(n8554) );
  OR2_X1 U7929 ( .A1(n8762), .A2(n8554), .ZN(n8529) );
  INV_X1 U7930 ( .A(n8529), .ZN(n6194) );
  INV_X2 U7931 ( .A(n8554), .ZN(n8532) );
  OR2_X2 U7932 ( .A1(n8762), .A2(n8532), .ZN(n8215) );
  NAND2_X1 U7933 ( .A1(n8762), .A2(n8532), .ZN(n8216) );
  NAND2_X1 U7934 ( .A1(n7668), .A2(n4560), .ZN(n6165) );
  OR2_X1 U7935 ( .A1(n4474), .A2(n7669), .ZN(n6164) );
  NAND2_X2 U7936 ( .A1(n6165), .A2(n6164), .ZN(n8756) );
  NAND2_X1 U7937 ( .A1(n6166), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6167) );
  INV_X1 U7938 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U7939 ( .A1(n6199), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7940 ( .A1(n4298), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6168) );
  OAI211_X1 U7941 ( .C1(n10301), .C2(n6202), .A(n6169), .B(n6168), .ZN(n6170)
         );
  INV_X1 U7942 ( .A(n6170), .ZN(n6171) );
  NAND2_X1 U7943 ( .A1(n7571), .A2(n4560), .ZN(n6174) );
  OR2_X1 U7944 ( .A1(n4474), .A2(n7654), .ZN(n6173) );
  NAND2_X1 U7945 ( .A1(n6175), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7946 ( .A1(n6177), .A2(n6176), .ZN(n8559) );
  NAND2_X1 U7947 ( .A1(n8559), .A2(n6216), .ZN(n6182) );
  INV_X1 U7948 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n8768) );
  NAND2_X1 U7949 ( .A1(n4298), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7950 ( .A1(n6199), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6178) );
  OAI211_X1 U7951 ( .C1(n8768), .C2(n6202), .A(n6179), .B(n6178), .ZN(n6180)
         );
  INV_X1 U7952 ( .A(n6180), .ZN(n6181) );
  AOI22_X1 U7953 ( .A1(n8756), .A2(n8520), .B1(n8529), .B2(n8551), .ZN(n6183)
         );
  INV_X1 U7954 ( .A(n6185), .ZN(n6184) );
  INV_X1 U7955 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U7956 ( .A1(n6185), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7957 ( .A1(n6197), .A2(n6186), .ZN(n8526) );
  NAND2_X1 U7958 ( .A1(n8526), .A2(n6216), .ZN(n6191) );
  INV_X1 U7959 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U7960 ( .A1(n6199), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U7961 ( .A1(n4297), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6187) );
  OAI211_X1 U7962 ( .C1(n8750), .C2(n6202), .A(n6188), .B(n6187), .ZN(n6189)
         );
  INV_X1 U7963 ( .A(n6189), .ZN(n6190) );
  NAND2_X1 U7964 ( .A1(n7707), .A2(n4560), .ZN(n6193) );
  OR2_X1 U7965 ( .A1(n4474), .A2(n7717), .ZN(n6192) );
  NOR2_X1 U7966 ( .A1(n8756), .A2(n8520), .ZN(n8514) );
  NOR2_X1 U7967 ( .A1(n8769), .A2(n8572), .ZN(n6390) );
  NOR2_X1 U7968 ( .A1(n6194), .A2(n6390), .ZN(n8513) );
  NOR2_X1 U7969 ( .A1(n8512), .A2(n8513), .ZN(n6195) );
  AOI211_X1 U7970 ( .C1(n8533), .C2(n7834), .A(n8514), .B(n6195), .ZN(n6196)
         );
  NAND2_X1 U7971 ( .A1(n8751), .A2(n8259), .ZN(n6337) );
  NAND2_X1 U7972 ( .A1(n6332), .A2(n6337), .ZN(n6206) );
  NAND2_X1 U7973 ( .A1(n6197), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7974 ( .A1(n7753), .A2(n6198), .ZN(n8504) );
  NAND2_X1 U7975 ( .A1(n8504), .A2(n6216), .ZN(n6205) );
  INV_X1 U7976 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n10328) );
  NAND2_X1 U7977 ( .A1(n6199), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7978 ( .A1(n4297), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6200) );
  OAI211_X1 U7979 ( .C1(n10328), .C2(n6202), .A(n6201), .B(n6200), .ZN(n6203)
         );
  INV_X1 U7980 ( .A(n6203), .ZN(n6204) );
  XNOR2_X1 U7981 ( .A(n8505), .B(n8519), .ZN(n8068) );
  XNOR2_X1 U7982 ( .A(n6206), .B(n8068), .ZN(n6212) );
  NAND2_X1 U7983 ( .A1(n6207), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6208) );
  INV_X1 U7984 ( .A(n8242), .ZN(n6210) );
  NAND2_X1 U7985 ( .A1(n6213), .A2(n6210), .ZN(n8039) );
  NAND2_X1 U7986 ( .A1(n6259), .A2(n8255), .ZN(n6211) );
  NAND2_X1 U7987 ( .A1(n6212), .A2(n8640), .ZN(n6226) );
  INV_X1 U7988 ( .A(n6578), .ZN(n8251) );
  NAND2_X1 U7989 ( .A1(n8251), .A2(n8477), .ZN(n6215) );
  NAND2_X1 U7990 ( .A1(n5858), .A2(n6215), .ZN(n6855) );
  INV_X1 U7991 ( .A(n7753), .ZN(n6217) );
  NAND2_X1 U7992 ( .A1(n6217), .A2(n6216), .ZN(n8027) );
  NAND2_X1 U7993 ( .A1(n4298), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6220) );
  NAND2_X1 U7994 ( .A1(n6057), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6219) );
  OAI211_X1 U7995 ( .C1(n6420), .C2(n5957), .A(n6220), .B(n6219), .ZN(n6221)
         );
  INV_X1 U7996 ( .A(n6221), .ZN(n6222) );
  INV_X1 U7997 ( .A(n6855), .ZN(n6824) );
  NAND2_X1 U7998 ( .A1(n6226), .A2(n6225), .ZN(n8510) );
  AOI21_X1 U7999 ( .B1(n10144), .B2(n8505), .A(n8510), .ZN(n6314) );
  OR2_X1 U8000 ( .A1(n8222), .A2(n8241), .ZN(n6814) );
  OAI21_X2 U8001 ( .B1(n6227), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U8002 ( .A1(n6241), .A2(n6242), .ZN(n6228) );
  NAND2_X1 U8003 ( .A1(n6232), .A2(n6231), .ZN(n6233) );
  XNOR2_X2 U8004 ( .A(n6230), .B(n6229), .ZN(n6244) );
  INV_X1 U8005 ( .A(n6244), .ZN(n6240) );
  NAND2_X1 U8006 ( .A1(n6235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6236) );
  MUX2_X1 U8007 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6236), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6238) );
  NOR2_X1 U8008 ( .A1(n6243), .A2(n7671), .ZN(n6239) );
  XNOR2_X1 U8009 ( .A(n6243), .B(P2_B_REG_SCAN_IN), .ZN(n6245) );
  NAND2_X1 U8010 ( .A1(n6245), .A2(n6244), .ZN(n6247) );
  NAND2_X1 U8011 ( .A1(n6247), .A2(n6246), .ZN(n6261) );
  NOR2_X1 U8012 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .ZN(
        n6251) );
  NOR4_X1 U8013 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n6250) );
  NOR4_X1 U8014 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6249) );
  NOR4_X1 U8015 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n6248) );
  NAND4_X1 U8016 ( .A1(n6251), .A2(n6250), .A3(n6249), .A4(n6248), .ZN(n6257)
         );
  NOR4_X1 U8017 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6255) );
  NOR4_X1 U8018 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6254) );
  NOR4_X1 U8019 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6253) );
  NOR4_X1 U8020 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6252) );
  NAND4_X1 U8021 ( .A1(n6255), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(n6256)
         );
  NOR2_X1 U8022 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  NAND3_X1 U8023 ( .A1(n6814), .A2(n6820), .A3(n6303), .ZN(n6401) );
  NOR2_X1 U8024 ( .A1(n6401), .A2(n6399), .ZN(n6267) );
  NAND2_X1 U8025 ( .A1(n8487), .A2(n8255), .ZN(n6298) );
  OR2_X1 U8026 ( .A1(n6298), .A2(n8242), .ZN(n6260) );
  NAND2_X1 U8027 ( .A1(n8222), .A2(n6260), .ZN(n6265) );
  NAND2_X1 U8028 ( .A1(n6243), .A2(n7671), .ZN(n6485) );
  OAI21_X2 U8029 ( .B1(n6261), .B2(P2_D_REG_0__SCAN_IN), .A(n6485), .ZN(n6266)
         );
  OR2_X1 U8030 ( .A1(n6261), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6263) );
  NAND2_X1 U8031 ( .A1(n6244), .A2(n7671), .ZN(n6262) );
  NAND2_X1 U8032 ( .A1(n8808), .A2(n6265), .ZN(n6264) );
  OAI21_X1 U8033 ( .B1(n6265), .B2(n6266), .A(n6264), .ZN(n6404) );
  INV_X2 U8034 ( .A(n6266), .ZN(n6848) );
  NAND2_X1 U8035 ( .A1(n8808), .A2(n6848), .ZN(n6308) );
  MUX2_X1 U8036 ( .A(n6268), .B(n6314), .S(n10168), .Z(n6302) );
  AND2_X1 U8037 ( .A1(n7423), .A2(n7452), .ZN(n6278) );
  OR2_X1 U8038 ( .A1(n7429), .A2(n7455), .ZN(n8135) );
  NAND2_X1 U8039 ( .A1(n7349), .A2(n8273), .ZN(n8134) );
  OAI211_X1 U8040 ( .C1(n6278), .C2(n8106), .A(n8135), .B(n8134), .ZN(n6279)
         );
  INV_X1 U8041 ( .A(n6279), .ZN(n7403) );
  AND2_X1 U8042 ( .A1(n7403), .A2(n8110), .ZN(n6276) );
  NAND2_X2 U8043 ( .A1(n6270), .A2(n6269), .ZN(n8100) );
  NAND2_X1 U8044 ( .A1(n6271), .A2(n10132), .ZN(n8102) );
  INV_X1 U8045 ( .A(n8093), .ZN(n8111) );
  INV_X1 U8046 ( .A(n6272), .ZN(n8090) );
  INV_X1 U8047 ( .A(n8278), .ZN(n6273) );
  NAND2_X1 U8048 ( .A1(n6273), .A2(n6850), .ZN(n8087) );
  OAI21_X2 U8049 ( .B1(n7135), .B2(n8087), .A(n8088), .ZN(n6920) );
  NAND2_X1 U8050 ( .A1(n8090), .A2(n6920), .ZN(n6921) );
  AND2_X1 U8051 ( .A1(n8093), .A2(n8094), .ZN(n6274) );
  NAND2_X1 U8052 ( .A1(n6921), .A2(n6274), .ZN(n7112) );
  INV_X1 U8053 ( .A(n8276), .ZN(n7009) );
  NAND2_X1 U8054 ( .A1(n7009), .A2(n7119), .ZN(n8103) );
  AND2_X1 U8055 ( .A1(n8104), .A2(n6277), .ZN(n8114) );
  INV_X1 U8056 ( .A(n6278), .ZN(n8127) );
  OR2_X1 U8057 ( .A1(n7401), .A2(n6279), .ZN(n6282) );
  NAND2_X1 U8058 ( .A1(n7429), .A2(n7455), .ZN(n8128) );
  INV_X1 U8059 ( .A(n8128), .ZN(n6280) );
  NOR2_X1 U8060 ( .A1(n8043), .A2(n6280), .ZN(n6281) );
  NAND3_X1 U8061 ( .A1(n6283), .A2(n6282), .A3(n6281), .ZN(n7407) );
  INV_X1 U8062 ( .A(n8148), .ZN(n6284) );
  INV_X1 U8063 ( .A(n8268), .ZN(n8152) );
  OR2_X1 U8064 ( .A1(n8153), .A2(n8152), .ZN(n8155) );
  NAND2_X1 U8065 ( .A1(n7658), .A2(n8155), .ZN(n7633) );
  NAND2_X1 U8066 ( .A1(n8157), .A2(n7888), .ZN(n6285) );
  NAND2_X1 U8067 ( .A1(n7633), .A2(n6285), .ZN(n6287) );
  OR2_X1 U8068 ( .A1(n8157), .A2(n7888), .ZN(n6286) );
  NOR2_X1 U8069 ( .A1(n7839), .A2(n7950), .ZN(n8165) );
  NAND2_X1 U8070 ( .A1(n7839), .A2(n7950), .ZN(n7697) );
  INV_X1 U8071 ( .A(n8176), .ZN(n6288) );
  OAI21_X1 U8072 ( .B1(n7729), .B2(n6288), .A(n8169), .ZN(n6289) );
  INV_X1 U8073 ( .A(n6289), .ZN(n7724) );
  NAND2_X1 U8074 ( .A1(n7724), .A2(n8065), .ZN(n7723) );
  NAND2_X1 U8075 ( .A1(n8595), .A2(n8594), .ZN(n6293) );
  NAND2_X1 U8076 ( .A1(n8194), .A2(n8596), .ZN(n8192) );
  INV_X1 U8077 ( .A(n8188), .ZN(n8184) );
  AND2_X1 U8078 ( .A1(n8595), .A2(n8184), .ZN(n6291) );
  NOR2_X1 U8079 ( .A1(n8192), .A2(n6291), .ZN(n6292) );
  OAI21_X1 U8080 ( .B1(n8626), .B2(n6293), .A(n6292), .ZN(n6294) );
  NAND2_X1 U8081 ( .A1(n6294), .A2(n8201), .ZN(n8579) );
  INV_X1 U8082 ( .A(n8775), .ZN(n6295) );
  NAND2_X1 U8083 ( .A1(n8769), .A2(n7850), .ZN(n8204) );
  INV_X1 U8084 ( .A(n8553), .ZN(n8582) );
  NAND2_X1 U8085 ( .A1(n8775), .A2(n8582), .ZN(n8562) );
  NAND2_X1 U8086 ( .A1(n8560), .A2(n4991), .ZN(n6297) );
  INV_X2 U8087 ( .A(n8520), .ZN(n7991) );
  NAND2_X1 U8088 ( .A1(n8751), .A2(n8533), .ZN(n8224) );
  XNOR2_X1 U8089 ( .A(n6329), .B(n8068), .ZN(n8508) );
  INV_X1 U8090 ( .A(n6298), .ZN(n6300) );
  INV_X1 U8091 ( .A(n8241), .ZN(n6299) );
  NAND2_X1 U8092 ( .A1(n8245), .A2(n7288), .ZN(n10127) );
  NAND2_X1 U8093 ( .A1(n10168), .A2(n10153), .ZN(n8716) );
  NAND2_X1 U8094 ( .A1(n6302), .A2(n6301), .ZN(P2_U3487) );
  NOR2_X1 U8095 ( .A1(n8808), .A2(n6307), .ZN(n6304) );
  NAND2_X1 U8096 ( .A1(n4397), .A2(n8255), .ZN(n6309) );
  NAND2_X1 U8097 ( .A1(n6309), .A2(n8222), .ZN(n6305) );
  INV_X1 U8098 ( .A(n8245), .ZN(n6306) );
  NAND2_X1 U8099 ( .A1(n6807), .A2(n8671), .ZN(n6810) );
  NAND2_X1 U8100 ( .A1(n6858), .A2(n6810), .ZN(n6313) );
  NOR2_X1 U8101 ( .A1(n6308), .A2(n6307), .ZN(n6811) );
  NAND2_X1 U8102 ( .A1(n6811), .A2(n6820), .ZN(n6826) );
  INV_X1 U8103 ( .A(n6309), .ZN(n6310) );
  NAND2_X1 U8104 ( .A1(n6310), .A2(n6847), .ZN(n6817) );
  AND2_X1 U8105 ( .A1(n6817), .A2(n6856), .ZN(n6311) );
  MUX2_X1 U8106 ( .A(n10328), .B(n6314), .S(n10155), .Z(n6316) );
  INV_X1 U8107 ( .A(n10153), .ZN(n10133) );
  NAND2_X1 U8108 ( .A1(n6316), .A2(n6315), .ZN(P2_U3455) );
  INV_X1 U8109 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6325) );
  XNOR2_X1 U8110 ( .A(n6317), .B(n9259), .ZN(n9607) );
  NAND2_X1 U8111 ( .A1(n9384), .A2(n9267), .ZN(n7547) );
  INV_X1 U8112 ( .A(n6318), .ZN(n9624) );
  INV_X1 U8113 ( .A(n6362), .ZN(n6319) );
  AOI211_X1 U8114 ( .C1(n8981), .C2(n9624), .A(n9832), .B(n6319), .ZN(n9608)
         );
  OAI211_X1 U8115 ( .C1(n6321), .C2(n9259), .A(n9846), .B(n6320), .ZN(n6324)
         );
  OR2_X1 U8116 ( .A1(n9031), .A2(n9810), .ZN(n6323) );
  NAND2_X1 U8117 ( .A1(n9456), .A2(n9841), .ZN(n6322) );
  AND2_X1 U8118 ( .A1(n6323), .A2(n6322), .ZN(n8977) );
  NAND2_X1 U8119 ( .A1(n6324), .A2(n8977), .ZN(n9614) );
  AOI211_X1 U8120 ( .C1(n9607), .C2(n10113), .A(n9608), .B(n9614), .ZN(n9867)
         );
  MUX2_X1 U8121 ( .A(n6325), .B(n9867), .S(n10348), .Z(n6328) );
  NAND2_X1 U8122 ( .A1(n8981), .A2(n6326), .ZN(n6327) );
  NAND2_X1 U8123 ( .A1(n6328), .A2(n6327), .ZN(P1_U3517) );
  INV_X1 U8124 ( .A(n8519), .ZN(n8078) );
  INV_X1 U8125 ( .A(n8505), .ZN(n8239) );
  NAND2_X1 U8126 ( .A1(n8815), .A2(n4560), .ZN(n6331) );
  INV_X1 U8127 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8817) );
  OR2_X1 U8128 ( .A1(n4474), .A2(n8817), .ZN(n6330) );
  NAND2_X1 U8129 ( .A1(n6331), .A2(n6330), .ZN(n6419) );
  OR2_X2 U8130 ( .A1(n6419), .A2(n7818), .ZN(n8233) );
  NAND2_X1 U8131 ( .A1(n6419), .A2(n7818), .ZN(n8032) );
  OAI211_X1 U8132 ( .C1(n8239), .C2(n8078), .A(n8227), .B(n6337), .ZN(n6342)
         );
  INV_X1 U8133 ( .A(n8227), .ZN(n6334) );
  NOR2_X1 U8134 ( .A1(n8505), .A2(n8519), .ZN(n6339) );
  INV_X1 U8135 ( .A(n6339), .ZN(n6333) );
  NAND3_X1 U8136 ( .A1(n6343), .A2(n6334), .A3(n6333), .ZN(n6341) );
  INV_X1 U8137 ( .A(n6337), .ZN(n6335) );
  OAI21_X1 U8138 ( .B1(n6335), .B2(n8519), .A(n8505), .ZN(n6336) );
  OAI211_X1 U8139 ( .C1(n8078), .C2(n6337), .A(n6334), .B(n6336), .ZN(n6338)
         );
  OAI21_X1 U8140 ( .B1(n6334), .B2(n6339), .A(n6338), .ZN(n6340) );
  OAI211_X1 U8141 ( .C1(n6343), .C2(n6342), .A(n6341), .B(n6340), .ZN(n6344)
         );
  INV_X1 U8142 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8143 ( .A1(n4295), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6347) );
  INV_X1 U8144 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6345) );
  OR2_X1 U8145 ( .A1(n8022), .A2(n6345), .ZN(n6346) );
  OAI211_X1 U8146 ( .C1(n5957), .C2(n6348), .A(n6347), .B(n6346), .ZN(n6349)
         );
  INV_X1 U8147 ( .A(n6349), .ZN(n6350) );
  NAND2_X1 U8148 ( .A1(n8027), .A2(n6350), .ZN(n8258) );
  AOI21_X1 U8149 ( .B1(P2_B_REG_SCAN_IN), .B2(n5858), .A(n8658), .ZN(n8497) );
  AOI22_X1 U8150 ( .A1(n8573), .A2(n8519), .B1(n8258), .B2(n8497), .ZN(n6351)
         );
  OR2_X1 U8151 ( .A1(n7752), .A2(n10127), .ZN(n6352) );
  NAND2_X1 U8152 ( .A1(n7760), .A2(n6352), .ZN(n6418) );
  NAND2_X1 U8153 ( .A1(n6418), .A2(n10155), .ZN(n6355) );
  NOR2_X2 U8154 ( .A1(n10156), .A2(n10150), .ZN(n8801) );
  NAND2_X1 U8155 ( .A1(n6355), .A2(n6354), .ZN(P2_U3456) );
  NAND2_X1 U8156 ( .A1(n6356), .A2(n9262), .ZN(n6357) );
  OAI211_X1 U8157 ( .C1(n6359), .C2(n9262), .A(n6358), .B(n9846), .ZN(n6361)
         );
  OAI22_X1 U8158 ( .A1(n9199), .A2(n9808), .B1(n7022), .B2(n9810), .ZN(n6360)
         );
  INV_X1 U8159 ( .A(n6360), .ZN(n9043) );
  NAND2_X1 U8160 ( .A1(n6361), .A2(n9043), .ZN(n7749) );
  AOI21_X1 U8161 ( .B1(n6362), .B2(n9045), .A(n9832), .ZN(n6363) );
  AND2_X1 U8162 ( .A1(n6363), .A2(n4374), .ZN(n7745) );
  NOR2_X1 U8163 ( .A1(n7749), .A2(n7745), .ZN(n6364) );
  NAND2_X1 U8164 ( .A1(n6368), .A2(n10348), .ZN(n6367) );
  AOI21_X1 U8165 ( .B1(n10346), .B2(P1_REG0_REG_28__SCAN_IN), .A(n6365), .ZN(
        n6366) );
  NAND2_X1 U8166 ( .A1(n6367), .A2(n6366), .ZN(P1_U3518) );
  NAND2_X1 U8167 ( .A1(n6368), .A2(n10117), .ZN(n6373) );
  INV_X1 U8168 ( .A(n9899), .ZN(n6370) );
  NAND2_X1 U8169 ( .A1(n10118), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6369) );
  INV_X1 U8170 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U8171 ( .A1(n6373), .A2(n6372), .ZN(P1_U3550) );
  OR2_X1 U8172 ( .A1(n9370), .A2(n9943), .ZN(n6374) );
  INV_X1 U8173 ( .A(n6377), .ZN(n6375) );
  NOR2_X1 U8174 ( .A1(n6375), .A2(n9943), .ZN(n6376) );
  AND2_X1 U8175 ( .A1(n9370), .A2(n6376), .ZN(n6380) );
  OR3_X1 U8176 ( .A1(n9370), .A2(n9943), .A3(n6377), .ZN(n6378) );
  INV_X1 U8177 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U8178 ( .A1(n10118), .A2(n6385), .ZN(n6386) );
  OAI21_X1 U8179 ( .B1(n6412), .B2(n10118), .A(n6386), .ZN(n6388) );
  NAND2_X1 U8180 ( .A1(n6388), .A2(n6387), .ZN(P1_U3551) );
  INV_X1 U8181 ( .A(n6390), .ZN(n6391) );
  NAND2_X1 U8182 ( .A1(n6389), .A2(n6391), .ZN(n8552) );
  INV_X1 U8183 ( .A(n8551), .ZN(n6392) );
  AND2_X1 U8184 ( .A1(n8552), .A2(n6392), .ZN(n6394) );
  AND2_X1 U8185 ( .A1(n6392), .A2(n8212), .ZN(n6393) );
  NAND2_X1 U8186 ( .A1(n8552), .A2(n6393), .ZN(n8539) );
  INV_X1 U8187 ( .A(n8760), .ZN(n6407) );
  INV_X1 U8188 ( .A(n8762), .ZN(n8531) );
  NOR2_X1 U8189 ( .A1(n8531), .A2(n8671), .ZN(n6400) );
  OR2_X1 U8190 ( .A1(n6400), .A2(n4995), .ZN(n6406) );
  INV_X1 U8191 ( .A(n6401), .ZN(n6402) );
  OAI21_X1 U8192 ( .B1(n8808), .B2(n6848), .A(n6402), .ZN(n6403) );
  XNOR2_X1 U8193 ( .A(n6408), .B(n8212), .ZN(n8763) );
  NAND2_X1 U8194 ( .A1(n8245), .A2(n6213), .ZN(n6924) );
  NAND2_X1 U8195 ( .A1(n7648), .A2(n6924), .ZN(n6409) );
  AOI22_X1 U8196 ( .A1(n8763), .A2(n8678), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8681), .ZN(n6410) );
  NAND2_X1 U8197 ( .A1(n6412), .A2(n10348), .ZN(n6417) );
  NOR2_X1 U8198 ( .A1(n10348), .A2(n10311), .ZN(n6414) );
  NAND2_X1 U8199 ( .A1(n6417), .A2(n6416), .ZN(P1_U3519) );
  NAND2_X1 U8200 ( .A1(n6418), .A2(n10168), .ZN(n6424) );
  INV_X1 U8201 ( .A(n6419), .ZN(n7755) );
  NOR2_X1 U8202 ( .A1(n10168), .A2(n6420), .ZN(n6421) );
  NAND2_X1 U8203 ( .A1(n6424), .A2(n6423), .ZN(P2_U3488) );
  NOR2_X1 U8204 ( .A1(n6677), .A2(P1_U3086), .ZN(n6425) );
  INV_X1 U8205 ( .A(n6486), .ZN(n6426) );
  NAND2_X1 U8206 ( .A1(n8222), .A2(n6813), .ZN(n6427) );
  NAND2_X1 U8207 ( .A1(n6427), .A2(n7392), .ZN(n6579) );
  NAND2_X1 U8208 ( .A1(n6579), .A2(n5858), .ZN(n6428) );
  NAND2_X1 U8209 ( .A1(n6428), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  INV_X1 U8210 ( .A(n6429), .ZN(n6440) );
  AOI22_X1 U8211 ( .A1(n6548), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n9990), .ZN(n6431) );
  OAI21_X1 U8212 ( .B1(n6440), .B2(n9993), .A(n6431), .ZN(P1_U3351) );
  AOI22_X1 U8213 ( .A1(n9514), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9990), .ZN(n6432) );
  OAI21_X1 U8214 ( .B1(n6436), .B2(n9993), .A(n6432), .ZN(P1_U3349) );
  INV_X1 U8215 ( .A(n9990), .ZN(n9995) );
  INV_X1 U8216 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6433) );
  OAI222_X1 U8217 ( .A1(n9995), .A2(n6433), .B1(n9993), .B2(n6461), .C1(n6509), 
        .C2(P1_U3086), .ZN(P1_U3354) );
  INV_X1 U8218 ( .A(n6887), .ZN(n6966) );
  NAND2_X1 U8219 ( .A1(n4543), .A2(P2_U3151), .ZN(n8822) );
  INV_X2 U8220 ( .A(n8820), .ZN(n8816) );
  OAI222_X1 U8221 ( .A1(P2_U3151), .A2(n6966), .B1(n8822), .B2(n6455), .C1(
        n5097), .C2(n8816), .ZN(P2_U3290) );
  OAI222_X1 U8222 ( .A1(n8816), .A2(n6434), .B1(n8822), .B2(n6458), .C1(n6762), 
        .C2(P2_U3151), .ZN(P2_U3292) );
  INV_X1 U8223 ( .A(n7095), .ZN(n7088) );
  INV_X1 U8224 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6435) );
  OAI222_X1 U8225 ( .A1(P2_U3151), .A2(n7088), .B1(n8822), .B2(n6436), .C1(
        n6435), .C2(n8816), .ZN(P2_U3289) );
  INV_X1 U8226 ( .A(n6437), .ZN(n6451) );
  OAI222_X1 U8227 ( .A1(n8816), .A2(n6438), .B1(n8822), .B2(n6451), .C1(
        P2_U3151), .C2(n6659), .ZN(P2_U3293) );
  INV_X1 U8228 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6439) );
  OAI222_X1 U8229 ( .A1(P2_U3151), .A2(n6881), .B1(n8822), .B2(n6440), .C1(
        n6439), .C2(n8816), .ZN(P2_U3291) );
  INV_X1 U8230 ( .A(n6441), .ZN(n6447) );
  OAI222_X1 U8231 ( .A1(P2_U3151), .A2(n7098), .B1(n8822), .B2(n6447), .C1(
        n10205), .C2(n8816), .ZN(P2_U3288) );
  INV_X1 U8232 ( .A(n6442), .ZN(n6444) );
  AOI22_X1 U8233 ( .A1(n9540), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n9990), .ZN(n6443) );
  OAI21_X1 U8234 ( .B1(n6444), .B2(n9993), .A(n6443), .ZN(P1_U3347) );
  INV_X1 U8235 ( .A(n7297), .ZN(n7306) );
  OAI222_X1 U8236 ( .A1(n8816), .A2(n5151), .B1(n8822), .B2(n6444), .C1(
        P2_U3151), .C2(n7306), .ZN(P2_U3287) );
  AOI22_X1 U8237 ( .A1(n6779), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9990), .ZN(n6445) );
  OAI21_X1 U8238 ( .B1(n6465), .B2(n9993), .A(n6445), .ZN(P1_U3345) );
  INV_X1 U8239 ( .A(n9993), .ZN(n7395) );
  AOI22_X1 U8240 ( .A1(n9527), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9990), .ZN(n6446) );
  OAI21_X1 U8241 ( .B1(n6447), .B2(n9993), .A(n6446), .ZN(P1_U3348) );
  INV_X1 U8242 ( .A(n6448), .ZN(n9449) );
  OR2_X1 U8243 ( .A1(n6678), .A2(n10066), .ZN(n9452) );
  NAND2_X1 U8244 ( .A1(n9449), .A2(n9452), .ZN(n6468) );
  AOI21_X1 U8245 ( .B1(n9237), .B2(n6678), .A(n6449), .ZN(n6467) );
  INV_X1 U8246 ( .A(n6467), .ZN(n6450) );
  AND2_X1 U8247 ( .A1(n6468), .A2(n6450), .ZN(n10033) );
  NOR2_X1 U8248 ( .A1(n10033), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8249 ( .A(n6530), .ZN(n6452) );
  OAI222_X1 U8250 ( .A1(n10066), .A2(n6452), .B1(n9993), .B2(n6451), .C1(n9995), .C2(n5044), .ZN(P1_U3353) );
  INV_X1 U8251 ( .A(n6453), .ZN(n6463) );
  OAI222_X1 U8252 ( .A1(n9995), .A2(n6454), .B1(n9993), .B2(n6463), .C1(n6636), 
        .C2(n10066), .ZN(P1_U3346) );
  INV_X1 U8253 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6456) );
  OAI222_X1 U8254 ( .A1(n9995), .A2(n6456), .B1(n9993), .B2(n6455), .C1(n6551), 
        .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U8255 ( .A(n9488), .ZN(n6457) );
  OAI222_X1 U8256 ( .A1(n9995), .A2(n6459), .B1(n9993), .B2(n6458), .C1(n6457), 
        .C2(n10066), .ZN(P1_U3352) );
  INV_X1 U8257 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10258) );
  NOR2_X1 U8258 ( .A1(n6484), .A2(n10258), .ZN(P2_U3239) );
  INV_X1 U8259 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U8260 ( .A1(n6484), .A2(n10234), .ZN(P2_U3234) );
  INV_X1 U8261 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8262 ( .A1(n9075), .A2(P1_U3973), .ZN(n6460) );
  OAI21_X1 U8263 ( .B1(n6567), .B2(P1_U3973), .A(n6460), .ZN(P1_U3567) );
  INV_X1 U8264 ( .A(n8822), .ZN(n7391) );
  INV_X1 U8265 ( .A(n7391), .ZN(n7670) );
  OAI222_X1 U8266 ( .A1(n8816), .A2(n5039), .B1(n7670), .B2(n6461), .C1(n6606), 
        .C2(P2_U3151), .ZN(P2_U3294) );
  OAI222_X1 U8267 ( .A1(P2_U3151), .A2(n7300), .B1(n7670), .B2(n6463), .C1(
        n6462), .C2(n8816), .ZN(P2_U3286) );
  INV_X1 U8268 ( .A(n8295), .ZN(n8279) );
  INV_X1 U8269 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6464) );
  OAI222_X1 U8270 ( .A1(P2_U3151), .A2(n8279), .B1(n7670), .B2(n6465), .C1(
        n6464), .C2(n8816), .ZN(P2_U3285) );
  NAND2_X1 U8271 ( .A1(n9376), .A2(P1_U3973), .ZN(n6466) );
  OAI21_X1 U8272 ( .B1(P1_U3973), .B2(n8028), .A(n6466), .ZN(P1_U3585) );
  INV_X1 U8273 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U8274 ( .A1(n6468), .A2(n6467), .ZN(n6518) );
  INV_X1 U8275 ( .A(n6518), .ZN(n6471) );
  INV_X1 U8276 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10097) );
  AOI21_X1 U8277 ( .B1(n6514), .B2(n10097), .A(n7763), .ZN(n6499) );
  OAI21_X1 U8278 ( .B1(n6514), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6499), .ZN(
        n6469) );
  XNOR2_X1 U8279 ( .A(n6469), .B(n4469), .ZN(n6470) );
  AOI22_X1 U8280 ( .A1(n6471), .A2(n6470), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10066), .ZN(n6472) );
  OAI21_X1 U8281 ( .B1(n10070), .B2(n6473), .A(n6472), .ZN(P1_U3243) );
  INV_X1 U8282 ( .A(n6474), .ZN(n6479) );
  AOI22_X1 U8283 ( .A1(n9559), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9990), .ZN(n6475) );
  OAI21_X1 U8284 ( .B1(n6479), .B2(n9993), .A(n6475), .ZN(P1_U3344) );
  NAND2_X1 U8285 ( .A1(n6476), .A2(P2_U3893), .ZN(n6477) );
  OAI21_X1 U8286 ( .B1(P2_U3893), .B2(n5044), .A(n6477), .ZN(P2_U3493) );
  AND2_X1 U8287 ( .A1(n6478), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8288 ( .A1(n6478), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8289 ( .A1(n6478), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8290 ( .A1(n6478), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8291 ( .A1(n6478), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8292 ( .A1(n6478), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8293 ( .A1(n6478), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8294 ( .A1(n6478), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8295 ( .A1(n6478), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8296 ( .A1(n6478), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8297 ( .A1(n6478), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  INV_X1 U8298 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6480) );
  INV_X1 U8299 ( .A(n8305), .ZN(n8298) );
  OAI222_X1 U8300 ( .A1(n8816), .A2(n6480), .B1(n7670), .B2(n6479), .C1(
        P2_U3151), .C2(n8298), .ZN(P2_U3284) );
  INV_X1 U8301 ( .A(n8338), .ZN(n8329) );
  INV_X1 U8302 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6481) );
  OAI222_X1 U8303 ( .A1(P2_U3151), .A2(n8329), .B1(n7670), .B2(n6482), .C1(
        n6481), .C2(n8816), .ZN(P2_U3283) );
  INV_X1 U8304 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6483) );
  INV_X1 U8305 ( .A(n6788), .ZN(n6991) );
  OAI222_X1 U8306 ( .A1(n9995), .A2(n6483), .B1(n9993), .B2(n6482), .C1(n6991), 
        .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U8307 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6488) );
  INV_X1 U8308 ( .A(n6485), .ZN(n6487) );
  AOI22_X1 U8309 ( .A1(n6478), .A2(n6488), .B1(n6487), .B2(n6486), .ZN(
        P2_U3376) );
  AND2_X1 U8310 ( .A1(n6478), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8311 ( .A1(n6478), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8312 ( .A1(n6478), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8313 ( .A1(n6478), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8314 ( .A1(n6478), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8315 ( .A1(n6478), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8316 ( .A1(n6478), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8317 ( .A1(n6478), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8318 ( .A1(n6478), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8319 ( .A1(n6478), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8320 ( .A1(n6478), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8321 ( .A1(n6478), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8322 ( .A1(n6478), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8323 ( .A1(n6478), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8324 ( .A1(n6478), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8325 ( .A1(n6478), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8326 ( .A1(n6478), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  INV_X1 U8327 ( .A(n6489), .ZN(n6568) );
  AOI22_X1 U8328 ( .A1(n9576), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9990), .ZN(n6490) );
  OAI21_X1 U8329 ( .B1(n6568), .B2(n9993), .A(n6490), .ZN(P1_U3342) );
  NAND2_X1 U8330 ( .A1(n4289), .A2(n10090), .ZN(n6492) );
  INV_X1 U8331 ( .A(n6677), .ZN(n6495) );
  NAND2_X1 U8332 ( .A1(n6495), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6494) );
  OAI211_X2 U8333 ( .C1(n4301), .C2(n9443), .A(n7260), .B(n6677), .ZN(n6709)
         );
  INV_X2 U8334 ( .A(n6709), .ZN(n8952) );
  NAND2_X1 U8335 ( .A1(n9474), .A2(n8952), .ZN(n6497) );
  NAND2_X1 U8336 ( .A1(n6497), .A2(n6496), .ZN(n6691) );
  XNOR2_X1 U8337 ( .A(n6692), .B(n6691), .ZN(n6722) );
  NOR2_X1 U8338 ( .A1(n7763), .A2(n6514), .ZN(n6501) );
  INV_X2 U8339 ( .A(P1_U3973), .ZN(n9473) );
  AND2_X1 U8340 ( .A1(n4469), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9476) );
  INV_X1 U8341 ( .A(n9476), .ZN(n6498) );
  OR2_X1 U8342 ( .A1(n7763), .A2(n7708), .ZN(n9448) );
  OAI22_X1 U8343 ( .A1(n6499), .A2(n4469), .B1(n6498), .B2(n9448), .ZN(n6500)
         );
  AOI211_X1 U8344 ( .C1(n6722), .C2(n6501), .A(n9473), .B(n6500), .ZN(n6536)
         );
  MUX2_X1 U8345 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n5524), .S(n6548), .Z(n6506)
         );
  INV_X1 U8346 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7178) );
  XNOR2_X1 U8347 ( .A(n9488), .B(n7178), .ZN(n9494) );
  INV_X1 U8348 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10077) );
  MUX2_X1 U8349 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10077), .S(n6530), .Z(n6526)
         );
  XNOR2_X1 U8350 ( .A(n6509), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9477) );
  NAND2_X1 U8351 ( .A1(n9477), .A2(n9476), .ZN(n9475) );
  NAND2_X1 U8352 ( .A1(n5061), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6502) );
  NAND2_X1 U8353 ( .A1(n9475), .A2(n6502), .ZN(n6525) );
  NAND2_X1 U8354 ( .A1(n6526), .A2(n6525), .ZN(n6524) );
  NAND2_X1 U8355 ( .A1(n6530), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U8356 ( .A1(n6524), .A2(n6503), .ZN(n9493) );
  NAND2_X1 U8357 ( .A1(n9494), .A2(n9493), .ZN(n9492) );
  NAND2_X1 U8358 ( .A1(n9488), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6504) );
  NAND2_X1 U8359 ( .A1(n9492), .A2(n6504), .ZN(n6505) );
  INV_X1 U8360 ( .A(n10060), .ZN(n10048) );
  NAND2_X1 U8361 ( .A1(n6505), .A2(n6506), .ZN(n6538) );
  OAI211_X1 U8362 ( .C1(n6506), .C2(n6505), .A(n10048), .B(n6538), .ZN(n6522)
         );
  INV_X1 U8363 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6507) );
  MUX2_X1 U8364 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6507), .S(n6548), .Z(n6516)
         );
  INV_X1 U8365 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6508) );
  XNOR2_X1 U8366 ( .A(n9488), .B(n6508), .ZN(n9491) );
  XNOR2_X1 U8367 ( .A(n6509), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n9480) );
  AND2_X1 U8368 ( .A1(n4469), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9479) );
  NAND2_X1 U8369 ( .A1(n9480), .A2(n9479), .ZN(n9478) );
  NAND2_X1 U8370 ( .A1(n5061), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U8371 ( .A1(n9478), .A2(n6510), .ZN(n6528) );
  INV_X1 U8372 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6511) );
  MUX2_X1 U8373 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6511), .S(n6530), .Z(n6529)
         );
  NAND2_X1 U8374 ( .A1(n6528), .A2(n6529), .ZN(n6527) );
  NAND2_X1 U8375 ( .A1(n6530), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U8376 ( .A1(n6527), .A2(n6512), .ZN(n9490) );
  NAND2_X1 U8377 ( .A1(n9491), .A2(n9490), .ZN(n9489) );
  NAND2_X1 U8378 ( .A1(n9488), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6513) );
  NAND2_X1 U8379 ( .A1(n9489), .A2(n6513), .ZN(n6515) );
  NAND2_X1 U8380 ( .A1(n6515), .A2(n6516), .ZN(n6550) );
  OAI211_X1 U8381 ( .C1(n6516), .C2(n6515), .A(n10047), .B(n6550), .ZN(n6521)
         );
  AND2_X1 U8382 ( .A1(n10066), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9120) );
  AOI21_X1 U8383 ( .B1(n10033), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n9120), .ZN(
        n6520) );
  NAND2_X1 U8384 ( .A1(n4409), .A2(n6548), .ZN(n6519) );
  NAND4_X1 U8385 ( .A1(n6522), .A2(n6521), .A3(n6520), .A4(n6519), .ZN(n6523)
         );
  OR2_X1 U8386 ( .A1(n6536), .A2(n6523), .ZN(P1_U3247) );
  OAI211_X1 U8387 ( .C1(n6526), .C2(n6525), .A(n10048), .B(n6524), .ZN(n6534)
         );
  AOI22_X1 U8388 ( .A1(n10033), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10066), .ZN(n6533) );
  OAI211_X1 U8389 ( .C1(n6529), .C2(n6528), .A(n10047), .B(n6527), .ZN(n6532)
         );
  NAND2_X1 U8390 ( .A1(n4409), .A2(n6530), .ZN(n6531) );
  NAND4_X1 U8391 ( .A1(n6534), .A2(n6533), .A3(n6532), .A4(n6531), .ZN(n6535)
         );
  OR2_X1 U8392 ( .A1(n6536), .A2(n6535), .ZN(P1_U3245) );
  INV_X1 U8393 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6635) );
  XNOR2_X1 U8394 ( .A(n6636), .B(n6635), .ZN(n6546) );
  NAND2_X1 U8395 ( .A1(n6548), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8396 ( .A1(n6538), .A2(n6537), .ZN(n9506) );
  XNOR2_X1 U8397 ( .A(n6551), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n9507) );
  NAND2_X1 U8398 ( .A1(n9506), .A2(n9507), .ZN(n9505) );
  NAND2_X1 U8399 ( .A1(n9501), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8400 ( .A1(n9505), .A2(n6539), .ZN(n9516) );
  INV_X1 U8401 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7342) );
  MUX2_X1 U8402 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7342), .S(n9514), .Z(n9517)
         );
  NAND2_X1 U8403 ( .A1(n9516), .A2(n9517), .ZN(n9515) );
  NAND2_X1 U8404 ( .A1(n9514), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6540) );
  NAND2_X1 U8405 ( .A1(n9515), .A2(n6540), .ZN(n9529) );
  INV_X1 U8406 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6541) );
  XNOR2_X1 U8407 ( .A(n9527), .B(n6541), .ZN(n9530) );
  NAND2_X1 U8408 ( .A1(n9529), .A2(n9530), .ZN(n9528) );
  NAND2_X1 U8409 ( .A1(n9527), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6542) );
  NAND2_X1 U8410 ( .A1(n9528), .A2(n6542), .ZN(n9542) );
  INV_X1 U8411 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n9854) );
  XNOR2_X1 U8412 ( .A(n9540), .B(n9854), .ZN(n9543) );
  NAND2_X1 U8413 ( .A1(n9542), .A2(n9543), .ZN(n9541) );
  NAND2_X1 U8414 ( .A1(n9540), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6543) );
  NAND2_X1 U8415 ( .A1(n9541), .A2(n6543), .ZN(n6545) );
  INV_X1 U8416 ( .A(n6638), .ZN(n6544) );
  AOI21_X1 U8417 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6566) );
  INV_X1 U8418 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n6547) );
  NAND2_X1 U8419 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n9134) );
  OAI21_X1 U8420 ( .B1(n10070), .B2(n6547), .A(n9134), .ZN(n6563) );
  NAND2_X1 U8421 ( .A1(n6548), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U8422 ( .A1(n6550), .A2(n6549), .ZN(n9503) );
  XNOR2_X1 U8423 ( .A(n6551), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9504) );
  NAND2_X1 U8424 ( .A1(n9503), .A2(n9504), .ZN(n9502) );
  NAND2_X1 U8425 ( .A1(n9501), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6552) );
  NAND2_X1 U8426 ( .A1(n9502), .A2(n6552), .ZN(n9519) );
  INV_X1 U8427 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U8428 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6553), .S(n9514), .Z(n9520)
         );
  NAND2_X1 U8429 ( .A1(n9519), .A2(n9520), .ZN(n9518) );
  NAND2_X1 U8430 ( .A1(n9514), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6554) );
  NAND2_X1 U8431 ( .A1(n9518), .A2(n6554), .ZN(n9532) );
  INV_X1 U8432 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6555) );
  XNOR2_X1 U8433 ( .A(n9527), .B(n6555), .ZN(n9533) );
  NAND2_X1 U8434 ( .A1(n9532), .A2(n9533), .ZN(n9531) );
  NAND2_X1 U8435 ( .A1(n9527), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U8436 ( .A1(n9531), .A2(n6556), .ZN(n9546) );
  INV_X1 U8437 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6557) );
  XNOR2_X1 U8438 ( .A(n9540), .B(n6557), .ZN(n9545) );
  NAND2_X1 U8439 ( .A1(n9546), .A2(n9545), .ZN(n9544) );
  NAND2_X1 U8440 ( .A1(n9540), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U8441 ( .A1(n9544), .A2(n6558), .ZN(n6560) );
  INV_X1 U8442 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6629) );
  XNOR2_X1 U8443 ( .A(n6636), .B(n6629), .ZN(n6559) );
  NAND2_X1 U8444 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  AOI21_X1 U8445 ( .B1(n6631), .B2(n6561), .A(n10055), .ZN(n6562) );
  AOI211_X1 U8446 ( .C1(n4409), .C2(n6564), .A(n6563), .B(n6562), .ZN(n6565)
         );
  OAI21_X1 U8447 ( .B1(n6566), .B2(n10060), .A(n6565), .ZN(P1_U3252) );
  INV_X1 U8448 ( .A(n8355), .ZN(n8341) );
  OAI222_X1 U8449 ( .A1(P2_U3151), .A2(n8341), .B1(n7670), .B2(n6568), .C1(
        n8816), .C2(n6567), .ZN(P2_U3282) );
  NAND2_X1 U8450 ( .A1(n6579), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6569) );
  MUX2_X1 U8451 ( .A(n8457), .B(n6569), .S(n6578), .Z(n6571) );
  INV_X1 U8452 ( .A(n7392), .ZN(n6572) );
  NOR2_X1 U8453 ( .A1(n6813), .A2(n6572), .ZN(n6573) );
  NOR2_X1 U8454 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5870), .ZN(n6577) );
  INV_X1 U8455 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U8456 ( .A1(n6598), .A2(n6603), .ZN(n6597) );
  AOI211_X1 U8457 ( .C1(n6575), .C2(n6597), .A(n8482), .B(n6608), .ZN(n6576)
         );
  AOI211_X1 U8458 ( .C1(n8484), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6577), .B(
        n6576), .ZN(n6592) );
  NOR2_X1 U8459 ( .A1(n6578), .A2(P2_U3151), .ZN(n8819) );
  INV_X1 U8460 ( .A(n6606), .ZN(n6581) );
  NAND2_X1 U8461 ( .A1(n6603), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6580) );
  AND2_X1 U8462 ( .A1(n6585), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6611) );
  NAND2_X1 U8463 ( .A1(n6582), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6613) );
  OAI21_X1 U8464 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(n6582), .A(n6613), .ZN(
        n6590) );
  INV_X1 U8465 ( .A(n6596), .ZN(n6583) );
  INV_X1 U8466 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7137) );
  NOR2_X1 U8467 ( .A1(n6584), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6586) );
  NAND2_X1 U8468 ( .A1(n6585), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6618) );
  AOI21_X1 U8469 ( .B1(n7137), .B2(n6587), .A(n6620), .ZN(n6588) );
  NOR2_X1 U8470 ( .A1(n8495), .A2(n6588), .ZN(n6589) );
  AOI21_X1 U8471 ( .B1(n8492), .B2(n6590), .A(n6589), .ZN(n6591) );
  OAI211_X1 U8472 ( .C1(n6606), .C2(n8488), .A(n6592), .B(n6591), .ZN(P2_U3183) );
  INV_X1 U8473 ( .A(n6593), .ZN(n6604) );
  AOI22_X1 U8474 ( .A1(n10006), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n9990), .ZN(n6594) );
  OAI21_X1 U8475 ( .B1(n6604), .B2(n9993), .A(n6594), .ZN(P1_U3341) );
  MUX2_X1 U8476 ( .A(n6726), .B(n8637), .S(P2_U3893), .Z(n6595) );
  INV_X1 U8477 ( .A(n6595), .ZN(P2_U3508) );
  INV_X1 U8478 ( .A(n8482), .ZN(n8436) );
  NOR2_X1 U8479 ( .A1(n6596), .A2(n8436), .ZN(n6600) );
  AOI21_X1 U8480 ( .B1(n6598), .B2(n6603), .A(n6597), .ZN(n6599) );
  OAI22_X1 U8481 ( .A1(n6600), .A2(n6599), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6843), .ZN(n6601) );
  AOI21_X1 U8482 ( .B1(n8484), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n6601), .ZN(
        n6602) );
  OAI21_X1 U8483 ( .B1(n6603), .B2(n8488), .A(n6602), .ZN(P2_U3182) );
  INV_X1 U8484 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6605) );
  INV_X1 U8485 ( .A(n8378), .ZN(n8391) );
  OAI222_X1 U8486 ( .A1(n8816), .A2(n6605), .B1(n7670), .B2(n6604), .C1(
        P2_U3151), .C2(n8391), .ZN(P2_U3281) );
  MUX2_X1 U8487 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6214), .Z(n6648) );
  XNOR2_X1 U8488 ( .A(n6648), .B(n6659), .ZN(n6609) );
  AOI211_X1 U8489 ( .C1(n6610), .C2(n6609), .A(n8482), .B(n6647), .ZN(n6627)
         );
  INV_X1 U8490 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10331) );
  XNOR2_X1 U8491 ( .A(n6659), .B(n10331), .ZN(n6615) );
  INV_X1 U8492 ( .A(n6611), .ZN(n6612) );
  NAND2_X1 U8493 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  NAND2_X1 U8494 ( .A1(n6614), .A2(n6615), .ZN(n6661) );
  OAI21_X1 U8495 ( .B1(n6615), .B2(n6614), .A(n6661), .ZN(n6616) );
  NAND2_X1 U8496 ( .A1(n8492), .A2(n6616), .ZN(n6617) );
  OAI21_X1 U8497 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n5850), .A(n6617), .ZN(n6626) );
  INV_X1 U8498 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6624) );
  XNOR2_X1 U8499 ( .A(n6659), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6622) );
  INV_X1 U8500 ( .A(n6618), .ZN(n6619) );
  NOR2_X1 U8501 ( .A1(n6620), .A2(n6619), .ZN(n6621) );
  NOR2_X1 U8502 ( .A1(n6621), .A2(n6622), .ZN(n6653) );
  AOI21_X1 U8503 ( .B1(n6622), .B2(n6621), .A(n6653), .ZN(n6623) );
  OAI22_X1 U8504 ( .A1(n8371), .A2(n6624), .B1(n8495), .B2(n6623), .ZN(n6625)
         );
  NOR3_X1 U8505 ( .A1(n6627), .A2(n6626), .A3(n6625), .ZN(n6628) );
  OAI21_X1 U8506 ( .B1(n6659), .B2(n8488), .A(n6628), .ZN(P2_U3184) );
  XNOR2_X1 U8507 ( .A(n6779), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U8508 ( .A1(n6636), .A2(n6629), .ZN(n6630) );
  NAND2_X1 U8509 ( .A1(n6631), .A2(n6630), .ZN(n6633) );
  INV_X1 U8510 ( .A(n6771), .ZN(n6632) );
  AOI211_X1 U8511 ( .C1(n6634), .C2(n6633), .A(n10055), .B(n6632), .ZN(n6646)
         );
  XNOR2_X1 U8512 ( .A(n6779), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U8513 ( .A1(n6636), .A2(n6635), .ZN(n6637) );
  NAND2_X1 U8514 ( .A1(n6638), .A2(n6637), .ZN(n6640) );
  INV_X1 U8515 ( .A(n6781), .ZN(n6639) );
  AOI211_X1 U8516 ( .C1(n6641), .C2(n6640), .A(n10060), .B(n6639), .ZN(n6645)
         );
  INV_X1 U8517 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U8518 ( .A1(n4409), .A2(n6779), .ZN(n6642) );
  NAND2_X1 U8519 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9016) );
  OAI211_X1 U8520 ( .C1(n6643), .C2(n10070), .A(n6642), .B(n9016), .ZN(n6644)
         );
  OR3_X1 U8521 ( .A1(n6646), .A2(n6645), .A3(n6644), .ZN(P1_U3253) );
  MUX2_X1 U8522 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8405), .Z(n6763) );
  XOR2_X1 U8523 ( .A(n6762), .B(n6763), .Z(n6649) );
  OAI21_X1 U8524 ( .B1(n6650), .B2(n6649), .A(n6761), .ZN(n6651) );
  NAND2_X1 U8525 ( .A1(n6651), .A2(n8436), .ZN(n6669) );
  INV_X1 U8526 ( .A(n8495), .ZN(n8345) );
  NOR2_X1 U8527 ( .A1(n6653), .A2(n6652), .ZN(n6655) );
  INV_X1 U8528 ( .A(n6762), .ZN(n6654) );
  NOR2_X1 U8529 ( .A1(n6655), .A2(n6654), .ZN(n6752) );
  NAND2_X1 U8530 ( .A1(n6657), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6753) );
  OAI21_X1 U8531 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n6657), .A(n6753), .ZN(
        n6658) );
  AOI22_X1 U8532 ( .A1(n8484), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(n8345), .B2(
        n6658), .ZN(n6667) );
  NAND2_X1 U8533 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U8534 ( .A1(n6659), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8535 ( .A1(n6661), .A2(n6660), .ZN(n6662) );
  NAND2_X1 U8536 ( .A1(n6662), .A2(n6762), .ZN(n6747) );
  OR2_X1 U8537 ( .A1(n6662), .A2(n6762), .ZN(n6663) );
  OAI21_X1 U8538 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n6664), .A(n6750), .ZN(
        n6665) );
  NAND2_X1 U8539 ( .A1(n8492), .A2(n6665), .ZN(n6666) );
  AND3_X1 U8540 ( .A1(n6667), .A2(n6889), .A3(n6666), .ZN(n6668) );
  OAI211_X1 U8541 ( .C1(n8488), .C2(n6762), .A(n6669), .B(n6668), .ZN(P2_U3185) );
  INV_X1 U8542 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U8543 ( .A1(n9474), .A2(n7265), .ZN(n9400) );
  NAND2_X1 U8544 ( .A1(n7254), .A2(n9400), .ZN(n10087) );
  OAI21_X1 U8545 ( .B1(n9846), .B2(n10113), .A(n10087), .ZN(n6670) );
  OR2_X1 U8546 ( .A1(n5509), .A2(n9810), .ZN(n10092) );
  OAI211_X1 U8547 ( .C1(n7265), .C2(n10085), .A(n6670), .B(n10092), .ZN(n9945)
         );
  NAND2_X1 U8548 ( .A1(n9945), .A2(n10348), .ZN(n6671) );
  OAI21_X1 U8549 ( .B1(n10348), .B2(n10262), .A(n6671), .ZN(P1_U3453) );
  OAI211_X1 U8550 ( .C1(n6675), .C2(n6674), .A(n6673), .B(n6672), .ZN(n6695)
         );
  INV_X1 U8551 ( .A(n9940), .ZN(n10110) );
  NAND2_X1 U8552 ( .A1(n6695), .A2(n10110), .ZN(n6680) );
  INV_X1 U8553 ( .A(n6676), .ZN(n6679) );
  NAND4_X1 U8554 ( .A1(n6680), .A2(n6679), .A3(n6678), .A4(n6677), .ZN(n6681)
         );
  NAND2_X1 U8555 ( .A1(n6681), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6683) );
  NAND3_X1 U8556 ( .A1(n6695), .A2(n6699), .A3(P1_STATE_REG_SCAN_IN), .ZN(
        n6682) );
  NAND2_X1 U8557 ( .A1(n9210), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6719) );
  INV_X1 U8558 ( .A(n6719), .ZN(n6706) );
  INV_X1 U8559 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7266) );
  NAND2_X4 U8560 ( .A1(n6688), .A2(n9394), .ZN(n8964) );
  XNOR2_X1 U8561 ( .A(n6689), .B(n8964), .ZN(n6712) );
  OAI22_X1 U8562 ( .A1(n5509), .A2(n6709), .B1(n10101), .B2(n4293), .ZN(n6710)
         );
  XNOR2_X1 U8563 ( .A(n6712), .B(n6710), .ZN(n6694) );
  NOR2_X1 U8564 ( .A1(n6694), .A2(n6693), .ZN(n6697) );
  NOR2_X1 U8565 ( .A1(n6695), .A2(n9449), .ZN(n6698) );
  NOR2_X1 U8566 ( .A1(n9940), .A2(n9237), .ZN(n6696) );
  OAI21_X1 U8567 ( .B1(n6697), .B2(n6714), .A(n9196), .ZN(n6705) );
  INV_X1 U8568 ( .A(n6698), .ZN(n6701) );
  OR2_X1 U8569 ( .A1(n6701), .A2(n9443), .ZN(n9167) );
  NAND2_X1 U8570 ( .A1(n9202), .A2(n9841), .ZN(n9212) );
  INV_X1 U8571 ( .A(n9212), .ZN(n9015) );
  NAND2_X1 U8572 ( .A1(n9202), .A2(n9843), .ZN(n9209) );
  INV_X1 U8573 ( .A(n6699), .ZN(n6700) );
  OR2_X1 U8574 ( .A1(n6701), .A2(n6700), .ZN(n6702) );
  OAI22_X1 U8575 ( .A1(n9209), .A2(n5518), .B1(n9205), .B2(n10101), .ZN(n6703)
         );
  AOI21_X1 U8576 ( .B1(n9015), .B2(n9474), .A(n6703), .ZN(n6704) );
  OAI211_X1 U8577 ( .C1(n6706), .C2(n7266), .A(n6705), .B(n6704), .ZN(P1_U3222) );
  NAND2_X1 U8578 ( .A1(n10073), .A2(n4289), .ZN(n6707) );
  OAI21_X1 U8579 ( .B1(n5518), .B2(n4293), .A(n6707), .ZN(n6708) );
  XNOR2_X1 U8580 ( .A(n6708), .B(n9034), .ZN(n6732) );
  OAI22_X1 U8581 ( .A1(n5518), .A2(n8947), .B1(n6801), .B2(n4293), .ZN(n6731)
         );
  INV_X1 U8582 ( .A(n6710), .ZN(n6711) );
  XOR2_X1 U8583 ( .A(n6734), .B(n6733), .Z(n6718) );
  AOI22_X1 U8584 ( .A1(n9843), .A2(n9471), .B1(n6715), .B2(n9841), .ZN(n6796)
         );
  OAI22_X1 U8585 ( .A1(n9205), .A2(n6801), .B1(n6796), .B2(n9167), .ZN(n6716)
         );
  AOI21_X1 U8586 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6719), .A(n6716), .ZN(
        n6717) );
  OAI21_X1 U8587 ( .B1(n6718), .B2(n9217), .A(n6717), .ZN(P1_U3237) );
  INV_X1 U8588 ( .A(n9209), .ZN(n9180) );
  AOI22_X1 U8589 ( .A1(n9180), .A2(n6715), .B1(n10090), .B2(n9215), .ZN(n6721)
         );
  NAND2_X1 U8590 ( .A1(n6719), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6720) );
  OAI211_X1 U8591 ( .C1(n6722), .C2(n9217), .A(n6721), .B(n6720), .ZN(P1_U3232) );
  INV_X1 U8592 ( .A(n6723), .ZN(n6725) );
  OAI222_X1 U8593 ( .A1(n8816), .A2(n6724), .B1(n7670), .B2(n6725), .C1(
        P2_U3151), .C2(n4765), .ZN(P2_U3278) );
  INV_X1 U8594 ( .A(n10045), .ZN(n9583) );
  OAI222_X1 U8595 ( .A1(n9995), .A2(n6726), .B1(n9993), .B2(n6725), .C1(n10066), .C2(n9583), .ZN(P1_U3338) );
  INV_X1 U8596 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6728) );
  INV_X1 U8597 ( .A(n6727), .ZN(n6729) );
  INV_X1 U8598 ( .A(n8402), .ZN(n8388) );
  OAI222_X1 U8599 ( .A1(n8816), .A2(n6728), .B1(n7670), .B2(n6729), .C1(
        P2_U3151), .C2(n8388), .ZN(P2_U3280) );
  OAI222_X1 U8600 ( .A1(n9995), .A2(n6730), .B1(n9993), .B2(n6729), .C1(
        P1_U3086), .C2(n10015), .ZN(P1_U3340) );
  OAI22_X1 U8601 ( .A1(n6956), .A2(n4293), .B1(n10111), .B2(n8922), .ZN(n6735)
         );
  XNOR2_X1 U8602 ( .A(n6735), .B(n8964), .ZN(n7037) );
  OAI22_X1 U8603 ( .A1(n6956), .A2(n8947), .B1(n10111), .B2(n4294), .ZN(n7035)
         );
  XNOR2_X1 U8604 ( .A(n7037), .B(n7035), .ZN(n7038) );
  XOR2_X1 U8605 ( .A(n7039), .B(n7038), .Z(n6741) );
  NAND2_X1 U8606 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(n10066), .ZN(n9485) );
  OAI21_X1 U8607 ( .B1(n9205), .B2(n10111), .A(n9485), .ZN(n6738) );
  OAI22_X1 U8608 ( .A1(n6736), .A2(n9209), .B1(n9212), .B2(n5518), .ZN(n6737)
         );
  AOI211_X1 U8609 ( .C1(n6739), .C2(n9165), .A(n6738), .B(n6737), .ZN(n6740)
         );
  OAI21_X1 U8610 ( .B1(n6741), .B2(n9217), .A(n6740), .ZN(P1_U3218) );
  INV_X1 U8611 ( .A(n6742), .ZN(n6745) );
  AOI22_X1 U8612 ( .A1(n8475), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n8820), .ZN(n6743) );
  OAI21_X1 U8613 ( .B1(n6745), .B2(n7670), .A(n6743), .ZN(P2_U3277) );
  AOI22_X1 U8614 ( .A1(n10065), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9990), .ZN(n6744) );
  OAI21_X1 U8615 ( .B1(n6745), .B2(n9993), .A(n6744), .ZN(P1_U3337) );
  INV_X1 U8616 ( .A(n6747), .ZN(n6746) );
  XNOR2_X1 U8617 ( .A(n6881), .B(n10162), .ZN(n6748) );
  NOR2_X1 U8618 ( .A1(n6746), .A2(n6748), .ZN(n6751) );
  INV_X1 U8619 ( .A(n6874), .ZN(n6749) );
  AOI21_X1 U8620 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6760) );
  INV_X1 U8621 ( .A(n8492), .ZN(n7302) );
  INV_X1 U8622 ( .A(n6752), .ZN(n6754) );
  XNOR2_X1 U8623 ( .A(n6881), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6755) );
  AOI21_X1 U8624 ( .B1(n6753), .B2(n6754), .A(n6755), .ZN(n6870) );
  INV_X1 U8625 ( .A(n6870), .ZN(n6757) );
  NAND3_X1 U8626 ( .A1(n6753), .A2(n6755), .A3(n6754), .ZN(n6756) );
  AOI21_X1 U8627 ( .B1(n6757), .B2(n6756), .A(n8495), .ZN(n6758) );
  AOI21_X1 U8628 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(n8484), .A(n6758), .ZN(
        n6759) );
  NAND2_X1 U8629 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6943) );
  OAI211_X1 U8630 ( .C1(n6760), .C2(n7302), .A(n6759), .B(n6943), .ZN(n6767)
         );
  MUX2_X1 U8631 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8405), .Z(n6882) );
  XNOR2_X1 U8632 ( .A(n6882), .B(n6881), .ZN(n6765) );
  AOI211_X1 U8633 ( .C1(n6765), .C2(n6764), .A(n8482), .B(n6880), .ZN(n6766)
         );
  AOI211_X1 U8634 ( .C1(n8373), .C2(n6768), .A(n6767), .B(n6766), .ZN(n6769)
         );
  INV_X1 U8635 ( .A(n6769), .ZN(P2_U3186) );
  XNOR2_X1 U8636 ( .A(n6788), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U8637 ( .A1(n6779), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U8638 ( .A1(n6771), .A2(n6770), .ZN(n9552) );
  INV_X1 U8639 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6772) );
  XNOR2_X1 U8640 ( .A(n9559), .B(n6772), .ZN(n9551) );
  NAND2_X1 U8641 ( .A1(n9552), .A2(n9551), .ZN(n9550) );
  NAND2_X1 U8642 ( .A1(n9559), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6773) );
  NAND2_X1 U8643 ( .A1(n9550), .A2(n6773), .ZN(n6775) );
  INV_X1 U8644 ( .A(n6986), .ZN(n6774) );
  AOI21_X1 U8645 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n6790) );
  INV_X1 U8646 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n6778) );
  AND2_X1 U8647 ( .A1(n10066), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9074) );
  INV_X1 U8648 ( .A(n9074), .ZN(n6777) );
  OAI21_X1 U8649 ( .B1(n10070), .B2(n6778), .A(n6777), .ZN(n6787) );
  NAND2_X1 U8650 ( .A1(n6779), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6780) );
  INV_X1 U8651 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7443) );
  XNOR2_X1 U8652 ( .A(n9559), .B(n7443), .ZN(n9554) );
  NAND2_X1 U8653 ( .A1(n9555), .A2(n9554), .ZN(n9553) );
  NAND2_X1 U8654 ( .A1(n9559), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6782) );
  XNOR2_X1 U8655 ( .A(n6788), .B(P1_REG2_REG_12__SCAN_IN), .ZN(n6783) );
  NAND2_X1 U8656 ( .A1(n6784), .A2(n6783), .ZN(n6785) );
  AOI21_X1 U8657 ( .B1(n6993), .B2(n6785), .A(n10060), .ZN(n6786) );
  AOI211_X1 U8658 ( .C1(n4409), .C2(n6788), .A(n6787), .B(n6786), .ZN(n6789)
         );
  OAI21_X1 U8659 ( .B1(n6790), .B2(n10055), .A(n6789), .ZN(P1_U3255) );
  OR2_X1 U8660 ( .A1(n6791), .A2(n9242), .ZN(n6792) );
  NAND2_X1 U8661 ( .A1(n6793), .A2(n6792), .ZN(n10072) );
  OAI21_X1 U8662 ( .B1(n6801), .B2(n7263), .A(n9782), .ZN(n6794) );
  NOR2_X1 U8663 ( .A1(n6794), .A2(n7177), .ZN(n10075) );
  XOR2_X1 U8664 ( .A(n6795), .B(n9242), .Z(n6798) );
  INV_X1 U8665 ( .A(n6796), .ZN(n6797) );
  AOI21_X1 U8666 ( .B1(n6798), .B2(n9846), .A(n6797), .ZN(n10083) );
  INV_X1 U8667 ( .A(n10083), .ZN(n6799) );
  AOI211_X1 U8668 ( .C1(n10113), .C2(n10072), .A(n10075), .B(n6799), .ZN(n6805) );
  INV_X1 U8669 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6800) );
  OAI22_X1 U8670 ( .A1(n9981), .A2(n6801), .B1(n10348), .B2(n6800), .ZN(n6802)
         );
  INV_X1 U8671 ( .A(n6802), .ZN(n6803) );
  OAI21_X1 U8672 ( .B1(n6805), .B2(n10346), .A(n6803), .ZN(P1_U3459) );
  AOI22_X1 U8673 ( .A1(n9899), .A2(n10073), .B1(n10118), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6804) );
  OAI21_X1 U8674 ( .B1(n6805), .B2(n10118), .A(n6804), .ZN(P1_U3524) );
  INV_X1 U8675 ( .A(n6817), .ZN(n6806) );
  NAND2_X1 U8676 ( .A1(n6858), .A2(n6806), .ZN(n6809) );
  OR2_X1 U8677 ( .A1(n6826), .A2(n6807), .ZN(n6808) );
  INV_X1 U8678 ( .A(n6850), .ZN(n6844) );
  NAND2_X1 U8679 ( .A1(n8278), .A2(n6844), .ZN(n8082) );
  AND2_X1 U8680 ( .A1(n8087), .A2(n8082), .ZN(n8044) );
  INV_X1 U8681 ( .A(n6810), .ZN(n6812) );
  OR2_X1 U8682 ( .A1(n6812), .A2(n6811), .ZN(n6816) );
  AND3_X1 U8683 ( .A1(n6814), .A2(n6813), .A3(n7392), .ZN(n6815) );
  OAI211_X1 U8684 ( .C1(n6819), .C2(n6817), .A(n6816), .B(n6815), .ZN(n6818)
         );
  NAND2_X1 U8685 ( .A1(n6818), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6823) );
  INV_X1 U8686 ( .A(n6819), .ZN(n6821) );
  INV_X1 U8687 ( .A(n6820), .ZN(n8807) );
  NOR2_X1 U8688 ( .A1(n6856), .A2(n8807), .ZN(n8252) );
  NAND2_X1 U8689 ( .A1(n6821), .A2(n8252), .ZN(n6822) );
  NAND2_X1 U8690 ( .A1(n7953), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6867) );
  NAND2_X1 U8691 ( .A1(n6867), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6829) );
  NOR2_X1 U8692 ( .A1(n6856), .A2(n6824), .ZN(n6825) );
  OR2_X1 U8693 ( .A1(n6826), .A2(n10150), .ZN(n6827) );
  AOI22_X1 U8694 ( .A1(n7984), .A2(n8277), .B1(n7998), .B2(n6850), .ZN(n6828)
         );
  OAI211_X1 U8695 ( .C1(n8000), .C2(n8044), .A(n6829), .B(n6828), .ZN(P2_U3172) );
  INV_X1 U8696 ( .A(n8424), .ZN(n8438) );
  INV_X1 U8697 ( .A(n6062), .ZN(n6831) );
  OAI222_X1 U8698 ( .A1(P2_U3151), .A2(n8438), .B1(n7670), .B2(n6831), .C1(
        n6830), .C2(n8816), .ZN(P2_U3279) );
  INV_X1 U8699 ( .A(n10037), .ZN(n9574) );
  OAI222_X1 U8700 ( .A1(n9995), .A2(n6832), .B1(n9993), .B2(n6831), .C1(n9574), 
        .C2(n10066), .ZN(P1_U3339) );
  INV_X1 U8701 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6838) );
  NOR2_X1 U8702 ( .A1(n10153), .A2(n8640), .ZN(n6833) );
  OR2_X1 U8703 ( .A1(n8044), .A2(n6833), .ZN(n6836) );
  OR2_X1 U8704 ( .A1(n6928), .A2(n8658), .ZN(n6839) );
  OAI21_X1 U8705 ( .B1(n6844), .B2(n10150), .A(n6839), .ZN(n6834) );
  INV_X1 U8706 ( .A(n6834), .ZN(n6835) );
  NAND2_X1 U8707 ( .A1(n6836), .A2(n6835), .ZN(n8741) );
  NAND2_X1 U8708 ( .A1(n10155), .A2(n8741), .ZN(n6837) );
  OAI21_X1 U8709 ( .B1(n10155), .B2(n6838), .A(n6837), .ZN(P2_U3390) );
  NAND2_X1 U8710 ( .A1(n10150), .A2(n6856), .ZN(n6840) );
  OAI21_X1 U8711 ( .B1(n8044), .B2(n6840), .A(n6839), .ZN(n6841) );
  MUX2_X1 U8712 ( .A(P2_REG2_REG_0__SCAN_IN), .B(n6841), .S(n8663), .Z(n6846)
         );
  NOR2_X2 U8713 ( .A1(n6842), .A2(n8671), .ZN(n8666) );
  OAI22_X1 U8714 ( .A1(n8630), .A2(n6844), .B1(n6843), .B2(n8643), .ZN(n6845)
         );
  OR2_X1 U8715 ( .A1(n6846), .A2(n6845), .ZN(P2_U3233) );
  NAND2_X1 U8716 ( .A1(n6847), .A2(n8245), .ZN(n6849) );
  INV_X2 U8717 ( .A(n6854), .ZN(n6893) );
  OAI21_X1 U8718 ( .B1(n6893), .B2(n6850), .A(n8087), .ZN(n6863) );
  XNOR2_X1 U8719 ( .A(n6895), .B(n5880), .ZN(n6897) );
  XOR2_X1 U8720 ( .A(n6898), .B(n6897), .Z(n6862) );
  NOR2_X1 U8721 ( .A1(n6856), .A2(n6855), .ZN(n6857) );
  AND2_X2 U8722 ( .A1(n6858), .A2(n6857), .ZN(n8007) );
  AOI22_X1 U8723 ( .A1(n7984), .A2(n6271), .B1(n8007), .B2(n8277), .ZN(n6859)
         );
  OAI21_X1 U8724 ( .B1(n10126), .B2(n8015), .A(n6859), .ZN(n6860) );
  AOI21_X1 U8725 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6867), .A(n6860), .ZN(
        n6861) );
  OAI21_X1 U8726 ( .B1(n6862), .B2(n8000), .A(n6861), .ZN(P2_U3177) );
  XOR2_X1 U8727 ( .A(n6864), .B(n6863), .Z(n6869) );
  AOI22_X1 U8728 ( .A1(n7984), .A2(n6476), .B1(n8007), .B2(n8278), .ZN(n6865)
         );
  OAI21_X1 U8729 ( .B1(n10122), .B2(n8015), .A(n6865), .ZN(n6866) );
  AOI21_X1 U8730 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6867), .A(n6866), .ZN(
        n6868) );
  OAI21_X1 U8731 ( .B1(n8000), .B2(n6869), .A(n6868), .ZN(P2_U3162) );
  INV_X1 U8732 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6879) );
  INV_X1 U8733 ( .A(n6979), .ZN(n6872) );
  OAI21_X1 U8734 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n4415), .A(n6872), .ZN(
        n6877) );
  NAND2_X1 U8735 ( .A1(n6881), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U8736 ( .A1(n6874), .A2(n6873), .ZN(n6875) );
  NAND2_X1 U8737 ( .A1(n6875), .A2(n6966), .ZN(n6971) );
  OAI21_X1 U8738 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n4416), .A(n6972), .ZN(
        n6876) );
  AOI22_X1 U8739 ( .A1(n6877), .A2(n8345), .B1(n8492), .B2(n6876), .ZN(n6878)
         );
  NAND2_X1 U8740 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7027) );
  OAI211_X1 U8741 ( .C1(n8371), .C2(n6879), .A(n6878), .B(n7027), .ZN(n6886)
         );
  MUX2_X1 U8742 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8405), .Z(n6967) );
  XOR2_X1 U8743 ( .A(n6887), .B(n6967), .Z(n6883) );
  AOI211_X1 U8744 ( .C1(n6884), .C2(n6883), .A(n8482), .B(n6965), .ZN(n6885)
         );
  AOI211_X1 U8745 ( .C1(n8373), .C2(n6887), .A(n6886), .B(n6885), .ZN(n6888)
         );
  INV_X1 U8746 ( .A(n6888), .ZN(P2_U3187) );
  INV_X1 U8747 ( .A(n6889), .ZN(n6890) );
  AOI21_X1 U8748 ( .B1(n8007), .B2(n6476), .A(n6890), .ZN(n6892) );
  OAI211_X1 U8749 ( .C1(n7009), .C2(n8009), .A(n6892), .B(n6891), .ZN(n6902)
         );
  INV_X4 U8750 ( .A(n6893), .ZN(n7813) );
  XNOR2_X1 U8751 ( .A(n7813), .B(n10132), .ZN(n6937) );
  XNOR2_X1 U8752 ( .A(n6937), .B(n6894), .ZN(n6900) );
  INV_X1 U8753 ( .A(n6895), .ZN(n6896) );
  AOI211_X1 U8754 ( .C1(n6900), .C2(n6899), .A(n8000), .B(n6938), .ZN(n6901)
         );
  AOI211_X1 U8755 ( .C1(n7130), .C2(n8011), .A(n6902), .B(n6901), .ZN(n6903)
         );
  INV_X1 U8756 ( .A(n6903), .ZN(P2_U3158) );
  OAI21_X1 U8757 ( .B1(n6904), .B2(n9243), .A(n6905), .ZN(n7544) );
  INV_X1 U8758 ( .A(n6953), .ZN(n6906) );
  AOI211_X1 U8759 ( .C1(n7054), .C2(n6906), .A(n9832), .B(n5133), .ZN(n7538)
         );
  NAND2_X1 U8760 ( .A1(n6907), .A2(n9846), .ZN(n6914) );
  INV_X1 U8761 ( .A(n9243), .ZN(n6909) );
  AOI21_X1 U8762 ( .B1(n6908), .B2(n9280), .A(n6909), .ZN(n6913) );
  NAND2_X1 U8763 ( .A1(n9468), .A2(n9843), .ZN(n6911) );
  NAND2_X1 U8764 ( .A1(n9470), .A2(n9841), .ZN(n6910) );
  NAND2_X1 U8765 ( .A1(n6911), .A2(n6910), .ZN(n7053) );
  INV_X1 U8766 ( .A(n7053), .ZN(n6912) );
  OAI21_X1 U8767 ( .B1(n6914), .B2(n6913), .A(n6912), .ZN(n7537) );
  AOI211_X1 U8768 ( .C1(n10113), .C2(n7544), .A(n7538), .B(n7537), .ZN(n6919)
         );
  AOI22_X1 U8769 ( .A1(n9899), .A2(n7054), .B1(n10118), .B2(
        P1_REG1_REG_5__SCAN_IN), .ZN(n6915) );
  OAI21_X1 U8770 ( .B1(n6919), .B2(n10118), .A(n6915), .ZN(P1_U3527) );
  INV_X1 U8771 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n6916) );
  OAI22_X1 U8772 ( .A1(n9981), .A2(n7542), .B1(n10348), .B2(n6916), .ZN(n6917)
         );
  INV_X1 U8773 ( .A(n6917), .ZN(n6918) );
  OAI21_X1 U8774 ( .B1(n6919), .B2(n10346), .A(n6918), .ZN(P1_U3468) );
  INV_X1 U8775 ( .A(n6920), .ZN(n6923) );
  INV_X1 U8776 ( .A(n6921), .ZN(n6922) );
  AOI21_X1 U8777 ( .B1(n6923), .B2(n6272), .A(n6922), .ZN(n10128) );
  INV_X1 U8778 ( .A(n6924), .ZN(n6925) );
  AND2_X1 U8779 ( .A1(n8663), .A2(n6925), .ZN(n7757) );
  INV_X1 U8780 ( .A(n7757), .ZN(n7019) );
  INV_X1 U8781 ( .A(n7135), .ZN(n8050) );
  INV_X1 U8782 ( .A(n6926), .ZN(n6927) );
  NOR2_X1 U8783 ( .A1(n8050), .A2(n6927), .ZN(n7133) );
  AOI211_X1 U8784 ( .C1(n6928), .C2(n10122), .A(n6272), .B(n7133), .ZN(n6931)
         );
  INV_X1 U8785 ( .A(n6929), .ZN(n6930) );
  OAI21_X1 U8786 ( .B1(n6931), .B2(n6930), .A(n8640), .ZN(n6933) );
  AOI22_X1 U8787 ( .A1(n8277), .A2(n8573), .B1(n8571), .B2(n6271), .ZN(n6932)
         );
  OAI211_X1 U8788 ( .C1(n10128), .C2(n7648), .A(n6933), .B(n6932), .ZN(n10130)
         );
  OAI22_X1 U8789 ( .A1(n8643), .A2(n5850), .B1(n10126), .B2(n8671), .ZN(n6934)
         );
  NOR2_X1 U8790 ( .A1(n10130), .A2(n6934), .ZN(n6935) );
  MUX2_X1 U8791 ( .A(n5847), .B(n6935), .S(n8663), .Z(n6936) );
  OAI21_X1 U8792 ( .B1(n10128), .B2(n7019), .A(n6936), .ZN(P2_U3231) );
  INV_X1 U8793 ( .A(n7119), .ZN(n10139) );
  XNOR2_X1 U8794 ( .A(n7813), .B(n10139), .ZN(n7023) );
  XNOR2_X1 U8795 ( .A(n7023), .B(n8276), .ZN(n6941) );
  INV_X1 U8796 ( .A(n6937), .ZN(n6939) );
  AOI21_X1 U8797 ( .B1(n6271), .B2(n6939), .A(n6938), .ZN(n6940) );
  OAI21_X1 U8798 ( .B1(n6941), .B2(n6940), .A(n7024), .ZN(n6942) );
  NAND2_X1 U8799 ( .A1(n6942), .A2(n8003), .ZN(n6948) );
  INV_X1 U8800 ( .A(n6943), .ZN(n6944) );
  AOI21_X1 U8801 ( .B1(n8007), .B2(n6271), .A(n6944), .ZN(n6945) );
  OAI21_X1 U8802 ( .B1(n7075), .B2(n8009), .A(n6945), .ZN(n6946) );
  AOI21_X1 U8803 ( .B1(n7119), .B2(n7998), .A(n6946), .ZN(n6947) );
  OAI211_X1 U8804 ( .C1(n7117), .C2(n7953), .A(n6948), .B(n6947), .ZN(P2_U3170) );
  AND2_X1 U8805 ( .A1(n6949), .A2(n6950), .ZN(n7182) );
  NOR2_X1 U8806 ( .A1(n7182), .A2(n6951), .ZN(n6952) );
  INV_X1 U8807 ( .A(n5763), .ZN(n9246) );
  XNOR2_X1 U8808 ( .A(n6952), .B(n9246), .ZN(n7327) );
  AOI211_X1 U8809 ( .C1(n9123), .C2(n7176), .A(n9832), .B(n6953), .ZN(n7333)
         );
  INV_X1 U8810 ( .A(n9275), .ZN(n6954) );
  OAI21_X1 U8811 ( .B1(n6954), .B2(n9281), .A(n5763), .ZN(n6955) );
  AOI21_X1 U8812 ( .B1(n6955), .B2(n6908), .A(n9761), .ZN(n6959) );
  OR2_X1 U8813 ( .A1(n6956), .A2(n9808), .ZN(n6958) );
  NAND2_X1 U8814 ( .A1(n9469), .A2(n9843), .ZN(n6957) );
  NAND2_X1 U8815 ( .A1(n6958), .A2(n6957), .ZN(n9121) );
  OR2_X1 U8816 ( .A1(n6959), .A2(n9121), .ZN(n7328) );
  AOI211_X1 U8817 ( .C1(n10113), .C2(n7327), .A(n7333), .B(n7328), .ZN(n6964)
         );
  INV_X1 U8818 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6960) );
  OAI22_X1 U8819 ( .A1(n9981), .A2(n7330), .B1(n10348), .B2(n6960), .ZN(n6961)
         );
  INV_X1 U8820 ( .A(n6961), .ZN(n6962) );
  OAI21_X1 U8821 ( .B1(n6964), .B2(n10346), .A(n6962), .ZN(P1_U3465) );
  AOI22_X1 U8822 ( .A1(n9899), .A2(n9123), .B1(n10118), .B2(
        P1_REG1_REG_4__SCAN_IN), .ZN(n6963) );
  OAI21_X1 U8823 ( .B1(n6964), .B2(n10118), .A(n6963), .ZN(P1_U3526) );
  MUX2_X1 U8824 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8405), .Z(n7089) );
  XNOR2_X1 U8825 ( .A(n7089), .B(n7095), .ZN(n6968) );
  OAI21_X1 U8826 ( .B1(n6969), .B2(n6968), .A(n7087), .ZN(n6970) );
  NAND2_X1 U8827 ( .A1(n6970), .A2(n8436), .ZN(n6984) );
  INV_X1 U8828 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6976) );
  NAND3_X1 U8829 ( .A1(n6972), .A2(n4417), .A3(n6971), .ZN(n6973) );
  NAND2_X1 U8830 ( .A1(n7091), .A2(n6973), .ZN(n6974) );
  NAND2_X1 U8831 ( .A1(n8492), .A2(n6974), .ZN(n6975) );
  NAND2_X1 U8832 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7080) );
  OAI211_X1 U8833 ( .C1(n8371), .C2(n6976), .A(n6975), .B(n7080), .ZN(n6982)
         );
  XNOR2_X1 U8834 ( .A(n7095), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n6977) );
  OR3_X1 U8835 ( .A1(n6979), .A2(n6978), .A3(n6977), .ZN(n6980) );
  AOI21_X1 U8836 ( .B1(n7097), .B2(n6980), .A(n8495), .ZN(n6981) );
  AOI211_X1 U8837 ( .C1(n8373), .C2(n7095), .A(n6982), .B(n6981), .ZN(n6983)
         );
  NAND2_X1 U8838 ( .A1(n6984), .A2(n6983), .ZN(P2_U3188) );
  XNOR2_X1 U8839 ( .A(n9576), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n6989) );
  INV_X1 U8840 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U8841 ( .A1(n6991), .A2(n10248), .ZN(n6985) );
  NAND2_X1 U8842 ( .A1(n6986), .A2(n6985), .ZN(n6988) );
  INV_X1 U8843 ( .A(n9578), .ZN(n6987) );
  AOI211_X1 U8844 ( .C1(n6989), .C2(n6988), .A(n10055), .B(n6987), .ZN(n7002)
         );
  XNOR2_X1 U8845 ( .A(n9576), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n6996) );
  INV_X1 U8846 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8847 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  NAND2_X1 U8848 ( .A1(n6993), .A2(n6992), .ZN(n6995) );
  INV_X1 U8849 ( .A(n9564), .ZN(n6994) );
  AOI211_X1 U8850 ( .C1(n6996), .C2(n6995), .A(n10060), .B(n6994), .ZN(n7001)
         );
  INV_X1 U8851 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n6999) );
  NAND2_X1 U8852 ( .A1(n4409), .A2(n9576), .ZN(n6998) );
  AND2_X1 U8853 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9159) );
  INV_X1 U8854 ( .A(n9159), .ZN(n6997) );
  OAI211_X1 U8855 ( .C1(n6999), .C2(n10070), .A(n6998), .B(n6997), .ZN(n7000)
         );
  OR3_X1 U8856 ( .A1(n7002), .A2(n7001), .A3(n7000), .ZN(P1_U3256) );
  INV_X1 U8857 ( .A(n7003), .ZN(n7005) );
  OAI222_X1 U8858 ( .A1(n9995), .A2(n7004), .B1(n9993), .B2(n7005), .C1(n10066), .C2(n9765), .ZN(P1_U3336) );
  OAI222_X1 U8859 ( .A1(n8816), .A2(n7006), .B1(n7670), .B2(n7005), .C1(n8487), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  XNOR2_X1 U8860 ( .A(n7007), .B(n8049), .ZN(n10146) );
  INV_X1 U8861 ( .A(n10146), .ZN(n7020) );
  INV_X1 U8862 ( .A(n7648), .ZN(n7015) );
  OAI22_X1 U8863 ( .A1(n7009), .A2(n8656), .B1(n8123), .B2(n8658), .ZN(n7014)
         );
  NAND2_X1 U8864 ( .A1(n7011), .A2(n8049), .ZN(n7012) );
  AOI21_X1 U8865 ( .B1(n7010), .B2(n7012), .A(n8653), .ZN(n7013) );
  AOI211_X1 U8866 ( .C1(n10146), .C2(n7015), .A(n7014), .B(n7013), .ZN(n10148)
         );
  MUX2_X1 U8867 ( .A(n4754), .B(n10148), .S(n6405), .Z(n7018) );
  INV_X1 U8868 ( .A(n7034), .ZN(n7016) );
  AOI22_X1 U8869 ( .A1(n8666), .A2(n10143), .B1(n8677), .B2(n7016), .ZN(n7017)
         );
  OAI211_X1 U8870 ( .C1(n7020), .C2(n7019), .A(n7018), .B(n7017), .ZN(P2_U3228) );
  NAND2_X1 U8871 ( .A1(n9473), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7021) );
  OAI21_X1 U8872 ( .B1(n7022), .B2(n9473), .A(n7021), .ZN(P1_U3583) );
  XNOR2_X1 U8873 ( .A(n7813), .B(n7025), .ZN(n7074) );
  XNOR2_X1 U8874 ( .A(n7074), .B(n8275), .ZN(n7076) );
  XNOR2_X1 U8875 ( .A(n7077), .B(n7076), .ZN(n7026) );
  NAND2_X1 U8876 ( .A1(n7026), .A2(n8003), .ZN(n7033) );
  INV_X1 U8877 ( .A(n7027), .ZN(n7028) );
  AOI21_X1 U8878 ( .B1(n8007), .B2(n8276), .A(n7028), .ZN(n7030) );
  NAND2_X1 U8879 ( .A1(n7998), .A2(n10143), .ZN(n7029) );
  OAI211_X1 U8880 ( .C1(n8123), .C2(n8009), .A(n7030), .B(n7029), .ZN(n7031)
         );
  INV_X1 U8881 ( .A(n7031), .ZN(n7032) );
  OAI211_X1 U8882 ( .C1(n7034), .C2(n7953), .A(n7033), .B(n7032), .ZN(P2_U3167) );
  INV_X1 U8883 ( .A(n7035), .ZN(n7036) );
  AND2_X1 U8884 ( .A1(n9470), .A2(n8952), .ZN(n7041) );
  AOI21_X1 U8885 ( .B1(n9123), .B2(n7040), .A(n7041), .ZN(n7045) );
  NAND2_X1 U8886 ( .A1(n9470), .A2(n7040), .ZN(n7042) );
  OAI21_X1 U8887 ( .B1(n7330), .B2(n8922), .A(n7042), .ZN(n7043) );
  XNOR2_X1 U8888 ( .A(n7043), .B(n8964), .ZN(n7044) );
  NOR2_X1 U8889 ( .A1(n7044), .A2(n7045), .ZN(n7046) );
  AOI21_X1 U8890 ( .B1(n7045), .B2(n7044), .A(n7046), .ZN(n9118) );
  INV_X1 U8891 ( .A(n7046), .ZN(n7047) );
  OAI22_X1 U8892 ( .A1(n7542), .A2(n8922), .B1(n7051), .B2(n4293), .ZN(n7048)
         );
  XNOR2_X1 U8893 ( .A(n7048), .B(n9034), .ZN(n7049) );
  NAND2_X1 U8894 ( .A1(n5009), .A2(n7210), .ZN(n7052) );
  OAI22_X1 U8895 ( .A1(n7542), .A2(n4293), .B1(n7051), .B2(n8947), .ZN(n7208)
         );
  XNOR2_X1 U8896 ( .A(n7052), .B(n7208), .ZN(n7059) );
  INV_X1 U8897 ( .A(n7539), .ZN(n7057) );
  AOI22_X1 U8898 ( .A1(n9202), .A2(n7053), .B1(P1_REG3_REG_5__SCAN_IN), .B2(
        n10066), .ZN(n7056) );
  NAND2_X1 U8899 ( .A1(n9215), .A2(n7054), .ZN(n7055) );
  OAI211_X1 U8900 ( .C1(n9210), .C2(n7057), .A(n7056), .B(n7055), .ZN(n7058)
         );
  AOI21_X1 U8901 ( .B1(n7059), .B2(n9196), .A(n7058), .ZN(n7060) );
  INV_X1 U8902 ( .A(n7060), .ZN(P1_U3227) );
  OAI21_X1 U8903 ( .B1(n7061), .B2(n7199), .A(n7062), .ZN(n7337) );
  INV_X1 U8904 ( .A(n7198), .ZN(n7063) );
  AOI211_X1 U8905 ( .C1(n7317), .C2(n7064), .A(n9832), .B(n7063), .ZN(n7345)
         );
  XOR2_X1 U8906 ( .A(n7065), .B(n7199), .Z(n7068) );
  NAND2_X1 U8907 ( .A1(n9469), .A2(n9841), .ZN(n7067) );
  NAND2_X1 U8908 ( .A1(n9467), .A2(n9843), .ZN(n7066) );
  AND2_X1 U8909 ( .A1(n7067), .A2(n7066), .ZN(n7319) );
  OAI21_X1 U8910 ( .B1(n7068), .B2(n9761), .A(n7319), .ZN(n7338) );
  AOI211_X1 U8911 ( .C1(n10113), .C2(n7337), .A(n7345), .B(n7338), .ZN(n7073)
         );
  AOI22_X1 U8912 ( .A1(n9899), .A2(n7317), .B1(n10118), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n7069) );
  OAI21_X1 U8913 ( .B1(n7073), .B2(n10118), .A(n7069), .ZN(P1_U3528) );
  INV_X1 U8914 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7070) );
  OAI22_X1 U8915 ( .A1(n9981), .A2(n7339), .B1(n10348), .B2(n7070), .ZN(n7071)
         );
  INV_X1 U8916 ( .A(n7071), .ZN(n7072) );
  OAI21_X1 U8917 ( .B1(n7073), .B2(n10346), .A(n7072), .ZN(P1_U3471) );
  XNOR2_X1 U8918 ( .A(n7809), .B(n10151), .ZN(n7419) );
  XNOR2_X1 U8919 ( .A(n7419), .B(n8274), .ZN(n7078) );
  OAI211_X1 U8920 ( .C1(n7079), .C2(n7078), .A(n7421), .B(n8003), .ZN(n7086)
         );
  INV_X1 U8921 ( .A(n7080), .ZN(n7081) );
  AOI21_X1 U8922 ( .B1(n8007), .B2(n8275), .A(n7081), .ZN(n7083) );
  NAND2_X1 U8923 ( .A1(n7998), .A2(n8122), .ZN(n7082) );
  OAI211_X1 U8924 ( .C1(n7423), .C2(n8009), .A(n7083), .B(n7082), .ZN(n7084)
         );
  INV_X1 U8925 ( .A(n7084), .ZN(n7085) );
  OAI211_X1 U8926 ( .C1(n7170), .C2(n7953), .A(n7086), .B(n7085), .ZN(P2_U3179) );
  MUX2_X1 U8927 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8405), .Z(n7141) );
  XNOR2_X1 U8928 ( .A(n7141), .B(n7143), .ZN(n7144) );
  XOR2_X1 U8929 ( .A(n7144), .B(n7145), .Z(n7106) );
  OR2_X1 U8930 ( .A1(n7095), .A2(n10166), .ZN(n7090) );
  NAND2_X1 U8931 ( .A1(n7091), .A2(n7090), .ZN(n7092) );
  NAND2_X1 U8932 ( .A1(n7092), .A2(n7098), .ZN(n7150) );
  OAI21_X1 U8933 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n7093), .A(n7147), .ZN(
        n7104) );
  NAND2_X1 U8934 ( .A1(n8484), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7094) );
  NAND2_X1 U8935 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7450) );
  OAI211_X1 U8936 ( .C1(n8488), .C2(n7098), .A(n7094), .B(n7450), .ZN(n7103)
         );
  INV_X1 U8937 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7169) );
  NAND2_X1 U8938 ( .A1(n7088), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7096) );
  NAND2_X1 U8939 ( .A1(n7097), .A2(n7096), .ZN(n7099) );
  AOI21_X1 U8940 ( .B1(n10245), .B2(n7100), .A(n7158), .ZN(n7101) );
  NOR2_X1 U8941 ( .A1(n7101), .A2(n8495), .ZN(n7102) );
  AOI211_X1 U8942 ( .C1(n8492), .C2(n7104), .A(n7103), .B(n7102), .ZN(n7105)
         );
  OAI21_X1 U8943 ( .B1(n7106), .B2(n8482), .A(n7105), .ZN(P2_U3189) );
  INV_X1 U8944 ( .A(n7107), .ZN(n7109) );
  OAI222_X1 U8945 ( .A1(n9995), .A2(n7108), .B1(n9993), .B2(n7109), .C1(n9267), 
        .C2(P1_U3086), .ZN(P1_U3335) );
  OAI222_X1 U8946 ( .A1(n8816), .A2(n7110), .B1(P2_U3151), .B2(n8242), .C1(
        n8822), .C2(n7109), .ZN(P2_U3275) );
  AND2_X1 U8947 ( .A1(n7112), .A2(n7111), .ZN(n7113) );
  XNOR2_X1 U8948 ( .A(n7113), .B(n8100), .ZN(n10141) );
  INV_X1 U8949 ( .A(n10141), .ZN(n7122) );
  INV_X1 U8950 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7116) );
  XOR2_X1 U8951 ( .A(n7114), .B(n8100), .Z(n7115) );
  AOI222_X1 U8952 ( .A1(n6271), .A2(n8573), .B1(n8640), .B2(n7115), .C1(n8275), 
        .C2(n8571), .ZN(n10138) );
  MUX2_X1 U8953 ( .A(n7116), .B(n10138), .S(n6405), .Z(n7121) );
  INV_X1 U8954 ( .A(n7117), .ZN(n7118) );
  AOI22_X1 U8955 ( .A1(n8666), .A2(n7119), .B1(n8677), .B2(n7118), .ZN(n7120)
         );
  OAI211_X1 U8956 ( .C1(n7122), .C2(n8669), .A(n7121), .B(n7120), .ZN(P2_U3229) );
  NAND2_X1 U8957 ( .A1(n6921), .A2(n8094), .ZN(n7124) );
  NAND2_X1 U8958 ( .A1(n7124), .A2(n8048), .ZN(n7126) );
  NAND3_X1 U8959 ( .A1(n6921), .A2(n8094), .A3(n7123), .ZN(n7125) );
  AND2_X1 U8960 ( .A1(n7126), .A2(n7125), .ZN(n10134) );
  INV_X1 U8961 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7129) );
  XOR2_X1 U8962 ( .A(n7127), .B(n8048), .Z(n7128) );
  AOI222_X1 U8963 ( .A1(n7128), .A2(n8640), .B1(n8276), .B2(n8571), .C1(n6476), 
        .C2(n8573), .ZN(n10131) );
  MUX2_X1 U8964 ( .A(n7129), .B(n10131), .S(n6405), .Z(n7132) );
  OAI211_X1 U8965 ( .C1(n10134), .C2(n8669), .A(n7132), .B(n7131), .ZN(
        P2_U3230) );
  XNOR2_X1 U8966 ( .A(n8050), .B(n8087), .ZN(n10120) );
  INV_X1 U8967 ( .A(n7133), .ZN(n7134) );
  OAI21_X1 U8968 ( .B1(n7135), .B2(n6926), .A(n7134), .ZN(n7136) );
  AOI222_X1 U8969 ( .A1(n7136), .A2(n8640), .B1(n6476), .B2(n8571), .C1(n8278), 
        .C2(n8573), .ZN(n10121) );
  MUX2_X1 U8970 ( .A(n7137), .B(n10121), .S(n8663), .Z(n7140) );
  AOI22_X1 U8971 ( .A1(n8666), .A2(n7138), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8677), .ZN(n7139) );
  OAI211_X1 U8972 ( .C1(n10120), .C2(n8669), .A(n7140), .B(n7139), .ZN(
        P2_U3232) );
  MUX2_X1 U8973 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8405), .Z(n7307) );
  XOR2_X1 U8974 ( .A(n7297), .B(n7307), .Z(n7308) );
  INV_X1 U8975 ( .A(n7141), .ZN(n7142) );
  XOR2_X1 U8976 ( .A(n7308), .B(n7309), .Z(n7162) );
  INV_X1 U8977 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7146) );
  NAND2_X1 U8978 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7427) );
  OAI21_X1 U8979 ( .B1(n8371), .B2(n7146), .A(n7427), .ZN(n7154) );
  NAND2_X1 U8980 ( .A1(n7147), .A2(n7150), .ZN(n7148) );
  XNOR2_X1 U8981 ( .A(n7297), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7149) );
  NAND2_X1 U8982 ( .A1(n7148), .A2(n7149), .ZN(n7299) );
  INV_X1 U8983 ( .A(n7149), .ZN(n7151) );
  NAND3_X1 U8984 ( .A1(n7147), .A2(n7151), .A3(n7150), .ZN(n7152) );
  AOI21_X1 U8985 ( .B1(n7299), .B2(n7152), .A(n7302), .ZN(n7153) );
  AOI211_X1 U8986 ( .C1(n8373), .C2(n7297), .A(n7154), .B(n7153), .ZN(n7161)
         );
  XNOR2_X1 U8987 ( .A(n7297), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7156) );
  NOR3_X1 U8988 ( .A1(n7158), .A2(n7157), .A3(n7156), .ZN(n7159) );
  OAI21_X1 U8989 ( .B1(n4412), .B2(n7159), .A(n8345), .ZN(n7160) );
  OAI211_X1 U8990 ( .C1(n7162), .C2(n8482), .A(n7161), .B(n7160), .ZN(P2_U3190) );
  NAND2_X1 U8991 ( .A1(n7007), .A2(n8110), .ZN(n7402) );
  NAND2_X1 U8992 ( .A1(n7402), .A2(n8104), .ZN(n7164) );
  INV_X1 U8993 ( .A(n7163), .ZN(n8045) );
  XNOR2_X1 U8994 ( .A(n7164), .B(n8045), .ZN(n10154) );
  INV_X1 U8995 ( .A(n10154), .ZN(n7174) );
  NAND3_X1 U8996 ( .A1(n7010), .A2(n8045), .A3(n7166), .ZN(n7167) );
  NAND2_X1 U8997 ( .A1(n7165), .A2(n7167), .ZN(n7168) );
  AOI222_X1 U8998 ( .A1(n7168), .A2(n8640), .B1(n8275), .B2(n8573), .C1(n8273), 
        .C2(n8571), .ZN(n10149) );
  MUX2_X1 U8999 ( .A(n7169), .B(n10149), .S(n8663), .Z(n7173) );
  INV_X1 U9000 ( .A(n7170), .ZN(n7171) );
  AOI22_X1 U9001 ( .A1(n8666), .A2(n8122), .B1(n8677), .B2(n7171), .ZN(n7172)
         );
  OAI211_X1 U9002 ( .C1(n8669), .C2(n7174), .A(n7173), .B(n7172), .ZN(P2_U3227) );
  XNOR2_X1 U9003 ( .A(n9282), .B(n6950), .ZN(n7175) );
  AOI222_X1 U9004 ( .A1(n9846), .A2(n7175), .B1(n9472), .B2(n9841), .C1(n9470), 
        .C2(n9843), .ZN(n10116) );
  OAI211_X1 U9005 ( .C1(n7177), .C2(n10111), .A(n9782), .B(n7176), .ZN(n10109)
         );
  NOR2_X1 U9006 ( .A1(n9783), .A2(n10109), .ZN(n7180) );
  OAI22_X1 U9007 ( .A1(n9855), .A2(n7178), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9852), .ZN(n7179) );
  AOI211_X1 U9008 ( .C1(n10074), .C2(n7181), .A(n7180), .B(n7179), .ZN(n7185)
         );
  INV_X1 U9009 ( .A(n7182), .ZN(n7183) );
  OAI21_X1 U9010 ( .B1(n6950), .B2(n6949), .A(n7183), .ZN(n10114) );
  NAND2_X1 U9011 ( .A1(n10114), .A2(n10071), .ZN(n7184) );
  OAI211_X1 U9012 ( .C1(n10116), .C2(n10084), .A(n7185), .B(n7184), .ZN(
        P1_U3290) );
  INV_X1 U9013 ( .A(n10127), .ZN(n10145) );
  NAND2_X1 U9014 ( .A1(n7402), .A2(n8114), .ZN(n7187) );
  INV_X1 U9015 ( .A(n8125), .ZN(n8046) );
  AOI21_X1 U9016 ( .B1(n7187), .B2(n8106), .A(n8046), .ZN(n7271) );
  INV_X1 U9017 ( .A(n8106), .ZN(n8115) );
  NOR2_X1 U9018 ( .A1(n8125), .A2(n8115), .ZN(n7186) );
  AND2_X1 U9019 ( .A1(n7187), .A2(n7186), .ZN(n7188) );
  OR2_X1 U9020 ( .A1(n7271), .A2(n7188), .ZN(n7190) );
  INV_X1 U9021 ( .A(n7190), .ZN(n7353) );
  XNOR2_X1 U9022 ( .A(n7189), .B(n8125), .ZN(n7193) );
  OR2_X1 U9023 ( .A1(n7190), .A2(n7648), .ZN(n7192) );
  AOI22_X1 U9024 ( .A1(n8274), .A2(n8573), .B1(n8571), .B2(n8272), .ZN(n7191)
         );
  OAI211_X1 U9025 ( .C1(n8653), .C2(n7193), .A(n7192), .B(n7191), .ZN(n7350)
         );
  AOI21_X1 U9026 ( .B1(n10145), .B2(n7353), .A(n7350), .ZN(n7314) );
  INV_X1 U9027 ( .A(n8801), .ZN(n8747) );
  OAI22_X1 U9028 ( .A1(n8747), .A2(n7349), .B1(n5944), .B2(n10155), .ZN(n7194)
         );
  INV_X1 U9029 ( .A(n7194), .ZN(n7195) );
  OAI21_X1 U9030 ( .B1(n7314), .B2(n10156), .A(n7195), .ZN(P2_U3411) );
  OAI21_X1 U9031 ( .B1(n7196), .B2(n7232), .A(n7197), .ZN(n7534) );
  AOI211_X1 U9032 ( .C1(n7221), .C2(n7198), .A(n9832), .B(n7230), .ZN(n7528)
         );
  OAI21_X1 U9033 ( .B1(n7065), .B2(n7199), .A(n9284), .ZN(n7235) );
  XNOR2_X1 U9034 ( .A(n7235), .B(n7232), .ZN(n7202) );
  NAND2_X1 U9035 ( .A1(n9468), .A2(n9841), .ZN(n7200) );
  OAI21_X1 U9036 ( .B1(n9137), .B2(n9810), .A(n7200), .ZN(n7220) );
  INV_X1 U9037 ( .A(n7220), .ZN(n7201) );
  OAI21_X1 U9038 ( .B1(n7202), .B2(n9761), .A(n7201), .ZN(n7527) );
  AOI211_X1 U9039 ( .C1(n10113), .C2(n7534), .A(n7528), .B(n7527), .ZN(n7207)
         );
  AOI22_X1 U9040 ( .A1(n9899), .A2(n7221), .B1(n10118), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n7203) );
  OAI21_X1 U9041 ( .B1(n7207), .B2(n10118), .A(n7203), .ZN(P1_U3529) );
  INV_X1 U9042 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7204) );
  OAI22_X1 U9043 ( .A1(n9981), .A2(n7532), .B1(n10348), .B2(n7204), .ZN(n7205)
         );
  INV_X1 U9044 ( .A(n7205), .ZN(n7206) );
  OAI21_X1 U9045 ( .B1(n7207), .B2(n10346), .A(n7206), .ZN(P1_U3474) );
  INV_X1 U9046 ( .A(n7208), .ZN(n7209) );
  NAND2_X1 U9047 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  AND2_X2 U9048 ( .A1(n5009), .A2(n7211), .ZN(n7320) );
  OAI22_X1 U9049 ( .A1(n7339), .A2(n8922), .B1(n7212), .B2(n4294), .ZN(n7213)
         );
  XNOR2_X1 U9050 ( .A(n7213), .B(n9034), .ZN(n7216) );
  NAND2_X1 U9051 ( .A1(n9468), .A2(n8952), .ZN(n7214) );
  OAI21_X1 U9052 ( .B1(n7339), .B2(n4294), .A(n7214), .ZN(n7215) );
  XNOR2_X1 U9053 ( .A(n7216), .B(n7215), .ZN(n7321) );
  OAI22_X1 U9054 ( .A1(n7532), .A2(n8922), .B1(n7218), .B2(n4293), .ZN(n7217)
         );
  XNOR2_X1 U9055 ( .A(n7217), .B(n9034), .ZN(n7578) );
  OAI22_X1 U9056 ( .A1(n7532), .A2(n4294), .B1(n7218), .B2(n8947), .ZN(n7577)
         );
  INV_X1 U9057 ( .A(n7577), .ZN(n7580) );
  XNOR2_X1 U9058 ( .A(n7578), .B(n7580), .ZN(n7219) );
  XNOR2_X1 U9059 ( .A(n7581), .B(n7219), .ZN(n7226) );
  INV_X1 U9060 ( .A(n7529), .ZN(n7224) );
  AOI22_X1 U9061 ( .A1(n9202), .A2(n7220), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7223) );
  NAND2_X1 U9062 ( .A1(n9215), .A2(n7221), .ZN(n7222) );
  OAI211_X1 U9063 ( .C1(n9210), .C2(n7224), .A(n7223), .B(n7222), .ZN(n7225)
         );
  AOI21_X1 U9064 ( .B1(n7226), .B2(n9196), .A(n7225), .ZN(n7227) );
  INV_X1 U9065 ( .A(n7227), .ZN(P1_U3213) );
  OAI21_X1 U9066 ( .B1(n7228), .B2(n7236), .A(n7229), .ZN(n9858) );
  OAI21_X1 U9067 ( .B1(n7230), .B2(n7244), .A(n9782), .ZN(n7231) );
  NOR2_X1 U9068 ( .A1(n7231), .A2(n7379), .ZN(n9859) );
  INV_X1 U9069 ( .A(n7232), .ZN(n9288) );
  INV_X1 U9070 ( .A(n7233), .ZN(n7234) );
  AOI21_X1 U9071 ( .B1(n7235), .B2(n9288), .A(n7234), .ZN(n7238) );
  INV_X1 U9072 ( .A(n7236), .ZN(n7237) );
  NAND2_X1 U9073 ( .A1(n7238), .A2(n7237), .ZN(n7382) );
  OAI211_X1 U9074 ( .C1(n7238), .C2(n7237), .A(n7382), .B(n9846), .ZN(n7241)
         );
  NAND2_X1 U9075 ( .A1(n9467), .A2(n9841), .ZN(n7239) );
  OAI21_X1 U9076 ( .B1(n8828), .B2(n9810), .A(n7239), .ZN(n7589) );
  INV_X1 U9077 ( .A(n7589), .ZN(n7240) );
  NAND2_X1 U9078 ( .A1(n7241), .A2(n7240), .ZN(n9851) );
  AOI211_X1 U9079 ( .C1(n10113), .C2(n9858), .A(n9859), .B(n9851), .ZN(n7247)
         );
  AOI22_X1 U9080 ( .A1(n9899), .A2(n9857), .B1(n10118), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7242) );
  OAI21_X1 U9081 ( .B1(n7247), .B2(n10118), .A(n7242), .ZN(P1_U3530) );
  INV_X1 U9082 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7243) );
  OAI22_X1 U9083 ( .A1(n9981), .A2(n7244), .B1(n10348), .B2(n7243), .ZN(n7245)
         );
  INV_X1 U9084 ( .A(n7245), .ZN(n7246) );
  OAI21_X1 U9085 ( .B1(n7247), .B2(n10346), .A(n7246), .ZN(P1_U3477) );
  INV_X1 U9086 ( .A(n6125), .ZN(n7249) );
  OAI222_X1 U9087 ( .A1(n9995), .A2(n7248), .B1(n9993), .B2(n7249), .C1(n6686), 
        .C2(n10066), .ZN(P1_U3334) );
  OAI222_X1 U9088 ( .A1(n8816), .A2(n7250), .B1(P2_U3151), .B2(n6847), .C1(
        n8822), .C2(n7249), .ZN(P2_U3274) );
  INV_X1 U9089 ( .A(n7252), .ZN(n7253) );
  AOI21_X1 U9090 ( .B1(n7251), .B2(n7254), .A(n7253), .ZN(n7259) );
  AOI22_X1 U9091 ( .A1(n9472), .A2(n9843), .B1(n9841), .B2(n9474), .ZN(n7258)
         );
  OAI21_X1 U9092 ( .B1(n7251), .B2(n7256), .A(n7255), .ZN(n10104) );
  INV_X1 U9093 ( .A(n9815), .ZN(n7438) );
  NAND2_X1 U9094 ( .A1(n10104), .A2(n7438), .ZN(n7257) );
  OAI211_X1 U9095 ( .C1(n7259), .C2(n9761), .A(n7258), .B(n7257), .ZN(n10102)
         );
  INV_X1 U9096 ( .A(n7260), .ZN(n7261) );
  NAND2_X1 U9097 ( .A1(n9855), .A2(n7261), .ZN(n9824) );
  INV_X1 U9098 ( .A(n9824), .ZN(n7262) );
  AOI22_X1 U9099 ( .A1(n10102), .A2(n9855), .B1(n7262), .B2(n10104), .ZN(n7269) );
  INV_X1 U9100 ( .A(n7263), .ZN(n7264) );
  OAI211_X1 U9101 ( .C1(n10101), .C2(n7265), .A(n7264), .B(n9782), .ZN(n10100)
         );
  OAI22_X1 U9102 ( .A1(n9783), .A2(n10100), .B1(n7266), .B2(n9852), .ZN(n7267)
         );
  AOI21_X1 U9103 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n10084), .A(n7267), .ZN(
        n7268) );
  OAI211_X1 U9104 ( .C1(n10101), .C2(n9836), .A(n7269), .B(n7268), .ZN(
        P1_U3292) );
  INV_X1 U9105 ( .A(n8134), .ZN(n7270) );
  NOR2_X1 U9106 ( .A1(n7271), .A2(n7270), .ZN(n7272) );
  AND2_X1 U9107 ( .A1(n8135), .A2(n8128), .ZN(n8053) );
  XNOR2_X1 U9108 ( .A(n7272), .B(n8053), .ZN(n7525) );
  XNOR2_X1 U9109 ( .A(n7273), .B(n8053), .ZN(n7274) );
  OAI222_X1 U9110 ( .A1(n8658), .A2(n7560), .B1(n8656), .B2(n7423), .C1(n7274), 
        .C2(n8653), .ZN(n7522) );
  AOI21_X1 U9111 ( .B1(n10153), .B2(n7525), .A(n7522), .ZN(n7398) );
  AOI22_X1 U9112 ( .A1(n8801), .A2(n7429), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10156), .ZN(n7275) );
  OAI21_X1 U9113 ( .B1(n7398), .B2(n10156), .A(n7275), .ZN(P2_U3414) );
  OAI21_X1 U9114 ( .B1(n7276), .B2(n9250), .A(n7277), .ZN(n7505) );
  AOI211_X1 U9115 ( .C1(n9019), .C2(n7378), .A(n9832), .B(n4398), .ZN(n7506)
         );
  INV_X1 U9116 ( .A(n7278), .ZN(n7279) );
  AOI21_X1 U9117 ( .B1(n9250), .B2(n7280), .A(n7279), .ZN(n7281) );
  OAI222_X1 U9118 ( .A1(n9810), .A2(n9072), .B1(n9808), .B2(n8828), .C1(n9761), 
        .C2(n7281), .ZN(n7511) );
  AOI211_X1 U9119 ( .C1(n10113), .C2(n7505), .A(n7506), .B(n7511), .ZN(n7284)
         );
  AOI22_X1 U9120 ( .A1(n9899), .A2(n9019), .B1(n10118), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7282) );
  OAI21_X1 U9121 ( .B1(n7284), .B2(n10118), .A(n7282), .ZN(P1_U3532) );
  AOI22_X1 U9122 ( .A1(n6326), .A2(n9019), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n10346), .ZN(n7283) );
  OAI21_X1 U9123 ( .B1(n7284), .B2(n10346), .A(n7283), .ZN(P1_U3483) );
  INV_X1 U9124 ( .A(n7285), .ZN(n7289) );
  OAI222_X1 U9125 ( .A1(n9995), .A2(n7287), .B1(n9993), .B2(n7289), .C1(
        P1_U3086), .C2(n7286), .ZN(P1_U3333) );
  OAI222_X1 U9126 ( .A1(n8816), .A2(n7290), .B1(n7670), .B2(n7289), .C1(n7288), 
        .C2(P2_U3151), .ZN(P2_U3273) );
  INV_X1 U9127 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7295) );
  INV_X1 U9128 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7291) );
  NAND2_X1 U9129 ( .A1(n7292), .A2(n7300), .ZN(n7361) );
  AOI21_X1 U9130 ( .B1(n7295), .B2(n7294), .A(n7364), .ZN(n7313) );
  INV_X1 U9131 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7296) );
  NAND2_X1 U9132 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7561) );
  OAI21_X1 U9133 ( .B1(n8371), .B2(n7296), .A(n7561), .ZN(n7305) );
  OR2_X1 U9134 ( .A1(n7297), .A2(n7399), .ZN(n7298) );
  AOI21_X1 U9135 ( .B1(n7569), .B2(n7301), .A(n4396), .ZN(n7303) );
  NOR2_X1 U9136 ( .A1(n7303), .A2(n7302), .ZN(n7304) );
  AOI211_X1 U9137 ( .C1(n8373), .C2(n7357), .A(n7305), .B(n7304), .ZN(n7312)
         );
  MUX2_X1 U9138 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8405), .Z(n7355) );
  XNOR2_X1 U9139 ( .A(n7355), .B(n7357), .ZN(n7358) );
  XNOR2_X1 U9140 ( .A(n7359), .B(n7358), .ZN(n7310) );
  NAND2_X1 U9141 ( .A1(n7310), .A2(n8436), .ZN(n7311) );
  OAI211_X1 U9142 ( .C1(n7313), .C2(n8495), .A(n7312), .B(n7311), .ZN(P2_U3191) );
  INV_X1 U9143 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7315) );
  MUX2_X1 U9144 ( .A(n7315), .B(n7314), .S(n10168), .Z(n7316) );
  OAI21_X1 U9145 ( .B1(n7349), .B2(n8696), .A(n7316), .ZN(P2_U3466) );
  NAND2_X1 U9146 ( .A1(n9215), .A2(n7317), .ZN(n7318) );
  NAND2_X1 U9147 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9511) );
  OAI211_X1 U9148 ( .C1(n7319), .C2(n9167), .A(n7318), .B(n9511), .ZN(n7325)
         );
  XOR2_X1 U9149 ( .A(n7322), .B(n7321), .Z(n7323) );
  NOR2_X1 U9150 ( .A1(n7323), .A2(n9217), .ZN(n7324) );
  AOI211_X1 U9151 ( .C1(n7340), .C2(n9165), .A(n7325), .B(n7324), .ZN(n7326)
         );
  INV_X1 U9152 ( .A(n7326), .ZN(P1_U3239) );
  INV_X1 U9153 ( .A(n7327), .ZN(n7336) );
  NAND2_X1 U9154 ( .A1(n7328), .A2(n9855), .ZN(n7335) );
  INV_X1 U9155 ( .A(n9122), .ZN(n7329) );
  OAI22_X1 U9156 ( .A1(n9855), .A2(n5524), .B1(n7329), .B2(n9852), .ZN(n7332)
         );
  NOR2_X1 U9157 ( .A1(n9836), .A2(n7330), .ZN(n7331) );
  AOI211_X1 U9158 ( .C1(n7333), .C2(n10076), .A(n7332), .B(n7331), .ZN(n7334)
         );
  OAI211_X1 U9159 ( .C1(n7336), .C2(n9850), .A(n7335), .B(n7334), .ZN(P1_U3289) );
  INV_X1 U9160 ( .A(n7337), .ZN(n7348) );
  NAND2_X1 U9161 ( .A1(n7338), .A2(n9855), .ZN(n7347) );
  NOR2_X1 U9162 ( .A1(n9836), .A2(n7339), .ZN(n7344) );
  INV_X1 U9163 ( .A(n7340), .ZN(n7341) );
  OAI22_X1 U9164 ( .A1(n9855), .A2(n7342), .B1(n7341), .B2(n9852), .ZN(n7343)
         );
  AOI211_X1 U9165 ( .C1(n7345), .C2(n10076), .A(n7344), .B(n7343), .ZN(n7346)
         );
  OAI211_X1 U9166 ( .C1(n7348), .C2(n9850), .A(n7347), .B(n7346), .ZN(P1_U3287) );
  OAI22_X1 U9167 ( .A1(n8630), .A2(n7349), .B1(n7449), .B2(n8643), .ZN(n7352)
         );
  MUX2_X1 U9168 ( .A(n7350), .B(P2_REG2_REG_7__SCAN_IN), .S(n8681), .Z(n7351)
         );
  AOI211_X1 U9169 ( .C1(n7353), .C2(n7757), .A(n7352), .B(n7351), .ZN(n7354)
         );
  INV_X1 U9170 ( .A(n7354), .ZN(P2_U3226) );
  MUX2_X1 U9171 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8405), .Z(n8280) );
  XOR2_X1 U9172 ( .A(n8295), .B(n8280), .Z(n8281) );
  INV_X1 U9173 ( .A(n7355), .ZN(n7356) );
  XOR2_X1 U9174 ( .A(n8282), .B(n8281), .Z(n7375) );
  INV_X1 U9175 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7360) );
  NAND2_X1 U9176 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n7689) );
  OAI21_X1 U9177 ( .B1(n8371), .B2(n7360), .A(n7689), .ZN(n7367) );
  INV_X1 U9178 ( .A(n7361), .ZN(n7363) );
  XNOR2_X1 U9179 ( .A(n8295), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n7362) );
  OR3_X1 U9180 ( .A1(n7364), .A2(n7363), .A3(n7362), .ZN(n7365) );
  AOI21_X1 U9181 ( .B1(n8285), .B2(n7365), .A(n8495), .ZN(n7366) );
  AOI211_X1 U9182 ( .C1(n8373), .C2(n8295), .A(n7367), .B(n7366), .ZN(n7374)
         );
  XNOR2_X1 U9183 ( .A(n8295), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n7369) );
  NOR3_X1 U9184 ( .A1(n4396), .A2(n4783), .A3(n7369), .ZN(n7372) );
  NAND2_X1 U9185 ( .A1(n7370), .A2(n7369), .ZN(n8297) );
  INV_X1 U9186 ( .A(n8297), .ZN(n7371) );
  OAI21_X1 U9187 ( .B1(n7372), .B2(n7371), .A(n8492), .ZN(n7373) );
  OAI211_X1 U9188 ( .C1(n7375), .C2(n8482), .A(n7374), .B(n7373), .ZN(P2_U3192) );
  OAI21_X1 U9189 ( .B1(n7376), .B2(n7384), .A(n7377), .ZN(n7490) );
  OAI211_X1 U9190 ( .C1(n9142), .C2(n7379), .A(n7378), .B(n9782), .ZN(n7380)
         );
  OAI21_X1 U9191 ( .B1(n9178), .B2(n9810), .A(n7380), .ZN(n7486) );
  NAND2_X1 U9192 ( .A1(n7382), .A2(n7381), .ZN(n7383) );
  XOR2_X1 U9193 ( .A(n7384), .B(n7383), .Z(n7385) );
  OAI22_X1 U9194 ( .A1(n7385), .A2(n9761), .B1(n9137), .B2(n9808), .ZN(n7485)
         );
  AOI211_X1 U9195 ( .C1(n10113), .C2(n7490), .A(n7486), .B(n7485), .ZN(n7390)
         );
  INV_X1 U9196 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7386) );
  OAI22_X1 U9197 ( .A1(n9981), .A2(n9142), .B1(n10348), .B2(n7386), .ZN(n7387)
         );
  INV_X1 U9198 ( .A(n7387), .ZN(n7388) );
  OAI21_X1 U9199 ( .B1(n7390), .B2(n10346), .A(n7388), .ZN(P1_U3480) );
  AOI22_X1 U9200 ( .A1(n9899), .A2(n8830), .B1(n10118), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7389) );
  OAI21_X1 U9201 ( .B1(n7390), .B2(n10118), .A(n7389), .ZN(P1_U3531) );
  NAND2_X1 U9202 ( .A1(n7396), .A2(n7391), .ZN(n7393) );
  OR2_X1 U9203 ( .A1(n7392), .A2(P2_U3151), .ZN(n8254) );
  OAI211_X1 U9204 ( .C1(n7394), .C2(n8816), .A(n7393), .B(n8254), .ZN(P2_U3272) );
  NAND2_X1 U9205 ( .A1(n7396), .A2(n7395), .ZN(n7397) );
  OAI211_X1 U9206 ( .C1(n10231), .C2(n9995), .A(n7397), .B(n9452), .ZN(
        P1_U3332) );
  INV_X1 U9207 ( .A(n7429), .ZN(n7521) );
  MUX2_X1 U9208 ( .A(n7399), .B(n7398), .S(n10168), .Z(n7400) );
  OAI21_X1 U9209 ( .B1(n7521), .B2(n8696), .A(n7400), .ZN(P2_U3467) );
  NAND2_X1 U9210 ( .A1(n7402), .A2(n7401), .ZN(n7404) );
  NAND2_X1 U9211 ( .A1(n7404), .A2(n7403), .ZN(n7405) );
  NAND2_X1 U9212 ( .A1(n7405), .A2(n8128), .ZN(n7406) );
  NAND2_X1 U9213 ( .A1(n7406), .A2(n8043), .ZN(n7409) );
  CLKBUF_X1 U9214 ( .A(n7407), .Z(n7408) );
  NAND2_X1 U9215 ( .A1(n7409), .A2(n7408), .ZN(n7417) );
  INV_X1 U9216 ( .A(n7417), .ZN(n7620) );
  AND2_X1 U9217 ( .A1(n7411), .A2(n7410), .ZN(n7413) );
  OAI21_X1 U9218 ( .B1(n7413), .B2(n8043), .A(n7412), .ZN(n7414) );
  NAND2_X1 U9219 ( .A1(n7414), .A2(n8640), .ZN(n7416) );
  AOI22_X1 U9220 ( .A1(n8571), .A2(n8270), .B1(n8573), .B2(n7557), .ZN(n7415)
         );
  OAI211_X1 U9221 ( .C1(n7417), .C2(n7648), .A(n7416), .B(n7415), .ZN(n7617)
         );
  AOI21_X1 U9222 ( .B1(n10145), .B2(n7620), .A(n7617), .ZN(n7568) );
  AOI22_X1 U9223 ( .A1(n8801), .A2(n7567), .B1(n10156), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n7418) );
  OAI21_X1 U9224 ( .B1(n7568), .B2(n10156), .A(n7418), .ZN(P2_U3417) );
  XNOR2_X1 U9225 ( .A(n7809), .B(n7452), .ZN(n7422) );
  INV_X1 U9226 ( .A(n7422), .ZN(n7424) );
  XNOR2_X1 U9227 ( .A(n7422), .B(n8273), .ZN(n7458) );
  XNOR2_X1 U9228 ( .A(n7429), .B(n7813), .ZN(n7556) );
  XNOR2_X1 U9229 ( .A(n7556), .B(n7557), .ZN(n7425) );
  XNOR2_X1 U9230 ( .A(n7555), .B(n7425), .ZN(n7426) );
  NAND2_X1 U9231 ( .A1(n7426), .A2(n8003), .ZN(n7434) );
  INV_X1 U9232 ( .A(n7427), .ZN(n7428) );
  AOI21_X1 U9233 ( .B1(n8007), .B2(n8273), .A(n7428), .ZN(n7431) );
  NAND2_X1 U9234 ( .A1(n7998), .A2(n7429), .ZN(n7430) );
  OAI211_X1 U9235 ( .C1(n7560), .C2(n8009), .A(n7431), .B(n7430), .ZN(n7432)
         );
  INV_X1 U9236 ( .A(n7432), .ZN(n7433) );
  OAI211_X1 U9237 ( .C1(n7520), .C2(n7953), .A(n7434), .B(n7433), .ZN(P2_U3161) );
  OAI21_X1 U9238 ( .B1(n7436), .B2(n9241), .A(n7435), .ZN(n7551) );
  INV_X1 U9239 ( .A(n7551), .ZN(n7448) );
  NAND2_X1 U9240 ( .A1(n7278), .A2(n9303), .ZN(n7437) );
  XNOR2_X1 U9241 ( .A(n7437), .B(n9241), .ZN(n7441) );
  NAND2_X1 U9242 ( .A1(n7551), .A2(n7438), .ZN(n7440) );
  AOI22_X1 U9243 ( .A1(n9841), .A2(n9464), .B1(n9842), .B2(n9843), .ZN(n7439)
         );
  OAI211_X1 U9244 ( .C1(n9761), .C2(n7441), .A(n7440), .B(n7439), .ZN(n7549)
         );
  NAND2_X1 U9245 ( .A1(n7549), .A2(n9855), .ZN(n7447) );
  INV_X1 U9246 ( .A(n7442), .ZN(n9177) );
  OAI22_X1 U9247 ( .A1(n9855), .A2(n7443), .B1(n9177), .B2(n9852), .ZN(n7445)
         );
  OAI211_X1 U9248 ( .C1(n5201), .C2(n4398), .A(n7499), .B(n9782), .ZN(n7548)
         );
  NOR2_X1 U9249 ( .A1(n7548), .A2(n9783), .ZN(n7444) );
  AOI211_X1 U9250 ( .C1(n10074), .C2(n8845), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OAI211_X1 U9251 ( .C1(n7448), .C2(n9824), .A(n7447), .B(n7446), .ZN(P1_U3282) );
  INV_X1 U9252 ( .A(n7449), .ZN(n7462) );
  INV_X1 U9253 ( .A(n7450), .ZN(n7451) );
  AOI21_X1 U9254 ( .B1(n8007), .B2(n8274), .A(n7451), .ZN(n7454) );
  NAND2_X1 U9255 ( .A1(n7998), .A2(n7452), .ZN(n7453) );
  OAI211_X1 U9256 ( .C1(n7455), .C2(n8009), .A(n7454), .B(n7453), .ZN(n7461)
         );
  AOI21_X1 U9257 ( .B1(n7458), .B2(n7457), .A(n7456), .ZN(n7459) );
  NOR2_X1 U9258 ( .A1(n7459), .A2(n8000), .ZN(n7460) );
  AOI211_X1 U9259 ( .C1(n7462), .C2(n8011), .A(n7461), .B(n7460), .ZN(n7463)
         );
  INV_X1 U9260 ( .A(n7463), .ZN(P2_U3153) );
  INV_X1 U9261 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10178) );
  INV_X1 U9262 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10069) );
  INV_X1 U9263 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10052) );
  INV_X1 U9264 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n7464) );
  AOI22_X1 U9265 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10052), .B2(n7464), .ZN(n10181) );
  INV_X1 U9266 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10257) );
  INV_X1 U9267 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7465) );
  AOI22_X1 U9268 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10257), .B2(n7465), .ZN(n10184) );
  NOR2_X1 U9269 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7466) );
  AOI21_X1 U9270 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7466), .ZN(n10187) );
  NOR2_X1 U9271 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7467) );
  AOI21_X1 U9272 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7467), .ZN(n10190) );
  NOR2_X1 U9273 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7468) );
  AOI21_X1 U9274 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7468), .ZN(n10193) );
  NOR2_X1 U9275 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7469) );
  AOI21_X1 U9276 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7469), .ZN(n10196) );
  NOR2_X1 U9277 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7470) );
  AOI21_X1 U9278 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7470), .ZN(n10199) );
  NOR2_X1 U9279 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n7471) );
  AOI21_X1 U9280 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7471), .ZN(n10202) );
  NOR2_X1 U9281 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7472) );
  AOI21_X1 U9282 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7472), .ZN(n10359) );
  NOR2_X1 U9283 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7473) );
  AOI21_X1 U9284 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7473), .ZN(n10365) );
  NOR2_X1 U9285 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7474) );
  AOI21_X1 U9286 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7474), .ZN(n10362) );
  NOR2_X1 U9287 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7475) );
  AOI21_X1 U9288 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7475), .ZN(n10353) );
  NOR2_X1 U9289 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7476) );
  AOI21_X1 U9290 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7476), .ZN(n10356) );
  AND2_X1 U9291 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7477) );
  NOR2_X1 U9292 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7477), .ZN(n10170) );
  INV_X1 U9293 ( .A(n10170), .ZN(n10171) );
  INV_X1 U9294 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10173) );
  NAND3_X1 U9295 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U9296 ( .A1(n10173), .A2(n10172), .ZN(n10169) );
  NAND2_X1 U9297 ( .A1(n10171), .A2(n10169), .ZN(n10368) );
  NAND2_X1 U9298 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7478) );
  OAI21_X1 U9299 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7478), .ZN(n10367) );
  NOR2_X1 U9300 ( .A1(n10368), .A2(n10367), .ZN(n10366) );
  AOI21_X1 U9301 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10366), .ZN(n10371) );
  NAND2_X1 U9302 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7479) );
  OAI21_X1 U9303 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n7479), .ZN(n10370) );
  NOR2_X1 U9304 ( .A1(n10371), .A2(n10370), .ZN(n10369) );
  AOI21_X1 U9305 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10369), .ZN(n10374) );
  NOR2_X1 U9306 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7480) );
  AOI21_X1 U9307 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7480), .ZN(n10373) );
  NAND2_X1 U9308 ( .A1(n10374), .A2(n10373), .ZN(n10372) );
  OAI21_X1 U9309 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10372), .ZN(n10355) );
  NAND2_X1 U9310 ( .A1(n10356), .A2(n10355), .ZN(n10354) );
  OAI21_X1 U9311 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10354), .ZN(n10352) );
  NAND2_X1 U9312 ( .A1(n10353), .A2(n10352), .ZN(n10351) );
  OAI21_X1 U9313 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10351), .ZN(n10361) );
  NAND2_X1 U9314 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  OAI21_X1 U9315 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10360), .ZN(n10364) );
  NAND2_X1 U9316 ( .A1(n10365), .A2(n10364), .ZN(n10363) );
  OAI21_X1 U9317 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10363), .ZN(n10358) );
  NAND2_X1 U9318 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  OAI21_X1 U9319 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10357), .ZN(n10201) );
  NAND2_X1 U9320 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  OAI21_X1 U9321 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10200), .ZN(n10198) );
  NAND2_X1 U9322 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  OAI21_X1 U9323 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10197), .ZN(n10195) );
  NAND2_X1 U9324 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  OAI21_X1 U9325 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10194), .ZN(n10192) );
  NAND2_X1 U9326 ( .A1(n10193), .A2(n10192), .ZN(n10191) );
  OAI21_X1 U9327 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10191), .ZN(n10189) );
  NAND2_X1 U9328 ( .A1(n10190), .A2(n10189), .ZN(n10188) );
  OAI21_X1 U9329 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10188), .ZN(n10186) );
  NAND2_X1 U9330 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  OAI21_X1 U9331 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10185), .ZN(n10183) );
  NAND2_X1 U9332 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  OAI21_X1 U9333 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10182), .ZN(n10180) );
  NAND2_X1 U9334 ( .A1(n10181), .A2(n10180), .ZN(n10179) );
  OAI21_X1 U9335 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10179), .ZN(n7481) );
  OR2_X1 U9336 ( .A1(n10069), .A2(n7481), .ZN(n10177) );
  NAND2_X1 U9337 ( .A1(n10178), .A2(n10177), .ZN(n10174) );
  NAND2_X1 U9338 ( .A1(n10069), .A2(n7481), .ZN(n10176) );
  NAND2_X1 U9339 ( .A1(n10174), .A2(n10176), .ZN(n7484) );
  XNOR2_X1 U9340 ( .A(n7482), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7483) );
  XNOR2_X1 U9341 ( .A(n7484), .B(n7483), .ZN(ADD_1068_U4) );
  INV_X1 U9342 ( .A(n7485), .ZN(n7492) );
  NAND2_X1 U9343 ( .A1(n7486), .A2(n10076), .ZN(n7488) );
  AOI22_X1 U9344 ( .A1(n10084), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9135), .B2(
        n10094), .ZN(n7487) );
  OAI211_X1 U9345 ( .C1(n9142), .C2(n9836), .A(n7488), .B(n7487), .ZN(n7489)
         );
  AOI21_X1 U9346 ( .B1(n7490), .B2(n10071), .A(n7489), .ZN(n7491) );
  OAI21_X1 U9347 ( .B1(n7492), .B2(n10084), .A(n7491), .ZN(P1_U3284) );
  OAI21_X1 U9348 ( .B1(n7493), .B2(n9240), .A(n7494), .ZN(n7516) );
  INV_X1 U9349 ( .A(n7516), .ZN(n7504) );
  INV_X1 U9350 ( .A(n7495), .ZN(n7496) );
  AOI21_X1 U9351 ( .B1(n9240), .B2(n7497), .A(n7496), .ZN(n7498) );
  OAI222_X1 U9352 ( .A1(n9810), .A2(n9809), .B1(n9808), .B2(n9072), .C1(n9761), 
        .C2(n7498), .ZN(n7514) );
  AOI211_X1 U9353 ( .C1(n8856), .C2(n7499), .A(n9832), .B(n9830), .ZN(n7515)
         );
  NAND2_X1 U9354 ( .A1(n7515), .A2(n10076), .ZN(n7501) );
  AOI22_X1 U9355 ( .A1(n10084), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n9070), .B2(
        n10094), .ZN(n7500) );
  OAI211_X1 U9356 ( .C1(n4793), .C2(n9836), .A(n7501), .B(n7500), .ZN(n7502)
         );
  AOI21_X1 U9357 ( .B1(n7514), .B2(n9855), .A(n7502), .ZN(n7503) );
  OAI21_X1 U9358 ( .B1(n7504), .B2(n9850), .A(n7503), .ZN(P1_U3281) );
  INV_X1 U9359 ( .A(n7505), .ZN(n7513) );
  INV_X1 U9360 ( .A(n9019), .ZN(n7509) );
  NAND2_X1 U9361 ( .A1(n7506), .A2(n10076), .ZN(n7508) );
  AOI22_X1 U9362 ( .A1(n10084), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n9014), .B2(
        n10094), .ZN(n7507) );
  OAI211_X1 U9363 ( .C1(n7509), .C2(n9836), .A(n7508), .B(n7507), .ZN(n7510)
         );
  AOI21_X1 U9364 ( .B1(n7511), .B2(n9855), .A(n7510), .ZN(n7512) );
  OAI21_X1 U9365 ( .B1(n7513), .B2(n9850), .A(n7512), .ZN(P1_U3283) );
  AOI211_X1 U9366 ( .C1(n10113), .C2(n7516), .A(n7515), .B(n7514), .ZN(n7519)
         );
  AOI22_X1 U9367 ( .A1(n8856), .A2(n9899), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n10118), .ZN(n7517) );
  OAI21_X1 U9368 ( .B1(n7519), .B2(n10118), .A(n7517), .ZN(P1_U3534) );
  AOI22_X1 U9369 ( .A1(n8856), .A2(n6326), .B1(P1_REG0_REG_12__SCAN_IN), .B2(
        n10346), .ZN(n7518) );
  OAI21_X1 U9370 ( .B1(n7519), .B2(n10346), .A(n7518), .ZN(P1_U3489) );
  OAI22_X1 U9371 ( .A1(n8630), .A2(n7521), .B1(n7520), .B2(n8643), .ZN(n7524)
         );
  MUX2_X1 U9372 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7522), .S(n8663), .Z(n7523)
         );
  AOI211_X1 U9373 ( .C1(n8678), .C2(n7525), .A(n7524), .B(n7523), .ZN(n7526)
         );
  INV_X1 U9374 ( .A(n7526), .ZN(P2_U3225) );
  INV_X1 U9375 ( .A(n7527), .ZN(n7536) );
  NAND2_X1 U9376 ( .A1(n7528), .A2(n10076), .ZN(n7531) );
  AOI22_X1 U9377 ( .A1(n10084), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7529), .B2(
        n10094), .ZN(n7530) );
  OAI211_X1 U9378 ( .C1(n7532), .C2(n9836), .A(n7531), .B(n7530), .ZN(n7533)
         );
  AOI21_X1 U9379 ( .B1(n7534), .B2(n10071), .A(n7533), .ZN(n7535) );
  OAI21_X1 U9380 ( .B1(n7536), .B2(n10084), .A(n7535), .ZN(P1_U3286) );
  INV_X1 U9381 ( .A(n7537), .ZN(n7546) );
  NAND2_X1 U9382 ( .A1(n7538), .A2(n10076), .ZN(n7541) );
  AOI22_X1 U9383 ( .A1(n10084), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7539), .B2(
        n10094), .ZN(n7540) );
  OAI211_X1 U9384 ( .C1(n7542), .C2(n9836), .A(n7541), .B(n7540), .ZN(n7543)
         );
  AOI21_X1 U9385 ( .B1(n10071), .B2(n7544), .A(n7543), .ZN(n7545) );
  OAI21_X1 U9386 ( .B1(n10084), .B2(n7546), .A(n7545), .ZN(P1_U3288) );
  INV_X1 U9387 ( .A(n7547), .ZN(n10105) );
  OAI21_X1 U9388 ( .B1(n5201), .B2(n10110), .A(n7548), .ZN(n7550) );
  AOI211_X1 U9389 ( .C1(n10105), .C2(n7551), .A(n7550), .B(n7549), .ZN(n7554)
         );
  NAND2_X1 U9390 ( .A1(n10118), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7552) );
  OAI21_X1 U9391 ( .B1(n7554), .B2(n10118), .A(n7552), .ZN(P1_U3533) );
  NAND2_X1 U9392 ( .A1(n10346), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7553) );
  OAI21_X1 U9393 ( .B1(n7554), .B2(n10346), .A(n7553), .ZN(P1_U3486) );
  NAND2_X1 U9394 ( .A1(n7556), .A2(n7557), .ZN(n7558) );
  XNOR2_X1 U9395 ( .A(n7567), .B(n7813), .ZN(n7685) );
  XNOR2_X1 U9396 ( .A(n7685), .B(n7560), .ZN(n7686) );
  XNOR2_X1 U9397 ( .A(n7687), .B(n7686), .ZN(n7566) );
  NAND2_X1 U9398 ( .A1(n8007), .A2(n8272), .ZN(n7562) );
  OAI211_X1 U9399 ( .C1(n7882), .C2(n8009), .A(n7562), .B(n7561), .ZN(n7564)
         );
  NOR2_X1 U9400 ( .A1(n7953), .A2(n7615), .ZN(n7563) );
  AOI211_X1 U9401 ( .C1(n7567), .C2(n7998), .A(n7564), .B(n7563), .ZN(n7565)
         );
  OAI21_X1 U9402 ( .B1(n7566), .B2(n8000), .A(n7565), .ZN(P2_U3171) );
  INV_X1 U9403 ( .A(n7567), .ZN(n7616) );
  MUX2_X1 U9404 ( .A(n7569), .B(n7568), .S(n10168), .Z(n7570) );
  OAI21_X1 U9405 ( .B1(n7616), .B2(n8696), .A(n7570), .ZN(P2_U3468) );
  INV_X1 U9406 ( .A(n7571), .ZN(n7655) );
  OAI222_X1 U9407 ( .A1(n9995), .A2(n7573), .B1(n10066), .B2(n7572), .C1(n7655), .C2(n9993), .ZN(P1_U3331) );
  NAND2_X1 U9408 ( .A1(n8457), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7574) );
  OAI21_X1 U9409 ( .B1(n7818), .B2(n8457), .A(n7574), .ZN(P2_U3520) );
  NAND2_X1 U9410 ( .A1(n9857), .A2(n7040), .ZN(n7576) );
  NAND2_X1 U9411 ( .A1(n9466), .A2(n8952), .ZN(n7575) );
  NAND2_X1 U9412 ( .A1(n7576), .A2(n7575), .ZN(n8839) );
  INV_X1 U9413 ( .A(n7578), .ZN(n7579) );
  INV_X1 U9414 ( .A(n8844), .ZN(n7585) );
  NAND2_X1 U9415 ( .A1(n9857), .A2(n4290), .ZN(n7583) );
  NAND2_X1 U9416 ( .A1(n9466), .A2(n7040), .ZN(n7582) );
  NAND2_X1 U9417 ( .A1(n7583), .A2(n7582), .ZN(n7584) );
  XNOR2_X1 U9418 ( .A(n7584), .B(n9034), .ZN(n8831) );
  INV_X1 U9419 ( .A(n8831), .ZN(n8841) );
  NAND2_X1 U9420 ( .A1(n7585), .A2(n8841), .ZN(n9128) );
  OAI21_X1 U9421 ( .B1(n7585), .B2(n8841), .A(n9128), .ZN(n7586) );
  NOR2_X1 U9422 ( .A1(n7586), .A2(n8839), .ZN(n9131) );
  AOI21_X1 U9423 ( .B1(n8839), .B2(n7586), .A(n9131), .ZN(n7594) );
  INV_X1 U9424 ( .A(n7587), .ZN(n9853) );
  NAND2_X1 U9425 ( .A1(n10066), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9537) );
  INV_X1 U9426 ( .A(n9537), .ZN(n7588) );
  AOI21_X1 U9427 ( .B1(n9202), .B2(n7589), .A(n7588), .ZN(n7591) );
  NAND2_X1 U9428 ( .A1(n9215), .A2(n9857), .ZN(n7590) );
  OAI211_X1 U9429 ( .C1(n9210), .C2(n9853), .A(n7591), .B(n7590), .ZN(n7592)
         );
  INV_X1 U9430 ( .A(n7592), .ZN(n7593) );
  OAI21_X1 U9431 ( .B1(n7594), .B2(n9217), .A(n7593), .ZN(P1_U3221) );
  NAND2_X1 U9432 ( .A1(n7597), .A2(n7596), .ZN(n7598) );
  NAND2_X1 U9433 ( .A1(n7598), .A2(n8058), .ZN(n7599) );
  NAND3_X1 U9434 ( .A1(n7595), .A2(n8640), .A3(n7599), .ZN(n7601) );
  AOI22_X1 U9435 ( .A1(n8571), .A2(n8268), .B1(n8573), .B2(n8270), .ZN(n7600)
         );
  MUX2_X1 U9436 ( .A(n7610), .B(n7602), .S(n10165), .Z(n7605) );
  XNOR2_X1 U9437 ( .A(n7603), .B(n8058), .ZN(n7609) );
  AOI22_X1 U9438 ( .A1(n7609), .A2(n8734), .B1(n8733), .B2(n7971), .ZN(n7604)
         );
  NAND2_X1 U9439 ( .A1(n7605), .A2(n7604), .ZN(P2_U3470) );
  MUX2_X1 U9440 ( .A(n7610), .B(n7606), .S(n10156), .Z(n7608) );
  AOI22_X1 U9441 ( .A1(n7609), .A2(n8802), .B1(n8801), .B2(n7971), .ZN(n7607)
         );
  NAND2_X1 U9442 ( .A1(n7608), .A2(n7607), .ZN(P2_U3423) );
  INV_X1 U9443 ( .A(n7609), .ZN(n7614) );
  INV_X1 U9444 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8290) );
  MUX2_X1 U9445 ( .A(n7610), .B(n8290), .S(n8681), .Z(n7613) );
  INV_X1 U9446 ( .A(n7611), .ZN(n7975) );
  AOI22_X1 U9447 ( .A1(n8666), .A2(n7971), .B1(n8677), .B2(n7975), .ZN(n7612)
         );
  OAI211_X1 U9448 ( .C1(n7614), .C2(n8669), .A(n7613), .B(n7612), .ZN(P2_U3222) );
  OAI22_X1 U9449 ( .A1(n8630), .A2(n7616), .B1(n7615), .B2(n8643), .ZN(n7619)
         );
  MUX2_X1 U9450 ( .A(n7617), .B(P2_REG2_REG_9__SCAN_IN), .S(n8681), .Z(n7618)
         );
  AOI211_X1 U9451 ( .C1(n7620), .C2(n7757), .A(n7619), .B(n7618), .ZN(n7621)
         );
  INV_X1 U9452 ( .A(n7621), .ZN(P2_U3224) );
  NAND2_X1 U9453 ( .A1(n7595), .A2(n7622), .ZN(n7624) );
  AND2_X1 U9454 ( .A1(n7624), .A2(n7623), .ZN(n7625) );
  NAND2_X1 U9455 ( .A1(n7625), .A2(n8059), .ZN(n7626) );
  NAND2_X1 U9456 ( .A1(n7627), .A2(n7626), .ZN(n7628) );
  NAND2_X1 U9457 ( .A1(n7628), .A2(n8640), .ZN(n7630) );
  AOI22_X1 U9458 ( .A1(n8571), .A2(n8266), .B1(n8573), .B2(n8268), .ZN(n7629)
         );
  NAND2_X1 U9459 ( .A1(n7630), .A2(n7629), .ZN(n7675) );
  INV_X1 U9460 ( .A(n8157), .ZN(n7631) );
  OAI22_X1 U9461 ( .A1(n7631), .A2(n8671), .B1(n7954), .B2(n8643), .ZN(n7632)
         );
  OAI21_X1 U9462 ( .B1(n7675), .B2(n7632), .A(n8663), .ZN(n7636) );
  CLKBUF_X1 U9463 ( .A(n7633), .Z(n7634) );
  XNOR2_X1 U9464 ( .A(n7634), .B(n6032), .ZN(n7677) );
  AOI22_X1 U9465 ( .A1(n7677), .A2(n8678), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8681), .ZN(n7635) );
  NAND2_X1 U9466 ( .A1(n7636), .A2(n7635), .ZN(P2_U3220) );
  INV_X1 U9467 ( .A(n7637), .ZN(n7640) );
  OAI222_X1 U9468 ( .A1(P2_U3151), .A2(n6244), .B1(n8822), .B2(n7640), .C1(
        n7638), .C2(n8816), .ZN(P2_U3270) );
  OAI222_X1 U9469 ( .A1(P1_U3086), .A2(n7641), .B1(n9993), .B2(n7640), .C1(
        n7639), .C2(n9995), .ZN(P1_U3330) );
  NOR2_X1 U9470 ( .A1(n8132), .A2(n4696), .ZN(n8056) );
  XNOR2_X1 U9471 ( .A(n7642), .B(n8056), .ZN(n7649) );
  INV_X1 U9472 ( .A(n7649), .ZN(n7683) );
  XOR2_X1 U9473 ( .A(n7644), .B(n8056), .Z(n7645) );
  NAND2_X1 U9474 ( .A1(n7645), .A2(n8640), .ZN(n7647) );
  AOI22_X1 U9475 ( .A1(n8573), .A2(n8271), .B1(n8269), .B2(n8571), .ZN(n7646)
         );
  OAI211_X1 U9476 ( .C1(n7649), .C2(n7648), .A(n7647), .B(n7646), .ZN(n7680)
         );
  AOI21_X1 U9477 ( .B1(n10145), .B2(n7683), .A(n7680), .ZN(n7652) );
  MUX2_X1 U9478 ( .A(n7650), .B(n7652), .S(n10155), .Z(n7651) );
  OAI21_X1 U9479 ( .B1(n7767), .B2(n8747), .A(n7651), .ZN(P2_U3420) );
  MUX2_X1 U9480 ( .A(n8294), .B(n7652), .S(n10168), .Z(n7653) );
  OAI21_X1 U9481 ( .B1(n7767), .B2(n8696), .A(n7653), .ZN(P2_U3469) );
  OAI222_X1 U9482 ( .A1(P2_U3151), .A2(n6243), .B1(n7670), .B2(n7655), .C1(
        n7654), .C2(n8816), .ZN(P2_U3271) );
  OR2_X1 U9483 ( .A1(n7656), .A2(n8150), .ZN(n7657) );
  NAND2_X1 U9484 ( .A1(n7658), .A2(n7657), .ZN(n7715) );
  NAND2_X1 U9485 ( .A1(n7595), .A2(n7659), .ZN(n7660) );
  XOR2_X1 U9486 ( .A(n7660), .B(n8150), .Z(n7661) );
  OAI222_X1 U9487 ( .A1(n8658), .A2(n7888), .B1(n8656), .B2(n7884), .C1(n7661), 
        .C2(n8653), .ZN(n7710) );
  NAND2_X1 U9488 ( .A1(n7710), .A2(n8663), .ZN(n7664) );
  INV_X1 U9489 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8333) );
  OAI22_X1 U9490 ( .A1(n8663), .A2(n8333), .B1(n7892), .B2(n8643), .ZN(n7662)
         );
  AOI21_X1 U9491 ( .B1(n8153), .B2(n8666), .A(n7662), .ZN(n7663) );
  OAI211_X1 U9492 ( .C1(n7715), .C2(n8669), .A(n7664), .B(n7663), .ZN(P2_U3221) );
  MUX2_X1 U9493 ( .A(n7675), .B(P2_REG0_REG_13__SCAN_IN), .S(n10156), .Z(n7665) );
  INV_X1 U9494 ( .A(n7665), .ZN(n7667) );
  AOI22_X1 U9495 ( .A1(n7677), .A2(n8802), .B1(n8801), .B2(n8157), .ZN(n7666)
         );
  NAND2_X1 U9496 ( .A1(n7667), .A2(n7666), .ZN(P2_U3429) );
  INV_X1 U9497 ( .A(n7668), .ZN(n7673) );
  OAI222_X1 U9498 ( .A1(P2_U3151), .A2(n7671), .B1(n7670), .B2(n7673), .C1(
        n7669), .C2(n8816), .ZN(P2_U3269) );
  OAI222_X1 U9499 ( .A1(n10066), .A2(n7674), .B1(n9993), .B2(n7673), .C1(n7672), .C2(n9995), .ZN(P1_U3329) );
  INV_X1 U9500 ( .A(n7675), .ZN(n7676) );
  MUX2_X1 U9501 ( .A(n7676), .B(n4789), .S(n10165), .Z(n7679) );
  AOI22_X1 U9502 ( .A1(n7677), .A2(n8734), .B1(n8733), .B2(n8157), .ZN(n7678)
         );
  NAND2_X1 U9503 ( .A1(n7679), .A2(n7678), .ZN(P2_U3472) );
  OAI22_X1 U9504 ( .A1(n8630), .A2(n7767), .B1(n7691), .B2(n8643), .ZN(n7682)
         );
  MUX2_X1 U9505 ( .A(n7680), .B(P2_REG2_REG_10__SCAN_IN), .S(n8681), .Z(n7681)
         );
  AOI211_X1 U9506 ( .C1(n7757), .C2(n7683), .A(n7682), .B(n7681), .ZN(n7684)
         );
  INV_X1 U9507 ( .A(n7684), .ZN(P2_U3223) );
  XNOR2_X1 U9508 ( .A(n7883), .B(n7882), .ZN(n7688) );
  NOR2_X1 U9509 ( .A1(n7688), .A2(n5002), .ZN(n7881) );
  AOI21_X1 U9510 ( .B1(n5002), .B2(n7688), .A(n7881), .ZN(n7695) );
  NAND2_X1 U9511 ( .A1(n8007), .A2(n8271), .ZN(n7690) );
  OAI211_X1 U9512 ( .C1(n7884), .C2(n8009), .A(n7690), .B(n7689), .ZN(n7693)
         );
  NOR2_X1 U9513 ( .A1(n7953), .A2(n7691), .ZN(n7692) );
  AOI211_X1 U9514 ( .C1(n7770), .C2(n7998), .A(n7693), .B(n7692), .ZN(n7694)
         );
  OAI21_X1 U9515 ( .B1(n7695), .B2(n8000), .A(n7694), .ZN(P2_U3157) );
  INV_X1 U9516 ( .A(n7697), .ZN(n8164) );
  XNOR2_X1 U9517 ( .A(n7696), .B(n8163), .ZN(n7698) );
  AOI222_X1 U9518 ( .A1(n7698), .A2(n8640), .B1(n8265), .B2(n8571), .C1(n8267), 
        .C2(n8573), .ZN(n8673) );
  MUX2_X1 U9519 ( .A(n7699), .B(n8673), .S(n10155), .Z(n7703) );
  XNOR2_X1 U9520 ( .A(n7701), .B(n8163), .ZN(n8679) );
  AOI22_X1 U9521 ( .A1(n8679), .A2(n8802), .B1(n8801), .B2(n7839), .ZN(n7702)
         );
  NAND2_X1 U9522 ( .A1(n7703), .A2(n7702), .ZN(P2_U3432) );
  MUX2_X1 U9523 ( .A(n7704), .B(n8673), .S(n10168), .Z(n7706) );
  AOI22_X1 U9524 ( .A1(n8679), .A2(n8734), .B1(n8733), .B2(n7839), .ZN(n7705)
         );
  NAND2_X1 U9525 ( .A1(n7706), .A2(n7705), .ZN(P2_U3473) );
  INV_X1 U9526 ( .A(n7707), .ZN(n7716) );
  OAI222_X1 U9527 ( .A1(n9995), .A2(n7709), .B1(n9993), .B2(n7716), .C1(n7708), 
        .C2(P1_U3086), .ZN(P1_U3328) );
  AOI21_X1 U9528 ( .B1(n10144), .B2(n8153), .A(n7710), .ZN(n7713) );
  MUX2_X1 U9529 ( .A(n7711), .B(n7713), .S(n10155), .Z(n7712) );
  OAI21_X1 U9530 ( .B1(n7715), .B2(n8790), .A(n7712), .ZN(P2_U3426) );
  MUX2_X1 U9531 ( .A(n8337), .B(n7713), .S(n10168), .Z(n7714) );
  OAI21_X1 U9532 ( .B1(n8716), .B2(n7715), .A(n7714), .ZN(P2_U3471) );
  OAI222_X1 U9533 ( .A1(n8816), .A2(n7717), .B1(P2_U3151), .B2(n8405), .C1(
        n8822), .C2(n7716), .ZN(P2_U3268) );
  INV_X1 U9534 ( .A(n7718), .ZN(n7719) );
  AOI21_X1 U9535 ( .B1(n7719), .B2(n8065), .A(n8653), .ZN(n7722) );
  OAI22_X1 U9536 ( .A1(n8637), .A2(n8658), .B1(n7838), .B2(n8656), .ZN(n7720)
         );
  AOI21_X1 U9537 ( .B1(n7722), .B2(n7721), .A(n7720), .ZN(n8740) );
  OAI21_X1 U9538 ( .B1(n8065), .B2(n7724), .A(n7723), .ZN(n8738) );
  INV_X1 U9539 ( .A(n8737), .ZN(n7726) );
  AOI22_X1 U9540 ( .A1(n8681), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8677), .B2(
        n7910), .ZN(n7725) );
  OAI21_X1 U9541 ( .B1(n7726), .B2(n8630), .A(n7725), .ZN(n7727) );
  AOI21_X1 U9542 ( .B1(n8738), .B2(n8678), .A(n7727), .ZN(n7728) );
  OAI21_X1 U9543 ( .B1(n8740), .B2(n8681), .A(n7728), .ZN(P2_U3217) );
  XNOR2_X1 U9544 ( .A(n7729), .B(n8061), .ZN(n7744) );
  INV_X1 U9545 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n7735) );
  INV_X1 U9546 ( .A(n7730), .ZN(n7731) );
  INV_X1 U9547 ( .A(n8061), .ZN(n8167) );
  AOI21_X1 U9548 ( .B1(n7731), .B2(n8167), .A(n8653), .ZN(n7734) );
  OAI22_X1 U9549 ( .A1(n8657), .A2(n8658), .B1(n7950), .B2(n8656), .ZN(n7732)
         );
  AOI21_X1 U9550 ( .B1(n7734), .B2(n7733), .A(n7732), .ZN(n7740) );
  MUX2_X1 U9551 ( .A(n7735), .B(n7740), .S(n10155), .Z(n7737) );
  NAND2_X1 U9552 ( .A1(n8002), .A2(n8801), .ZN(n7736) );
  OAI211_X1 U9553 ( .C1(n7744), .C2(n8790), .A(n7737), .B(n7736), .ZN(P2_U3435) );
  MUX2_X1 U9554 ( .A(n4728), .B(n7740), .S(n6405), .Z(n7739) );
  AOI22_X1 U9555 ( .A1(n8002), .A2(n8666), .B1(n8677), .B2(n8012), .ZN(n7738)
         );
  OAI211_X1 U9556 ( .C1(n7744), .C2(n8669), .A(n7739), .B(n7738), .ZN(P2_U3218) );
  INV_X1 U9557 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n7741) );
  MUX2_X1 U9558 ( .A(n7741), .B(n7740), .S(n10168), .Z(n7743) );
  NAND2_X1 U9559 ( .A1(n8002), .A2(n8733), .ZN(n7742) );
  OAI211_X1 U9560 ( .C1(n8716), .C2(n7744), .A(n7743), .B(n7742), .ZN(P2_U3474) );
  NAND2_X1 U9561 ( .A1(n7745), .A2(n10076), .ZN(n7747) );
  AOI22_X1 U9562 ( .A1(n9041), .A2(n10094), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n10084), .ZN(n7746) );
  OAI211_X1 U9563 ( .C1(n4808), .C2(n9836), .A(n7747), .B(n7746), .ZN(n7748)
         );
  AOI21_X1 U9564 ( .B1(n7749), .B2(n9855), .A(n7748), .ZN(n7750) );
  OAI21_X1 U9565 ( .B1(n7751), .B2(n9850), .A(n7750), .ZN(P1_U3265) );
  INV_X1 U9566 ( .A(n7752), .ZN(n7758) );
  NOR2_X1 U9567 ( .A1(n7753), .A2(n8643), .ZN(n8499) );
  AOI21_X1 U9568 ( .B1(n8681), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8499), .ZN(
        n7754) );
  OAI21_X1 U9569 ( .B1(n7755), .B2(n8630), .A(n7754), .ZN(n7756) );
  AOI21_X1 U9570 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7759) );
  OAI21_X1 U9571 ( .B1(n7760), .B2(n8681), .A(n7759), .ZN(P2_U3204) );
  INV_X1 U9572 ( .A(n7761), .ZN(n8823) );
  OAI222_X1 U9573 ( .A1(n7763), .A2(P1_U3086), .B1(n9993), .B2(n8823), .C1(
        n7762), .C2(n9995), .ZN(P1_U3327) );
  XNOR2_X1 U9574 ( .A(n8519), .B(n7772), .ZN(n7764) );
  XNOR2_X1 U9575 ( .A(n8505), .B(n7764), .ZN(n7821) );
  INV_X1 U9576 ( .A(n7821), .ZN(n7765) );
  NAND2_X1 U9577 ( .A1(n7765), .A2(n8003), .ZN(n7826) );
  XNOR2_X1 U9578 ( .A(n8058), .B(n7772), .ZN(n7968) );
  NAND2_X1 U9579 ( .A1(n5002), .A2(n8270), .ZN(n7766) );
  NOR3_X1 U9580 ( .A1(n7767), .A2(n8270), .A3(n7809), .ZN(n7769) );
  AOI211_X1 U9581 ( .C1(n7884), .C2(n7809), .A(n7769), .B(n7768), .ZN(n7774)
         );
  NOR3_X1 U9582 ( .A1(n7770), .A2(n7772), .A3(n8270), .ZN(n7771) );
  AOI211_X1 U9583 ( .C1(n7884), .C2(n7772), .A(n7771), .B(n8058), .ZN(n7773)
         );
  XNOR2_X1 U9584 ( .A(n8153), .B(n7813), .ZN(n7777) );
  XNOR2_X1 U9585 ( .A(n7777), .B(n8152), .ZN(n7886) );
  XNOR2_X1 U9586 ( .A(n8157), .B(n7772), .ZN(n7778) );
  NOR2_X1 U9587 ( .A1(n7778), .A2(n7888), .ZN(n7947) );
  XNOR2_X1 U9588 ( .A(n7839), .B(n7809), .ZN(n7779) );
  XNOR2_X1 U9589 ( .A(n7779), .B(n7950), .ZN(n7835) );
  INV_X1 U9590 ( .A(n7779), .ZN(n7780) );
  XNOR2_X1 U9591 ( .A(n8002), .B(n7813), .ZN(n7781) );
  XNOR2_X1 U9592 ( .A(n7781), .B(n7838), .ZN(n8005) );
  INV_X1 U9593 ( .A(n7781), .ZN(n7782) );
  XNOR2_X1 U9594 ( .A(n8737), .B(n7772), .ZN(n7916) );
  XNOR2_X1 U9595 ( .A(n8800), .B(n7809), .ZN(n7784) );
  NAND2_X1 U9596 ( .A1(n7784), .A2(n7783), .ZN(n7914) );
  OAI21_X1 U9597 ( .B1(n7916), .B2(n8657), .A(n7914), .ZN(n7787) );
  NAND3_X1 U9598 ( .A1(n7916), .A2(n8657), .A3(n7914), .ZN(n7786) );
  INV_X1 U9599 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U9600 ( .A1(n7785), .A2(n8637), .ZN(n7978) );
  XNOR2_X1 U9601 ( .A(n8711), .B(n7809), .ZN(n7794) );
  NAND2_X1 U9602 ( .A1(n7794), .A2(n8261), .ZN(n7867) );
  INV_X1 U9603 ( .A(n7867), .ZN(n7790) );
  XNOR2_X1 U9604 ( .A(n7854), .B(n7809), .ZN(n7858) );
  NAND2_X1 U9605 ( .A1(n7858), .A2(n8262), .ZN(n7938) );
  XNOR2_X1 U9606 ( .A(n8726), .B(n7809), .ZN(n7855) );
  NAND2_X1 U9607 ( .A1(n7855), .A2(n8263), .ZN(n7788) );
  INV_X1 U9608 ( .A(n7855), .ZN(n7791) );
  NAND2_X1 U9609 ( .A1(n7791), .A2(n8659), .ZN(n7859) );
  AOI21_X1 U9610 ( .B1(n8262), .B2(n7859), .A(n7858), .ZN(n7793) );
  NOR3_X1 U9611 ( .A1(n7855), .A2(n8262), .A3(n8263), .ZN(n7792) );
  OAI21_X1 U9612 ( .B1(n7793), .B2(n7792), .A(n7867), .ZN(n7796) );
  INV_X1 U9613 ( .A(n7794), .ZN(n7795) );
  NAND2_X1 U9614 ( .A1(n7795), .A2(n8621), .ZN(n7870) );
  XNOR2_X1 U9615 ( .A(n8706), .B(n7772), .ZN(n7798) );
  NAND2_X1 U9616 ( .A1(n7798), .A2(n8608), .ZN(n7802) );
  INV_X1 U9617 ( .A(n7798), .ZN(n7799) );
  NAND2_X1 U9618 ( .A1(n7799), .A2(n8260), .ZN(n7800) );
  AND2_X1 U9619 ( .A1(n7802), .A2(n7800), .ZN(n7871) );
  NAND2_X1 U9620 ( .A1(n7801), .A2(n7871), .ZN(n7873) );
  XNOR2_X1 U9621 ( .A(n8703), .B(n7813), .ZN(n7803) );
  XNOR2_X1 U9622 ( .A(n7803), .B(n8591), .ZN(n7960) );
  XNOR2_X1 U9623 ( .A(n8775), .B(n7809), .ZN(n7844) );
  XNOR2_X1 U9624 ( .A(n8769), .B(n7772), .ZN(n7805) );
  NAND2_X1 U9625 ( .A1(n7805), .A2(n7850), .ZN(n7808) );
  OAI21_X1 U9626 ( .B1(n7805), .B2(n7850), .A(n7808), .ZN(n7925) );
  AOI21_X1 U9627 ( .B1(n8553), .B2(n7844), .A(n7925), .ZN(n7806) );
  XNOR2_X1 U9628 ( .A(n8762), .B(n7809), .ZN(n7810) );
  XNOR2_X1 U9629 ( .A(n7810), .B(n8532), .ZN(n7898) );
  INV_X1 U9630 ( .A(n7810), .ZN(n7811) );
  NAND2_X1 U9631 ( .A1(n7811), .A2(n8532), .ZN(n7812) );
  XOR2_X1 U9632 ( .A(n7813), .B(n8756), .Z(n7992) );
  XNOR2_X1 U9633 ( .A(n7834), .B(n7772), .ZN(n7819) );
  NAND2_X1 U9634 ( .A1(n7819), .A2(n8259), .ZN(n7814) );
  OAI21_X1 U9635 ( .B1(n7819), .B2(n8259), .A(n7814), .ZN(n7828) );
  AND2_X1 U9636 ( .A1(n7821), .A2(n5006), .ZN(n7815) );
  NAND2_X1 U9637 ( .A1(n7830), .A2(n7815), .ZN(n7825) );
  AOI22_X1 U9638 ( .A1(n8504), .A2(n8011), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n7817) );
  NAND2_X1 U9639 ( .A1(n8259), .A2(n8007), .ZN(n7816) );
  OAI211_X1 U9640 ( .C1(n7818), .C2(n8009), .A(n7817), .B(n7816), .ZN(n7823)
         );
  INV_X1 U9641 ( .A(n7819), .ZN(n7820) );
  NOR4_X1 U9642 ( .A1(n7821), .A2(n7820), .A3(n8533), .A4(n8000), .ZN(n7822)
         );
  AOI211_X1 U9643 ( .C1(n8505), .C2(n7998), .A(n7823), .B(n7822), .ZN(n7824)
         );
  OAI211_X1 U9644 ( .C1(n7826), .C2(n7830), .A(n7825), .B(n7824), .ZN(P2_U3160) );
  INV_X1 U9645 ( .A(n8018), .ZN(n9994) );
  OAI222_X1 U9646 ( .A1(n8816), .A2(n8019), .B1(n8822), .B2(n9994), .C1(n7827), 
        .C2(P2_U3151), .ZN(P2_U3265) );
  INV_X1 U9647 ( .A(n8007), .ZN(n7986) );
  AOI22_X1 U9648 ( .A1(n8526), .A2(n8011), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n7831) );
  OAI21_X1 U9649 ( .B1(n7991), .B2(n7986), .A(n7831), .ZN(n7832) );
  AOI21_X1 U9650 ( .B1(n7984), .B2(n8519), .A(n7832), .ZN(n7833) );
  XOR2_X1 U9651 ( .A(n7836), .B(n7835), .Z(n7843) );
  NAND2_X1 U9652 ( .A1(n8007), .A2(n8267), .ZN(n7837) );
  NAND2_X1 U9653 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8369) );
  OAI211_X1 U9654 ( .C1(n7838), .C2(n8009), .A(n7837), .B(n8369), .ZN(n7841)
         );
  INV_X1 U9655 ( .A(n7839), .ZN(n8672) );
  NOR2_X1 U9656 ( .A1(n8672), .A2(n8015), .ZN(n7840) );
  AOI211_X1 U9657 ( .C1(n8676), .C2(n8011), .A(n7841), .B(n7840), .ZN(n7842)
         );
  OAI21_X1 U9658 ( .B1(n7843), .B2(n8000), .A(n7842), .ZN(P2_U3155) );
  INV_X1 U9659 ( .A(n7844), .ZN(n7845) );
  NAND2_X1 U9660 ( .A1(n7846), .A2(n7845), .ZN(n7926) );
  OAI21_X1 U9661 ( .B1(n7846), .B2(n7845), .A(n7926), .ZN(n7847) );
  NOR2_X1 U9662 ( .A1(n7847), .A2(n8553), .ZN(n7929) );
  AOI21_X1 U9663 ( .B1(n8553), .B2(n7847), .A(n7929), .ZN(n7853) );
  AOI22_X1 U9664 ( .A1(n8574), .A2(n8007), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n7849) );
  NAND2_X1 U9665 ( .A1(n8576), .A2(n8011), .ZN(n7848) );
  OAI211_X1 U9666 ( .C1(n7850), .C2(n8009), .A(n7849), .B(n7848), .ZN(n7851)
         );
  AOI21_X1 U9667 ( .B1(n8775), .B2(n7998), .A(n7851), .ZN(n7852) );
  OAI21_X1 U9668 ( .B1(n7853), .B2(n8000), .A(n7852), .ZN(P2_U3156) );
  INV_X1 U9669 ( .A(n7854), .ZN(n8720) );
  XNOR2_X1 U9670 ( .A(n7855), .B(n8659), .ZN(n7979) );
  NAND2_X1 U9671 ( .A1(n7856), .A2(n7979), .ZN(n7860) );
  INV_X1 U9672 ( .A(n7860), .ZN(n7982) );
  INV_X1 U9673 ( .A(n7859), .ZN(n7857) );
  NOR2_X1 U9674 ( .A1(n7982), .A2(n7857), .ZN(n7862) );
  XNOR2_X1 U9675 ( .A(n7858), .B(n8638), .ZN(n7861) );
  INV_X1 U9676 ( .A(n7869), .ZN(n7939) );
  OAI211_X1 U9677 ( .C1(n7862), .C2(n7861), .A(n7939), .B(n8003), .ZN(n7866)
         );
  NAND2_X1 U9678 ( .A1(n8007), .A2(n8263), .ZN(n7863) );
  NAND2_X1 U9679 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8485) );
  OAI211_X1 U9680 ( .C1(n8621), .C2(n8009), .A(n7863), .B(n8485), .ZN(n7864)
         );
  AOI21_X1 U9681 ( .B1(n8627), .B2(n8011), .A(n7864), .ZN(n7865) );
  OAI211_X1 U9682 ( .C1(n8720), .C2(n8015), .A(n7866), .B(n7865), .ZN(P2_U3159) );
  INV_X1 U9683 ( .A(n8706), .ZN(n7880) );
  INV_X1 U9684 ( .A(n7938), .ZN(n7868) );
  NAND2_X1 U9685 ( .A1(n7867), .A2(n7870), .ZN(n7936) );
  NOR3_X1 U9686 ( .A1(n7869), .A2(n7868), .A3(n7936), .ZN(n7941) );
  INV_X1 U9687 ( .A(n7870), .ZN(n7872) );
  NOR3_X1 U9688 ( .A1(n7941), .A2(n7872), .A3(n7871), .ZN(n7875) );
  INV_X1 U9689 ( .A(n7873), .ZN(n7874) );
  OAI21_X1 U9690 ( .B1(n7875), .B2(n7874), .A(n8003), .ZN(n7879) );
  AOI22_X1 U9691 ( .A1(n8574), .A2(n7984), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n7876) );
  OAI21_X1 U9692 ( .B1(n8621), .B2(n7986), .A(n7876), .ZN(n7877) );
  AOI21_X1 U9693 ( .B1(n8600), .B2(n8011), .A(n7877), .ZN(n7878) );
  OAI211_X1 U9694 ( .C1(n7880), .C2(n8015), .A(n7879), .B(n7878), .ZN(P2_U3163) );
  AOI21_X1 U9695 ( .B1(n7883), .B2(n7882), .A(n7881), .ZN(n7969) );
  NAND2_X1 U9696 ( .A1(n7969), .A2(n7968), .ZN(n7967) );
  OAI21_X1 U9697 ( .B1(n7884), .B2(n7968), .A(n7967), .ZN(n7885) );
  XOR2_X1 U9698 ( .A(n7886), .B(n7885), .Z(n7894) );
  NAND2_X1 U9699 ( .A1(n8153), .A2(n7998), .ZN(n7891) );
  NAND2_X1 U9700 ( .A1(n8007), .A2(n8269), .ZN(n7887) );
  NAND2_X1 U9701 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8308) );
  OAI211_X1 U9702 ( .C1(n7888), .C2(n8009), .A(n7887), .B(n8308), .ZN(n7889)
         );
  INV_X1 U9703 ( .A(n7889), .ZN(n7890) );
  OAI211_X1 U9704 ( .C1(n7892), .C2(n7953), .A(n7891), .B(n7890), .ZN(n7893)
         );
  AOI21_X1 U9705 ( .B1(n7894), .B2(n8003), .A(n7893), .ZN(n7895) );
  INV_X1 U9706 ( .A(n7895), .ZN(P2_U3164) );
  OAI21_X1 U9707 ( .B1(n7898), .B2(n7897), .A(n7896), .ZN(n7899) );
  NAND2_X1 U9708 ( .A1(n7899), .A2(n8003), .ZN(n7905) );
  INV_X1 U9709 ( .A(n7900), .ZN(n7902) );
  AOI22_X1 U9710 ( .A1(n8572), .A2(n8007), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n7901) );
  OAI21_X1 U9711 ( .B1(n7902), .B2(n7953), .A(n7901), .ZN(n7903) );
  AOI21_X1 U9712 ( .B1(n7984), .B2(n8520), .A(n7903), .ZN(n7904) );
  OAI211_X1 U9713 ( .C1(n8531), .C2(n8015), .A(n7905), .B(n7904), .ZN(P2_U3165) );
  XNOR2_X1 U9714 ( .A(n7916), .B(n8264), .ZN(n7907) );
  XNOR2_X1 U9715 ( .A(n7906), .B(n7907), .ZN(n7913) );
  NAND2_X1 U9716 ( .A1(n8007), .A2(n8265), .ZN(n7908) );
  NAND2_X1 U9717 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8406) );
  OAI211_X1 U9718 ( .C1(n8637), .C2(n8009), .A(n7908), .B(n8406), .ZN(n7909)
         );
  AOI21_X1 U9719 ( .B1(n7910), .B2(n8011), .A(n7909), .ZN(n7912) );
  NAND2_X1 U9720 ( .A1(n8737), .A2(n7998), .ZN(n7911) );
  OAI211_X1 U9721 ( .C1(n7913), .C2(n8000), .A(n7912), .B(n7911), .ZN(P2_U3166) );
  NAND2_X1 U9722 ( .A1(n7914), .A2(n7978), .ZN(n7919) );
  NOR2_X1 U9723 ( .A1(n7906), .A2(n8264), .ZN(n7917) );
  INV_X1 U9724 ( .A(n7906), .ZN(n7915) );
  OAI22_X1 U9725 ( .A1(n7917), .A2(n7916), .B1(n7915), .B2(n8657), .ZN(n7918)
         );
  NOR2_X1 U9726 ( .A1(n7918), .A2(n7919), .ZN(n7981) );
  AOI21_X1 U9727 ( .B1(n7919), .B2(n7918), .A(n7981), .ZN(n7924) );
  NAND2_X1 U9728 ( .A1(n8007), .A2(n8264), .ZN(n7920) );
  NAND2_X1 U9729 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U9730 ( .C1(n8659), .C2(n8009), .A(n7920), .B(n8433), .ZN(n7921)
         );
  AOI21_X1 U9731 ( .B1(n8665), .B2(n8011), .A(n7921), .ZN(n7923) );
  NAND2_X1 U9732 ( .A1(n8800), .A2(n7998), .ZN(n7922) );
  OAI211_X1 U9733 ( .C1(n7924), .C2(n8000), .A(n7923), .B(n7922), .ZN(P2_U3168) );
  INV_X1 U9734 ( .A(n8769), .ZN(n8697) );
  NAND2_X1 U9735 ( .A1(n7926), .A2(n7925), .ZN(n7928) );
  OAI21_X1 U9736 ( .B1(n7929), .B2(n7928), .A(n7927), .ZN(n7930) );
  NAND2_X1 U9737 ( .A1(n7930), .A2(n8003), .ZN(n7935) );
  INV_X1 U9738 ( .A(n8559), .ZN(n7932) );
  AOI22_X1 U9739 ( .A1(n8553), .A2(n8007), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n7931) );
  OAI21_X1 U9740 ( .B1(n7932), .B2(n7953), .A(n7931), .ZN(n7933) );
  AOI21_X1 U9741 ( .B1(n7984), .B2(n8554), .A(n7933), .ZN(n7934) );
  OAI211_X1 U9742 ( .C1(n8697), .C2(n8015), .A(n7935), .B(n7934), .ZN(P2_U3169) );
  INV_X1 U9743 ( .A(n8711), .ZN(n7946) );
  INV_X1 U9744 ( .A(n7936), .ZN(n7937) );
  AOI21_X1 U9745 ( .B1(n7939), .B2(n7938), .A(n7937), .ZN(n7940) );
  OAI21_X1 U9746 ( .B1(n7941), .B2(n7940), .A(n8003), .ZN(n7945) );
  AOI22_X1 U9747 ( .A1(n8260), .A2(n7984), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n7942) );
  OAI21_X1 U9748 ( .B1(n8638), .B2(n7986), .A(n7942), .ZN(n7943) );
  AOI21_X1 U9749 ( .B1(n8613), .B2(n8011), .A(n7943), .ZN(n7944) );
  OAI211_X1 U9750 ( .C1(n7946), .C2(n8015), .A(n7945), .B(n7944), .ZN(P2_U3173) );
  NOR2_X1 U9751 ( .A1(n7947), .A2(n4410), .ZN(n7948) );
  XNOR2_X1 U9752 ( .A(n7949), .B(n7948), .ZN(n7957) );
  NAND2_X1 U9753 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8347) );
  OAI21_X1 U9754 ( .B1(n8009), .B2(n7950), .A(n8347), .ZN(n7951) );
  AOI21_X1 U9755 ( .B1(n8007), .B2(n8268), .A(n7951), .ZN(n7952) );
  OAI21_X1 U9756 ( .B1(n7954), .B2(n7953), .A(n7952), .ZN(n7955) );
  AOI21_X1 U9757 ( .B1(n8157), .B2(n7998), .A(n7955), .ZN(n7956) );
  OAI21_X1 U9758 ( .B1(n7957), .B2(n8000), .A(n7956), .ZN(P2_U3174) );
  INV_X1 U9759 ( .A(n8703), .ZN(n7966) );
  OAI21_X1 U9760 ( .B1(n7960), .B2(n7959), .A(n7958), .ZN(n7961) );
  NAND2_X1 U9761 ( .A1(n7961), .A2(n8003), .ZN(n7965) );
  AOI22_X1 U9762 ( .A1(n8260), .A2(n8007), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n7962) );
  OAI21_X1 U9763 ( .B1(n8582), .B2(n8009), .A(n7962), .ZN(n7963) );
  AOI21_X1 U9764 ( .B1(n8583), .B2(n8011), .A(n7963), .ZN(n7964) );
  OAI211_X1 U9765 ( .C1(n7966), .C2(n8015), .A(n7965), .B(n7964), .ZN(P2_U3175) );
  OAI211_X1 U9766 ( .C1(n7969), .C2(n7968), .A(n7967), .B(n8003), .ZN(n7977)
         );
  NAND2_X1 U9767 ( .A1(n8007), .A2(n8270), .ZN(n7970) );
  NAND2_X1 U9768 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8283) );
  OAI211_X1 U9769 ( .C1(n8152), .C2(n8009), .A(n7970), .B(n8283), .ZN(n7974)
         );
  INV_X1 U9770 ( .A(n7971), .ZN(n7972) );
  NOR2_X1 U9771 ( .A1(n8015), .A2(n7972), .ZN(n7973) );
  AOI211_X1 U9772 ( .C1(n7975), .C2(n8011), .A(n7974), .B(n7973), .ZN(n7976)
         );
  NAND2_X1 U9773 ( .A1(n7977), .A2(n7976), .ZN(P2_U3176) );
  INV_X1 U9774 ( .A(n8726), .ZN(n7990) );
  INV_X1 U9775 ( .A(n7978), .ZN(n7980) );
  NOR3_X1 U9776 ( .A1(n7981), .A2(n7980), .A3(n7979), .ZN(n7983) );
  OAI21_X1 U9777 ( .B1(n7983), .B2(n7982), .A(n8003), .ZN(n7989) );
  AND2_X1 U9778 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8458) );
  AOI21_X1 U9779 ( .B1(n8262), .B2(n7984), .A(n8458), .ZN(n7985) );
  OAI21_X1 U9780 ( .B1(n7986), .B2(n8637), .A(n7985), .ZN(n7987) );
  AOI21_X1 U9781 ( .B1(n8642), .B2(n8011), .A(n7987), .ZN(n7988) );
  OAI211_X1 U9782 ( .C1(n7990), .C2(n8015), .A(n7989), .B(n7988), .ZN(P2_U3178) );
  XNOR2_X1 U9783 ( .A(n7992), .B(n7991), .ZN(n7993) );
  XNOR2_X1 U9784 ( .A(n7994), .B(n7993), .ZN(n8001) );
  AOI22_X1 U9785 ( .A1(n8545), .A2(n8011), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n7996) );
  NAND2_X1 U9786 ( .A1(n8554), .A2(n8007), .ZN(n7995) );
  OAI211_X1 U9787 ( .C1(n8533), .C2(n8009), .A(n7996), .B(n7995), .ZN(n7997)
         );
  AOI21_X1 U9788 ( .B1(n8756), .B2(n7998), .A(n7997), .ZN(n7999) );
  OAI21_X1 U9789 ( .B1(n8001), .B2(n8000), .A(n7999), .ZN(P2_U3180) );
  INV_X1 U9790 ( .A(n8002), .ZN(n8016) );
  OAI211_X1 U9791 ( .C1(n8006), .C2(n8005), .A(n8004), .B(n8003), .ZN(n8014)
         );
  NAND2_X1 U9792 ( .A1(n8007), .A2(n8266), .ZN(n8008) );
  NAND2_X1 U9793 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8386) );
  OAI211_X1 U9794 ( .C1(n8657), .C2(n8009), .A(n8008), .B(n8386), .ZN(n8010)
         );
  AOI21_X1 U9795 ( .B1(n8012), .B2(n8011), .A(n8010), .ZN(n8013) );
  OAI211_X1 U9796 ( .C1(n8016), .C2(n8015), .A(n8014), .B(n8013), .ZN(P2_U3181) );
  NAND2_X1 U9797 ( .A1(n8018), .A2(n4560), .ZN(n8021) );
  OR2_X1 U9798 ( .A1(n4474), .A2(n8019), .ZN(n8020) );
  AND2_X2 U9799 ( .A1(n8021), .A2(n8020), .ZN(n8748) );
  INV_X1 U9800 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8684) );
  NAND2_X1 U9801 ( .A1(n6057), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8024) );
  INV_X1 U9802 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8501) );
  OR2_X1 U9803 ( .A1(n8022), .A2(n8501), .ZN(n8023) );
  OAI211_X1 U9804 ( .C1(n5957), .C2(n8684), .A(n8024), .B(n8023), .ZN(n8025)
         );
  INV_X1 U9805 ( .A(n8025), .ZN(n8026) );
  NAND2_X1 U9806 ( .A1(n8809), .A2(n4560), .ZN(n8031) );
  OR2_X1 U9807 ( .A1(n4474), .A2(n8028), .ZN(n8030) );
  AOI21_X1 U9808 ( .B1(n8748), .B2(n8076), .A(n8742), .ZN(n8033) );
  INV_X1 U9809 ( .A(n8748), .ZN(n8035) );
  INV_X1 U9810 ( .A(n8258), .ZN(n8034) );
  NAND2_X1 U9811 ( .A1(n8035), .A2(n8034), .ZN(n8073) );
  NAND2_X1 U9812 ( .A1(n8073), .A2(n8032), .ZN(n8230) );
  NOR2_X1 U9813 ( .A1(n8033), .A2(n8230), .ZN(n8037) );
  NOR2_X1 U9814 ( .A1(n8035), .A2(n8034), .ZN(n8072) );
  NOR2_X1 U9815 ( .A1(n8040), .A2(n8039), .ZN(n8250) );
  INV_X1 U9816 ( .A(n8562), .ZN(n8041) );
  NAND2_X1 U9817 ( .A1(n8079), .A2(n8042), .ZN(n8172) );
  INV_X1 U9818 ( .A(n8043), .ZN(n8055) );
  NAND3_X1 U9819 ( .A1(n8045), .A2(n8044), .A3(n8100), .ZN(n8047) );
  OR2_X1 U9820 ( .A1(n8047), .A2(n8046), .ZN(n8052) );
  NAND4_X1 U9821 ( .A1(n8090), .A2(n8050), .A3(n8049), .A4(n8048), .ZN(n8051)
         );
  NOR2_X1 U9822 ( .A1(n8052), .A2(n8051), .ZN(n8054) );
  AND4_X1 U9823 ( .A1(n8056), .A2(n8055), .A3(n8054), .A4(n8053), .ZN(n8057)
         );
  NAND4_X1 U9824 ( .A1(n8059), .A2(n8058), .A3(n8057), .A4(n8150), .ZN(n8060)
         );
  OR4_X1 U9825 ( .A1(n8172), .A2(n8061), .A3(n8163), .A4(n8060), .ZN(n8063) );
  NAND2_X1 U9826 ( .A1(n8173), .A2(n8062), .ZN(n8181) );
  NOR2_X1 U9827 ( .A1(n8063), .A2(n8181), .ZN(n8064) );
  NAND4_X1 U9828 ( .A1(n8611), .A2(n8625), .A3(n8065), .A4(n8064), .ZN(n8066)
         );
  INV_X1 U9829 ( .A(n8067), .ZN(n8218) );
  NAND2_X1 U9830 ( .A1(n8199), .A2(n8204), .ZN(n8563) );
  INV_X1 U9831 ( .A(n8072), .ZN(n8234) );
  NOR2_X1 U9832 ( .A1(n8742), .A2(n8076), .ZN(n8231) );
  INV_X1 U9833 ( .A(n8231), .ZN(n8069) );
  NAND2_X1 U9834 ( .A1(n8742), .A2(n8076), .ZN(n8236) );
  INV_X1 U9835 ( .A(n8236), .ZN(n8070) );
  NAND2_X1 U9836 ( .A1(n8243), .A2(n4397), .ZN(n8249) );
  AOI21_X1 U9837 ( .B1(n8235), .B2(n8073), .A(n8072), .ZN(n8074) );
  NAND2_X1 U9838 ( .A1(n8074), .A2(n8498), .ZN(n8077) );
  INV_X1 U9839 ( .A(n8074), .ZN(n8075) );
  AOI22_X1 U9840 ( .A1(n8077), .A2(n8742), .B1(n8076), .B2(n8075), .ZN(n8240)
         );
  MUX2_X1 U9841 ( .A(n8078), .B(n8239), .S(n8222), .Z(n8228) );
  INV_X1 U9842 ( .A(n8079), .ZN(n8175) );
  NAND2_X1 U9843 ( .A1(n8082), .A2(n6213), .ZN(n8081) );
  NAND2_X1 U9844 ( .A1(n8081), .A2(n8222), .ZN(n8085) );
  NAND2_X1 U9845 ( .A1(n8080), .A2(n8083), .ZN(n8084) );
  NAND2_X1 U9846 ( .A1(n8085), .A2(n8084), .ZN(n8086) );
  OAI21_X1 U9847 ( .B1(n6213), .B2(n8087), .A(n8086), .ZN(n8089) );
  OAI211_X1 U9848 ( .C1(n8235), .C2(n8080), .A(n8091), .B(n8090), .ZN(n8099)
         );
  NAND2_X1 U9849 ( .A1(n8102), .A2(n8092), .ZN(n8096) );
  NAND2_X1 U9850 ( .A1(n8094), .A2(n8093), .ZN(n8095) );
  MUX2_X1 U9851 ( .A(n8096), .B(n8095), .S(n8222), .Z(n8097) );
  INV_X1 U9852 ( .A(n8097), .ZN(n8098) );
  NAND2_X1 U9853 ( .A1(n8099), .A2(n8098), .ZN(n8101) );
  NAND2_X1 U9854 ( .A1(n8101), .A2(n8100), .ZN(n8112) );
  INV_X1 U9855 ( .A(n8102), .ZN(n8105) );
  OAI211_X1 U9856 ( .C1(n8112), .C2(n8105), .A(n8104), .B(n8103), .ZN(n8107)
         );
  NAND3_X1 U9857 ( .A1(n8107), .A2(n8106), .A3(n8110), .ZN(n8108) );
  NAND2_X1 U9858 ( .A1(n10139), .A2(n8276), .ZN(n8109) );
  OAI211_X1 U9859 ( .C1(n8112), .C2(n8111), .A(n8110), .B(n8109), .ZN(n8113)
         );
  NAND2_X1 U9860 ( .A1(n8128), .A2(n8129), .ZN(n8133) );
  NAND2_X1 U9861 ( .A1(n8133), .A2(n8222), .ZN(n8121) );
  AND2_X1 U9862 ( .A1(n8135), .A2(n8139), .ZN(n8120) );
  NAND2_X1 U9863 ( .A1(n8121), .A2(n8120), .ZN(n8131) );
  NAND3_X1 U9864 ( .A1(n8123), .A2(n8122), .A3(n8222), .ZN(n8124) );
  NAND2_X1 U9865 ( .A1(n8125), .A2(n8124), .ZN(n8126) );
  AND2_X1 U9866 ( .A1(n8128), .A2(n8127), .ZN(n8130) );
  OAI211_X1 U9867 ( .C1(n8131), .C2(n8130), .A(n8129), .B(n8143), .ZN(n8141)
         );
  INV_X1 U9868 ( .A(n8132), .ZN(n8144) );
  INV_X1 U9869 ( .A(n8133), .ZN(n8137) );
  NAND2_X1 U9870 ( .A1(n8135), .A2(n8134), .ZN(n8136) );
  NAND2_X1 U9871 ( .A1(n8137), .A2(n8136), .ZN(n8138) );
  NAND3_X1 U9872 ( .A1(n8144), .A2(n8139), .A3(n8138), .ZN(n8140) );
  MUX2_X1 U9873 ( .A(n8141), .B(n8140), .S(n8222), .Z(n8142) );
  NAND2_X1 U9874 ( .A1(n8148), .A2(n8143), .ZN(n8146) );
  NAND2_X1 U9875 ( .A1(n8147), .A2(n8144), .ZN(n8145) );
  MUX2_X1 U9876 ( .A(n8146), .B(n8145), .S(n8235), .Z(n8151) );
  MUX2_X1 U9877 ( .A(n8148), .B(n8147), .S(n8222), .Z(n8149) );
  NAND2_X1 U9878 ( .A1(n8153), .A2(n8152), .ZN(n8154) );
  MUX2_X1 U9879 ( .A(n8155), .B(n8154), .S(n8222), .Z(n8156) );
  MUX2_X1 U9880 ( .A(n8267), .B(n8157), .S(n8235), .Z(n8158) );
  INV_X1 U9881 ( .A(n8158), .ZN(n8159) );
  INV_X1 U9882 ( .A(n8161), .ZN(n8162) );
  MUX2_X1 U9883 ( .A(n8165), .B(n8164), .S(n8222), .Z(n8166) );
  NAND3_X1 U9884 ( .A1(n8178), .A2(n8179), .A3(n8169), .ZN(n8170) );
  INV_X1 U9885 ( .A(n8171), .ZN(n8654) );
  MUX2_X1 U9886 ( .A(n8175), .B(n8174), .S(n8235), .Z(n8187) );
  NAND3_X1 U9887 ( .A1(n8178), .A2(n8177), .A3(n8176), .ZN(n8180) );
  NAND3_X1 U9888 ( .A1(n8180), .A2(n8179), .A3(n8222), .ZN(n8182) );
  AOI21_X1 U9889 ( .B1(n8183), .B2(n8182), .A(n8181), .ZN(n8185) );
  OR2_X1 U9890 ( .A1(n8185), .A2(n8184), .ZN(n8186) );
  AND2_X1 U9891 ( .A1(n8596), .A2(n8188), .ZN(n8190) );
  AND2_X1 U9892 ( .A1(n8611), .A2(n8594), .ZN(n8189) );
  MUX2_X1 U9893 ( .A(n8190), .B(n8189), .S(n8222), .Z(n8191) );
  NAND2_X1 U9894 ( .A1(n8192), .A2(n8222), .ZN(n8193) );
  INV_X1 U9895 ( .A(n8590), .ZN(n8598) );
  NAND2_X1 U9896 ( .A1(n8201), .A2(n8595), .ZN(n8195) );
  NAND2_X1 U9897 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  NAND4_X1 U9898 ( .A1(n6296), .A2(n8235), .A3(n8199), .A4(n8198), .ZN(n8214)
         );
  NAND3_X1 U9899 ( .A1(n8202), .A2(n4541), .A3(n8201), .ZN(n8213) );
  OAI211_X1 U9900 ( .C1(n8206), .C2(n8572), .A(n8697), .B(n8222), .ZN(n8210)
         );
  NAND2_X1 U9901 ( .A1(n8562), .A2(n8572), .ZN(n8205) );
  NAND3_X1 U9902 ( .A1(n8205), .A2(n8769), .A3(n8235), .ZN(n8209) );
  OR3_X1 U9903 ( .A1(n8562), .A2(n8572), .A3(n8222), .ZN(n8208) );
  NAND3_X1 U9904 ( .A1(n8206), .A2(n8572), .A3(n8222), .ZN(n8207) );
  NAND4_X1 U9905 ( .A1(n8210), .A2(n8209), .A3(n8208), .A4(n8207), .ZN(n8211)
         );
  MUX2_X1 U9906 ( .A(n8216), .B(n8215), .S(n8235), .Z(n8217) );
  INV_X1 U9907 ( .A(n8540), .ZN(n8546) );
  MUX2_X1 U9908 ( .A(n8219), .B(n8218), .S(n8235), .Z(n8220) );
  MUX2_X1 U9909 ( .A(n8224), .B(n8223), .S(n8222), .Z(n8225) );
  INV_X1 U9910 ( .A(n8225), .ZN(n8226) );
  OAI21_X1 U9911 ( .B1(n8227), .B2(n8228), .A(n8229), .ZN(n8238) );
  INV_X1 U9912 ( .A(n8238), .ZN(n8232) );
  NAND4_X1 U9913 ( .A1(n8236), .A2(n8235), .A3(n8234), .A4(n8233), .ZN(n8237)
         );
  NOR3_X1 U9914 ( .A1(n8243), .A2(n6259), .A3(n8242), .ZN(n8244) );
  AOI211_X2 U9915 ( .C1(n8246), .C2(n8245), .A(n8244), .B(n8254), .ZN(n8247)
         );
  NAND3_X1 U9916 ( .A1(n8252), .A2(n8251), .A3(n8405), .ZN(n8253) );
  OAI211_X1 U9917 ( .C1(n8255), .C2(n8254), .A(n8253), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8256) );
  NAND2_X1 U9918 ( .A1(n8257), .A2(n8256), .ZN(P2_U3296) );
  MUX2_X1 U9919 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8498), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U9920 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8258), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U9921 ( .A(n8519), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8457), .Z(
        P2_U3519) );
  MUX2_X1 U9922 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8259), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9923 ( .A(n8520), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8457), .Z(
        P2_U3517) );
  MUX2_X1 U9924 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8554), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9925 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8572), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U9926 ( .A(n8553), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8457), .Z(
        P2_U3514) );
  MUX2_X1 U9927 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8574), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9928 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8260), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8261), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8262), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U9931 ( .A(n8263), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8457), .Z(
        P2_U3509) );
  MUX2_X1 U9932 ( .A(n8264), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8457), .Z(
        P2_U3507) );
  MUX2_X1 U9933 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8265), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9934 ( .A(n8266), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8457), .Z(
        P2_U3505) );
  MUX2_X1 U9935 ( .A(n8267), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8457), .Z(
        P2_U3504) );
  MUX2_X1 U9936 ( .A(n8268), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8457), .Z(
        P2_U3503) );
  MUX2_X1 U9937 ( .A(n8269), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8457), .Z(
        P2_U3502) );
  MUX2_X1 U9938 ( .A(n8270), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8457), .Z(
        P2_U3501) );
  MUX2_X1 U9939 ( .A(n8271), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8457), .Z(
        P2_U3500) );
  MUX2_X1 U9940 ( .A(n8272), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8457), .Z(
        P2_U3499) );
  MUX2_X1 U9941 ( .A(n8273), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8457), .Z(
        P2_U3498) );
  MUX2_X1 U9942 ( .A(n8274), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8457), .Z(
        P2_U3497) );
  MUX2_X1 U9943 ( .A(n8275), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8457), .Z(
        P2_U3496) );
  MUX2_X1 U9944 ( .A(n8276), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8457), .Z(
        P2_U3495) );
  MUX2_X1 U9945 ( .A(n6271), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8457), .Z(
        P2_U3494) );
  MUX2_X1 U9946 ( .A(n8277), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8457), .Z(
        P2_U3492) );
  MUX2_X1 U9947 ( .A(n8278), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8457), .Z(
        P2_U3491) );
  MUX2_X1 U9948 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8405), .Z(n8303) );
  XNOR2_X1 U9949 ( .A(n8303), .B(n8305), .ZN(n8306) );
  XOR2_X1 U9950 ( .A(n8307), .B(n8306), .Z(n8302) );
  INV_X1 U9951 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8284) );
  OAI21_X1 U9952 ( .B1(n8371), .B2(n8284), .A(n8283), .ZN(n8293) );
  INV_X1 U9953 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8286) );
  NAND2_X1 U9954 ( .A1(n8287), .A2(n8298), .ZN(n8310) );
  AOI21_X1 U9955 ( .B1(n8290), .B2(n8289), .A(n8313), .ZN(n8291) );
  NOR2_X1 U9956 ( .A1(n8291), .A2(n8495), .ZN(n8292) );
  AOI211_X1 U9957 ( .C1(n8373), .C2(n8305), .A(n8293), .B(n8292), .ZN(n8301)
         );
  OR2_X1 U9958 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  OAI21_X1 U9959 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n4408), .A(n8317), .ZN(
        n8299) );
  NAND2_X1 U9960 ( .A1(n8299), .A2(n8492), .ZN(n8300) );
  OAI211_X1 U9961 ( .C1(n8302), .C2(n8482), .A(n8301), .B(n8300), .ZN(P2_U3193) );
  MUX2_X1 U9962 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8405), .Z(n8330) );
  XOR2_X1 U9963 ( .A(n8330), .B(n8338), .Z(n8331) );
  INV_X1 U9964 ( .A(n8303), .ZN(n8304) );
  XOR2_X1 U9965 ( .A(n8332), .B(n8331), .Z(n8328) );
  INV_X1 U9966 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8309) );
  OAI21_X1 U9967 ( .B1(n8371), .B2(n8309), .A(n8308), .ZN(n8316) );
  INV_X1 U9968 ( .A(n8310), .ZN(n8312) );
  XNOR2_X1 U9969 ( .A(n8338), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8311) );
  OR3_X1 U9970 ( .A1(n8313), .A2(n8312), .A3(n8311), .ZN(n8314) );
  AOI21_X1 U9971 ( .B1(n8335), .B2(n8314), .A(n8495), .ZN(n8315) );
  AOI211_X1 U9972 ( .C1(n8373), .C2(n8338), .A(n8316), .B(n8315), .ZN(n8327)
         );
  INV_X1 U9973 ( .A(n8317), .ZN(n8319) );
  INV_X1 U9974 ( .A(n8320), .ZN(n8318) );
  XNOR2_X1 U9975 ( .A(n8338), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8322) );
  NOR3_X1 U9976 ( .A1(n8319), .A2(n8318), .A3(n8322), .ZN(n8325) );
  NAND2_X1 U9977 ( .A1(n8321), .A2(n8320), .ZN(n8323) );
  NAND2_X1 U9978 ( .A1(n8323), .A2(n8322), .ZN(n8340) );
  INV_X1 U9979 ( .A(n8340), .ZN(n8324) );
  OAI21_X1 U9980 ( .B1(n8325), .B2(n8324), .A(n8492), .ZN(n8326) );
  OAI211_X1 U9981 ( .C1(n8328), .C2(n8482), .A(n8327), .B(n8326), .ZN(P2_U3194) );
  MUX2_X1 U9982 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8405), .Z(n8353) );
  XNOR2_X1 U9983 ( .A(n8353), .B(n8355), .ZN(n8356) );
  XOR2_X1 U9984 ( .A(n8356), .B(n8357), .Z(n8352) );
  OAI21_X1 U9985 ( .B1(n4403), .B2(P2_REG2_REG_13__SCAN_IN), .A(n8365), .ZN(
        n8346) );
  OR2_X1 U9986 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  NAND2_X1 U9987 ( .A1(n8340), .A2(n8339), .ZN(n8342) );
  OAI21_X1 U9988 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n4395), .A(n8359), .ZN(
        n8344) );
  AOI22_X1 U9989 ( .A1(n8346), .A2(n8345), .B1(n8492), .B2(n8344), .ZN(n8351)
         );
  INV_X1 U9990 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8348) );
  OAI21_X1 U9991 ( .B1(n8371), .B2(n8348), .A(n8347), .ZN(n8349) );
  AOI21_X1 U9992 ( .B1(n8355), .B2(n8373), .A(n8349), .ZN(n8350) );
  OAI211_X1 U9993 ( .C1(n8352), .C2(n8482), .A(n8351), .B(n8350), .ZN(P2_U3195) );
  MUX2_X1 U9994 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8405), .Z(n8383) );
  XOR2_X1 U9995 ( .A(n8378), .B(n8383), .Z(n8384) );
  INV_X1 U9996 ( .A(n8353), .ZN(n8354) );
  XOR2_X1 U9997 ( .A(n8384), .B(n8385), .Z(n8376) );
  NAND3_X1 U9998 ( .A1(n8359), .A2(n4418), .A3(n8358), .ZN(n8360) );
  NAND2_X1 U9999 ( .A1(n8393), .A2(n8360), .ZN(n8368) );
  NAND2_X1 U10000 ( .A1(n8365), .A2(n8363), .ZN(n8361) );
  XNOR2_X1 U10001 ( .A(n8378), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n8362) );
  NAND2_X1 U10002 ( .A1(n8361), .A2(n8362), .ZN(n8379) );
  INV_X1 U10003 ( .A(n8362), .ZN(n8364) );
  NAND3_X1 U10004 ( .A1(n8365), .A2(n8364), .A3(n8363), .ZN(n8366) );
  AOI21_X1 U10005 ( .B1(n8379), .B2(n8366), .A(n8495), .ZN(n8367) );
  AOI21_X1 U10006 ( .B1(n8492), .B2(n8368), .A(n8367), .ZN(n8375) );
  INV_X1 U10007 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8370) );
  OAI21_X1 U10008 ( .B1(n8371), .B2(n8370), .A(n8369), .ZN(n8372) );
  AOI21_X1 U10009 ( .B1(n8378), .B2(n8373), .A(n8372), .ZN(n8374) );
  OAI211_X1 U10010 ( .C1(n8376), .C2(n8482), .A(n8375), .B(n8374), .ZN(
        P2_U3196) );
  NAND2_X1 U10011 ( .A1(n8380), .A2(n8388), .ZN(n8408) );
  OAI21_X1 U10012 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n4332), .A(n8409), .ZN(
        n8382) );
  INV_X1 U10013 ( .A(n8382), .ZN(n8399) );
  MUX2_X1 U10014 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8405), .Z(n8400) );
  XNOR2_X1 U10015 ( .A(n8400), .B(n8402), .ZN(n8403) );
  XNOR2_X1 U10016 ( .A(n8404), .B(n8403), .ZN(n8390) );
  NAND2_X1 U10017 ( .A1(n8484), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n8387) );
  OAI211_X1 U10018 ( .C1(n8488), .C2(n8388), .A(n8387), .B(n8386), .ZN(n8389)
         );
  AOI21_X1 U10019 ( .B1(n8390), .B2(n8436), .A(n8389), .ZN(n8398) );
  NAND2_X1 U10020 ( .A1(n8391), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8392) );
  AOI21_X1 U10021 ( .B1(n8394), .B2(n8402), .A(n8414), .ZN(n8395) );
  NAND2_X1 U10022 ( .A1(n8395), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8418) );
  OAI21_X1 U10023 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n8395), .A(n8418), .ZN(
        n8396) );
  NAND2_X1 U10024 ( .A1(n8396), .A2(n8492), .ZN(n8397) );
  OAI211_X1 U10025 ( .C1(n8399), .C2(n8495), .A(n8398), .B(n8397), .ZN(
        P2_U3197) );
  INV_X1 U10026 ( .A(n8400), .ZN(n8401) );
  AOI22_X1 U10027 ( .A1(n8404), .A2(n8403), .B1(n8402), .B2(n8401), .ZN(n8432)
         );
  MUX2_X1 U10028 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8405), .Z(n8430) );
  XOR2_X1 U10029 ( .A(n8424), .B(n8430), .Z(n8431) );
  XNOR2_X1 U10030 ( .A(n8432), .B(n8431), .ZN(n8413) );
  NAND2_X1 U10031 ( .A1(n8484), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n8407) );
  OAI211_X1 U10032 ( .C1(n8488), .C2(n8438), .A(n8407), .B(n8406), .ZN(n8412)
         );
  NAND3_X1 U10033 ( .A1(n8409), .A2(n4419), .A3(n8408), .ZN(n8410) );
  AOI21_X1 U10034 ( .B1(n8422), .B2(n8410), .A(n8495), .ZN(n8411) );
  AOI211_X1 U10035 ( .C1(n8436), .C2(n8413), .A(n8412), .B(n8411), .ZN(n8421)
         );
  INV_X1 U10036 ( .A(n8414), .ZN(n8416) );
  INV_X1 U10037 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8415) );
  XNOR2_X1 U10038 ( .A(n8424), .B(n8415), .ZN(n8417) );
  AND3_X1 U10039 ( .A1(n8418), .A2(n8417), .A3(n8416), .ZN(n8419) );
  OAI21_X1 U10040 ( .B1(n4766), .B2(n8419), .A(n8492), .ZN(n8420) );
  NAND2_X1 U10041 ( .A1(n8421), .A2(n8420), .ZN(P2_U3198) );
  INV_X1 U10042 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8664) );
  INV_X1 U10043 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8423) );
  INV_X1 U10044 ( .A(n8425), .ZN(n8426) );
  NAND2_X1 U10045 ( .A1(n8426), .A2(n8451), .ZN(n8427) );
  INV_X1 U10046 ( .A(n8447), .ZN(n8428) );
  AOI21_X1 U10047 ( .B1(n8664), .B2(n8429), .A(n8428), .ZN(n8443) );
  MUX2_X1 U10048 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n8405), .Z(n8449) );
  XNOR2_X1 U10049 ( .A(n8449), .B(n8451), .ZN(n8452) );
  XNOR2_X1 U10050 ( .A(n8453), .B(n8452), .ZN(n8437) );
  NAND2_X1 U10051 ( .A1(n8484), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8434) );
  OAI211_X1 U10052 ( .C1(n8488), .C2(n4765), .A(n8434), .B(n8433), .ZN(n8435)
         );
  AOI21_X1 U10053 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8442) );
  OAI21_X1 U10054 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n8439), .A(n8463), .ZN(
        n8440) );
  NAND2_X1 U10055 ( .A1(n8440), .A2(n8492), .ZN(n8441) );
  OAI211_X1 U10056 ( .C1(n8443), .C2(n8495), .A(n8442), .B(n8441), .ZN(
        P2_U3199) );
  INV_X1 U10057 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8645) );
  OR2_X1 U10058 ( .A1(n8475), .A2(n8645), .ZN(n8466) );
  NAND2_X1 U10059 ( .A1(n8475), .A2(n8645), .ZN(n8444) );
  NAND2_X1 U10060 ( .A1(n8466), .A2(n8444), .ZN(n8445) );
  AND3_X1 U10061 ( .A1(n8447), .A2(n8446), .A3(n8445), .ZN(n8448) );
  INV_X1 U10062 ( .A(n8449), .ZN(n8450) );
  AOI22_X1 U10063 ( .A1(n8453), .A2(n8452), .B1(n8451), .B2(n8450), .ZN(n8455)
         );
  MUX2_X1 U10064 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8405), .Z(n8454) );
  NAND2_X1 U10065 ( .A1(n8455), .A2(n8454), .ZN(n8474) );
  INV_X1 U10066 ( .A(n8474), .ZN(n8456) );
  INV_X1 U10067 ( .A(n8459), .ZN(n8462) );
  INV_X1 U10068 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8731) );
  OR2_X1 U10069 ( .A1(n8475), .A2(n8731), .ZN(n8469) );
  NAND2_X1 U10070 ( .A1(n8475), .A2(n8731), .ZN(n8460) );
  NAND2_X1 U10071 ( .A1(n8469), .A2(n8460), .ZN(n8461) );
  AOI21_X1 U10072 ( .B1(n8463), .B2(n8462), .A(n8461), .ZN(n8471) );
  AND3_X1 U10073 ( .A1(n8463), .A2(n8462), .A3(n8461), .ZN(n8464) );
  OAI21_X1 U10074 ( .B1(n8471), .B2(n8464), .A(n8492), .ZN(n8465) );
  XNOR2_X1 U10075 ( .A(n6259), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n8478) );
  XNOR2_X1 U10076 ( .A(n8468), .B(n8478), .ZN(n8496) );
  INV_X1 U10077 ( .A(n8469), .ZN(n8470) );
  NOR2_X1 U10078 ( .A1(n8471), .A2(n8470), .ZN(n8473) );
  XNOR2_X1 U10079 ( .A(n8487), .B(n8723), .ZN(n8479) );
  INV_X1 U10080 ( .A(n8479), .ZN(n8472) );
  XNOR2_X1 U10081 ( .A(n8473), .B(n8472), .ZN(n8493) );
  MUX2_X1 U10082 ( .A(n8479), .B(n8478), .S(n8477), .Z(n8480) );
  XNOR2_X1 U10083 ( .A(n8481), .B(n8480), .ZN(n8483) );
  NAND2_X1 U10084 ( .A1(n8484), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n8486) );
  OAI211_X1 U10085 ( .C1(n8488), .C2(n8487), .A(n8486), .B(n8485), .ZN(n8489)
         );
  INV_X1 U10086 ( .A(n8489), .ZN(n8490) );
  AOI21_X1 U10087 ( .B1(n8493), .B2(n8492), .A(n8491), .ZN(n8494) );
  OAI21_X1 U10088 ( .B1(n8496), .B2(n8495), .A(n8494), .ZN(P2_U3201) );
  NAND2_X1 U10089 ( .A1(n8742), .A2(n8666), .ZN(n8500) );
  AOI21_X1 U10090 ( .B1(n8743), .B2(n8663), .A(n8499), .ZN(n8503) );
  OAI211_X1 U10091 ( .C1(n8501), .C2(n8663), .A(n8500), .B(n8503), .ZN(
        P2_U3202) );
  NAND2_X1 U10092 ( .A1(n8681), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8502) );
  OAI211_X1 U10093 ( .C1(n8748), .C2(n8630), .A(n8503), .B(n8502), .ZN(
        P2_U3203) );
  AOI22_X1 U10094 ( .A1(n8504), .A2(n8677), .B1(n8681), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8507) );
  NAND2_X1 U10095 ( .A1(n8505), .A2(n8666), .ZN(n8506) );
  OAI211_X1 U10096 ( .C1(n8508), .C2(n8669), .A(n8507), .B(n8506), .ZN(n8509)
         );
  INV_X1 U10097 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8525) );
  NOR2_X2 U10098 ( .A1(n8515), .A2(n8514), .ZN(n8518) );
  XNOR2_X1 U10099 ( .A(n8518), .B(n8517), .ZN(n8524) );
  AOI21_X1 U10100 ( .B1(n8524), .B2(n8640), .A(n8523), .ZN(n8749) );
  MUX2_X1 U10101 ( .A(n8525), .B(n8749), .S(n8663), .Z(n8528) );
  AOI22_X1 U10102 ( .A1(n8751), .A2(n8666), .B1(n8677), .B2(n8526), .ZN(n8527)
         );
  INV_X1 U10103 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U10104 ( .A1(n8529), .A2(n8640), .ZN(n8530) );
  NOR2_X1 U10105 ( .A1(n8540), .A2(n8530), .ZN(n8538) );
  NAND4_X1 U10106 ( .A1(n8540), .A2(n8532), .A3(n8531), .A4(n8640), .ZN(n8536)
         );
  OAI22_X1 U10107 ( .A1(n8533), .A2(n8658), .B1(n8532), .B2(n8656), .ZN(n8534)
         );
  INV_X1 U10108 ( .A(n8534), .ZN(n8535) );
  NAND2_X1 U10109 ( .A1(n8536), .A2(n8535), .ZN(n8537) );
  AOI21_X1 U10110 ( .B1(n8539), .B2(n8538), .A(n8537), .ZN(n8543) );
  INV_X1 U10111 ( .A(n8539), .ZN(n8541) );
  NAND3_X1 U10112 ( .A1(n8541), .A2(n8640), .A3(n8540), .ZN(n8542) );
  AOI22_X1 U10113 ( .A1(n8756), .A2(n8666), .B1(n8677), .B2(n8545), .ZN(n8549)
         );
  XNOR2_X1 U10114 ( .A(n8547), .B(n8546), .ZN(n8757) );
  NAND2_X1 U10115 ( .A1(n8757), .A2(n8678), .ZN(n8548) );
  NAND3_X1 U10116 ( .A1(n8550), .A2(n8549), .A3(n8548), .ZN(P2_U3207) );
  NOR2_X1 U10117 ( .A1(n8697), .A2(n8671), .ZN(n8558) );
  NOR2_X1 U10118 ( .A1(n8552), .A2(n8551), .ZN(n8557) );
  OAI21_X1 U10119 ( .B1(n6389), .B2(n8563), .A(n8640), .ZN(n8556) );
  AOI22_X1 U10120 ( .A1(n8554), .A2(n8571), .B1(n8573), .B2(n8553), .ZN(n8555)
         );
  OAI21_X1 U10121 ( .B1(n8557), .B2(n8556), .A(n8555), .ZN(n8766) );
  AOI211_X1 U10122 ( .C1(n8677), .C2(n8559), .A(n8558), .B(n8766), .ZN(n8567)
         );
  NAND2_X1 U10123 ( .A1(n8561), .A2(n8562), .ZN(n8564) );
  XNOR2_X1 U10124 ( .A(n8564), .B(n8563), .ZN(n8772) );
  INV_X1 U10125 ( .A(n8772), .ZN(n8565) );
  AOI22_X1 U10126 ( .A1(n8565), .A2(n8678), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8681), .ZN(n8566) );
  OAI21_X1 U10127 ( .B1(n8567), .B2(n8681), .A(n8566), .ZN(P2_U3209) );
  XOR2_X1 U10128 ( .A(n8568), .B(n8570), .Z(n8778) );
  XNOR2_X1 U10129 ( .A(n8569), .B(n8570), .ZN(n8575) );
  AOI222_X1 U10130 ( .A1(n8575), .A2(n8640), .B1(n8574), .B2(n8573), .C1(n8572), .C2(n8571), .ZN(n8773) );
  MUX2_X1 U10131 ( .A(n10286), .B(n8773), .S(n6405), .Z(n8578) );
  AOI22_X1 U10132 ( .A1(n8775), .A2(n8666), .B1(n8677), .B2(n8576), .ZN(n8577)
         );
  OAI211_X1 U10133 ( .C1(n8778), .C2(n8669), .A(n8578), .B(n8577), .ZN(
        P2_U3210) );
  XNOR2_X1 U10134 ( .A(n8579), .B(n4541), .ZN(n8782) );
  XNOR2_X1 U10135 ( .A(n8580), .B(n4541), .ZN(n8581) );
  OAI222_X1 U10136 ( .A1(n8658), .A2(n8582), .B1(n8656), .B2(n8608), .C1(n8581), .C2(n8653), .ZN(n8702) );
  NAND2_X1 U10137 ( .A1(n8702), .A2(n8663), .ZN(n8588) );
  INV_X1 U10138 ( .A(n8583), .ZN(n8585) );
  INV_X1 U10139 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8584) );
  OAI22_X1 U10140 ( .A1(n8585), .A2(n8643), .B1(n8663), .B2(n8584), .ZN(n8586)
         );
  AOI21_X1 U10141 ( .B1(n8703), .B2(n8666), .A(n8586), .ZN(n8587) );
  OAI211_X1 U10142 ( .C1(n8782), .C2(n8669), .A(n8588), .B(n8587), .ZN(
        P2_U3211) );
  XNOR2_X1 U10143 ( .A(n8589), .B(n8590), .ZN(n8593) );
  OAI22_X1 U10144 ( .A1(n8591), .A2(n8658), .B1(n8621), .B2(n8656), .ZN(n8592)
         );
  AOI21_X1 U10145 ( .B1(n8593), .B2(n8640), .A(n8592), .ZN(n8708) );
  NAND2_X1 U10146 ( .A1(n8626), .A2(n8625), .ZN(n8717) );
  NAND2_X1 U10147 ( .A1(n8717), .A2(n8594), .ZN(n8612) );
  INV_X1 U10148 ( .A(n8595), .ZN(n8597) );
  OAI21_X1 U10149 ( .B1(n8612), .B2(n8597), .A(n8596), .ZN(n8599) );
  XNOR2_X1 U10150 ( .A(n8599), .B(n8598), .ZN(n8785) );
  NAND2_X1 U10151 ( .A1(n8706), .A2(n8666), .ZN(n8602) );
  AOI22_X1 U10152 ( .A1(n8600), .A2(n8677), .B1(n8681), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n8601) );
  NAND2_X1 U10153 ( .A1(n8602), .A2(n8601), .ZN(n8603) );
  AOI21_X1 U10154 ( .B1(n8785), .B2(n8678), .A(n8603), .ZN(n8604) );
  OAI21_X1 U10155 ( .B1(n8708), .B2(n8681), .A(n8604), .ZN(P2_U3212) );
  NAND2_X1 U10156 ( .A1(n8605), .A2(n8611), .ZN(n8606) );
  NAND2_X1 U10157 ( .A1(n8607), .A2(n8606), .ZN(n8610) );
  OAI22_X1 U10158 ( .A1(n8608), .A2(n8658), .B1(n8638), .B2(n8656), .ZN(n8609)
         );
  AOI21_X1 U10159 ( .B1(n8610), .B2(n8640), .A(n8609), .ZN(n8713) );
  XNOR2_X1 U10160 ( .A(n8612), .B(n8611), .ZN(n8791) );
  AOI22_X1 U10161 ( .A1(n8681), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8613), .B2(
        n8677), .ZN(n8615) );
  NAND2_X1 U10162 ( .A1(n8711), .A2(n8666), .ZN(n8614) );
  OAI211_X1 U10163 ( .C1(n8791), .C2(n8669), .A(n8615), .B(n8614), .ZN(n8616)
         );
  INV_X1 U10164 ( .A(n8616), .ZN(n8617) );
  OAI21_X1 U10165 ( .B1(n8713), .B2(n8681), .A(n8617), .ZN(P2_U3213) );
  NAND2_X1 U10166 ( .A1(n8619), .A2(n8625), .ZN(n8620) );
  NAND3_X1 U10167 ( .A1(n8618), .A2(n8640), .A3(n8620), .ZN(n8624) );
  OAI22_X1 U10168 ( .A1(n8621), .A2(n8658), .B1(n8659), .B2(n8656), .ZN(n8622)
         );
  INV_X1 U10169 ( .A(n8622), .ZN(n8623) );
  NAND2_X1 U10170 ( .A1(n8624), .A2(n8623), .ZN(n8722) );
  OR2_X1 U10171 ( .A1(n8626), .A2(n8625), .ZN(n8718) );
  NAND3_X1 U10172 ( .A1(n8718), .A2(n8678), .A3(n8717), .ZN(n8629) );
  AOI22_X1 U10173 ( .A1(n8681), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8677), .B2(
        n8627), .ZN(n8628) );
  OAI211_X1 U10174 ( .C1(n8720), .C2(n8630), .A(n8629), .B(n8628), .ZN(n8631)
         );
  AOI21_X1 U10175 ( .B1(n8722), .B2(n8663), .A(n8631), .ZN(n8632) );
  INV_X1 U10176 ( .A(n8632), .ZN(P2_U3214) );
  NAND2_X1 U10177 ( .A1(n8633), .A2(n8634), .ZN(n8635) );
  NAND2_X1 U10178 ( .A1(n8636), .A2(n8635), .ZN(n8641) );
  OAI22_X1 U10179 ( .A1(n8638), .A2(n8658), .B1(n8637), .B2(n8656), .ZN(n8639)
         );
  AOI21_X1 U10180 ( .B1(n8641), .B2(n8640), .A(n8639), .ZN(n8730) );
  INV_X1 U10181 ( .A(n8642), .ZN(n8644) );
  OAI22_X1 U10182 ( .A1(n6405), .A2(n8645), .B1(n8644), .B2(n8643), .ZN(n8646)
         );
  AOI21_X1 U10183 ( .B1(n8726), .B2(n8666), .A(n8646), .ZN(n8650) );
  NAND2_X1 U10184 ( .A1(n8648), .A2(n6092), .ZN(n8725) );
  NAND3_X1 U10185 ( .A1(n8647), .A2(n8725), .A3(n8678), .ZN(n8649) );
  OAI211_X1 U10186 ( .C1(n8730), .C2(n8681), .A(n8650), .B(n8649), .ZN(
        P2_U3215) );
  XNOR2_X1 U10187 ( .A(n8651), .B(n8654), .ZN(n8803) );
  INV_X1 U10188 ( .A(n8803), .ZN(n8670) );
  INV_X1 U10189 ( .A(n8652), .ZN(n8655) );
  AOI21_X1 U10190 ( .B1(n8655), .B2(n8654), .A(n8653), .ZN(n8662) );
  OAI22_X1 U10191 ( .A1(n8659), .A2(n8658), .B1(n8657), .B2(n8656), .ZN(n8660)
         );
  AOI21_X1 U10192 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n8798) );
  MUX2_X1 U10193 ( .A(n8664), .B(n8798), .S(n8663), .Z(n8668) );
  AOI22_X1 U10194 ( .A1(n8800), .A2(n8666), .B1(n8677), .B2(n8665), .ZN(n8667)
         );
  OAI211_X1 U10195 ( .C1(n8670), .C2(n8669), .A(n8668), .B(n8667), .ZN(
        P2_U3216) );
  NOR2_X1 U10196 ( .A1(n8672), .A2(n8671), .ZN(n8675) );
  INV_X1 U10197 ( .A(n8673), .ZN(n8674) );
  AOI211_X1 U10198 ( .C1(n8677), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8682)
         );
  AOI22_X1 U10199 ( .A1(n8679), .A2(n8678), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n8681), .ZN(n8680) );
  OAI21_X1 U10200 ( .B1(n8682), .B2(n8681), .A(n8680), .ZN(P2_U3219) );
  NAND2_X1 U10201 ( .A1(n8742), .A2(n8733), .ZN(n8683) );
  NAND2_X1 U10202 ( .A1(n8743), .A2(n10168), .ZN(n8686) );
  OAI211_X1 U10203 ( .C1(n10168), .C2(n8684), .A(n8683), .B(n8686), .ZN(
        P2_U3490) );
  NAND2_X1 U10204 ( .A1(n10165), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8685) );
  OAI211_X1 U10205 ( .C1(n8748), .C2(n8696), .A(n8686), .B(n8685), .ZN(
        P2_U3489) );
  INV_X1 U10206 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8687) );
  MUX2_X1 U10207 ( .A(n8687), .B(n8749), .S(n10168), .Z(n8689) );
  NAND2_X1 U10208 ( .A1(n8751), .A2(n8733), .ZN(n8688) );
  INV_X1 U10209 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8690) );
  AOI22_X1 U10210 ( .A1(n8757), .A2(n8734), .B1(n8733), .B2(n8756), .ZN(n8691)
         );
  NAND2_X1 U10211 ( .A1(n8692), .A2(n8691), .ZN(P2_U3485) );
  INV_X1 U10212 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8693) );
  MUX2_X1 U10213 ( .A(n8693), .B(n8760), .S(n10168), .Z(n8695) );
  AOI22_X1 U10214 ( .A1(n8763), .A2(n8734), .B1(n8733), .B2(n8762), .ZN(n8694)
         );
  NAND2_X1 U10215 ( .A1(n8695), .A2(n8694), .ZN(P2_U3484) );
  MUX2_X1 U10216 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8766), .S(n10168), .Z(
        n8699) );
  OAI22_X1 U10217 ( .A1(n8772), .A2(n8716), .B1(n8697), .B2(n8696), .ZN(n8698)
         );
  OR2_X1 U10218 ( .A1(n8699), .A2(n8698), .ZN(P2_U3483) );
  MUX2_X1 U10219 ( .A(n10330), .B(n8773), .S(n10168), .Z(n8701) );
  NAND2_X1 U10220 ( .A1(n8775), .A2(n8733), .ZN(n8700) );
  OAI211_X1 U10221 ( .C1(n8778), .C2(n8716), .A(n8701), .B(n8700), .ZN(
        P2_U3482) );
  INV_X1 U10222 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8704) );
  AOI21_X1 U10223 ( .B1(n10144), .B2(n8703), .A(n8702), .ZN(n8779) );
  MUX2_X1 U10224 ( .A(n8704), .B(n8779), .S(n10168), .Z(n8705) );
  OAI21_X1 U10225 ( .B1(n8782), .B2(n8716), .A(n8705), .ZN(P2_U3481) );
  NAND2_X1 U10226 ( .A1(n8706), .A2(n10144), .ZN(n8707) );
  NAND2_X1 U10227 ( .A1(n8708), .A2(n8707), .ZN(n8783) );
  MUX2_X1 U10228 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8783), .S(n10168), .Z(
        n8709) );
  AOI21_X1 U10229 ( .B1(n8734), .B2(n8785), .A(n8709), .ZN(n8710) );
  INV_X1 U10230 ( .A(n8710), .ZN(P2_U3480) );
  NAND2_X1 U10231 ( .A1(n8711), .A2(n10144), .ZN(n8712) );
  NAND2_X1 U10232 ( .A1(n8713), .A2(n8712), .ZN(n8787) );
  MUX2_X1 U10233 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8787), .S(n10168), .Z(
        n8714) );
  INV_X1 U10234 ( .A(n8714), .ZN(n8715) );
  OAI21_X1 U10235 ( .B1(n8791), .B2(n8716), .A(n8715), .ZN(P2_U3479) );
  NAND3_X1 U10236 ( .A1(n8718), .A2(n10153), .A3(n8717), .ZN(n8719) );
  OAI21_X1 U10237 ( .B1(n8720), .B2(n10150), .A(n8719), .ZN(n8721) );
  NOR2_X1 U10238 ( .A1(n8722), .A2(n8721), .ZN(n8792) );
  MUX2_X1 U10239 ( .A(n8723), .B(n8792), .S(n10168), .Z(n8724) );
  INV_X1 U10240 ( .A(n8724), .ZN(P2_U3478) );
  NAND3_X1 U10241 ( .A1(n8647), .A2(n8725), .A3(n10153), .ZN(n8728) );
  NAND2_X1 U10242 ( .A1(n8726), .A2(n10144), .ZN(n8727) );
  AND2_X1 U10243 ( .A1(n8728), .A2(n8727), .ZN(n8729) );
  AND2_X1 U10244 ( .A1(n8730), .A2(n8729), .ZN(n8795) );
  MUX2_X1 U10245 ( .A(n8731), .B(n8795), .S(n10168), .Z(n8732) );
  INV_X1 U10246 ( .A(n8732), .ZN(P2_U3477) );
  MUX2_X1 U10247 ( .A(n4758), .B(n8798), .S(n10168), .Z(n8736) );
  AOI22_X1 U10248 ( .A1(n8803), .A2(n8734), .B1(n8733), .B2(n8800), .ZN(n8735)
         );
  NAND2_X1 U10249 ( .A1(n8736), .A2(n8735), .ZN(P2_U3476) );
  AOI22_X1 U10250 ( .A1(n8738), .A2(n10153), .B1(n10144), .B2(n8737), .ZN(
        n8739) );
  NAND2_X1 U10251 ( .A1(n8740), .A2(n8739), .ZN(n8806) );
  MUX2_X1 U10252 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8806), .S(n10168), .Z(
        P2_U3475) );
  MUX2_X1 U10253 ( .A(n8741), .B(P2_REG1_REG_0__SCAN_IN), .S(n10165), .Z(
        P2_U3459) );
  INV_X1 U10254 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U10255 ( .A1(n8742), .A2(n8801), .ZN(n8744) );
  NAND2_X1 U10256 ( .A1(n8743), .A2(n10155), .ZN(n8746) );
  OAI211_X1 U10257 ( .C1(n10314), .C2(n10155), .A(n8744), .B(n8746), .ZN(
        P2_U3458) );
  NAND2_X1 U10258 ( .A1(n10156), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8745) );
  OAI211_X1 U10259 ( .C1(n8748), .C2(n8747), .A(n8746), .B(n8745), .ZN(
        P2_U3457) );
  MUX2_X1 U10260 ( .A(n8750), .B(n8749), .S(n10155), .Z(n8753) );
  NAND2_X1 U10261 ( .A1(n8751), .A2(n8801), .ZN(n8752) );
  AOI22_X1 U10262 ( .A1(n8757), .A2(n8802), .B1(n8801), .B2(n8756), .ZN(n8758)
         );
  NAND2_X1 U10263 ( .A1(n8759), .A2(n8758), .ZN(P2_U3453) );
  INV_X1 U10264 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n8761) );
  MUX2_X1 U10265 ( .A(n8761), .B(n8760), .S(n10155), .Z(n8765) );
  AOI22_X1 U10266 ( .A1(n8763), .A2(n8802), .B1(n8801), .B2(n8762), .ZN(n8764)
         );
  NAND2_X1 U10267 ( .A1(n8765), .A2(n8764), .ZN(P2_U3452) );
  INV_X1 U10268 ( .A(n8766), .ZN(n8767) );
  MUX2_X1 U10269 ( .A(n8768), .B(n8767), .S(n10155), .Z(n8771) );
  NAND2_X1 U10270 ( .A1(n8769), .A2(n8801), .ZN(n8770) );
  OAI211_X1 U10271 ( .C1(n8772), .C2(n8790), .A(n8771), .B(n8770), .ZN(
        P2_U3451) );
  INV_X1 U10272 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n8774) );
  MUX2_X1 U10273 ( .A(n8774), .B(n8773), .S(n10155), .Z(n8777) );
  NAND2_X1 U10274 ( .A1(n8775), .A2(n8801), .ZN(n8776) );
  OAI211_X1 U10275 ( .C1(n8778), .C2(n8790), .A(n8777), .B(n8776), .ZN(
        P2_U3450) );
  MUX2_X1 U10276 ( .A(n8780), .B(n8779), .S(n10155), .Z(n8781) );
  OAI21_X1 U10277 ( .B1(n8782), .B2(n8790), .A(n8781), .ZN(P2_U3449) );
  MUX2_X1 U10278 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8783), .S(n10155), .Z(
        n8784) );
  AOI21_X1 U10279 ( .B1(n8785), .B2(n8802), .A(n8784), .ZN(n8786) );
  INV_X1 U10280 ( .A(n8786), .ZN(P2_U3448) );
  MUX2_X1 U10281 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8787), .S(n10155), .Z(
        n8788) );
  INV_X1 U10282 ( .A(n8788), .ZN(n8789) );
  OAI21_X1 U10283 ( .B1(n8791), .B2(n8790), .A(n8789), .ZN(P2_U3447) );
  INV_X1 U10284 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8793) );
  MUX2_X1 U10285 ( .A(n8793), .B(n8792), .S(n10155), .Z(n8794) );
  INV_X1 U10286 ( .A(n8794), .ZN(P2_U3446) );
  MUX2_X1 U10287 ( .A(n8796), .B(n8795), .S(n10155), .Z(n8797) );
  INV_X1 U10288 ( .A(n8797), .ZN(P2_U3444) );
  INV_X1 U10289 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8799) );
  MUX2_X1 U10290 ( .A(n8799), .B(n8798), .S(n10155), .Z(n8805) );
  AOI22_X1 U10291 ( .A1(n8803), .A2(n8802), .B1(n8801), .B2(n8800), .ZN(n8804)
         );
  NAND2_X1 U10292 ( .A1(n8805), .A2(n8804), .ZN(P2_U3441) );
  MUX2_X1 U10293 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8806), .S(n10155), .Z(
        P2_U3438) );
  MUX2_X1 U10294 ( .A(n8808), .B(P2_D_REG_1__SCAN_IN), .S(n8807), .Z(P2_U3377)
         );
  INV_X1 U10295 ( .A(n8809), .ZN(n9989) );
  INV_X1 U10296 ( .A(n8810), .ZN(n8812) );
  NOR4_X1 U10297 ( .A1(n8812), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8811), .A4(
        P2_U3151), .ZN(n8813) );
  AOI21_X1 U10298 ( .B1(n8820), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8813), .ZN(
        n8814) );
  OAI21_X1 U10299 ( .B1(n9989), .B2(n8822), .A(n8814), .ZN(P2_U3264) );
  INV_X1 U10300 ( .A(n8815), .ZN(n9998) );
  OAI222_X1 U10301 ( .A1(n8822), .A2(n9998), .B1(P2_U3151), .B2(n8818), .C1(
        n8817), .C2(n8816), .ZN(P2_U3266) );
  AOI21_X1 U10302 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n8820), .A(n8819), .ZN(
        n8821) );
  OAI21_X1 U10303 ( .B1(n8823), .B2(n8822), .A(n8821), .ZN(P2_U3267) );
  MUX2_X1 U10304 ( .A(n8824), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10305 ( .A1(n8830), .A2(n4290), .ZN(n8826) );
  NAND2_X1 U10306 ( .A1(n9465), .A2(n7040), .ZN(n8825) );
  NAND2_X1 U10307 ( .A1(n8826), .A2(n8825), .ZN(n8827) );
  XNOR2_X1 U10308 ( .A(n8827), .B(n9034), .ZN(n8836) );
  NOR2_X1 U10309 ( .A1(n8828), .A2(n8947), .ZN(n8829) );
  AOI21_X1 U10310 ( .B1(n8830), .B2(n7040), .A(n8829), .ZN(n8837) );
  XNOR2_X1 U10311 ( .A(n8836), .B(n8837), .ZN(n9129) );
  NAND2_X1 U10312 ( .A1(n8831), .A2(n8839), .ZN(n8832) );
  NAND2_X1 U10313 ( .A1(n9129), .A2(n8832), .ZN(n9008) );
  AOI22_X1 U10314 ( .A1(n9019), .A2(n7040), .B1(n8952), .B2(n9464), .ZN(n9007)
         );
  NAND2_X1 U10315 ( .A1(n9019), .A2(n4290), .ZN(n8834) );
  NAND2_X1 U10316 ( .A1(n9464), .A2(n7040), .ZN(n8833) );
  NAND2_X1 U10317 ( .A1(n8834), .A2(n8833), .ZN(n8835) );
  XNOR2_X1 U10318 ( .A(n8835), .B(n8964), .ZN(n9011) );
  INV_X1 U10319 ( .A(n8836), .ZN(n8838) );
  AND2_X1 U10320 ( .A1(n8838), .A2(n8837), .ZN(n9010) );
  INV_X1 U10321 ( .A(n8839), .ZN(n8840) );
  NAND2_X1 U10322 ( .A1(n8841), .A2(n8840), .ZN(n9009) );
  NOR2_X1 U10323 ( .A1(n9008), .A2(n9009), .ZN(n8842) );
  AOI22_X1 U10324 ( .A1(n8845), .A2(n4290), .B1(n7040), .B2(n9463), .ZN(n8846)
         );
  XNOR2_X1 U10325 ( .A(n8846), .B(n8964), .ZN(n8848) );
  OAI22_X1 U10326 ( .A1(n5201), .A2(n4294), .B1(n9072), .B2(n8947), .ZN(n8847)
         );
  NOR2_X1 U10327 ( .A1(n8848), .A2(n8847), .ZN(n9067) );
  AOI21_X1 U10328 ( .B1(n8848), .B2(n8847), .A(n9067), .ZN(n9173) );
  INV_X1 U10329 ( .A(n9011), .ZN(n8850) );
  NAND2_X1 U10330 ( .A1(n8856), .A2(n4290), .ZN(n8853) );
  OR2_X1 U10331 ( .A1(n9157), .A2(n4294), .ZN(n8852) );
  NAND2_X1 U10332 ( .A1(n8853), .A2(n8852), .ZN(n8854) );
  XNOR2_X1 U10333 ( .A(n8854), .B(n8964), .ZN(n8858) );
  NOR2_X1 U10334 ( .A1(n9157), .A2(n8947), .ZN(n8855) );
  AOI21_X1 U10335 ( .B1(n8856), .B2(n4480), .A(n8855), .ZN(n8857) );
  NAND2_X1 U10336 ( .A1(n8858), .A2(n8857), .ZN(n8860) );
  OR2_X1 U10337 ( .A1(n8858), .A2(n8857), .ZN(n8859) );
  AND2_X1 U10338 ( .A1(n8860), .A2(n8859), .ZN(n9066) );
  NAND2_X1 U10339 ( .A1(n9939), .A2(n4290), .ZN(n8862) );
  NAND2_X1 U10340 ( .A1(n9075), .A2(n7040), .ZN(n8861) );
  NAND2_X1 U10341 ( .A1(n8862), .A2(n8861), .ZN(n8863) );
  XNOR2_X1 U10342 ( .A(n8863), .B(n8964), .ZN(n8864) );
  OAI22_X1 U10343 ( .A1(n9837), .A2(n4293), .B1(n9809), .B2(n8947), .ZN(n8865)
         );
  XNOR2_X1 U10344 ( .A(n8864), .B(n8865), .ZN(n9154) );
  NAND2_X1 U10345 ( .A1(n8864), .A2(n8866), .ZN(n8867) );
  NAND2_X1 U10346 ( .A1(n5616), .A2(n4290), .ZN(n8869) );
  OR2_X1 U10347 ( .A1(n9211), .A2(n4294), .ZN(n8868) );
  NAND2_X1 U10348 ( .A1(n8869), .A2(n8868), .ZN(n8870) );
  XNOR2_X1 U10349 ( .A(n8870), .B(n8964), .ZN(n8985) );
  NOR2_X1 U10350 ( .A1(n9211), .A2(n8947), .ZN(n8871) );
  AOI21_X1 U10351 ( .B1(n5616), .B2(n4480), .A(n8871), .ZN(n8984) );
  OR2_X1 U10352 ( .A1(n8985), .A2(n8984), .ZN(n8873) );
  AND2_X1 U10353 ( .A1(n8985), .A2(n8984), .ZN(n8872) );
  NAND2_X1 U10354 ( .A1(n9929), .A2(n4290), .ZN(n8875) );
  NAND2_X1 U10355 ( .A1(n9773), .A2(n4480), .ZN(n8874) );
  NAND2_X1 U10356 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  XNOR2_X1 U10357 ( .A(n8876), .B(n9034), .ZN(n8883) );
  NAND2_X1 U10358 ( .A1(n9929), .A2(n4480), .ZN(n8878) );
  NAND2_X1 U10359 ( .A1(n9773), .A2(n8952), .ZN(n8877) );
  NAND2_X1 U10360 ( .A1(n8878), .A2(n8877), .ZN(n9208) );
  OR2_X1 U10361 ( .A1(n8883), .A2(n9208), .ZN(n8879) );
  OAI22_X1 U10362 ( .A1(n9307), .A2(n8922), .B1(n9764), .B2(n4294), .ZN(n8880)
         );
  XNOR2_X1 U10363 ( .A(n8880), .B(n9034), .ZN(n8882) );
  OAI22_X1 U10364 ( .A1(n9307), .A2(n4293), .B1(n9764), .B2(n8947), .ZN(n8881)
         );
  NOR2_X1 U10365 ( .A1(n8882), .A2(n8881), .ZN(n8886) );
  AOI21_X1 U10366 ( .B1(n8882), .B2(n8881), .A(n8886), .ZN(n9092) );
  INV_X1 U10367 ( .A(n8883), .ZN(n9088) );
  NAND2_X1 U10368 ( .A1(n8883), .A2(n9208), .ZN(n8884) );
  NAND2_X1 U10369 ( .A1(n8885), .A2(n5003), .ZN(n9093) );
  INV_X1 U10370 ( .A(n8886), .ZN(n8887) );
  NAND2_X1 U10371 ( .A1(n9919), .A2(n4290), .ZN(n8889) );
  NAND2_X1 U10372 ( .A1(n9772), .A2(n4480), .ZN(n8888) );
  NAND2_X1 U10373 ( .A1(n8889), .A2(n8888), .ZN(n8890) );
  XNOR2_X1 U10374 ( .A(n8890), .B(n8964), .ZN(n8891) );
  OAI22_X1 U10375 ( .A1(n9108), .A2(n4294), .B1(n9742), .B2(n8947), .ZN(n8892)
         );
  XNOR2_X1 U10376 ( .A(n8891), .B(n8892), .ZN(n9101) );
  INV_X1 U10377 ( .A(n8892), .ZN(n8893) );
  NAND2_X1 U10378 ( .A1(n9747), .A2(n4290), .ZN(n8896) );
  NAND2_X1 U10379 ( .A1(n9730), .A2(n4480), .ZN(n8895) );
  NAND2_X1 U10380 ( .A1(n8896), .A2(n8895), .ZN(n8897) );
  XNOR2_X1 U10381 ( .A(n8897), .B(n9034), .ZN(n8901) );
  NAND2_X1 U10382 ( .A1(n9747), .A2(n4480), .ZN(n8899) );
  NAND2_X1 U10383 ( .A1(n9730), .A2(n8952), .ZN(n8898) );
  NAND2_X1 U10384 ( .A1(n8899), .A2(n8898), .ZN(n8900) );
  NAND2_X1 U10385 ( .A1(n8901), .A2(n8900), .ZN(n9183) );
  NAND2_X1 U10386 ( .A1(n9908), .A2(n4290), .ZN(n8904) );
  NAND2_X1 U10387 ( .A1(n9462), .A2(n4480), .ZN(n8903) );
  NAND2_X1 U10388 ( .A1(n8904), .A2(n8903), .ZN(n8905) );
  XNOR2_X1 U10389 ( .A(n8905), .B(n8964), .ZN(n8908) );
  AND2_X1 U10390 ( .A1(n9462), .A2(n8952), .ZN(n8906) );
  AOI21_X1 U10391 ( .B1(n9908), .B2(n4480), .A(n8906), .ZN(n8907) );
  NOR2_X1 U10392 ( .A1(n8908), .A2(n8907), .ZN(n9024) );
  NAND2_X1 U10393 ( .A1(n8908), .A2(n8907), .ZN(n9022) );
  OAI22_X1 U10394 ( .A1(n9717), .A2(n8922), .B1(n9056), .B2(n4293), .ZN(n8909)
         );
  XNOR2_X1 U10395 ( .A(n8909), .B(n9034), .ZN(n8911) );
  OAI22_X1 U10396 ( .A1(n9717), .A2(n4294), .B1(n9056), .B2(n8947), .ZN(n8910)
         );
  NOR2_X1 U10397 ( .A1(n8911), .A2(n8910), .ZN(n8912) );
  AOI21_X1 U10398 ( .B1(n8911), .B2(n8910), .A(n8912), .ZN(n9145) );
  INV_X1 U10399 ( .A(n8912), .ZN(n8913) );
  NAND2_X1 U10400 ( .A1(n9968), .A2(n4290), .ZN(n8915) );
  NAND2_X1 U10401 ( .A1(n9461), .A2(n4480), .ZN(n8914) );
  NAND2_X1 U10402 ( .A1(n8915), .A2(n8914), .ZN(n8916) );
  XNOR2_X1 U10403 ( .A(n8916), .B(n8964), .ZN(n8920) );
  OAI22_X1 U10404 ( .A1(n9697), .A2(n4294), .B1(n8917), .B2(n8947), .ZN(n8918)
         );
  XNOR2_X1 U10405 ( .A(n8920), .B(n8918), .ZN(n9053) );
  INV_X1 U10406 ( .A(n8918), .ZN(n8919) );
  NAND2_X1 U10407 ( .A1(n8920), .A2(n8919), .ZN(n8921) );
  OAI22_X1 U10408 ( .A1(n9965), .A2(n8922), .B1(n9055), .B2(n4293), .ZN(n8923)
         );
  XNOR2_X1 U10409 ( .A(n8923), .B(n9034), .ZN(n8993) );
  OR2_X1 U10410 ( .A1(n9965), .A2(n4294), .ZN(n8925) );
  OR2_X1 U10411 ( .A1(n9055), .A2(n8947), .ZN(n8924) );
  NAND2_X1 U10412 ( .A1(n8925), .A2(n8924), .ZN(n9164) );
  NAND2_X1 U10413 ( .A1(n9667), .A2(n4290), .ZN(n8927) );
  NAND2_X1 U10414 ( .A1(n9459), .A2(n4480), .ZN(n8926) );
  NAND2_X1 U10415 ( .A1(n8927), .A2(n8926), .ZN(n8928) );
  XNOR2_X1 U10416 ( .A(n8928), .B(n8964), .ZN(n8931) );
  AND2_X1 U10417 ( .A1(n9459), .A2(n8952), .ZN(n8929) );
  AOI21_X1 U10418 ( .B1(n9667), .B2(n4480), .A(n8929), .ZN(n8930) );
  NAND2_X1 U10419 ( .A1(n8931), .A2(n8930), .ZN(n9111) );
  OAI21_X1 U10420 ( .B1(n8931), .B2(n8930), .A(n9111), .ZN(n8995) );
  NAND2_X1 U10421 ( .A1(n9652), .A2(n4290), .ZN(n8935) );
  NAND2_X1 U10422 ( .A1(n9458), .A2(n4480), .ZN(n8934) );
  NAND2_X1 U10423 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  XNOR2_X1 U10424 ( .A(n8936), .B(n8964), .ZN(n8938) );
  AND2_X1 U10425 ( .A1(n9458), .A2(n8952), .ZN(n8937) );
  AOI21_X1 U10426 ( .B1(n9652), .B2(n4480), .A(n8937), .ZN(n8939) );
  NAND2_X1 U10427 ( .A1(n8938), .A2(n8939), .ZN(n8943) );
  INV_X1 U10428 ( .A(n8938), .ZN(n8941) );
  INV_X1 U10429 ( .A(n8939), .ZN(n8940) );
  NAND2_X1 U10430 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  NAND2_X1 U10431 ( .A1(n9637), .A2(n4290), .ZN(n8945) );
  NAND2_X1 U10432 ( .A1(n9457), .A2(n4480), .ZN(n8944) );
  NAND2_X1 U10433 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  XNOR2_X1 U10434 ( .A(n8946), .B(n8964), .ZN(n8954) );
  OAI22_X1 U10435 ( .A1(n9955), .A2(n4293), .B1(n9198), .B2(n8947), .ZN(n8955)
         );
  XNOR2_X1 U10436 ( .A(n8954), .B(n8955), .ZN(n9080) );
  NAND2_X1 U10437 ( .A1(n9950), .A2(n4290), .ZN(n8950) );
  NAND2_X1 U10438 ( .A1(n9456), .A2(n4480), .ZN(n8949) );
  NAND2_X1 U10439 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  XNOR2_X1 U10440 ( .A(n8951), .B(n8964), .ZN(n8958) );
  AND2_X1 U10441 ( .A1(n9456), .A2(n8952), .ZN(n8953) );
  AOI21_X1 U10442 ( .B1(n9950), .B2(n4480), .A(n8953), .ZN(n8959) );
  XNOR2_X1 U10443 ( .A(n8958), .B(n8959), .ZN(n9192) );
  INV_X1 U10444 ( .A(n8954), .ZN(n8956) );
  NOR2_X1 U10445 ( .A1(n8956), .A2(n8955), .ZN(n9193) );
  NOR2_X1 U10446 ( .A1(n9192), .A2(n9193), .ZN(n8957) );
  INV_X1 U10447 ( .A(n8958), .ZN(n8961) );
  INV_X1 U10448 ( .A(n8959), .ZN(n8960) );
  NAND2_X1 U10449 ( .A1(n8961), .A2(n8960), .ZN(n8972) );
  NAND2_X1 U10450 ( .A1(n8981), .A2(n4290), .ZN(n8963) );
  NAND2_X1 U10451 ( .A1(n9455), .A2(n4480), .ZN(n8962) );
  NAND2_X1 U10452 ( .A1(n8963), .A2(n8962), .ZN(n8965) );
  XNOR2_X1 U10453 ( .A(n8965), .B(n8964), .ZN(n8968) );
  INV_X1 U10454 ( .A(n8968), .ZN(n8970) );
  NOR2_X1 U10455 ( .A1(n9199), .A2(n8947), .ZN(n8966) );
  AOI21_X1 U10456 ( .B1(n8981), .B2(n4480), .A(n8966), .ZN(n8967) );
  INV_X1 U10457 ( .A(n8967), .ZN(n8969) );
  AOI21_X1 U10458 ( .B1(n8970), .B2(n8969), .A(n9046), .ZN(n8971) );
  AOI21_X1 U10459 ( .B1(n9195), .B2(n8972), .A(n8971), .ZN(n8976) );
  INV_X1 U10460 ( .A(n8971), .ZN(n8974) );
  INV_X1 U10461 ( .A(n8972), .ZN(n8973) );
  NOR2_X1 U10462 ( .A1(n8974), .A2(n8973), .ZN(n8975) );
  OAI21_X1 U10463 ( .B1(n8976), .B2(n9040), .A(n9196), .ZN(n8983) );
  NOR2_X1 U10464 ( .A1(n8977), .A2(n9167), .ZN(n8980) );
  OAI22_X1 U10465 ( .A1(n9609), .A2(n9210), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8978), .ZN(n8979) );
  AOI211_X1 U10466 ( .C1(n8981), .C2(n9215), .A(n8980), .B(n8979), .ZN(n8982)
         );
  NAND2_X1 U10467 ( .A1(n8983), .A2(n8982), .ZN(P1_U3214) );
  XNOR2_X1 U10468 ( .A(n8985), .B(n8984), .ZN(n8986) );
  XNOR2_X1 U10469 ( .A(n8987), .B(n8986), .ZN(n8991) );
  AOI22_X1 U10470 ( .A1(n9015), .A2(n9075), .B1(n9165), .B2(n9819), .ZN(n8988)
         );
  NAND2_X1 U10471 ( .A1(n10066), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10012) );
  OAI211_X1 U10472 ( .C1(n9811), .C2(n9209), .A(n8988), .B(n10012), .ZN(n8989)
         );
  AOI21_X1 U10473 ( .B1(n5616), .B2(n9215), .A(n8989), .ZN(n8990) );
  OAI21_X1 U10474 ( .B1(n8991), .B2(n9217), .A(n8990), .ZN(P1_U3215) );
  INV_X1 U10475 ( .A(n9667), .ZN(n9961) );
  INV_X1 U10476 ( .A(n8993), .ZN(n8994) );
  NAND2_X1 U10477 ( .A1(n8992), .A2(n8994), .ZN(n8996) );
  OAI21_X1 U10478 ( .B1(n8992), .B2(n8994), .A(n8996), .ZN(n9163) );
  NOR2_X1 U10479 ( .A1(n9163), .A2(n9164), .ZN(n9162) );
  INV_X1 U10480 ( .A(n8995), .ZN(n8998) );
  INV_X1 U10481 ( .A(n8996), .ZN(n8997) );
  INV_X1 U10482 ( .A(n9112), .ZN(n9000) );
  OAI21_X1 U10483 ( .B1(n9001), .B2(n9000), .A(n9196), .ZN(n9006) );
  NOR2_X1 U10484 ( .A1(n9669), .A2(n9210), .ZN(n9004) );
  NOR2_X1 U10485 ( .A1(n9055), .A2(n9808), .ZN(n9002) );
  AOI21_X1 U10486 ( .B1(n9458), .B2(n9843), .A(n9002), .ZN(n9661) );
  NOR2_X1 U10487 ( .A1(n9661), .A2(n9167), .ZN(n9003) );
  AOI211_X1 U10488 ( .C1(P1_REG3_REG_23__SCAN_IN), .C2(P1_U3086), .A(n9004), 
        .B(n9003), .ZN(n9005) );
  AOI21_X1 U10489 ( .B1(n8844), .B2(n9009), .A(n9008), .ZN(n9132) );
  OR2_X1 U10490 ( .A1(n9132), .A2(n9010), .ZN(n9012) );
  NAND2_X1 U10491 ( .A1(n9012), .A2(n9011), .ZN(n9171) );
  OAI21_X1 U10492 ( .B1(n9012), .B2(n9011), .A(n9171), .ZN(n9013) );
  NOR2_X1 U10493 ( .A1(n9013), .A2(n8849), .ZN(n9174) );
  AOI21_X1 U10494 ( .B1(n8849), .B2(n9013), .A(n9174), .ZN(n9021) );
  AOI22_X1 U10495 ( .A1(n9015), .A2(n9465), .B1(n9165), .B2(n9014), .ZN(n9017)
         );
  OAI211_X1 U10496 ( .C1(n9072), .C2(n9209), .A(n9017), .B(n9016), .ZN(n9018)
         );
  AOI21_X1 U10497 ( .B1(n9019), .B2(n9215), .A(n9018), .ZN(n9020) );
  OAI21_X1 U10498 ( .B1(n9021), .B2(n9217), .A(n9020), .ZN(P1_U3217) );
  INV_X1 U10499 ( .A(n9022), .ZN(n9023) );
  NOR2_X1 U10500 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  XNOR2_X1 U10501 ( .A(n9026), .B(n9025), .ZN(n9030) );
  OAI22_X1 U10502 ( .A1(n9056), .A2(n9209), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10261), .ZN(n9028) );
  OAI22_X1 U10503 ( .A1(n9212), .A2(n9763), .B1(n9210), .B2(n9724), .ZN(n9027)
         );
  AOI211_X1 U10504 ( .C1(n9908), .C2(n9215), .A(n9028), .B(n9027), .ZN(n9029)
         );
  OAI21_X1 U10505 ( .B1(n9030), .B2(n9217), .A(n9029), .ZN(P1_U3219) );
  INV_X1 U10506 ( .A(n9046), .ZN(n9039) );
  NAND2_X1 U10507 ( .A1(n9045), .A2(n4480), .ZN(n9033) );
  OR2_X1 U10508 ( .A1(n9031), .A2(n8947), .ZN(n9032) );
  NAND2_X1 U10509 ( .A1(n9033), .A2(n9032), .ZN(n9035) );
  XNOR2_X1 U10510 ( .A(n9035), .B(n9034), .ZN(n9037) );
  AOI22_X1 U10511 ( .A1(n9045), .A2(n4290), .B1(n4480), .B2(n9454), .ZN(n9036)
         );
  XNOR2_X1 U10512 ( .A(n9037), .B(n9036), .ZN(n9047) );
  INV_X1 U10513 ( .A(n9047), .ZN(n9038) );
  NAND3_X1 U10514 ( .A1(n9040), .A2(n9196), .A3(n9047), .ZN(n9050) );
  AOI22_X1 U10515 ( .A1(n9041), .A2(n9165), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        n10066), .ZN(n9042) );
  OAI21_X1 U10516 ( .B1(n9043), .B2(n9167), .A(n9042), .ZN(n9044) );
  AOI21_X1 U10517 ( .B1(n9045), .B2(n9215), .A(n9044), .ZN(n9049) );
  NAND3_X1 U10518 ( .A1(n9047), .A2(n9046), .A3(n9196), .ZN(n9048) );
  OAI21_X1 U10519 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9054) );
  NAND2_X1 U10520 ( .A1(n9054), .A2(n9196), .ZN(n9063) );
  INV_X1 U10521 ( .A(n9694), .ZN(n9061) );
  OR2_X1 U10522 ( .A1(n9055), .A2(n9810), .ZN(n9058) );
  OR2_X1 U10523 ( .A1(n9056), .A2(n9808), .ZN(n9057) );
  NAND2_X1 U10524 ( .A1(n9058), .A2(n9057), .ZN(n9705) );
  INV_X1 U10525 ( .A(n9705), .ZN(n9059) );
  OAI22_X1 U10526 ( .A1(n9059), .A2(n9167), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10233), .ZN(n9060) );
  AOI21_X1 U10527 ( .B1(n9061), .B2(n9165), .A(n9060), .ZN(n9062) );
  OAI211_X1 U10528 ( .C1(n9697), .C2(n9205), .A(n9063), .B(n9062), .ZN(
        P1_U3223) );
  INV_X1 U10529 ( .A(n9064), .ZN(n9069) );
  NOR3_X1 U10530 ( .A1(n9175), .A2(n9067), .A3(n9066), .ZN(n9068) );
  OAI21_X1 U10531 ( .B1(n9069), .B2(n9068), .A(n9196), .ZN(n9077) );
  INV_X1 U10532 ( .A(n9070), .ZN(n9071) );
  OAI22_X1 U10533 ( .A1(n9212), .A2(n9072), .B1(n9210), .B2(n9071), .ZN(n9073)
         );
  AOI211_X1 U10534 ( .C1(n9180), .C2(n9075), .A(n9074), .B(n9073), .ZN(n9076)
         );
  OAI211_X1 U10535 ( .C1(n4793), .C2(n9205), .A(n9077), .B(n9076), .ZN(
        P1_U3224) );
  OAI21_X1 U10536 ( .B1(n9080), .B2(n9079), .A(n9078), .ZN(n9081) );
  NAND2_X1 U10537 ( .A1(n9081), .A2(n9196), .ZN(n9086) );
  AOI22_X1 U10538 ( .A1(n9456), .A2(n9843), .B1(n9841), .B2(n9458), .ZN(n9632)
         );
  INV_X1 U10539 ( .A(n9632), .ZN(n9084) );
  OAI22_X1 U10540 ( .A1(n9639), .A2(n9210), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9082), .ZN(n9083) );
  AOI21_X1 U10541 ( .B1(n9084), .B2(n9202), .A(n9083), .ZN(n9085) );
  OAI211_X1 U10542 ( .C1(n9955), .C2(n9205), .A(n9086), .B(n9085), .ZN(
        P1_U3225) );
  INV_X1 U10543 ( .A(n9087), .ZN(n9089) );
  NAND2_X1 U10544 ( .A1(n9089), .A2(n9088), .ZN(n9090) );
  OAI21_X1 U10545 ( .B1(n9089), .B2(n9088), .A(n9090), .ZN(n9207) );
  NOR2_X1 U10546 ( .A1(n9207), .A2(n9208), .ZN(n9206) );
  INV_X1 U10547 ( .A(n9090), .ZN(n9091) );
  NOR3_X1 U10548 ( .A1(n9206), .A2(n9092), .A3(n9091), .ZN(n9095) );
  INV_X1 U10549 ( .A(n9093), .ZN(n9094) );
  OAI21_X1 U10550 ( .B1(n9095), .B2(n9094), .A(n9196), .ZN(n9098) );
  AND2_X1 U10551 ( .A1(n10066), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10032) );
  OAI22_X1 U10552 ( .A1(n9212), .A2(n9811), .B1(n9210), .B2(n9780), .ZN(n9096)
         );
  AOI211_X1 U10553 ( .C1(n9180), .C2(n9772), .A(n10032), .B(n9096), .ZN(n9097)
         );
  OAI211_X1 U10554 ( .C1(n9307), .C2(n9205), .A(n9098), .B(n9097), .ZN(
        P1_U3226) );
  OAI21_X1 U10555 ( .B1(n9101), .B2(n9100), .A(n4479), .ZN(n9102) );
  NAND2_X1 U10556 ( .A1(n9102), .A2(n9196), .ZN(n9107) );
  NAND2_X1 U10557 ( .A1(n10066), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10050) );
  INV_X1 U10558 ( .A(n10050), .ZN(n9105) );
  INV_X1 U10559 ( .A(n9103), .ZN(n9755) );
  OAI22_X1 U10560 ( .A1(n9212), .A2(n9764), .B1(n9210), .B2(n9755), .ZN(n9104)
         );
  AOI211_X1 U10561 ( .C1(n9180), .C2(n9730), .A(n9105), .B(n9104), .ZN(n9106)
         );
  OAI211_X1 U10562 ( .C1(n9108), .C2(n9205), .A(n9107), .B(n9106), .ZN(
        P1_U3228) );
  AOI22_X1 U10563 ( .A1(n9457), .A2(n9843), .B1(n9841), .B2(n9459), .ZN(n9649)
         );
  AOI22_X1 U10564 ( .A1(n9653), .A2(n9165), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9109) );
  OAI21_X1 U10565 ( .B1(n9649), .B2(n9167), .A(n9109), .ZN(n9116) );
  NAND3_X1 U10566 ( .A1(n9112), .A2(n9111), .A3(n4818), .ZN(n9113) );
  AOI21_X1 U10567 ( .B1(n9114), .B2(n9113), .A(n9217), .ZN(n9115) );
  OAI211_X1 U10568 ( .C1(n9119), .C2(n9118), .A(n9117), .B(n9196), .ZN(n9127)
         );
  AOI21_X1 U10569 ( .B1(n9202), .B2(n9121), .A(n9120), .ZN(n9126) );
  NAND2_X1 U10570 ( .A1(n9165), .A2(n9122), .ZN(n9125) );
  NAND2_X1 U10571 ( .A1(n9215), .A2(n9123), .ZN(n9124) );
  NAND4_X1 U10572 ( .A1(n9127), .A2(n9126), .A3(n9125), .A4(n9124), .ZN(
        P1_U3230) );
  INV_X1 U10573 ( .A(n9128), .ZN(n9130) );
  NOR3_X1 U10574 ( .A1(n9131), .A2(n9130), .A3(n9129), .ZN(n9133) );
  OAI21_X1 U10575 ( .B1(n9133), .B2(n9132), .A(n9196), .ZN(n9141) );
  INV_X1 U10576 ( .A(n9134), .ZN(n9139) );
  INV_X1 U10577 ( .A(n9135), .ZN(n9136) );
  OAI22_X1 U10578 ( .A1(n9212), .A2(n9137), .B1(n9210), .B2(n9136), .ZN(n9138)
         );
  AOI211_X1 U10579 ( .C1(n9180), .C2(n9464), .A(n9139), .B(n9138), .ZN(n9140)
         );
  OAI211_X1 U10580 ( .C1(n9142), .C2(n9205), .A(n9141), .B(n9140), .ZN(
        P1_U3231) );
  OAI21_X1 U10581 ( .B1(n9145), .B2(n9144), .A(n9143), .ZN(n9146) );
  NAND2_X1 U10582 ( .A1(n9146), .A2(n9196), .ZN(n9151) );
  AND2_X1 U10583 ( .A1(n9462), .A2(n9841), .ZN(n9147) );
  AOI21_X1 U10584 ( .B1(n9461), .B2(n9843), .A(n9147), .ZN(n9710) );
  OAI22_X1 U10585 ( .A1(n9710), .A2(n9167), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9148), .ZN(n9149) );
  AOI21_X1 U10586 ( .B1(n9715), .B2(n9165), .A(n9149), .ZN(n9150) );
  OAI211_X1 U10587 ( .C1(n9717), .C2(n9205), .A(n9151), .B(n9150), .ZN(
        P1_U3233) );
  OAI21_X1 U10588 ( .B1(n9154), .B2(n9153), .A(n9152), .ZN(n9155) );
  NAND2_X1 U10589 ( .A1(n9155), .A2(n9196), .ZN(n9161) );
  INV_X1 U10590 ( .A(n9834), .ZN(n9156) );
  OAI22_X1 U10591 ( .A1(n9212), .A2(n9157), .B1(n9210), .B2(n9156), .ZN(n9158)
         );
  AOI211_X1 U10592 ( .C1(n9180), .C2(n9844), .A(n9159), .B(n9158), .ZN(n9160)
         );
  OAI211_X1 U10593 ( .C1(n9837), .C2(n9205), .A(n9161), .B(n9160), .ZN(
        P1_U3234) );
  AOI21_X1 U10594 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9170) );
  AOI22_X1 U10595 ( .A1(n9459), .A2(n9843), .B1(n9841), .B2(n9461), .ZN(n9681)
         );
  AOI22_X1 U10596 ( .A1(n9685), .A2(n9165), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9166) );
  OAI21_X1 U10597 ( .B1(n9681), .B2(n9167), .A(n9166), .ZN(n9168) );
  AOI21_X1 U10598 ( .B1(n9683), .B2(n9215), .A(n9168), .ZN(n9169) );
  OAI21_X1 U10599 ( .B1(n9170), .B2(n9217), .A(n9169), .ZN(P1_U3235) );
  INV_X1 U10600 ( .A(n9171), .ZN(n9172) );
  NOR3_X1 U10601 ( .A1(n9174), .A2(n9173), .A3(n9172), .ZN(n9176) );
  OAI21_X1 U10602 ( .B1(n9176), .B2(n9175), .A(n9196), .ZN(n9182) );
  AND2_X1 U10603 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9558) );
  OAI22_X1 U10604 ( .A1(n9212), .A2(n9178), .B1(n9210), .B2(n9177), .ZN(n9179)
         );
  AOI211_X1 U10605 ( .C1(n9180), .C2(n9842), .A(n9558), .B(n9179), .ZN(n9181)
         );
  OAI211_X1 U10606 ( .C1(n5201), .C2(n9205), .A(n9182), .B(n9181), .ZN(
        P1_U3236) );
  NAND2_X1 U10607 ( .A1(n4402), .A2(n9183), .ZN(n9184) );
  XNOR2_X1 U10608 ( .A(n9185), .B(n9184), .ZN(n9191) );
  OAI22_X1 U10609 ( .A1(n9209), .A2(n9743), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9186), .ZN(n9189) );
  INV_X1 U10610 ( .A(n9748), .ZN(n9187) );
  OAI22_X1 U10611 ( .A1(n9212), .A2(n9742), .B1(n9210), .B2(n9187), .ZN(n9188)
         );
  AOI211_X1 U10612 ( .C1(n9747), .C2(n9215), .A(n9189), .B(n9188), .ZN(n9190)
         );
  OAI21_X1 U10613 ( .B1(n9191), .B2(n9217), .A(n9190), .ZN(P1_U3238) );
  INV_X1 U10614 ( .A(n9078), .ZN(n9194) );
  OAI21_X1 U10615 ( .B1(n9194), .B2(n9193), .A(n9192), .ZN(n9197) );
  NAND3_X1 U10616 ( .A1(n9197), .A2(n9196), .A3(n9195), .ZN(n9204) );
  OAI22_X1 U10617 ( .A1(n9199), .A2(n9810), .B1(n9198), .B2(n9808), .ZN(n9617)
         );
  OAI22_X1 U10618 ( .A1(n9622), .A2(n9210), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9200), .ZN(n9201) );
  AOI21_X1 U10619 ( .B1(n9617), .B2(n9202), .A(n9201), .ZN(n9203) );
  OAI211_X1 U10620 ( .C1(n9625), .C2(n9205), .A(n9204), .B(n9203), .ZN(
        P1_U3240) );
  AOI21_X1 U10621 ( .B1(n9208), .B2(n9207), .A(n9206), .ZN(n9218) );
  NAND2_X1 U10622 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10025)
         );
  OAI21_X1 U10623 ( .B1(n9209), .B2(n9764), .A(n10025), .ZN(n9214) );
  OAI22_X1 U10624 ( .A1(n9212), .A2(n9211), .B1(n9210), .B2(n9790), .ZN(n9213)
         );
  AOI211_X1 U10625 ( .C1(n9929), .C2(n9215), .A(n9214), .B(n9213), .ZN(n9216)
         );
  OAI21_X1 U10626 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(P1_U3241) );
  NAND2_X1 U10627 ( .A1(n9358), .A2(n4363), .ZN(n9363) );
  INV_X1 U10628 ( .A(n9230), .ZN(n9437) );
  OAI211_X1 U10629 ( .C1(n5776), .C2(n9348), .A(n9351), .B(n4322), .ZN(n9221)
         );
  NAND2_X1 U10630 ( .A1(n9221), .A2(n9352), .ZN(n9222) );
  AND2_X1 U10631 ( .A1(n9222), .A2(n9362), .ZN(n9228) );
  INV_X1 U10632 ( .A(n9228), .ZN(n9434) );
  NOR2_X1 U10633 ( .A1(n9223), .A2(n9434), .ZN(n9232) );
  NAND2_X1 U10634 ( .A1(n9349), .A2(n9257), .ZN(n9347) );
  INV_X1 U10635 ( .A(n9347), .ZN(n9225) );
  NAND3_X1 U10636 ( .A1(n9352), .A2(n9225), .A3(n9224), .ZN(n9227) );
  NAND2_X1 U10637 ( .A1(n9361), .A2(n9226), .ZN(n9360) );
  AOI21_X1 U10638 ( .B1(n9228), .B2(n9227), .A(n9360), .ZN(n9231) );
  NAND2_X1 U10639 ( .A1(n9359), .A2(n9357), .ZN(n9367) );
  INV_X1 U10640 ( .A(n9377), .ZN(n9229) );
  INV_X1 U10641 ( .A(n9234), .ZN(n9233) );
  INV_X1 U10642 ( .A(n9376), .ZN(n9385) );
  NAND2_X1 U10643 ( .A1(n9233), .A2(n4996), .ZN(n9236) );
  AOI21_X1 U10644 ( .B1(n9236), .B2(n4804), .A(n9235), .ZN(n9238) );
  NAND2_X1 U10645 ( .A1(n9391), .A2(n9385), .ZN(n9393) );
  OAI211_X1 U10646 ( .C1(n9238), .C2(n9438), .A(n9237), .B(n9393), .ZN(n9266)
         );
  INV_X1 U10647 ( .A(n9241), .ZN(n9252) );
  NOR2_X1 U10648 ( .A1(n9243), .A2(n9242), .ZN(n9247) );
  NOR2_X1 U10649 ( .A1(n10087), .A2(n4299), .ZN(n9245) );
  NOR2_X1 U10650 ( .A1(n6950), .A2(n7251), .ZN(n9244) );
  NAND4_X1 U10651 ( .A1(n9247), .A2(n9246), .A3(n9245), .A4(n9244), .ZN(n9248)
         );
  NOR3_X1 U10652 ( .A1(n9250), .A2(n9249), .A3(n9248), .ZN(n9251) );
  NAND4_X1 U10653 ( .A1(n5773), .A2(n9252), .A3(n9412), .A4(n9251), .ZN(n9253)
         );
  NOR2_X1 U10654 ( .A1(n9827), .A2(n9253), .ZN(n9254) );
  NAND4_X1 U10655 ( .A1(n9796), .A2(n9807), .A3(n9760), .A4(n9254), .ZN(n9255)
         );
  NOR2_X1 U10656 ( .A1(n9740), .A2(n9255), .ZN(n9256) );
  NAND4_X1 U10657 ( .A1(n9713), .A2(n9778), .A3(n9729), .A4(n9256), .ZN(n9258)
         );
  AND4_X1 U10658 ( .A1(n9259), .A2(n9635), .A3(n4992), .A4(n9664), .ZN(n9261)
         );
  INV_X1 U10659 ( .A(n9620), .ZN(n9260) );
  NAND3_X1 U10660 ( .A1(n9262), .A2(n9261), .A3(n9260), .ZN(n9263) );
  OR3_X1 U10661 ( .A1(n4327), .A2(n9370), .A3(n9263), .ZN(n9265) );
  NOR2_X1 U10662 ( .A1(n9602), .A2(n9383), .ZN(n9381) );
  INV_X1 U10663 ( .A(n9381), .ZN(n9264) );
  NAND2_X1 U10664 ( .A1(n9393), .A2(n9264), .ZN(n9440) );
  NAND2_X1 U10665 ( .A1(n4335), .A2(n9395), .ZN(n9269) );
  AOI21_X1 U10666 ( .B1(n9384), .B2(n4300), .A(n9267), .ZN(n9268) );
  INV_X1 U10667 ( .A(n9327), .ZN(n9311) );
  AND2_X1 U10668 ( .A1(n9764), .A2(n9384), .ZN(n9270) );
  AOI22_X1 U10669 ( .A1(n9929), .A2(n9270), .B1(n9382), .B2(n9797), .ZN(n9272)
         );
  INV_X1 U10670 ( .A(n9270), .ZN(n9271) );
  OAI22_X1 U10671 ( .A1(n9311), .A2(n9272), .B1(n9773), .B2(n9271), .ZN(n9314)
         );
  AND2_X1 U10672 ( .A1(n9403), .A2(n9402), .ZN(n9274) );
  NAND2_X1 U10673 ( .A1(n9286), .A2(n9280), .ZN(n9273) );
  AOI21_X1 U10674 ( .B1(n9275), .B2(n9274), .A(n9273), .ZN(n9399) );
  NAND4_X1 U10675 ( .A1(n9288), .A2(n9382), .A3(n9276), .A4(n9406), .ZN(n9291)
         );
  NAND2_X1 U10676 ( .A1(n9284), .A2(n9382), .ZN(n9277) );
  OAI211_X1 U10677 ( .C1(n9278), .C2(n9382), .A(n9288), .B(n9277), .ZN(n9290)
         );
  NAND3_X1 U10678 ( .A1(n9283), .A2(n9406), .A3(n9403), .ZN(n9289) );
  INV_X1 U10679 ( .A(n9284), .ZN(n9285) );
  NOR2_X1 U10680 ( .A1(n9285), .A2(n9382), .ZN(n9287) );
  MUX2_X1 U10681 ( .A(n9293), .B(n9292), .S(n9384), .Z(n9300) );
  INV_X1 U10682 ( .A(n9294), .ZN(n9295) );
  NOR2_X1 U10683 ( .A1(n9296), .A2(n9295), .ZN(n9297) );
  MUX2_X1 U10684 ( .A(n9298), .B(n9297), .S(n9384), .Z(n9299) );
  NAND2_X1 U10685 ( .A1(n9319), .A2(n9303), .ZN(n9414) );
  INV_X1 U10686 ( .A(n9929), .ZN(n9793) );
  NOR2_X1 U10687 ( .A1(n9764), .A2(n9811), .ZN(n9305) );
  AOI211_X1 U10688 ( .C1(n9793), .C2(n9305), .A(n9382), .B(n9307), .ZN(n9313)
         );
  NAND3_X1 U10689 ( .A1(n9306), .A2(n9764), .A3(n9304), .ZN(n9308) );
  AOI211_X1 U10690 ( .C1(n9764), .C2(n9311), .A(n9384), .B(n9310), .ZN(n9312)
         );
  AOI21_X1 U10691 ( .B1(n9317), .B2(n9316), .A(n9315), .ZN(n9321) );
  NAND2_X1 U10692 ( .A1(n9318), .A2(n9409), .ZN(n9320) );
  OAI211_X1 U10693 ( .C1(n9321), .C2(n9320), .A(n9416), .B(n9319), .ZN(n9323)
         );
  NAND2_X1 U10694 ( .A1(n9323), .A2(n9322), .ZN(n9325) );
  INV_X1 U10695 ( .A(n9419), .ZN(n9324) );
  AOI211_X1 U10696 ( .C1(n9325), .C2(n9417), .A(n9324), .B(n9804), .ZN(n9329)
         );
  INV_X1 U10697 ( .A(n9758), .ZN(n9328) );
  NAND2_X1 U10698 ( .A1(n9327), .A2(n9326), .ZN(n9422) );
  NAND2_X1 U10699 ( .A1(n9333), .A2(n9332), .ZN(n9336) );
  INV_X1 U10700 ( .A(n9334), .ZN(n9335) );
  AND2_X1 U10701 ( .A1(n9338), .A2(n9337), .ZN(n9425) );
  NAND2_X1 U10702 ( .A1(n9340), .A2(n9339), .ZN(n9429) );
  AOI21_X1 U10703 ( .B1(n9341), .B2(n9425), .A(n9429), .ZN(n9343) );
  NAND2_X1 U10704 ( .A1(n9700), .A2(n9428), .ZN(n9342) );
  MUX2_X1 U10705 ( .A(n9345), .B(n9344), .S(n9384), .Z(n9346) );
  AOI21_X1 U10706 ( .B1(n4322), .B2(n9348), .A(n9382), .ZN(n9350) );
  INV_X1 U10707 ( .A(n9351), .ZN(n9354) );
  INV_X1 U10708 ( .A(n9352), .ZN(n9353) );
  MUX2_X1 U10709 ( .A(n9354), .B(n9353), .S(n9384), .Z(n9355) );
  NOR2_X1 U10710 ( .A1(n4955), .A2(n9362), .ZN(n9364) );
  OAI21_X1 U10711 ( .B1(n9368), .B2(n9367), .A(n9366), .ZN(n9369) );
  INV_X1 U10712 ( .A(n9378), .ZN(n9373) );
  NAND2_X1 U10713 ( .A1(n9377), .A2(n9384), .ZN(n9372) );
  OAI22_X1 U10714 ( .A1(n9384), .A2(n9373), .B1(n9372), .B2(n9602), .ZN(n9375)
         );
  NOR2_X1 U10715 ( .A1(n4804), .A2(n9384), .ZN(n9374) );
  OAI21_X1 U10716 ( .B1(n9377), .B2(n9382), .A(n9376), .ZN(n9380) );
  NOR2_X1 U10717 ( .A1(n9378), .A2(n9384), .ZN(n9379) );
  NOR4_X1 U10718 ( .A1(n4327), .A2(n9381), .A3(n9380), .A4(n9379), .ZN(n9389)
         );
  NOR3_X1 U10719 ( .A1(n9383), .A2(n9385), .A3(n9382), .ZN(n9387) );
  INV_X1 U10720 ( .A(n9383), .ZN(n9453) );
  NOR3_X1 U10721 ( .A1(n9453), .A2(n9385), .A3(n9384), .ZN(n9386) );
  MUX2_X1 U10722 ( .A(n9387), .B(n9386), .S(n9602), .Z(n9388) );
  NAND3_X1 U10723 ( .A1(n9398), .A2(n9395), .A3(n4299), .ZN(n9447) );
  NOR2_X1 U10724 ( .A1(n9393), .A2(n9765), .ZN(n9397) );
  AOI211_X1 U10725 ( .C1(n9438), .C2(n9395), .A(n4301), .B(n9394), .ZN(n9396)
         );
  OAI21_X1 U10726 ( .B1(n9398), .B2(n9397), .A(n9396), .ZN(n9445) );
  INV_X1 U10727 ( .A(n9399), .ZN(n9408) );
  AND4_X1 U10728 ( .A1(n9402), .A2(n9401), .A3(n9400), .A4(n4299), .ZN(n9405)
         );
  AND3_X1 U10729 ( .A1(n9405), .A2(n9404), .A3(n9403), .ZN(n9407) );
  OAI21_X1 U10730 ( .B1(n9408), .B2(n9407), .A(n9406), .ZN(n9413) );
  NAND2_X1 U10731 ( .A1(n9410), .A2(n9409), .ZN(n9411) );
  AOI21_X1 U10732 ( .B1(n9413), .B2(n9412), .A(n9411), .ZN(n9415) );
  OAI21_X1 U10733 ( .B1(n9415), .B2(n9414), .A(n4401), .ZN(n9418) );
  NAND3_X1 U10734 ( .A1(n9418), .A2(n9417), .A3(n9416), .ZN(n9420) );
  AND3_X1 U10735 ( .A1(n9420), .A2(n9304), .A3(n9419), .ZN(n9423) );
  OAI211_X1 U10736 ( .C1(n9423), .C2(n9422), .A(n9421), .B(n9306), .ZN(n9424)
         );
  NAND2_X1 U10737 ( .A1(n9424), .A2(n9758), .ZN(n9427) );
  INV_X1 U10738 ( .A(n9425), .ZN(n9426) );
  AOI21_X1 U10739 ( .B1(n9427), .B2(n4400), .A(n9426), .ZN(n9430) );
  OAI21_X1 U10740 ( .B1(n9430), .B2(n9429), .A(n9428), .ZN(n9431) );
  NAND2_X1 U10741 ( .A1(n9432), .A2(n9431), .ZN(n9433) );
  NOR2_X1 U10742 ( .A1(n9434), .A2(n9433), .ZN(n9436) );
  AOI21_X1 U10743 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9441) );
  INV_X1 U10744 ( .A(n9438), .ZN(n9439) );
  OAI21_X1 U10745 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9442) );
  MUX2_X1 U10746 ( .A(n10088), .B(n9443), .S(n9442), .Z(n9444) );
  NAND2_X1 U10747 ( .A1(n9445), .A2(n9444), .ZN(n9446) );
  NOR3_X1 U10748 ( .A1(n9449), .A2(n10086), .A3(n9448), .ZN(n9451) );
  OAI21_X1 U10749 ( .B1(n9452), .B2(n4301), .A(P1_B_REG_SCAN_IN), .ZN(n9450)
         );
  MUX2_X1 U10750 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9453), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10751 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9454), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10752 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9455), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10753 ( .A(n9456), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9473), .Z(
        P1_U3580) );
  MUX2_X1 U10754 ( .A(n9457), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9473), .Z(
        P1_U3579) );
  MUX2_X1 U10755 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9458), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10756 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9459), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10757 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9460), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10758 ( .A(n9461), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9473), .Z(
        P1_U3575) );
  MUX2_X1 U10759 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9731), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10760 ( .A(n9462), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9473), .Z(
        P1_U3573) );
  MUX2_X1 U10761 ( .A(n9730), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9473), .Z(
        P1_U3572) );
  MUX2_X1 U10762 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9772), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10763 ( .A(n9797), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9473), .Z(
        P1_U3570) );
  MUX2_X1 U10764 ( .A(n9773), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9473), .Z(
        P1_U3569) );
  MUX2_X1 U10765 ( .A(n9844), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9473), .Z(
        P1_U3568) );
  MUX2_X1 U10766 ( .A(n9842), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9473), .Z(
        P1_U3566) );
  MUX2_X1 U10767 ( .A(n9463), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9473), .Z(
        P1_U3565) );
  MUX2_X1 U10768 ( .A(n9464), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9473), .Z(
        P1_U3564) );
  MUX2_X1 U10769 ( .A(n9465), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9473), .Z(
        P1_U3563) );
  MUX2_X1 U10770 ( .A(n9466), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9473), .Z(
        P1_U3562) );
  MUX2_X1 U10771 ( .A(n9467), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9473), .Z(
        P1_U3561) );
  MUX2_X1 U10772 ( .A(n9468), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9473), .Z(
        P1_U3560) );
  MUX2_X1 U10773 ( .A(n9469), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9473), .Z(
        P1_U3559) );
  MUX2_X1 U10774 ( .A(n9470), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9473), .Z(
        P1_U3558) );
  MUX2_X1 U10775 ( .A(n9471), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9473), .Z(
        P1_U3557) );
  MUX2_X1 U10776 ( .A(n9472), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9473), .Z(
        P1_U3556) );
  MUX2_X1 U10777 ( .A(n6715), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9473), .Z(
        P1_U3555) );
  MUX2_X1 U10778 ( .A(n9474), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9473), .Z(
        P1_U3554) );
  OAI211_X1 U10779 ( .C1(n9477), .C2(n9476), .A(n10048), .B(n9475), .ZN(n9484)
         );
  OAI211_X1 U10780 ( .C1(n9480), .C2(n9479), .A(n10047), .B(n9478), .ZN(n9483)
         );
  AOI22_X1 U10781 ( .A1(n10033), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10066), .ZN(n9482) );
  NAND2_X1 U10782 ( .A1(n4409), .A2(n5061), .ZN(n9481) );
  NAND4_X1 U10783 ( .A1(n9484), .A2(n9483), .A3(n9482), .A4(n9481), .ZN(
        P1_U3244) );
  INV_X1 U10784 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9486) );
  OAI21_X1 U10785 ( .B1(n10070), .B2(n9486), .A(n9485), .ZN(n9487) );
  AOI21_X1 U10786 ( .B1(n9488), .B2(n4409), .A(n9487), .ZN(n9497) );
  OAI211_X1 U10787 ( .C1(n9491), .C2(n9490), .A(n10047), .B(n9489), .ZN(n9496)
         );
  OAI211_X1 U10788 ( .C1(n9494), .C2(n9493), .A(n10048), .B(n9492), .ZN(n9495)
         );
  NAND3_X1 U10789 ( .A1(n9497), .A2(n9496), .A3(n9495), .ZN(P1_U3246) );
  INV_X1 U10790 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9499) );
  NAND2_X1 U10791 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9498) );
  OAI21_X1 U10792 ( .B1(n10070), .B2(n9499), .A(n9498), .ZN(n9500) );
  AOI21_X1 U10793 ( .B1(n9501), .B2(n4409), .A(n9500), .ZN(n9510) );
  OAI211_X1 U10794 ( .C1(n9504), .C2(n9503), .A(n10047), .B(n9502), .ZN(n9509)
         );
  OAI211_X1 U10795 ( .C1(n9507), .C2(n9506), .A(n10048), .B(n9505), .ZN(n9508)
         );
  NAND3_X1 U10796 ( .A1(n9510), .A2(n9509), .A3(n9508), .ZN(P1_U3248) );
  INV_X1 U10797 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9512) );
  OAI21_X1 U10798 ( .B1(n10070), .B2(n9512), .A(n9511), .ZN(n9513) );
  AOI21_X1 U10799 ( .B1(n9514), .B2(n4409), .A(n9513), .ZN(n9523) );
  OAI211_X1 U10800 ( .C1(n9517), .C2(n9516), .A(n10048), .B(n9515), .ZN(n9522)
         );
  OAI211_X1 U10801 ( .C1(n9520), .C2(n9519), .A(n10047), .B(n9518), .ZN(n9521)
         );
  NAND3_X1 U10802 ( .A1(n9523), .A2(n9522), .A3(n9521), .ZN(P1_U3249) );
  INV_X1 U10803 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U10804 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(n10066), .ZN(n9524) );
  OAI21_X1 U10805 ( .B1(n10070), .B2(n9525), .A(n9524), .ZN(n9526) );
  AOI21_X1 U10806 ( .B1(n9527), .B2(n4409), .A(n9526), .ZN(n9536) );
  OAI211_X1 U10807 ( .C1(n9530), .C2(n9529), .A(n10048), .B(n9528), .ZN(n9535)
         );
  OAI211_X1 U10808 ( .C1(n9533), .C2(n9532), .A(n10047), .B(n9531), .ZN(n9534)
         );
  NAND3_X1 U10809 ( .A1(n9536), .A2(n9535), .A3(n9534), .ZN(P1_U3250) );
  INV_X1 U10810 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9538) );
  OAI21_X1 U10811 ( .B1(n10070), .B2(n9538), .A(n9537), .ZN(n9539) );
  AOI21_X1 U10812 ( .B1(n9540), .B2(n4409), .A(n9539), .ZN(n9549) );
  OAI211_X1 U10813 ( .C1(n9543), .C2(n9542), .A(n10048), .B(n9541), .ZN(n9548)
         );
  OAI211_X1 U10814 ( .C1(n9546), .C2(n9545), .A(n9544), .B(n10047), .ZN(n9547)
         );
  NAND3_X1 U10815 ( .A1(n9549), .A2(n9548), .A3(n9547), .ZN(P1_U3251) );
  OAI211_X1 U10816 ( .C1(n9552), .C2(n9551), .A(n9550), .B(n10047), .ZN(n9562)
         );
  OAI211_X1 U10817 ( .C1(n9555), .C2(n9554), .A(n9553), .B(n10048), .ZN(n9561)
         );
  INV_X1 U10818 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9556) );
  NOR2_X1 U10819 ( .A1(n10070), .A2(n9556), .ZN(n9557) );
  AOI211_X1 U10820 ( .C1(n4409), .C2(n9559), .A(n9558), .B(n9557), .ZN(n9560)
         );
  NAND3_X1 U10821 ( .A1(n9562), .A2(n9561), .A3(n9560), .ZN(P1_U3254) );
  NAND2_X1 U10822 ( .A1(n9576), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9563) );
  NAND2_X1 U10823 ( .A1(n9564), .A2(n9563), .ZN(n10003) );
  NAND2_X1 U10824 ( .A1(n10006), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9565) );
  OAI21_X1 U10825 ( .B1(n10006), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9565), .ZN(
        n9566) );
  INV_X1 U10826 ( .A(n9566), .ZN(n10002) );
  NOR2_X1 U10827 ( .A1(n9567), .A2(n10015), .ZN(n9568) );
  INV_X1 U10828 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10020) );
  XNOR2_X1 U10829 ( .A(n10015), .B(n9567), .ZN(n10021) );
  NOR2_X1 U10830 ( .A1(n10020), .A2(n10021), .ZN(n10019) );
  NAND2_X1 U10831 ( .A1(n10037), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9569) );
  OAI21_X1 U10832 ( .B1(n10037), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9569), .ZN(
        n10029) );
  NOR2_X1 U10833 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  XNOR2_X1 U10834 ( .A(n10045), .B(n10312), .ZN(n10041) );
  NAND2_X1 U10835 ( .A1(n10042), .A2(n10041), .ZN(n9571) );
  NAND2_X1 U10836 ( .A1(n9583), .A2(n10312), .ZN(n9570) );
  NAND2_X1 U10837 ( .A1(n9571), .A2(n9570), .ZN(n10061) );
  NAND2_X1 U10838 ( .A1(n10065), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9572) );
  OAI21_X1 U10839 ( .B1(n10065), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9572), .ZN(
        n10062) );
  NAND2_X1 U10840 ( .A1(n10058), .A2(n9572), .ZN(n9573) );
  XNOR2_X1 U10841 ( .A(n9573), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9591) );
  INV_X1 U10842 ( .A(n9591), .ZN(n9589) );
  INV_X1 U10843 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9575) );
  AOI22_X1 U10844 ( .A1(n10037), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n9575), 
        .B2(n9574), .ZN(n10036) );
  NAND2_X1 U10845 ( .A1(n9576), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9577) );
  NAND2_X1 U10846 ( .A1(n9578), .A2(n9577), .ZN(n10001) );
  INV_X1 U10847 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9936) );
  XNOR2_X1 U10848 ( .A(n10006), .B(n9936), .ZN(n10000) );
  AOI21_X1 U10849 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10006), .A(n10009), 
        .ZN(n9579) );
  NOR2_X1 U10850 ( .A1(n9579), .A2(n10015), .ZN(n9580) );
  XNOR2_X1 U10851 ( .A(n10015), .B(n9579), .ZN(n10018) );
  NOR2_X1 U10852 ( .A1(n10017), .A2(n10018), .ZN(n10016) );
  NOR2_X1 U10853 ( .A1(n9580), .A2(n10016), .ZN(n10035) );
  NAND2_X1 U10854 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  OR2_X1 U10855 ( .A1(n10037), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U10856 ( .A1(n10034), .A2(n9581), .ZN(n10044) );
  INV_X1 U10857 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9582) );
  XNOR2_X1 U10858 ( .A(n10045), .B(n9582), .ZN(n10043) );
  NAND2_X1 U10859 ( .A1(n10044), .A2(n10043), .ZN(n9585) );
  NAND2_X1 U10860 ( .A1(n9583), .A2(n9582), .ZN(n9584) );
  NAND2_X1 U10861 ( .A1(n9585), .A2(n9584), .ZN(n10056) );
  NAND2_X1 U10862 ( .A1(n10065), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9586) );
  OAI21_X1 U10863 ( .B1(n10065), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9586), .ZN(
        n10057) );
  NAND2_X1 U10864 ( .A1(n10053), .A2(n9586), .ZN(n9587) );
  XNOR2_X1 U10865 ( .A(n9587), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9590) );
  AOI21_X1 U10866 ( .B1(n9590), .B2(n10047), .A(n4409), .ZN(n9588) );
  OAI21_X1 U10867 ( .B1(n9589), .B2(n10060), .A(n9588), .ZN(n9593) );
  OAI22_X1 U10868 ( .A1(n9591), .A2(n10060), .B1(n9590), .B2(n10055), .ZN(
        n9592) );
  NAND2_X1 U10869 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9594) );
  NAND2_X1 U10870 ( .A1(n9596), .A2(n10076), .ZN(n9599) );
  INV_X1 U10871 ( .A(n9864), .ZN(n9597) );
  NOR2_X1 U10872 ( .A1(n10084), .A2(n9597), .ZN(n9604) );
  AOI21_X1 U10873 ( .B1(P1_REG2_REG_31__SCAN_IN), .B2(n10084), .A(n9604), .ZN(
        n9598) );
  OAI211_X1 U10874 ( .C1(n9600), .C2(n9836), .A(n9599), .B(n9598), .ZN(
        P1_U3263) );
  NAND2_X1 U10875 ( .A1(n9865), .A2(n10076), .ZN(n9606) );
  AOI21_X1 U10876 ( .B1(n10084), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9604), .ZN(
        n9605) );
  OAI211_X1 U10877 ( .C1(n4804), .C2(n9836), .A(n9606), .B(n9605), .ZN(
        P1_U3264) );
  INV_X1 U10878 ( .A(n9607), .ZN(n9616) );
  NAND2_X1 U10879 ( .A1(n9608), .A2(n10076), .ZN(n9612) );
  INV_X1 U10880 ( .A(n9609), .ZN(n9610) );
  AOI22_X1 U10881 ( .A1(n9610), .A2(n10094), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10084), .ZN(n9611) );
  OAI211_X1 U10882 ( .C1(n9870), .C2(n9836), .A(n9612), .B(n9611), .ZN(n9613)
         );
  AOI21_X1 U10883 ( .B1(n9614), .B2(n9855), .A(n9613), .ZN(n9615) );
  OAI21_X1 U10884 ( .B1(n9616), .B2(n9850), .A(n9615), .ZN(P1_U3266) );
  AOI21_X1 U10885 ( .B1(n9618), .B2(n9846), .A(n9617), .ZN(n9872) );
  OR2_X1 U10886 ( .A1(n9873), .A2(n9850), .ZN(n9629) );
  OAI22_X1 U10887 ( .A1(n9622), .A2(n9852), .B1(n9621), .B2(n9855), .ZN(n9627)
         );
  OAI211_X1 U10888 ( .C1(n9625), .C2(n9623), .A(n9624), .B(n9782), .ZN(n9871)
         );
  NOR2_X1 U10889 ( .A1(n9871), .A2(n9783), .ZN(n9626) );
  AOI211_X1 U10890 ( .C1(n10074), .C2(n9950), .A(n9627), .B(n9626), .ZN(n9628)
         );
  OAI211_X1 U10891 ( .C1(n9872), .C2(n10084), .A(n9629), .B(n9628), .ZN(
        P1_U3267) );
  OAI211_X1 U10892 ( .C1(n9631), .C2(n9635), .A(n9630), .B(n9846), .ZN(n9633)
         );
  NAND2_X1 U10893 ( .A1(n9633), .A2(n9632), .ZN(n9875) );
  INV_X1 U10894 ( .A(n9875), .ZN(n9644) );
  XNOR2_X1 U10895 ( .A(n9634), .B(n9635), .ZN(n9877) );
  NAND2_X1 U10896 ( .A1(n9877), .A2(n10071), .ZN(n9643) );
  INV_X1 U10897 ( .A(n9651), .ZN(n9636) );
  AOI211_X1 U10898 ( .C1(n9637), .C2(n9636), .A(n9832), .B(n9623), .ZN(n9876)
         );
  NOR2_X1 U10899 ( .A1(n9955), .A2(n9836), .ZN(n9641) );
  OAI22_X1 U10900 ( .A1(n9639), .A2(n9852), .B1(n9638), .B2(n9855), .ZN(n9640)
         );
  AOI211_X1 U10901 ( .C1(n9876), .C2(n10076), .A(n9641), .B(n9640), .ZN(n9642)
         );
  OAI211_X1 U10902 ( .C1(n10084), .C2(n9644), .A(n9643), .B(n9642), .ZN(
        P1_U3268) );
  XNOR2_X1 U10903 ( .A(n9645), .B(n9646), .ZN(n9882) );
  INV_X1 U10904 ( .A(n9882), .ZN(n9658) );
  OAI211_X1 U10905 ( .C1(n9648), .C2(n5778), .A(n9846), .B(n9647), .ZN(n9650)
         );
  NAND2_X1 U10906 ( .A1(n9650), .A2(n9649), .ZN(n9880) );
  AOI211_X1 U10907 ( .C1(n9652), .C2(n9665), .A(n9832), .B(n9651), .ZN(n9881)
         );
  NAND2_X1 U10908 ( .A1(n9881), .A2(n10076), .ZN(n9655) );
  AOI22_X1 U10909 ( .A1(n9653), .A2(n10094), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n10084), .ZN(n9654) );
  OAI211_X1 U10910 ( .C1(n4798), .C2(n9836), .A(n9655), .B(n9654), .ZN(n9656)
         );
  AOI21_X1 U10911 ( .B1(n9855), .B2(n9880), .A(n9656), .ZN(n9657) );
  OAI21_X1 U10912 ( .B1(n9658), .B2(n9850), .A(n9657), .ZN(P1_U3269) );
  XNOR2_X1 U10913 ( .A(n9659), .B(n9664), .ZN(n9660) );
  NAND2_X1 U10914 ( .A1(n9660), .A2(n9846), .ZN(n9662) );
  NAND2_X1 U10915 ( .A1(n9662), .A2(n9661), .ZN(n9885) );
  INV_X1 U10916 ( .A(n9885), .ZN(n9674) );
  XNOR2_X1 U10917 ( .A(n9663), .B(n9664), .ZN(n9887) );
  NAND2_X1 U10918 ( .A1(n9887), .A2(n10071), .ZN(n9673) );
  INV_X1 U10919 ( .A(n9665), .ZN(n9666) );
  AOI211_X1 U10920 ( .C1(n9667), .C2(n4378), .A(n9832), .B(n9666), .ZN(n9886)
         );
  NOR2_X1 U10921 ( .A1(n9961), .A2(n9836), .ZN(n9671) );
  OAI22_X1 U10922 ( .A1(n9669), .A2(n9852), .B1(n9668), .B2(n9855), .ZN(n9670)
         );
  AOI211_X1 U10923 ( .C1(n9886), .C2(n10076), .A(n9671), .B(n9670), .ZN(n9672)
         );
  OAI211_X1 U10924 ( .C1(n10084), .C2(n9674), .A(n9673), .B(n9672), .ZN(
        P1_U3270) );
  NAND2_X1 U10925 ( .A1(n9675), .A2(n9676), .ZN(n9692) );
  NAND2_X1 U10926 ( .A1(n9692), .A2(n9703), .ZN(n9691) );
  NAND2_X1 U10927 ( .A1(n9691), .A2(n9677), .ZN(n9678) );
  XOR2_X1 U10928 ( .A(n9680), .B(n9678), .Z(n9892) );
  INV_X1 U10929 ( .A(n9892), .ZN(n9690) );
  XNOR2_X1 U10930 ( .A(n9679), .B(n9680), .ZN(n9682) );
  OAI21_X1 U10931 ( .B1(n9682), .B2(n9761), .A(n9681), .ZN(n9890) );
  AOI21_X1 U10932 ( .B1(n9696), .B2(n9683), .A(n9832), .ZN(n9684) );
  AND2_X1 U10933 ( .A1(n9684), .A2(n4378), .ZN(n9891) );
  NAND2_X1 U10934 ( .A1(n9891), .A2(n10076), .ZN(n9687) );
  AOI22_X1 U10935 ( .A1(n9685), .A2(n10094), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10084), .ZN(n9686) );
  OAI211_X1 U10936 ( .C1(n9965), .C2(n9836), .A(n9687), .B(n9686), .ZN(n9688)
         );
  AOI21_X1 U10937 ( .B1(n9890), .B2(n9855), .A(n9688), .ZN(n9689) );
  OAI21_X1 U10938 ( .B1(n9690), .B2(n9850), .A(n9689), .ZN(P1_U3271) );
  OAI21_X1 U10939 ( .B1(n9692), .B2(n9703), .A(n9691), .ZN(n9897) );
  OAI22_X1 U10940 ( .A1(n9694), .A2(n9852), .B1(n9855), .B2(n9693), .ZN(n9699)
         );
  OAI211_X1 U10941 ( .C1(n9695), .C2(n9697), .A(n9782), .B(n9696), .ZN(n9895)
         );
  NOR2_X1 U10942 ( .A1(n9895), .A2(n9783), .ZN(n9698) );
  AOI211_X1 U10943 ( .C1(n10074), .C2(n9968), .A(n9699), .B(n9698), .ZN(n9708)
         );
  INV_X1 U10944 ( .A(n9700), .ZN(n9702) );
  OAI21_X1 U10945 ( .B1(n9709), .B2(n9702), .A(n9701), .ZN(n9704) );
  XNOR2_X1 U10946 ( .A(n9704), .B(n9703), .ZN(n9706) );
  AOI21_X1 U10947 ( .B1(n9706), .B2(n9846), .A(n9705), .ZN(n9896) );
  OR2_X1 U10948 ( .A1(n9896), .A2(n10084), .ZN(n9707) );
  OAI211_X1 U10949 ( .C1(n9897), .C2(n9850), .A(n9708), .B(n9707), .ZN(
        P1_U3272) );
  XOR2_X1 U10950 ( .A(n9713), .B(n9709), .Z(n9711) );
  OAI21_X1 U10951 ( .B1(n9711), .B2(n9761), .A(n9710), .ZN(n9901) );
  INV_X1 U10952 ( .A(n9901), .ZN(n9721) );
  NAND2_X1 U10953 ( .A1(n9712), .A2(n9713), .ZN(n9904) );
  NAND3_X1 U10954 ( .A1(n9675), .A2(n10071), .A3(n9904), .ZN(n9720) );
  INV_X1 U10955 ( .A(n9723), .ZN(n9714) );
  AOI211_X1 U10956 ( .C1(n9903), .C2(n9714), .A(n9832), .B(n9695), .ZN(n9902)
         );
  AOI22_X1 U10957 ( .A1(n10084), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9715), 
        .B2(n10094), .ZN(n9716) );
  OAI21_X1 U10958 ( .B1(n9717), .B2(n9836), .A(n9716), .ZN(n9718) );
  AOI21_X1 U10959 ( .B1(n9902), .B2(n10076), .A(n9718), .ZN(n9719) );
  OAI211_X1 U10960 ( .C1(n10084), .C2(n9721), .A(n9720), .B(n9719), .ZN(
        P1_U3273) );
  XOR2_X1 U10961 ( .A(n9722), .B(n9729), .Z(n9911) );
  AOI211_X1 U10962 ( .C1(n9908), .C2(n9745), .A(n9832), .B(n9723), .ZN(n9907)
         );
  INV_X1 U10963 ( .A(n9724), .ZN(n9725) );
  AOI22_X1 U10964 ( .A1(n10084), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9725), 
        .B2(n10094), .ZN(n9726) );
  OAI21_X1 U10965 ( .B1(n4802), .B2(n9836), .A(n9726), .ZN(n9734) );
  OAI21_X1 U10966 ( .B1(n9729), .B2(n9728), .A(n9727), .ZN(n9732) );
  AOI222_X1 U10967 ( .A1(n9846), .A2(n9732), .B1(n9731), .B2(n9843), .C1(n9730), .C2(n9841), .ZN(n9910) );
  NOR2_X1 U10968 ( .A1(n9910), .A2(n10084), .ZN(n9733) );
  AOI211_X1 U10969 ( .C1(n9907), .C2(n10076), .A(n9734), .B(n9733), .ZN(n9735)
         );
  OAI21_X1 U10970 ( .B1(n9850), .B2(n9911), .A(n9735), .ZN(P1_U3274) );
  XOR2_X1 U10971 ( .A(n9736), .B(n9740), .Z(n9914) );
  INV_X1 U10972 ( .A(n9914), .ZN(n9753) );
  INV_X1 U10973 ( .A(n9738), .ZN(n9739) );
  AOI21_X1 U10974 ( .B1(n9740), .B2(n9737), .A(n9739), .ZN(n9741) );
  OAI222_X1 U10975 ( .A1(n9810), .A2(n9743), .B1(n9808), .B2(n9742), .C1(n9761), .C2(n9741), .ZN(n9912) );
  INV_X1 U10976 ( .A(n9745), .ZN(n9746) );
  AOI211_X1 U10977 ( .C1(n9747), .C2(n9744), .A(n9832), .B(n9746), .ZN(n9913)
         );
  NAND2_X1 U10978 ( .A1(n9913), .A2(n10076), .ZN(n9750) );
  AOI22_X1 U10979 ( .A1(n10084), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9748), 
        .B2(n10094), .ZN(n9749) );
  OAI211_X1 U10980 ( .C1(n4803), .C2(n9836), .A(n9750), .B(n9749), .ZN(n9751)
         );
  AOI21_X1 U10981 ( .B1(n9912), .B2(n9855), .A(n9751), .ZN(n9752) );
  OAI21_X1 U10982 ( .B1(n9753), .B2(n9850), .A(n9752), .ZN(P1_U3275) );
  XOR2_X1 U10983 ( .A(n9754), .B(n9760), .Z(n9921) );
  OAI22_X1 U10984 ( .A1(n9855), .A2(n10312), .B1(n9755), .B2(n9852), .ZN(n9768) );
  INV_X1 U10985 ( .A(n9744), .ZN(n9756) );
  AOI211_X1 U10986 ( .C1(n9919), .C2(n4323), .A(n9832), .B(n9756), .ZN(n9918)
         );
  NAND2_X1 U10987 ( .A1(n9770), .A2(n9758), .ZN(n9759) );
  XOR2_X1 U10988 ( .A(n9760), .B(n9759), .Z(n9762) );
  OAI222_X1 U10989 ( .A1(n9808), .A2(n9764), .B1(n9810), .B2(n9763), .C1(n9762), .C2(n9761), .ZN(n9917) );
  AOI21_X1 U10990 ( .B1(n9918), .B2(n9765), .A(n9917), .ZN(n9766) );
  NOR2_X1 U10991 ( .A1(n9766), .A2(n10084), .ZN(n9767) );
  AOI211_X1 U10992 ( .C1(n10074), .C2(n9919), .A(n9768), .B(n9767), .ZN(n9769)
         );
  OAI21_X1 U10993 ( .B1(n9850), .B2(n9921), .A(n9769), .ZN(P1_U3276) );
  OAI21_X1 U10994 ( .B1(n9778), .B2(n9771), .A(n9770), .ZN(n9774) );
  AOI222_X1 U10995 ( .A1(n9846), .A2(n9774), .B1(n9773), .B2(n9841), .C1(n9772), .C2(n9843), .ZN(n9926) );
  NAND2_X1 U10996 ( .A1(n9777), .A2(n9776), .ZN(n9779) );
  NAND2_X1 U10997 ( .A1(n9779), .A2(n9778), .ZN(n9922) );
  NAND3_X1 U10998 ( .A1(n9775), .A2(n9922), .A3(n10071), .ZN(n9787) );
  INV_X1 U10999 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9781) );
  OAI22_X1 U11000 ( .A1(n9855), .A2(n9781), .B1(n9780), .B2(n9852), .ZN(n9785)
         );
  OAI211_X1 U11001 ( .C1(n9307), .C2(n9789), .A(n4323), .B(n9782), .ZN(n9925)
         );
  NOR2_X1 U11002 ( .A1(n9925), .A2(n9783), .ZN(n9784) );
  AOI211_X1 U11003 ( .C1(n10074), .C2(n9923), .A(n9785), .B(n9784), .ZN(n9786)
         );
  OAI211_X1 U11004 ( .C1(n10084), .C2(n9926), .A(n9787), .B(n9786), .ZN(
        P1_U3277) );
  XNOR2_X1 U11005 ( .A(n9788), .B(n9796), .ZN(n9932) );
  AOI211_X1 U11006 ( .C1(n9929), .C2(n9817), .A(n9832), .B(n9789), .ZN(n9928)
         );
  INV_X1 U11007 ( .A(n9790), .ZN(n9791) );
  AOI22_X1 U11008 ( .A1(n10084), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9791), 
        .B2(n10094), .ZN(n9792) );
  OAI21_X1 U11009 ( .B1(n9793), .B2(n9836), .A(n9792), .ZN(n9800) );
  OAI21_X1 U11010 ( .B1(n9796), .B2(n9795), .A(n9794), .ZN(n9798) );
  AOI222_X1 U11011 ( .A1(n9846), .A2(n9798), .B1(n9797), .B2(n9843), .C1(n9844), .C2(n9841), .ZN(n9931) );
  NOR2_X1 U11012 ( .A1(n9931), .A2(n10084), .ZN(n9799) );
  AOI211_X1 U11013 ( .C1(n9928), .C2(n10076), .A(n9800), .B(n9799), .ZN(n9801)
         );
  OAI21_X1 U11014 ( .B1(n9932), .B2(n9850), .A(n9801), .ZN(P1_U3278) );
  OAI21_X1 U11015 ( .B1(n9802), .B2(n9804), .A(n9803), .ZN(n9935) );
  INV_X1 U11016 ( .A(n9935), .ZN(n9825) );
  OAI21_X1 U11017 ( .B1(n9807), .B2(n9806), .A(n9805), .ZN(n9813) );
  OAI22_X1 U11018 ( .A1(n9811), .A2(n9810), .B1(n9809), .B2(n9808), .ZN(n9812)
         );
  AOI21_X1 U11019 ( .B1(n9813), .B2(n9846), .A(n9812), .ZN(n9814) );
  OAI21_X1 U11020 ( .B1(n9825), .B2(n9815), .A(n9814), .ZN(n9933) );
  NAND2_X1 U11021 ( .A1(n9933), .A2(n9855), .ZN(n9823) );
  INV_X1 U11022 ( .A(n9817), .ZN(n9818) );
  AOI211_X1 U11023 ( .C1(n5616), .C2(n9816), .A(n9818), .B(n9832), .ZN(n9934)
         );
  INV_X1 U11024 ( .A(n5616), .ZN(n9982) );
  AOI22_X1 U11025 ( .A1(n10084), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9819), 
        .B2(n10094), .ZN(n9820) );
  OAI21_X1 U11026 ( .B1(n9982), .B2(n9836), .A(n9820), .ZN(n9821) );
  AOI21_X1 U11027 ( .B1(n9934), .B2(n10076), .A(n9821), .ZN(n9822) );
  OAI211_X1 U11028 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(
        P1_U3279) );
  OAI21_X1 U11029 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9829) );
  INV_X1 U11030 ( .A(n9829), .ZN(n9944) );
  INV_X1 U11031 ( .A(n9830), .ZN(n9833) );
  INV_X1 U11032 ( .A(n9816), .ZN(n9831) );
  AOI211_X1 U11033 ( .C1(n9939), .C2(n9833), .A(n9832), .B(n9831), .ZN(n9938)
         );
  AOI22_X1 U11034 ( .A1(n10084), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9834), 
        .B2(n10094), .ZN(n9835) );
  OAI21_X1 U11035 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9848) );
  OAI21_X1 U11036 ( .B1(n9840), .B2(n9839), .A(n9838), .ZN(n9845) );
  AOI222_X1 U11037 ( .A1(n9846), .A2(n9845), .B1(n9844), .B2(n9843), .C1(n9842), .C2(n9841), .ZN(n9942) );
  NOR2_X1 U11038 ( .A1(n9942), .A2(n10084), .ZN(n9847) );
  AOI211_X1 U11039 ( .C1(n9938), .C2(n10076), .A(n9848), .B(n9847), .ZN(n9849)
         );
  OAI21_X1 U11040 ( .B1(n9944), .B2(n9850), .A(n9849), .ZN(P1_U3280) );
  NAND2_X1 U11041 ( .A1(n9851), .A2(n9855), .ZN(n9863) );
  OAI22_X1 U11042 ( .A1(n9855), .A2(n9854), .B1(n9853), .B2(n9852), .ZN(n9856)
         );
  AOI21_X1 U11043 ( .B1(n10074), .B2(n9857), .A(n9856), .ZN(n9862) );
  NAND2_X1 U11044 ( .A1(n9858), .A2(n10071), .ZN(n9861) );
  NAND2_X1 U11045 ( .A1(n9859), .A2(n10076), .ZN(n9860) );
  NAND4_X1 U11046 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(
        P1_U3285) );
  INV_X1 U11047 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10318) );
  NOR2_X1 U11048 ( .A1(n9865), .A2(n9864), .ZN(n9946) );
  MUX2_X1 U11049 ( .A(n10318), .B(n9946), .S(n10117), .Z(n9866) );
  OAI21_X1 U11050 ( .B1(n4804), .B2(n6370), .A(n9866), .ZN(P1_U3552) );
  OAI21_X1 U11051 ( .B1(n9870), .B2(n6370), .A(n9869), .ZN(P1_U3549) );
  INV_X1 U11052 ( .A(n9874), .ZN(P1_U3548) );
  INV_X1 U11053 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9878) );
  AOI211_X1 U11054 ( .C1(n9877), .C2(n10113), .A(n9876), .B(n9875), .ZN(n9952)
         );
  MUX2_X1 U11055 ( .A(n9878), .B(n9952), .S(n10117), .Z(n9879) );
  OAI21_X1 U11056 ( .B1(n9955), .B2(n6370), .A(n9879), .ZN(P1_U3547) );
  INV_X1 U11057 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9883) );
  AOI211_X1 U11058 ( .C1(n9882), .C2(n10113), .A(n9881), .B(n9880), .ZN(n9956)
         );
  MUX2_X1 U11059 ( .A(n9883), .B(n9956), .S(n10117), .Z(n9884) );
  OAI21_X1 U11060 ( .B1(n4798), .B2(n6370), .A(n9884), .ZN(P1_U3546) );
  INV_X1 U11061 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9888) );
  AOI211_X1 U11062 ( .C1(n9887), .C2(n10113), .A(n9886), .B(n9885), .ZN(n9958)
         );
  MUX2_X1 U11063 ( .A(n9888), .B(n9958), .S(n10117), .Z(n9889) );
  OAI21_X1 U11064 ( .B1(n9961), .B2(n6370), .A(n9889), .ZN(P1_U3545) );
  INV_X1 U11065 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9893) );
  AOI211_X1 U11066 ( .C1(n9892), .C2(n10113), .A(n9891), .B(n9890), .ZN(n9962)
         );
  MUX2_X1 U11067 ( .A(n9893), .B(n9962), .S(n10117), .Z(n9894) );
  OAI21_X1 U11068 ( .B1(n9965), .B2(n6370), .A(n9894), .ZN(P1_U3544) );
  OAI211_X1 U11069 ( .C1(n9897), .C2(n9943), .A(n9896), .B(n9895), .ZN(n9966)
         );
  MUX2_X1 U11070 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9966), .S(n10117), .Z(
        n9898) );
  AOI21_X1 U11071 ( .B1(n9899), .B2(n9968), .A(n9898), .ZN(n9900) );
  INV_X1 U11072 ( .A(n9900), .ZN(P1_U3543) );
  AOI211_X1 U11073 ( .C1(n9940), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9906)
         );
  NAND3_X1 U11074 ( .A1(n9675), .A2(n10113), .A3(n9904), .ZN(n9905) );
  NAND2_X1 U11075 ( .A1(n9906), .A2(n9905), .ZN(n9970) );
  MUX2_X1 U11076 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9970), .S(n10117), .Z(
        P1_U3542) );
  AOI21_X1 U11077 ( .B1(n9940), .B2(n9908), .A(n9907), .ZN(n9909) );
  OAI211_X1 U11078 ( .C1(n9911), .C2(n9943), .A(n9910), .B(n9909), .ZN(n9971)
         );
  MUX2_X1 U11079 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9971), .S(n10117), .Z(
        P1_U3541) );
  INV_X1 U11080 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9915) );
  AOI211_X1 U11081 ( .C1(n9914), .C2(n10113), .A(n9913), .B(n9912), .ZN(n9972)
         );
  MUX2_X1 U11082 ( .A(n9915), .B(n9972), .S(n10117), .Z(n9916) );
  OAI21_X1 U11083 ( .B1(n4803), .B2(n6370), .A(n9916), .ZN(P1_U3540) );
  AOI211_X1 U11084 ( .C1(n9940), .C2(n9919), .A(n9918), .B(n9917), .ZN(n9920)
         );
  OAI21_X1 U11085 ( .B1(n9921), .B2(n9943), .A(n9920), .ZN(n9975) );
  MUX2_X1 U11086 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9975), .S(n10117), .Z(
        P1_U3539) );
  NAND3_X1 U11087 ( .A1(n9775), .A2(n9922), .A3(n10113), .ZN(n9927) );
  NAND2_X1 U11088 ( .A1(n9923), .A2(n9940), .ZN(n9924) );
  NAND4_X1 U11089 ( .A1(n9927), .A2(n9926), .A3(n9925), .A4(n9924), .ZN(n9976)
         );
  MUX2_X1 U11090 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9976), .S(n10117), .Z(
        P1_U3538) );
  AOI21_X1 U11091 ( .B1(n9940), .B2(n9929), .A(n9928), .ZN(n9930) );
  OAI211_X1 U11092 ( .C1(n9932), .C2(n9943), .A(n9931), .B(n9930), .ZN(n9977)
         );
  MUX2_X1 U11093 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9977), .S(n10117), .Z(
        P1_U3537) );
  AOI211_X1 U11094 ( .C1(n10105), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9978)
         );
  MUX2_X1 U11095 ( .A(n9936), .B(n9978), .S(n10117), .Z(n9937) );
  OAI21_X1 U11096 ( .B1(n9982), .B2(n6370), .A(n9937), .ZN(P1_U3536) );
  AOI21_X1 U11097 ( .B1(n9940), .B2(n9939), .A(n9938), .ZN(n9941) );
  OAI211_X1 U11098 ( .C1(n9944), .C2(n9943), .A(n9942), .B(n9941), .ZN(n9983)
         );
  MUX2_X1 U11099 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9983), .S(n10117), .Z(
        P1_U3535) );
  MUX2_X1 U11100 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9945), .S(n10117), .Z(
        P1_U3522) );
  INV_X1 U11101 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9947) );
  MUX2_X1 U11102 ( .A(n9947), .B(n9946), .S(n10348), .Z(n9948) );
  OAI21_X1 U11103 ( .B1(n4804), .B2(n9981), .A(n9948), .ZN(P1_U3520) );
  INV_X1 U11104 ( .A(n9951), .ZN(P1_U3516) );
  INV_X1 U11105 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9953) );
  MUX2_X1 U11106 ( .A(n9953), .B(n9952), .S(n10348), .Z(n9954) );
  OAI21_X1 U11107 ( .B1(n9955), .B2(n9981), .A(n9954), .ZN(P1_U3515) );
  MUX2_X1 U11108 ( .A(n10317), .B(n9956), .S(n10348), .Z(n9957) );
  OAI21_X1 U11109 ( .B1(n4798), .B2(n9981), .A(n9957), .ZN(P1_U3514) );
  INV_X1 U11110 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9959) );
  MUX2_X1 U11111 ( .A(n9959), .B(n9958), .S(n10348), .Z(n9960) );
  OAI21_X1 U11112 ( .B1(n9961), .B2(n9981), .A(n9960), .ZN(P1_U3513) );
  INV_X1 U11113 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n9963) );
  MUX2_X1 U11114 ( .A(n9963), .B(n9962), .S(n10348), .Z(n9964) );
  OAI21_X1 U11115 ( .B1(n9965), .B2(n9981), .A(n9964), .ZN(P1_U3512) );
  MUX2_X1 U11116 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9966), .S(n10348), .Z(
        n9967) );
  AOI21_X1 U11117 ( .B1(n6326), .B2(n9968), .A(n9967), .ZN(n9969) );
  INV_X1 U11118 ( .A(n9969), .ZN(P1_U3511) );
  MUX2_X1 U11119 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9970), .S(n10348), .Z(
        P1_U3510) );
  MUX2_X1 U11120 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9971), .S(n10348), .Z(
        P1_U3509) );
  INV_X1 U11121 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U11122 ( .A(n9973), .B(n9972), .S(n10348), .Z(n9974) );
  OAI21_X1 U11123 ( .B1(n4803), .B2(n9981), .A(n9974), .ZN(P1_U3507) );
  MUX2_X1 U11124 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9975), .S(n10348), .Z(
        P1_U3504) );
  MUX2_X1 U11125 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9976), .S(n10348), .Z(
        P1_U3501) );
  MUX2_X1 U11126 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9977), .S(n10348), .Z(
        P1_U3498) );
  INV_X1 U11127 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9979) );
  MUX2_X1 U11128 ( .A(n9979), .B(n9978), .S(n10348), .Z(n9980) );
  OAI21_X1 U11129 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(P1_U3495) );
  MUX2_X1 U11130 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9983), .S(n10348), .Z(
        P1_U3492) );
  MUX2_X1 U11131 ( .A(n9984), .B(P1_D_REG_1__SCAN_IN), .S(n10099), .Z(P1_U3440) );
  MUX2_X1 U11132 ( .A(n9985), .B(P1_D_REG_0__SCAN_IN), .S(n10099), .Z(P1_U3439) );
  NOR4_X1 U11133 ( .A1(n9986), .A2(P1_IR_REG_30__SCAN_IN), .A3(n5035), .A4(
        n10066), .ZN(n9987) );
  AOI21_X1 U11134 ( .B1(n9990), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9987), .ZN(
        n9988) );
  OAI21_X1 U11135 ( .B1(n9989), .B2(n9993), .A(n9988), .ZN(P1_U3324) );
  AOI22_X1 U11136 ( .A1(n9991), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9990), .ZN(n9992) );
  OAI21_X1 U11137 ( .B1(n9994), .B2(n9993), .A(n9992), .ZN(P1_U3325) );
  OAI222_X1 U11138 ( .A1(n9993), .A2(n9998), .B1(P1_U3086), .B2(n9997), .C1(
        n9996), .C2(n9995), .ZN(P1_U3326) );
  MUX2_X1 U11139 ( .A(n9999), .B(n4469), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11140 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11141 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11142 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10014) );
  OAI21_X1 U11143 ( .B1(n10001), .B2(n10000), .A(n10047), .ZN(n10010) );
  OAI21_X1 U11144 ( .B1(n10003), .B2(n10002), .A(n10048), .ZN(n10004) );
  OR2_X1 U11145 ( .A1(n10005), .A2(n10004), .ZN(n10008) );
  NAND2_X1 U11146 ( .A1(n4409), .A2(n10006), .ZN(n10007) );
  OAI211_X1 U11147 ( .C1(n10010), .C2(n10009), .A(n10008), .B(n10007), .ZN(
        n10011) );
  INV_X1 U11148 ( .A(n10011), .ZN(n10013) );
  OAI211_X1 U11149 ( .C1(n10070), .C2(n10014), .A(n10013), .B(n10012), .ZN(
        P1_U3257) );
  INV_X1 U11150 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10027) );
  INV_X1 U11151 ( .A(n10015), .ZN(n10024) );
  AOI211_X1 U11152 ( .C1(n10018), .C2(n10017), .A(n10016), .B(n10055), .ZN(
        n10023) );
  AOI211_X1 U11153 ( .C1(n10021), .C2(n10020), .A(n10019), .B(n10060), .ZN(
        n10022) );
  AOI211_X1 U11154 ( .C1(n4409), .C2(n10024), .A(n10023), .B(n10022), .ZN(
        n10026) );
  OAI211_X1 U11155 ( .C1(n10070), .C2(n10027), .A(n10026), .B(n10025), .ZN(
        P1_U3258) );
  AOI211_X1 U11156 ( .C1(n10030), .C2(n10029), .A(n10028), .B(n10060), .ZN(
        n10031) );
  AOI211_X1 U11157 ( .C1(n10033), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n10032), 
        .B(n10031), .ZN(n10040) );
  OAI21_X1 U11158 ( .B1(n10036), .B2(n10035), .A(n10034), .ZN(n10038) );
  AOI22_X1 U11159 ( .A1(n10038), .A2(n10047), .B1(n10037), .B2(n4409), .ZN(
        n10039) );
  NAND2_X1 U11160 ( .A1(n10040), .A2(n10039), .ZN(P1_U3259) );
  XNOR2_X1 U11161 ( .A(n10042), .B(n10041), .ZN(n10049) );
  XNOR2_X1 U11162 ( .A(n10044), .B(n10043), .ZN(n10046) );
  AOI222_X1 U11163 ( .A1(n10049), .A2(n10048), .B1(n10047), .B2(n10046), .C1(
        n10045), .C2(n4409), .ZN(n10051) );
  OAI211_X1 U11164 ( .C1(n10070), .C2(n10052), .A(n10051), .B(n10050), .ZN(
        P1_U3260) );
  INV_X1 U11165 ( .A(n10053), .ZN(n10054) );
  AOI211_X1 U11166 ( .C1(n10057), .C2(n10056), .A(n10055), .B(n10054), .ZN(
        n10064) );
  INV_X1 U11167 ( .A(n10058), .ZN(n10059) );
  AOI211_X1 U11168 ( .C1(n10062), .C2(n10061), .A(n10060), .B(n10059), .ZN(
        n10063) );
  AOI211_X1 U11169 ( .C1(n4409), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10068) );
  NAND2_X1 U11170 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(n10066), .ZN(n10067) );
  OAI211_X1 U11171 ( .C1(n10070), .C2(n10069), .A(n10068), .B(n10067), .ZN(
        P1_U3261) );
  NAND2_X1 U11172 ( .A1(n10072), .A2(n10071), .ZN(n10081) );
  NAND2_X1 U11173 ( .A1(n10074), .A2(n10073), .ZN(n10080) );
  AOI22_X1 U11174 ( .A1(n10076), .A2(n10075), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10094), .ZN(n10079) );
  OR2_X1 U11175 ( .A1(n9855), .A2(n10077), .ZN(n10078) );
  AND4_X1 U11176 ( .A1(n10081), .A2(n10080), .A3(n10079), .A4(n10078), .ZN(
        n10082) );
  OAI21_X1 U11177 ( .B1(n10084), .B2(n10083), .A(n10082), .ZN(P1_U3291) );
  NAND3_X1 U11178 ( .A1(n10087), .A2(n10086), .A3(n10085), .ZN(n10093) );
  NAND3_X1 U11179 ( .A1(n10090), .A2(n10089), .A3(n10088), .ZN(n10091) );
  NAND3_X1 U11180 ( .A1(n10093), .A2(n10092), .A3(n10091), .ZN(n10095) );
  AOI22_X1 U11181 ( .A1(n9855), .A2(n10095), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10094), .ZN(n10096) );
  OAI21_X1 U11182 ( .B1(n10097), .B2(n9855), .A(n10096), .ZN(P1_U3293) );
  AND2_X1 U11183 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10099), .ZN(P1_U3294) );
  AND2_X1 U11184 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10099), .ZN(P1_U3295) );
  AND2_X1 U11185 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10099), .ZN(P1_U3296) );
  AND2_X1 U11186 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10099), .ZN(P1_U3297) );
  AND2_X1 U11187 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10099), .ZN(P1_U3298) );
  AND2_X1 U11188 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10099), .ZN(P1_U3299) );
  AND2_X1 U11189 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10099), .ZN(P1_U3300) );
  AND2_X1 U11190 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10099), .ZN(P1_U3301) );
  AND2_X1 U11191 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10099), .ZN(P1_U3302) );
  AND2_X1 U11192 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10099), .ZN(P1_U3303) );
  AND2_X1 U11193 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10099), .ZN(P1_U3304) );
  AND2_X1 U11194 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10099), .ZN(P1_U3305) );
  INV_X1 U11195 ( .A(n10099), .ZN(n10098) );
  INV_X1 U11196 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U11197 ( .A1(n10098), .A2(n10327), .ZN(P1_U3306) );
  AND2_X1 U11198 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10099), .ZN(P1_U3307) );
  AND2_X1 U11199 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10099), .ZN(P1_U3308) );
  AND2_X1 U11200 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10099), .ZN(P1_U3309) );
  AND2_X1 U11201 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10099), .ZN(P1_U3310) );
  AND2_X1 U11202 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10099), .ZN(P1_U3311) );
  AND2_X1 U11203 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10099), .ZN(P1_U3312) );
  AND2_X1 U11204 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10099), .ZN(P1_U3313) );
  AND2_X1 U11205 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10099), .ZN(P1_U3314) );
  AND2_X1 U11206 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10099), .ZN(P1_U3315) );
  AND2_X1 U11207 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10099), .ZN(P1_U3316) );
  INV_X1 U11208 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U11209 ( .A1(n10098), .A2(n10271), .ZN(P1_U3317) );
  AND2_X1 U11210 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10099), .ZN(P1_U3318) );
  AND2_X1 U11211 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10099), .ZN(P1_U3319) );
  AND2_X1 U11212 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10099), .ZN(P1_U3320) );
  AND2_X1 U11213 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10099), .ZN(P1_U3321) );
  INV_X1 U11214 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10272) );
  NOR2_X1 U11215 ( .A1(n10098), .A2(n10272), .ZN(P1_U3322) );
  AND2_X1 U11216 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10099), .ZN(P1_U3323) );
  OAI21_X1 U11217 ( .B1(n10101), .B2(n10110), .A(n10100), .ZN(n10103) );
  AOI211_X1 U11218 ( .C1(n10105), .C2(n10104), .A(n10103), .B(n10102), .ZN(
        n10108) );
  INV_X1 U11219 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10106) );
  AOI22_X1 U11220 ( .A1(n10348), .A2(n10108), .B1(n10106), .B2(n10346), .ZN(
        P1_U3456) );
  INV_X1 U11221 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11222 ( .A1(n10117), .A2(n10108), .B1(n10107), .B2(n10118), .ZN(
        P1_U3523) );
  OAI21_X1 U11223 ( .B1(n10111), .B2(n10110), .A(n10109), .ZN(n10112) );
  AOI21_X1 U11224 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10115) );
  NAND2_X1 U11225 ( .A1(n10116), .A2(n10115), .ZN(n10347) );
  OAI22_X1 U11226 ( .A1(n10118), .A2(n10347), .B1(P1_REG1_REG_3__SCAN_IN), 
        .B2(n10117), .ZN(n10119) );
  INV_X1 U11227 ( .A(n10119), .ZN(P1_U3525) );
  INV_X1 U11228 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10125) );
  INV_X1 U11229 ( .A(n10120), .ZN(n10124) );
  OAI21_X1 U11230 ( .B1(n10122), .B2(n10150), .A(n10121), .ZN(n10123) );
  AOI21_X1 U11231 ( .B1(n10153), .B2(n10124), .A(n10123), .ZN(n10158) );
  AOI22_X1 U11232 ( .A1(n10156), .A2(n10125), .B1(n10158), .B2(n10155), .ZN(
        P2_U3393) );
  OAI22_X1 U11233 ( .A1(n10128), .A2(n10127), .B1(n10126), .B2(n10150), .ZN(
        n10129) );
  NOR2_X1 U11234 ( .A1(n10130), .A2(n10129), .ZN(n10159) );
  AOI22_X1 U11235 ( .A1(n10156), .A2(n5851), .B1(n10159), .B2(n10155), .ZN(
        P2_U3396) );
  INV_X1 U11236 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10137) );
  INV_X1 U11237 ( .A(n10131), .ZN(n10136) );
  OAI22_X1 U11238 ( .A1(n10134), .A2(n10133), .B1(n10132), .B2(n10150), .ZN(
        n10135) );
  NOR2_X1 U11239 ( .A1(n10136), .A2(n10135), .ZN(n10161) );
  AOI22_X1 U11240 ( .A1(n10156), .A2(n10137), .B1(n10161), .B2(n10155), .ZN(
        P2_U3399) );
  INV_X1 U11241 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10142) );
  OAI21_X1 U11242 ( .B1(n10139), .B2(n10150), .A(n10138), .ZN(n10140) );
  AOI21_X1 U11243 ( .B1(n10153), .B2(n10141), .A(n10140), .ZN(n10163) );
  AOI22_X1 U11244 ( .A1(n10156), .A2(n10142), .B1(n10163), .B2(n10155), .ZN(
        P2_U3402) );
  AOI22_X1 U11245 ( .A1(n10146), .A2(n10145), .B1(n10144), .B2(n10143), .ZN(
        n10147) );
  AND2_X1 U11246 ( .A1(n10148), .A2(n10147), .ZN(n10164) );
  AOI22_X1 U11247 ( .A1(n10156), .A2(n5918), .B1(n10164), .B2(n10155), .ZN(
        P2_U3405) );
  OAI21_X1 U11248 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10152) );
  AOI21_X1 U11249 ( .B1(n10154), .B2(n10153), .A(n10152), .ZN(n10167) );
  AOI22_X1 U11250 ( .A1(n10156), .A2(n5924), .B1(n10167), .B2(n10155), .ZN(
        P2_U3408) );
  AOI22_X1 U11251 ( .A1(n10168), .A2(n10158), .B1(n10157), .B2(n10165), .ZN(
        P2_U3460) );
  AOI22_X1 U11252 ( .A1(n10168), .A2(n10159), .B1(n10331), .B2(n10165), .ZN(
        P2_U3461) );
  AOI22_X1 U11253 ( .A1(n10168), .A2(n10161), .B1(n10160), .B2(n10165), .ZN(
        P2_U3462) );
  AOI22_X1 U11254 ( .A1(n10168), .A2(n10163), .B1(n10162), .B2(n10165), .ZN(
        P2_U3463) );
  AOI22_X1 U11255 ( .A1(n10168), .A2(n10164), .B1(n4776), .B2(n10165), .ZN(
        P2_U3464) );
  INV_X1 U11256 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10166) );
  AOI22_X1 U11257 ( .A1(n10168), .A2(n10167), .B1(n10166), .B2(n10165), .ZN(
        P2_U3465) );
  OAI222_X1 U11258 ( .A1(n10173), .A2(n10172), .B1(n10173), .B2(n10171), .C1(
        n10170), .C2(n10169), .ZN(ADD_1068_U5) );
  XOR2_X1 U11259 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11260 ( .A(n10176), .ZN(n10175) );
  OAI222_X1 U11261 ( .A1(n10178), .A2(n10177), .B1(n10178), .B2(n10176), .C1(
        n10175), .C2(n10174), .ZN(ADD_1068_U55) );
  OAI21_X1 U11262 ( .B1(n10181), .B2(n10180), .A(n10179), .ZN(ADD_1068_U56) );
  OAI21_X1 U11263 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1068_U57) );
  OAI21_X1 U11264 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(ADD_1068_U58) );
  OAI21_X1 U11265 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(ADD_1068_U59) );
  OAI21_X1 U11266 ( .B1(n10193), .B2(n10192), .A(n10191), .ZN(ADD_1068_U60) );
  OAI21_X1 U11267 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(ADD_1068_U61) );
  OAI21_X1 U11268 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(ADD_1068_U62) );
  OAI21_X1 U11269 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(ADD_1068_U63) );
  NAND4_X1 U11270 ( .A1(SI_28_), .A2(P1_DATAO_REG_4__SCAN_IN), .A3(
        P1_REG3_REG_8__SCAN_IN), .A4(n5896), .ZN(n10210) );
  INV_X1 U11271 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10203) );
  NAND4_X1 U11272 ( .A1(n10203), .A2(P2_D_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_23__SCAN_IN), .A4(P1_REG0_REG_3__SCAN_IN), .ZN(n10209) );
  NAND4_X1 U11273 ( .A1(n10205), .A2(n10204), .A3(n10301), .A4(SI_15_), .ZN(
        n10208) );
  INV_X1 U11274 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10287) );
  NAND4_X1 U11275 ( .A1(n10206), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n7443), 
        .A4(n10287), .ZN(n10207) );
  NOR4_X1 U11276 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10345) );
  NOR4_X1 U11277 ( .A1(P1_REG2_REG_1__SCAN_IN), .A2(P2_REG1_REG_23__SCAN_IN), 
        .A3(n10211), .A4(n10331), .ZN(n10215) );
  NOR4_X1 U11278 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), 
        .A3(P2_REG1_REG_29__SCAN_IN), .A4(n10328), .ZN(n10214) );
  NOR4_X1 U11279 ( .A1(P1_REG0_REG_19__SCAN_IN), .A2(n10317), .A3(n10327), 
        .A4(n10318), .ZN(n10213) );
  NOR4_X1 U11280 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P1_REG0_REG_29__SCAN_IN), 
        .A3(P1_REG2_REG_17__SCAN_IN), .A4(P2_REG0_REG_31__SCAN_IN), .ZN(n10212) );
  NAND4_X1 U11281 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10229) );
  NOR4_X1 U11282 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .A4(P2_REG1_REG_11__SCAN_IN), .ZN(n10219)
         );
  NOR4_X1 U11283 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .A3(P1_REG2_REG_10__SCAN_IN), .A4(n10262), .ZN(n10218) );
  INV_X1 U11284 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10246) );
  AND4_X1 U11285 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P2_REG2_REG_7__SCAN_IN), 
        .A3(n10216), .A4(n10246), .ZN(n10217) );
  NAND4_X1 U11286 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10219), .A3(n10218), .A4(
        n10217), .ZN(n10220) );
  NOR4_X1 U11287 ( .A1(n10272), .A2(n10220), .A3(n10234), .A4(
        P1_D_REG_8__SCAN_IN), .ZN(n10222) );
  NOR4_X1 U11288 ( .A1(n10231), .A2(n10233), .A3(P1_REG2_REG_20__SCAN_IN), 
        .A4(P1_REG1_REG_12__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U11289 ( .A1(n10222), .A2(n10221), .ZN(n10228) );
  NOR4_X1 U11290 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), 
        .A3(P1_IR_REG_10__SCAN_IN), .A4(P1_IR_REG_26__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U11291 ( .A1(n10223), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U11292 ( .A1(n10225), .A2(P2_REG1_REG_20__SCAN_IN), .A3(
        P2_REG3_REG_27__SCAN_IN), .A4(n10224), .ZN(n10227) );
  NAND4_X1 U11293 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n5851), .A3(n10243), .A4(
        n10257), .ZN(n10226) );
  NOR4_X1 U11294 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10344) );
  AOI22_X1 U11295 ( .A1(n10231), .A2(keyinput42), .B1(keyinput35), .B2(
        P2_U3151), .ZN(n10230) );
  OAI221_X1 U11296 ( .B1(n10231), .B2(keyinput42), .C1(P2_U3151), .C2(
        keyinput35), .A(n10230), .ZN(n10241) );
  AOI22_X1 U11297 ( .A1(n5667), .A2(keyinput32), .B1(n10233), .B2(keyinput9), 
        .ZN(n10232) );
  OAI221_X1 U11298 ( .B1(n5667), .B2(keyinput32), .C1(n10233), .C2(keyinput9), 
        .A(n10232), .ZN(n10240) );
  XOR2_X1 U11299 ( .A(n10234), .B(keyinput40), .Z(n10238) );
  XNOR2_X1 U11300 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput29), .ZN(n10237) );
  XNOR2_X1 U11301 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput19), .ZN(n10236) );
  XNOR2_X1 U11302 ( .A(P2_REG1_REG_7__SCAN_IN), .B(keyinput22), .ZN(n10235) );
  NAND4_X1 U11303 ( .A1(n10238), .A2(n10237), .A3(n10236), .A4(n10235), .ZN(
        n10239) );
  NOR3_X1 U11304 ( .A1(n10241), .A2(n10240), .A3(n10239), .ZN(n10285) );
  AOI22_X1 U11305 ( .A1(n5851), .A2(keyinput48), .B1(n10243), .B2(keyinput6), 
        .ZN(n10242) );
  OAI221_X1 U11306 ( .B1(n5851), .B2(keyinput48), .C1(n10243), .C2(keyinput6), 
        .A(n10242), .ZN(n10255) );
  AOI22_X1 U11307 ( .A1(n10246), .A2(keyinput55), .B1(keyinput56), .B2(n10245), 
        .ZN(n10244) );
  OAI221_X1 U11308 ( .B1(n10246), .B2(keyinput55), .C1(n10245), .C2(keyinput56), .A(n10244), .ZN(n10254) );
  AOI22_X1 U11309 ( .A1(n10249), .A2(keyinput5), .B1(n10248), .B2(keyinput3), 
        .ZN(n10247) );
  OAI221_X1 U11310 ( .B1(n10249), .B2(keyinput5), .C1(n10248), .C2(keyinput3), 
        .A(n10247), .ZN(n10253) );
  XNOR2_X1 U11311 ( .A(P2_REG2_REG_25__SCAN_IN), .B(keyinput0), .ZN(n10251) );
  XNOR2_X1 U11312 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput47), .ZN(n10250) );
  NAND2_X1 U11313 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  NOR4_X1 U11314 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10284) );
  AOI22_X1 U11315 ( .A1(n10258), .A2(keyinput20), .B1(keyinput43), .B2(n10257), 
        .ZN(n10256) );
  OAI221_X1 U11316 ( .B1(n10258), .B2(keyinput20), .C1(n10257), .C2(keyinput43), .A(n10256), .ZN(n10269) );
  INV_X1 U11317 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U11318 ( .A1(n10261), .A2(keyinput37), .B1(keyinput7), .B2(n10260), 
        .ZN(n10259) );
  OAI221_X1 U11319 ( .B1(n10261), .B2(keyinput37), .C1(n10260), .C2(keyinput7), 
        .A(n10259), .ZN(n10268) );
  XOR2_X1 U11320 ( .A(n10262), .B(keyinput57), .Z(n10266) );
  XNOR2_X1 U11321 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput36), .ZN(n10265)
         );
  XNOR2_X1 U11322 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput51), .ZN(n10264) );
  XNOR2_X1 U11323 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(keyinput2), .ZN(n10263)
         );
  NAND4_X1 U11324 ( .A1(n10266), .A2(n10265), .A3(n10264), .A4(n10263), .ZN(
        n10267) );
  NOR3_X1 U11325 ( .A1(n10269), .A2(n10268), .A3(n10267), .ZN(n10283) );
  AOI22_X1 U11326 ( .A1(n10272), .A2(keyinput23), .B1(keyinput25), .B2(n10271), 
        .ZN(n10270) );
  OAI221_X1 U11327 ( .B1(n10272), .B2(keyinput23), .C1(n10271), .C2(keyinput25), .A(n10270), .ZN(n10281) );
  XNOR2_X1 U11328 ( .A(n10273), .B(keyinput49), .ZN(n10280) );
  XOR2_X1 U11329 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(keyinput59), .Z(n10279) );
  XNOR2_X1 U11330 ( .A(P2_REG1_REG_11__SCAN_IN), .B(keyinput8), .ZN(n10277) );
  XNOR2_X1 U11331 ( .A(P2_IR_REG_26__SCAN_IN), .B(keyinput15), .ZN(n10276) );
  XNOR2_X1 U11332 ( .A(P2_REG1_REG_20__SCAN_IN), .B(keyinput28), .ZN(n10275)
         );
  XNOR2_X1 U11333 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput24), .ZN(n10274) );
  NAND4_X1 U11334 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10278) );
  NOR4_X1 U11335 ( .A1(n10281), .A2(n10280), .A3(n10279), .A4(n10278), .ZN(
        n10282) );
  NAND4_X1 U11336 ( .A1(n10285), .A2(n10284), .A3(n10283), .A4(n10282), .ZN(
        n10343) );
  INV_X1 U11337 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n10286) );
  XOR2_X1 U11338 ( .A(n10286), .B(keyinput34), .Z(n10291) );
  XOR2_X1 U11339 ( .A(n10287), .B(keyinput27), .Z(n10290) );
  XNOR2_X1 U11340 ( .A(SI_8_), .B(keyinput1), .ZN(n10289) );
  XNOR2_X1 U11341 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput17), .ZN(n10288)
         );
  NAND4_X1 U11342 ( .A1(n10291), .A2(n10290), .A3(n10289), .A4(n10288), .ZN(
        n10297) );
  XNOR2_X1 U11343 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput53), .ZN(n10295) );
  XNOR2_X1 U11344 ( .A(P1_REG0_REG_13__SCAN_IN), .B(keyinput63), .ZN(n10294)
         );
  XNOR2_X1 U11345 ( .A(P2_REG0_REG_8__SCAN_IN), .B(keyinput38), .ZN(n10293) );
  XNOR2_X1 U11346 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput58), .ZN(n10292)
         );
  NAND4_X1 U11347 ( .A1(n10295), .A2(n10294), .A3(n10293), .A4(n10292), .ZN(
        n10296) );
  NOR2_X1 U11348 ( .A1(n10297), .A2(n10296), .ZN(n10341) );
  AOI22_X1 U11349 ( .A1(n5391), .A2(keyinput11), .B1(keyinput33), .B2(n5896), 
        .ZN(n10298) );
  OAI221_X1 U11350 ( .B1(n5391), .B2(keyinput11), .C1(n5896), .C2(keyinput33), 
        .A(n10298), .ZN(n10309) );
  AOI22_X1 U11351 ( .A1(n10301), .A2(keyinput4), .B1(n10300), .B2(keyinput31), 
        .ZN(n10299) );
  OAI221_X1 U11352 ( .B1(n10301), .B2(keyinput4), .C1(n10300), .C2(keyinput31), 
        .A(n10299), .ZN(n10308) );
  INV_X1 U11353 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10302) );
  XOR2_X1 U11354 ( .A(n10302), .B(keyinput41), .Z(n10306) );
  XOR2_X1 U11355 ( .A(n7443), .B(keyinput39), .Z(n10305) );
  XNOR2_X1 U11356 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput60), .ZN(n10304) );
  XNOR2_X1 U11357 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput14), .ZN(n10303) );
  NAND4_X1 U11358 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10307) );
  NOR3_X1 U11359 ( .A1(n10309), .A2(n10308), .A3(n10307), .ZN(n10340) );
  AOI22_X1 U11360 ( .A1(n10312), .A2(keyinput18), .B1(n10311), .B2(keyinput54), 
        .ZN(n10310) );
  OAI221_X1 U11361 ( .B1(n10312), .B2(keyinput18), .C1(n10311), .C2(keyinput54), .A(n10310), .ZN(n10324) );
  AOI22_X1 U11362 ( .A1(n10315), .A2(keyinput16), .B1(keyinput26), .B2(n10314), 
        .ZN(n10313) );
  OAI221_X1 U11363 ( .B1(n10315), .B2(keyinput16), .C1(n10314), .C2(keyinput26), .A(n10313), .ZN(n10323) );
  AOI22_X1 U11364 ( .A1(n10318), .A2(keyinput52), .B1(n10317), .B2(keyinput12), 
        .ZN(n10316) );
  OAI221_X1 U11365 ( .B1(n10318), .B2(keyinput52), .C1(n10317), .C2(keyinput12), .A(n10316), .ZN(n10322) );
  XNOR2_X1 U11366 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(keyinput44), .ZN(n10320)
         );
  XNOR2_X1 U11367 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput45), .ZN(n10319) );
  NAND2_X1 U11368 ( .A1(n10320), .A2(n10319), .ZN(n10321) );
  NOR4_X1 U11369 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10339) );
  AOI22_X1 U11370 ( .A1(n6420), .A2(keyinput21), .B1(n5044), .B2(keyinput13), 
        .ZN(n10325) );
  OAI221_X1 U11371 ( .B1(n6420), .B2(keyinput21), .C1(n5044), .C2(keyinput13), 
        .A(n10325), .ZN(n10337) );
  AOI22_X1 U11372 ( .A1(n10328), .A2(keyinput62), .B1(n10327), .B2(keyinput61), 
        .ZN(n10326) );
  OAI221_X1 U11373 ( .B1(n10328), .B2(keyinput62), .C1(n10327), .C2(keyinput61), .A(n10326), .ZN(n10336) );
  AOI22_X1 U11374 ( .A1(n10331), .A2(keyinput50), .B1(n10330), .B2(keyinput46), 
        .ZN(n10329) );
  OAI221_X1 U11375 ( .B1(n10331), .B2(keyinput50), .C1(n10330), .C2(keyinput46), .A(n10329), .ZN(n10335) );
  XNOR2_X1 U11376 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput10), .ZN(n10333) );
  XNOR2_X1 U11377 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput30), .ZN(n10332) );
  NAND2_X1 U11378 ( .A1(n10333), .A2(n10332), .ZN(n10334) );
  NOR4_X1 U11379 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10338) );
  NAND4_X1 U11380 ( .A1(n10341), .A2(n10340), .A3(n10339), .A4(n10338), .ZN(
        n10342) );
  AOI211_X1 U11381 ( .C1(n10345), .C2(n10344), .A(n10343), .B(n10342), .ZN(
        n10350) );
  AOI22_X1 U11382 ( .A1(n10348), .A2(n10347), .B1(P1_REG0_REG_3__SCAN_IN), 
        .B2(n10346), .ZN(n10349) );
  XNOR2_X1 U11383 ( .A(n10350), .B(n10349), .ZN(P1_U3462) );
  OAI21_X1 U11384 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(ADD_1068_U50) );
  OAI21_X1 U11385 ( .B1(n10356), .B2(n10355), .A(n10354), .ZN(ADD_1068_U51) );
  OAI21_X1 U11386 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(ADD_1068_U47) );
  OAI21_X1 U11387 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(ADD_1068_U49) );
  OAI21_X1 U11388 ( .B1(n10365), .B2(n10364), .A(n10363), .ZN(ADD_1068_U48) );
  AOI21_X1 U11389 ( .B1(n10368), .B2(n10367), .A(n10366), .ZN(ADD_1068_U54) );
  AOI21_X1 U11390 ( .B1(n10371), .B2(n10370), .A(n10369), .ZN(ADD_1068_U53) );
  OAI21_X1 U11391 ( .B1(n10374), .B2(n10373), .A(n10372), .ZN(ADD_1068_U52) );
  NAND2_X1 U4806 ( .A1(n4431), .A2(n6677), .ZN(n8922) );
  CLKBUF_X1 U4807 ( .A(n6685), .Z(n4299) );
  CLKBUF_X1 U4811 ( .A(n8999), .Z(n9112) );
  NAND2_X1 U4815 ( .A1(n6491), .A2(n6677), .ZN(n8948) );
endmodule

