

module b21_C_SARLock_k_64_4 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, 
        ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, 
        ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, 
        ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, 
        U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, 
        P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, 
        P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, 
        P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, 
        P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, 
        P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, 
        P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, 
        P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, 
        P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, 
        P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, 
        P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, 
        P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, 
        P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, 
        P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, 
        P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, 
        P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, 
        P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, 
        P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, 
        P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, 
        P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, 
        P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, 
        P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, 
        P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, 
        P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, 
        P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, 
        P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, 
        P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, 
        P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, 
        P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, 
        P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, 
        P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, 
        P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, 
        P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, 
        P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, 
        P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, 
        P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, 
        P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, 
        P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000;

  OR2_X1 U4750 ( .A1(n7949), .A2(n7948), .ZN(n4279) );
  AND2_X1 U4751 ( .A1(n9051), .A2(n9015), .ZN(n9029) );
  AOI21_X1 U4752 ( .B1(n8527), .B2(n8534), .A(n4377), .ZN(n8513) );
  INV_X1 U4753 ( .A(n5651), .ZN(n6045) );
  BUF_X2 U4756 ( .A(n5621), .Z(n6152) );
  CLKBUF_X2 U4757 ( .A(n5236), .Z(n7683) );
  NAND2_X1 U4758 ( .A1(n9697), .A2(n6358), .ZN(n7726) );
  NAND2_X1 U4759 ( .A1(n4895), .A2(n4503), .ZN(n6851) );
  AND2_X2 U4760 ( .A1(n7981), .A2(n8720), .ZN(n5621) );
  XNOR2_X1 U4761 ( .A(n6049), .B(P2_IR_REG_22__SCAN_IN), .ZN(n5580) );
  CLKBUF_X2 U4762 ( .A(n5184), .Z(n6567) );
  NAND2_X1 U4763 ( .A1(n4865), .A2(n4866), .ZN(n9584) );
  NOR2_X2 U4764 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4828) );
  CLKBUF_X3 U4765 ( .A(n5651), .Z(n6024) );
  NAND2_X1 U4766 ( .A1(n8079), .A2(n4386), .ZN(n8169) );
  AND2_X1 U4768 ( .A1(n8503), .A2(n8497), .ZN(n8498) );
  NAND2_X1 U4769 ( .A1(n9806), .A2(n7592), .ZN(n9805) );
  XNOR2_X1 U4770 ( .A(n8868), .B(n6397), .ZN(n7770) );
  NAND2_X1 U4771 ( .A1(n7865), .A2(n7863), .ZN(n7776) );
  INV_X1 U4772 ( .A(n8817), .ZN(n9748) );
  AND3_X1 U4773 ( .A1(n4912), .A2(n4913), .A3(n4670), .ZN(n9730) );
  INV_X1 U4774 ( .A(n6335), .ZN(n6775) );
  NAND2_X1 U4775 ( .A1(n7966), .A2(n5846), .ZN(n7971) );
  NAND2_X1 U4776 ( .A1(n5562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5560) );
  OR2_X1 U4777 ( .A1(n5585), .A2(n4559), .ZN(n4558) );
  NAND2_X2 U4778 ( .A1(n5040), .A2(n5039), .ZN(n7705) );
  CLKBUF_X3 U4779 ( .A(n4940), .Z(n7680) );
  OAI21_X1 U4780 ( .B1(n6671), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6668), .ZN(
        n6985) );
  OAI21_X1 U4781 ( .B1(n4967), .B2(n6629), .A(n4885), .ZN(n7080) );
  NAND4_X2 U4782 ( .A1(n4860), .A2(n4859), .A3(n4858), .A4(n4857), .ZN(n6363)
         );
  AND4_X2 U4783 ( .A1(n5715), .A2(n5550), .A3(n5781), .A4(n5782), .ZN(n4268)
         );
  INV_X4 U4784 ( .A(n8017), .ZN(n4244) );
  NAND2_X4 U4785 ( .A1(n5536), .A2(n6927), .ZN(n4266) );
  NAND4_X2 U4786 ( .A1(n4883), .A2(n4882), .A3(n4881), .A4(n4880), .ZN(n6346)
         );
  XNOR2_X2 U4787 ( .A(n5963), .B(n5961), .ZN(n8183) );
  OAI222_X1 U4788 ( .A1(P2_U3152), .A2(n7981), .B1(n8719), .B2(n9412), .C1(
        n7980), .C2(n8722), .ZN(P2_U3328) );
  NOR2_X2 U4789 ( .A1(n9807), .A2(n9928), .ZN(n4599) );
  NAND2_X2 U4790 ( .A1(n5145), .A2(n5144), .ZN(n7673) );
  XNOR2_X2 U4791 ( .A(n5074), .B(n4822), .ZN(n6664) );
  OAI21_X2 U4792 ( .B1(n6289), .B2(n4744), .A(n7040), .ZN(n5651) );
  NAND2_X2 U4793 ( .A1(n5303), .A2(n5302), .ZN(n9216) );
  XNOR2_X1 U4794 ( .A(n7705), .B(n8864), .ZN(n9674) );
  OR2_X1 U4795 ( .A1(n8971), .A2(n8972), .ZN(n8974) );
  NAND2_X1 U4796 ( .A1(n9043), .A2(n9042), .ZN(n9041) );
  AOI211_X1 U4797 ( .C1(n9244), .C2(n9203), .A(n9202), .B(n9201), .ZN(n9204)
         );
  NAND2_X1 U4798 ( .A1(n4260), .A2(n4245), .ZN(n8792) );
  AOI21_X1 U4799 ( .B1(n9051), .B2(n5392), .A(n4823), .ZN(n9000) );
  NAND2_X2 U4800 ( .A1(n7695), .A2(n9085), .ZN(n9097) );
  NAND2_X1 U4801 ( .A1(n7561), .A2(n5834), .ZN(n5848) );
  AND2_X1 U4802 ( .A1(n4258), .A2(n6416), .ZN(n6421) );
  NAND2_X1 U4803 ( .A1(n7088), .A2(n7087), .ZN(n4258) );
  NAND2_X2 U4804 ( .A1(n5508), .A2(n7847), .ZN(n7845) );
  OAI21_X1 U4805 ( .B1(n5030), .B2(n5029), .A(n5028), .ZN(n5050) );
  NAND2_X1 U4806 ( .A1(n7185), .A2(n8817), .ZN(n7831) );
  NAND2_X1 U4807 ( .A1(n7799), .A2(n7197), .ZN(n9694) );
  XNOR2_X1 U4808 ( .A(n4265), .B(n6361), .ZN(n6368) );
  NAND2_X2 U4809 ( .A1(n7726), .A2(n7723), .ZN(n7764) );
  AND2_X1 U4810 ( .A1(n6342), .A2(n4247), .ZN(n6374) );
  INV_X1 U4811 ( .A(n8867), .ZN(n7185) );
  INV_X1 U4812 ( .A(n7941), .ZN(n7943) );
  NAND3_X1 U4813 ( .A1(n4918), .A2(n4917), .A3(n4916), .ZN(n8869) );
  INV_X1 U4814 ( .A(n6363), .ZN(n9697) );
  INV_X2 U4815 ( .A(n6357), .ZN(n4247) );
  INV_X1 U4816 ( .A(n6830), .ZN(n6112) );
  AND2_X1 U4817 ( .A1(n9413), .A2(n4856), .ZN(n4934) );
  NAND2_X1 U4818 ( .A1(n4854), .A2(n4856), .ZN(n4940) );
  INV_X1 U4819 ( .A(n4853), .ZN(n4856) );
  INV_X1 U4820 ( .A(n5622), .ZN(n5610) );
  MUX2_X1 U4821 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4861), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n4863) );
  OAI21_X1 U4822 ( .B1(n5447), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5462) );
  INV_X4 U4823 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U4824 ( .A(n8626), .ZN(n4593) );
  OAI21_X1 U4825 ( .B1(n4594), .B2(n8533), .A(n8006), .ZN(n8626) );
  NAND2_X1 U4826 ( .A1(n8824), .A2(n6520), .ZN(n8828) );
  XNOR2_X1 U4827 ( .A(n8001), .B(n4475), .ZN(n4594) );
  AND2_X1 U4828 ( .A1(n4592), .A2(n4362), .ZN(n4591) );
  NAND2_X1 U4829 ( .A1(n8743), .A2(n8744), .ZN(n8824) );
  NAND2_X1 U4830 ( .A1(n8773), .A2(n6509), .ZN(n8743) );
  NAND2_X1 U4831 ( .A1(n4792), .A2(n8725), .ZN(n8773) );
  NAND2_X1 U4832 ( .A1(n9041), .A2(n4296), .ZN(n9025) );
  NAND2_X1 U4833 ( .A1(n8791), .A2(n8794), .ZN(n6502) );
  NAND2_X1 U4834 ( .A1(n4263), .A2(n6497), .ZN(n8791) );
  INV_X1 U4835 ( .A(n4263), .ZN(n4260) );
  AND2_X1 U4836 ( .A1(n9003), .A2(n4552), .ZN(n8978) );
  NOR2_X1 U4837 ( .A1(n8627), .A2(n4326), .ZN(n4362) );
  NAND2_X1 U4838 ( .A1(n8733), .A2(n6496), .ZN(n4263) );
  OR2_X1 U4839 ( .A1(n9000), .A2(n8999), .ZN(n9003) );
  NOR2_X2 U4840 ( .A1(n9180), .A2(n8984), .ZN(n8966) );
  AOI21_X1 U4841 ( .B1(n6475), .B2(n4405), .A(n6489), .ZN(n4409) );
  OR2_X2 U4842 ( .A1(n9096), .A2(n9097), .ZN(n9094) );
  NAND2_X1 U4843 ( .A1(n8765), .A2(n6471), .ZN(n8804) );
  NAND2_X1 U4844 ( .A1(n4543), .A2(n4546), .ZN(n9096) );
  NAND2_X1 U4845 ( .A1(n6085), .A2(n6084), .ZN(n8630) );
  NAND3_X1 U4846 ( .A1(n4251), .A2(n4389), .A3(n4249), .ZN(n8765) );
  NAND2_X1 U4847 ( .A1(n7652), .A2(n7872), .ZN(n7651) );
  XNOR2_X1 U4848 ( .A(n5430), .B(n5429), .ZN(n8721) );
  NAND2_X1 U4849 ( .A1(n9151), .A2(n5241), .ZN(n9150) );
  NAND2_X1 U4850 ( .A1(n4250), .A2(n6464), .ZN(n4249) );
  OR2_X1 U4851 ( .A1(n8838), .A2(n4390), .ZN(n4251) );
  NAND3_X1 U4852 ( .A1(n7971), .A2(n7972), .A3(n5866), .ZN(n8122) );
  INV_X1 U4853 ( .A(n8839), .ZN(n4250) );
  NAND2_X1 U4854 ( .A1(n4379), .A2(n4381), .ZN(n7972) );
  NAND2_X1 U4855 ( .A1(n4252), .A2(n6456), .ZN(n8839) );
  NAND2_X1 U4856 ( .A1(n9805), .A2(n7593), .ZN(n7594) );
  NAND2_X1 U4857 ( .A1(n5848), .A2(n5847), .ZN(n7966) );
  INV_X1 U4858 ( .A(n6497), .ZN(n4245) );
  NAND2_X1 U4859 ( .A1(n7424), .A2(n4308), .ZN(n4393) );
  OAI21_X1 U4860 ( .B1(n9510), .B2(n7760), .A(n7761), .ZN(n7498) );
  NAND2_X1 U4861 ( .A1(n4269), .A2(n4396), .ZN(n4397) );
  NAND2_X1 U4862 ( .A1(n5296), .A2(n5295), .ZN(n5315) );
  NAND2_X1 U4863 ( .A1(n4258), .A2(n4257), .ZN(n4259) );
  NAND2_X1 U4864 ( .A1(n5169), .A2(n5168), .ZN(n8851) );
  AND2_X1 U4865 ( .A1(n4320), .A2(n6416), .ZN(n4257) );
  NAND2_X1 U4866 ( .A1(n5193), .A2(n5192), .ZN(n8762) );
  NAND2_X1 U4867 ( .A1(n5821), .A2(n5820), .ZN(n7620) );
  OAI21_X1 U4868 ( .B1(n5222), .B2(n4647), .A(n4644), .ZN(n5267) );
  NAND2_X1 U4869 ( .A1(n7009), .A2(n4799), .ZN(n4388) );
  NAND2_X1 U4870 ( .A1(n5080), .A2(n5079), .ZN(n7459) );
  NAND2_X1 U4871 ( .A1(n5124), .A2(n5123), .ZN(n9486) );
  NAND2_X1 U4872 ( .A1(n5102), .A2(n5101), .ZN(n7507) );
  AND2_X1 U4873 ( .A1(n7706), .A2(n7835), .ZN(n7839) );
  OR2_X1 U4874 ( .A1(n6415), .A2(n6414), .ZN(n6416) );
  NAND2_X1 U4875 ( .A1(n5135), .A2(n5134), .ZN(n5137) );
  NAND2_X1 U4876 ( .A1(n5018), .A2(n5017), .ZN(n7313) );
  NAND2_X1 U4877 ( .A1(n4993), .A2(n4992), .ZN(n7130) );
  INV_X1 U4878 ( .A(n6399), .ZN(n4246) );
  NAND2_X1 U4879 ( .A1(n6687), .A2(n6351), .ZN(n6695) );
  AND2_X1 U4880 ( .A1(n7204), .A2(n9745), .ZN(n7323) );
  NAND3_X1 U4881 ( .A1(n6765), .A2(n6792), .A3(n5609), .ZN(n8064) );
  NAND2_X1 U4882 ( .A1(n6349), .A2(n6348), .ZN(n6686) );
  AND2_X1 U4883 ( .A1(n5686), .A2(n5685), .ZN(n7109) );
  INV_X1 U4884 ( .A(n6374), .ZN(n6440) );
  INV_X1 U4885 ( .A(n8869), .ZN(n9699) );
  NAND4_X2 U4886 ( .A1(n4946), .A2(n4945), .A3(n4944), .A4(n4943), .ZN(n8868)
         );
  NAND2_X1 U4887 ( .A1(n5451), .A2(n5450), .ZN(n9701) );
  NAND3_X1 U4888 ( .A1(n4903), .A2(n4902), .A3(n4901), .ZN(n8870) );
  NAND2_X1 U4889 ( .A1(n5534), .A2(n6842), .ZN(n6339) );
  NAND2_X1 U4890 ( .A1(n4952), .A2(n4951), .ZN(n4972) );
  OR2_X1 U4891 ( .A1(n4940), .A2(n4855), .ZN(n4858) );
  INV_X1 U4892 ( .A(n6114), .ZN(n6759) );
  AND4_X1 U4893 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), .ZN(n7020)
         );
  AND3_X1 U4894 ( .A1(n5634), .A2(n5633), .A3(n5632), .ZN(n9818) );
  NAND4_X1 U4895 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5624), .ZN(n8236)
         );
  NAND2_X1 U4896 ( .A1(n4568), .A2(n4276), .ZN(n6807) );
  NAND2_X1 U4897 ( .A1(n4853), .A2(n4854), .ZN(n5236) );
  XNOR2_X1 U4898 ( .A(n4256), .B(P1_IR_REG_19__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U4899 ( .A1(n6334), .A2(n6590), .ZN(n8017) );
  NAND2_X1 U4900 ( .A1(n5474), .A2(n4392), .ZN(n6590) );
  INV_X1 U4901 ( .A(n4253), .ZN(n4256) );
  AND2_X2 U4902 ( .A1(n9413), .A2(n4853), .ZN(n4935) );
  NAND2_X4 U4903 ( .A1(n7959), .A2(n9584), .ZN(n4967) );
  INV_X1 U4904 ( .A(n9413), .ZN(n4854) );
  AOI21_X1 U4905 ( .B1(n5207), .B2(P1_IR_REG_31__SCAN_IN), .A(n4254), .ZN(
        n4253) );
  OAI21_X1 U4906 ( .B1(n5207), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5253) );
  AND2_X2 U4907 ( .A1(n5565), .A2(n5564), .ZN(n5640) );
  AND2_X1 U4908 ( .A1(n4851), .A2(n9407), .ZN(n9413) );
  NAND2_X1 U4909 ( .A1(n5471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5463) );
  OR2_X1 U4910 ( .A1(n5469), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5471) );
  XNOR2_X1 U4911 ( .A(n5462), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7956) );
  NAND2_X1 U4912 ( .A1(n5563), .A2(n5562), .ZN(n8720) );
  MUX2_X1 U4913 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5561), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n5563) );
  INV_X2 U4914 ( .A(n8715), .ZN(n8719) );
  AND2_X1 U4915 ( .A1(n4248), .A2(n5057), .ZN(n5099) );
  NOR2_X1 U4916 ( .A1(n5036), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n4248) );
  NAND2_X2 U4917 ( .A1(n6567), .A2(P1_U3084), .ZN(n6758) );
  NAND2_X1 U4918 ( .A1(n5252), .A2(n4255), .ZN(n4254) );
  NOR2_X1 U4919 ( .A1(n4957), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n4989) );
  NAND3_X1 U4920 ( .A1(n8959), .A2(n4350), .A3(n4349), .ZN(n4867) );
  AND4_X1 U4921 ( .A1(n5549), .A2(n5547), .A3(n5548), .A4(n5546), .ZN(n4783)
         );
  XNOR2_X1 U4922 ( .A(n4521), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6639) );
  INV_X1 U4923 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4830) );
  INV_X1 U4924 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5444) );
  INV_X1 U4925 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4349) );
  INV_X1 U4926 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U4927 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), 
        .ZN(n4255) );
  INV_X2 U4928 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND3_X1 U4929 ( .A1(n6349), .A2(n6348), .A3(n6350), .ZN(n6687) );
  INV_X1 U4930 ( .A(n4248), .ZN(n5037) );
  OAI21_X2 U4931 ( .B1(n7665), .B2(n7668), .A(n7666), .ZN(n4252) );
  NOR2_X2 U4932 ( .A1(n6454), .A2(n6453), .ZN(n7665) );
  NOR2_X2 U4933 ( .A1(n4252), .A2(n6456), .ZN(n8838) );
  NAND2_X1 U4934 ( .A1(n6454), .A2(n6453), .ZN(n7666) );
  NAND2_X2 U4935 ( .A1(n4259), .A2(n4802), .ZN(n7424) );
  OAI21_X1 U4936 ( .B1(n4263), .B2(n4262), .A(n4261), .ZN(n6505) );
  NAND2_X1 U4937 ( .A1(n8794), .A2(n4245), .ZN(n4261) );
  NOR2_X1 U4938 ( .A1(n8794), .A2(n4245), .ZN(n4262) );
  OR2_X1 U4939 ( .A1(n4264), .A2(n6399), .ZN(n6400) );
  XNOR2_X2 U4940 ( .A(n4264), .B(n4246), .ZN(n7009) );
  NAND2_X1 U4941 ( .A1(n6393), .A2(n6392), .ZN(n4264) );
  AND2_X1 U4942 ( .A1(n9669), .A2(n9760), .ZN(n9671) );
  NOR2_X2 U4943 ( .A1(n7154), .A2(n7313), .ZN(n9669) );
  NAND2_X1 U4944 ( .A1(n5534), .A2(n7393), .ZN(n5536) );
  NOR2_X2 U4945 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5589) );
  NAND2_X2 U4946 ( .A1(n5584), .A2(n5583), .ZN(n6092) );
  NAND4_X2 U4947 ( .A1(n4828), .A2(n4829), .A3(n4831), .A4(n4830), .ZN(n4957)
         );
  NOR2_X4 U4948 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n4829) );
  INV_X1 U4949 ( .A(n4266), .ZN(n4265) );
  OR2_X2 U4950 ( .A1(n8993), .A2(n8982), .ZN(n8984) );
  NAND2_X1 U4951 ( .A1(n6590), .A2(n6927), .ZN(n6357) );
  OR2_X1 U4952 ( .A1(n9203), .A2(n5390), .ZN(n9017) );
  NAND2_X1 U4953 ( .A1(n9203), .A2(n5390), .ZN(n9016) );
  NAND2_X1 U4954 ( .A1(n9097), .A2(n5524), .ZN(n4720) );
  NAND2_X1 U4955 ( .A1(n4623), .A2(n4622), .ZN(n6142) );
  AOI21_X1 U4956 ( .B1(n4625), .B2(n4627), .A(n4339), .ZN(n4622) );
  NAND2_X1 U4957 ( .A1(n5411), .A2(n4625), .ZN(n4623) );
  INV_X1 U4958 ( .A(n4935), .ZN(n5231) );
  NOR2_X1 U4959 ( .A1(n4712), .A2(n7786), .ZN(n4711) );
  INV_X1 U4960 ( .A(n5529), .ZN(n4712) );
  OAI211_X1 U4961 ( .C1(n4977), .C2(n6575), .A(n4877), .B(n4876), .ZN(n6358)
         );
  NAND2_X1 U4962 ( .A1(n4455), .A2(n4454), .ZN(n4453) );
  NAND2_X1 U4963 ( .A1(n7898), .A2(n7941), .ZN(n4455) );
  AOI211_X1 U4964 ( .C1(n7899), .C2(n7943), .A(n9097), .B(n4547), .ZN(n4454)
         );
  NAND2_X1 U4965 ( .A1(n4466), .A2(n4467), .ZN(n4464) );
  AOI21_X1 U4966 ( .B1(n4470), .B2(n4270), .A(n4466), .ZN(n4465) );
  OR2_X1 U4967 ( .A1(n8618), .A2(n6166), .ZN(n6287) );
  OR2_X1 U4968 ( .A1(n8982), .A2(n9001), .ZN(n7928) );
  INV_X1 U4969 ( .A(n4691), .ZN(n4690) );
  NAND2_X1 U4970 ( .A1(n5050), .A2(n4323), .ZN(n5052) );
  INV_X1 U4971 ( .A(n6012), .ZN(n6010) );
  OR2_X1 U4972 ( .A1(n7620), .A2(n8225), .ZN(n7989) );
  NAND2_X1 U4973 ( .A1(n7255), .A2(n7260), .ZN(n7356) );
  NAND2_X1 U4974 ( .A1(n5557), .A2(n4787), .ZN(n4786) );
  INV_X1 U4975 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4787) );
  NOR2_X1 U4976 ( .A1(n4411), .A2(n4407), .ZN(n4406) );
  NOR2_X1 U4977 ( .A1(n4408), .A2(n4414), .ZN(n4407) );
  NAND2_X1 U4978 ( .A1(n8982), .A2(n9001), .ZN(n7929) );
  NAND2_X1 U4979 ( .A1(n7928), .A2(n7929), .ZN(n8975) );
  OR2_X1 U4980 ( .A1(n9191), .A2(n8025), .ZN(n7924) );
  NOR2_X1 U4981 ( .A1(n9196), .A2(n8856), .ZN(n7786) );
  OR2_X1 U4982 ( .A1(n9216), .A2(n9100), .ZN(n7906) );
  NAND2_X1 U4983 ( .A1(n4696), .A2(n4698), .ZN(n7628) );
  INV_X1 U4984 ( .A(n4699), .ZN(n4698) );
  OAI21_X1 U4985 ( .B1(n5515), .B2(n4700), .A(n5514), .ZN(n4699) );
  NAND2_X1 U4986 ( .A1(n5396), .A2(n5395), .ZN(n5411) );
  AOI21_X1 U4987 ( .B1(n4636), .B2(n4322), .A(n4634), .ZN(n4633) );
  NAND2_X1 U4988 ( .A1(n5333), .A2(n5332), .ZN(n5335) );
  OAI21_X1 U4989 ( .B1(n5267), .B2(n5266), .A(n5265), .ZN(n5282) );
  AND2_X1 U4990 ( .A1(n5283), .A2(n5272), .ZN(n5281) );
  AND2_X1 U4991 ( .A1(n5205), .A2(n5188), .ZN(n5203) );
  NAND2_X1 U4992 ( .A1(n5181), .A2(n5163), .ZN(n5182) );
  OR2_X1 U4993 ( .A1(n5736), .A2(n5735), .ZN(n5754) );
  NAND2_X1 U4994 ( .A1(n5580), .A2(n8377), .ZN(n6811) );
  AND2_X1 U4995 ( .A1(n5960), .A2(n5959), .ZN(n8106) );
  INV_X1 U4996 ( .A(n7981), .ZN(n5564) );
  NOR2_X1 U4997 ( .A1(n9451), .A2(n9450), .ZN(n9449) );
  NAND2_X1 U4998 ( .A1(n8642), .A2(n8111), .ZN(n8421) );
  OR2_X1 U4999 ( .A1(n8661), .A2(n8106), .ZN(n6259) );
  OR2_X1 U5000 ( .A1(n8671), .A2(n8101), .ZN(n8515) );
  AND2_X1 U5001 ( .A1(n7616), .A2(n4287), .ZN(n4781) );
  INV_X1 U5002 ( .A(n6087), .ZN(n9866) );
  INV_X1 U5003 ( .A(n9021), .ZN(n8025) );
  AOI21_X1 U5004 ( .B1(n6346), .B2(n4244), .A(n6345), .ZN(n6689) );
  INV_X1 U5005 ( .A(n7683), .ZN(n5419) );
  INV_X1 U5006 ( .A(n4940), .ZN(n5420) );
  OR2_X1 U5007 ( .A1(n9203), .A2(n9054), .ZN(n5529) );
  INV_X1 U5008 ( .A(n9028), .ZN(n4713) );
  NAND2_X1 U5009 ( .A1(n4536), .A2(n4539), .ZN(n9050) );
  AOI21_X1 U5010 ( .B1(n9069), .B2(n4541), .A(n4540), .ZN(n4539) );
  NAND2_X1 U5011 ( .A1(n9094), .A2(n4537), .ZN(n4536) );
  INV_X1 U5012 ( .A(n7906), .ZN(n4541) );
  AOI21_X1 U5013 ( .B1(n4719), .B2(n5525), .A(n4273), .ZN(n4718) );
  NAND2_X1 U5014 ( .A1(n4930), .A2(n9695), .ZN(n4933) );
  NAND2_X1 U5015 ( .A1(n5437), .A2(n5436), .ZN(n9180) );
  AND2_X1 U5016 ( .A1(n4819), .A2(n4847), .ZN(n4817) );
  OAI21_X1 U5017 ( .B1(n4708), .B2(n5447), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4864) );
  NAND2_X1 U5018 ( .A1(n4709), .A2(n4818), .ZN(n4708) );
  CLKBUF_X1 U5019 ( .A(n5534), .Z(n5254) );
  NAND2_X1 U5020 ( .A1(n5996), .A2(n5995), .ZN(n8646) );
  NAND2_X1 U5021 ( .A1(n7567), .A2(n5713), .ZN(n5996) );
  XNOR2_X1 U5022 ( .A(n4374), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U5023 ( .A1(n8949), .A2(n4375), .ZN(n4374) );
  OR2_X1 U5024 ( .A1(n8950), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n4375) );
  AOI21_X1 U5025 ( .B1(n5459), .B2(n9701), .A(n5458), .ZN(n9182) );
  AND2_X1 U5026 ( .A1(n6307), .A2(n6288), .ZN(n4461) );
  INV_X1 U5027 ( .A(n4450), .ZN(n4449) );
  OAI21_X1 U5028 ( .B1(n7844), .B2(n7943), .A(n7846), .ZN(n4450) );
  MUX2_X1 U5029 ( .A(n6237), .B(n6236), .S(n6279), .Z(n6238) );
  AOI21_X1 U5030 ( .B1(n4459), .B2(n4289), .A(n4456), .ZN(n6240) );
  NOR2_X1 U5031 ( .A1(n7868), .A2(n7943), .ZN(n4447) );
  OAI21_X1 U5032 ( .B1(n7869), .B2(n7941), .A(n7870), .ZN(n4446) );
  NAND2_X1 U5033 ( .A1(n4484), .A2(n4482), .ZN(n4481) );
  NOR2_X1 U5034 ( .A1(n8482), .A2(n4483), .ZN(n4482) );
  INV_X1 U5035 ( .A(n6266), .ZN(n4665) );
  AND2_X1 U5036 ( .A1(n6274), .A2(n6273), .ZN(n4476) );
  NAND2_X1 U5037 ( .A1(n4366), .A2(n4365), .ZN(n6274) );
  NAND2_X1 U5038 ( .A1(n6272), .A2(n6288), .ZN(n4365) );
  OR2_X1 U5039 ( .A1(n6271), .A2(n4367), .ZN(n4366) );
  AND2_X1 U5040 ( .A1(n6270), .A2(n6267), .ZN(n4659) );
  NAND2_X1 U5041 ( .A1(n4663), .A2(n4661), .ZN(n4660) );
  AND2_X1 U5042 ( .A1(n4278), .A2(n6021), .ZN(n4725) );
  NOR2_X1 U5043 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5546) );
  NOR2_X1 U5044 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5551) );
  OR3_X1 U5045 ( .A1(n7911), .A2(n7699), .A3(n7698), .ZN(n7814) );
  AND2_X1 U5046 ( .A1(n7845), .A2(n4693), .ZN(n4688) );
  NAND2_X1 U5047 ( .A1(n5221), .A2(n5225), .ZN(n4648) );
  NAND2_X1 U5048 ( .A1(n5033), .A2(n9357), .ZN(n5051) );
  NAND2_X1 U5049 ( .A1(n5012), .A2(n5011), .ZN(n5028) );
  NAND2_X1 U5050 ( .A1(n6087), .A2(n7372), .ZN(n4744) );
  AND2_X1 U5051 ( .A1(n8625), .A2(n4578), .ZN(n4577) );
  NAND2_X1 U5052 ( .A1(n6280), .A2(n4582), .ZN(n4578) );
  OR2_X1 U5053 ( .A1(n4579), .A2(n4577), .ZN(n4576) );
  INV_X1 U5054 ( .A(n4580), .ZN(n4579) );
  OAI22_X1 U5055 ( .A1(n6284), .A2(n4581), .B1(n8383), .B2(n7372), .ZN(n4580)
         );
  NAND2_X1 U5056 ( .A1(n4582), .A2(n6280), .ZN(n4581) );
  NAND2_X1 U5057 ( .A1(n4473), .A2(n6280), .ZN(n4583) );
  INV_X1 U5058 ( .A(n6285), .ZN(n4364) );
  INV_X1 U5059 ( .A(n6287), .ZN(n4493) );
  AND2_X1 U5060 ( .A1(n4435), .A2(n8326), .ZN(n4432) );
  OR2_X1 U5061 ( .A1(n8630), .A2(n8045), .ZN(n6273) );
  NOR2_X1 U5062 ( .A1(n8642), .A2(n4759), .ZN(n4758) );
  INV_X1 U5063 ( .A(n8111), .ZN(n4759) );
  OR2_X1 U5064 ( .A1(n8642), .A2(n8111), .ZN(n6270) );
  OR2_X1 U5065 ( .A1(n5998), .A2(n5997), .ZN(n6012) );
  NOR2_X1 U5066 ( .A1(n8646), .A2(n4610), .ZN(n4609) );
  INV_X1 U5067 ( .A(n4611), .ZN(n4610) );
  XNOR2_X1 U5068 ( .A(n8646), .B(n8472), .ZN(n7997) );
  OR2_X1 U5069 ( .A1(n8650), .A2(n8220), .ZN(n6264) );
  INV_X1 U5070 ( .A(n8504), .ZN(n6134) );
  OR2_X1 U5071 ( .A1(n8681), .A2(n8224), .ZN(n4766) );
  NOR2_X1 U5072 ( .A1(n8569), .A2(n4768), .ZN(n4767) );
  INV_X1 U5073 ( .A(n4769), .ZN(n4768) );
  NOR2_X1 U5074 ( .A1(n8584), .A2(n4770), .ZN(n4769) );
  INV_X1 U5075 ( .A(n4824), .ZN(n4770) );
  XNOR2_X1 U5076 ( .A(n7976), .B(n4668), .ZN(n6224) );
  NAND2_X1 U5077 ( .A1(n6222), .A2(n6221), .ZN(n6120) );
  OR2_X1 U5078 ( .A1(n9928), .A2(n7600), .ZN(n6307) );
  INV_X1 U5079 ( .A(n6303), .ZN(n4566) );
  OAI21_X1 U5080 ( .B1(n6304), .B2(n4566), .A(n6293), .ZN(n4565) );
  INV_X1 U5081 ( .A(n7169), .ZN(n4761) );
  NAND2_X1 U5082 ( .A1(n4570), .A2(n4569), .ZN(n7171) );
  NAND2_X1 U5083 ( .A1(n4309), .A2(n6118), .ZN(n4569) );
  NAND2_X1 U5084 ( .A1(n7045), .A2(n4357), .ZN(n4570) );
  NAND2_X1 U5085 ( .A1(n7411), .A2(n7372), .ZN(n6087) );
  INV_X1 U5086 ( .A(n5569), .ZN(n4486) );
  NOR2_X1 U5087 ( .A1(n5556), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n4487) );
  INV_X1 U5088 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4350) );
  INV_X1 U5089 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4378) );
  INV_X1 U5090 ( .A(n4811), .ZN(n4810) );
  NAND2_X1 U5091 ( .A1(n7290), .A2(n4809), .ZN(n4808) );
  INV_X1 U5092 ( .A(n7933), .ZN(n7791) );
  AND2_X1 U5093 ( .A1(n5391), .A2(n9017), .ZN(n7915) );
  NOR2_X1 U5094 ( .A1(n9111), .A2(n4550), .ZN(n4549) );
  INV_X1 U5095 ( .A(n4549), .ZN(n4548) );
  INV_X1 U5096 ( .A(n7892), .ZN(n4545) );
  OR2_X1 U5097 ( .A1(n9223), .A2(n8795), .ZN(n7695) );
  NAND2_X1 U5098 ( .A1(n4707), .A2(n9486), .ZN(n4704) );
  NOR2_X1 U5099 ( .A1(n9486), .A2(n4707), .ZN(n4706) );
  OR2_X1 U5100 ( .A1(n7673), .A2(n9495), .ZN(n7865) );
  OR2_X1 U5101 ( .A1(n5082), .A2(n5081), .ZN(n5105) );
  INV_X1 U5102 ( .A(n9674), .ZN(n4525) );
  NAND2_X1 U5103 ( .A1(n4529), .A2(n7835), .ZN(n4526) );
  NAND2_X1 U5104 ( .A1(n7706), .A2(n4530), .ZN(n4529) );
  OR2_X1 U5105 ( .A1(n4531), .A2(n7833), .ZN(n4530) );
  NAND2_X1 U5106 ( .A1(n7835), .A2(n7830), .ZN(n4527) );
  NOR2_X1 U5107 ( .A1(n5501), .A2(n4678), .ZN(n4673) );
  INV_X1 U5108 ( .A(n5503), .ZN(n4678) );
  INV_X1 U5109 ( .A(n7839), .ZN(n5504) );
  NAND2_X1 U5110 ( .A1(n4995), .A2(n4994), .ZN(n5020) );
  AND2_X1 U5111 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n4994) );
  INV_X1 U5112 ( .A(n4998), .ZN(n4995) );
  INV_X1 U5113 ( .A(n9730), .ZN(n6375) );
  NAND2_X1 U5114 ( .A1(n5496), .A2(n6375), .ZN(n7799) );
  NAND2_X1 U5115 ( .A1(n9730), .A2(n8870), .ZN(n7197) );
  NAND2_X1 U5116 ( .A1(n6146), .A2(n6145), .ZN(n6157) );
  OR2_X1 U5117 ( .A1(n6142), .A2(n6141), .ZN(n6146) );
  NOR2_X1 U5118 ( .A1(n5352), .A2(n4641), .ZN(n4640) );
  INV_X1 U5119 ( .A(n5334), .ZN(n4641) );
  OAI21_X1 U5120 ( .B1(n5315), .B2(n5314), .A(n5313), .ZN(n5333) );
  AND2_X1 U5121 ( .A1(n5334), .A2(n5320), .ZN(n5332) );
  NAND2_X1 U5122 ( .A1(n5206), .A2(n5205), .ZN(n5222) );
  AOI21_X1 U5123 ( .B1(n4653), .B2(n4655), .A(n4651), .ZN(n4650) );
  NAND2_X1 U5124 ( .A1(n4613), .A2(n4616), .ZN(n5114) );
  AOI21_X1 U5125 ( .B1(n4617), .B2(n4619), .A(n4328), .ZN(n4616) );
  NAND2_X1 U5126 ( .A1(n5112), .A2(n5097), .ZN(n5113) );
  XNOR2_X1 U5127 ( .A(n5091), .B(n5076), .ZN(n5090) );
  XNOR2_X1 U5128 ( .A(n5008), .B(SI_7_), .ZN(n5005) );
  NAND2_X1 U5129 ( .A1(n4986), .A2(n4985), .ZN(n5007) );
  INV_X1 U5130 ( .A(n4981), .ZN(n4982) );
  NOR2_X1 U5131 ( .A1(n6555), .A2(n4385), .ZN(n4384) );
  INV_X1 U5132 ( .A(n5801), .ZN(n4385) );
  NAND2_X1 U5133 ( .A1(n6150), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U5134 ( .A1(n5970), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5979) );
  AND2_X1 U5135 ( .A1(n5933), .A2(n5919), .ZN(n4386) );
  NAND2_X1 U5136 ( .A1(n6150), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5758) );
  INV_X1 U5137 ( .A(n5754), .ZN(n5752) );
  NAND2_X1 U5138 ( .A1(n5895), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n5910) );
  INV_X1 U5139 ( .A(n5847), .ZN(n4381) );
  INV_X1 U5140 ( .A(n5848), .ZN(n4379) );
  NAND2_X1 U5141 ( .A1(n4741), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U5142 ( .A1(n6150), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6001) );
  INV_X1 U5143 ( .A(n5640), .ZN(n6038) );
  AND4_X1 U5144 ( .A1(n5726), .A2(n5725), .A3(n5724), .A4(n5723), .ZN(n7262)
         );
  AND4_X1 U5145 ( .A1(n5678), .A2(n5677), .A3(n5676), .A4(n5675), .ZN(n7118)
         );
  NOR2_X1 U5146 ( .A1(n9449), .A2(n4286), .ZN(n6741) );
  OR2_X1 U5147 ( .A1(n6741), .A2(n6740), .ZN(n4419) );
  NOR2_X1 U5148 ( .A1(n6888), .A2(n4324), .ZN(n8246) );
  OR2_X1 U5149 ( .A1(n8246), .A2(n8247), .ZN(n4425) );
  OR2_X1 U5150 ( .A1(n8287), .A2(n8286), .ZN(n4423) );
  AND2_X1 U5151 ( .A1(n4423), .A2(n4422), .ZN(n8299) );
  NAND2_X1 U5152 ( .A1(n8284), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n4422) );
  OR2_X1 U5153 ( .A1(n8299), .A2(n8300), .ZN(n4421) );
  NAND2_X1 U5154 ( .A1(n6139), .A2(n6138), .ZN(n8628) );
  AND2_X1 U5155 ( .A1(n8422), .A2(n8421), .ZN(n6137) );
  NOR2_X1 U5156 ( .A1(n4758), .A2(n4757), .ZN(n4756) );
  INV_X1 U5157 ( .A(n7998), .ZN(n4757) );
  NAND2_X1 U5158 ( .A1(n4755), .A2(n4754), .ZN(n4753) );
  INV_X1 U5159 ( .A(n4758), .ZN(n4755) );
  INV_X1 U5160 ( .A(n8439), .ZN(n4754) );
  OR2_X1 U5161 ( .A1(n8646), .A2(n8472), .ZN(n7998) );
  NAND2_X1 U5162 ( .A1(n8454), .A2(n7997), .ZN(n8458) );
  NOR2_X1 U5163 ( .A1(n8650), .A2(n8656), .ZN(n4611) );
  AOI21_X1 U5164 ( .B1(n4774), .B2(n8479), .A(n4307), .ZN(n4772) );
  INV_X1 U5165 ( .A(n4774), .ZN(n4773) );
  NOR2_X1 U5166 ( .A1(n8469), .A2(n4775), .ZN(n4774) );
  INV_X1 U5167 ( .A(n4825), .ZN(n4775) );
  AND2_X1 U5168 ( .A1(n6264), .A2(n6266), .ZN(n8469) );
  NAND2_X1 U5169 ( .A1(n6135), .A2(n6134), .ZN(n8508) );
  AND2_X1 U5170 ( .A1(n8671), .A2(n8223), .ZN(n4377) );
  AND2_X1 U5171 ( .A1(n6130), .A2(n6251), .ZN(n4590) );
  INV_X1 U5172 ( .A(n8534), .ZN(n6130) );
  AND2_X1 U5173 ( .A1(n5944), .A2(n5943), .ZN(n8539) );
  OR2_X1 U5174 ( .A1(n8681), .A2(n8138), .ZN(n8554) );
  NAND2_X1 U5175 ( .A1(n8568), .A2(n8569), .ZN(n8567) );
  AND2_X1 U5176 ( .A1(n8554), .A2(n6242), .ZN(n8569) );
  OR2_X1 U5177 ( .A1(n8596), .A2(n8137), .ZN(n4824) );
  NAND2_X1 U5178 ( .A1(n8591), .A2(n4769), .ZN(n4771) );
  OR2_X1 U5179 ( .A1(n7594), .A2(n7598), .ZN(n4782) );
  NAND2_X1 U5180 ( .A1(n6150), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5844) );
  AND2_X1 U5181 ( .A1(n7989), .A2(n6121), .ZN(n7616) );
  INV_X1 U5182 ( .A(n6120), .ZN(n7598) );
  NAND2_X1 U5183 ( .A1(n5789), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5806) );
  INV_X1 U5184 ( .A(n5790), .ZN(n5789) );
  NOR2_X1 U5185 ( .A1(n7396), .A2(n4777), .ZN(n4776) );
  CLKBUF_X1 U5186 ( .A(n7356), .Z(n7256) );
  AND4_X1 U5187 ( .A1(n5706), .A2(n5705), .A3(n5704), .A4(n5703), .ZN(n8088)
         );
  AND4_X1 U5188 ( .A1(n5664), .A2(n5663), .A3(n5662), .A4(n5661), .ZN(n8157)
         );
  NAND2_X1 U5189 ( .A1(n6150), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U5190 ( .A1(n6871), .A2(n6300), .ZN(n4584) );
  INV_X1 U5191 ( .A(n8571), .ZN(n8536) );
  NAND2_X1 U5192 ( .A1(n6113), .A2(n9865), .ZN(n9827) );
  NAND2_X1 U5193 ( .A1(n6165), .A2(n6164), .ZN(n8618) );
  NAND2_X1 U5194 ( .A1(n5951), .A2(n5950), .ZN(n8661) );
  INV_X1 U5195 ( .A(n8524), .ZN(n8668) );
  INV_X1 U5196 ( .A(n8039), .ZN(n9893) );
  OAI22_X1 U5197 ( .A1(n5628), .A2(n6575), .B1(n6574), .B2(n6710), .ZN(n4567)
         );
  NAND3_X1 U5198 ( .A1(n4486), .A2(n4785), .A3(n4487), .ZN(n4788) );
  NOR2_X1 U5199 ( .A1(n4786), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4785) );
  INV_X1 U5200 ( .A(n4788), .ZN(n5581) );
  NOR2_X1 U5201 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n4742) );
  OR3_X1 U5202 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n5630) );
  AND2_X1 U5203 ( .A1(n7568), .A2(n7580), .ZN(n4392) );
  NAND2_X1 U5204 ( .A1(n5304), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5324) );
  INV_X1 U5205 ( .A(n5305), .ZN(n5304) );
  INV_X1 U5206 ( .A(n8866), .ZN(n7292) );
  OR2_X1 U5207 ( .A1(n6568), .A2(n5587), .ZN(n4501) );
  NAND2_X1 U5208 ( .A1(n4410), .A2(n4409), .ZN(n8734) );
  OAI21_X1 U5209 ( .B1(n6476), .B2(n4408), .A(n4406), .ZN(n4410) );
  NOR2_X1 U5210 ( .A1(n4411), .A2(n6481), .ZN(n4405) );
  NAND2_X1 U5211 ( .A1(n4398), .A2(n4397), .ZN(n7546) );
  NAND2_X1 U5212 ( .A1(n4400), .A2(n4399), .ZN(n4398) );
  INV_X1 U5213 ( .A(n7424), .ZN(n4400) );
  NAND2_X1 U5214 ( .A1(n4791), .A2(n6460), .ZN(n8753) );
  NOR2_X1 U5215 ( .A1(n7349), .A2(n4805), .ZN(n4804) );
  INV_X1 U5216 ( .A(n4807), .ZN(n4805) );
  NAND2_X1 U5217 ( .A1(n6464), .A2(n4391), .ZN(n4390) );
  INV_X1 U5218 ( .A(n4789), .ZN(n4389) );
  OR2_X1 U5219 ( .A1(n9582), .A2(n9581), .ZN(n4513) );
  NAND2_X1 U5220 ( .A1(n4513), .A2(n4512), .ZN(n4511) );
  NAND2_X1 U5221 ( .A1(n9592), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4512) );
  AND2_X1 U5222 ( .A1(n4511), .A2(n4510), .ZN(n9423) );
  INV_X1 U5223 ( .A(n9424), .ZN(n4510) );
  OAI22_X1 U5224 ( .A1(n6987), .A2(n6986), .B1(P1_REG1_REG_7__SCAN_IN), .B2(
        n6996), .ZN(n8872) );
  OAI21_X1 U5225 ( .B1(n6997), .B2(n6998), .A(n4514), .ZN(n8878) );
  OR2_X1 U5226 ( .A1(n6996), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U5227 ( .A1(n9616), .A2(n4517), .ZN(n9629) );
  AND2_X1 U5228 ( .A1(n9620), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4517) );
  NOR2_X1 U5229 ( .A1(n9628), .A2(n9629), .ZN(n9627) );
  AOI21_X1 U5230 ( .B1(n8939), .B2(P1_REG1_REG_17__SCAN_IN), .A(n8930), .ZN(
        n8931) );
  OR3_X1 U5231 ( .A1(n5417), .A2(n5416), .A3(n8022), .ZN(n5539) );
  NAND2_X1 U5232 ( .A1(n9003), .A2(n7924), .ZN(n8976) );
  NOR2_X1 U5233 ( .A1(n9196), .A2(n9033), .ZN(n9010) );
  OR2_X1 U5234 ( .A1(n7786), .A2(n7785), .ZN(n9008) );
  INV_X1 U5235 ( .A(n8856), .ZN(n9031) );
  AND2_X1 U5236 ( .A1(n9017), .A2(n9016), .ZN(n9028) );
  NAND2_X1 U5237 ( .A1(n7747), .A2(n9015), .ZN(n9042) );
  NAND2_X1 U5238 ( .A1(n4542), .A2(n7906), .ZN(n9070) );
  NAND2_X1 U5239 ( .A1(n9094), .A2(n7903), .ZN(n4542) );
  INV_X1 U5240 ( .A(n4718), .ZN(n4717) );
  AOI21_X1 U5241 ( .B1(n4718), .B2(n4720), .A(n4716), .ZN(n4715) );
  INV_X1 U5242 ( .A(n9087), .ZN(n4716) );
  OR2_X1 U5243 ( .A1(n7941), .A2(n7957), .ZN(n9247) );
  INV_X1 U5244 ( .A(n9112), .ZN(n4723) );
  CLKBUF_X1 U5245 ( .A(n9110), .Z(n9112) );
  NAND2_X1 U5246 ( .A1(n9150), .A2(n7892), .ZN(n9135) );
  NAND2_X1 U5247 ( .A1(n9135), .A2(n9136), .ZN(n9134) );
  AND2_X1 U5248 ( .A1(n9144), .A2(n9133), .ZN(n9128) );
  NAND2_X1 U5249 ( .A1(n7651), .A2(n5518), .ZN(n9160) );
  NOR2_X1 U5250 ( .A1(n5507), .A2(n4694), .ZN(n4693) );
  INV_X1 U5251 ( .A(n5506), .ZN(n4694) );
  NAND2_X1 U5252 ( .A1(n4695), .A2(n4291), .ZN(n4691) );
  NAND2_X1 U5253 ( .A1(n7203), .A2(n7766), .ZN(n7192) );
  OR2_X1 U5254 ( .A1(n9688), .A2(n6375), .ZN(n9689) );
  INV_X1 U5255 ( .A(n6570), .ZN(n4671) );
  AOI21_X2 U5256 ( .B1(n4444), .B2(n7723), .A(n4443), .ZN(n9695) );
  INV_X1 U5257 ( .A(n7726), .ZN(n4443) );
  NAND2_X1 U5258 ( .A1(n7222), .A2(n9724), .ZN(n9688) );
  NOR2_X1 U5259 ( .A1(n6851), .A2(n7080), .ZN(n7222) );
  INV_X1 U5260 ( .A(n9698), .ZN(n9152) );
  NAND2_X1 U5261 ( .A1(n5360), .A2(n5359), .ZN(n9203) );
  NAND2_X1 U5262 ( .A1(n5274), .A2(n5273), .ZN(n9226) );
  XNOR2_X1 U5263 ( .A(n6157), .B(n6156), .ZN(n6160) );
  NAND2_X1 U5264 ( .A1(n4865), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4861) );
  XNOR2_X1 U5265 ( .A(n5291), .B(n5292), .ZN(n7335) );
  OAI21_X1 U5266 ( .B1(n5137), .B2(n4655), .A(n4653), .ZN(n5204) );
  NAND2_X1 U5267 ( .A1(n4652), .A2(n5157), .ZN(n5183) );
  XNOR2_X1 U5268 ( .A(n5007), .B(n5005), .ZN(n4361) );
  INV_X1 U5269 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4831) );
  OR2_X1 U5270 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4910) );
  NAND2_X1 U5271 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4521) );
  NAND2_X1 U5272 ( .A1(n6023), .A2(n6022), .ZN(n8636) );
  NAND2_X1 U5273 ( .A1(n7648), .A2(n5713), .ZN(n6023) );
  AND4_X1 U5274 ( .A1(n5811), .A2(n5810), .A3(n5809), .A4(n5808), .ZN(n7619)
         );
  INV_X1 U5275 ( .A(n9818), .ZN(n6115) );
  NAND2_X1 U5276 ( .A1(n5908), .A2(n5907), .ZN(n8677) );
  NAND2_X1 U5277 ( .A1(n4346), .A2(n8118), .ZN(n4345) );
  NAND2_X1 U5278 ( .A1(n5734), .A2(n5733), .ZN(n7354) );
  AND2_X1 U5279 ( .A1(n5673), .A2(n5657), .ZN(n4743) );
  INV_X1 U5280 ( .A(n6956), .ZN(n5673) );
  NAND2_X1 U5281 ( .A1(n6091), .A2(n6082), .ZN(n8216) );
  INV_X1 U5282 ( .A(n8190), .ZN(n8214) );
  NAND2_X1 U5283 ( .A1(n6171), .A2(n6810), .ZN(n4358) );
  NAND2_X1 U5284 ( .A1(n6322), .A2(n6321), .ZN(n6323) );
  NAND2_X1 U5285 ( .A1(n4490), .A2(n4489), .ZN(n4488) );
  NAND2_X1 U5286 ( .A1(n6030), .A2(n6029), .ZN(n8219) );
  NOR2_X1 U5287 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4557) );
  AND2_X1 U5288 ( .A1(n6532), .A2(n8829), .ZN(n4816) );
  NAND2_X1 U5289 ( .A1(n5257), .A2(n5256), .ZN(n9232) );
  NAND2_X1 U5290 ( .A1(n7009), .A2(n7011), .ZN(n7010) );
  NAND2_X1 U5291 ( .A1(n5338), .A2(n5337), .ZN(n9206) );
  NAND2_X1 U5292 ( .A1(n5368), .A2(n5367), .ZN(n9054) );
  NAND2_X1 U5293 ( .A1(n5347), .A2(n5346), .ZN(n9072) );
  OR2_X1 U5294 ( .A1(n9046), .A2(n5231), .ZN(n5347) );
  NAND2_X1 U5295 ( .A1(n5331), .A2(n5330), .ZN(n9088) );
  AND2_X1 U5296 ( .A1(n4915), .A2(n4914), .ZN(n4917) );
  OR2_X1 U5297 ( .A1(n5231), .A2(n7207), .ZN(n4918) );
  NAND2_X1 U5298 ( .A1(n4934), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4882) );
  OR2_X1 U5299 ( .A1(n4940), .A2(n4878), .ZN(n4883) );
  OR2_X1 U5300 ( .A1(n5236), .A2(n4879), .ZN(n4881) );
  NOR2_X1 U5301 ( .A1(n8938), .A2(n4520), .ZN(n8940) );
  AND2_X1 U5302 ( .A1(n8939), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4520) );
  NAND2_X1 U5303 ( .A1(n8953), .A2(n8952), .ZN(n4372) );
  INV_X1 U5304 ( .A(n8956), .ZN(n4373) );
  NAND2_X1 U5305 ( .A1(n7678), .A2(n7677), .ZN(n9177) );
  NAND2_X1 U5306 ( .A1(n9684), .A2(n6546), .ZN(n9710) );
  AND2_X1 U5307 ( .A1(n9684), .A2(n5538), .ZN(n9692) );
  INV_X1 U5308 ( .A(n4352), .ZN(n4351) );
  NAND2_X1 U5309 ( .A1(n9180), .A2(n9244), .ZN(n4497) );
  INV_X1 U5310 ( .A(n5254), .ZN(n7953) );
  INV_X2 U5311 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8959) );
  NAND2_X1 U5312 ( .A1(n4478), .A2(n4477), .ZN(n6191) );
  OAI211_X1 U5313 ( .C1(n6220), .C2(n6288), .A(n4460), .B(n7598), .ZN(n4459)
         );
  OAI21_X1 U5314 ( .B1(n6216), .B2(n6215), .A(n4461), .ZN(n4460) );
  NAND2_X1 U5315 ( .A1(n4458), .A2(n4457), .ZN(n4456) );
  INV_X1 U5316 ( .A(n8597), .ZN(n4457) );
  INV_X1 U5317 ( .A(n6231), .ZN(n4458) );
  NAND2_X1 U5318 ( .A1(n4448), .A2(n7851), .ZN(n7852) );
  NAND2_X1 U5319 ( .A1(n4451), .A2(n4449), .ZN(n4448) );
  AND2_X1 U5320 ( .A1(n6249), .A2(n6288), .ZN(n4483) );
  OAI21_X1 U5321 ( .B1(n6244), .B2(n6243), .A(n4298), .ZN(n6246) );
  NAND2_X1 U5322 ( .A1(n4445), .A2(n7878), .ZN(n7890) );
  NAND2_X1 U5323 ( .A1(n4368), .A2(n6279), .ZN(n4367) );
  NAND2_X1 U5324 ( .A1(n8636), .A2(n8406), .ZN(n4368) );
  NOR2_X1 U5325 ( .A1(n6265), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U5326 ( .A1(n4480), .A2(n4293), .ZN(n4479) );
  NOR2_X1 U5327 ( .A1(n8455), .A2(n4662), .ZN(n4661) );
  NOR2_X1 U5328 ( .A1(n6266), .A2(n6279), .ZN(n4662) );
  AOI21_X1 U5329 ( .B1(n4476), .B2(n6275), .A(n4306), .ZN(n4466) );
  NOR2_X1 U5330 ( .A1(n8630), .A2(n6288), .ZN(n4474) );
  INV_X1 U5331 ( .A(n4476), .ZN(n4467) );
  NAND2_X1 U5332 ( .A1(n4468), .A2(n4270), .ZN(n4463) );
  OAI21_X1 U5333 ( .B1(n4469), .B2(n4476), .A(n4475), .ZN(n4468) );
  NAND2_X1 U5334 ( .A1(n4335), .A2(n6444), .ZN(n4812) );
  NAND2_X1 U5335 ( .A1(n4453), .A2(n7905), .ZN(n4452) );
  NAND2_X1 U5336 ( .A1(n4294), .A2(n4473), .ZN(n4472) );
  INV_X1 U5337 ( .A(n6176), .ZN(n4571) );
  INV_X1 U5338 ( .A(n4812), .ZN(n4395) );
  OAI21_X1 U5339 ( .B1(n7547), .B2(n4812), .A(n7570), .ZN(n4811) );
  OR2_X1 U5340 ( .A1(n9211), .A2(n8796), .ZN(n7690) );
  NAND2_X1 U5341 ( .A1(n4702), .A2(n4705), .ZN(n4700) );
  NOR2_X1 U5342 ( .A1(n4703), .A2(n5515), .ZN(n4701) );
  INV_X1 U5343 ( .A(n4626), .ZN(n4625) );
  OAI21_X1 U5344 ( .B1(n5410), .B2(n4627), .A(n5429), .ZN(n4626) );
  INV_X1 U5345 ( .A(n5412), .ZN(n4627) );
  NAND2_X1 U5346 ( .A1(n4846), .A2(n4821), .ZN(n4820) );
  INV_X1 U5347 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4821) );
  INV_X1 U5348 ( .A(n5393), .ZN(n4634) );
  INV_X1 U5349 ( .A(n5203), .ZN(n4651) );
  NAND2_X1 U5350 ( .A1(n5161), .A2(n5160), .ZN(n5181) );
  NOR2_X1 U5351 ( .A1(n4618), .A2(n4615), .ZN(n4614) );
  INV_X1 U5352 ( .A(n5051), .ZN(n4615) );
  INV_X1 U5353 ( .A(n4619), .ZN(n4618) );
  NOR2_X1 U5354 ( .A1(n5092), .A2(n4620), .ZN(n4619) );
  INV_X1 U5355 ( .A(n5075), .ZN(n4620) );
  INV_X1 U5356 ( .A(n5090), .ZN(n5092) );
  INV_X1 U5357 ( .A(n4822), .ZN(n4617) );
  NAND2_X1 U5358 ( .A1(n5095), .A2(n5094), .ZN(n5112) );
  INV_X1 U5359 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5057) );
  INV_X1 U5360 ( .A(n4728), .ZN(n4727) );
  OAI21_X1 U5361 ( .B1(n4271), .B2(n4729), .A(n8043), .ZN(n4728) );
  NAND2_X1 U5362 ( .A1(n6150), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5725) );
  NOR2_X1 U5363 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5715) );
  INV_X1 U5364 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5781) );
  OR2_X1 U5365 ( .A1(n8656), .A2(n8506), .ZN(n6263) );
  NAND2_X1 U5366 ( .A1(n8553), .A2(n4603), .ZN(n4602) );
  NAND2_X1 U5367 ( .A1(n5838), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5860) );
  OR2_X1 U5368 ( .A1(n5823), .A2(n5822), .ZN(n5840) );
  OR2_X1 U5369 ( .A1(n5806), .A2(n7282), .ZN(n5823) );
  INV_X1 U5370 ( .A(n7355), .ZN(n4777) );
  AND2_X1 U5371 ( .A1(n4599), .A2(n4595), .ZN(n8611) );
  NOR2_X1 U5372 ( .A1(n7614), .A2(n7620), .ZN(n4595) );
  INV_X1 U5373 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5552) );
  NOR2_X1 U5374 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5547) );
  NOR2_X1 U5375 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5548) );
  INV_X1 U5376 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5782) );
  OR2_X1 U5377 ( .A1(n5732), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5785) );
  AND2_X1 U5378 ( .A1(n5551), .A2(n5589), .ZN(n5647) );
  INV_X1 U5379 ( .A(n8784), .ZN(n4411) );
  NAND2_X1 U5380 ( .A1(n7455), .A2(n4403), .ZN(n4396) );
  NAND2_X1 U5381 ( .A1(n4404), .A2(n6431), .ZN(n4403) );
  INV_X1 U5382 ( .A(n6430), .ZN(n4404) );
  INV_X1 U5383 ( .A(n6420), .ZN(n4809) );
  NAND2_X1 U5384 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  INV_X1 U5385 ( .A(n8841), .ZN(n4391) );
  AND2_X1 U5386 ( .A1(n9177), .A2(n7756), .ZN(n7933) );
  NAND2_X1 U5387 ( .A1(n4642), .A2(n4336), .ZN(n7796) );
  OAI21_X1 U5388 ( .B1(n7814), .B2(n7749), .A(n7812), .ZN(n7750) );
  AND2_X1 U5389 ( .A1(n5139), .A2(n5138), .ZN(n5190) );
  INV_X1 U5390 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5138) );
  AND2_X1 U5391 ( .A1(n8892), .A2(n4522), .ZN(n7518) );
  NAND2_X1 U5392 ( .A1(n8887), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5393 ( .A1(n7979), .A2(n7684), .ZN(n4642) );
  OR2_X1 U5394 ( .A1(n9180), .A2(n7938), .ZN(n7753) );
  NOR2_X1 U5395 ( .A1(n9060), .A2(n4538), .ZN(n4537) );
  INV_X1 U5396 ( .A(n7903), .ZN(n4538) );
  INV_X1 U5397 ( .A(n7690), .ZN(n4540) );
  NAND2_X1 U5398 ( .A1(n9049), .A2(n4508), .ZN(n4507) );
  OR2_X1 U5399 ( .A1(n9206), .A2(n9032), .ZN(n7747) );
  NAND2_X1 U5400 ( .A1(n9206), .A2(n9032), .ZN(n9015) );
  AND2_X1 U5401 ( .A1(n7907), .A2(n9085), .ZN(n7903) );
  NOR2_X1 U5402 ( .A1(n9211), .A2(n9216), .ZN(n4508) );
  NAND2_X1 U5403 ( .A1(n4685), .A2(n7881), .ZN(n4684) );
  INV_X1 U5404 ( .A(n5519), .ZN(n4685) );
  NOR2_X1 U5405 ( .A1(n4686), .A2(n4681), .ZN(n4680) );
  INV_X1 U5406 ( .A(n5518), .ZN(n4681) );
  OR2_X1 U5407 ( .A1(n8762), .A2(n9165), .ZN(n7877) );
  NAND2_X1 U5408 ( .A1(n5170), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5195) );
  INV_X1 U5409 ( .A(n5172), .ZN(n5170) );
  NOR2_X1 U5410 ( .A1(n8851), .A2(n7673), .ZN(n4499) );
  OAI21_X1 U5411 ( .B1(n9494), .B2(n4535), .A(n4532), .ZN(n7632) );
  AOI21_X1 U5412 ( .B1(n5153), .B2(n4534), .A(n4533), .ZN(n4532) );
  INV_X1 U5413 ( .A(n7865), .ZN(n4533) );
  NAND2_X1 U5414 ( .A1(n4360), .A2(n7631), .ZN(n7630) );
  OR2_X1 U5415 ( .A1(n5126), .A2(n5125), .ZN(n5146) );
  NAND2_X1 U5416 ( .A1(n5103), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5126) );
  INV_X1 U5417 ( .A(n5105), .ZN(n5103) );
  NAND2_X1 U5418 ( .A1(n4687), .A2(n4689), .ZN(n9505) );
  AOI21_X1 U5419 ( .B1(n7845), .B2(n4690), .A(n4297), .ZN(n4689) );
  NAND2_X1 U5420 ( .A1(n5064), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5082) );
  NAND2_X1 U5421 ( .A1(n5019), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5042) );
  INV_X1 U5422 ( .A(n5020), .ZN(n5019) );
  INV_X1 U5423 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5041) );
  OR2_X1 U5424 ( .A1(n5042), .A2(n5041), .ZN(n5065) );
  NAND2_X1 U5425 ( .A1(n4554), .A2(n7728), .ZN(n7829) );
  INV_X1 U5426 ( .A(n8870), .ZN(n5496) );
  NOR2_X1 U5427 ( .A1(n4820), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n4819) );
  INV_X1 U5428 ( .A(n4820), .ZN(n4818) );
  INV_X1 U5429 ( .A(n5351), .ZN(n4638) );
  INV_X1 U5430 ( .A(n4637), .ZN(n4636) );
  OAI21_X1 U5431 ( .B1(n4640), .B2(n4322), .A(n5369), .ZN(n4637) );
  NAND2_X1 U5432 ( .A1(n4284), .A2(n5448), .ZN(n4710) );
  NAND2_X1 U5433 ( .A1(n4643), .A2(n4325), .ZN(n5296) );
  AOI21_X1 U5434 ( .B1(n4646), .B2(n4645), .A(n4330), .ZN(n4644) );
  INV_X1 U5435 ( .A(n5225), .ZN(n4645) );
  NAND2_X1 U5436 ( .A1(n4656), .A2(n5157), .ZN(n4655) );
  INV_X1 U5437 ( .A(n5182), .ZN(n4656) );
  INV_X1 U5438 ( .A(n4654), .ZN(n4653) );
  OAI21_X1 U5439 ( .B1(n4657), .B2(n4655), .A(n5181), .ZN(n4654) );
  NOR2_X1 U5440 ( .A1(n5158), .A2(n4658), .ZN(n4657) );
  INV_X1 U5441 ( .A(n5136), .ZN(n4658) );
  INV_X1 U5442 ( .A(n5154), .ZN(n5158) );
  XNOR2_X1 U5443 ( .A(n5155), .B(SI_14_), .ZN(n5154) );
  OAI21_X2 U5444 ( .B1(n5114), .B2(n5113), .A(n5112), .ZN(n5135) );
  AND2_X1 U5445 ( .A1(n5136), .A2(n5119), .ZN(n5134) );
  NAND2_X1 U5446 ( .A1(n5028), .A2(n5014), .ZN(n5029) );
  XNOR2_X1 U5447 ( .A(n4984), .B(SI_6_), .ZN(n4981) );
  INV_X1 U5448 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4925) );
  OAI21_X1 U5449 ( .B1(n5184), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n4370), .ZN(
        n4906) );
  NAND2_X1 U5450 ( .A1(n5184), .A2(n4874), .ZN(n4370) );
  OR2_X1 U5451 ( .A1(n5979), .A2(n8151), .ZN(n5998) );
  INV_X1 U5452 ( .A(n5987), .ZN(n5988) );
  NAND2_X1 U5453 ( .A1(n7234), .A2(n5742), .ZN(n7231) );
  NAND2_X1 U5454 ( .A1(n8074), .A2(n5915), .ZN(n8079) );
  INV_X1 U5455 ( .A(n5954), .ZN(n5952) );
  INV_X1 U5456 ( .A(n5742), .ZN(n4739) );
  INV_X1 U5457 ( .A(n7232), .ZN(n4740) );
  INV_X1 U5458 ( .A(n5764), .ZN(n4736) );
  AND2_X1 U5459 ( .A1(n6827), .A2(n5605), .ZN(n6767) );
  AND2_X1 U5460 ( .A1(n8136), .A2(n5871), .ZN(n4380) );
  AOI21_X1 U5461 ( .B1(n4579), .B2(n4583), .A(n4575), .ZN(n4574) );
  AND2_X1 U5462 ( .A1(n4577), .A2(n6277), .ZN(n4575) );
  CLKBUF_X1 U5463 ( .A(n5603), .Z(n6171) );
  NOR2_X1 U5464 ( .A1(n9866), .A2(n6289), .ZN(n4489) );
  NAND2_X1 U5465 ( .A1(n4491), .A2(n7309), .ZN(n6321) );
  NAND2_X1 U5466 ( .A1(n4493), .A2(n6279), .ZN(n4492) );
  NAND2_X1 U5467 ( .A1(n4363), .A2(n4288), .ZN(n6286) );
  OR2_X1 U5468 ( .A1(n8398), .A2(n6038), .ZN(n6044) );
  AND3_X1 U5469 ( .A1(n5928), .A2(n5927), .A3(n5926), .ZN(n8101) );
  NAND2_X1 U5470 ( .A1(n6150), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5826) );
  NAND2_X1 U5471 ( .A1(n5621), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5567) );
  AND2_X1 U5472 ( .A1(n4425), .A2(n4424), .ZN(n8260) );
  NAND2_X1 U5473 ( .A1(n8244), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n4424) );
  NOR2_X1 U5474 ( .A1(n8260), .A2(n8261), .ZN(n8259) );
  NOR2_X1 U5475 ( .A1(n6973), .A2(n4427), .ZN(n6975) );
  AND2_X1 U5476 ( .A1(n6974), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U5477 ( .A1(n6976), .A2(n6975), .ZN(n7140) );
  NOR2_X1 U5478 ( .A1(n7140), .A2(n4426), .ZN(n7144) );
  AND2_X1 U5479 ( .A1(n7141), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4426) );
  NAND2_X1 U5480 ( .A1(n7144), .A2(n7143), .ZN(n7278) );
  NAND2_X1 U5481 ( .A1(n4433), .A2(n4431), .ZN(n8313) );
  NOR2_X1 U5482 ( .A1(n4435), .A2(n8326), .ZN(n4434) );
  NAND2_X1 U5483 ( .A1(n7381), .A2(n9472), .ZN(n4435) );
  NOR2_X1 U5484 ( .A1(n8351), .A2(n4343), .ZN(n8353) );
  NAND2_X1 U5485 ( .A1(n8353), .A2(n8352), .ZN(n8370) );
  NOR2_X1 U5486 ( .A1(n8396), .A2(n8628), .ZN(n8388) );
  OR3_X1 U5487 ( .A1(n6036), .A2(n8046), .A3(n6104), .ZN(n6094) );
  INV_X1 U5488 ( .A(n7999), .ZN(n4745) );
  OR2_X1 U5489 ( .A1(n8630), .A2(n8414), .ZN(n8396) );
  AOI21_X1 U5490 ( .B1(n4750), .B2(n4748), .A(n4302), .ZN(n4747) );
  INV_X1 U5491 ( .A(n4756), .ZN(n4748) );
  OR2_X1 U5492 ( .A1(n8636), .A2(n8430), .ZN(n8414) );
  NAND2_X1 U5493 ( .A1(n8498), .A2(n4608), .ZN(n8430) );
  AND2_X1 U5494 ( .A1(n4609), .A2(n8434), .ZN(n4608) );
  NAND2_X1 U5495 ( .A1(n6270), .A2(n8421), .ZN(n8439) );
  NAND2_X1 U5496 ( .A1(n4587), .A2(n4586), .ZN(n8470) );
  NAND2_X1 U5497 ( .A1(n4589), .A2(n6250), .ZN(n4586) );
  NAND2_X1 U5498 ( .A1(n8498), .A2(n8491), .ZN(n8485) );
  NAND2_X1 U5499 ( .A1(n6259), .A2(n6245), .ZN(n8504) );
  NAND2_X1 U5500 ( .A1(n5922), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5937) );
  INV_X1 U5501 ( .A(n5924), .ZN(n5922) );
  OR2_X1 U5502 ( .A1(n5937), .A2(n8107), .ZN(n5954) );
  NAND2_X1 U5503 ( .A1(n4600), .A2(n4601), .ZN(n8547) );
  NOR2_X1 U5504 ( .A1(n8681), .A2(n4602), .ZN(n4601) );
  INV_X1 U5505 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5506 ( .B1(n8569), .B2(n7992), .A(n4766), .ZN(n4765) );
  OAI21_X1 U5507 ( .B1(n8585), .B2(n6126), .A(n6236), .ZN(n8568) );
  NOR3_X1 U5508 ( .A1(n8593), .A2(n8687), .A3(n8681), .ZN(n8563) );
  NOR2_X1 U5509 ( .A1(n7614), .A2(n4597), .ZN(n4596) );
  NAND2_X1 U5510 ( .A1(n9467), .A2(n9463), .ZN(n4597) );
  INV_X1 U5511 ( .A(n6224), .ZN(n8608) );
  AOI21_X1 U5512 ( .B1(n4781), .B2(n7598), .A(n4780), .ZN(n4779) );
  INV_X1 U5513 ( .A(n7989), .ZN(n4780) );
  AND2_X1 U5514 ( .A1(n6307), .A2(n6306), .ZN(n9804) );
  AOI21_X1 U5515 ( .B1(n4564), .B2(n4566), .A(n4562), .ZN(n4561) );
  INV_X1 U5516 ( .A(n4565), .ZN(n4564) );
  AND2_X1 U5517 ( .A1(n7365), .A2(n9910), .ZN(n7405) );
  NAND2_X1 U5518 ( .A1(n7261), .A2(n6304), .ZN(n4563) );
  NOR2_X1 U5519 ( .A1(n7267), .A2(n7354), .ZN(n7365) );
  NOR2_X1 U5520 ( .A1(n7251), .A2(n4761), .ZN(n4760) );
  NAND2_X1 U5521 ( .A1(n4607), .A2(n4606), .ZN(n7267) );
  INV_X1 U5522 ( .A(n7177), .ZN(n4607) );
  NAND2_X1 U5523 ( .A1(n7113), .A2(n9893), .ZN(n7177) );
  NOR2_X1 U5524 ( .A1(n7047), .A2(n9883), .ZN(n7113) );
  NAND2_X1 U5525 ( .A1(n4585), .A2(n4584), .ZN(n7025) );
  AND2_X1 U5526 ( .A1(n6299), .A2(n6175), .ZN(n4585) );
  NOR2_X1 U5527 ( .A1(n9843), .A2(n6807), .ZN(n6874) );
  AND2_X1 U5528 ( .A1(n9851), .A2(n6762), .ZN(n7048) );
  AOI211_X1 U5529 ( .C1(n8396), .C2(n8628), .A(n8388), .B(n9921), .ZN(n8627)
         );
  OR2_X1 U5530 ( .A1(n8629), .A2(n9888), .ZN(n4592) );
  NAND2_X1 U5531 ( .A1(n5921), .A2(n5920), .ZN(n8671) );
  AND2_X1 U5532 ( .A1(n9866), .A2(n6328), .ZN(n9927) );
  NAND2_X1 U5533 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n4559) );
  INV_X1 U5534 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U5535 ( .A1(n5572), .A2(n5571), .ZN(n5576) );
  NAND2_X1 U5536 ( .A1(n4667), .A2(n4666), .ZN(n5601) );
  AND2_X1 U5537 ( .A1(n4867), .A2(n4868), .ZN(n4666) );
  NAND2_X1 U5538 ( .A1(n5232), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5259) );
  INV_X1 U5539 ( .A(n5233), .ZN(n5232) );
  NAND2_X1 U5540 ( .A1(n5194), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5213) );
  INV_X1 U5541 ( .A(n5195), .ZN(n5194) );
  NAND2_X1 U5542 ( .A1(n5323), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U5543 ( .A1(n4794), .A2(n4793), .ZN(n4792) );
  NAND2_X1 U5544 ( .A1(n4795), .A2(n8726), .ZN(n4793) );
  XNOR2_X1 U5545 ( .A(n6383), .B(n6362), .ZN(n6389) );
  NAND2_X1 U5546 ( .A1(n6382), .A2(n6381), .ZN(n6383) );
  NAND2_X1 U5547 ( .A1(n8869), .A2(n4244), .ZN(n6382) );
  OR2_X1 U5548 ( .A1(n7290), .A2(n4809), .ZN(n4807) );
  NAND2_X1 U5549 ( .A1(n6421), .A2(n4808), .ZN(n4806) );
  AND2_X1 U5550 ( .A1(n4417), .A2(n8801), .ZN(n4414) );
  AND2_X1 U5551 ( .A1(n4303), .A2(n4417), .ZN(n4408) );
  OR2_X1 U5552 ( .A1(n7426), .A2(n7425), .ZN(n6430) );
  NAND2_X1 U5553 ( .A1(n4803), .A2(n4283), .ZN(n4802) );
  INV_X1 U5554 ( .A(n4804), .ZN(n4803) );
  NAND2_X1 U5555 ( .A1(n4936), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n4998) );
  OR2_X1 U5556 ( .A1(n9177), .A2(n7756), .ZN(n7955) );
  XNOR2_X1 U5557 ( .A(n6639), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n9570) );
  AOI21_X1 U5558 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6642), .A(n9420), .ZN(
        n9602) );
  NAND2_X1 U5559 ( .A1(n4516), .A2(n4515), .ZN(n6997) );
  NAND2_X1 U5560 ( .A1(n6671), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4515) );
  INV_X1 U5561 ( .A(n6670), .ZN(n4516) );
  NAND2_X1 U5562 ( .A1(n8878), .A2(n8877), .ZN(n8876) );
  AOI21_X1 U5563 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n8880), .A(n8871), .ZN(
        n9612) );
  NOR2_X1 U5564 ( .A1(n9627), .A2(n4327), .ZN(n9645) );
  NAND2_X1 U5565 ( .A1(n9645), .A2(n9646), .ZN(n9644) );
  XNOR2_X1 U5566 ( .A(n7518), .B(n9653), .ZN(n9656) );
  NAND2_X1 U5567 ( .A1(n9656), .A2(n7539), .ZN(n9655) );
  XNOR2_X1 U5568 ( .A(n4518), .B(n8947), .ZN(n8955) );
  OR2_X1 U5569 ( .A1(n8946), .A2(n4519), .ZN(n4518) );
  AND2_X1 U5570 ( .A1(n8950), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4519) );
  NAND2_X1 U5571 ( .A1(n4642), .A2(n7685), .ZN(n8967) );
  INV_X1 U5572 ( .A(n8975), .ZN(n8972) );
  INV_X1 U5573 ( .A(n7924), .ZN(n4553) );
  OR2_X1 U5574 ( .A1(n8986), .A2(n5231), .ZN(n5427) );
  INV_X1 U5575 ( .A(n9008), .ZN(n9019) );
  NAND2_X1 U5576 ( .A1(n9021), .A2(n9152), .ZN(n4355) );
  OR2_X1 U5577 ( .A1(n5361), .A2(n8746), .ZN(n5381) );
  OR2_X1 U5578 ( .A1(n5340), .A2(n5339), .ZN(n5361) );
  INV_X1 U5579 ( .A(n9072), .ZN(n9032) );
  NOR2_X1 U5580 ( .A1(n9101), .A2(n4506), .ZN(n9062) );
  INV_X1 U5581 ( .A(n4508), .ZN(n4506) );
  NOR2_X1 U5582 ( .A1(n9101), .A2(n9216), .ZN(n9080) );
  NAND2_X1 U5583 ( .A1(n5275), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5287) );
  INV_X1 U5584 ( .A(n5277), .ZN(n5275) );
  OR2_X1 U5585 ( .A1(n5287), .A2(n8737), .ZN(n5305) );
  AOI21_X1 U5586 ( .B1(n4549), .B2(n9127), .A(n4547), .ZN(n4546) );
  NOR2_X1 U5587 ( .A1(n4548), .A2(n4545), .ZN(n4544) );
  AOI21_X1 U5588 ( .B1(n9162), .B2(n9161), .A(n4344), .ZN(n9151) );
  INV_X1 U5589 ( .A(n7692), .ZN(n4344) );
  NAND2_X1 U5590 ( .A1(n9488), .A2(n4272), .ZN(n9169) );
  AND2_X1 U5591 ( .A1(n9488), .A2(n4499), .ZN(n7657) );
  AND2_X1 U5592 ( .A1(n9488), .A2(n9536), .ZN(n7642) );
  NAND2_X1 U5593 ( .A1(n9492), .A2(n5153), .ZN(n7532) );
  OAI21_X1 U5594 ( .B1(n7498), .B2(n7712), .A(n7860), .ZN(n9494) );
  NAND2_X1 U5595 ( .A1(n9494), .A2(n9493), .ZN(n9492) );
  AND2_X1 U5596 ( .A1(n7855), .A2(n7860), .ZN(n7774) );
  INV_X1 U5597 ( .A(n8861), .ZN(n9511) );
  NAND2_X1 U5598 ( .A1(n5049), .A2(n7837), .ZN(n7298) );
  AOI21_X1 U5599 ( .B1(n4526), .B2(n4527), .A(n4525), .ZN(n4524) );
  NAND2_X1 U5600 ( .A1(n7159), .A2(n5506), .ZN(n9668) );
  NAND2_X1 U5601 ( .A1(n4528), .A2(n7830), .ZN(n7841) );
  NAND2_X1 U5602 ( .A1(n4442), .A2(n4441), .ZN(n4528) );
  AND2_X1 U5603 ( .A1(n7828), .A2(n7833), .ZN(n4441) );
  NAND2_X1 U5604 ( .A1(n4676), .A2(n4675), .ZN(n7160) );
  AOI21_X1 U5605 ( .B1(n7131), .B2(n4678), .A(n4301), .ZN(n4675) );
  NAND2_X1 U5606 ( .A1(n5502), .A2(n4677), .ZN(n4676) );
  AND2_X1 U5607 ( .A1(n4442), .A2(n7828), .ZN(n7122) );
  OR3_X1 U5608 ( .A1(n6785), .A2(n6781), .A3(n6534), .ZN(n6935) );
  NAND2_X1 U5609 ( .A1(n9181), .A2(n9526), .ZN(n4376) );
  NAND2_X1 U5610 ( .A1(n5403), .A2(n5402), .ZN(n9191) );
  NAND2_X1 U5611 ( .A1(n5378), .A2(n5377), .ZN(n9196) );
  NAND2_X1 U5612 ( .A1(n7579), .A2(n7684), .ZN(n5378) );
  INV_X1 U5613 ( .A(n9759), .ZN(n9244) );
  XNOR2_X1 U5614 ( .A(n6160), .B(SI_30_), .ZN(n7979) );
  XNOR2_X1 U5615 ( .A(n6142), .B(n5434), .ZN(n8717) );
  NAND2_X1 U5616 ( .A1(n4624), .A2(n5412), .ZN(n5430) );
  XNOR2_X1 U5617 ( .A(n5411), .B(n5410), .ZN(n7648) );
  XNOR2_X1 U5618 ( .A(n5394), .B(n5393), .ZN(n7579) );
  OAI21_X1 U5619 ( .B1(n5335), .B2(n4322), .A(n4636), .ZN(n5394) );
  NAND2_X1 U5620 ( .A1(n4639), .A2(n5351), .ZN(n5371) );
  NAND2_X1 U5621 ( .A1(n5335), .A2(n4640), .ZN(n4639) );
  XNOR2_X1 U5622 ( .A(n5333), .B(n5332), .ZN(n7449) );
  XNOR2_X1 U5623 ( .A(n5315), .B(n5314), .ZN(n7392) );
  XNOR2_X1 U5624 ( .A(n5159), .B(n5154), .ZN(n6756) );
  NAND2_X1 U5625 ( .A1(n5137), .A2(n5136), .ZN(n5159) );
  XNOR2_X1 U5626 ( .A(n5135), .B(n5134), .ZN(n6684) );
  NAND2_X1 U5627 ( .A1(n4621), .A2(n5075), .ZN(n5093) );
  NAND2_X1 U5628 ( .A1(n5074), .A2(n4822), .ZN(n4621) );
  XNOR2_X1 U5629 ( .A(n5050), .B(n4323), .ZN(n6616) );
  XNOR2_X1 U5630 ( .A(n4973), .B(SI_5_), .ZN(n4971) );
  XNOR2_X1 U5631 ( .A(n4949), .B(SI_4_), .ZN(n4947) );
  XNOR2_X1 U5632 ( .A(n4921), .B(SI_3_), .ZN(n4919) );
  XNOR2_X1 U5633 ( .A(n4906), .B(SI_2_), .ZN(n4905) );
  AND2_X1 U5634 ( .A1(n5711), .A2(n5692), .ZN(n4387) );
  NAND2_X1 U5635 ( .A1(n6942), .A2(n5692), .ZN(n8035) );
  NAND2_X1 U5636 ( .A1(n5696), .A2(n5695), .ZN(n8039) );
  NAND2_X1 U5637 ( .A1(n4726), .A2(n6021), .ZN(n8044) );
  NAND2_X1 U5638 ( .A1(n4731), .A2(n4271), .ZN(n4726) );
  AND4_X1 U5639 ( .A1(n5741), .A2(n5740), .A3(n5739), .A4(n5738), .ZN(n7359)
         );
  NAND2_X1 U5640 ( .A1(n7231), .A2(n7232), .ZN(n7244) );
  OAI21_X1 U5641 ( .B1(n7234), .B2(n4740), .A(n4737), .ZN(n7339) );
  AND3_X1 U5642 ( .A1(n5900), .A2(n5899), .A3(n5898), .ZN(n8138) );
  NAND2_X1 U5643 ( .A1(n6150), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5898) );
  AND4_X1 U5644 ( .A1(n5775), .A2(n5774), .A3(n5773), .A4(n5772), .ZN(n7588)
         );
  OR2_X1 U5645 ( .A1(n8216), .A2(n6828), .ZN(n8194) );
  NAND2_X1 U5646 ( .A1(n5858), .A2(n5857), .ZN(n8692) );
  NAND2_X1 U5647 ( .A1(n8079), .A2(n5919), .ZN(n8171) );
  NAND2_X1 U5648 ( .A1(n7443), .A2(n5801), .ZN(n6556) );
  AND4_X1 U5649 ( .A1(n5759), .A2(n5758), .A3(n5757), .A4(n5756), .ZN(n7404)
         );
  AND4_X1 U5650 ( .A1(n5795), .A2(n5794), .A3(n5793), .A4(n5792), .ZN(n7600)
         );
  NAND2_X1 U5651 ( .A1(n6766), .A2(n6767), .ZN(n6765) );
  NAND2_X1 U5652 ( .A1(n4731), .A2(n8117), .ZN(n8207) );
  NAND2_X1 U5653 ( .A1(n7971), .A2(n7972), .ZN(n8124) );
  NAND2_X1 U5654 ( .A1(n4669), .A2(n5837), .ZN(n7976) );
  NAND2_X1 U5655 ( .A1(n6883), .A2(n5713), .ZN(n4669) );
  INV_X1 U5656 ( .A(n8216), .ZN(n8181) );
  NAND2_X1 U5657 ( .A1(n6150), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6149) );
  OR2_X1 U5658 ( .A1(n8432), .A2(n6038), .ZN(n6018) );
  NAND2_X1 U5659 ( .A1(n6004), .A2(n6003), .ZN(n8472) );
  NAND4_X2 U5660 ( .A1(n5598), .A2(n5597), .A3(n5596), .A4(n5595), .ZN(n6829)
         );
  INV_X1 U5661 ( .A(n4419), .ZN(n6739) );
  AND2_X1 U5662 ( .A1(n4419), .A2(n4418), .ZN(n6721) );
  NAND2_X1 U5663 ( .A1(n6723), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n4418) );
  INV_X1 U5664 ( .A(n4425), .ZN(n8245) );
  INV_X1 U5665 ( .A(n4423), .ZN(n8285) );
  INV_X1 U5666 ( .A(n4421), .ZN(n8298) );
  AND2_X1 U5667 ( .A1(n4421), .A2(n4420), .ZN(n6900) );
  NAND2_X1 U5668 ( .A1(n8297), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4420) );
  XNOR2_X1 U5669 ( .A(n4428), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U5670 ( .A1(n8370), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U5671 ( .A1(n8360), .A2(n4430), .ZN(n4429) );
  INV_X1 U5672 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n4430) );
  INV_X1 U5673 ( .A(n8618), .ZN(n8384) );
  NAND2_X1 U5674 ( .A1(n4752), .A2(n4753), .ZN(n8413) );
  NAND2_X1 U5675 ( .A1(n8498), .A2(n4611), .ZN(n8450) );
  NAND2_X1 U5676 ( .A1(n8484), .A2(n4825), .ZN(n8463) );
  NAND2_X1 U5677 ( .A1(n8508), .A2(n4588), .ZN(n8478) );
  AND2_X1 U5678 ( .A1(n5936), .A2(n5935), .ZN(n8524) );
  NAND2_X1 U5679 ( .A1(n6129), .A2(n6251), .ZN(n8535) );
  AND2_X1 U5680 ( .A1(n4771), .A2(n7992), .ZN(n8562) );
  NAND2_X1 U5681 ( .A1(n8591), .A2(n4824), .ZN(n8580) );
  NAND2_X1 U5682 ( .A1(n4782), .A2(n4781), .ZN(n7990) );
  NAND2_X1 U5683 ( .A1(n7597), .A2(n6221), .ZN(n7617) );
  NAND2_X1 U5684 ( .A1(n5788), .A2(n5787), .ZN(n9928) );
  NAND2_X1 U5685 ( .A1(n7256), .A2(n7355), .ZN(n7395) );
  NAND2_X1 U5686 ( .A1(n4762), .A2(n7169), .ZN(n7250) );
  NAND2_X1 U5687 ( .A1(n7045), .A2(n7044), .ZN(n4572) );
  NAND2_X1 U5688 ( .A1(n4584), .A2(n6175), .ZN(n7101) );
  OR3_X1 U5689 ( .A1(n7052), .A2(n7051), .A3(n8377), .ZN(n9819) );
  INV_X1 U5690 ( .A(n6807), .ZN(n7068) );
  INV_X1 U5691 ( .A(n9839), .ZN(n9814) );
  OR2_X1 U5692 ( .A1(n8495), .A2(n7041), .ZN(n8604) );
  NOR2_X1 U5693 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5582) );
  INV_X1 U5694 ( .A(n5585), .ZN(n6060) );
  INV_X1 U5695 ( .A(n5580), .ZN(n7411) );
  NAND2_X1 U5696 ( .A1(n5575), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4383) );
  INV_X1 U5697 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6579) );
  INV_X1 U5698 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6573) );
  INV_X1 U5699 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6571) );
  INV_X1 U5700 ( .A(n8862), .ZN(n7499) );
  INV_X1 U5701 ( .A(n6475), .ZN(n4415) );
  NAND2_X1 U5702 ( .A1(n6476), .A2(n8801), .ZN(n4416) );
  NAND2_X1 U5703 ( .A1(n6421), .A2(n6420), .ZN(n7289) );
  OAI21_X1 U5704 ( .B1(n4967), .B2(n6639), .A(n4500), .ZN(n4503) );
  NAND2_X1 U5705 ( .A1(n4967), .A2(n4501), .ZN(n4500) );
  NAND2_X1 U5706 ( .A1(n8753), .A2(n6464), .ZN(n8766) );
  NAND2_X1 U5707 ( .A1(n4798), .A2(n4797), .ZN(n4796) );
  XNOR2_X1 U5708 ( .A(n6389), .B(n6388), .ZN(n6860) );
  NAND2_X1 U5709 ( .A1(n4412), .A2(n4413), .ZN(n8783) );
  NAND2_X1 U5710 ( .A1(n6475), .A2(n4417), .ZN(n4413) );
  AOI21_X1 U5711 ( .B1(n6476), .B2(n4414), .A(n4408), .ZN(n4412) );
  NAND2_X1 U5712 ( .A1(n8783), .A2(n8784), .ZN(n8782) );
  NAND2_X1 U5713 ( .A1(n7545), .A2(n6444), .ZN(n7572) );
  NAND2_X1 U5714 ( .A1(n4402), .A2(n6431), .ZN(n7456) );
  NAND2_X1 U5715 ( .A1(n7424), .A2(n6430), .ZN(n4402) );
  NAND2_X1 U5716 ( .A1(n5230), .A2(n5229), .ZN(n9236) );
  AND2_X1 U5717 ( .A1(n6539), .A2(n9589), .ZN(n8831) );
  NAND2_X1 U5718 ( .A1(n8814), .A2(n8815), .ZN(n8813) );
  NAND2_X1 U5719 ( .A1(n7010), .A2(n6400), .ZN(n8814) );
  INV_X1 U5720 ( .A(n8844), .ZN(n8833) );
  INV_X1 U5721 ( .A(n8807), .ZN(n8843) );
  INV_X1 U5722 ( .A(n8837), .ZN(n8850) );
  AND2_X1 U5723 ( .A1(n7955), .A2(n4631), .ZN(n4630) );
  NOR2_X1 U5724 ( .A1(n7393), .A2(n7794), .ZN(n4631) );
  NAND2_X1 U5725 ( .A1(n4440), .A2(n4299), .ZN(n4437) );
  NOR2_X1 U5726 ( .A1(n4632), .A2(n7964), .ZN(n4440) );
  AND2_X1 U5727 ( .A1(n4629), .A2(n7965), .ZN(n4628) );
  OR2_X1 U5728 ( .A1(n7958), .A2(n7957), .ZN(n4629) );
  NAND2_X1 U5729 ( .A1(n5388), .A2(n5387), .ZN(n8856) );
  OR2_X1 U5730 ( .A1(n9011), .A2(n5231), .ZN(n5388) );
  INV_X1 U5731 ( .A(n4513), .ZN(n9580) );
  INV_X1 U5732 ( .A(n4511), .ZN(n9425) );
  NOR2_X1 U5733 ( .A1(n9423), .A2(n4509), .ZN(n9598) );
  AND2_X1 U5734 ( .A1(n6642), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n4509) );
  AOI21_X1 U5735 ( .B1(n6657), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6652), .ZN(
        n6632) );
  NOR2_X1 U5736 ( .A1(n8907), .A2(n8906), .ZN(n8910) );
  NOR2_X1 U5737 ( .A1(n8940), .A2(n8941), .ZN(n8946) );
  INV_X1 U5738 ( .A(n8967), .ZN(n9523) );
  AOI21_X1 U5739 ( .B1(n4356), .B2(n9701), .A(n4353), .ZN(n9199) );
  NAND2_X1 U5740 ( .A1(n4355), .A2(n4354), .ZN(n4353) );
  XNOR2_X1 U5741 ( .A(n9020), .B(n9019), .ZN(n4356) );
  NAND2_X1 U5742 ( .A1(n9054), .A2(n9154), .ZN(n4354) );
  NAND2_X1 U5743 ( .A1(n9025), .A2(n5529), .ZN(n9009) );
  NAND2_X1 U5744 ( .A1(n9041), .A2(n5528), .ZN(n9027) );
  NAND2_X1 U5745 ( .A1(n9070), .A2(n9069), .ZN(n9068) );
  NAND2_X1 U5746 ( .A1(n4714), .A2(n4718), .ZN(n9079) );
  NAND2_X1 U5747 ( .A1(n9112), .A2(n4719), .ZN(n4714) );
  OR2_X1 U5748 ( .A1(n9247), .A2(n5492), .ZN(n9105) );
  NAND2_X1 U5749 ( .A1(n4721), .A2(n4719), .ZN(n9093) );
  NAND2_X1 U5750 ( .A1(n4723), .A2(n4722), .ZN(n4721) );
  NAND2_X1 U5751 ( .A1(n9134), .A2(n7891), .ZN(n9120) );
  AOI21_X1 U5752 ( .B1(n9160), .B2(n5519), .A(n4686), .ZN(n4682) );
  OR2_X1 U5753 ( .A1(n7497), .A2(n4705), .ZN(n4697) );
  INV_X1 U5754 ( .A(n7459), .ZN(n9552) );
  NAND2_X1 U5755 ( .A1(n7301), .A2(n7845), .ZN(n7300) );
  NAND2_X1 U5756 ( .A1(n4692), .A2(n4691), .ZN(n7301) );
  NAND2_X1 U5757 ( .A1(n7159), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U5758 ( .A1(n7320), .A2(n5503), .ZN(n7132) );
  NAND2_X1 U5759 ( .A1(n7192), .A2(n4826), .ZN(n9742) );
  AND2_X1 U5760 ( .A1(n4933), .A2(n4932), .ZN(n7183) );
  NAND2_X1 U5761 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  INV_X1 U5762 ( .A(n9710), .ZN(n9107) );
  INV_X1 U5763 ( .A(n9105), .ZN(n9707) );
  XNOR2_X1 U5764 ( .A(n6163), .B(n6162), .ZN(n9405) );
  MUX2_X1 U5765 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4849), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n4851) );
  AND2_X1 U5766 ( .A1(n5226), .A2(n5209), .ZN(n8939) );
  INV_X1 U5767 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6609) );
  NOR2_X1 U5768 ( .A1(n4991), .A2(n4990), .ZN(n6996) );
  AND2_X1 U5769 ( .A1(n4829), .A2(n4828), .ZN(n4926) );
  XNOR2_X1 U5770 ( .A(n4875), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9592) );
  NOR2_X1 U5771 ( .A1(n7488), .A2(n9990), .ZN(n9981) );
  OAI21_X1 U5772 ( .B1(n4346), .B2(n4285), .A(n4345), .ZN(n8119) );
  NAND2_X1 U5773 ( .A1(n8161), .A2(n5657), .ZN(n6955) );
  OAI21_X1 U5774 ( .B1(n6326), .B2(n6327), .A(n6325), .ZN(n6333) );
  AOI21_X1 U5775 ( .B1(n4816), .B2(n4281), .A(n4329), .ZN(n4814) );
  INV_X1 U5776 ( .A(n4816), .ZN(n4815) );
  OAI22_X1 U5777 ( .A1(n4373), .A2(n7953), .B1(n8951), .B2(n4371), .ZN(n8958)
         );
  NAND2_X1 U5778 ( .A1(n4372), .A2(n7953), .ZN(n4371) );
  AOI21_X1 U5779 ( .B1(n9181), .B2(n9692), .A(n5542), .ZN(n5543) );
  OAI21_X1 U5780 ( .B1(n4496), .B2(n4495), .A(n4334), .ZN(P1_U3520) );
  INV_X1 U5781 ( .A(n9255), .ZN(n4496) );
  NAND2_X1 U5782 ( .A1(n5805), .A2(n5804), .ZN(n7614) );
  NAND2_X1 U5783 ( .A1(n5892), .A2(n5891), .ZN(n8681) );
  OR2_X1 U5784 ( .A1(n6463), .A2(n6462), .ZN(n6464) );
  NAND2_X1 U5785 ( .A1(n6438), .A2(n6437), .ZN(n4269) );
  INV_X1 U5786 ( .A(n9493), .ZN(n4534) );
  OR2_X1 U5787 ( .A1(n6277), .A2(n6279), .ZN(n4270) );
  AND2_X1 U5788 ( .A1(n6304), .A2(n6303), .ZN(n7258) );
  NOR2_X1 U5789 ( .A1(n8206), .A2(n4730), .ZN(n4271) );
  AND2_X1 U5790 ( .A1(n4499), .A2(n9531), .ZN(n4272) );
  INV_X1 U5791 ( .A(n7881), .ZN(n4686) );
  AND2_X1 U5792 ( .A1(n9223), .A2(n9121), .ZN(n4273) );
  INV_X1 U5793 ( .A(n6284), .ZN(n4473) );
  AND3_X1 U5794 ( .A1(n5551), .A2(n5552), .A3(n5589), .ZN(n4274) );
  NAND2_X1 U5795 ( .A1(n6263), .A2(n6250), .ZN(n8482) );
  INV_X1 U5796 ( .A(n8403), .ZN(n8394) );
  AND2_X1 U5797 ( .A1(n4750), .A2(n8403), .ZN(n4275) );
  AND2_X1 U5798 ( .A1(n7896), .A2(n7891), .ZN(n9136) );
  INV_X1 U5799 ( .A(n9136), .ZN(n9127) );
  OR2_X1 U5800 ( .A1(n5629), .A2(n6576), .ZN(n4276) );
  OAI21_X1 U5801 ( .B1(n7954), .B2(n7953), .A(n7957), .ZN(n4632) );
  NOR3_X1 U5802 ( .A1(n8681), .A2(n4602), .A3(n8671), .ZN(n4277) );
  NOR2_X1 U5803 ( .A1(n8114), .A2(n4733), .ZN(n4278) );
  AND2_X1 U5804 ( .A1(n4272), .A2(n4498), .ZN(n4280) );
  INV_X1 U5805 ( .A(n4439), .ZN(n4438) );
  NOR2_X1 U5806 ( .A1(n4628), .A2(n7964), .ZN(n4439) );
  NAND2_X1 U5807 ( .A1(n4806), .A2(n4807), .ZN(n7348) );
  AND2_X1 U5808 ( .A1(n6524), .A2(n6523), .ZN(n4281) );
  AND2_X1 U5809 ( .A1(n4599), .A2(n4598), .ZN(n4282) );
  OR2_X1 U5810 ( .A1(n5580), .A2(n6172), .ZN(n6279) );
  INV_X1 U5811 ( .A(n8815), .ZN(n4801) );
  NAND2_X1 U5812 ( .A1(n6759), .A2(n6830), .ZN(n6297) );
  XNOR2_X1 U5813 ( .A(n9211), .B(n9088), .ZN(n9069) );
  INV_X1 U5814 ( .A(n4954), .ZN(n5015) );
  NAND2_X1 U5815 ( .A1(n6424), .A2(n6423), .ZN(n4283) );
  AND2_X1 U5816 ( .A1(n7313), .A2(n9676), .ZN(n7737) );
  NAND2_X1 U5817 ( .A1(n5466), .A2(n4819), .ZN(n4865) );
  INV_X1 U5818 ( .A(n4470), .ZN(n4469) );
  AOI21_X1 U5819 ( .B1(n4476), .B2(n6275), .A(n4471), .ZN(n4470) );
  NAND2_X1 U5820 ( .A1(n8234), .A2(n7060), .ZN(n6294) );
  NAND2_X1 U5821 ( .A1(n5415), .A2(n5414), .ZN(n8982) );
  AND2_X1 U5822 ( .A1(n4845), .A2(n4844), .ZN(n4284) );
  OR3_X1 U5823 ( .A1(n4730), .A2(n8216), .A3(n8114), .ZN(n4285) );
  AND2_X1 U5824 ( .A1(n9453), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4286) );
  INV_X1 U5825 ( .A(n6281), .ZN(n4582) );
  NAND2_X1 U5826 ( .A1(n7614), .A2(n8226), .ZN(n4287) );
  INV_X1 U5827 ( .A(n4977), .ZN(n4672) );
  OR2_X1 U5828 ( .A1(n8687), .A2(n8570), .ZN(n7992) );
  INV_X1 U5829 ( .A(n7891), .ZN(n4550) );
  OR2_X1 U5830 ( .A1(n6290), .A2(n6288), .ZN(n4288) );
  AND3_X1 U5831 ( .A1(n6224), .A2(n6122), .A3(n6223), .ZN(n4289) );
  INV_X1 U5832 ( .A(n6292), .ZN(n4562) );
  INV_X1 U5833 ( .A(n7372), .ZN(n6319) );
  XNOR2_X1 U5834 ( .A(n4383), .B(n4382), .ZN(n7372) );
  INV_X1 U5835 ( .A(n7131), .ZN(n4674) );
  INV_X1 U5836 ( .A(n5513), .ZN(n4707) );
  OAI22_X1 U5837 ( .A1(n8992), .A2(n7922), .B1(n9191), .B2(n9021), .ZN(n8971)
         );
  NAND2_X1 U5838 ( .A1(n6280), .A2(n6281), .ZN(n8002) );
  INV_X1 U5839 ( .A(n8002), .ZN(n4475) );
  AOI21_X1 U5840 ( .B1(n7979), .B2(n5713), .A(n6147), .ZN(n8625) );
  OR2_X1 U5841 ( .A1(n6250), .A2(n6288), .ZN(n4290) );
  NOR2_X1 U5842 ( .A1(n7705), .A2(n8864), .ZN(n4291) );
  NOR2_X1 U5843 ( .A1(n7416), .A2(n9675), .ZN(n7848) );
  AND2_X1 U5844 ( .A1(n5993), .A2(n4725), .ZN(n4292) );
  NAND2_X1 U5845 ( .A1(n7924), .A2(n7925), .ZN(n8999) );
  AND2_X1 U5846 ( .A1(n6262), .A2(n6264), .ZN(n4293) );
  NAND2_X1 U5847 ( .A1(n8390), .A2(n6167), .ZN(n4294) );
  NAND2_X1 U5848 ( .A1(n8498), .A2(n4609), .ZN(n4612) );
  AND2_X1 U5849 ( .A1(n4721), .A2(n5524), .ZN(n4295) );
  INV_X1 U5850 ( .A(n5525), .ZN(n4722) );
  INV_X1 U5851 ( .A(n6481), .ZN(n4417) );
  NAND2_X1 U5852 ( .A1(n5322), .A2(n5321), .ZN(n9211) );
  AND2_X1 U5853 ( .A1(n4713), .A2(n5528), .ZN(n4296) );
  INV_X1 U5854 ( .A(n8656), .ZN(n8491) );
  NAND2_X1 U5855 ( .A1(n5967), .A2(n5966), .ZN(n8656) );
  INV_X1 U5856 ( .A(n8650), .ZN(n8467) );
  NAND2_X1 U5857 ( .A1(n5969), .A2(n5968), .ZN(n8650) );
  INV_X1 U5858 ( .A(n4703), .ZN(n4702) );
  OAI21_X1 U5859 ( .B1(n4706), .B2(n7708), .A(n4704), .ZN(n4703) );
  INV_X1 U5860 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4382) );
  INV_X1 U5861 ( .A(n8117), .ZN(n4730) );
  NOR2_X1 U5862 ( .A1(n7416), .A2(n8863), .ZN(n4297) );
  INV_X1 U5863 ( .A(n5507), .ZN(n4695) );
  INV_X1 U5864 ( .A(n4505), .ZN(n9044) );
  NOR2_X1 U5865 ( .A1(n9101), .A2(n4507), .ZN(n4505) );
  OR2_X1 U5866 ( .A1(n9226), .A2(n9099), .ZN(n7900) );
  INV_X1 U5867 ( .A(n7900), .ZN(n4547) );
  AND2_X1 U5868 ( .A1(n6260), .A2(n8515), .ZN(n4298) );
  NAND2_X1 U5869 ( .A1(n7951), .A2(n7953), .ZN(n4299) );
  NOR2_X1 U5870 ( .A1(n5120), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5139) );
  OR2_X1 U5871 ( .A1(n8630), .A2(n4471), .ZN(n4300) );
  AND2_X1 U5872 ( .A1(n7292), .A2(n9755), .ZN(n4301) );
  NOR2_X1 U5873 ( .A1(n8636), .A2(n8219), .ZN(n4302) );
  AND2_X1 U5874 ( .A1(n7982), .A2(n7983), .ZN(n4303) );
  NAND2_X1 U5875 ( .A1(n7952), .A2(n7953), .ZN(n4304) );
  AND2_X1 U5876 ( .A1(n6317), .A2(n6288), .ZN(n4305) );
  OR2_X1 U5877 ( .A1(n6271), .A2(n4474), .ZN(n4306) );
  INV_X1 U5878 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5448) );
  OAI21_X1 U5879 ( .B1(n4747), .B2(n8394), .A(n4300), .ZN(n4746) );
  OAI21_X1 U5880 ( .B1(n6460), .B2(n4790), .A(n8767), .ZN(n4789) );
  NAND2_X1 U5881 ( .A1(n8483), .A2(n8482), .ZN(n8484) );
  NOR2_X1 U5882 ( .A1(n7996), .A2(n8650), .ZN(n4307) );
  AND2_X1 U5883 ( .A1(n4395), .A2(n4397), .ZN(n4308) );
  OR2_X1 U5884 ( .A1(n8628), .A2(n8405), .ZN(n6280) );
  INV_X1 U5885 ( .A(n4750), .ZN(n4749) );
  AND2_X1 U5886 ( .A1(n4753), .A2(n4751), .ZN(n4750) );
  INV_X1 U5887 ( .A(n4589), .ZN(n4588) );
  NAND2_X1 U5888 ( .A1(n8479), .A2(n6259), .ZN(n4589) );
  NAND2_X1 U5889 ( .A1(n7753), .A2(n7821), .ZN(n7759) );
  OR2_X1 U5890 ( .A1(n6117), .A2(n4571), .ZN(n4309) );
  AND2_X1 U5891 ( .A1(n4415), .A2(n4416), .ZN(n4310) );
  AND2_X1 U5892 ( .A1(n9182), .A2(n4497), .ZN(n4311) );
  AND2_X1 U5893 ( .A1(n4795), .A2(n6503), .ZN(n4312) );
  OR2_X1 U5894 ( .A1(n5990), .A2(n5991), .ZN(n4313) );
  AND2_X1 U5895 ( .A1(n6134), .A2(n6250), .ZN(n4314) );
  AND2_X1 U5896 ( .A1(n5993), .A2(n4278), .ZN(n4315) );
  AND2_X1 U5897 ( .A1(n6122), .A2(n6221), .ZN(n4316) );
  AND2_X1 U5898 ( .A1(n4742), .A2(n4382), .ZN(n4317) );
  INV_X1 U5899 ( .A(n6021), .ZN(n4729) );
  NOR2_X1 U5900 ( .A1(n8975), .A2(n4553), .ZN(n4552) );
  AND2_X1 U5901 ( .A1(n8484), .A2(n4774), .ZN(n4318) );
  AOI21_X1 U5902 ( .B1(n4552), .B2(n8999), .A(n5428), .ZN(n4551) );
  AND2_X1 U5903 ( .A1(n8508), .A2(n6259), .ZN(n4319) );
  AND2_X1 U5904 ( .A1(n4283), .A2(n4808), .ZN(n4320) );
  INV_X1 U5905 ( .A(n8642), .ZN(n8434) );
  NAND2_X1 U5906 ( .A1(n6009), .A2(n6008), .ZN(n8642) );
  INV_X1 U5907 ( .A(n4401), .ZN(n4399) );
  NAND2_X1 U5908 ( .A1(n6431), .A2(n4269), .ZN(n4401) );
  INV_X1 U5909 ( .A(n6464), .ZN(n4790) );
  OR2_X1 U5910 ( .A1(n4439), .A2(n4304), .ZN(n4321) );
  INV_X2 U5911 ( .A(n5629), .ZN(n5887) );
  INV_X1 U5912 ( .A(n8126), .ZN(n4668) );
  OR2_X1 U5913 ( .A1(n5370), .A2(n4638), .ZN(n4322) );
  AND2_X1 U5914 ( .A1(n5051), .A2(n5035), .ZN(n4323) );
  XNOR2_X1 U5915 ( .A(n8636), .B(n8219), .ZN(n8422) );
  INV_X1 U5916 ( .A(n8422), .ZN(n4751) );
  INV_X1 U5917 ( .A(n4720), .ZN(n4719) );
  AND2_X1 U5918 ( .A1(n6044), .A2(n6043), .ZN(n8045) );
  INV_X1 U5919 ( .A(n8045), .ZN(n4471) );
  INV_X1 U5920 ( .A(n4682), .ZN(n9143) );
  NAND2_X1 U5921 ( .A1(n4697), .A2(n4702), .ZN(n7531) );
  XNOR2_X1 U5922 ( .A(n5463), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5474) );
  AND2_X1 U5923 ( .A1(n6889), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4324) );
  AND2_X1 U5924 ( .A1(n5292), .A2(n5283), .ZN(n4325) );
  INV_X1 U5925 ( .A(n7830), .ZN(n4531) );
  INV_X1 U5926 ( .A(n8726), .ZN(n4797) );
  NAND2_X1 U5927 ( .A1(n7546), .A2(n7547), .ZN(n7545) );
  AND2_X1 U5928 ( .A1(n8628), .A2(n9927), .ZN(n4326) );
  AND2_X1 U5929 ( .A1(n7001), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4327) );
  OR2_X1 U5930 ( .A1(n8610), .A2(n8692), .ZN(n8593) );
  NOR2_X1 U5931 ( .A1(n8593), .A2(n8687), .ZN(n4605) );
  AND2_X1 U5932 ( .A1(n5091), .A2(SI_11_), .ZN(n4328) );
  INV_X1 U5933 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6576) );
  OR2_X1 U5934 ( .A1(n6536), .A2(n6552), .ZN(n4329) );
  AND2_X1 U5935 ( .A1(n5245), .A2(SI_18_), .ZN(n4330) );
  INV_X1 U5936 ( .A(n4647), .ZN(n4646) );
  NAND2_X1 U5937 ( .A1(n4648), .A2(n5243), .ZN(n4647) );
  AND2_X1 U5938 ( .A1(n6533), .A2(n8829), .ZN(n4331) );
  AND2_X1 U5939 ( .A1(n8122), .A2(n5871), .ZN(n4332) );
  AND2_X1 U5940 ( .A1(n4782), .A2(n4287), .ZN(n4333) );
  OR2_X1 U5941 ( .A1(n6817), .A2(n7050), .ZN(n9950) );
  INV_X1 U5942 ( .A(n9767), .ZN(n4495) );
  INV_X1 U5943 ( .A(n8853), .ZN(n8829) );
  INV_X1 U5944 ( .A(n7614), .ZN(n4598) );
  INV_X1 U5945 ( .A(n8681), .ZN(n4604) );
  INV_X1 U5946 ( .A(n5621), .ZN(n5674) );
  NAND2_X1 U5947 ( .A1(n5875), .A2(n5874), .ZN(n8687) );
  INV_X1 U5948 ( .A(n8687), .ZN(n4603) );
  NAND2_X1 U5949 ( .A1(n4486), .A2(n4487), .ZN(n4485) );
  NAND2_X1 U5950 ( .A1(n7953), .A2(n6340), .ZN(n7941) );
  OR2_X1 U5951 ( .A1(n9767), .A2(n5438), .ZN(n4334) );
  NAND2_X1 U5952 ( .A1(n4572), .A2(n6176), .ZN(n7116) );
  NAND2_X1 U5953 ( .A1(n4563), .A2(n6303), .ZN(n7357) );
  AND2_X1 U5954 ( .A1(n6205), .A2(n6204), .ZN(n7251) );
  NAND2_X1 U5955 ( .A1(n5211), .A2(n5210), .ZN(n9243) );
  INV_X1 U5956 ( .A(n9243), .ZN(n4498) );
  OR2_X1 U5957 ( .A1(n6451), .A2(n6450), .ZN(n4335) );
  NOR2_X1 U5958 ( .A1(n5569), .A2(n5556), .ZN(n6053) );
  NAND2_X1 U5959 ( .A1(n5502), .A2(n5501), .ZN(n7320) );
  INV_X1 U5960 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5574) );
  AND2_X1 U5961 ( .A1(n8855), .A2(n7685), .ZN(n4336) );
  AND2_X1 U5962 ( .A1(n4806), .A2(n4804), .ZN(n4337) );
  OR2_X1 U5963 ( .A1(n6421), .A2(n6420), .ZN(n4338) );
  AND2_X1 U5964 ( .A1(n5432), .A2(n5431), .ZN(n4339) );
  AND2_X1 U5965 ( .A1(n7385), .A2(n8319), .ZN(n4340) );
  AND2_X1 U5966 ( .A1(n9866), .A2(n7309), .ZN(n4341) );
  NAND4_X1 U5967 ( .A1(n5566), .A2(n5567), .A3(n5568), .A4(n4784), .ZN(n6830)
         );
  INV_X1 U5968 ( .A(n8094), .ZN(n4606) );
  AND2_X1 U5969 ( .A1(n6765), .A2(n5609), .ZN(n4342) );
  INV_X1 U5970 ( .A(n8443), .ZN(n8377) );
  AND2_X1 U5971 ( .A1(n8357), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4343) );
  INV_X1 U5972 ( .A(n6639), .ZN(n4502) );
  INV_X1 U5973 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4494) );
  NAND2_X2 U5974 ( .A1(n6567), .A2(P2_U3152), .ZN(n8722) );
  NAND2_X1 U5975 ( .A1(n4351), .A2(n4311), .ZN(n9255) );
  NAND2_X1 U5976 ( .A1(n4976), .A2(n4975), .ZN(n4983) );
  OAI21_X1 U5977 ( .B1(n9183), .B2(n9529), .A(n4376), .ZN(n4352) );
  OAI21_X2 U5978 ( .B1(n4717), .B2(n9110), .A(n4715), .ZN(n9078) );
  NAND2_X1 U5979 ( .A1(n4479), .A2(n4664), .ZN(n4663) );
  NAND2_X1 U5980 ( .A1(n4481), .A2(n4290), .ZN(n4480) );
  NAND2_X1 U5981 ( .A1(n6248), .A2(n6279), .ZN(n4484) );
  NAND2_X1 U5982 ( .A1(n6286), .A2(n4492), .ZN(n4491) );
  NAND2_X1 U5983 ( .A1(n4660), .A2(n4659), .ZN(n6269) );
  OAI21_X1 U5984 ( .B1(n6283), .B2(n4305), .A(n4364), .ZN(n4363) );
  NAND2_X1 U5985 ( .A1(n4555), .A2(n7847), .ZN(n9510) );
  NAND2_X1 U5986 ( .A1(n8144), .A2(n4313), .ZN(n5993) );
  NAND2_X1 U5987 ( .A1(n4732), .A2(n5994), .ZN(n4346) );
  NAND2_X1 U5988 ( .A1(n7232), .A2(n4739), .ZN(n4738) );
  NAND2_X1 U5989 ( .A1(n6554), .A2(n5830), .ZN(n7561) );
  OAI21_X1 U5990 ( .B1(n7653), .B2(n5517), .A(n7877), .ZN(n9162) );
  NAND2_X1 U5991 ( .A1(n5073), .A2(n5508), .ZN(n4555) );
  XNOR2_X1 U5992 ( .A(n4347), .B(n7790), .ZN(n5459) );
  NAND2_X1 U5993 ( .A1(n4348), .A2(n4551), .ZN(n4347) );
  NAND2_X1 U5994 ( .A1(n9000), .A2(n4552), .ZN(n4348) );
  NAND2_X1 U5995 ( .A1(n7634), .A2(n7701), .ZN(n7653) );
  INV_X1 U5996 ( .A(n5153), .ZN(n4535) );
  NAND2_X1 U5997 ( .A1(n8408), .A2(n6273), .ZN(n8001) );
  AND2_X1 U5998 ( .A1(n6118), .A2(n7044), .ZN(n4357) );
  INV_X1 U5999 ( .A(n8505), .ZN(n6135) );
  NAND2_X1 U6000 ( .A1(n7170), .A2(n6204), .ZN(n7261) );
  AND2_X1 U6001 ( .A1(n4359), .A2(n4358), .ZN(n6327) );
  XNOR2_X1 U6002 ( .A(n6170), .B(n8443), .ZN(n4359) );
  AOI21_X2 U6003 ( .B1(n8605), .B2(n6224), .A(n6226), .ZN(n8598) );
  NAND2_X1 U6004 ( .A1(n4904), .A2(n4905), .ZN(n4909) );
  NAND2_X1 U6005 ( .A1(n4873), .A2(n4872), .ZN(n4904) );
  NAND2_X1 U6006 ( .A1(n6124), .A2(n6232), .ZN(n8585) );
  NAND2_X1 U6007 ( .A1(n7597), .A2(n4316), .ZN(n6123) );
  AOI21_X1 U6008 ( .B1(n6169), .B2(n6168), .A(n6285), .ZN(n6170) );
  NAND2_X1 U6009 ( .A1(n5052), .A2(n5051), .ZN(n5074) );
  NAND3_X1 U6010 ( .A1(n4378), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4667) );
  NAND2_X1 U6011 ( .A1(n8974), .A2(n5532), .ZN(n5533) );
  NAND2_X2 U6012 ( .A1(n5512), .A2(n5511), .ZN(n7497) );
  INV_X1 U6013 ( .A(n7628), .ZN(n4360) );
  OAI21_X1 U6014 ( .B1(n9505), .B2(n9552), .A(n7499), .ZN(n5510) );
  NOR2_X1 U6015 ( .A1(n4674), .A2(n4673), .ZN(n4677) );
  AOI21_X2 U6016 ( .B1(n8609), .B2(n8608), .A(n7991), .ZN(n8592) );
  OAI22_X2 U6017 ( .A1(n8545), .A2(n7993), .B1(n8553), .B2(n8537), .ZN(n8527)
         );
  INV_X1 U6018 ( .A(n6321), .ZN(n4490) );
  OAI211_X1 U6019 ( .C1(n6276), .C2(n4465), .A(n4463), .B(n4464), .ZN(n4462)
         );
  OAI211_X1 U6020 ( .C1(n4321), .C2(n4279), .A(n4436), .B(n4369), .ZN(P1_U3240) );
  NAND2_X1 U6021 ( .A1(n4437), .A2(n4438), .ZN(n4369) );
  NOR2_X1 U6022 ( .A1(n5586), .A2(n4557), .ZN(n4556) );
  NAND2_X1 U6023 ( .A1(n8513), .A2(n4827), .ZN(n7995) );
  NAND2_X1 U6024 ( .A1(n7168), .A2(n7167), .ZN(n4762) );
  NAND2_X1 U6025 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  NAND2_X1 U6026 ( .A1(n6869), .A2(n6870), .ZN(n7019) );
  NAND2_X1 U6027 ( .A1(n4593), .A2(n4591), .ZN(n8698) );
  NAND2_X1 U6028 ( .A1(n5282), .A2(n5281), .ZN(n4643) );
  NAND2_X1 U6029 ( .A1(n6323), .A2(n4488), .ZN(n6326) );
  AOI21_X1 U6030 ( .B1(n4462), .B2(n6282), .A(n4472), .ZN(n6283) );
  NAND2_X1 U6031 ( .A1(n4635), .A2(n4633), .ZN(n5396) );
  INV_X1 U6032 ( .A(n5184), .ZN(n5587) );
  NAND2_X4 U6033 ( .A1(n4667), .A2(n4867), .ZN(n5184) );
  NAND2_X1 U6034 ( .A1(n7630), .A2(n5516), .ZN(n7652) );
  NOR2_X2 U6035 ( .A1(n5989), .A2(n5988), .ZN(n8144) );
  NAND2_X2 U6036 ( .A1(n5965), .A2(n5964), .ZN(n5989) );
  NAND2_X1 U6037 ( .A1(n8122), .A2(n4380), .ZN(n8135) );
  NAND3_X1 U6038 ( .A1(n9866), .A2(n7309), .A3(n8443), .ZN(n5603) );
  OR2_X1 U6039 ( .A1(n6112), .A2(n6828), .ZN(n5608) );
  INV_X2 U6040 ( .A(n5603), .ZN(n6828) );
  NAND2_X1 U6041 ( .A1(n7443), .A2(n4384), .ZN(n6554) );
  NAND2_X1 U6042 ( .A1(n8087), .A2(n5712), .ZN(n5727) );
  NAND2_X1 U6043 ( .A1(n4387), .A2(n6942), .ZN(n8087) );
  NAND3_X1 U6044 ( .A1(n4274), .A2(n4783), .A3(n4268), .ZN(n5569) );
  NAND4_X1 U6045 ( .A1(n4274), .A2(n4783), .A3(n5570), .A4(n4268), .ZN(n5889)
         );
  OAI211_X2 U6046 ( .C1(n6400), .C2(n4801), .A(n4388), .B(n6409), .ZN(n7088)
         );
  OAI21_X1 U6047 ( .B1(n8838), .B2(n8841), .A(n8839), .ZN(n8752) );
  NAND3_X1 U6048 ( .A1(n4393), .A2(n4394), .A3(n4810), .ZN(n6454) );
  NAND3_X1 U6049 ( .A1(n4395), .A2(n4397), .A3(n4401), .ZN(n4394) );
  AOI21_X1 U6050 ( .B1(n7384), .B2(n4340), .A(n4434), .ZN(n4433) );
  NAND2_X1 U6051 ( .A1(n7384), .A2(n7385), .ZN(n8311) );
  NAND2_X1 U6052 ( .A1(n8311), .A2(n4435), .ZN(n8318) );
  NOR2_X1 U6053 ( .A1(n8313), .A2(n9466), .ZN(n8320) );
  NAND2_X1 U6054 ( .A1(n8311), .A2(n4432), .ZN(n4431) );
  NAND3_X1 U6055 ( .A1(n4279), .A2(n4438), .A3(n4630), .ZN(n4436) );
  NAND3_X1 U6056 ( .A1(n4554), .A2(n7728), .A3(n4980), .ZN(n4442) );
  INV_X1 U6057 ( .A(n7215), .ZN(n4444) );
  OAI21_X1 U6058 ( .B1(n4447), .B2(n4446), .A(n7875), .ZN(n4445) );
  NAND3_X1 U6059 ( .A1(n7843), .A2(n7943), .A3(n7842), .ZN(n4451) );
  AOI21_X1 U6060 ( .B1(n4452), .B2(n7910), .A(n7909), .ZN(n7918) );
  NAND3_X1 U6061 ( .A1(n7959), .A2(n9584), .A3(n9592), .ZN(n4876) );
  INV_X2 U6062 ( .A(n4967), .ZN(n5255) );
  NAND2_X2 U6063 ( .A1(n4863), .A2(n4862), .ZN(n7959) );
  NAND2_X1 U6064 ( .A1(n6174), .A2(n6288), .ZN(n4478) );
  INV_X1 U6065 ( .A(n6191), .ZN(n6195) );
  NAND3_X1 U6066 ( .A1(n6294), .A2(n7024), .A3(n6279), .ZN(n4477) );
  AND2_X1 U6067 ( .A1(n6294), .A2(n7024), .ZN(n6173) );
  NAND2_X2 U6068 ( .A1(n5565), .A2(n7981), .ZN(n5622) );
  XNOR2_X2 U6069 ( .A(n5560), .B(n4494), .ZN(n7981) );
  NOR2_X2 U6070 ( .A1(n9689), .A2(n7210), .ZN(n7204) );
  NAND2_X1 U6071 ( .A1(n9488), .A2(n4280), .ZN(n9167) );
  NAND2_X1 U6072 ( .A1(n4967), .A2(n6567), .ZN(n4977) );
  INV_X1 U6073 ( .A(n4504), .ZN(n9033) );
  NOR3_X2 U6074 ( .A1(n9101), .A2(n9203), .A3(n4507), .ZN(n4504) );
  NAND2_X1 U6075 ( .A1(n4524), .A2(n4523), .ZN(n5049) );
  NAND2_X1 U6076 ( .A1(n7122), .A2(n4526), .ZN(n4523) );
  OAI21_X1 U6077 ( .B1(n7122), .B2(n4527), .A(n4526), .ZN(n9673) );
  INV_X1 U6078 ( .A(n7632), .ZN(n5180) );
  NAND2_X1 U6079 ( .A1(n4247), .A2(n6851), .ZN(n6336) );
  NAND2_X1 U6080 ( .A1(n9150), .A2(n4544), .ZN(n4543) );
  NAND3_X1 U6081 ( .A1(n4933), .A2(n4932), .A3(n7732), .ZN(n4554) );
  NOR2_X2 U6082 ( .A1(n5447), .A2(n4710), .ZN(n5466) );
  NAND2_X2 U6083 ( .A1(n4558), .A2(n4556), .ZN(n8004) );
  NAND2_X1 U6084 ( .A1(n4560), .A2(n4561), .ZN(n7401) );
  NAND2_X1 U6085 ( .A1(n7261), .A2(n4564), .ZN(n4560) );
  INV_X1 U6086 ( .A(n4567), .ZN(n4568) );
  NAND2_X1 U6087 ( .A1(n8237), .A2(n7068), .ZN(n6181) );
  NAND2_X1 U6088 ( .A1(n8001), .A2(n4576), .ZN(n4573) );
  NAND2_X1 U6089 ( .A1(n4573), .A2(n4574), .ZN(n6169) );
  NAND2_X1 U6090 ( .A1(n6135), .A2(n4314), .ZN(n4587) );
  OR2_X2 U6091 ( .A1(n7596), .A2(n6120), .ZN(n7597) );
  NAND2_X1 U6092 ( .A1(n6129), .A2(n4590), .ZN(n8514) );
  NAND2_X1 U6093 ( .A1(n8514), .A2(n6132), .ZN(n6133) );
  NAND2_X1 U6094 ( .A1(n6119), .A2(n6307), .ZN(n7596) );
  NAND2_X1 U6095 ( .A1(n6298), .A2(n9827), .ZN(n9832) );
  NAND2_X1 U6096 ( .A1(n8402), .A2(n8394), .ZN(n8408) );
  NAND2_X1 U6097 ( .A1(n6112), .A2(n6114), .ZN(n6298) );
  NOR2_X2 U6098 ( .A1(n4485), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5585) );
  NOR2_X2 U6099 ( .A1(n4485), .A2(n4786), .ZN(n5586) );
  NAND2_X1 U6100 ( .A1(n4596), .A2(n4599), .ZN(n8610) );
  INV_X1 U6101 ( .A(n4599), .ZN(n9808) );
  INV_X1 U6102 ( .A(n8593), .ZN(n4600) );
  NAND2_X1 U6103 ( .A1(n4277), .A2(n4600), .ZN(n8528) );
  INV_X1 U6104 ( .A(n4605), .ZN(n8581) );
  INV_X1 U6105 ( .A(n4612), .ZN(n8449) );
  NAND2_X1 U6106 ( .A1(n5052), .A2(n4614), .ZN(n4613) );
  NAND2_X1 U6107 ( .A1(n5411), .A2(n5410), .ZN(n4624) );
  NAND2_X1 U6108 ( .A1(n5335), .A2(n4636), .ZN(n4635) );
  NAND2_X1 U6109 ( .A1(n5335), .A2(n5334), .ZN(n5353) );
  NAND2_X1 U6110 ( .A1(n4643), .A2(n5283), .ZN(n5291) );
  OAI21_X1 U6111 ( .B1(n5222), .B2(n5221), .A(n5225), .ZN(n5244) );
  NAND2_X1 U6112 ( .A1(n5137), .A2(n4653), .ZN(n4649) );
  NAND2_X1 U6113 ( .A1(n4649), .A2(n4650), .ZN(n5206) );
  NAND2_X1 U6114 ( .A1(n5137), .A2(n4657), .ZN(n4652) );
  NAND2_X1 U6115 ( .A1(n4679), .A2(n4683), .ZN(n5521) );
  NAND2_X1 U6116 ( .A1(n7651), .A2(n4680), .ZN(n4679) );
  AND2_X1 U6117 ( .A1(n9149), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U6118 ( .A1(n7159), .A2(n4688), .ZN(n4687) );
  NAND2_X1 U6119 ( .A1(n7497), .A2(n4701), .ZN(n4696) );
  NAND2_X1 U6120 ( .A1(n7497), .A2(n5513), .ZN(n9485) );
  NOR2_X1 U6121 ( .A1(n9486), .A2(n8860), .ZN(n4705) );
  INV_X1 U6122 ( .A(n4710), .ZN(n4709) );
  NAND2_X1 U6123 ( .A1(n9025), .A2(n4711), .ZN(n5530) );
  NAND2_X1 U6124 ( .A1(n5994), .A2(n4315), .ZN(n4731) );
  NAND2_X1 U6125 ( .A1(n4724), .A2(n4727), .ZN(n6035) );
  NAND2_X1 U6126 ( .A1(n5994), .A2(n4292), .ZN(n4724) );
  AND2_X1 U6127 ( .A1(n5993), .A2(n5992), .ZN(n4732) );
  INV_X1 U6128 ( .A(n5992), .ZN(n4733) );
  NAND2_X1 U6129 ( .A1(n8064), .A2(n5620), .ZN(n5639) );
  NAND2_X1 U6130 ( .A1(n7234), .A2(n4737), .ZN(n4734) );
  NAND2_X1 U6131 ( .A1(n4734), .A2(n4735), .ZN(n5780) );
  AOI21_X1 U6132 ( .B1(n4737), .B2(n4740), .A(n4736), .ZN(n4735) );
  AND2_X1 U6133 ( .A1(n7245), .A2(n4738), .ZN(n4737) );
  NAND2_X1 U6134 ( .A1(n5572), .A2(n4742), .ZN(n5575) );
  NAND2_X1 U6135 ( .A1(n5572), .A2(n4317), .ZN(n4741) );
  NAND2_X1 U6136 ( .A1(n6953), .A2(n5688), .ZN(n6942) );
  NAND2_X1 U6137 ( .A1(n8161), .A2(n4743), .ZN(n6953) );
  OAI21_X1 U6138 ( .B1(n7999), .B2(n4749), .A(n4747), .ZN(n8395) );
  NAND2_X1 U6139 ( .A1(n7999), .A2(n7998), .ZN(n8429) );
  AOI21_X2 U6140 ( .B1(n4745), .B2(n4275), .A(n4746), .ZN(n8000) );
  NAND2_X1 U6141 ( .A1(n7999), .A2(n4756), .ZN(n4752) );
  NAND2_X1 U6142 ( .A1(n4762), .A2(n4760), .ZN(n7254) );
  NAND2_X1 U6143 ( .A1(n8591), .A2(n4767), .ZN(n4763) );
  NAND2_X1 U6144 ( .A1(n4763), .A2(n4764), .ZN(n8545) );
  INV_X1 U6145 ( .A(n4771), .ZN(n8579) );
  OAI21_X2 U6146 ( .B1(n8483), .B2(n4773), .A(n4772), .ZN(n8447) );
  NAND2_X1 U6147 ( .A1(n7356), .A2(n4776), .ZN(n7399) );
  NAND2_X1 U6148 ( .A1(n7594), .A2(n4781), .ZN(n4778) );
  NAND2_X1 U6149 ( .A1(n4778), .A2(n4779), .ZN(n8609) );
  INV_X1 U6150 ( .A(n4782), .ZN(n7615) );
  NAND3_X1 U6151 ( .A1(n4268), .A2(n4783), .A3(n5647), .ZN(n5849) );
  NAND3_X1 U6152 ( .A1(n5565), .A2(n5564), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n4784) );
  NAND2_X1 U6153 ( .A1(n4788), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5561) );
  INV_X1 U6154 ( .A(n8752), .ZN(n4791) );
  NAND2_X1 U6155 ( .A1(n6505), .A2(n6504), .ZN(n8725) );
  NAND3_X1 U6156 ( .A1(n8792), .A2(n6502), .A3(n6503), .ZN(n4798) );
  NAND3_X1 U6157 ( .A1(n8792), .A2(n6502), .A3(n4312), .ZN(n4794) );
  NAND2_X1 U6158 ( .A1(n4796), .A2(n8725), .ZN(n8776) );
  INV_X1 U6159 ( .A(n8775), .ZN(n4795) );
  NOR2_X1 U6160 ( .A1(n4801), .A2(n4800), .ZN(n4799) );
  INV_X1 U6161 ( .A(n7011), .ZN(n4800) );
  NAND2_X1 U6162 ( .A1(n8828), .A2(n4331), .ZN(n4813) );
  OAI211_X1 U6163 ( .C1(n8828), .C2(n4815), .A(n4814), .B(n4813), .ZN(P1_U3212) );
  NAND2_X1 U6164 ( .A1(n8828), .A2(n6533), .ZN(n8032) );
  NAND2_X1 U6165 ( .A1(n5466), .A2(n4846), .ZN(n5464) );
  NAND2_X1 U6166 ( .A1(n5466), .A2(n4817), .ZN(n4862) );
  NAND3_X1 U6167 ( .A1(n4829), .A2(n4828), .A3(n4830), .ZN(n4955) );
  XNOR2_X1 U6168 ( .A(n5371), .B(n5370), .ZN(n7567) );
  OAI21_X1 U6169 ( .B1(n6160), .B2(n6159), .A(n6158), .ZN(n6163) );
  NAND2_X1 U6170 ( .A1(n5610), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5596) );
  OR2_X1 U6171 ( .A1(n9188), .A2(n9529), .ZN(n9189) );
  OR2_X1 U6172 ( .A1(n5545), .A2(n5544), .ZN(P1_U3355) );
  CLKBUF_X1 U6173 ( .A(n8135), .Z(n8193) );
  INV_X1 U6174 ( .A(n5889), .ZN(n5572) );
  AND2_X1 U6175 ( .A1(n6719), .A2(n8004), .ZN(n9787) );
  INV_X1 U6176 ( .A(n5592), .ZN(n5594) );
  NAND2_X1 U6177 ( .A1(n4934), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4889) );
  NAND2_X1 U6178 ( .A1(n4934), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U6179 ( .A1(n6360), .A2(n6359), .ZN(n6361) );
  AND2_X2 U6180 ( .A1(n5564), .A2(n8720), .ZN(n5623) );
  INV_X1 U6181 ( .A(n8720), .ZN(n5565) );
  NAND2_X1 U6182 ( .A1(n8734), .A2(n8735), .ZN(n8733) );
  NAND2_X1 U6183 ( .A1(n4967), .A2(n9419), .ZN(n4885) );
  AND2_X2 U6184 ( .A1(n4967), .A2(n5587), .ZN(n4954) );
  NAND2_X1 U6185 ( .A1(n8183), .A2(n8182), .ZN(n5965) );
  INV_X1 U6186 ( .A(n6353), .ZN(n6697) );
  NAND2_X1 U6187 ( .A1(n8592), .A2(n8597), .ZN(n8591) );
  OAI21_X1 U6188 ( .B1(n9183), .B2(n9176), .A(n5543), .ZN(n5544) );
  NAND2_X1 U6189 ( .A1(n6358), .A2(n4247), .ZN(n6359) );
  INV_X1 U6190 ( .A(n6358), .ZN(n9724) );
  XNOR2_X2 U6192 ( .A(n5989), .B(n5987), .ZN(n8052) );
  AND2_X1 U6193 ( .A1(n5976), .A2(n5975), .ZN(n8220) );
  INV_X1 U6194 ( .A(n8220), .ZN(n7996) );
  AND2_X1 U6195 ( .A1(n5075), .A2(n5056), .ZN(n4822) );
  NOR2_X1 U6196 ( .A1(n7688), .A2(n7915), .ZN(n4823) );
  OR2_X1 U6197 ( .A1(n8491), .A2(n8506), .ZN(n4825) );
  AND2_X1 U6198 ( .A1(n5499), .A2(n7191), .ZN(n4826) );
  AND2_X1 U6199 ( .A1(n5427), .A2(n5426), .ZN(n9001) );
  INV_X1 U6200 ( .A(n6705), .ZN(n6325) );
  INV_X1 U6201 ( .A(n9804), .ZN(n7592) );
  OR2_X1 U6202 ( .A1(n8524), .A2(n8539), .ZN(n4827) );
  INV_X1 U6203 ( .A(n9149), .ZN(n5241) );
  OR2_X1 U6204 ( .A1(n6817), .A2(n6800), .ZN(n9935) );
  INV_X1 U6205 ( .A(n5501), .ZN(n4980) );
  MUX2_X1 U6206 ( .A(n6230), .B(n6229), .S(n6279), .Z(n6231) );
  INV_X1 U6207 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4832) );
  INV_X1 U6208 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5550) );
  INV_X1 U6209 ( .A(n5840), .ZN(n5838) );
  INV_X1 U6210 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9331) );
  INV_X1 U6211 ( .A(n5977), .ZN(n5970) );
  OAI22_X1 U6212 ( .A1(n5628), .A2(n6568), .B1(n6710), .B2(n6727), .ZN(n5592)
         );
  NOR2_X1 U6213 ( .A1(n8384), .A2(n8383), .ZN(n6285) );
  INV_X1 U6214 ( .A(n5896), .ZN(n5895) );
  INV_X1 U6215 ( .A(n5860), .ZN(n5859) );
  INV_X1 U6216 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5557) );
  INV_X1 U6217 ( .A(n5324), .ZN(n5323) );
  INV_X1 U6218 ( .A(n5065), .ZN(n5064) );
  INV_X1 U6219 ( .A(n9001), .ZN(n5531) );
  INV_X1 U6220 ( .A(n5005), .ZN(n5006) );
  AND2_X1 U6221 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5697) );
  OR2_X1 U6222 ( .A1(n5629), .A2(n6569), .ZN(n5593) );
  NAND2_X1 U6223 ( .A1(n5658), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5701) );
  INV_X1 U6224 ( .A(n8125), .ZN(n5866) );
  NAND2_X1 U6225 ( .A1(n6829), .A2(n9865), .ZN(n9835) );
  NAND2_X1 U6226 ( .A1(n5952), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5977) );
  OR2_X1 U6227 ( .A1(n8146), .A2(n8149), .ZN(n5992) );
  NAND2_X1 U6228 ( .A1(n6010), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U6229 ( .A1(n5859), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5876) );
  INV_X1 U6230 ( .A(n8755), .ZN(n6460) );
  INV_X1 U6231 ( .A(n4938), .ZN(n4936) );
  INV_X1 U6232 ( .A(n5381), .ZN(n5379) );
  OR2_X1 U6233 ( .A1(n5146), .A2(n7670), .ZN(n5172) );
  NAND2_X1 U6234 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n4938) );
  AOI22_X1 U6235 ( .A1(n5531), .A2(n9154), .B1(n8961), .B2(n8855), .ZN(n5457)
         );
  INV_X1 U6236 ( .A(n7631), .ZN(n7870) );
  INV_X1 U6237 ( .A(SI_9_), .ZN(n9357) );
  INV_X1 U6238 ( .A(n8034), .ZN(n5711) );
  NAND2_X1 U6239 ( .A1(n5752), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5770) );
  OR2_X1 U6240 ( .A1(n5876), .A2(n8139), .ZN(n5896) );
  NAND2_X1 U6241 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5659) );
  OR2_X1 U6242 ( .A1(n5770), .A2(n5769), .ZN(n5790) );
  AND2_X1 U6243 ( .A1(n6012), .A2(n5999), .ZN(n8451) );
  OR2_X1 U6244 ( .A1(n5910), .A2(n5909), .ZN(n5924) );
  NOR2_X1 U6245 ( .A1(n4668), .A2(n7976), .ZN(n7991) );
  NAND2_X1 U6246 ( .A1(n7094), .A2(n7021), .ZN(n7022) );
  INV_X1 U6247 ( .A(n7976), .ZN(n9463) );
  AND2_X1 U6248 ( .A1(n6811), .A2(n6810), .ZN(n8533) );
  AND2_X1 U6249 ( .A1(n6066), .A2(n6065), .ZN(n6799) );
  NOR2_X1 U6250 ( .A1(n5581), .A2(n5582), .ZN(n5583) );
  AND2_X1 U6251 ( .A1(n8804), .A2(n8802), .ZN(n6475) );
  XNOR2_X1 U6252 ( .A(n6338), .B(n4266), .ZN(n6353) );
  OR2_X1 U6253 ( .A1(n5213), .A2(n5212), .ZN(n5233) );
  NAND2_X1 U6254 ( .A1(n7426), .A2(n7425), .ZN(n6431) );
  OR2_X1 U6255 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  OR2_X1 U6256 ( .A1(n6538), .A2(n9589), .ZN(n8807) );
  NAND2_X1 U6257 ( .A1(n5379), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5417) );
  AND2_X1 U6258 ( .A1(n5381), .A2(n5362), .ZN(n9035) );
  OR2_X1 U6259 ( .A1(n5259), .A2(n5258), .ZN(n5277) );
  INV_X1 U6260 ( .A(n5457), .ZN(n5458) );
  OR3_X1 U6261 ( .A1(n6838), .A2(n6362), .A3(n7953), .ZN(n9704) );
  INV_X1 U6262 ( .A(n8198), .ZN(n8209) );
  AND2_X1 U6263 ( .A1(n5985), .A2(n5984), .ZN(n8506) );
  AND4_X1 U6264 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(n8126)
         );
  AND2_X1 U6265 ( .A1(n6734), .A2(n6092), .ZN(n9454) );
  INV_X1 U6266 ( .A(n8373), .ZN(n9784) );
  INV_X1 U6267 ( .A(n8447), .ZN(n8448) );
  AND2_X1 U6268 ( .A1(n6620), .A2(n6093), .ZN(n8571) );
  NAND2_X1 U6269 ( .A1(n7039), .A2(n9814), .ZN(n9815) );
  INV_X1 U6270 ( .A(n4341), .ZN(n9921) );
  AND2_X1 U6271 ( .A1(n7605), .A2(n9473), .ZN(n9888) );
  OR2_X1 U6272 ( .A1(n6799), .A2(n6798), .ZN(n6817) );
  AND2_X1 U6273 ( .A1(n6706), .A2(n9864), .ZN(n9851) );
  AND2_X1 U6274 ( .A1(n5693), .A2(n5684), .ZN(n8258) );
  INV_X1 U6275 ( .A(n9517), .ZN(n9684) );
  AND2_X1 U6276 ( .A1(n9704), .A2(n9247), .ZN(n9529) );
  AND2_X1 U6277 ( .A1(n6780), .A2(n6779), .ZN(n6787) );
  AND2_X1 U6278 ( .A1(n5061), .A2(n5077), .ZN(n7001) );
  XNOR2_X1 U6279 ( .A(n4871), .B(n4870), .ZN(n4894) );
  OR3_X1 U6280 ( .A1(n7513), .A2(n7582), .A3(n7587), .ZN(n6706) );
  AOI21_X1 U6281 ( .B1(n6109), .B2(n8630), .A(n6108), .ZN(n6110) );
  INV_X1 U6282 ( .A(n8661), .ZN(n8503) );
  OR2_X1 U6283 ( .A1(n6331), .A2(n6330), .ZN(n6332) );
  AND2_X1 U6284 ( .A1(n6018), .A2(n6017), .ZN(n8111) );
  AND4_X1 U6285 ( .A1(n5865), .A2(n5864), .A3(n5863), .A4(n5862), .ZN(n8137)
         );
  INV_X1 U6286 ( .A(n9454), .ZN(n9789) );
  INV_X1 U6287 ( .A(n9815), .ZN(n9840) );
  AND2_X1 U6288 ( .A1(n6324), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9864) );
  XNOR2_X1 U6289 ( .A(n6052), .B(n6051), .ZN(n7513) );
  INV_X1 U6290 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6676) );
  INV_X1 U6291 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6611) );
  AND2_X1 U6292 ( .A1(n6535), .A2(n9105), .ZN(n8837) );
  NAND2_X1 U6293 ( .A1(n5409), .A2(n5408), .ZN(n9021) );
  AND2_X1 U6294 ( .A1(n7640), .A2(n7639), .ZN(n9253) );
  INV_X1 U6295 ( .A(n9684), .ZN(n9708) );
  AND2_X1 U6296 ( .A1(n6935), .A2(n9105), .ZN(n9517) );
  INV_X1 U6297 ( .A(n9783), .ZN(n9780) );
  INV_X1 U6298 ( .A(n9722), .ZN(n9723) );
  INV_X1 U6299 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6665) );
  NOR2_X1 U6300 ( .A1(n9981), .A2(n9980), .ZN(n9979) );
  NAND2_X1 U6301 ( .A1(n6333), .A2(n6332), .ZN(P2_U3244) );
  INV_X1 U6302 ( .A(n4957), .ZN(n4842) );
  INV_X2 U6303 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5208) );
  NAND2_X1 U6304 ( .A1(n5208), .A2(n4832), .ZN(n5251) );
  INV_X1 U6305 ( .A(n5251), .ZN(n4834) );
  NOR2_X1 U6306 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n4833) );
  NAND4_X1 U6307 ( .A1(n4834), .A2(n4833), .A3(n5059), .A4(n9331), .ZN(n4840)
         );
  NOR2_X1 U6308 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4838) );
  NOR2_X1 U6309 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4837) );
  NOR2_X1 U6310 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4836) );
  NOR2_X1 U6311 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n4835) );
  NAND4_X1 U6312 ( .A1(n4838), .A2(n4837), .A3(n4836), .A4(n4835), .ZN(n4839)
         );
  NOR2_X1 U6313 ( .A1(n4840), .A2(n4839), .ZN(n4841) );
  NAND2_X1 U6314 ( .A1(n4842), .A2(n4841), .ZN(n5447) );
  INV_X1 U6315 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U6316 ( .A1(n5444), .A2(n4843), .ZN(n5460) );
  INV_X1 U6317 ( .A(n5460), .ZN(n4845) );
  NOR2_X1 U6318 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n4844) );
  INV_X1 U6319 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4846) );
  INV_X1 U6320 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4847) );
  NOR2_X2 U6321 ( .A1(n4862), .A2(P1_IR_REG_29__SCAN_IN), .ZN(n4850) );
  OR2_X2 U6322 ( .A1(n4850), .A2(n9406), .ZN(n4848) );
  XNOR2_X2 U6323 ( .A(n4848), .B(P1_IR_REG_30__SCAN_IN), .ZN(n4853) );
  NAND2_X1 U6324 ( .A1(n4862), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4849) );
  INV_X1 U6325 ( .A(n4850), .ZN(n9407) );
  INV_X1 U6326 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n4852) );
  OR2_X1 U6327 ( .A1(n5236), .A2(n4852), .ZN(n4860) );
  NAND2_X1 U6328 ( .A1(n4935), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n4859) );
  INV_X1 U6329 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n4855) );
  MUX2_X1 U6330 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4864), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n4866) );
  NAND3_X1 U6331 ( .A1(n5184), .A2(SI_0_), .A3(P2_DATAO_REG_0__SCAN_IN), .ZN(
        n4869) );
  AND2_X1 U6332 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4868) );
  NAND2_X1 U6333 ( .A1(n4869), .A2(n5601), .ZN(n4871) );
  INV_X1 U6334 ( .A(SI_1_), .ZN(n4870) );
  MUX2_X1 U6335 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5184), .Z(n4893) );
  NAND2_X1 U6336 ( .A1(n4894), .A2(n4893), .ZN(n4873) );
  NAND2_X1 U6337 ( .A1(n4871), .A2(SI_1_), .ZN(n4872) );
  INV_X1 U6338 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4874) );
  XNOR2_X1 U6339 ( .A(n4904), .B(n4905), .ZN(n6575) );
  NAND2_X1 U6340 ( .A1(n4954), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4877) );
  NAND2_X1 U6341 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n4910), .ZN(n4875) );
  NAND2_X1 U6342 ( .A1(n6363), .A2(n9724), .ZN(n7723) );
  INV_X1 U6343 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n4878) );
  INV_X1 U6344 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n4879) );
  NAND2_X1 U6345 ( .A1(n4935), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4880) );
  INV_X1 U6346 ( .A(n6346), .ZN(n4886) );
  NAND2_X1 U6347 ( .A1(n6567), .A2(SI_0_), .ZN(n4884) );
  XNOR2_X1 U6348 ( .A(n4884), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U6349 ( .A1(n4886), .A2(n7080), .ZN(n6847) );
  INV_X1 U6350 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4887) );
  OR2_X1 U6351 ( .A1(n5236), .A2(n4887), .ZN(n4892) );
  NAND2_X1 U6352 ( .A1(n4935), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n4891) );
  INV_X1 U6353 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n4888) );
  OR2_X1 U6354 ( .A1(n4940), .A2(n4888), .ZN(n4890) );
  NAND4_X2 U6355 ( .A1(n4892), .A2(n4891), .A3(n4890), .A4(n4889), .ZN(n6335)
         );
  XNOR2_X1 U6356 ( .A(n4894), .B(n4893), .ZN(n6568) );
  NAND2_X1 U6357 ( .A1(n4954), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4895) );
  NAND2_X1 U6358 ( .A1(n6775), .A2(n6851), .ZN(n4896) );
  NAND2_X1 U6359 ( .A1(n6847), .A2(n4896), .ZN(n7725) );
  INV_X1 U6360 ( .A(n6851), .ZN(n6930) );
  NAND2_X1 U6361 ( .A1(n6335), .A2(n6930), .ZN(n7722) );
  NAND2_X1 U6362 ( .A1(n7725), .A2(n7722), .ZN(n7215) );
  INV_X1 U6363 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n4897) );
  OR2_X1 U6364 ( .A1(n5236), .A2(n4897), .ZN(n4899) );
  NAND2_X1 U6365 ( .A1(n4934), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n4898) );
  AND2_X1 U6366 ( .A1(n4899), .A2(n4898), .ZN(n4903) );
  INV_X1 U6367 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4900) );
  OR2_X1 U6368 ( .A1(n4940), .A2(n4900), .ZN(n4902) );
  INV_X1 U6369 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U6370 ( .A1(n4935), .A2(n9706), .ZN(n4901) );
  INV_X1 U6371 ( .A(n4906), .ZN(n4907) );
  NAND2_X1 U6372 ( .A1(n4907), .A2(SI_2_), .ZN(n4908) );
  NAND2_X1 U6373 ( .A1(n4909), .A2(n4908), .ZN(n4920) );
  INV_X1 U6374 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U6375 ( .A(n6571), .B(n6564), .S(n5184), .Z(n4921) );
  XNOR2_X1 U6376 ( .A(n4920), .B(n4919), .ZN(n6570) );
  NAND2_X1 U6377 ( .A1(n4954), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4913) );
  OAI21_X1 U6378 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(n4910), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n4911) );
  XNOR2_X1 U6379 ( .A(n4911), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6642) );
  NAND2_X1 U6380 ( .A1(n5255), .A2(n6642), .ZN(n4912) );
  OAI21_X1 U6381 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n4938), .ZN(n7207) );
  NAND2_X1 U6382 ( .A1(n5420), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n4915) );
  NAND2_X1 U6383 ( .A1(n4934), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4914) );
  INV_X1 U6384 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7208) );
  OR2_X1 U6385 ( .A1(n7683), .A2(n7208), .ZN(n4916) );
  NAND2_X1 U6386 ( .A1(n4920), .A2(n4919), .ZN(n4924) );
  INV_X1 U6387 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6388 ( .A1(n4922), .A2(SI_3_), .ZN(n4923) );
  NAND2_X1 U6389 ( .A1(n4924), .A2(n4923), .ZN(n4948) );
  MUX2_X1 U6390 ( .A(n6573), .B(n4925), .S(n5184), .Z(n4949) );
  XNOR2_X1 U6391 ( .A(n4948), .B(n4947), .ZN(n6572) );
  NAND2_X1 U6392 ( .A1(n4954), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n4929) );
  INV_X1 U6393 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9406) );
  OR2_X1 U6394 ( .A1(n4926), .A2(n9406), .ZN(n4927) );
  XNOR2_X1 U6395 ( .A(n4927), .B(P1_IR_REG_4__SCAN_IN), .ZN(n9600) );
  NAND2_X1 U6396 ( .A1(n5255), .A2(n9600), .ZN(n4928) );
  OAI211_X1 U6397 ( .C1(n4977), .C2(n6572), .A(n4929), .B(n4928), .ZN(n7210)
         );
  NAND2_X1 U6398 ( .A1(n9699), .A2(n7210), .ZN(n7729) );
  AND2_X1 U6399 ( .A1(n7799), .A2(n7729), .ZN(n4930) );
  INV_X1 U6400 ( .A(n7729), .ZN(n4931) );
  INV_X1 U6401 ( .A(n7210), .ZN(n9735) );
  NAND2_X1 U6402 ( .A1(n8869), .A2(n9735), .ZN(n7800) );
  AND2_X1 U6403 ( .A1(n7800), .A2(n7197), .ZN(n7798) );
  OR2_X1 U6404 ( .A1(n4931), .A2(n7798), .ZN(n4932) );
  NAND2_X1 U6405 ( .A1(n4267), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4946) );
  INV_X1 U6406 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6407 ( .A1(n4938), .A2(n4937), .ZN(n4939) );
  AND2_X1 U6408 ( .A1(n4998), .A2(n4939), .ZN(n7187) );
  NAND2_X1 U6409 ( .A1(n4935), .A2(n7187), .ZN(n4945) );
  INV_X1 U6410 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n4941) );
  OR2_X1 U6411 ( .A1(n7680), .A2(n4941), .ZN(n4944) );
  INV_X1 U6412 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n4942) );
  OR2_X1 U6413 ( .A1(n5236), .A2(n4942), .ZN(n4943) );
  NAND2_X1 U6414 ( .A1(n4948), .A2(n4947), .ZN(n4952) );
  INV_X1 U6415 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6416 ( .A1(n4950), .A2(SI_4_), .ZN(n4951) );
  INV_X1 U6417 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n4953) );
  MUX2_X1 U6418 ( .A(n6579), .B(n4953), .S(n5184), .Z(n4973) );
  XNOR2_X1 U6419 ( .A(n4972), .B(n4971), .ZN(n6578) );
  NAND2_X1 U6420 ( .A1(n4954), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4960) );
  NAND2_X1 U6421 ( .A1(n4955), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4956) );
  MUX2_X1 U6422 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4956), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n4958) );
  AND2_X1 U6423 ( .A1(n4958), .A2(n4957), .ZN(n6657) );
  NAND2_X1 U6424 ( .A1(n5255), .A2(n6657), .ZN(n4959) );
  OAI211_X1 U6425 ( .C1(n4977), .C2(n6578), .A(n4960), .B(n4959), .ZN(n6397)
         );
  INV_X1 U6426 ( .A(n6397), .ZN(n9745) );
  NAND2_X1 U6427 ( .A1(n8868), .A2(n9745), .ZN(n7732) );
  INV_X1 U6428 ( .A(n8868), .ZN(n4961) );
  NAND2_X1 U6429 ( .A1(n4961), .A2(n6397), .ZN(n7728) );
  NAND2_X1 U6430 ( .A1(n4267), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n4966) );
  XNOR2_X1 U6431 ( .A(n4998), .B(P1_REG3_REG_6__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U6432 ( .A1(n4935), .A2(n8819), .ZN(n4965) );
  INV_X1 U6433 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n4962) );
  OR2_X1 U6434 ( .A1(n7680), .A2(n4962), .ZN(n4964) );
  INV_X1 U6435 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6645) );
  OR2_X1 U6436 ( .A1(n7683), .A2(n6645), .ZN(n4963) );
  NAND4_X1 U6437 ( .A1(n4966), .A2(n4965), .A3(n4964), .A4(n4963), .ZN(n8867)
         );
  NAND2_X1 U6438 ( .A1(n4957), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4968) );
  MUX2_X1 U6439 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4968), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n4970) );
  INV_X1 U6440 ( .A(n4989), .ZN(n4969) );
  NAND2_X1 U6441 ( .A1(n4970), .A2(n4969), .ZN(n6644) );
  NAND2_X1 U6442 ( .A1(n4972), .A2(n4971), .ZN(n4976) );
  INV_X1 U6443 ( .A(n4973), .ZN(n4974) );
  NAND2_X1 U6444 ( .A1(n4974), .A2(SI_5_), .ZN(n4975) );
  MUX2_X1 U6445 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n5184), .Z(n4984) );
  XNOR2_X1 U6446 ( .A(n4983), .B(n4981), .ZN(n6583) );
  NAND2_X1 U6447 ( .A1(n6583), .A2(n4672), .ZN(n4979) );
  NAND2_X1 U6448 ( .A1(n5435), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4978) );
  OAI211_X1 U6449 ( .C1(n4967), .C2(n6644), .A(n4979), .B(n4978), .ZN(n8817)
         );
  NAND2_X1 U6450 ( .A1(n8867), .A2(n9748), .ZN(n7828) );
  NAND2_X1 U6451 ( .A1(n7831), .A2(n7828), .ZN(n5501) );
  NAND2_X1 U6452 ( .A1(n4983), .A2(n4982), .ZN(n4986) );
  NAND2_X1 U6453 ( .A1(n4984), .A2(SI_6_), .ZN(n4985) );
  MUX2_X1 U6454 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5184), .Z(n5008) );
  NAND2_X1 U6455 ( .A1(n4361), .A2(n7684), .ZN(n4993) );
  INV_X2 U6456 ( .A(n5015), .ZN(n5435) );
  NOR2_X1 U6457 ( .A1(n4989), .A2(n9406), .ZN(n4987) );
  MUX2_X1 U6458 ( .A(n9406), .B(n4987), .S(P1_IR_REG_7__SCAN_IN), .Z(n4991) );
  INV_X1 U6459 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U6460 ( .A1(n4989), .A2(n4988), .ZN(n5036) );
  INV_X1 U6461 ( .A(n5036), .ZN(n4990) );
  AOI22_X1 U6462 ( .A1(n5435), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5255), .B2(
        n6996), .ZN(n4992) );
  INV_X1 U6463 ( .A(n7130), .ZN(n9755) );
  NAND2_X1 U6464 ( .A1(n4267), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5004) );
  INV_X1 U6465 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n4997) );
  INV_X1 U6466 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n4996) );
  OAI21_X1 U6467 ( .B1(n4998), .B2(n4997), .A(n4996), .ZN(n4999) );
  AND2_X1 U6468 ( .A1(n5020), .A2(n4999), .ZN(n7124) );
  NAND2_X1 U6469 ( .A1(n4935), .A2(n7124), .ZN(n5003) );
  INV_X1 U6470 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5000) );
  OR2_X1 U6471 ( .A1(n7680), .A2(n5000), .ZN(n5002) );
  INV_X1 U6472 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7126) );
  OR2_X1 U6473 ( .A1(n7683), .A2(n7126), .ZN(n5001) );
  NAND4_X1 U6474 ( .A1(n5004), .A2(n5003), .A3(n5002), .A4(n5001), .ZN(n8866)
         );
  NAND2_X1 U6475 ( .A1(n9755), .A2(n8866), .ZN(n7833) );
  NAND2_X1 U6476 ( .A1(n7292), .A2(n7130), .ZN(n7830) );
  NAND2_X1 U6477 ( .A1(n5007), .A2(n5006), .ZN(n5010) );
  NAND2_X1 U6478 ( .A1(n5008), .A2(SI_7_), .ZN(n5009) );
  NAND2_X2 U6479 ( .A1(n5010), .A2(n5009), .ZN(n5030) );
  MUX2_X1 U6480 ( .A(n6611), .B(n6609), .S(n5184), .Z(n5012) );
  INV_X1 U6481 ( .A(SI_8_), .ZN(n5011) );
  INV_X1 U6482 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6483 ( .A1(n5013), .A2(SI_8_), .ZN(n5014) );
  XNOR2_X1 U6484 ( .A(n5030), .B(n5029), .ZN(n6608) );
  NAND2_X1 U6485 ( .A1(n6608), .A2(n7684), .ZN(n5018) );
  NAND2_X1 U6486 ( .A1(n5036), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5016) );
  XNOR2_X1 U6487 ( .A(n5016), .B(P1_IR_REG_8__SCAN_IN), .ZN(n8880) );
  AOI22_X1 U6488 ( .A1(n5435), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5255), .B2(
        n8880), .ZN(n5017) );
  INV_X1 U6489 ( .A(n7313), .ZN(n7155) );
  NAND2_X1 U6490 ( .A1(n4267), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5027) );
  INV_X1 U6491 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U6492 ( .A1(n5020), .A2(n9321), .ZN(n5021) );
  AND2_X1 U6493 ( .A1(n5042), .A2(n5021), .ZN(n7156) );
  NAND2_X1 U6494 ( .A1(n4935), .A2(n7156), .ZN(n5026) );
  INV_X1 U6495 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5022) );
  OR2_X1 U6496 ( .A1(n7680), .A2(n5022), .ZN(n5025) );
  INV_X1 U6497 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5023) );
  OR2_X1 U6498 ( .A1(n7683), .A2(n5023), .ZN(n5024) );
  NAND4_X1 U6499 ( .A1(n5027), .A2(n5026), .A3(n5025), .A4(n5024), .ZN(n8865)
         );
  NAND2_X1 U6500 ( .A1(n7155), .A2(n8865), .ZN(n7706) );
  INV_X1 U6501 ( .A(n8865), .ZN(n9676) );
  INV_X1 U6502 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5032) );
  INV_X1 U6503 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5031) );
  MUX2_X1 U6504 ( .A(n5032), .B(n5031), .S(n5184), .Z(n5033) );
  INV_X1 U6505 ( .A(n5033), .ZN(n5034) );
  NAND2_X1 U6506 ( .A1(n5034), .A2(SI_9_), .ZN(n5035) );
  NAND2_X1 U6507 ( .A1(n6616), .A2(n7684), .ZN(n5040) );
  NAND2_X1 U6508 ( .A1(n5037), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5038) );
  XNOR2_X1 U6509 ( .A(n5038), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U6510 ( .A1(n5435), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5255), .B2(
        n9620), .ZN(n5039) );
  NAND2_X1 U6511 ( .A1(n4267), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5048) );
  NAND2_X1 U6512 ( .A1(n5042), .A2(n5041), .ZN(n5043) );
  AND2_X1 U6513 ( .A1(n5065), .A2(n5043), .ZN(n9681) );
  NAND2_X1 U6514 ( .A1(n4935), .A2(n9681), .ZN(n5047) );
  INV_X1 U6515 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5044) );
  OR2_X1 U6516 ( .A1(n7680), .A2(n5044), .ZN(n5046) );
  INV_X1 U6517 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6999) );
  OR2_X1 U6518 ( .A1(n7683), .A2(n6999), .ZN(n5045) );
  NAND4_X1 U6519 ( .A1(n5048), .A2(n5047), .A3(n5046), .A4(n5045), .ZN(n8864)
         );
  INV_X1 U6520 ( .A(n8864), .ZN(n7704) );
  OR2_X1 U6521 ( .A1(n7705), .A2(n7704), .ZN(n7837) );
  INV_X1 U6522 ( .A(n7298), .ZN(n5073) );
  MUX2_X1 U6523 ( .A(n6676), .B(n6665), .S(n5184), .Z(n5054) );
  INV_X1 U6524 ( .A(SI_10_), .ZN(n5053) );
  NAND2_X1 U6525 ( .A1(n5054), .A2(n5053), .ZN(n5075) );
  INV_X1 U6526 ( .A(n5054), .ZN(n5055) );
  NAND2_X1 U6527 ( .A1(n5055), .A2(SI_10_), .ZN(n5056) );
  NAND2_X1 U6528 ( .A1(n6664), .A2(n7684), .ZN(n5063) );
  NOR2_X1 U6529 ( .A1(n5099), .A2(n9406), .ZN(n5058) );
  NAND2_X1 U6530 ( .A1(n5058), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n5061) );
  INV_X1 U6531 ( .A(n5058), .ZN(n5060) );
  NAND2_X1 U6532 ( .A1(n5060), .A2(n5059), .ZN(n5077) );
  AOI22_X1 U6533 ( .A1(n5435), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5255), .B2(
        n7001), .ZN(n5062) );
  NAND2_X2 U6534 ( .A1(n5063), .A2(n5062), .ZN(n7416) );
  NAND2_X1 U6535 ( .A1(n4267), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5072) );
  INV_X1 U6536 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7429) );
  NAND2_X1 U6537 ( .A1(n5065), .A2(n7429), .ZN(n5066) );
  AND2_X1 U6538 ( .A1(n5082), .A2(n5066), .ZN(n7430) );
  NAND2_X1 U6539 ( .A1(n4935), .A2(n7430), .ZN(n5071) );
  INV_X1 U6540 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5067) );
  OR2_X1 U6541 ( .A1(n7680), .A2(n5067), .ZN(n5070) );
  INV_X1 U6542 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5068) );
  OR2_X1 U6543 ( .A1(n7683), .A2(n5068), .ZN(n5069) );
  NAND4_X1 U6544 ( .A1(n5072), .A2(n5071), .A3(n5070), .A4(n5069), .ZN(n8863)
         );
  INV_X1 U6545 ( .A(n8863), .ZN(n9675) );
  NAND2_X1 U6546 ( .A1(n7416), .A2(n9675), .ZN(n7847) );
  MUX2_X1 U6547 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n5184), .Z(n5091) );
  INV_X1 U6548 ( .A(SI_11_), .ZN(n5076) );
  XNOR2_X1 U6549 ( .A(n5093), .B(n5090), .ZN(n6666) );
  NAND2_X1 U6550 ( .A1(n6666), .A2(n7684), .ZN(n5080) );
  NAND2_X1 U6551 ( .A1(n5077), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U6552 ( .A(n5078), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9640) );
  AOI22_X1 U6553 ( .A1(n5435), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5255), .B2(
        n9640), .ZN(n5079) );
  NAND2_X1 U6554 ( .A1(n4267), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n5089) );
  INV_X1 U6555 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U6556 ( .A1(n5082), .A2(n5081), .ZN(n5083) );
  AND2_X1 U6557 ( .A1(n5105), .A2(n5083), .ZN(n9516) );
  NAND2_X1 U6558 ( .A1(n4935), .A2(n9516), .ZN(n5088) );
  INV_X1 U6559 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6560 ( .A1(n7680), .A2(n5084), .ZN(n5087) );
  INV_X1 U6561 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5085) );
  OR2_X1 U6562 ( .A1(n5236), .A2(n5085), .ZN(n5086) );
  NAND4_X1 U6563 ( .A1(n5089), .A2(n5088), .A3(n5087), .A4(n5086), .ZN(n8862)
         );
  AND2_X1 U6564 ( .A1(n7459), .A2(n7499), .ZN(n7760) );
  OR2_X1 U6565 ( .A1(n7459), .A2(n7499), .ZN(n7761) );
  INV_X1 U6566 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6681) );
  INV_X1 U6567 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6683) );
  MUX2_X1 U6568 ( .A(n6681), .B(n6683), .S(n5184), .Z(n5095) );
  INV_X1 U6569 ( .A(SI_12_), .ZN(n5094) );
  INV_X1 U6570 ( .A(n5095), .ZN(n5096) );
  NAND2_X1 U6571 ( .A1(n5096), .A2(SI_12_), .ZN(n5097) );
  XNOR2_X1 U6572 ( .A(n5114), .B(n5113), .ZN(n6680) );
  NAND2_X1 U6573 ( .A1(n6680), .A2(n7684), .ZN(n5102) );
  NOR2_X1 U6574 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5098) );
  NAND2_X1 U6575 ( .A1(n5099), .A2(n5098), .ZN(n5120) );
  NAND2_X1 U6576 ( .A1(n5120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5100) );
  XNOR2_X1 U6577 ( .A(n5100), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7524) );
  AOI22_X1 U6578 ( .A1(n5435), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5255), .B2(
        n7524), .ZN(n5101) );
  INV_X1 U6579 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6580 ( .A1(n5105), .A2(n5104), .ZN(n5106) );
  AND2_X1 U6581 ( .A1(n5126), .A2(n5106), .ZN(n7503) );
  NAND2_X1 U6582 ( .A1(n4935), .A2(n7503), .ZN(n5111) );
  NAND2_X1 U6583 ( .A1(n4267), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n5110) );
  INV_X1 U6584 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7516) );
  OR2_X1 U6585 ( .A1(n7683), .A2(n7516), .ZN(n5109) );
  INV_X1 U6586 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5107) );
  OR2_X1 U6587 ( .A1(n7680), .A2(n5107), .ZN(n5108) );
  NAND4_X1 U6588 ( .A1(n5111), .A2(n5110), .A3(n5109), .A4(n5108), .ZN(n8861)
         );
  NOR2_X1 U6589 ( .A1(n7507), .A2(n9511), .ZN(n7712) );
  NAND2_X1 U6590 ( .A1(n7507), .A2(n9511), .ZN(n7860) );
  INV_X1 U6591 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6703) );
  INV_X1 U6592 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5115) );
  MUX2_X1 U6593 ( .A(n6703), .B(n5115), .S(n5184), .Z(n5117) );
  INV_X1 U6594 ( .A(SI_13_), .ZN(n5116) );
  NAND2_X1 U6595 ( .A1(n5117), .A2(n5116), .ZN(n5136) );
  INV_X1 U6596 ( .A(n5117), .ZN(n5118) );
  NAND2_X1 U6597 ( .A1(n5118), .A2(SI_13_), .ZN(n5119) );
  NAND2_X1 U6598 ( .A1(n6684), .A2(n7684), .ZN(n5124) );
  INV_X1 U6599 ( .A(n5139), .ZN(n5121) );
  NAND2_X1 U6600 ( .A1(n5121), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U6601 ( .A(n5122), .B(P1_IR_REG_13__SCAN_IN), .ZN(n8887) );
  AOI22_X1 U6602 ( .A1(n5435), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5255), .B2(
        n8887), .ZN(n5123) );
  NAND2_X1 U6603 ( .A1(n4267), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5133) );
  INV_X1 U6604 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5125) );
  NAND2_X1 U6605 ( .A1(n5126), .A2(n5125), .ZN(n5127) );
  AND2_X1 U6606 ( .A1(n5146), .A2(n5127), .ZN(n9500) );
  NAND2_X1 U6607 ( .A1(n4935), .A2(n9500), .ZN(n5132) );
  INV_X1 U6608 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5128) );
  OR2_X1 U6609 ( .A1(n7680), .A2(n5128), .ZN(n5131) );
  INV_X1 U6610 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n5129) );
  OR2_X1 U6611 ( .A1(n7683), .A2(n5129), .ZN(n5130) );
  NAND4_X1 U6612 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n8860)
         );
  XNOR2_X1 U6613 ( .A(n9486), .B(n8860), .ZN(n9493) );
  INV_X1 U6614 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6791) );
  INV_X1 U6615 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6757) );
  MUX2_X1 U6616 ( .A(n6791), .B(n6757), .S(n5184), .Z(n5155) );
  NAND2_X1 U6617 ( .A1(n6756), .A2(n7684), .ZN(n5145) );
  NOR2_X1 U6618 ( .A1(n5190), .A2(n9406), .ZN(n5140) );
  NAND2_X1 U6619 ( .A1(n5140), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5143) );
  INV_X1 U6620 ( .A(n5140), .ZN(n5142) );
  INV_X1 U6621 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6622 ( .A1(n5142), .A2(n5141), .ZN(n5164) );
  AND2_X1 U6623 ( .A1(n5143), .A2(n5164), .ZN(n9653) );
  AOI22_X1 U6624 ( .A1(n9653), .A2(n5255), .B1(n5435), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n5144) );
  NAND2_X1 U6625 ( .A1(n4267), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n5152) );
  INV_X1 U6626 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U6627 ( .A1(n5146), .A2(n7670), .ZN(n5147) );
  AND2_X1 U6628 ( .A1(n5172), .A2(n5147), .ZN(n7538) );
  NAND2_X1 U6629 ( .A1(n4935), .A2(n7538), .ZN(n5151) );
  INV_X1 U6630 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7539) );
  OR2_X1 U6631 ( .A1(n7683), .A2(n7539), .ZN(n5150) );
  INV_X1 U6632 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5148) );
  OR2_X1 U6633 ( .A1(n7680), .A2(n5148), .ZN(n5149) );
  NAND4_X1 U6634 ( .A1(n5152), .A2(n5151), .A3(n5150), .A4(n5149), .ZN(n8859)
         );
  INV_X1 U6635 ( .A(n8859), .ZN(n9495) );
  NAND2_X1 U6636 ( .A1(n7673), .A2(n9495), .ZN(n7863) );
  INV_X1 U6637 ( .A(n8860), .ZN(n7708) );
  AND2_X1 U6638 ( .A1(n9486), .A2(n7708), .ZN(n7856) );
  NOR2_X1 U6639 ( .A1(n7776), .A2(n7856), .ZN(n5153) );
  INV_X1 U6640 ( .A(n5155), .ZN(n5156) );
  NAND2_X1 U6641 ( .A1(n5156), .A2(SI_14_), .ZN(n5157) );
  INV_X1 U6642 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6886) );
  INV_X1 U6643 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6884) );
  MUX2_X1 U6644 ( .A(n6886), .B(n6884), .S(n5184), .Z(n5161) );
  INV_X1 U6645 ( .A(SI_15_), .ZN(n5160) );
  INV_X1 U6646 ( .A(n5161), .ZN(n5162) );
  NAND2_X1 U6647 ( .A1(n5162), .A2(SI_15_), .ZN(n5163) );
  XNOR2_X1 U6648 ( .A(n5183), .B(n5182), .ZN(n6883) );
  NAND2_X1 U6649 ( .A1(n6883), .A2(n7684), .ZN(n5169) );
  NAND2_X1 U6650 ( .A1(n5164), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5166) );
  INV_X1 U6651 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U6652 ( .A(n5166), .B(n5165), .ZN(n8905) );
  OAI22_X1 U6653 ( .A1(n8905), .A2(n4967), .B1(n5015), .B2(n6884), .ZN(n5167)
         );
  INV_X1 U6654 ( .A(n5167), .ZN(n5168) );
  NAND2_X1 U6655 ( .A1(n4267), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5179) );
  INV_X1 U6656 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6657 ( .A1(n5172), .A2(n5171), .ZN(n5173) );
  AND2_X1 U6658 ( .A1(n5195), .A2(n5173), .ZN(n8845) );
  NAND2_X1 U6659 ( .A1(n4935), .A2(n8845), .ZN(n5178) );
  INV_X1 U6660 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5174) );
  OR2_X1 U6661 ( .A1(n7680), .A2(n5174), .ZN(n5177) );
  INV_X1 U6662 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n5175) );
  OR2_X1 U6663 ( .A1(n5236), .A2(n5175), .ZN(n5176) );
  NAND4_X1 U6664 ( .A1(n5179), .A2(n5178), .A3(n5177), .A4(n5176), .ZN(n8858)
         );
  INV_X1 U6665 ( .A(n8858), .ZN(n8757) );
  OR2_X1 U6666 ( .A1(n8851), .A2(n8757), .ZN(n7718) );
  NAND2_X1 U6667 ( .A1(n8851), .A2(n8757), .ZN(n7701) );
  NAND2_X1 U6668 ( .A1(n7718), .A2(n7701), .ZN(n7631) );
  NAND2_X1 U6669 ( .A1(n5180), .A2(n7870), .ZN(n7634) );
  INV_X1 U6670 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6926) );
  INV_X1 U6671 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6941) );
  MUX2_X1 U6672 ( .A(n6926), .B(n6941), .S(n5184), .Z(n5186) );
  INV_X1 U6673 ( .A(SI_16_), .ZN(n5185) );
  NAND2_X1 U6674 ( .A1(n5186), .A2(n5185), .ZN(n5205) );
  INV_X1 U6675 ( .A(n5186), .ZN(n5187) );
  NAND2_X1 U6676 ( .A1(n5187), .A2(SI_16_), .ZN(n5188) );
  XNOR2_X1 U6677 ( .A(n5204), .B(n5203), .ZN(n6925) );
  NAND2_X1 U6678 ( .A1(n6925), .A2(n7684), .ZN(n5193) );
  NOR2_X1 U6679 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5189) );
  NAND2_X1 U6680 ( .A1(n5190), .A2(n5189), .ZN(n5207) );
  NAND2_X1 U6681 ( .A1(n5207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5191) );
  XNOR2_X1 U6682 ( .A(n5191), .B(P1_IR_REG_16__SCAN_IN), .ZN(n8921) );
  AOI22_X1 U6683 ( .A1(n8921), .A2(n5255), .B1(n5435), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5192) );
  NAND2_X1 U6684 ( .A1(n4267), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5202) );
  INV_X1 U6685 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U6686 ( .A1(n5195), .A2(n8756), .ZN(n5196) );
  AND2_X1 U6687 ( .A1(n5213), .A2(n5196), .ZN(n8758) );
  NAND2_X1 U6688 ( .A1(n4935), .A2(n8758), .ZN(n5201) );
  INV_X1 U6689 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5197) );
  OR2_X1 U6690 ( .A1(n7680), .A2(n5197), .ZN(n5200) );
  INV_X1 U6691 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n5198) );
  OR2_X1 U6692 ( .A1(n5236), .A2(n5198), .ZN(n5199) );
  NAND4_X1 U6693 ( .A1(n5202), .A2(n5201), .A3(n5200), .A4(n5199), .ZN(n8857)
         );
  INV_X1 U6694 ( .A(n8857), .ZN(n9165) );
  AND2_X1 U6695 ( .A1(n8762), .A2(n9165), .ZN(n5517) );
  INV_X1 U6696 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6963) );
  INV_X1 U6697 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9359) );
  MUX2_X1 U6698 ( .A(n6963), .B(n9359), .S(n6567), .Z(n5223) );
  XNOR2_X1 U6699 ( .A(n5223), .B(SI_17_), .ZN(n5220) );
  XNOR2_X1 U6700 ( .A(n5222), .B(n5220), .ZN(n6962) );
  NAND2_X1 U6701 ( .A1(n6962), .A2(n7684), .ZN(n5211) );
  NAND2_X1 U6702 ( .A1(n5253), .A2(n5208), .ZN(n5226) );
  OR2_X1 U6703 ( .A1(n5253), .A2(n5208), .ZN(n5209) );
  AOI22_X1 U6704 ( .A1(n8939), .A2(n5255), .B1(n5435), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6705 ( .A1(n4267), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n5219) );
  INV_X1 U6706 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5212) );
  NAND2_X1 U6707 ( .A1(n5213), .A2(n5212), .ZN(n5214) );
  AND2_X1 U6708 ( .A1(n5233), .A2(n5214), .ZN(n9171) );
  NAND2_X1 U6709 ( .A1(n4935), .A2(n9171), .ZN(n5218) );
  INV_X1 U6710 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9362) );
  OR2_X1 U6711 ( .A1(n7680), .A2(n9362), .ZN(n5217) );
  INV_X1 U6712 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5215) );
  OR2_X1 U6713 ( .A1(n7683), .A2(n5215), .ZN(n5216) );
  NAND4_X1 U6714 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n9155)
         );
  OR2_X1 U6715 ( .A1(n9243), .A2(n9155), .ZN(n5519) );
  NAND2_X1 U6716 ( .A1(n9243), .A2(n9155), .ZN(n7881) );
  NAND2_X1 U6717 ( .A1(n5519), .A2(n7881), .ZN(n9161) );
  INV_X1 U6718 ( .A(n9155), .ZN(n8806) );
  OR2_X1 U6719 ( .A1(n9243), .A2(n8806), .ZN(n7692) );
  INV_X1 U6720 ( .A(n5220), .ZN(n5221) );
  INV_X1 U6721 ( .A(n5223), .ZN(n5224) );
  NAND2_X1 U6722 ( .A1(n5224), .A2(SI_17_), .ZN(n5225) );
  MUX2_X1 U6723 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6567), .Z(n5245) );
  XNOR2_X1 U6724 ( .A(n5245), .B(SI_18_), .ZN(n5242) );
  XNOR2_X1 U6725 ( .A(n5244), .B(n5242), .ZN(n7084) );
  NAND2_X1 U6726 ( .A1(n7084), .A2(n7684), .ZN(n5230) );
  NAND2_X1 U6727 ( .A1(n5226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5227) );
  XNOR2_X1 U6728 ( .A(n5227), .B(P1_IR_REG_18__SCAN_IN), .ZN(n8950) );
  INV_X1 U6729 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9380) );
  NOR2_X1 U6730 ( .A1(n5015), .A2(n9380), .ZN(n5228) );
  AOI21_X1 U6731 ( .B1(n8950), .B2(n5255), .A(n5228), .ZN(n5229) );
  INV_X1 U6732 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8805) );
  NAND2_X1 U6733 ( .A1(n5233), .A2(n8805), .ZN(n5234) );
  NAND2_X1 U6734 ( .A1(n5259), .A2(n5234), .ZN(n9145) );
  OR2_X1 U6735 ( .A1(n5231), .A2(n9145), .ZN(n5240) );
  NAND2_X1 U6736 ( .A1(n5420), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5239) );
  NAND2_X1 U6737 ( .A1(n4267), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5238) );
  INV_X1 U6738 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5235) );
  OR2_X1 U6739 ( .A1(n5236), .A2(n5235), .ZN(n5237) );
  NAND4_X1 U6740 ( .A1(n5240), .A2(n5239), .A3(n5238), .A4(n5237), .ZN(n9138)
         );
  INV_X1 U6741 ( .A(n9138), .ZN(n9166) );
  OR2_X1 U6742 ( .A1(n9236), .A2(n9166), .ZN(n7885) );
  NAND2_X1 U6743 ( .A1(n9236), .A2(n9166), .ZN(n7892) );
  NAND2_X1 U6744 ( .A1(n7885), .A2(n7892), .ZN(n9149) );
  INV_X1 U6745 ( .A(n5242), .ZN(n5243) );
  INV_X1 U6746 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7166) );
  INV_X1 U6747 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n5246) );
  MUX2_X1 U6748 ( .A(n7166), .B(n5246), .S(n6567), .Z(n5248) );
  INV_X1 U6749 ( .A(SI_19_), .ZN(n5247) );
  NAND2_X1 U6750 ( .A1(n5248), .A2(n5247), .ZN(n5265) );
  INV_X1 U6751 ( .A(n5248), .ZN(n5249) );
  NAND2_X1 U6752 ( .A1(n5249), .A2(SI_19_), .ZN(n5250) );
  NAND2_X1 U6753 ( .A1(n5265), .A2(n5250), .ZN(n5266) );
  XNOR2_X1 U6754 ( .A(n5267), .B(n5266), .ZN(n7107) );
  NAND2_X1 U6755 ( .A1(n7107), .A2(n7684), .ZN(n5257) );
  NAND2_X1 U6756 ( .A1(n5251), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5252) );
  AOI22_X1 U6757 ( .A1(n7953), .A2(n5255), .B1(P2_DATAO_REG_19__SCAN_IN), .B2(
        n5435), .ZN(n5256) );
  INV_X1 U6758 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6759 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  NAND2_X1 U6760 ( .A1(n5277), .A2(n5260), .ZN(n9130) );
  NAND2_X1 U6761 ( .A1(n4267), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n5262) );
  NAND2_X1 U6762 ( .A1(n5420), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5261) );
  AND2_X1 U6763 ( .A1(n5262), .A2(n5261), .ZN(n5264) );
  INV_X1 U6764 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8947) );
  OR2_X1 U6765 ( .A1(n7683), .A2(n8947), .ZN(n5263) );
  OAI211_X1 U6766 ( .C1(n9130), .C2(n5231), .A(n5264), .B(n5263), .ZN(n9153)
         );
  INV_X1 U6767 ( .A(n9153), .ZN(n8808) );
  OR2_X1 U6768 ( .A1(n9232), .A2(n8808), .ZN(n7896) );
  NAND2_X1 U6769 ( .A1(n9232), .A2(n8808), .ZN(n7891) );
  INV_X1 U6770 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7311) );
  INV_X1 U6771 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n5268) );
  MUX2_X1 U6772 ( .A(n7311), .B(n5268), .S(n6567), .Z(n5270) );
  INV_X1 U6773 ( .A(SI_20_), .ZN(n5269) );
  NAND2_X1 U6774 ( .A1(n5270), .A2(n5269), .ZN(n5283) );
  INV_X1 U6775 ( .A(n5270), .ZN(n5271) );
  NAND2_X1 U6776 ( .A1(n5271), .A2(SI_20_), .ZN(n5272) );
  XNOR2_X1 U6777 ( .A(n5282), .B(n5281), .ZN(n7229) );
  NAND2_X1 U6778 ( .A1(n7229), .A2(n7684), .ZN(n5274) );
  NAND2_X1 U6779 ( .A1(n4954), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5273) );
  INV_X1 U6780 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n9360) );
  INV_X1 U6781 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6782 ( .A1(n5277), .A2(n5276), .ZN(n5278) );
  NAND2_X1 U6783 ( .A1(n5287), .A2(n5278), .ZN(n8785) );
  OR2_X1 U6784 ( .A1(n8785), .A2(n5231), .ZN(n5280) );
  AOI22_X1 U6785 ( .A1(n4267), .A2(P1_REG1_REG_20__SCAN_IN), .B1(n5419), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n5279) );
  OAI211_X1 U6786 ( .C1(n7680), .C2(n9360), .A(n5280), .B(n5279), .ZN(n9137)
         );
  INV_X1 U6787 ( .A(n9137), .ZN(n9099) );
  XNOR2_X1 U6788 ( .A(n9226), .B(n9099), .ZN(n9111) );
  INV_X1 U6789 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7374) );
  INV_X1 U6790 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n5284) );
  MUX2_X1 U6791 ( .A(n7374), .B(n5284), .S(n6567), .Z(n5293) );
  XNOR2_X1 U6792 ( .A(n5293), .B(SI_21_), .ZN(n5292) );
  NAND2_X1 U6793 ( .A1(n7335), .A2(n7684), .ZN(n5286) );
  NAND2_X1 U6794 ( .A1(n5435), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5285) );
  NAND2_X2 U6795 ( .A1(n5286), .A2(n5285), .ZN(n9223) );
  INV_X1 U6796 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U6797 ( .A1(n5287), .A2(n8737), .ZN(n5288) );
  NAND2_X1 U6798 ( .A1(n5305), .A2(n5288), .ZN(n9104) );
  AOI22_X1 U6799 ( .A1(n4267), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n5419), .B2(
        P1_REG2_REG_21__SCAN_IN), .ZN(n5290) );
  NAND2_X1 U6800 ( .A1(n5420), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5289) );
  OAI211_X1 U6801 ( .C1(n9104), .C2(n5231), .A(n5290), .B(n5289), .ZN(n9121)
         );
  INV_X1 U6802 ( .A(n9121), .ZN(n8795) );
  NAND2_X1 U6803 ( .A1(n9223), .A2(n8795), .ZN(n9085) );
  INV_X1 U6804 ( .A(n5293), .ZN(n5294) );
  NAND2_X1 U6805 ( .A1(n5294), .A2(SI_21_), .ZN(n5295) );
  INV_X1 U6806 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7413) );
  INV_X1 U6807 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n5297) );
  MUX2_X1 U6808 ( .A(n7413), .B(n5297), .S(n6567), .Z(n5299) );
  INV_X1 U6809 ( .A(SI_22_), .ZN(n5298) );
  NAND2_X1 U6810 ( .A1(n5299), .A2(n5298), .ZN(n5313) );
  INV_X1 U6811 ( .A(n5299), .ZN(n5300) );
  NAND2_X1 U6812 ( .A1(n5300), .A2(SI_22_), .ZN(n5301) );
  NAND2_X1 U6813 ( .A1(n5313), .A2(n5301), .ZN(n5314) );
  NAND2_X1 U6814 ( .A1(n7392), .A2(n7684), .ZN(n5303) );
  NAND2_X1 U6815 ( .A1(n5435), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5302) );
  INV_X1 U6816 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9379) );
  NAND2_X1 U6817 ( .A1(n5305), .A2(n9379), .ZN(n5306) );
  NAND2_X1 U6818 ( .A1(n5324), .A2(n5306), .ZN(n9081) );
  OR2_X1 U6819 ( .A1(n9081), .A2(n5231), .ZN(n5312) );
  INV_X1 U6820 ( .A(n4267), .ZN(n5424) );
  INV_X1 U6821 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5309) );
  NAND2_X1 U6822 ( .A1(n5420), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6823 ( .A1(n5419), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5307) );
  OAI211_X1 U6824 ( .C1(n5424), .C2(n5309), .A(n5308), .B(n5307), .ZN(n5310)
         );
  INV_X1 U6825 ( .A(n5310), .ZN(n5311) );
  NAND2_X1 U6826 ( .A1(n5312), .A2(n5311), .ZN(n9071) );
  INV_X1 U6827 ( .A(n9071), .ZN(n9100) );
  NAND2_X1 U6828 ( .A1(n9216), .A2(n9100), .ZN(n7907) );
  INV_X1 U6829 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5316) );
  INV_X1 U6830 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9319) );
  MUX2_X1 U6831 ( .A(n5316), .B(n9319), .S(n6567), .Z(n5318) );
  INV_X1 U6832 ( .A(SI_23_), .ZN(n5317) );
  NAND2_X1 U6833 ( .A1(n5318), .A2(n5317), .ZN(n5334) );
  INV_X1 U6834 ( .A(n5318), .ZN(n5319) );
  NAND2_X1 U6835 ( .A1(n5319), .A2(SI_23_), .ZN(n5320) );
  NAND2_X1 U6836 ( .A1(n7449), .A2(n7684), .ZN(n5322) );
  NAND2_X1 U6837 ( .A1(n5435), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5321) );
  INV_X1 U6838 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8728) );
  NAND2_X1 U6839 ( .A1(n5324), .A2(n8728), .ZN(n5325) );
  NAND2_X1 U6840 ( .A1(n5340), .A2(n5325), .ZN(n9064) );
  OR2_X1 U6841 ( .A1(n9064), .A2(n5231), .ZN(n5331) );
  INV_X1 U6842 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5328) );
  NAND2_X1 U6843 ( .A1(n5420), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6844 ( .A1(n5419), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5326) );
  OAI211_X1 U6845 ( .C1(n5424), .C2(n5328), .A(n5327), .B(n5326), .ZN(n5329)
         );
  INV_X1 U6846 ( .A(n5329), .ZN(n5330) );
  INV_X1 U6847 ( .A(n9088), .ZN(n8796) );
  INV_X1 U6848 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7511) );
  INV_X1 U6849 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5336) );
  MUX2_X1 U6850 ( .A(n7511), .B(n5336), .S(n6567), .Z(n5349) );
  XNOR2_X1 U6851 ( .A(n5349), .B(SI_24_), .ZN(n5348) );
  XNOR2_X1 U6852 ( .A(n5353), .B(n5348), .ZN(n7463) );
  NAND2_X1 U6853 ( .A1(n7463), .A2(n7684), .ZN(n5338) );
  NAND2_X1 U6854 ( .A1(n5435), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5337) );
  INV_X1 U6855 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6856 ( .A1(n5340), .A2(n5339), .ZN(n5341) );
  NAND2_X1 U6857 ( .A1(n5361), .A2(n5341), .ZN(n9046) );
  INV_X1 U6858 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5344) );
  NAND2_X1 U6859 ( .A1(n5419), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6860 ( .A1(n5420), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5342) );
  OAI211_X1 U6861 ( .C1(n5424), .C2(n5344), .A(n5343), .B(n5342), .ZN(n5345)
         );
  INV_X1 U6862 ( .A(n5345), .ZN(n5346) );
  OR2_X2 U6863 ( .A1(n9050), .A2(n9042), .ZN(n9051) );
  INV_X1 U6864 ( .A(n5348), .ZN(n5352) );
  INV_X1 U6865 ( .A(n5349), .ZN(n5350) );
  NAND2_X1 U6866 ( .A1(n5350), .A2(SI_24_), .ZN(n5351) );
  INV_X1 U6867 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7584) );
  INV_X1 U6868 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5354) );
  MUX2_X1 U6869 ( .A(n7584), .B(n5354), .S(n6567), .Z(n5356) );
  INV_X1 U6870 ( .A(SI_25_), .ZN(n5355) );
  NAND2_X1 U6871 ( .A1(n5356), .A2(n5355), .ZN(n5369) );
  INV_X1 U6872 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U6873 ( .A1(n5357), .A2(SI_25_), .ZN(n5358) );
  NAND2_X1 U6874 ( .A1(n5369), .A2(n5358), .ZN(n5370) );
  NAND2_X1 U6875 ( .A1(n7567), .A2(n7684), .ZN(n5360) );
  NAND2_X1 U6876 ( .A1(n5435), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5359) );
  INV_X1 U6877 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U6878 ( .A1(n5361), .A2(n8746), .ZN(n5362) );
  NAND2_X1 U6879 ( .A1(n9035), .A2(n4935), .ZN(n5368) );
  INV_X1 U6880 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n5365) );
  NAND2_X1 U6881 ( .A1(n4267), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5364) );
  NAND2_X1 U6882 ( .A1(n5419), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5363) );
  OAI211_X1 U6883 ( .C1(n7680), .C2(n5365), .A(n5364), .B(n5363), .ZN(n5366)
         );
  INV_X1 U6884 ( .A(n5366), .ZN(n5367) );
  INV_X1 U6885 ( .A(n9054), .ZN(n5390) );
  INV_X1 U6886 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7585) );
  INV_X1 U6887 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5372) );
  MUX2_X1 U6888 ( .A(n7585), .B(n5372), .S(n6567), .Z(n5374) );
  INV_X1 U6889 ( .A(SI_26_), .ZN(n5373) );
  NAND2_X1 U6890 ( .A1(n5374), .A2(n5373), .ZN(n5395) );
  INV_X1 U6891 ( .A(n5374), .ZN(n5375) );
  NAND2_X1 U6892 ( .A1(n5375), .A2(SI_26_), .ZN(n5376) );
  AND2_X1 U6893 ( .A1(n5395), .A2(n5376), .ZN(n5393) );
  NAND2_X1 U6894 ( .A1(n5435), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5377) );
  INV_X1 U6895 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5380) );
  NAND2_X1 U6896 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  NAND2_X1 U6897 ( .A1(n5417), .A2(n5382), .ZN(n9011) );
  INV_X1 U6898 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5385) );
  NAND2_X1 U6899 ( .A1(n5419), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6900 ( .A1(n5420), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5383) );
  OAI211_X1 U6901 ( .C1(n5424), .C2(n5385), .A(n5384), .B(n5383), .ZN(n5386)
         );
  INV_X1 U6902 ( .A(n5386), .ZN(n5387) );
  NAND2_X1 U6903 ( .A1(n9196), .A2(n9031), .ZN(n7919) );
  AND2_X1 U6904 ( .A1(n9016), .A2(n7919), .ZN(n5389) );
  AND2_X1 U6905 ( .A1(n5389), .A2(n9015), .ZN(n5392) );
  INV_X1 U6906 ( .A(n7919), .ZN(n7688) );
  OR2_X1 U6907 ( .A1(n9196), .A2(n9031), .ZN(n5391) );
  INV_X1 U6908 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7664) );
  INV_X1 U6909 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5397) );
  MUX2_X1 U6910 ( .A(n7664), .B(n5397), .S(n6567), .Z(n5399) );
  INV_X1 U6911 ( .A(SI_27_), .ZN(n5398) );
  NAND2_X1 U6912 ( .A1(n5399), .A2(n5398), .ZN(n5412) );
  INV_X1 U6913 ( .A(n5399), .ZN(n5400) );
  NAND2_X1 U6914 ( .A1(n5400), .A2(SI_27_), .ZN(n5401) );
  AND2_X1 U6915 ( .A1(n5412), .A2(n5401), .ZN(n5410) );
  NAND2_X1 U6916 ( .A1(n7648), .A2(n7684), .ZN(n5403) );
  NAND2_X1 U6917 ( .A1(n5435), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5402) );
  XNOR2_X1 U6918 ( .A(n5417), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U6919 ( .A1(n8996), .A2(n4935), .ZN(n5409) );
  INV_X1 U6920 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6921 ( .A1(n5420), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6922 ( .A1(n5419), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5404) );
  OAI211_X1 U6923 ( .C1(n5424), .C2(n5406), .A(n5405), .B(n5404), .ZN(n5407)
         );
  INV_X1 U6924 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U6925 ( .A1(n9191), .A2(n8025), .ZN(n7925) );
  INV_X1 U6926 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8723) );
  INV_X1 U6927 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5413) );
  MUX2_X1 U6928 ( .A(n8723), .B(n5413), .S(n6567), .Z(n5432) );
  XNOR2_X1 U6929 ( .A(n5432), .B(SI_28_), .ZN(n5429) );
  NAND2_X1 U6930 ( .A1(n8721), .A2(n7684), .ZN(n5415) );
  NAND2_X1 U6931 ( .A1(n4954), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5414) );
  INV_X1 U6932 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5416) );
  INV_X1 U6933 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8022) );
  OAI21_X1 U6934 ( .B1(n5417), .B2(n5416), .A(n8022), .ZN(n5418) );
  NAND2_X1 U6935 ( .A1(n5418), .A2(n5539), .ZN(n8986) );
  INV_X1 U6936 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5423) );
  NAND2_X1 U6937 ( .A1(n5419), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U6938 ( .A1(n5420), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5421) );
  OAI211_X1 U6939 ( .C1(n5424), .C2(n5423), .A(n5422), .B(n5421), .ZN(n5425)
         );
  INV_X1 U6940 ( .A(n5425), .ZN(n5426) );
  INV_X1 U6941 ( .A(n7929), .ZN(n5428) );
  INV_X1 U6942 ( .A(SI_28_), .ZN(n5431) );
  INV_X1 U6943 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8718) );
  INV_X1 U6944 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n5433) );
  MUX2_X1 U6945 ( .A(n8718), .B(n5433), .S(n6567), .Z(n6143) );
  XNOR2_X1 U6946 ( .A(n6143), .B(SI_29_), .ZN(n5434) );
  NAND2_X1 U6947 ( .A1(n8717), .A2(n7684), .ZN(n5437) );
  NAND2_X1 U6948 ( .A1(n5435), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5436) );
  INV_X1 U6949 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5441) );
  NAND2_X1 U6950 ( .A1(n4267), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5440) );
  INV_X1 U6951 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n5438) );
  OR2_X1 U6952 ( .A1(n7680), .A2(n5438), .ZN(n5439) );
  OAI211_X1 U6953 ( .C1(n5441), .C2(n7683), .A(n5440), .B(n5439), .ZN(n5442)
         );
  INV_X1 U6954 ( .A(n5442), .ZN(n5443) );
  OAI21_X1 U6955 ( .B1(n5539), .B2(n5231), .A(n5443), .ZN(n8979) );
  INV_X1 U6956 ( .A(n8979), .ZN(n7938) );
  NAND2_X1 U6957 ( .A1(n9180), .A2(n7938), .ZN(n7821) );
  NAND2_X1 U6958 ( .A1(n5462), .A2(n5444), .ZN(n5445) );
  NAND2_X1 U6959 ( .A1(n5445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U6960 ( .A(n5446), .B(P1_IR_REG_22__SCAN_IN), .ZN(n7393) );
  OR2_X1 U6961 ( .A1(n5254), .A2(n6340), .ZN(n5451) );
  NAND2_X1 U6962 ( .A1(n5447), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5449) );
  XNOR2_X1 U6963 ( .A(n5449), .B(n5448), .ZN(n6842) );
  INV_X1 U6964 ( .A(n6842), .ZN(n7957) );
  NAND2_X1 U6965 ( .A1(n7956), .A2(n7957), .ZN(n5450) );
  NAND2_X1 U6966 ( .A1(n7393), .A2(n7956), .ZN(n6589) );
  NOR2_X2 U6967 ( .A1(n7959), .A2(n6589), .ZN(n9154) );
  INV_X1 U6968 ( .A(n6589), .ZN(n7950) );
  NAND2_X1 U6969 ( .A1(n7959), .A2(n7950), .ZN(n9698) );
  INV_X1 U6970 ( .A(P1_B_REG_SCAN_IN), .ZN(n7963) );
  NOR2_X1 U6971 ( .A1(n9584), .A2(n7963), .ZN(n5452) );
  NOR2_X1 U6972 ( .A1(n9698), .A2(n5452), .ZN(n8961) );
  INV_X1 U6973 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n5456) );
  NAND2_X1 U6974 ( .A1(n4267), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n5455) );
  INV_X1 U6975 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n5453) );
  OR2_X1 U6976 ( .A1(n7680), .A2(n5453), .ZN(n5454) );
  OAI211_X1 U6977 ( .C1(n7683), .C2(n5456), .A(n5455), .B(n5454), .ZN(n8855)
         );
  NAND2_X1 U6978 ( .A1(n6339), .A2(n7950), .ZN(n6542) );
  NAND2_X1 U6979 ( .A1(n5460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5461) );
  NAND2_X1 U6980 ( .A1(n5462), .A2(n5461), .ZN(n5469) );
  NAND2_X1 U6981 ( .A1(n5464), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U6982 ( .A(n5465), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7580) );
  INV_X1 U6983 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6984 ( .A1(n5467), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5468) );
  XNOR2_X1 U6985 ( .A(n5468), .B(P1_IR_REG_25__SCAN_IN), .ZN(n7568) );
  NAND2_X1 U6986 ( .A1(n5469), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6987 ( .A1(n5471), .A2(n5470), .ZN(n7452) );
  AND2_X1 U6988 ( .A1(n7452), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5472) );
  NAND2_X1 U6989 ( .A1(n6590), .A2(n5472), .ZN(n7960) );
  INV_X1 U6990 ( .A(n7960), .ZN(n9402) );
  NAND2_X1 U6991 ( .A1(n6542), .A2(n9402), .ZN(n6785) );
  INV_X1 U6992 ( .A(n7568), .ZN(n5473) );
  NAND2_X1 U6993 ( .A1(n5473), .A2(P1_B_REG_SCAN_IN), .ZN(n5475) );
  MUX2_X1 U6994 ( .A(n5475), .B(P1_B_REG_SCAN_IN), .S(n5474), .Z(n5476) );
  NAND2_X1 U6995 ( .A1(n5476), .A2(n7580), .ZN(n9403) );
  INV_X1 U6996 ( .A(n9403), .ZN(n5478) );
  INV_X1 U6997 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5477) );
  NAND2_X1 U6998 ( .A1(n5478), .A2(n5477), .ZN(n5481) );
  INV_X1 U6999 ( .A(n5474), .ZN(n5480) );
  INV_X1 U7000 ( .A(n7580), .ZN(n5479) );
  NAND2_X1 U7001 ( .A1(n5480), .A2(n5479), .ZN(n9404) );
  NAND2_X1 U7002 ( .A1(n5481), .A2(n9404), .ZN(n6784) );
  INV_X1 U7003 ( .A(n6784), .ZN(n6781) );
  OAI22_X1 U7004 ( .A1(n9403), .A2(P1_D_REG_1__SCAN_IN), .B1(n7580), .B2(n7568), .ZN(n6777) );
  NOR4_X1 U7005 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5490) );
  NOR4_X1 U7006 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5489) );
  INV_X1 U7007 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n9715) );
  INV_X1 U7008 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9719) );
  INV_X1 U7009 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n9714) );
  INV_X1 U7010 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n9721) );
  NAND4_X1 U7011 ( .A1(n9715), .A2(n9719), .A3(n9714), .A4(n9721), .ZN(n5487)
         );
  NOR4_X1 U7012 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5485) );
  NOR4_X1 U7013 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n5484) );
  NOR4_X1 U7014 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5483) );
  NOR4_X1 U7015 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5482) );
  NAND4_X1 U7016 ( .A1(n5485), .A2(n5484), .A3(n5483), .A4(n5482), .ZN(n5486)
         );
  NOR4_X1 U7017 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5487), .A4(n5486), .ZN(n5488) );
  AND3_X1 U7018 ( .A1(n5490), .A2(n5489), .A3(n5488), .ZN(n5491) );
  NOR2_X1 U7019 ( .A1(n9403), .A2(n5491), .ZN(n6776) );
  OR2_X1 U7020 ( .A1(n6777), .A2(n6776), .ZN(n6534) );
  OR2_X1 U7021 ( .A1(n7960), .A2(n7956), .ZN(n5492) );
  NOR2_X1 U7022 ( .A1(n9182), .A2(n9708), .ZN(n5545) );
  NAND2_X1 U7023 ( .A1(n6335), .A2(n6851), .ZN(n6839) );
  NAND2_X1 U7024 ( .A1(n6346), .A2(n7080), .ZN(n6841) );
  NAND2_X1 U7025 ( .A1(n6839), .A2(n6841), .ZN(n5493) );
  NAND2_X1 U7026 ( .A1(n6775), .A2(n6930), .ZN(n6840) );
  NAND2_X1 U7027 ( .A1(n5493), .A2(n6840), .ZN(n7217) );
  NAND2_X1 U7028 ( .A1(n7764), .A2(n7217), .ZN(n5495) );
  NAND2_X1 U7029 ( .A1(n9697), .A2(n9724), .ZN(n5494) );
  NAND2_X1 U7030 ( .A1(n5495), .A2(n5494), .ZN(n9687) );
  NAND2_X1 U7031 ( .A1(n9687), .A2(n9694), .ZN(n5498) );
  NAND2_X1 U7032 ( .A1(n5496), .A2(n9730), .ZN(n5497) );
  NAND2_X1 U7033 ( .A1(n5498), .A2(n5497), .ZN(n7203) );
  NAND2_X1 U7034 ( .A1(n7729), .A2(n7800), .ZN(n7766) );
  INV_X1 U7035 ( .A(n7770), .ZN(n5499) );
  NAND2_X1 U7036 ( .A1(n9699), .A2(n9735), .ZN(n7191) );
  NAND2_X1 U7037 ( .A1(n8868), .A2(n6397), .ZN(n5500) );
  NAND2_X1 U7038 ( .A1(n9742), .A2(n5500), .ZN(n7321) );
  INV_X1 U7039 ( .A(n7321), .ZN(n5502) );
  NAND2_X1 U7040 ( .A1(n7185), .A2(n9748), .ZN(n5503) );
  NAND2_X1 U7041 ( .A1(n7830), .A2(n7833), .ZN(n7131) );
  INV_X1 U7042 ( .A(n7160), .ZN(n5505) );
  INV_X1 U7043 ( .A(n7737), .ZN(n7835) );
  NAND2_X1 U7044 ( .A1(n5505), .A2(n5504), .ZN(n7159) );
  NAND2_X1 U7045 ( .A1(n7313), .A2(n8865), .ZN(n5506) );
  AND2_X1 U7046 ( .A1(n7705), .A2(n8864), .ZN(n5507) );
  INV_X1 U7047 ( .A(n7848), .ZN(n5508) );
  NAND2_X1 U7048 ( .A1(n9505), .A2(n9552), .ZN(n5509) );
  NAND2_X1 U7049 ( .A1(n5510), .A2(n5509), .ZN(n7495) );
  INV_X1 U7050 ( .A(n7495), .ZN(n5512) );
  INV_X1 U7051 ( .A(n7712), .ZN(n7855) );
  INV_X1 U7052 ( .A(n7774), .ZN(n5511) );
  NAND2_X1 U7053 ( .A1(n7507), .A2(n8861), .ZN(n5513) );
  AND2_X1 U7054 ( .A1(n7673), .A2(n8859), .ZN(n5515) );
  OR2_X1 U7055 ( .A1(n7673), .A2(n8859), .ZN(n5514) );
  NAND2_X1 U7056 ( .A1(n8851), .A2(n8858), .ZN(n5516) );
  INV_X1 U7057 ( .A(n5517), .ZN(n7876) );
  NAND2_X1 U7058 ( .A1(n7877), .A2(n7876), .ZN(n7872) );
  NAND2_X1 U7059 ( .A1(n8762), .A2(n8857), .ZN(n5518) );
  NAND2_X1 U7060 ( .A1(n9236), .A2(n9138), .ZN(n5520) );
  NAND2_X1 U7061 ( .A1(n5521), .A2(n5520), .ZN(n9126) );
  NAND2_X1 U7062 ( .A1(n9126), .A2(n9127), .ZN(n5523) );
  NAND2_X1 U7063 ( .A1(n9232), .A2(n9153), .ZN(n5522) );
  NAND2_X1 U7064 ( .A1(n5523), .A2(n5522), .ZN(n9110) );
  AND2_X1 U7065 ( .A1(n9226), .A2(n9137), .ZN(n5525) );
  OR2_X1 U7066 ( .A1(n9226), .A2(n9137), .ZN(n5524) );
  INV_X1 U7067 ( .A(n9097), .ZN(n7781) );
  NAND2_X1 U7068 ( .A1(n7906), .A2(n7907), .ZN(n9087) );
  NAND2_X1 U7069 ( .A1(n9216), .A2(n9071), .ZN(n5526) );
  NAND2_X1 U7070 ( .A1(n9078), .A2(n5526), .ZN(n9061) );
  INV_X1 U7071 ( .A(n9069), .ZN(n9060) );
  NAND2_X1 U7072 ( .A1(n9061), .A2(n9060), .ZN(n9059) );
  NAND2_X1 U7073 ( .A1(n9211), .A2(n9088), .ZN(n5527) );
  NAND2_X1 U7074 ( .A1(n9059), .A2(n5527), .ZN(n9043) );
  NAND2_X1 U7075 ( .A1(n9206), .A2(n9072), .ZN(n5528) );
  NAND2_X1 U7076 ( .A1(n9196), .A2(n8856), .ZN(n7784) );
  NAND2_X1 U7077 ( .A1(n5530), .A2(n7784), .ZN(n8992) );
  INV_X1 U7078 ( .A(n8999), .ZN(n7922) );
  INV_X1 U7079 ( .A(n8982), .ZN(n9184) );
  NAND2_X1 U7080 ( .A1(n8982), .A2(n5531), .ZN(n5532) );
  XNOR2_X2 U7081 ( .A(n5533), .B(n7759), .ZN(n9183) );
  INV_X1 U7082 ( .A(n5536), .ZN(n5535) );
  NAND2_X1 U7083 ( .A1(n7956), .A2(n6842), .ZN(n6927) );
  INV_X1 U7084 ( .A(n6927), .ZN(n6334) );
  AND2_X1 U7085 ( .A1(n5535), .A2(n6334), .ZN(n6838) );
  NOR2_X1 U7086 ( .A1(n6838), .A2(n6362), .ZN(n5537) );
  NAND2_X1 U7087 ( .A1(n9684), .A2(n5537), .ZN(n9176) );
  INV_X1 U7088 ( .A(n9191), .ZN(n8998) );
  NAND2_X1 U7089 ( .A1(n7323), .A2(n9748), .ZN(n7325) );
  OR2_X2 U7090 ( .A1(n7325), .A2(n7130), .ZN(n7154) );
  INV_X1 U7091 ( .A(n7705), .ZN(n9760) );
  INV_X1 U7092 ( .A(n7416), .ZN(n7435) );
  NAND2_X1 U7093 ( .A1(n9671), .A2(n7435), .ZN(n7302) );
  OR2_X2 U7094 ( .A1(n7302), .A2(n7459), .ZN(n9506) );
  OR2_X2 U7095 ( .A1(n9506), .A2(n7507), .ZN(n9487) );
  NOR2_X2 U7096 ( .A1(n9487), .A2(n9486), .ZN(n9488) );
  INV_X1 U7097 ( .A(n7673), .ZN(n9536) );
  INV_X1 U7098 ( .A(n8851), .ZN(n9248) );
  INV_X1 U7099 ( .A(n8762), .ZN(n9531) );
  NOR2_X1 U7100 ( .A1(n9167), .A2(n9236), .ZN(n9144) );
  INV_X1 U7101 ( .A(n9232), .ZN(n9133) );
  INV_X1 U7102 ( .A(n9226), .ZN(n9118) );
  NAND2_X1 U7103 ( .A1(n9128), .A2(n9118), .ZN(n9113) );
  OR2_X2 U7104 ( .A1(n9113), .A2(n9223), .ZN(n9101) );
  INV_X1 U7105 ( .A(n9211), .ZN(n9067) );
  INV_X1 U7106 ( .A(n9206), .ZN(n9049) );
  NAND2_X1 U7107 ( .A1(n8998), .A2(n9010), .ZN(n8993) );
  AOI21_X1 U7108 ( .B1(n9180), .B2(n8984), .A(n8966), .ZN(n9181) );
  INV_X1 U7109 ( .A(n7956), .ZN(n7794) );
  AND2_X1 U7110 ( .A1(n6340), .A2(n7794), .ZN(n6843) );
  INV_X1 U7111 ( .A(n6843), .ZN(n6772) );
  NOR2_X1 U7112 ( .A1(n6339), .A2(n6772), .ZN(n5538) );
  INV_X1 U7113 ( .A(n9180), .ZN(n7939) );
  AND2_X1 U7114 ( .A1(n6843), .A2(n7957), .ZN(n6546) );
  INV_X1 U7115 ( .A(n5539), .ZN(n5540) );
  AOI22_X1 U7116 ( .A1(n5540), .A2(n9707), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9708), .ZN(n5541) );
  OAI21_X1 U7117 ( .B1(n7939), .B2(n9710), .A(n5541), .ZN(n5542) );
  NOR2_X1 U7118 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5549) );
  NOR2_X1 U7119 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5555) );
  NOR2_X1 U7120 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5554) );
  NOR2_X1 U7121 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5553) );
  NAND4_X1 U7122 ( .A1(n5555), .A2(n5554), .A3(n5553), .A4(n6051), .ZN(n5556)
         );
  INV_X1 U7123 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5558) );
  INV_X1 U7124 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U7125 ( .A1(n5581), .A2(n5559), .ZN(n5562) );
  NAND2_X1 U7126 ( .A1(n5623), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7127 ( .A1(n5610), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5566) );
  INV_X1 U7128 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5570) );
  INV_X1 U7129 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5571) );
  INV_X1 U7130 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U7131 ( .A1(n5576), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5577) );
  XNOR2_X1 U7132 ( .A(n5577), .B(n5573), .ZN(n7309) );
  INV_X1 U7133 ( .A(n7309), .ZN(n6806) );
  NAND2_X1 U7134 ( .A1(n5889), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5578) );
  MUX2_X1 U7135 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5578), .S(
        P2_IR_REG_19__SCAN_IN), .Z(n5579) );
  NAND2_X1 U7136 ( .A1(n5579), .A2(n5576), .ZN(n8443) );
  INV_X1 U7137 ( .A(n6811), .ZN(n6289) );
  NAND2_X1 U7138 ( .A1(n6319), .A2(n7309), .ZN(n7040) );
  OR3_X1 U7139 ( .A1(n5586), .A2(n5558), .A3(n6055), .ZN(n5584) );
  NAND2_X4 U7140 ( .A1(n6092), .A2(n8004), .ZN(n6710) );
  NAND2_X2 U7141 ( .A1(n6710), .A2(n5587), .ZN(n5628) );
  NAND2_X1 U7142 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5588) );
  MUX2_X1 U7143 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5588), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5591) );
  INV_X1 U7144 ( .A(n5589), .ZN(n5590) );
  NAND2_X1 U7145 ( .A1(n5591), .A2(n5590), .ZN(n6727) );
  NAND2_X2 U7146 ( .A1(n6710), .A2(n6567), .ZN(n5629) );
  INV_X1 U7147 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6569) );
  NAND2_X2 U7148 ( .A1(n5593), .A2(n5594), .ZN(n6114) );
  XNOR2_X1 U7149 ( .A(n5651), .B(n6114), .ZN(n5606) );
  XNOR2_X1 U7150 ( .A(n5608), .B(n5606), .ZN(n6766) );
  NAND2_X1 U7151 ( .A1(n5621), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7152 ( .A1(n5640), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7153 ( .A1(n5623), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5595) );
  INV_X1 U7154 ( .A(SI_0_), .ZN(n5600) );
  INV_X1 U7155 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5599) );
  OAI21_X1 U7156 ( .B1(n6567), .B2(n5600), .A(n5599), .ZN(n5602) );
  AND2_X1 U7157 ( .A1(n5602), .A2(n5601), .ZN(n8724) );
  MUX2_X1 U7158 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8724), .S(n6710), .Z(n9865) );
  INV_X1 U7159 ( .A(n9835), .ZN(n5604) );
  NAND2_X1 U7160 ( .A1(n5604), .A2(n6171), .ZN(n6827) );
  INV_X1 U7161 ( .A(n9865), .ZN(n6833) );
  NAND2_X1 U7162 ( .A1(n6833), .A2(n6045), .ZN(n5605) );
  INV_X1 U7163 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U7164 ( .A1(n5608), .A2(n5607), .ZN(n5609) );
  NAND2_X1 U7165 ( .A1(n5640), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7166 ( .A1(n5610), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7167 ( .A1(n5621), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5612) );
  NAND2_X1 U7168 ( .A1(n5623), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5611) );
  AND4_X2 U7169 ( .A1(n5614), .A2(n5613), .A3(n5612), .A4(n5611), .ZN(n8060)
         );
  NOR2_X1 U7170 ( .A1(n8060), .A2(n6828), .ZN(n5616) );
  INV_X1 U7171 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6055) );
  OR2_X1 U7172 ( .A1(n5589), .A2(n6055), .ZN(n5615) );
  XNOR2_X1 U7173 ( .A(n5615), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9453) );
  INV_X1 U7174 ( .A(n9453), .ZN(n6574) );
  XNOR2_X1 U7175 ( .A(n6807), .B(n5651), .ZN(n5617) );
  NAND2_X1 U7176 ( .A1(n5616), .A2(n5617), .ZN(n5620) );
  INV_X1 U7177 ( .A(n5616), .ZN(n5618) );
  INV_X1 U7178 ( .A(n5617), .ZN(n8061) );
  NAND2_X1 U7179 ( .A1(n5618), .A2(n8061), .ZN(n5619) );
  AND2_X1 U7180 ( .A1(n5620), .A2(n5619), .ZN(n6792) );
  NAND2_X1 U7181 ( .A1(n5621), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5627) );
  INV_X1 U7182 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U7183 ( .A1(n5640), .A2(n8070), .ZN(n5626) );
  INV_X2 U7184 ( .A(n5622), .ZN(n6150) );
  NAND2_X1 U7185 ( .A1(n6150), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7186 ( .A1(n5623), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5624) );
  AND2_X1 U7187 ( .A1(n8236), .A2(n6171), .ZN(n5636) );
  OR2_X1 U7188 ( .A1(n5628), .A2(n6570), .ZN(n5634) );
  OR2_X1 U7189 ( .A1(n5629), .A2(n6571), .ZN(n5633) );
  INV_X2 U7190 ( .A(n6710), .ZN(n5906) );
  NAND2_X1 U7191 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5630), .ZN(n5631) );
  XNOR2_X1 U7192 ( .A(n5631), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U7193 ( .A1(n5906), .A2(n6723), .ZN(n5632) );
  XNOR2_X1 U7194 ( .A(n9818), .B(n6045), .ZN(n5635) );
  NAND2_X1 U7195 ( .A1(n5636), .A2(n5635), .ZN(n5652) );
  INV_X1 U7196 ( .A(n5635), .ZN(n8164) );
  INV_X1 U7197 ( .A(n5636), .ZN(n5637) );
  NAND2_X1 U7198 ( .A1(n8164), .A2(n5637), .ZN(n5638) );
  AND2_X1 U7199 ( .A1(n5652), .A2(n5638), .ZN(n8062) );
  NAND2_X1 U7200 ( .A1(n5639), .A2(n8062), .ZN(n8065) );
  INV_X1 U7201 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7202 ( .A1(n5641), .A2(n8070), .ZN(n5642) );
  AND2_X1 U7203 ( .A1(n5642), .A2(n5659), .ZN(n8160) );
  NAND2_X1 U7204 ( .A1(n5640), .A2(n8160), .ZN(n5646) );
  NAND2_X1 U7205 ( .A1(n6150), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U7206 ( .A1(n5623), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7207 ( .A1(n6152), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5643) );
  OR2_X1 U7208 ( .A1(n7020), .A2(n6828), .ZN(n5656) );
  OR2_X1 U7209 ( .A1(n5647), .A2(n6055), .ZN(n5648) );
  XNOR2_X1 U7210 ( .A(n5648), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6889) );
  INV_X1 U7211 ( .A(n6889), .ZN(n6911) );
  OR2_X1 U7212 ( .A1(n5628), .A2(n6572), .ZN(n5650) );
  OR2_X1 U7213 ( .A1(n5629), .A2(n6573), .ZN(n5649) );
  OAI211_X1 U7214 ( .C1(n6710), .C2(n6911), .A(n5650), .B(n5649), .ZN(n7098)
         );
  XNOR2_X1 U7215 ( .A(n7098), .B(n6024), .ZN(n5654) );
  XNOR2_X1 U7216 ( .A(n5656), .B(n5654), .ZN(n8163) );
  AND2_X1 U7217 ( .A1(n8163), .A2(n5652), .ZN(n5653) );
  NAND2_X1 U7218 ( .A1(n8065), .A2(n5653), .ZN(n8161) );
  INV_X1 U7219 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U7220 ( .A1(n5656), .A2(n5655), .ZN(n5657) );
  INV_X1 U7221 ( .A(n5659), .ZN(n5658) );
  INV_X1 U7222 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8242) );
  NAND2_X1 U7223 ( .A1(n5659), .A2(n8242), .ZN(n5660) );
  AND2_X1 U7224 ( .A1(n5701), .A2(n5660), .ZN(n7058) );
  NAND2_X1 U7225 ( .A1(n5640), .A2(n7058), .ZN(n5664) );
  NAND2_X1 U7226 ( .A1(n5623), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7227 ( .A1(n6152), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5661) );
  NOR2_X1 U7228 ( .A1(n8157), .A2(n6828), .ZN(n5669) );
  INV_X1 U7229 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5665) );
  NAND2_X1 U7230 ( .A1(n5647), .A2(n5665), .ZN(n5666) );
  NAND2_X1 U7231 ( .A1(n5666), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5680) );
  XNOR2_X1 U7232 ( .A(n5680), .B(P2_IR_REG_5__SCAN_IN), .ZN(n8244) );
  INV_X1 U7233 ( .A(n8244), .ZN(n6577) );
  OR2_X1 U7234 ( .A1(n5628), .A2(n6578), .ZN(n5668) );
  OR2_X1 U7235 ( .A1(n5629), .A2(n6579), .ZN(n5667) );
  OAI211_X1 U7236 ( .C1(n6710), .C2(n6577), .A(n5668), .B(n5667), .ZN(n7031)
         );
  XNOR2_X1 U7237 ( .A(n7031), .B(n6024), .ZN(n6944) );
  NAND2_X1 U7238 ( .A1(n5669), .A2(n6944), .ZN(n5687) );
  INV_X1 U7239 ( .A(n5669), .ZN(n5671) );
  INV_X1 U7240 ( .A(n6944), .ZN(n5670) );
  NAND2_X1 U7241 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  NAND2_X1 U7242 ( .A1(n5687), .A2(n5672), .ZN(n6956) );
  XNOR2_X1 U7243 ( .A(n5701), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n6947) );
  NAND2_X1 U7244 ( .A1(n5640), .A2(n6947), .ZN(n5678) );
  NAND2_X1 U7245 ( .A1(n6150), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7246 ( .A1(n5623), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U7247 ( .A1(n6152), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5675) );
  OR2_X1 U7248 ( .A1(n7118), .A2(n6828), .ZN(n5691) );
  INV_X2 U7249 ( .A(n5628), .ZN(n5713) );
  NAND2_X1 U7250 ( .A1(n6583), .A2(n5713), .ZN(n5686) );
  INV_X1 U7251 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7252 ( .A1(n5680), .A2(n5679), .ZN(n5681) );
  NAND2_X1 U7253 ( .A1(n5681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5683) );
  INV_X1 U7254 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5682) );
  NAND2_X1 U7255 ( .A1(n5683), .A2(n5682), .ZN(n5693) );
  OR2_X1 U7256 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  AOI22_X1 U7257 ( .A1(n5887), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5906), .B2(
        n8258), .ZN(n5685) );
  XNOR2_X1 U7258 ( .A(n7109), .B(n6045), .ZN(n5689) );
  XNOR2_X1 U7259 ( .A(n5691), .B(n5689), .ZN(n6943) );
  AND2_X1 U7260 ( .A1(n6943), .A2(n5687), .ZN(n5688) );
  INV_X1 U7261 ( .A(n5689), .ZN(n5690) );
  NAND2_X1 U7262 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  NAND2_X1 U7263 ( .A1(n4361), .A2(n5713), .ZN(n5696) );
  NAND2_X1 U7264 ( .A1(n5693), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5694) );
  XNOR2_X1 U7265 ( .A(n5694), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8271) );
  AOI22_X1 U7266 ( .A1(n5887), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5906), .B2(
        n8271), .ZN(n5695) );
  XNOR2_X1 U7267 ( .A(n8039), .B(n6024), .ZN(n5707) );
  INV_X1 U7268 ( .A(n5701), .ZN(n5698) );
  NAND2_X1 U7269 ( .A1(n5698), .A2(n5697), .ZN(n5721) );
  INV_X1 U7270 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5700) );
  INV_X1 U7271 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5699) );
  OAI21_X1 U7272 ( .B1(n5701), .B2(n5700), .A(n5699), .ZN(n5702) );
  AND2_X1 U7273 ( .A1(n5721), .A2(n5702), .ZN(n8038) );
  NAND2_X1 U7274 ( .A1(n5640), .A2(n8038), .ZN(n5706) );
  NAND2_X1 U7275 ( .A1(n6150), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U7276 ( .A1(n5623), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7277 ( .A1(n6152), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5703) );
  NOR2_X1 U7278 ( .A1(n8088), .A2(n6828), .ZN(n5708) );
  NAND2_X1 U7279 ( .A1(n5707), .A2(n5708), .ZN(n5712) );
  INV_X1 U7280 ( .A(n5707), .ZN(n8089) );
  INV_X1 U7281 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U7282 ( .A1(n8089), .A2(n5709), .ZN(n5710) );
  NAND2_X1 U7283 ( .A1(n5712), .A2(n5710), .ZN(n8034) );
  NAND2_X1 U7284 ( .A1(n6608), .A2(n5713), .ZN(n5719) );
  NOR2_X1 U7285 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5714) );
  AND2_X1 U7286 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  NAND2_X1 U7287 ( .A1(n5647), .A2(n5716), .ZN(n5732) );
  NAND2_X1 U7288 ( .A1(n5732), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5717) );
  XNOR2_X1 U7289 ( .A(n5717), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8284) );
  AOI22_X1 U7290 ( .A1(n5887), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5906), .B2(
        n8284), .ZN(n5718) );
  NAND2_X1 U7291 ( .A1(n5719), .A2(n5718), .ZN(n8094) );
  XNOR2_X1 U7292 ( .A(n8094), .B(n6045), .ZN(n5728) );
  INV_X1 U7293 ( .A(n5721), .ZN(n5720) );
  NAND2_X1 U7294 ( .A1(n5720), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5736) );
  INV_X1 U7295 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9342) );
  NAND2_X1 U7296 ( .A1(n5721), .A2(n9342), .ZN(n5722) );
  AND2_X1 U7297 ( .A1(n5736), .A2(n5722), .ZN(n8093) );
  NAND2_X1 U7298 ( .A1(n5640), .A2(n8093), .ZN(n5726) );
  NAND2_X1 U7299 ( .A1(n6151), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U7300 ( .A1(n6152), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5723) );
  NOR2_X1 U7301 ( .A1(n7262), .A2(n6828), .ZN(n5729) );
  XNOR2_X1 U7302 ( .A(n5728), .B(n5729), .ZN(n8085) );
  NAND2_X1 U7303 ( .A1(n5727), .A2(n8085), .ZN(n8090) );
  INV_X1 U7304 ( .A(n5728), .ZN(n5730) );
  NAND2_X1 U7305 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  NAND2_X1 U7306 ( .A1(n8090), .A2(n5731), .ZN(n7234) );
  NAND2_X1 U7307 ( .A1(n6616), .A2(n5713), .ZN(n5734) );
  NAND2_X1 U7308 ( .A1(n5785), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5746) );
  XNOR2_X1 U7309 ( .A(n5746), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8297) );
  AOI22_X1 U7310 ( .A1(n5887), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5906), .B2(
        n8297), .ZN(n5733) );
  XNOR2_X1 U7311 ( .A(n7354), .B(n6045), .ZN(n5743) );
  INV_X1 U7312 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7313 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  AND2_X1 U7314 ( .A1(n5754), .A2(n5737), .ZN(n7269) );
  NAND2_X1 U7315 ( .A1(n5640), .A2(n7269), .ZN(n5741) );
  NAND2_X1 U7316 ( .A1(n6150), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U7317 ( .A1(n6151), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7318 ( .A1(n6152), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5738) );
  OR2_X1 U7319 ( .A1(n7359), .A2(n6828), .ZN(n5744) );
  NAND2_X1 U7320 ( .A1(n5743), .A2(n5744), .ZN(n5742) );
  INV_X1 U7321 ( .A(n5743), .ZN(n7236) );
  INV_X1 U7322 ( .A(n5744), .ZN(n5745) );
  NAND2_X1 U7323 ( .A1(n7236), .A2(n5745), .ZN(n7232) );
  NAND2_X1 U7324 ( .A1(n6664), .A2(n5713), .ZN(n5751) );
  INV_X1 U7325 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5783) );
  NAND2_X1 U7326 ( .A1(n5746), .A2(n5783), .ZN(n5747) );
  NAND2_X1 U7327 ( .A1(n5747), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7328 ( .A1(n5748), .A2(n5782), .ZN(n5765) );
  OR2_X1 U7329 ( .A1(n5748), .A2(n5782), .ZN(n5749) );
  AND2_X1 U7330 ( .A1(n5765), .A2(n5749), .ZN(n6974) );
  AOI22_X1 U7331 ( .A1(n5887), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5906), .B2(
        n6974), .ZN(n5750) );
  NAND2_X1 U7332 ( .A1(n5751), .A2(n5750), .ZN(n7397) );
  XNOR2_X1 U7333 ( .A(n7397), .B(n6024), .ZN(n5760) );
  INV_X1 U7334 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7335 ( .A1(n5754), .A2(n5753), .ZN(n5755) );
  AND2_X1 U7336 ( .A1(n5770), .A2(n5755), .ZN(n7367) );
  NAND2_X1 U7337 ( .A1(n5640), .A2(n7367), .ZN(n5759) );
  NAND2_X1 U7338 ( .A1(n6151), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U7339 ( .A1(n5621), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5756) );
  NOR2_X1 U7340 ( .A1(n7404), .A2(n6828), .ZN(n5761) );
  NAND2_X1 U7341 ( .A1(n5760), .A2(n5761), .ZN(n5764) );
  INV_X1 U7342 ( .A(n5760), .ZN(n7340) );
  INV_X1 U7343 ( .A(n5761), .ZN(n5762) );
  NAND2_X1 U7344 ( .A1(n7340), .A2(n5762), .ZN(n5763) );
  AND2_X1 U7345 ( .A1(n5764), .A2(n5763), .ZN(n7245) );
  NAND2_X1 U7346 ( .A1(n6666), .A2(n5713), .ZN(n5768) );
  NAND2_X1 U7347 ( .A1(n5765), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5766) );
  XNOR2_X1 U7348 ( .A(n5766), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7141) );
  AOI22_X1 U7349 ( .A1(n5887), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5906), .B2(
        n7141), .ZN(n5767) );
  NAND2_X1 U7350 ( .A1(n5768), .A2(n5767), .ZN(n7589) );
  XNOR2_X1 U7351 ( .A(n7589), .B(n6024), .ZN(n5776) );
  INV_X1 U7352 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U7353 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  AND2_X1 U7354 ( .A1(n5790), .A2(n5771), .ZN(n7406) );
  NAND2_X1 U7355 ( .A1(n5640), .A2(n7406), .ZN(n5775) );
  NAND2_X1 U7356 ( .A1(n6151), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U7357 ( .A1(n5621), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5772) );
  NOR2_X1 U7358 ( .A1(n7588), .A2(n6828), .ZN(n5777) );
  NAND2_X1 U7359 ( .A1(n5776), .A2(n5777), .ZN(n5796) );
  INV_X1 U7360 ( .A(n5776), .ZN(n7436) );
  INV_X1 U7361 ( .A(n5777), .ZN(n5778) );
  NAND2_X1 U7362 ( .A1(n7436), .A2(n5778), .ZN(n5779) );
  AND2_X1 U7363 ( .A1(n5796), .A2(n5779), .ZN(n7337) );
  NAND2_X1 U7364 ( .A1(n5780), .A2(n7337), .ZN(n7341) );
  NAND2_X1 U7365 ( .A1(n6680), .A2(n5713), .ZN(n5788) );
  NAND3_X1 U7366 ( .A1(n5783), .A2(n5782), .A3(n5781), .ZN(n5784) );
  NOR2_X1 U7367 ( .A1(n5785), .A2(n5784), .ZN(n5803) );
  OR2_X1 U7368 ( .A1(n5803), .A2(n6055), .ZN(n5786) );
  XNOR2_X1 U7369 ( .A(n5786), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7279) );
  AOI22_X1 U7370 ( .A1(n5887), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5906), .B2(
        n7279), .ZN(n5787) );
  XNOR2_X1 U7371 ( .A(n9928), .B(n6045), .ZN(n5800) );
  INV_X1 U7372 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7145) );
  NAND2_X1 U7373 ( .A1(n5790), .A2(n7145), .ZN(n5791) );
  AND2_X1 U7374 ( .A1(n5806), .A2(n5791), .ZN(n9803) );
  NAND2_X1 U7375 ( .A1(n5640), .A2(n9803), .ZN(n5795) );
  NAND2_X1 U7376 ( .A1(n6150), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5794) );
  NAND2_X1 U7377 ( .A1(n6151), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7378 ( .A1(n6152), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5792) );
  NOR2_X1 U7379 ( .A1(n7600), .A2(n6828), .ZN(n5798) );
  XNOR2_X1 U7380 ( .A(n5800), .B(n5798), .ZN(n7447) );
  AND2_X1 U7381 ( .A1(n7447), .A2(n5796), .ZN(n5797) );
  NAND2_X1 U7382 ( .A1(n7341), .A2(n5797), .ZN(n7443) );
  INV_X1 U7383 ( .A(n5798), .ZN(n5799) );
  NAND2_X1 U7384 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  NAND2_X1 U7385 ( .A1(n6684), .A2(n5713), .ZN(n5805) );
  INV_X1 U7386 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7387 ( .A1(n5803), .A2(n5802), .ZN(n5854) );
  NAND2_X1 U7388 ( .A1(n5854), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  XNOR2_X1 U7389 ( .A(n5816), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7383) );
  AOI22_X1 U7390 ( .A1(n5887), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5906), .B2(
        n7383), .ZN(n5804) );
  XNOR2_X1 U7391 ( .A(n7614), .B(n6024), .ZN(n5812) );
  INV_X1 U7392 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7282) );
  NAND2_X1 U7393 ( .A1(n5806), .A2(n7282), .ZN(n5807) );
  AND2_X1 U7394 ( .A1(n5823), .A2(n5807), .ZN(n7608) );
  NAND2_X1 U7395 ( .A1(n5640), .A2(n7608), .ZN(n5811) );
  NAND2_X1 U7396 ( .A1(n6150), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U7397 ( .A1(n6151), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5809) );
  NAND2_X1 U7398 ( .A1(n5621), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5808) );
  NOR2_X1 U7399 ( .A1(n7619), .A2(n6828), .ZN(n5813) );
  NAND2_X1 U7400 ( .A1(n5812), .A2(n5813), .ZN(n5829) );
  INV_X1 U7401 ( .A(n5812), .ZN(n7555) );
  INV_X1 U7402 ( .A(n5813), .ZN(n5814) );
  NAND2_X1 U7403 ( .A1(n7555), .A2(n5814), .ZN(n5815) );
  NAND2_X1 U7404 ( .A1(n5829), .A2(n5815), .ZN(n6555) );
  NAND2_X1 U7405 ( .A1(n6756), .A2(n5713), .ZN(n5821) );
  INV_X1 U7406 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5852) );
  NAND2_X1 U7407 ( .A1(n5816), .A2(n5852), .ZN(n5817) );
  NAND2_X1 U7408 ( .A1(n5817), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5818) );
  INV_X1 U7409 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U7410 ( .A1(n5818), .A2(n5851), .ZN(n5835) );
  OR2_X1 U7411 ( .A1(n5818), .A2(n5851), .ZN(n5819) );
  AND2_X1 U7412 ( .A1(n5835), .A2(n5819), .ZN(n8312) );
  AOI22_X1 U7413 ( .A1(n5887), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5906), .B2(
        n8312), .ZN(n5820) );
  XNOR2_X1 U7414 ( .A(n7620), .B(n6024), .ZN(n5831) );
  NAND2_X1 U7415 ( .A1(n6152), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5828) );
  INV_X1 U7416 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5822) );
  NAND2_X1 U7417 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  AND2_X1 U7418 ( .A1(n5840), .A2(n5824), .ZN(n7622) );
  NAND2_X1 U7419 ( .A1(n5640), .A2(n7622), .ZN(n5827) );
  NAND2_X1 U7420 ( .A1(n6151), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5825) );
  NAND4_X1 U7421 ( .A1(n5828), .A2(n5827), .A3(n5826), .A4(n5825), .ZN(n8225)
         );
  NAND2_X1 U7422 ( .A1(n8225), .A2(n6171), .ZN(n5832) );
  XNOR2_X1 U7423 ( .A(n5831), .B(n5832), .ZN(n7565) );
  AND2_X1 U7424 ( .A1(n7565), .A2(n5829), .ZN(n5830) );
  INV_X1 U7425 ( .A(n5831), .ZN(n5833) );
  NAND2_X1 U7426 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  NAND2_X1 U7427 ( .A1(n5835), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U7428 ( .A(n5836), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8326) );
  AOI22_X1 U7429 ( .A1(n5887), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5906), .B2(
        n8326), .ZN(n5837) );
  XNOR2_X1 U7430 ( .A(n7976), .B(n6045), .ZN(n5847) );
  INV_X1 U7431 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7432 ( .A1(n5840), .A2(n5839), .ZN(n5841) );
  AND2_X1 U7433 ( .A1(n5860), .A2(n5841), .ZN(n8612) );
  NAND2_X1 U7434 ( .A1(n5640), .A2(n8612), .ZN(n5845) );
  NAND2_X1 U7435 ( .A1(n6151), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7436 ( .A1(n5621), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5842) );
  NOR2_X1 U7437 ( .A1(n8126), .A2(n6828), .ZN(n5846) );
  NAND2_X1 U7438 ( .A1(n6925), .A2(n5713), .ZN(n5858) );
  INV_X1 U7439 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5850) );
  NAND3_X1 U7440 ( .A1(n5852), .A2(n5851), .A3(n5850), .ZN(n5853) );
  OAI21_X1 U7441 ( .B1(n5854), .B2(n5853), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5855) );
  MUX2_X1 U7442 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5855), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n5856) );
  AND2_X1 U7443 ( .A1(n5849), .A2(n5856), .ZN(n8335) );
  AOI22_X1 U7444 ( .A1(n5887), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5906), .B2(
        n8335), .ZN(n5857) );
  XNOR2_X1 U7445 ( .A(n8692), .B(n6024), .ZN(n5867) );
  INV_X1 U7446 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U7447 ( .A1(n5860), .A2(n8322), .ZN(n5861) );
  AND2_X1 U7448 ( .A1(n5876), .A2(n5861), .ZN(n8594) );
  NAND2_X1 U7449 ( .A1(n5640), .A2(n8594), .ZN(n5865) );
  NAND2_X1 U7450 ( .A1(n6150), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7451 ( .A1(n6151), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7452 ( .A1(n5621), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5862) );
  NOR2_X1 U7453 ( .A1(n8137), .A2(n6828), .ZN(n5868) );
  XNOR2_X1 U7454 ( .A(n5867), .B(n5868), .ZN(n8125) );
  INV_X1 U7455 ( .A(n5867), .ZN(n5870) );
  INV_X1 U7456 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U7457 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7458 ( .A1(n6962), .A2(n5713), .ZN(n5875) );
  NAND2_X1 U7459 ( .A1(n5849), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5872) );
  MUX2_X1 U7460 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5872), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n5873) );
  AND2_X1 U7461 ( .A1(n5873), .A2(n5569), .ZN(n8357) );
  AOI22_X1 U7462 ( .A1(n5887), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5906), .B2(
        n8357), .ZN(n5874) );
  XNOR2_X1 U7463 ( .A(n8687), .B(n6024), .ZN(n5882) );
  NAND2_X1 U7464 ( .A1(n6151), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5881) );
  INV_X1 U7465 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U7466 ( .A1(n5876), .A2(n8139), .ZN(n5877) );
  AND2_X1 U7467 ( .A1(n5896), .A2(n5877), .ZN(n8582) );
  NAND2_X1 U7468 ( .A1(n5640), .A2(n8582), .ZN(n5880) );
  NAND2_X1 U7469 ( .A1(n6150), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5879) );
  NAND2_X1 U7470 ( .A1(n5621), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5878) );
  NAND4_X1 U7471 ( .A1(n5881), .A2(n5880), .A3(n5879), .A4(n5878), .ZN(n8570)
         );
  AND2_X1 U7472 ( .A1(n8570), .A2(n6171), .ZN(n5883) );
  NAND2_X1 U7473 ( .A1(n5882), .A2(n5883), .ZN(n5886) );
  INV_X1 U7474 ( .A(n5882), .ZN(n8195) );
  INV_X1 U7475 ( .A(n5883), .ZN(n5884) );
  NAND2_X1 U7476 ( .A1(n8195), .A2(n5884), .ZN(n5885) );
  AND2_X1 U7477 ( .A1(n5886), .A2(n5885), .ZN(n8136) );
  NAND2_X1 U7478 ( .A1(n8135), .A2(n5886), .ZN(n5905) );
  NAND2_X1 U7479 ( .A1(n7084), .A2(n5713), .ZN(n5892) );
  NAND2_X1 U7480 ( .A1(n5569), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5888) );
  MUX2_X1 U7481 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5888), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n5890) );
  NAND2_X1 U7482 ( .A1(n5890), .A2(n5889), .ZN(n8360) );
  INV_X1 U7483 ( .A(n8360), .ZN(n8371) );
  AOI22_X1 U7484 ( .A1(n5887), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5906), .B2(
        n8371), .ZN(n5891) );
  XNOR2_X1 U7485 ( .A(n8681), .B(n6024), .ZN(n5901) );
  NAND2_X1 U7486 ( .A1(n6151), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n5894) );
  NAND2_X1 U7487 ( .A1(n6152), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5893) );
  AND2_X1 U7488 ( .A1(n5894), .A2(n5893), .ZN(n5900) );
  INV_X1 U7489 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8355) );
  NAND2_X1 U7490 ( .A1(n5896), .A2(n8355), .ZN(n5897) );
  NAND2_X1 U7491 ( .A1(n5910), .A2(n5897), .ZN(n8564) );
  OR2_X1 U7492 ( .A1(n8564), .A2(n6038), .ZN(n5899) );
  NOR2_X1 U7493 ( .A1(n8138), .A2(n6828), .ZN(n5902) );
  NAND2_X1 U7494 ( .A1(n5901), .A2(n5902), .ZN(n5914) );
  INV_X1 U7495 ( .A(n5901), .ZN(n8075) );
  INV_X1 U7496 ( .A(n5902), .ZN(n5903) );
  NAND2_X1 U7497 ( .A1(n8075), .A2(n5903), .ZN(n5904) );
  AND2_X1 U7498 ( .A1(n5914), .A2(n5904), .ZN(n8191) );
  NAND2_X1 U7499 ( .A1(n5905), .A2(n8191), .ZN(n8074) );
  NAND2_X1 U7500 ( .A1(n7107), .A2(n5713), .ZN(n5908) );
  AOI22_X1 U7501 ( .A1(n5887), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8377), .B2(
        n5906), .ZN(n5907) );
  XNOR2_X1 U7502 ( .A(n8677), .B(n6024), .ZN(n5916) );
  INV_X1 U7503 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7504 ( .A1(n5910), .A2(n5909), .ZN(n5911) );
  NAND2_X1 U7505 ( .A1(n5924), .A2(n5911), .ZN(n8550) );
  AOI22_X1 U7506 ( .A1(n6151), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n6152), .B2(
        P2_REG0_REG_19__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U7507 ( .A1(n6150), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5912) );
  OAI211_X1 U7508 ( .C1(n8550), .C2(n6038), .A(n5913), .B(n5912), .ZN(n8573)
         );
  NAND2_X1 U7509 ( .A1(n8573), .A2(n6171), .ZN(n5917) );
  XNOR2_X1 U7510 ( .A(n5916), .B(n5917), .ZN(n8083) );
  AND2_X1 U7511 ( .A1(n8083), .A2(n5914), .ZN(n5915) );
  INV_X1 U7512 ( .A(n5916), .ZN(n5918) );
  NAND2_X1 U7513 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  NAND2_X1 U7514 ( .A1(n7229), .A2(n5713), .ZN(n5921) );
  NAND2_X1 U7515 ( .A1(n5887), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5920) );
  XNOR2_X1 U7516 ( .A(n8671), .B(n6024), .ZN(n5929) );
  INV_X1 U7517 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7518 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  NAND2_X1 U7519 ( .A1(n5937), .A2(n5925), .ZN(n8173) );
  OR2_X1 U7520 ( .A1(n8173), .A2(n6038), .ZN(n5928) );
  AOI22_X1 U7521 ( .A1(n6151), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n6152), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5927) );
  NAND2_X1 U7522 ( .A1(n6150), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5926) );
  NOR2_X1 U7523 ( .A1(n8101), .A2(n6828), .ZN(n5930) );
  NAND2_X1 U7524 ( .A1(n5929), .A2(n5930), .ZN(n5934) );
  INV_X1 U7525 ( .A(n5929), .ZN(n8102) );
  INV_X1 U7526 ( .A(n5930), .ZN(n5931) );
  NAND2_X1 U7527 ( .A1(n8102), .A2(n5931), .ZN(n5932) );
  NAND2_X1 U7528 ( .A1(n5934), .A2(n5932), .ZN(n8172) );
  INV_X1 U7529 ( .A(n8172), .ZN(n5933) );
  NAND2_X1 U7530 ( .A1(n8169), .A2(n5934), .ZN(n5945) );
  NAND2_X1 U7531 ( .A1(n7335), .A2(n5713), .ZN(n5936) );
  NAND2_X1 U7532 ( .A1(n5887), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5935) );
  XNOR2_X1 U7533 ( .A(n8524), .B(n6024), .ZN(n5946) );
  INV_X1 U7534 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8107) );
  NAND2_X1 U7535 ( .A1(n5937), .A2(n8107), .ZN(n5938) );
  AND2_X1 U7536 ( .A1(n5954), .A2(n5938), .ZN(n8521) );
  NAND2_X1 U7537 ( .A1(n8521), .A2(n5640), .ZN(n5944) );
  INV_X1 U7538 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7539 ( .A1(n6151), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7540 ( .A1(n6152), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5939) );
  OAI211_X1 U7541 ( .C1(n5941), .C2(n5622), .A(n5940), .B(n5939), .ZN(n5942)
         );
  INV_X1 U7542 ( .A(n5942), .ZN(n5943) );
  NOR2_X1 U7543 ( .A1(n8539), .A2(n6828), .ZN(n5947) );
  XNOR2_X1 U7544 ( .A(n5946), .B(n5947), .ZN(n8099) );
  NAND2_X1 U7545 ( .A1(n5945), .A2(n8099), .ZN(n8103) );
  INV_X1 U7546 ( .A(n5946), .ZN(n5948) );
  NAND2_X1 U7547 ( .A1(n5948), .A2(n5947), .ZN(n5949) );
  NAND2_X1 U7548 ( .A1(n8103), .A2(n5949), .ZN(n5963) );
  NAND2_X1 U7549 ( .A1(n7392), .A2(n5713), .ZN(n5951) );
  NAND2_X1 U7550 ( .A1(n5887), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7551 ( .A(n8661), .B(n6045), .ZN(n5961) );
  INV_X1 U7552 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7553 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  NAND2_X1 U7554 ( .A1(n5977), .A2(n5955), .ZN(n8500) );
  OR2_X1 U7555 ( .A1(n8500), .A2(n6038), .ZN(n5960) );
  INV_X1 U7556 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9330) );
  NAND2_X1 U7557 ( .A1(n6151), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5957) );
  NAND2_X1 U7558 ( .A1(n6152), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5956) );
  OAI211_X1 U7559 ( .C1(n9330), .C2(n5622), .A(n5957), .B(n5956), .ZN(n5958)
         );
  INV_X1 U7560 ( .A(n5958), .ZN(n5959) );
  OR2_X1 U7561 ( .A1(n8106), .A2(n6828), .ZN(n8182) );
  INV_X1 U7562 ( .A(n5961), .ZN(n5962) );
  OR2_X1 U7563 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  NAND2_X1 U7564 ( .A1(n7449), .A2(n5713), .ZN(n5967) );
  NAND2_X1 U7565 ( .A1(n5887), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5966) );
  XNOR2_X1 U7566 ( .A(n8656), .B(n6024), .ZN(n5987) );
  NAND2_X1 U7567 ( .A1(n7463), .A2(n5713), .ZN(n5969) );
  NAND2_X1 U7568 ( .A1(n5887), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n5968) );
  XNOR2_X1 U7569 ( .A(n8650), .B(n6045), .ZN(n8146) );
  INV_X1 U7570 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U7571 ( .A1(n5979), .A2(n8151), .ZN(n5971) );
  NAND2_X1 U7572 ( .A1(n5998), .A2(n5971), .ZN(n8464) );
  OR2_X1 U7573 ( .A1(n8464), .A2(n6038), .ZN(n5976) );
  INV_X1 U7574 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U7575 ( .A1(n6151), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7576 ( .A1(n6152), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5972) );
  OAI211_X1 U7577 ( .C1(n9313), .C2(n5622), .A(n5973), .B(n5972), .ZN(n5974)
         );
  INV_X1 U7578 ( .A(n5974), .ZN(n5975) );
  INV_X1 U7579 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U7580 ( .A1(n5977), .A2(n8055), .ZN(n5978) );
  NAND2_X1 U7581 ( .A1(n5979), .A2(n5978), .ZN(n8488) );
  OR2_X1 U7582 ( .A1(n8488), .A2(n6038), .ZN(n5985) );
  INV_X1 U7583 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U7584 ( .A1(n6151), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7585 ( .A1(n6152), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5980) );
  OAI211_X1 U7586 ( .C1(n5982), .C2(n5622), .A(n5981), .B(n5980), .ZN(n5983)
         );
  INV_X1 U7587 ( .A(n5983), .ZN(n5984) );
  OR2_X1 U7588 ( .A1(n8506), .A2(n6828), .ZN(n8053) );
  AOI21_X1 U7589 ( .B1(n8146), .B2(n8220), .A(n8053), .ZN(n5986) );
  NAND2_X1 U7590 ( .A1(n8052), .A2(n5986), .ZN(n5994) );
  NOR2_X1 U7591 ( .A1(n8220), .A2(n6828), .ZN(n5991) );
  INV_X1 U7592 ( .A(n8146), .ZN(n5990) );
  INV_X1 U7593 ( .A(n5991), .ZN(n8149) );
  NAND2_X1 U7594 ( .A1(n5887), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5995) );
  XNOR2_X1 U7595 ( .A(n8646), .B(n6024), .ZN(n8115) );
  INV_X1 U7596 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7597 ( .A1(n5998), .A2(n5997), .ZN(n5999) );
  NAND2_X1 U7598 ( .A1(n8451), .A2(n5640), .ZN(n6004) );
  INV_X1 U7599 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9382) );
  NAND2_X1 U7600 ( .A1(n6151), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6000) );
  OAI211_X1 U7601 ( .C1(n5674), .C2(n9382), .A(n6001), .B(n6000), .ZN(n6002)
         );
  INV_X1 U7602 ( .A(n6002), .ZN(n6003) );
  AND2_X1 U7603 ( .A1(n8472), .A2(n6171), .ZN(n6005) );
  AND2_X1 U7604 ( .A1(n8115), .A2(n6005), .ZN(n8114) );
  INV_X1 U7605 ( .A(n8115), .ZN(n6007) );
  INV_X1 U7606 ( .A(n6005), .ZN(n6006) );
  NAND2_X1 U7607 ( .A1(n6007), .A2(n6006), .ZN(n8117) );
  NAND2_X1 U7608 ( .A1(n7579), .A2(n5713), .ZN(n6009) );
  NAND2_X1 U7609 ( .A1(n5887), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6008) );
  XNOR2_X1 U7610 ( .A(n8642), .B(n6024), .ZN(n6020) );
  INV_X1 U7611 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7612 ( .A1(n6012), .A2(n6011), .ZN(n6013) );
  NAND2_X1 U7613 ( .A1(n6036), .A2(n6013), .ZN(n8432) );
  INV_X1 U7614 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U7615 ( .A1(n6150), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7616 ( .A1(n6151), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6014) );
  OAI211_X1 U7617 ( .C1(n5674), .C2(n9369), .A(n6015), .B(n6014), .ZN(n6016)
         );
  INV_X1 U7618 ( .A(n6016), .ZN(n6017) );
  NOR2_X1 U7619 ( .A1(n8111), .A2(n6828), .ZN(n6019) );
  XNOR2_X1 U7620 ( .A(n6020), .B(n6019), .ZN(n8206) );
  NAND2_X1 U7621 ( .A1(n6020), .A2(n6019), .ZN(n6021) );
  NAND2_X1 U7622 ( .A1(n5887), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6022) );
  XNOR2_X1 U7623 ( .A(n8636), .B(n6024), .ZN(n6033) );
  XNOR2_X1 U7624 ( .A(n6036), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U7625 ( .A1(n8416), .A2(n5640), .ZN(n6030) );
  INV_X1 U7626 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6027) );
  NAND2_X1 U7627 ( .A1(n6151), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6026) );
  NAND2_X1 U7628 ( .A1(n6152), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6025) );
  OAI211_X1 U7629 ( .C1(n6027), .C2(n5622), .A(n6026), .B(n6025), .ZN(n6028)
         );
  INV_X1 U7630 ( .A(n6028), .ZN(n6029) );
  NAND2_X1 U7631 ( .A1(n8219), .A2(n6171), .ZN(n6031) );
  XNOR2_X1 U7632 ( .A(n6033), .B(n6031), .ZN(n8043) );
  INV_X1 U7633 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7634 ( .A1(n6033), .A2(n6032), .ZN(n6034) );
  NAND2_X1 U7635 ( .A1(n6035), .A2(n6034), .ZN(n6048) );
  INV_X1 U7636 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8046) );
  INV_X1 U7637 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7638 ( .B1(n6036), .B2(n8046), .A(n6104), .ZN(n6037) );
  NAND2_X1 U7639 ( .A1(n6037), .A2(n6094), .ZN(n8398) );
  INV_X1 U7640 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7641 ( .A1(n6151), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6040) );
  NAND2_X1 U7642 ( .A1(n6152), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6039) );
  OAI211_X1 U7643 ( .C1(n6041), .C2(n5622), .A(n6040), .B(n6039), .ZN(n6042)
         );
  INV_X1 U7644 ( .A(n6042), .ZN(n6043) );
  NOR2_X1 U7645 ( .A1(n8045), .A2(n6828), .ZN(n6046) );
  XNOR2_X1 U7646 ( .A(n6046), .B(n6045), .ZN(n6047) );
  XNOR2_X1 U7647 ( .A(n6048), .B(n6047), .ZN(n6090) );
  INV_X1 U7648 ( .A(n6090), .ZN(n6083) );
  NAND2_X1 U7649 ( .A1(n6049), .A2(n5574), .ZN(n6050) );
  NAND2_X1 U7650 ( .A1(n6050), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6079) );
  INV_X1 U7651 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6078) );
  NAND2_X1 U7652 ( .A1(n6079), .A2(n6078), .ZN(n6081) );
  NAND2_X1 U7653 ( .A1(n6081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6052) );
  XNOR2_X1 U7654 ( .A(n7513), .B(P2_B_REG_SCAN_IN), .ZN(n6058) );
  NOR2_X1 U7655 ( .A1(n6053), .A2(n6055), .ZN(n6054) );
  MUX2_X1 U7656 ( .A(n6055), .B(n6054), .S(P2_IR_REG_25__SCAN_IN), .Z(n6056)
         );
  INV_X1 U7657 ( .A(n6056), .ZN(n6057) );
  NAND2_X1 U7658 ( .A1(n6057), .A2(n4485), .ZN(n7582) );
  NAND2_X1 U7659 ( .A1(n6058), .A2(n7582), .ZN(n6063) );
  NAND2_X1 U7660 ( .A1(n4485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6059) );
  MUX2_X1 U7661 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6059), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6061) );
  NAND2_X1 U7662 ( .A1(n6061), .A2(n6060), .ZN(n7587) );
  INV_X1 U7663 ( .A(n7587), .ZN(n6062) );
  NAND2_X1 U7664 ( .A1(n6063), .A2(n6062), .ZN(n9852) );
  OR2_X1 U7665 ( .A1(n9852), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7666 ( .A1(n7513), .A2(n7587), .ZN(n9857) );
  NAND2_X1 U7667 ( .A1(n6064), .A2(n9857), .ZN(n7050) );
  OR2_X1 U7668 ( .A1(n9852), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6066) );
  AND2_X1 U7669 ( .A1(n7582), .A2(n7587), .ZN(n9863) );
  INV_X1 U7670 ( .A(n9863), .ZN(n6065) );
  NOR2_X1 U7671 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6070) );
  NOR4_X1 U7672 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6069) );
  NOR4_X1 U7673 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n6068) );
  NOR4_X1 U7674 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n6067) );
  NAND4_X1 U7675 ( .A1(n6070), .A2(n6069), .A3(n6068), .A4(n6067), .ZN(n6076)
         );
  NOR4_X1 U7676 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6074) );
  NOR4_X1 U7677 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6073) );
  NOR4_X1 U7678 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6072) );
  NOR4_X1 U7679 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_23__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6071) );
  NAND4_X1 U7680 ( .A1(n6074), .A2(n6073), .A3(n6072), .A4(n6071), .ZN(n6075)
         );
  NOR2_X1 U7681 ( .A1(n6076), .A2(n6075), .ZN(n6077) );
  OR2_X1 U7682 ( .A1(n9852), .A2(n6077), .ZN(n6797) );
  NAND2_X1 U7683 ( .A1(n6799), .A2(n6797), .ZN(n7038) );
  OR2_X1 U7684 ( .A1(n7050), .A2(n7038), .ZN(n6100) );
  OR2_X1 U7685 ( .A1(n6079), .A2(n6078), .ZN(n6080) );
  NAND2_X1 U7686 ( .A1(n6081), .A2(n6080), .ZN(n6324) );
  INV_X1 U7687 ( .A(n9851), .ZN(n6329) );
  NOR2_X1 U7688 ( .A1(n6100), .A2(n6329), .ZN(n6091) );
  AND2_X1 U7689 ( .A1(n7309), .A2(n8443), .ZN(n6101) );
  INV_X1 U7690 ( .A(n6101), .ZN(n6328) );
  NAND2_X1 U7691 ( .A1(n5580), .A2(n6319), .ZN(n6704) );
  INV_X1 U7692 ( .A(n6704), .ZN(n6620) );
  NOR2_X1 U7693 ( .A1(n9927), .A2(n6620), .ZN(n6082) );
  NOR2_X1 U7694 ( .A1(n6083), .A2(n8216), .ZN(n6086) );
  NAND2_X1 U7695 ( .A1(n8721), .A2(n5713), .ZN(n6085) );
  NAND2_X1 U7696 ( .A1(n5887), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6084) );
  INV_X1 U7697 ( .A(n8630), .ZN(n8401) );
  NAND2_X1 U7698 ( .A1(n6086), .A2(n8401), .ZN(n6111) );
  OR2_X1 U7699 ( .A1(n6087), .A2(n7309), .ZN(n8433) );
  INV_X1 U7700 ( .A(n8433), .ZN(n6089) );
  NAND2_X1 U7701 ( .A1(n9927), .A2(n8433), .ZN(n6796) );
  INV_X1 U7702 ( .A(n6796), .ZN(n6088) );
  AND2_X2 U7703 ( .A1(n9851), .A2(n6088), .ZN(n9839) );
  AOI21_X2 U7704 ( .B1(n6091), .B2(n6089), .A(n9839), .ZN(n8190) );
  OAI21_X1 U7705 ( .B1(n6090), .B2(n8216), .A(n8190), .ZN(n6109) );
  INV_X1 U7706 ( .A(n8219), .ZN(n8406) );
  NAND2_X1 U7707 ( .A1(n6091), .A2(n6101), .ZN(n8212) );
  INV_X1 U7708 ( .A(n6092), .ZN(n6093) );
  OR2_X1 U7709 ( .A1(n8212), .A2(n8536), .ZN(n8200) );
  INV_X1 U7710 ( .A(n6094), .ZN(n8007) );
  INV_X1 U7711 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7712 ( .A1(n6152), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7713 ( .A1(n6151), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6095) );
  OAI211_X1 U7714 ( .C1(n6097), .C2(n5622), .A(n6096), .B(n6095), .ZN(n6098)
         );
  AOI21_X1 U7715 ( .B1(n8007), .B2(n5640), .A(n6098), .ZN(n8405) );
  NAND2_X1 U7716 ( .A1(n6620), .A2(n6092), .ZN(n8538) );
  OR2_X1 U7717 ( .A1(n8212), .A2(n8538), .ZN(n8199) );
  OAI22_X1 U7718 ( .A1(n8406), .A2(n8200), .B1(n8405), .B2(n8199), .ZN(n6099)
         );
  INV_X1 U7719 ( .A(n6099), .ZN(n6107) );
  NAND2_X1 U7720 ( .A1(n6100), .A2(n6796), .ZN(n6763) );
  OR2_X1 U7721 ( .A1(n6704), .A2(n6101), .ZN(n6762) );
  AND3_X1 U7722 ( .A1(n6706), .A2(n6324), .A3(n6762), .ZN(n6102) );
  NAND2_X1 U7723 ( .A1(n6763), .A2(n6102), .ZN(n6103) );
  NAND2_X1 U7724 ( .A1(n6103), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8198) );
  OAI22_X1 U7725 ( .A1(n8398), .A2(n8198), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6104), .ZN(n6105) );
  INV_X1 U7726 ( .A(n6105), .ZN(n6106) );
  NAND2_X1 U7727 ( .A1(n6107), .A2(n6106), .ZN(n6108) );
  NAND2_X1 U7728 ( .A1(n6111), .A2(n6110), .ZN(P2_U3222) );
  NAND2_X1 U7729 ( .A1(n6319), .A2(n6806), .ZN(n6810) );
  INV_X1 U7730 ( .A(n6829), .ZN(n6113) );
  NAND2_X1 U7731 ( .A1(n9832), .A2(n6297), .ZN(n6809) );
  INV_X1 U7732 ( .A(n8060), .ZN(n8237) );
  NAND2_X1 U7733 ( .A1(n8060), .A2(n6807), .ZN(n6183) );
  NAND2_X1 U7734 ( .A1(n6181), .A2(n6183), .ZN(n6808) );
  OAI21_X1 U7735 ( .B1(n6809), .B2(n6808), .A(n6183), .ZN(n6871) );
  XNOR2_X1 U7736 ( .A(n8236), .B(n6115), .ZN(n6300) );
  INV_X1 U7737 ( .A(n8236), .ZN(n7103) );
  NAND2_X1 U7738 ( .A1(n7103), .A2(n6115), .ZN(n6175) );
  NAND2_X1 U7739 ( .A1(n7020), .A2(n7098), .ZN(n6299) );
  INV_X1 U7740 ( .A(n7020), .ZN(n8235) );
  INV_X1 U7741 ( .A(n7098), .ZN(n9877) );
  NAND2_X1 U7742 ( .A1(n8235), .A2(n9877), .ZN(n7024) );
  INV_X1 U7743 ( .A(n8157), .ZN(n8234) );
  INV_X1 U7744 ( .A(n7031), .ZN(n7060) );
  NAND2_X1 U7745 ( .A1(n7025), .A2(n6173), .ZN(n6116) );
  NAND2_X1 U7746 ( .A1(n8157), .A2(n7031), .ZN(n6295) );
  NAND2_X1 U7747 ( .A1(n6116), .A2(n6295), .ZN(n7045) );
  INV_X1 U7748 ( .A(n7118), .ZN(n8233) );
  INV_X2 U7749 ( .A(n7109), .ZN(n9883) );
  XNOR2_X1 U7750 ( .A(n8233), .B(n9883), .ZN(n7044) );
  NAND2_X1 U7751 ( .A1(n7118), .A2(n9883), .ZN(n6176) );
  AND2_X1 U7752 ( .A1(n8088), .A2(n8039), .ZN(n6117) );
  INV_X1 U7753 ( .A(n8088), .ZN(n8232) );
  NAND2_X1 U7754 ( .A1(n9893), .A2(n8232), .ZN(n6118) );
  OR2_X1 U7755 ( .A1(n8094), .A2(n7262), .ZN(n6205) );
  NAND2_X1 U7756 ( .A1(n8094), .A2(n7262), .ZN(n6204) );
  NAND2_X1 U7757 ( .A1(n7171), .A2(n7251), .ZN(n7170) );
  OR2_X1 U7758 ( .A1(n7354), .A2(n7359), .ZN(n6304) );
  NAND2_X1 U7759 ( .A1(n7354), .A2(n7359), .ZN(n6303) );
  OR2_X1 U7760 ( .A1(n7397), .A2(n7404), .ZN(n6293) );
  NAND2_X1 U7761 ( .A1(n7397), .A2(n7404), .ZN(n6292) );
  OR2_X1 U7762 ( .A1(n7589), .A2(n7588), .ZN(n6291) );
  NAND2_X1 U7763 ( .A1(n7401), .A2(n6291), .ZN(n9799) );
  NAND2_X1 U7764 ( .A1(n9928), .A2(n7600), .ZN(n6306) );
  NAND2_X1 U7765 ( .A1(n7589), .A2(n7588), .ZN(n9798) );
  AND2_X1 U7766 ( .A1(n6306), .A2(n9798), .ZN(n6218) );
  NAND2_X1 U7767 ( .A1(n9799), .A2(n6218), .ZN(n6119) );
  OR2_X1 U7768 ( .A1(n7614), .A2(n7619), .ZN(n6222) );
  NAND2_X1 U7769 ( .A1(n7614), .A2(n7619), .ZN(n6221) );
  NAND2_X1 U7770 ( .A1(n7620), .A2(n8225), .ZN(n6121) );
  INV_X1 U7771 ( .A(n7616), .ZN(n6122) );
  INV_X1 U7772 ( .A(n8225), .ZN(n7601) );
  OR2_X1 U7773 ( .A1(n7620), .A2(n7601), .ZN(n6228) );
  NAND2_X1 U7774 ( .A1(n6123), .A2(n6228), .ZN(n8605) );
  NOR2_X1 U7775 ( .A1(n7976), .A2(n8126), .ZN(n6226) );
  OR2_X1 U7776 ( .A1(n8692), .A2(n8137), .ZN(n6233) );
  NAND2_X1 U7777 ( .A1(n8598), .A2(n6233), .ZN(n6124) );
  NAND2_X1 U7778 ( .A1(n8692), .A2(n8137), .ZN(n6232) );
  NAND2_X1 U7779 ( .A1(n8687), .A2(n8570), .ZN(n6125) );
  NAND2_X1 U7780 ( .A1(n7992), .A2(n6125), .ZN(n8584) );
  INV_X1 U7781 ( .A(n8584), .ZN(n6126) );
  INV_X1 U7782 ( .A(n8570), .ZN(n8201) );
  OR2_X1 U7783 ( .A1(n8687), .A2(n8201), .ZN(n6236) );
  NAND2_X1 U7784 ( .A1(n8681), .A2(n8138), .ZN(n6242) );
  INV_X1 U7785 ( .A(n8573), .ZN(n8537) );
  OR2_X1 U7786 ( .A1(n8677), .A2(n8537), .ZN(n6254) );
  NAND2_X1 U7787 ( .A1(n8677), .A2(n8537), .ZN(n6251) );
  NAND2_X1 U7788 ( .A1(n6254), .A2(n6251), .ZN(n8555) );
  INV_X1 U7789 ( .A(n8554), .ZN(n6127) );
  NOR2_X1 U7790 ( .A1(n8555), .A2(n6127), .ZN(n6128) );
  NAND2_X1 U7791 ( .A1(n8567), .A2(n6128), .ZN(n6129) );
  NAND2_X1 U7792 ( .A1(n8671), .A2(n8101), .ZN(n6256) );
  NAND2_X1 U7793 ( .A1(n8515), .A2(n6256), .ZN(n8534) );
  OR2_X1 U7794 ( .A1(n8668), .A2(n8539), .ZN(n6260) );
  NAND2_X1 U7795 ( .A1(n8668), .A2(n8539), .ZN(n6255) );
  NAND2_X1 U7796 ( .A1(n6260), .A2(n6255), .ZN(n8517) );
  INV_X1 U7797 ( .A(n8515), .ZN(n6131) );
  NOR2_X1 U7798 ( .A1(n8517), .A2(n6131), .ZN(n6132) );
  NAND2_X1 U7799 ( .A1(n6133), .A2(n6255), .ZN(n8505) );
  NAND2_X1 U7800 ( .A1(n8661), .A2(n8106), .ZN(n6245) );
  NAND2_X1 U7801 ( .A1(n8656), .A2(n8506), .ZN(n6250) );
  INV_X1 U7802 ( .A(n8482), .ZN(n8479) );
  NAND2_X1 U7803 ( .A1(n8650), .A2(n8220), .ZN(n6266) );
  NAND2_X1 U7804 ( .A1(n8470), .A2(n8469), .ZN(n8468) );
  NAND2_X1 U7805 ( .A1(n8468), .A2(n6264), .ZN(n8454) );
  INV_X1 U7806 ( .A(n8472), .ZN(n8152) );
  NOR2_X1 U7807 ( .A1(n8646), .A2(n8152), .ZN(n8435) );
  NOR2_X1 U7808 ( .A1(n8439), .A2(n8435), .ZN(n6136) );
  NAND2_X1 U7809 ( .A1(n8458), .A2(n6136), .ZN(n8419) );
  NAND2_X1 U7810 ( .A1(n8419), .A2(n6137), .ZN(n8420) );
  OR2_X1 U7811 ( .A1(n8636), .A2(n8406), .ZN(n6272) );
  NAND2_X1 U7812 ( .A1(n8420), .A2(n6272), .ZN(n8402) );
  NAND2_X1 U7813 ( .A1(n8630), .A2(n8045), .ZN(n6278) );
  NAND2_X1 U7814 ( .A1(n6273), .A2(n6278), .ZN(n8403) );
  NAND2_X1 U7815 ( .A1(n8717), .A2(n5713), .ZN(n6139) );
  NAND2_X1 U7816 ( .A1(n5887), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7817 ( .A1(n8628), .A2(n8405), .ZN(n6281) );
  INV_X1 U7818 ( .A(SI_29_), .ZN(n6140) );
  AND2_X1 U7819 ( .A1(n6143), .A2(n6140), .ZN(n6141) );
  INV_X1 U7820 ( .A(n6143), .ZN(n6144) );
  NAND2_X1 U7821 ( .A1(n6144), .A2(SI_29_), .ZN(n6145) );
  MUX2_X1 U7822 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6567), .Z(n6156) );
  INV_X1 U7823 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n7980) );
  NOR2_X1 U7824 ( .A1(n5629), .A2(n7980), .ZN(n6147) );
  INV_X1 U7825 ( .A(n8625), .ZN(n8390) );
  INV_X1 U7826 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U7827 ( .A1(n6151), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6148) );
  OAI211_X1 U7828 ( .C1(n5674), .C2(n9356), .A(n6149), .B(n6148), .ZN(n8218)
         );
  AND2_X1 U7829 ( .A1(n8625), .A2(n8218), .ZN(n6284) );
  NAND2_X1 U7830 ( .A1(n6150), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7831 ( .A1(n6151), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7832 ( .A1(n6152), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6153) );
  AND3_X1 U7833 ( .A1(n6155), .A2(n6154), .A3(n6153), .ZN(n6166) );
  INV_X1 U7834 ( .A(n6166), .ZN(n8383) );
  INV_X1 U7835 ( .A(SI_30_), .ZN(n6159) );
  NAND2_X1 U7836 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  MUX2_X1 U7837 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6567), .Z(n6161) );
  XNOR2_X1 U7838 ( .A(n6161), .B(SI_31_), .ZN(n6162) );
  NAND2_X1 U7839 ( .A1(n9405), .A2(n5713), .ZN(n6165) );
  INV_X1 U7840 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8712) );
  OR2_X1 U7841 ( .A1(n5629), .A2(n8712), .ZN(n6164) );
  INV_X1 U7842 ( .A(n8218), .ZN(n6167) );
  NAND2_X1 U7843 ( .A1(n6287), .A2(n4294), .ZN(n6317) );
  INV_X1 U7844 ( .A(n6317), .ZN(n6168) );
  NAND2_X1 U7845 ( .A1(n6319), .A2(n8377), .ZN(n6172) );
  INV_X1 U7846 ( .A(n6279), .ZN(n6288) );
  INV_X1 U7847 ( .A(n6245), .ZN(n6249) );
  AND2_X1 U7848 ( .A1(n6295), .A2(n6299), .ZN(n6174) );
  NAND2_X1 U7849 ( .A1(n6299), .A2(n6175), .ZN(n6178) );
  NAND2_X1 U7850 ( .A1(n6295), .A2(n6176), .ZN(n6177) );
  AOI21_X1 U7851 ( .B1(n6191), .B2(n6178), .A(n6177), .ZN(n6189) );
  NAND2_X1 U7852 ( .A1(n6829), .A2(n6833), .ZN(n6296) );
  NAND2_X1 U7853 ( .A1(n6297), .A2(n6296), .ZN(n6179) );
  NAND3_X1 U7854 ( .A1(n6183), .A2(n6298), .A3(n6179), .ZN(n6180) );
  NAND2_X1 U7855 ( .A1(n6180), .A2(n6181), .ZN(n6186) );
  AND2_X1 U7856 ( .A1(n6296), .A2(n6319), .ZN(n6182) );
  OAI211_X1 U7857 ( .C1(n9832), .C2(n6182), .A(n6297), .B(n6181), .ZN(n6184)
         );
  NAND2_X1 U7858 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  MUX2_X1 U7859 ( .A(n6186), .B(n6185), .S(n6279), .Z(n6187) );
  NAND3_X1 U7860 ( .A1(n6187), .A2(n6191), .A3(n6300), .ZN(n6188) );
  OAI21_X1 U7861 ( .B1(n6189), .B2(n6288), .A(n6188), .ZN(n6190) );
  OR2_X1 U7862 ( .A1(n7118), .A2(n9883), .ZN(n6193) );
  NAND2_X1 U7863 ( .A1(n6190), .A2(n6193), .ZN(n6198) );
  NAND2_X1 U7864 ( .A1(n8236), .A2(n9818), .ZN(n6192) );
  AND2_X1 U7865 ( .A1(n7024), .A2(n6192), .ZN(n6194) );
  OAI211_X1 U7866 ( .C1(n6195), .C2(n6194), .A(n6294), .B(n6193), .ZN(n6196)
         );
  NAND2_X1 U7867 ( .A1(n6196), .A2(n6288), .ZN(n6197) );
  NAND2_X1 U7868 ( .A1(n6198), .A2(n6197), .ZN(n6200) );
  XNOR2_X1 U7869 ( .A(n8088), .B(n8039), .ZN(n7167) );
  INV_X1 U7870 ( .A(n7167), .ZN(n7117) );
  NAND3_X1 U7871 ( .A1(n7118), .A2(n6288), .A3(n9883), .ZN(n6199) );
  NAND3_X1 U7872 ( .A1(n6200), .A2(n7117), .A3(n6199), .ZN(n6203) );
  MUX2_X1 U7873 ( .A(n8232), .B(n8039), .S(n6279), .Z(n6201) );
  OAI21_X1 U7874 ( .B1(n9893), .B2(n8088), .A(n6201), .ZN(n6202) );
  NAND3_X1 U7875 ( .A1(n6203), .A2(n7251), .A3(n6202), .ZN(n6208) );
  MUX2_X1 U7876 ( .A(n6205), .B(n6204), .S(n6288), .Z(n6206) );
  AND2_X1 U7877 ( .A1(n6206), .A2(n6303), .ZN(n6207) );
  NAND2_X1 U7878 ( .A1(n6208), .A2(n6207), .ZN(n6211) );
  NAND3_X1 U7879 ( .A1(n6211), .A2(n6304), .A3(n6293), .ZN(n6209) );
  NAND3_X1 U7880 ( .A1(n6209), .A2(n9798), .A3(n6292), .ZN(n6214) );
  INV_X1 U7881 ( .A(n6304), .ZN(n6210) );
  AOI21_X1 U7882 ( .B1(n6211), .B2(n6303), .A(n6210), .ZN(n6212) );
  OAI211_X1 U7883 ( .C1(n6212), .C2(n4562), .A(n6291), .B(n6293), .ZN(n6213)
         );
  MUX2_X1 U7884 ( .A(n6214), .B(n6213), .S(n6279), .Z(n6219) );
  AND2_X1 U7885 ( .A1(n6219), .A2(n6291), .ZN(n6216) );
  INV_X1 U7886 ( .A(n6306), .ZN(n6215) );
  INV_X1 U7887 ( .A(n6307), .ZN(n6217) );
  AOI21_X1 U7888 ( .B1(n6219), .B2(n6218), .A(n6217), .ZN(n6220) );
  MUX2_X1 U7889 ( .A(n6222), .B(n6221), .S(n6279), .Z(n6223) );
  NAND3_X1 U7890 ( .A1(n6224), .A2(n7601), .A3(n7620), .ZN(n6225) );
  OAI21_X1 U7891 ( .B1(n9463), .B2(n4668), .A(n6225), .ZN(n6230) );
  INV_X1 U7892 ( .A(n6226), .ZN(n6227) );
  OAI21_X1 U7893 ( .B1(n8608), .B2(n6228), .A(n6227), .ZN(n6229) );
  NAND2_X1 U7894 ( .A1(n6233), .A2(n6232), .ZN(n8597) );
  MUX2_X1 U7895 ( .A(n6233), .B(n6232), .S(n6279), .Z(n6234) );
  NAND2_X1 U7896 ( .A1(n8584), .A2(n6234), .ZN(n6239) );
  INV_X1 U7897 ( .A(n6242), .ZN(n6235) );
  AOI21_X1 U7898 ( .B1(n8201), .B2(n8687), .A(n6235), .ZN(n6237) );
  OAI211_X1 U7899 ( .C1(n6240), .C2(n6239), .A(n6238), .B(n8554), .ZN(n6253)
         );
  INV_X1 U7900 ( .A(n6254), .ZN(n6241) );
  AOI21_X1 U7901 ( .B1(n6253), .B2(n6242), .A(n6241), .ZN(n6244) );
  NAND2_X1 U7902 ( .A1(n6256), .A2(n6251), .ZN(n6243) );
  NAND3_X1 U7903 ( .A1(n6246), .A2(n6255), .A3(n6245), .ZN(n6247) );
  NAND2_X1 U7904 ( .A1(n6247), .A2(n6259), .ZN(n6248) );
  INV_X1 U7905 ( .A(n6251), .ZN(n6252) );
  AOI21_X1 U7906 ( .B1(n6253), .B2(n8554), .A(n6252), .ZN(n6258) );
  NAND2_X1 U7907 ( .A1(n8515), .A2(n6254), .ZN(n6257) );
  OAI211_X1 U7908 ( .C1(n6258), .C2(n6257), .A(n6256), .B(n6255), .ZN(n6261)
         );
  NAND4_X1 U7909 ( .A1(n6261), .A2(n6288), .A3(n6260), .A4(n6259), .ZN(n6262)
         );
  AOI21_X1 U7910 ( .B1(n6264), .B2(n6263), .A(n6279), .ZN(n6265) );
  INV_X1 U7911 ( .A(n7997), .ZN(n8455) );
  INV_X1 U7912 ( .A(n8646), .ZN(n8453) );
  NAND3_X1 U7913 ( .A1(n8453), .A2(n6288), .A3(n8472), .ZN(n6267) );
  OAI21_X1 U7914 ( .B1(n8453), .B2(n8472), .A(n8421), .ZN(n6268) );
  AOI22_X1 U7915 ( .A1(n6269), .A2(n8421), .B1(n6279), .B2(n6268), .ZN(n6276)
         );
  OAI21_X1 U7916 ( .B1(n6288), .B2(n6270), .A(n8422), .ZN(n6275) );
  INV_X1 U7917 ( .A(n6278), .ZN(n6271) );
  INV_X1 U7918 ( .A(n6280), .ZN(n6277) );
  MUX2_X1 U7919 ( .A(n6281), .B(n6280), .S(n6279), .Z(n6282) );
  NOR2_X1 U7920 ( .A1(n6285), .A2(n6284), .ZN(n6290) );
  INV_X1 U7921 ( .A(n6290), .ZN(n6316) );
  INV_X1 U7922 ( .A(n8469), .ZN(n6313) );
  INV_X1 U7923 ( .A(n8555), .ZN(n8546) );
  NAND2_X1 U7924 ( .A1(n6291), .A2(n9798), .ZN(n7402) );
  AND2_X1 U7925 ( .A1(n6293), .A2(n6292), .ZN(n7396) );
  INV_X1 U7926 ( .A(n7396), .ZN(n7358) );
  NAND2_X1 U7927 ( .A1(n6295), .A2(n6294), .ZN(n7026) );
  NAND2_X1 U7928 ( .A1(n9827), .A2(n6296), .ZN(n9867) );
  NAND2_X1 U7929 ( .A1(n6298), .A2(n6297), .ZN(n6801) );
  OR4_X1 U7930 ( .A1(n6808), .A2(n9867), .A3(n6801), .A4(n7309), .ZN(n6301) );
  NAND2_X1 U7931 ( .A1(n6299), .A2(n7024), .ZN(n7100) );
  INV_X1 U7932 ( .A(n6300), .ZN(n6870) );
  NOR4_X1 U7933 ( .A1(n7026), .A2(n6301), .A3(n7100), .A4(n6870), .ZN(n6302)
         );
  NAND4_X1 U7934 ( .A1(n6302), .A2(n7251), .A3(n7117), .A4(n7044), .ZN(n6305)
         );
  INV_X1 U7935 ( .A(n7258), .ZN(n7260) );
  NOR4_X1 U7936 ( .A1(n7402), .A2(n7358), .A3(n6305), .A4(n7260), .ZN(n6308)
         );
  NAND3_X1 U7937 ( .A1(n7598), .A2(n6308), .A3(n9804), .ZN(n6309) );
  NOR4_X1 U7938 ( .A1(n8597), .A2(n8608), .A3(n7616), .A4(n6309), .ZN(n6310)
         );
  NAND4_X1 U7939 ( .A1(n8546), .A2(n8569), .A3(n6310), .A4(n8584), .ZN(n6311)
         );
  OR4_X1 U7940 ( .A1(n8504), .A2(n8517), .A3(n8534), .A4(n6311), .ZN(n6312) );
  NOR4_X1 U7941 ( .A1(n8439), .A2(n8482), .A3(n6313), .A4(n6312), .ZN(n6314)
         );
  NAND4_X1 U7942 ( .A1(n8394), .A2(n6314), .A3(n7997), .A4(n8422), .ZN(n6315)
         );
  NOR4_X1 U7943 ( .A1(n6317), .A2(n6316), .A3(n8002), .A4(n6315), .ZN(n6318)
         );
  XNOR2_X1 U7944 ( .A(n6318), .B(n8377), .ZN(n6320) );
  OAI22_X1 U7945 ( .A1(n6320), .A2(n6319), .B1(n6806), .B2(n6811), .ZN(n6322)
         );
  OR2_X1 U7946 ( .A1(n6324), .A2(P2_U3152), .ZN(n6705) );
  NOR4_X1 U7947 ( .A1(n6329), .A2(n8004), .A3(n6328), .A4(n8536), .ZN(n6331)
         );
  OAI21_X1 U7948 ( .B1(n6705), .B2(n5580), .A(P2_B_REG_SCAN_IN), .ZN(n6330) );
  NAND2_X1 U7949 ( .A1(n6335), .A2(n4244), .ZN(n6337) );
  NAND2_X1 U7950 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  INV_X1 U7951 ( .A(n6339), .ZN(n6341) );
  INV_X1 U7952 ( .A(n7393), .ZN(n6340) );
  NAND2_X1 U7953 ( .A1(n6374), .A2(n6335), .ZN(n6344) );
  NAND2_X1 U7954 ( .A1(n6851), .A2(n4244), .ZN(n6343) );
  NAND2_X1 U7955 ( .A1(n6344), .A2(n6343), .ZN(n6354) );
  NAND2_X1 U7956 ( .A1(n6353), .A2(n6354), .ZN(n6352) );
  INV_X1 U7957 ( .A(n7080), .ZN(n6771) );
  INV_X1 U7958 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6628) );
  OAI22_X1 U7959 ( .A1(n6771), .A2(n6357), .B1(n6590), .B2(n6628), .ZN(n6345)
         );
  INV_X1 U7960 ( .A(n6689), .ZN(n6350) );
  NAND2_X1 U7961 ( .A1(n6374), .A2(n6346), .ZN(n6349) );
  INV_X1 U7962 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6629) );
  NOR2_X1 U7963 ( .A1(n6590), .A2(n6629), .ZN(n6347) );
  AOI21_X1 U7964 ( .B1(n7080), .B2(n4244), .A(n6347), .ZN(n6348) );
  NAND2_X1 U7965 ( .A1(n6689), .A2(n4266), .ZN(n6351) );
  NAND2_X1 U7966 ( .A1(n6352), .A2(n6695), .ZN(n6356) );
  INV_X1 U7967 ( .A(n6354), .ZN(n6696) );
  NAND2_X1 U7968 ( .A1(n6697), .A2(n6696), .ZN(n6355) );
  NAND2_X1 U7969 ( .A1(n6356), .A2(n6355), .ZN(n6750) );
  INV_X1 U7970 ( .A(n4266), .ZN(n6362) );
  NAND2_X1 U7971 ( .A1(n6363), .A2(n4244), .ZN(n6360) );
  NAND2_X1 U7972 ( .A1(n6374), .A2(n6363), .ZN(n6365) );
  NAND2_X1 U7973 ( .A1(n6358), .A2(n4244), .ZN(n6364) );
  NAND2_X1 U7974 ( .A1(n6365), .A2(n6364), .ZN(n6366) );
  XNOR2_X1 U7975 ( .A(n6368), .B(n6366), .ZN(n6751) );
  NAND2_X1 U7976 ( .A1(n6750), .A2(n6751), .ZN(n6370) );
  INV_X1 U7977 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U7978 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  NAND2_X1 U7979 ( .A1(n6370), .A2(n6369), .ZN(n6821) );
  NAND2_X1 U7980 ( .A1(n8870), .A2(n4244), .ZN(n6372) );
  NAND2_X1 U7981 ( .A1(n6375), .A2(n4247), .ZN(n6371) );
  NAND2_X1 U7982 ( .A1(n6372), .A2(n6371), .ZN(n6373) );
  XNOR2_X1 U7983 ( .A(n6373), .B(n6362), .ZN(n6380) );
  INV_X2 U7984 ( .A(n6440), .ZN(n8013) );
  NAND2_X1 U7985 ( .A1(n8013), .A2(n8870), .ZN(n6377) );
  NAND2_X1 U7986 ( .A1(n6375), .A2(n4244), .ZN(n6376) );
  NAND2_X1 U7987 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  XNOR2_X1 U7988 ( .A(n6380), .B(n6378), .ZN(n6822) );
  NAND2_X1 U7989 ( .A1(n6821), .A2(n6822), .ZN(n6857) );
  INV_X1 U7990 ( .A(n6378), .ZN(n6379) );
  NAND2_X1 U7991 ( .A1(n6380), .A2(n6379), .ZN(n6858) );
  NAND2_X1 U7992 ( .A1(n7210), .A2(n4247), .ZN(n6381) );
  INV_X2 U7993 ( .A(n6440), .ZN(n6528) );
  NAND2_X1 U7994 ( .A1(n6528), .A2(n8869), .ZN(n6385) );
  NAND2_X1 U7995 ( .A1(n7210), .A2(n4244), .ZN(n6384) );
  NAND2_X1 U7996 ( .A1(n6385), .A2(n6384), .ZN(n6388) );
  INV_X1 U7997 ( .A(n6388), .ZN(n6386) );
  NAND2_X1 U7998 ( .A1(n6389), .A2(n6386), .ZN(n6391) );
  AND2_X1 U7999 ( .A1(n6858), .A2(n6391), .ZN(n6387) );
  NAND2_X1 U8000 ( .A1(n6857), .A2(n6387), .ZN(n6393) );
  INV_X1 U8001 ( .A(n6860), .ZN(n6390) );
  NAND2_X1 U8002 ( .A1(n6391), .A2(n6390), .ZN(n6392) );
  NAND2_X1 U8003 ( .A1(n8868), .A2(n4244), .ZN(n6395) );
  NAND2_X1 U8004 ( .A1(n6397), .A2(n4247), .ZN(n6394) );
  NAND2_X1 U8005 ( .A1(n6395), .A2(n6394), .ZN(n6396) );
  XNOR2_X1 U8006 ( .A(n6396), .B(n4266), .ZN(n6399) );
  AND2_X1 U8007 ( .A1(n6397), .A2(n4244), .ZN(n6398) );
  AOI21_X1 U8008 ( .B1(n6528), .B2(n8868), .A(n6398), .ZN(n7011) );
  NAND2_X1 U8009 ( .A1(n8867), .A2(n4244), .ZN(n6402) );
  NAND2_X1 U8010 ( .A1(n8817), .A2(n4247), .ZN(n6401) );
  NAND2_X1 U8011 ( .A1(n6402), .A2(n6401), .ZN(n6403) );
  XNOR2_X1 U8012 ( .A(n6403), .B(n6362), .ZN(n6408) );
  NAND2_X1 U8013 ( .A1(n8013), .A2(n8867), .ZN(n6405) );
  NAND2_X1 U8014 ( .A1(n8817), .A2(n4244), .ZN(n6404) );
  NAND2_X1 U8015 ( .A1(n6405), .A2(n6404), .ZN(n6406) );
  XNOR2_X1 U8016 ( .A(n6408), .B(n6406), .ZN(n8815) );
  INV_X1 U8017 ( .A(n6406), .ZN(n6407) );
  NAND2_X1 U8018 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  NAND2_X1 U8019 ( .A1(n8866), .A2(n4244), .ZN(n6411) );
  NAND2_X1 U8020 ( .A1(n7130), .A2(n4247), .ZN(n6410) );
  NAND2_X1 U8021 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  XNOR2_X1 U8022 ( .A(n6412), .B(n6362), .ZN(n6413) );
  OAI22_X1 U8023 ( .A1(n6440), .A2(n7292), .B1(n9755), .B2(n8017), .ZN(n6414)
         );
  XNOR2_X1 U8024 ( .A(n6413), .B(n6414), .ZN(n7087) );
  INV_X1 U8025 ( .A(n6413), .ZN(n6415) );
  NAND2_X1 U8026 ( .A1(n8013), .A2(n8865), .ZN(n6418) );
  NAND2_X1 U8027 ( .A1(n7313), .A2(n4244), .ZN(n6417) );
  NAND2_X1 U8028 ( .A1(n6418), .A2(n6417), .ZN(n6420) );
  AOI22_X1 U8029 ( .A1(n7313), .A2(n4247), .B1(n4244), .B2(n8865), .ZN(n6419)
         );
  XNOR2_X1 U8030 ( .A(n6419), .B(n4266), .ZN(n7290) );
  AOI22_X1 U8031 ( .A1(n7705), .A2(n4247), .B1(n4244), .B2(n8864), .ZN(n6422)
         );
  XNOR2_X1 U8032 ( .A(n6422), .B(n4266), .ZN(n6424) );
  AOI22_X1 U8033 ( .A1(n7705), .A2(n4244), .B1(n8013), .B2(n8864), .ZN(n6423)
         );
  XNOR2_X1 U8034 ( .A(n6424), .B(n6423), .ZN(n7349) );
  NAND2_X1 U8035 ( .A1(n7416), .A2(n4247), .ZN(n6426) );
  NAND2_X1 U8036 ( .A1(n8863), .A2(n4244), .ZN(n6425) );
  NAND2_X1 U8037 ( .A1(n6426), .A2(n6425), .ZN(n6427) );
  XNOR2_X1 U8038 ( .A(n6427), .B(n4266), .ZN(n7426) );
  NAND2_X1 U8039 ( .A1(n7416), .A2(n4244), .ZN(n6429) );
  NAND2_X1 U8040 ( .A1(n8013), .A2(n8863), .ZN(n6428) );
  NAND2_X1 U8041 ( .A1(n6429), .A2(n6428), .ZN(n7425) );
  NAND2_X1 U8042 ( .A1(n7459), .A2(n4247), .ZN(n6433) );
  NAND2_X1 U8043 ( .A1(n8862), .A2(n4244), .ZN(n6432) );
  NAND2_X1 U8044 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  XNOR2_X1 U8045 ( .A(n6434), .B(n4266), .ZN(n6438) );
  NOR2_X1 U8046 ( .A1(n6440), .A2(n7499), .ZN(n6435) );
  AOI21_X1 U8047 ( .B1(n7459), .B2(n4244), .A(n6435), .ZN(n6436) );
  XNOR2_X1 U8048 ( .A(n6438), .B(n6436), .ZN(n7455) );
  INV_X1 U8049 ( .A(n6436), .ZN(n6437) );
  AOI22_X1 U8050 ( .A1(n7507), .A2(n4247), .B1(n4244), .B2(n8861), .ZN(n6439)
         );
  XOR2_X1 U8051 ( .A(n4266), .B(n6439), .Z(n6442) );
  INV_X1 U8052 ( .A(n7507), .ZN(n9548) );
  OAI22_X1 U8053 ( .A1(n9548), .A2(n8017), .B1(n9511), .B2(n6440), .ZN(n6441)
         );
  NOR2_X1 U8054 ( .A1(n6442), .A2(n6441), .ZN(n6443) );
  AOI21_X1 U8055 ( .B1(n6442), .B2(n6441), .A(n6443), .ZN(n7547) );
  INV_X1 U8056 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8057 ( .A1(n9486), .A2(n4247), .ZN(n6446) );
  NAND2_X1 U8058 ( .A1(n8860), .A2(n4244), .ZN(n6445) );
  NAND2_X1 U8059 ( .A1(n6446), .A2(n6445), .ZN(n6447) );
  XNOR2_X1 U8060 ( .A(n6447), .B(n4266), .ZN(n6451) );
  NAND2_X1 U8061 ( .A1(n9486), .A2(n4244), .ZN(n6449) );
  NAND2_X1 U8062 ( .A1(n8013), .A2(n8860), .ZN(n6448) );
  NAND2_X1 U8063 ( .A1(n6449), .A2(n6448), .ZN(n6450) );
  NAND2_X1 U8064 ( .A1(n6451), .A2(n6450), .ZN(n7570) );
  AOI22_X1 U8065 ( .A1(n7673), .A2(n4247), .B1(n4244), .B2(n8859), .ZN(n6452)
         );
  XOR2_X1 U8066 ( .A(n4266), .B(n6452), .Z(n6453) );
  AOI22_X1 U8067 ( .A1(n7673), .A2(n4244), .B1(n8013), .B2(n8859), .ZN(n7668)
         );
  AOI22_X1 U8068 ( .A1(n8851), .A2(n4247), .B1(n4244), .B2(n8858), .ZN(n6455)
         );
  XOR2_X1 U8069 ( .A(n4266), .B(n6455), .Z(n6456) );
  AOI22_X1 U8070 ( .A1(n8851), .A2(n4244), .B1(n6528), .B2(n8858), .ZN(n8841)
         );
  AOI22_X1 U8071 ( .A1(n8762), .A2(n4244), .B1(n8013), .B2(n8857), .ZN(n6461)
         );
  NAND2_X1 U8072 ( .A1(n8762), .A2(n4247), .ZN(n6458) );
  NAND2_X1 U8073 ( .A1(n8857), .A2(n4244), .ZN(n6457) );
  NAND2_X1 U8074 ( .A1(n6458), .A2(n6457), .ZN(n6459) );
  XNOR2_X1 U8075 ( .A(n6459), .B(n4266), .ZN(n6463) );
  XOR2_X1 U8076 ( .A(n6461), .B(n6463), .Z(n8755) );
  INV_X1 U8077 ( .A(n6461), .ZN(n6462) );
  NAND2_X1 U8078 ( .A1(n9243), .A2(n4247), .ZN(n6466) );
  NAND2_X1 U8079 ( .A1(n9155), .A2(n4244), .ZN(n6465) );
  NAND2_X1 U8080 ( .A1(n6466), .A2(n6465), .ZN(n6467) );
  XNOR2_X1 U8081 ( .A(n6467), .B(n4266), .ZN(n6470) );
  AOI22_X1 U8082 ( .A1(n9243), .A2(n4244), .B1(n8013), .B2(n9155), .ZN(n6468)
         );
  XNOR2_X1 U8083 ( .A(n6470), .B(n6468), .ZN(n8767) );
  INV_X1 U8084 ( .A(n6468), .ZN(n6469) );
  INV_X1 U8085 ( .A(n8804), .ZN(n6473) );
  AOI22_X1 U8086 ( .A1(n9236), .A2(n4247), .B1(n4244), .B2(n9138), .ZN(n6472)
         );
  XOR2_X1 U8087 ( .A(n4266), .B(n6472), .Z(n6474) );
  NAND2_X1 U8088 ( .A1(n6473), .A2(n6474), .ZN(n6476) );
  AOI22_X1 U8089 ( .A1(n9236), .A2(n4244), .B1(n6528), .B2(n9138), .ZN(n8801)
         );
  INV_X1 U8090 ( .A(n6474), .ZN(n8802) );
  NAND2_X1 U8091 ( .A1(n9232), .A2(n4247), .ZN(n6478) );
  NAND2_X1 U8092 ( .A1(n9153), .A2(n4244), .ZN(n6477) );
  NAND2_X1 U8093 ( .A1(n6478), .A2(n6477), .ZN(n6479) );
  XNOR2_X1 U8094 ( .A(n6479), .B(n6362), .ZN(n7982) );
  AND2_X1 U8095 ( .A1(n8013), .A2(n9153), .ZN(n6480) );
  AOI21_X1 U8096 ( .B1(n9232), .B2(n4244), .A(n6480), .ZN(n7983) );
  NOR2_X1 U8097 ( .A1(n7982), .A2(n7983), .ZN(n6481) );
  NAND2_X1 U8098 ( .A1(n9226), .A2(n4247), .ZN(n6483) );
  NAND2_X1 U8099 ( .A1(n9137), .A2(n4244), .ZN(n6482) );
  NAND2_X1 U8100 ( .A1(n6483), .A2(n6482), .ZN(n6484) );
  XNOR2_X1 U8101 ( .A(n6484), .B(n4266), .ZN(n6488) );
  NAND2_X1 U8102 ( .A1(n9226), .A2(n4244), .ZN(n6486) );
  NAND2_X1 U8103 ( .A1(n9137), .A2(n6528), .ZN(n6485) );
  NAND2_X1 U8104 ( .A1(n6486), .A2(n6485), .ZN(n6487) );
  NOR2_X1 U8105 ( .A1(n6488), .A2(n6487), .ZN(n6489) );
  AOI21_X1 U8106 ( .B1(n6488), .B2(n6487), .A(n6489), .ZN(n8784) );
  NAND2_X1 U8107 ( .A1(n9223), .A2(n4247), .ZN(n6491) );
  NAND2_X1 U8108 ( .A1(n9121), .A2(n4244), .ZN(n6490) );
  NAND2_X1 U8109 ( .A1(n6491), .A2(n6490), .ZN(n6492) );
  XNOR2_X1 U8110 ( .A(n6492), .B(n4266), .ZN(n6493) );
  AOI22_X1 U8111 ( .A1(n9223), .A2(n4244), .B1(n6528), .B2(n9121), .ZN(n6494)
         );
  XNOR2_X1 U8112 ( .A(n6493), .B(n6494), .ZN(n8735) );
  INV_X1 U8113 ( .A(n6493), .ZN(n6495) );
  NAND2_X1 U8114 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  AOI22_X1 U8115 ( .A1(n9216), .A2(n4244), .B1(n6528), .B2(n9071), .ZN(n6497)
         );
  AOI22_X1 U8116 ( .A1(n9216), .A2(n4247), .B1(n4244), .B2(n9071), .ZN(n6498)
         );
  XOR2_X1 U8117 ( .A(n4266), .B(n6498), .Z(n8794) );
  NAND2_X1 U8118 ( .A1(n9211), .A2(n4247), .ZN(n6500) );
  NAND2_X1 U8119 ( .A1(n9088), .A2(n4244), .ZN(n6499) );
  NAND2_X1 U8120 ( .A1(n6500), .A2(n6499), .ZN(n6501) );
  XNOR2_X1 U8121 ( .A(n6501), .B(n6362), .ZN(n6503) );
  AOI22_X1 U8122 ( .A1(n9211), .A2(n4244), .B1(n8013), .B2(n9088), .ZN(n8726)
         );
  INV_X1 U8123 ( .A(n6503), .ZN(n6504) );
  AOI22_X1 U8124 ( .A1(n9206), .A2(n4247), .B1(n4244), .B2(n9072), .ZN(n6506)
         );
  XNOR2_X1 U8125 ( .A(n6506), .B(n4266), .ZN(n6508) );
  AOI22_X1 U8126 ( .A1(n9206), .A2(n4244), .B1(n6528), .B2(n9072), .ZN(n6507)
         );
  NAND2_X1 U8127 ( .A1(n6508), .A2(n6507), .ZN(n6509) );
  OAI21_X1 U8128 ( .B1(n6508), .B2(n6507), .A(n6509), .ZN(n8775) );
  NAND2_X1 U8129 ( .A1(n9203), .A2(n4247), .ZN(n6511) );
  NAND2_X1 U8130 ( .A1(n9054), .A2(n4244), .ZN(n6510) );
  NAND2_X1 U8131 ( .A1(n6511), .A2(n6510), .ZN(n6512) );
  XNOR2_X1 U8132 ( .A(n6512), .B(n4266), .ZN(n6519) );
  AOI22_X1 U8133 ( .A1(n9203), .A2(n4244), .B1(n6528), .B2(n9054), .ZN(n6517)
         );
  XNOR2_X1 U8134 ( .A(n6519), .B(n6517), .ZN(n8744) );
  NAND2_X1 U8135 ( .A1(n9196), .A2(n4247), .ZN(n6514) );
  NAND2_X1 U8136 ( .A1(n8856), .A2(n4244), .ZN(n6513) );
  NAND2_X1 U8137 ( .A1(n6514), .A2(n6513), .ZN(n6515) );
  XNOR2_X1 U8138 ( .A(n6515), .B(n6362), .ZN(n6521) );
  AND2_X1 U8139 ( .A1(n8856), .A2(n6528), .ZN(n6516) );
  AOI21_X1 U8140 ( .B1(n9196), .B2(n4244), .A(n6516), .ZN(n6522) );
  XNOR2_X1 U8141 ( .A(n6521), .B(n6522), .ZN(n8825) );
  INV_X1 U8142 ( .A(n6517), .ZN(n6518) );
  NOR2_X1 U8143 ( .A1(n6519), .A2(n6518), .ZN(n8826) );
  NOR2_X1 U8144 ( .A1(n8825), .A2(n8826), .ZN(n6520) );
  INV_X1 U8145 ( .A(n6521), .ZN(n6524) );
  INV_X1 U8146 ( .A(n6522), .ZN(n6523) );
  NAND2_X1 U8147 ( .A1(n9191), .A2(n4247), .ZN(n6526) );
  NAND2_X1 U8148 ( .A1(n9021), .A2(n4244), .ZN(n6525) );
  NAND2_X1 U8149 ( .A1(n6526), .A2(n6525), .ZN(n6527) );
  XNOR2_X1 U8150 ( .A(n6527), .B(n4265), .ZN(n6531) );
  AND2_X1 U8151 ( .A1(n9021), .A2(n6528), .ZN(n6529) );
  AOI21_X1 U8152 ( .B1(n9191), .B2(n4244), .A(n6529), .ZN(n6530) );
  NAND2_X1 U8153 ( .A1(n6531), .A2(n6530), .ZN(n8026) );
  OAI21_X1 U8154 ( .B1(n6531), .B2(n6530), .A(n8026), .ZN(n6532) );
  NOR2_X1 U8155 ( .A1(n6532), .A2(n4281), .ZN(n6533) );
  NAND2_X1 U8156 ( .A1(n6339), .A2(n6843), .ZN(n9759) );
  AND2_X1 U8157 ( .A1(n9759), .A2(n6589), .ZN(n6540) );
  OR2_X1 U8158 ( .A1(n6534), .A2(n6784), .ZN(n6541) );
  NOR2_X1 U8159 ( .A1(n6541), .A2(n7960), .ZN(n6537) );
  NAND2_X1 U8160 ( .A1(n6540), .A2(n6537), .ZN(n8853) );
  NAND2_X1 U8161 ( .A1(n6537), .A2(n6546), .ZN(n6535) );
  NOR2_X1 U8162 ( .A1(n8998), .A2(n8837), .ZN(n6536) );
  AND2_X1 U8163 ( .A1(n6537), .A2(n6838), .ZN(n6539) );
  INV_X1 U8164 ( .A(n6539), .ZN(n6538) );
  INV_X1 U8165 ( .A(n7959), .ZN(n9589) );
  AOI22_X1 U8166 ( .A1(n8856), .A2(n8831), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n6551) );
  INV_X1 U8167 ( .A(n6540), .ZN(n6544) );
  INV_X1 U8168 ( .A(n6541), .ZN(n6690) );
  AND3_X1 U8169 ( .A1(n6542), .A2(n6590), .A3(n7452), .ZN(n6543) );
  OAI21_X1 U8170 ( .B1(n6544), .B2(n6690), .A(n6543), .ZN(n6545) );
  NAND2_X1 U8171 ( .A1(n6545), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6549) );
  INV_X1 U8172 ( .A(n6838), .ZN(n7961) );
  INV_X1 U8173 ( .A(n6546), .ZN(n6929) );
  NAND2_X1 U8174 ( .A1(n7961), .A2(n6929), .ZN(n6547) );
  NAND2_X1 U8175 ( .A1(n6547), .A2(n9402), .ZN(n6691) );
  OR2_X1 U8176 ( .A1(n6691), .A2(n6690), .ZN(n6548) );
  NAND2_X1 U8177 ( .A1(n6549), .A2(n6548), .ZN(n8844) );
  NAND2_X1 U8178 ( .A1(n8996), .A2(n8844), .ZN(n6550) );
  OAI211_X1 U8179 ( .C1(n9001), .C2(n8807), .A(n6551), .B(n6550), .ZN(n6552)
         );
  INV_X1 U8180 ( .A(n7452), .ZN(n6553) );
  OR2_X1 U8181 ( .A1(n6590), .A2(n6553), .ZN(n6593) );
  NOR2_X1 U8182 ( .A1(n6593), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X1 U8183 ( .A(n9864), .ZN(n9858) );
  NOR2_X2 U8184 ( .A1(n6706), .A2(n9858), .ZN(P2_U3966) );
  INV_X1 U8185 ( .A(n6554), .ZN(n7557) );
  AOI211_X1 U8186 ( .C1(n6556), .C2(n6555), .A(n8216), .B(n7557), .ZN(n6561)
         );
  NOR2_X1 U8187 ( .A1(n4598), .A2(n8190), .ZN(n6560) );
  INV_X1 U8188 ( .A(n7608), .ZN(n6557) );
  OAI22_X1 U8189 ( .A1(n8198), .A2(n6557), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7282), .ZN(n6559) );
  OAI22_X1 U8190 ( .A1(n7601), .A2(n8199), .B1(n8200), .B2(n7600), .ZN(n6558)
         );
  OR4_X1 U8191 ( .A1(n6561), .A2(n6560), .A3(n6559), .A4(n6558), .ZN(P2_U3236)
         );
  NOR2_X2 U8192 ( .A1(n6567), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9416) );
  AOI22_X1 U8193 ( .A1(n9416), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n9592), .ZN(n6562) );
  OAI21_X1 U8194 ( .B1(n6575), .B2(n6758), .A(n6562), .ZN(P1_U3351) );
  INV_X1 U8195 ( .A(n9416), .ZN(n7086) );
  INV_X1 U8196 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6563) );
  OAI222_X1 U8197 ( .A1(n7086), .A2(n6563), .B1(n6758), .B2(n6568), .C1(
        P1_U3084), .C2(n4502), .ZN(P1_U3352) );
  INV_X1 U8198 ( .A(n6642), .ZN(n9428) );
  OAI222_X1 U8199 ( .A1(n7086), .A2(n6564), .B1(n6758), .B2(n6570), .C1(
        P1_U3084), .C2(n9428), .ZN(P1_U3350) );
  AOI22_X1 U8200 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9600), .B1(n9416), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6565) );
  OAI21_X1 U8201 ( .B1(n6572), .B2(n6758), .A(n6565), .ZN(P1_U3349) );
  AOI22_X1 U8202 ( .A1(n6657), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9416), .ZN(n6566) );
  OAI21_X1 U8203 ( .B1(n6578), .B2(n6758), .A(n6566), .ZN(P1_U3348) );
  NOR2_X1 U8204 ( .A1(n6567), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8715) );
  OAI222_X1 U8205 ( .A1(n8722), .A2(n6569), .B1(n8719), .B2(n6568), .C1(
        P2_U3152), .C2(n6727), .ZN(P2_U3357) );
  INV_X1 U8206 ( .A(n6723), .ZN(n6749) );
  OAI222_X1 U8207 ( .A1(n8722), .A2(n6571), .B1(n8719), .B2(n6570), .C1(
        P2_U3152), .C2(n6749), .ZN(P2_U3355) );
  OAI222_X1 U8208 ( .A1(n8722), .A2(n6573), .B1(n8719), .B2(n6572), .C1(
        P2_U3152), .C2(n6911), .ZN(P2_U3354) );
  OAI222_X1 U8209 ( .A1(n8722), .A2(n6576), .B1(n8719), .B2(n6575), .C1(
        P2_U3152), .C2(n6574), .ZN(P2_U3356) );
  OAI222_X1 U8210 ( .A1(n8722), .A2(n6579), .B1(n8719), .B2(n6578), .C1(
        P2_U3152), .C2(n6577), .ZN(P2_U3353) );
  INV_X1 U8211 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6582) );
  INV_X1 U8212 ( .A(n6777), .ZN(n6580) );
  NAND2_X1 U8213 ( .A1(n6580), .A2(n9402), .ZN(n6581) );
  OAI21_X1 U8214 ( .B1(n9402), .B2(n6582), .A(n6581), .ZN(P1_U3441) );
  INV_X1 U8215 ( .A(n6583), .ZN(n6585) );
  INV_X1 U8216 ( .A(n8722), .ZN(n7450) );
  AOI22_X1 U8217 ( .A1(n8258), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n7450), .ZN(n6584) );
  OAI21_X1 U8218 ( .B1(n6585), .B2(n8719), .A(n6584), .ZN(P2_U3352) );
  INV_X1 U8219 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9383) );
  OAI222_X1 U8220 ( .A1(n7086), .A2(n9383), .B1(n6758), .B2(n6585), .C1(
        P1_U3084), .C2(n6644), .ZN(P1_U3347) );
  INV_X1 U8221 ( .A(n4361), .ZN(n6588) );
  AOI22_X1 U8222 ( .A1(n8271), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n7450), .ZN(n6586) );
  OAI21_X1 U8223 ( .B1(n6588), .B2(n8719), .A(n6586), .ZN(P2_U3351) );
  AOI22_X1 U8224 ( .A1(n6996), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9416), .ZN(n6587) );
  OAI21_X1 U8225 ( .B1(n6588), .B2(n6758), .A(n6587), .ZN(P1_U3346) );
  NAND2_X1 U8226 ( .A1(n6590), .A2(n6589), .ZN(n6591) );
  NAND2_X1 U8227 ( .A1(n6591), .A2(n7452), .ZN(n6595) );
  NAND2_X1 U8228 ( .A1(n4967), .A2(n6595), .ZN(n6592) );
  NAND2_X1 U8229 ( .A1(n6592), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U8230 ( .A(P1_U3083), .ZN(n6594) );
  NAND2_X1 U8231 ( .A1(n6594), .A2(n6593), .ZN(n9667) );
  INV_X1 U8232 ( .A(n9667), .ZN(n8933) );
  NAND2_X1 U8233 ( .A1(n6628), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U8234 ( .A1(n6595), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6634) );
  INV_X1 U8235 ( .A(n6634), .ZN(n6601) );
  INV_X1 U8236 ( .A(n9584), .ZN(n7649) );
  NOR2_X1 U8237 ( .A1(n7959), .A2(n7649), .ZN(n6596) );
  NAND2_X1 U8238 ( .A1(n6601), .A2(n6596), .ZN(n9575) );
  OR2_X1 U8239 ( .A1(n9584), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6598) );
  AOI21_X1 U8240 ( .B1(n9589), .B2(n6598), .A(P1_IR_REG_0__SCAN_IN), .ZN(n9588) );
  INV_X1 U8241 ( .A(n9588), .ZN(n6602) );
  NAND2_X1 U8242 ( .A1(n9584), .A2(n6628), .ZN(n6597) );
  AND2_X1 U8243 ( .A1(n4967), .A2(n6597), .ZN(n6600) );
  NAND3_X1 U8244 ( .A1(n9589), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6598), .ZN(
        n6599) );
  NAND4_X1 U8245 ( .A1(n6602), .A2(n6601), .A3(n6600), .A4(n6599), .ZN(n6604)
         );
  NAND2_X1 U8246 ( .A1(P1_U3084), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6603) );
  OAI211_X1 U8247 ( .C1(n6605), .C2(n9575), .A(n6604), .B(n6603), .ZN(n6606)
         );
  AOI21_X1 U8248 ( .B1(n8933), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n6606), .ZN(
        n6607) );
  INV_X1 U8249 ( .A(n6607), .ZN(P1_U3241) );
  INV_X1 U8250 ( .A(n6608), .ZN(n6610) );
  INV_X1 U8251 ( .A(n8880), .ZN(n6995) );
  OAI222_X1 U8252 ( .A1(n7086), .A2(n6609), .B1(n6758), .B2(n6610), .C1(
        P1_U3084), .C2(n6995), .ZN(P1_U3345) );
  INV_X1 U8253 ( .A(n8284), .ZN(n6916) );
  OAI222_X1 U8254 ( .A1(n8722), .A2(n6611), .B1(n8719), .B2(n6610), .C1(
        P2_U3152), .C2(n6916), .ZN(P2_U3350) );
  INV_X1 U8255 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6613) );
  NAND2_X1 U8256 ( .A1(n6829), .A2(P2_U3966), .ZN(n6612) );
  OAI21_X1 U8257 ( .B1(P2_U3966), .B2(n6613), .A(n6612), .ZN(P2_U3552) );
  INV_X1 U8258 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6615) );
  NAND2_X1 U8259 ( .A1(n8383), .A2(P2_U3966), .ZN(n6614) );
  OAI21_X1 U8260 ( .B1(P2_U3966), .B2(n6615), .A(n6614), .ZN(P2_U3583) );
  INV_X1 U8261 ( .A(n6616), .ZN(n6619) );
  AOI22_X1 U8262 ( .A1(n8297), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n7450), .ZN(n6617) );
  OAI21_X1 U8263 ( .B1(n6619), .B2(n8719), .A(n6617), .ZN(P2_U3349) );
  AOI22_X1 U8264 ( .A1(n9620), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9416), .ZN(n6618) );
  OAI21_X1 U8265 ( .B1(n6619), .B2(n6758), .A(n6618), .ZN(P1_U3344) );
  NAND2_X1 U8266 ( .A1(n9851), .A2(n6620), .ZN(n6621) );
  NAND2_X1 U8267 ( .A1(n6621), .A2(n6710), .ZN(n6623) );
  OR2_X1 U8268 ( .A1(n9851), .A2(n6325), .ZN(n6622) );
  NAND2_X1 U8269 ( .A1(n6623), .A2(n6622), .ZN(n9437) );
  INV_X1 U8270 ( .A(n9437), .ZN(n9793) );
  NOR2_X1 U8271 ( .A1(n9793), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X2 U8272 ( .A(P2_U3966), .ZN(n8238) );
  NAND2_X1 U8273 ( .A1(n8238), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n6624) );
  OAI21_X1 U8274 ( .B1(n8137), .B2(n8238), .A(n6624), .ZN(P2_U3568) );
  INV_X1 U8275 ( .A(n6644), .ZN(n6671) );
  INV_X1 U8276 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9776) );
  AOI22_X1 U8277 ( .A1(n6671), .A2(P1_REG1_REG_6__SCAN_IN), .B1(n9776), .B2(
        n6644), .ZN(n6633) );
  NAND2_X1 U8278 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6657), .ZN(n6625) );
  OAI21_X1 U8279 ( .B1(n6657), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6625), .ZN(
        n6653) );
  NOR2_X1 U8280 ( .A1(P1_REG1_REG_4__SCAN_IN), .A2(n9600), .ZN(n6626) );
  AOI21_X1 U8281 ( .B1(n9600), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6626), .ZN(
        n9603) );
  NAND2_X1 U8282 ( .A1(n6639), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6627) );
  OAI21_X1 U8283 ( .B1(n6639), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6627), .ZN(
        n9567) );
  NOR3_X1 U8284 ( .A1(n6629), .A2(n6628), .A3(n9567), .ZN(n9566) );
  AOI21_X1 U8285 ( .B1(n6639), .B2(P1_REG1_REG_1__SCAN_IN), .A(n9566), .ZN(
        n9578) );
  NAND2_X1 U8286 ( .A1(P1_REG1_REG_2__SCAN_IN), .A2(n9592), .ZN(n6630) );
  OAI21_X1 U8287 ( .B1(n9592), .B2(P1_REG1_REG_2__SCAN_IN), .A(n6630), .ZN(
        n9577) );
  NOR2_X1 U8288 ( .A1(n9578), .A2(n9577), .ZN(n9576) );
  AOI21_X1 U8289 ( .B1(n9592), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9576), .ZN(
        n9422) );
  NAND2_X1 U8290 ( .A1(n6642), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U8291 ( .B1(n6642), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6631), .ZN(
        n9421) );
  NOR2_X1 U8292 ( .A1(n9422), .A2(n9421), .ZN(n9420) );
  NAND2_X1 U8293 ( .A1(n9603), .A2(n9602), .ZN(n9601) );
  OAI21_X1 U8294 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9600), .A(n9601), .ZN(
        n6654) );
  NOR2_X1 U8295 ( .A1(n6653), .A2(n6654), .ZN(n6652) );
  NAND2_X1 U8296 ( .A1(n6633), .A2(n6632), .ZN(n6668) );
  OAI21_X1 U8297 ( .B1(n6633), .B2(n6632), .A(n6668), .ZN(n6650) );
  INV_X1 U8298 ( .A(n9575), .ZN(n9661) );
  INV_X1 U8299 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6637) );
  OR2_X1 U8300 ( .A1(n6634), .A2(n9584), .ZN(n8948) );
  OR2_X1 U8301 ( .A1(n8948), .A2(n9589), .ZN(n9634) );
  INV_X1 U8302 ( .A(n9634), .ZN(n9654) );
  NAND2_X1 U8303 ( .A1(n9654), .A2(n6671), .ZN(n6636) );
  AND2_X1 U8304 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8818) );
  INV_X1 U8305 ( .A(n8818), .ZN(n6635) );
  OAI211_X1 U8306 ( .C1(n9667), .C2(n6637), .A(n6636), .B(n6635), .ZN(n6649)
         );
  NOR2_X1 U8307 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6657), .ZN(n6638) );
  AOI21_X1 U8308 ( .B1(n6657), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6638), .ZN(
        n6660) );
  NAND2_X1 U8309 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9583) );
  NOR2_X1 U8310 ( .A1(n9583), .A2(n9570), .ZN(n9569) );
  AOI21_X1 U8311 ( .B1(n6639), .B2(P1_REG2_REG_1__SCAN_IN), .A(n9569), .ZN(
        n9582) );
  NAND2_X1 U8312 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n9592), .ZN(n6640) );
  OAI21_X1 U8313 ( .B1(n9592), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6640), .ZN(
        n9581) );
  NAND2_X1 U8314 ( .A1(n6642), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6641) );
  OAI21_X1 U8315 ( .B1(n6642), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6641), .ZN(
        n9424) );
  NOR2_X1 U8316 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(n9600), .ZN(n6643) );
  AOI21_X1 U8317 ( .B1(n9600), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6643), .ZN(
        n9597) );
  NAND2_X1 U8318 ( .A1(n9598), .A2(n9597), .ZN(n9596) );
  OAI21_X1 U8319 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9600), .A(n9596), .ZN(
        n6659) );
  NAND2_X1 U8320 ( .A1(n6660), .A2(n6659), .ZN(n6658) );
  OAI21_X1 U8321 ( .B1(n6657), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6658), .ZN(
        n6647) );
  MUX2_X1 U8322 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6645), .S(n6644), .Z(n6646)
         );
  NOR2_X1 U8323 ( .A1(n6647), .A2(n6646), .ZN(n6670) );
  OR2_X1 U8324 ( .A1(n8948), .A2(n7959), .ZN(n9626) );
  AOI211_X1 U8325 ( .C1(n6647), .C2(n6646), .A(n6670), .B(n9626), .ZN(n6648)
         );
  AOI211_X1 U8326 ( .C1(n6650), .C2(n9661), .A(n6649), .B(n6648), .ZN(n6651)
         );
  INV_X1 U8327 ( .A(n6651), .ZN(P1_U3247) );
  NAND2_X1 U8328 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7012) );
  INV_X1 U8329 ( .A(n7012), .ZN(n6656) );
  AOI211_X1 U8330 ( .C1(n6654), .C2(n6653), .A(n6652), .B(n9575), .ZN(n6655)
         );
  AOI211_X1 U8331 ( .C1(n9654), .C2(n6657), .A(n6656), .B(n6655), .ZN(n6663)
         );
  INV_X1 U8332 ( .A(n9626), .ZN(n9662) );
  OAI21_X1 U8333 ( .B1(n6660), .B2(n6659), .A(n6658), .ZN(n6661) );
  AOI22_X1 U8334 ( .A1(n8933), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9662), .B2(
        n6661), .ZN(n6662) );
  NAND2_X1 U8335 ( .A1(n6663), .A2(n6662), .ZN(P1_U3246) );
  INV_X1 U8336 ( .A(n6664), .ZN(n6677) );
  INV_X1 U8337 ( .A(n7001), .ZN(n9633) );
  OAI222_X1 U8338 ( .A1(n6758), .A2(n6677), .B1(n9633), .B2(P1_U3084), .C1(
        n6665), .C2(n7086), .ZN(P1_U3343) );
  INV_X1 U8339 ( .A(n6666), .ZN(n6679) );
  AOI22_X1 U8340 ( .A1(n7141), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n7450), .ZN(n6667) );
  OAI21_X1 U8341 ( .B1(n6679), .B2(n8719), .A(n6667), .ZN(P2_U3347) );
  XNOR2_X1 U8342 ( .A(n6996), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6986) );
  XNOR2_X1 U8343 ( .A(n6985), .B(n6986), .ZN(n6675) );
  NAND2_X1 U8344 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7089) );
  INV_X1 U8345 ( .A(n7089), .ZN(n6669) );
  AOI21_X1 U8346 ( .B1(n8933), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6669), .ZN(
        n6674) );
  XNOR2_X1 U8347 ( .A(n6996), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6998) );
  XNOR2_X1 U8348 ( .A(n6998), .B(n6997), .ZN(n6672) );
  AOI22_X1 U8349 ( .A1(n6996), .A2(n9654), .B1(n9662), .B2(n6672), .ZN(n6673)
         );
  OAI211_X1 U8350 ( .C1(n6675), .C2(n9575), .A(n6674), .B(n6673), .ZN(P1_U3248) );
  INV_X1 U8351 ( .A(n6974), .ZN(n6924) );
  OAI222_X1 U8352 ( .A1(P2_U3152), .A2(n6924), .B1(n8719), .B2(n6677), .C1(
        n6676), .C2(n8722), .ZN(P2_U3348) );
  INV_X1 U8353 ( .A(n9640), .ZN(n6984) );
  INV_X1 U8354 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6678) );
  OAI222_X1 U8355 ( .A1(n6758), .A2(n6679), .B1(n6984), .B2(P1_U3084), .C1(
        n6678), .C2(n7086), .ZN(P1_U3342) );
  INV_X1 U8356 ( .A(n6680), .ZN(n6682) );
  INV_X1 U8357 ( .A(n7279), .ZN(n7152) );
  OAI222_X1 U8358 ( .A1(n8722), .A2(n6681), .B1(n8719), .B2(n6682), .C1(
        P2_U3152), .C2(n7152), .ZN(P2_U3346) );
  INV_X1 U8359 ( .A(n7524), .ZN(n7517) );
  OAI222_X1 U8360 ( .A1(n7086), .A2(n6683), .B1(n6758), .B2(n6682), .C1(
        P1_U3084), .C2(n7517), .ZN(P1_U3341) );
  INV_X1 U8361 ( .A(n6684), .ZN(n6702) );
  AOI22_X1 U8362 ( .A1(n8887), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9416), .ZN(n6685) );
  OAI21_X1 U8363 ( .B1(n6702), .B2(n6758), .A(n6685), .ZN(P1_U3340) );
  INV_X1 U8364 ( .A(n6687), .ZN(n6688) );
  AOI21_X1 U8365 ( .B1(n6689), .B2(n6686), .A(n6688), .ZN(n9585) );
  AOI21_X1 U8366 ( .B1(n6691), .B2(n9244), .A(n6690), .ZN(n6692) );
  OR2_X1 U8367 ( .A1(n6692), .A2(n6785), .ZN(n6752) );
  AOI22_X1 U8368 ( .A1(P1_REG3_REG_0__SCAN_IN), .A2(n6752), .B1(n8850), .B2(
        n7080), .ZN(n6694) );
  NAND2_X1 U8369 ( .A1(n8843), .A2(n6335), .ZN(n6693) );
  OAI211_X1 U8370 ( .C1(n9585), .C2(n8853), .A(n6694), .B(n6693), .ZN(P1_U3230) );
  XNOR2_X1 U8371 ( .A(n6695), .B(n6696), .ZN(n6698) );
  XNOR2_X1 U8372 ( .A(n6698), .B(n6697), .ZN(n6701) );
  AOI22_X1 U8373 ( .A1(P1_REG3_REG_1__SCAN_IN), .A2(n6752), .B1(n8850), .B2(
        n6851), .ZN(n6700) );
  AOI22_X1 U8374 ( .A1(n8843), .A2(n6363), .B1(n8831), .B2(n6346), .ZN(n6699)
         );
  OAI211_X1 U8375 ( .C1(n6701), .C2(n8853), .A(n6700), .B(n6699), .ZN(P1_U3220) );
  INV_X1 U8376 ( .A(n7383), .ZN(n7377) );
  OAI222_X1 U8377 ( .A1(n8722), .A2(n6703), .B1(n8719), .B2(n6702), .C1(n7377), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  NAND2_X1 U8378 ( .A1(n9851), .A2(n6704), .ZN(n6709) );
  OAI21_X1 U8379 ( .B1(n6706), .B2(P2_U3152), .A(n6705), .ZN(n6707) );
  INV_X1 U8380 ( .A(n6707), .ZN(n6708) );
  NAND2_X1 U8381 ( .A1(n6709), .A2(n6708), .ZN(n6711) );
  NAND2_X1 U8382 ( .A1(n6711), .A2(n6710), .ZN(n6718) );
  NAND2_X1 U8383 ( .A1(n6718), .A2(n8238), .ZN(n6734) );
  AND2_X1 U8384 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8159) );
  INV_X1 U8385 ( .A(n6727), .ZN(n9440) );
  NAND2_X1 U8386 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9434) );
  INV_X1 U8387 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6712) );
  NAND2_X1 U8388 ( .A1(n6727), .A2(n6712), .ZN(n6714) );
  NAND2_X1 U8389 ( .A1(n9440), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8390 ( .A1(n6714), .A2(n6713), .ZN(n9435) );
  NOR2_X1 U8391 ( .A1(n9434), .A2(n9435), .ZN(n9433) );
  AOI21_X1 U8392 ( .B1(n9440), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9433), .ZN(
        n9451) );
  NAND2_X1 U8393 ( .A1(n9453), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6715) );
  OAI21_X1 U8394 ( .B1(n9453), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6715), .ZN(
        n9450) );
  NAND2_X1 U8395 ( .A1(n6723), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6716) );
  OAI21_X1 U8396 ( .B1(n6723), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6716), .ZN(
        n6740) );
  NAND2_X1 U8397 ( .A1(n6889), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6717) );
  OAI21_X1 U8398 ( .B1(n6889), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6717), .ZN(
        n6720) );
  NOR2_X1 U8399 ( .A1(n6721), .A2(n6720), .ZN(n6888) );
  INV_X1 U8400 ( .A(n6718), .ZN(n6719) );
  INV_X1 U8401 ( .A(n9787), .ZN(n9448) );
  AOI211_X1 U8402 ( .C1(n6721), .C2(n6720), .A(n6888), .B(n9448), .ZN(n6722)
         );
  AOI211_X1 U8403 ( .C1(n9793), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n8159), .B(
        n6722), .ZN(n6738) );
  NAND2_X1 U8404 ( .A1(n6723), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6731) );
  INV_X1 U8405 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6724) );
  MUX2_X1 U8406 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6724), .S(n6723), .Z(n6745)
         );
  NAND2_X1 U8407 ( .A1(n9453), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6730) );
  INV_X1 U8408 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6725) );
  MUX2_X1 U8409 ( .A(n6725), .B(P2_REG2_REG_2__SCAN_IN), .S(n9453), .Z(n6726)
         );
  INV_X1 U8410 ( .A(n6726), .ZN(n9456) );
  NAND2_X1 U8411 ( .A1(n9440), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6729) );
  INV_X1 U8412 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6728) );
  MUX2_X1 U8413 ( .A(n6728), .B(P2_REG2_REG_1__SCAN_IN), .S(n6727), .Z(n9444)
         );
  NAND3_X1 U8414 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9444), .ZN(n9443) );
  NAND2_X1 U8415 ( .A1(n6729), .A2(n9443), .ZN(n9457) );
  NAND2_X1 U8416 ( .A1(n9456), .A2(n9457), .ZN(n9455) );
  NAND2_X1 U8417 ( .A1(n6730), .A2(n9455), .ZN(n6746) );
  NAND2_X1 U8418 ( .A1(n6745), .A2(n6746), .ZN(n6744) );
  NAND2_X1 U8419 ( .A1(n6731), .A2(n6744), .ZN(n6736) );
  INV_X1 U8420 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6732) );
  MUX2_X1 U8421 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6732), .S(n6889), .Z(n6735)
         );
  INV_X1 U8422 ( .A(n8004), .ZN(n6733) );
  NAND2_X1 U8423 ( .A1(n6734), .A2(n6733), .ZN(n9790) );
  OR2_X1 U8424 ( .A1(n9790), .A2(n6092), .ZN(n8373) );
  NAND2_X1 U8425 ( .A1(n6735), .A2(n6736), .ZN(n6910) );
  OAI211_X1 U8426 ( .C1(n6736), .C2(n6735), .A(n9784), .B(n6910), .ZN(n6737)
         );
  OAI211_X1 U8427 ( .C1(n9789), .C2(n6911), .A(n6738), .B(n6737), .ZN(P2_U3249) );
  AND2_X1 U8428 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6743) );
  AOI211_X1 U8429 ( .C1(n6741), .C2(n6740), .A(n6739), .B(n9448), .ZN(n6742)
         );
  AOI211_X1 U8430 ( .C1(n9793), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6743), .B(
        n6742), .ZN(n6748) );
  OAI211_X1 U8431 ( .C1(n6746), .C2(n6745), .A(n9784), .B(n6744), .ZN(n6747)
         );
  OAI211_X1 U8432 ( .C1(n9789), .C2(n6749), .A(n6748), .B(n6747), .ZN(P2_U3248) );
  XOR2_X1 U8433 ( .A(n6750), .B(n6751), .Z(n6755) );
  AOI22_X1 U8434 ( .A1(P1_REG3_REG_2__SCAN_IN), .A2(n6752), .B1(n8850), .B2(
        n6358), .ZN(n6754) );
  AOI22_X1 U8435 ( .A1(n8843), .A2(n8870), .B1(n8831), .B2(n6335), .ZN(n6753)
         );
  OAI211_X1 U8436 ( .C1(n6755), .C2(n8853), .A(n6754), .B(n6753), .ZN(P1_U3235) );
  INV_X1 U8437 ( .A(n6756), .ZN(n6790) );
  INV_X1 U8438 ( .A(n9653), .ZN(n7521) );
  OAI222_X1 U8439 ( .A1(n6758), .A2(n6790), .B1(n7521), .B2(P1_U3084), .C1(
        n6757), .C2(n7086), .ZN(P1_U3339) );
  INV_X1 U8440 ( .A(n8212), .ZN(n8129) );
  OR2_X1 U8441 ( .A1(n8060), .A2(n8538), .ZN(n6761) );
  NAND2_X1 U8442 ( .A1(n6829), .A2(n8571), .ZN(n6760) );
  AND2_X1 U8443 ( .A1(n6761), .A2(n6760), .ZN(n9833) );
  INV_X1 U8444 ( .A(n9833), .ZN(n6764) );
  AND2_X1 U8445 ( .A1(n6763), .A2(n7048), .ZN(n6832) );
  INV_X1 U8446 ( .A(n6832), .ZN(n6793) );
  INV_X1 U8447 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n9436) );
  AOI22_X1 U8448 ( .A1(n8129), .A2(n6764), .B1(n6793), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n6770) );
  OAI21_X1 U8449 ( .B1(n6767), .B2(n6766), .A(n6765), .ZN(n6768) );
  NAND2_X1 U8450 ( .A1(n8181), .A2(n6768), .ZN(n6769) );
  OAI211_X1 U8451 ( .C1(n6759), .C2(n8190), .A(n6770), .B(n6769), .ZN(P2_U3224) );
  INV_X1 U8452 ( .A(n6847), .ZN(n6773) );
  AND2_X1 U8453 ( .A1(n6346), .A2(n6771), .ZN(n7763) );
  OAI211_X1 U8454 ( .C1(n6773), .C2(n7763), .A(n7961), .B(n6772), .ZN(n6774)
         );
  OAI21_X1 U8455 ( .B1(n6775), .B2(n9698), .A(n6774), .ZN(n7079) );
  AOI21_X1 U8456 ( .B1(n7080), .B2(n6843), .A(n7079), .ZN(n6789) );
  OR2_X1 U8457 ( .A1(n9247), .A2(n7956), .ZN(n6780) );
  INV_X1 U8458 ( .A(n6776), .ZN(n6778) );
  AND2_X1 U8459 ( .A1(n6778), .A2(n6777), .ZN(n6779) );
  NOR2_X1 U8460 ( .A1(n6785), .A2(n6781), .ZN(n6782) );
  AND2_X2 U8461 ( .A1(n6787), .A2(n6782), .ZN(n9767) );
  NAND2_X1 U8462 ( .A1(n4495), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6783) );
  OAI21_X1 U8463 ( .B1(n6789), .B2(n4495), .A(n6783), .ZN(P1_U3454) );
  NOR2_X1 U8464 ( .A1(n6785), .A2(n6784), .ZN(n6786) );
  AND2_X2 U8465 ( .A1(n6787), .A2(n6786), .ZN(n9783) );
  NAND2_X1 U8466 ( .A1(n9780), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6788) );
  OAI21_X1 U8467 ( .B1(n6789), .B2(n9780), .A(n6788), .ZN(P1_U3523) );
  INV_X1 U8468 ( .A(n8312), .ZN(n7381) );
  OAI222_X1 U8469 ( .A1(n8722), .A2(n6791), .B1(n8719), .B2(n6790), .C1(n7381), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  OAI211_X1 U8470 ( .C1(n4342), .C2(n6792), .A(n8064), .B(n8181), .ZN(n6795)
         );
  OAI22_X1 U8471 ( .A1(n7103), .A2(n8538), .B1(n6112), .B2(n8536), .ZN(n6812)
         );
  AOI22_X1 U8472 ( .A1(n8129), .A2(n6812), .B1(n6793), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6794) );
  OAI211_X1 U8473 ( .C1(n7068), .C2(n8190), .A(n6795), .B(n6794), .ZN(P2_U3239) );
  NAND3_X1 U8474 ( .A1(n6797), .A2(n7048), .A3(n6796), .ZN(n6798) );
  INV_X1 U8475 ( .A(n7050), .ZN(n6800) );
  INV_X1 U8476 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6816) );
  NAND2_X1 U8477 ( .A1(n6801), .A2(n9835), .ZN(n9837) );
  NAND2_X1 U8478 ( .A1(n6112), .A2(n6759), .ZN(n6802) );
  NAND2_X1 U8479 ( .A1(n9837), .A2(n6802), .ZN(n6803) );
  NAND2_X1 U8480 ( .A1(n6803), .A2(n6808), .ZN(n6868) );
  OAI21_X1 U8481 ( .B1(n6803), .B2(n6808), .A(n6868), .ZN(n6804) );
  INV_X1 U8482 ( .A(n6804), .ZN(n7073) );
  XNOR2_X1 U8483 ( .A(n5580), .B(n7040), .ZN(n6805) );
  NAND2_X1 U8484 ( .A1(n6805), .A2(n8443), .ZN(n7605) );
  OR3_X1 U8485 ( .A1(n5580), .A2(n8443), .A3(n6806), .ZN(n9473) );
  NAND2_X1 U8486 ( .A1(n6759), .A2(n6833), .ZN(n9843) );
  AOI211_X1 U8487 ( .C1(n6807), .C2(n9843), .A(n9921), .B(n6874), .ZN(n7070)
         );
  AOI21_X1 U8488 ( .B1(n9927), .B2(n6807), .A(n7070), .ZN(n6814) );
  XNOR2_X1 U8489 ( .A(n6809), .B(n6808), .ZN(n6813) );
  INV_X1 U8490 ( .A(n8533), .ZN(n9830) );
  AOI21_X1 U8491 ( .B1(n6813), .B2(n9830), .A(n6812), .ZN(n7066) );
  OAI211_X1 U8492 ( .C1(n7073), .C2(n9888), .A(n6814), .B(n7066), .ZN(n6818)
         );
  NAND2_X1 U8493 ( .A1(n6818), .A2(n9937), .ZN(n6815) );
  OAI21_X1 U8494 ( .B1(n9937), .B2(n6816), .A(n6815), .ZN(P2_U3457) );
  INV_X1 U8495 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8496 ( .A1(n6818), .A2(n9952), .ZN(n6819) );
  OAI21_X1 U8497 ( .B1(n9952), .B2(n6820), .A(n6819), .ZN(P2_U3522) );
  XOR2_X1 U8498 ( .A(n6822), .B(n6821), .Z(n6826) );
  OAI22_X1 U8499 ( .A1(n9730), .A2(n8837), .B1(n8807), .B2(n9699), .ZN(n6824)
         );
  MUX2_X1 U8500 ( .A(n8844), .B(P1_U3084), .S(P1_REG3_REG_3__SCAN_IN), .Z(
        n6823) );
  AOI211_X1 U8501 ( .C1(n8831), .C2(n6363), .A(n6824), .B(n6823), .ZN(n6825)
         );
  OAI21_X1 U8502 ( .B1(n6826), .B2(n8853), .A(n6825), .ZN(P1_U3216) );
  INV_X1 U8503 ( .A(n6827), .ZN(n6837) );
  INV_X1 U8504 ( .A(n8194), .ZN(n8180) );
  AOI22_X1 U8505 ( .A1(n8180), .A2(n6829), .B1(n9865), .B2(n8181), .ZN(n6836)
         );
  INV_X1 U8506 ( .A(n8199), .ZN(n8175) );
  INV_X1 U8507 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6831) );
  OAI22_X1 U8508 ( .A1(n8190), .A2(n6833), .B1(n6832), .B2(n6831), .ZN(n6834)
         );
  AOI21_X1 U8509 ( .B1(n8175), .B2(n6830), .A(n6834), .ZN(n6835) );
  OAI21_X1 U8510 ( .B1(n6837), .B2(n6836), .A(n6835), .ZN(P2_U3234) );
  NAND2_X1 U8511 ( .A1(n6840), .A2(n6839), .ZN(n6848) );
  XNOR2_X1 U8512 ( .A(n6848), .B(n6841), .ZN(n6928) );
  NAND2_X1 U8513 ( .A1(n6851), .A2(n7080), .ZN(n6844) );
  AND2_X1 U8514 ( .A1(n6843), .A2(n6842), .ZN(n9526) );
  NAND2_X1 U8515 ( .A1(n6844), .A2(n9526), .ZN(n6845) );
  NOR2_X1 U8516 ( .A1(n7222), .A2(n6845), .ZN(n6937) );
  INV_X1 U8517 ( .A(n7722), .ZN(n6846) );
  NOR2_X1 U8518 ( .A1(n7725), .A2(n6846), .ZN(n7768) );
  OAI21_X1 U8519 ( .B1(n6848), .B2(n6847), .A(n9701), .ZN(n6850) );
  AOI22_X1 U8520 ( .A1(n9152), .A2(n6363), .B1(n6346), .B2(n9154), .ZN(n6849)
         );
  OAI21_X1 U8521 ( .B1(n7768), .B2(n6850), .A(n6849), .ZN(n6933) );
  AOI211_X1 U8522 ( .C1(n9244), .C2(n6851), .A(n6937), .B(n6933), .ZN(n6852)
         );
  OAI21_X1 U8523 ( .B1(n9529), .B2(n6928), .A(n6852), .ZN(n6854) );
  NAND2_X1 U8524 ( .A1(n6854), .A2(n9767), .ZN(n6853) );
  OAI21_X1 U8525 ( .B1(n9767), .B2(n4888), .A(n6853), .ZN(P1_U3457) );
  INV_X1 U8526 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6856) );
  NAND2_X1 U8527 ( .A1(n6854), .A2(n9783), .ZN(n6855) );
  OAI21_X1 U8528 ( .B1(n9783), .B2(n6856), .A(n6855), .ZN(P1_U3524) );
  NAND2_X1 U8529 ( .A1(n6857), .A2(n6858), .ZN(n6859) );
  XOR2_X1 U8530 ( .A(n6860), .B(n6859), .Z(n6866) );
  AOI22_X1 U8531 ( .A1(n8843), .A2(n8868), .B1(n8831), .B2(n8870), .ZN(n6865)
         );
  INV_X1 U8532 ( .A(n7207), .ZN(n6863) );
  INV_X1 U8533 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6861) );
  OAI22_X1 U8534 ( .A1(n8837), .A2(n9735), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6861), .ZN(n6862) );
  AOI21_X1 U8535 ( .B1(n6863), .B2(n8844), .A(n6862), .ZN(n6864) );
  OAI211_X1 U8536 ( .C1(n6866), .C2(n8853), .A(n6865), .B(n6864), .ZN(P1_U3228) );
  INV_X1 U8537 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8538 ( .A1(n8060), .A2(n7068), .ZN(n6867) );
  NAND2_X1 U8539 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  OAI21_X1 U8540 ( .B1(n6869), .B2(n6870), .A(n7019), .ZN(n9823) );
  INV_X1 U8541 ( .A(n9823), .ZN(n6877) );
  INV_X1 U8542 ( .A(n7605), .ZN(n7364) );
  XNOR2_X1 U8543 ( .A(n6871), .B(n6870), .ZN(n6872) );
  INV_X1 U8544 ( .A(n8538), .ZN(n8572) );
  AOI22_X1 U8545 ( .A1(n8571), .A2(n8237), .B1(n8235), .B2(n8572), .ZN(n8068)
         );
  OAI21_X1 U8546 ( .B1(n6872), .B2(n8533), .A(n8068), .ZN(n6873) );
  AOI21_X1 U8547 ( .B1(n7364), .B2(n9823), .A(n6873), .ZN(n9826) );
  INV_X1 U8548 ( .A(n6874), .ZN(n6875) );
  NAND2_X1 U8549 ( .A1(n6874), .A2(n9818), .ZN(n7029) );
  INV_X1 U8550 ( .A(n7029), .ZN(n7097) );
  AOI211_X1 U8551 ( .C1(n6115), .C2(n6875), .A(n9921), .B(n7097), .ZN(n9816)
         );
  AOI21_X1 U8552 ( .B1(n9927), .B2(n6115), .A(n9816), .ZN(n6876) );
  OAI211_X1 U8553 ( .C1(n6877), .C2(n9473), .A(n9826), .B(n6876), .ZN(n6880)
         );
  NAND2_X1 U8554 ( .A1(n6880), .A2(n9937), .ZN(n6878) );
  OAI21_X1 U8555 ( .B1(n9937), .B2(n6879), .A(n6878), .ZN(P2_U3460) );
  INV_X1 U8556 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U8557 ( .A1(n6880), .A2(n9952), .ZN(n6881) );
  OAI21_X1 U8558 ( .B1(n9952), .B2(n6882), .A(n6881), .ZN(P2_U3523) );
  INV_X1 U8559 ( .A(n6883), .ZN(n6885) );
  OAI222_X1 U8560 ( .A1(n7086), .A2(n6884), .B1(n6758), .B2(n6885), .C1(
        P1_U3084), .C2(n8905), .ZN(P1_U3338) );
  INV_X1 U8561 ( .A(n8326), .ZN(n8319) );
  OAI222_X1 U8562 ( .A1(n8722), .A2(n6886), .B1(n8719), .B2(n6885), .C1(
        P2_U3152), .C2(n8319), .ZN(P2_U3343) );
  NAND2_X1 U8563 ( .A1(n8238), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n6887) );
  OAI21_X1 U8564 ( .B1(n8111), .B2(n8238), .A(n6887), .ZN(P2_U3578) );
  AND2_X1 U8565 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7247) );
  OR2_X1 U8566 ( .A1(n8244), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8567 ( .A1(n8244), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U8568 ( .A1(n6891), .A2(n6890), .ZN(n8247) );
  OR2_X1 U8569 ( .A1(n8258), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6893) );
  NAND2_X1 U8570 ( .A1(n8258), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8571 ( .A1(n6893), .A2(n6892), .ZN(n8261) );
  AOI21_X1 U8572 ( .B1(n8258), .B2(P2_REG1_REG_6__SCAN_IN), .A(n8259), .ZN(
        n8273) );
  OR2_X1 U8573 ( .A1(n8271), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6895) );
  NAND2_X1 U8574 ( .A1(n8271), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6894) );
  NAND2_X1 U8575 ( .A1(n6895), .A2(n6894), .ZN(n8274) );
  NOR2_X1 U8576 ( .A1(n8273), .A2(n8274), .ZN(n8272) );
  AOI21_X1 U8577 ( .B1(n8271), .B2(P2_REG1_REG_7__SCAN_IN), .A(n8272), .ZN(
        n8287) );
  INV_X1 U8578 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6896) );
  MUX2_X1 U8579 ( .A(n6896), .B(P2_REG1_REG_8__SCAN_IN), .S(n8284), .Z(n8286)
         );
  INV_X1 U8580 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6897) );
  MUX2_X1 U8581 ( .A(n6897), .B(P2_REG1_REG_9__SCAN_IN), .S(n8297), .Z(n8300)
         );
  INV_X1 U8582 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6898) );
  MUX2_X1 U8583 ( .A(n6898), .B(P2_REG1_REG_10__SCAN_IN), .S(n6974), .Z(n6899)
         );
  NOR2_X1 U8584 ( .A1(n6900), .A2(n6899), .ZN(n6973) );
  AOI211_X1 U8585 ( .C1(n6900), .C2(n6899), .A(n6973), .B(n9448), .ZN(n6901)
         );
  AOI211_X1 U8586 ( .C1(n9793), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7247), .B(
        n6901), .ZN(n6923) );
  NAND2_X1 U8587 ( .A1(n8297), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6917) );
  INV_X1 U8588 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6902) );
  MUX2_X1 U8589 ( .A(n6902), .B(P2_REG2_REG_9__SCAN_IN), .S(n8297), .Z(n6903)
         );
  INV_X1 U8590 ( .A(n6903), .ZN(n8294) );
  INV_X1 U8591 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6915) );
  MUX2_X1 U8592 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6915), .S(n8284), .Z(n8281)
         );
  NAND2_X1 U8593 ( .A1(n8271), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6914) );
  INV_X1 U8594 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6904) );
  MUX2_X1 U8595 ( .A(n6904), .B(P2_REG2_REG_7__SCAN_IN), .S(n8271), .Z(n6905)
         );
  INV_X1 U8596 ( .A(n6905), .ZN(n8268) );
  NAND2_X1 U8597 ( .A1(n8258), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6913) );
  INV_X1 U8598 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6906) );
  MUX2_X1 U8599 ( .A(n6906), .B(P2_REG2_REG_6__SCAN_IN), .S(n8258), .Z(n6907)
         );
  INV_X1 U8600 ( .A(n6907), .ZN(n8254) );
  NAND2_X1 U8601 ( .A1(n8244), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6912) );
  INV_X1 U8602 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6908) );
  MUX2_X1 U8603 ( .A(n6908), .B(P2_REG2_REG_5__SCAN_IN), .S(n8244), .Z(n6909)
         );
  INV_X1 U8604 ( .A(n6909), .ZN(n8240) );
  OAI21_X1 U8605 ( .B1(n6911), .B2(n6732), .A(n6910), .ZN(n8241) );
  NAND2_X1 U8606 ( .A1(n8240), .A2(n8241), .ZN(n8239) );
  NAND2_X1 U8607 ( .A1(n6912), .A2(n8239), .ZN(n8255) );
  NAND2_X1 U8608 ( .A1(n8254), .A2(n8255), .ZN(n8253) );
  NAND2_X1 U8609 ( .A1(n6913), .A2(n8253), .ZN(n8269) );
  NAND2_X1 U8610 ( .A1(n8268), .A2(n8269), .ZN(n8267) );
  NAND2_X1 U8611 ( .A1(n6914), .A2(n8267), .ZN(n8282) );
  NAND2_X1 U8612 ( .A1(n8281), .A2(n8282), .ZN(n8280) );
  OAI21_X1 U8613 ( .B1(n6916), .B2(n6915), .A(n8280), .ZN(n8295) );
  NAND2_X1 U8614 ( .A1(n8294), .A2(n8295), .ZN(n8293) );
  NAND2_X1 U8615 ( .A1(n6917), .A2(n8293), .ZN(n6921) );
  INV_X1 U8616 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6918) );
  MUX2_X1 U8617 ( .A(n6918), .B(P2_REG2_REG_10__SCAN_IN), .S(n6974), .Z(n6919)
         );
  INV_X1 U8618 ( .A(n6919), .ZN(n6920) );
  NAND2_X1 U8619 ( .A1(n6920), .A2(n6921), .ZN(n6966) );
  OAI211_X1 U8620 ( .C1(n6921), .C2(n6920), .A(n9784), .B(n6966), .ZN(n6922)
         );
  OAI211_X1 U8621 ( .C1(n9789), .C2(n6924), .A(n6923), .B(n6922), .ZN(P2_U3255) );
  INV_X1 U8622 ( .A(n8335), .ZN(n8341) );
  INV_X1 U8623 ( .A(n6925), .ZN(n6940) );
  OAI222_X1 U8624 ( .A1(P2_U3152), .A2(n8341), .B1(n8719), .B2(n6940), .C1(
        n6926), .C2(n8722), .ZN(P2_U3342) );
  OR2_X1 U8625 ( .A1(n5254), .A2(n6927), .ZN(n7221) );
  AOI21_X1 U8626 ( .B1(n9704), .B2(n7221), .A(n6928), .ZN(n6934) );
  INV_X1 U8627 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6931) );
  OAI22_X1 U8628 ( .A1(n9105), .A2(n6931), .B1(n6930), .B2(n6929), .ZN(n6932)
         );
  NOR3_X1 U8629 ( .A1(n6934), .A2(n6933), .A3(n6932), .ZN(n6939) );
  INV_X1 U8630 ( .A(n6935), .ZN(n6936) );
  NAND2_X1 U8631 ( .A1(n6936), .A2(n5254), .ZN(n7660) );
  INV_X1 U8632 ( .A(n7660), .ZN(n9170) );
  AOI22_X1 U8633 ( .A1(n9170), .A2(n6937), .B1(n9517), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6938) );
  OAI21_X1 U8634 ( .B1(n6939), .B2(n9708), .A(n6938), .ZN(P1_U3290) );
  INV_X1 U8635 ( .A(n8921), .ZN(n8913) );
  OAI222_X1 U8636 ( .A1(n7086), .A2(n6941), .B1(n8913), .B2(P1_U3084), .C1(
        n6758), .C2(n6940), .ZN(P1_U3337) );
  OAI21_X1 U8637 ( .B1(n6943), .B2(n6953), .A(n6942), .ZN(n6951) );
  INV_X1 U8638 ( .A(n6943), .ZN(n6945) );
  NAND3_X1 U8639 ( .A1(n8180), .A2(n6945), .A3(n6944), .ZN(n6946) );
  AOI21_X1 U8640 ( .B1(n6946), .B2(n8200), .A(n8157), .ZN(n6950) );
  INV_X1 U8641 ( .A(n6947), .ZN(n7053) );
  AOI22_X1 U8642 ( .A1(n9883), .A2(n8214), .B1(n8175), .B2(n8232), .ZN(n6948)
         );
  NAND2_X1 U8643 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8256) );
  OAI211_X1 U8644 ( .C1(n7053), .C2(n8198), .A(n6948), .B(n8256), .ZN(n6949)
         );
  AOI211_X1 U8645 ( .C1(n6951), .C2(n8181), .A(n6950), .B(n6949), .ZN(n6952)
         );
  INV_X1 U8646 ( .A(n6952), .ZN(P2_U3241) );
  INV_X1 U8647 ( .A(n6953), .ZN(n6954) );
  AOI211_X1 U8648 ( .C1(n6956), .C2(n6955), .A(n8216), .B(n6954), .ZN(n6960)
         );
  AOI22_X1 U8649 ( .A1(n7031), .A2(n8214), .B1(n8175), .B2(n8233), .ZN(n6958)
         );
  AOI22_X1 U8650 ( .A1(n8209), .A2(n7058), .B1(P2_REG3_REG_5__SCAN_IN), .B2(
        P2_U3152), .ZN(n6957) );
  OAI211_X1 U8651 ( .C1(n7020), .C2(n8200), .A(n6958), .B(n6957), .ZN(n6959)
         );
  OR2_X1 U8652 ( .A1(n6960), .A2(n6959), .ZN(P2_U3229) );
  NAND2_X1 U8653 ( .A1(n8238), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6961) );
  OAI21_X1 U8654 ( .B1(n8405), .B2(n8238), .A(n6961), .ZN(P2_U3581) );
  INV_X1 U8655 ( .A(n8357), .ZN(n8348) );
  INV_X1 U8656 ( .A(n6962), .ZN(n6964) );
  OAI222_X1 U8657 ( .A1(P2_U3152), .A2(n8348), .B1(n8719), .B2(n6964), .C1(
        n6963), .C2(n8722), .ZN(P2_U3341) );
  INV_X1 U8658 ( .A(n8939), .ZN(n6965) );
  OAI222_X1 U8659 ( .A1(n7086), .A2(n9359), .B1(n6965), .B2(P1_U3084), .C1(
        n6758), .C2(n6964), .ZN(P1_U3336) );
  NAND2_X1 U8660 ( .A1(n6974), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6967) );
  NAND2_X1 U8661 ( .A1(n6967), .A2(n6966), .ZN(n6971) );
  INV_X1 U8662 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6968) );
  MUX2_X1 U8663 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n6968), .S(n7141), .Z(n6969)
         );
  INV_X1 U8664 ( .A(n6969), .ZN(n6970) );
  NOR2_X1 U8665 ( .A1(n6971), .A2(n6970), .ZN(n7135) );
  AOI21_X1 U8666 ( .B1(n6971), .B2(n6970), .A(n7135), .ZN(n6983) );
  INV_X1 U8667 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6972) );
  MUX2_X1 U8668 ( .A(n6972), .B(P2_REG1_REG_11__SCAN_IN), .S(n7141), .Z(n6976)
         );
  AOI21_X1 U8669 ( .B1(n6976), .B2(n6975), .A(n7140), .ZN(n6980) );
  INV_X1 U8670 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n6978) );
  NOR2_X1 U8671 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5769), .ZN(n7345) );
  INV_X1 U8672 ( .A(n7345), .ZN(n6977) );
  OAI21_X1 U8673 ( .B1(n9437), .B2(n6978), .A(n6977), .ZN(n6979) );
  AOI21_X1 U8674 ( .B1(n9787), .B2(n6980), .A(n6979), .ZN(n6982) );
  NAND2_X1 U8675 ( .A1(n9454), .A2(n7141), .ZN(n6981) );
  OAI211_X1 U8676 ( .C1(n6983), .C2(n8373), .A(n6982), .B(n6981), .ZN(P2_U3256) );
  INV_X1 U8677 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9557) );
  AOI22_X1 U8678 ( .A1(n9640), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n9557), .B2(
        n6984), .ZN(n9643) );
  INV_X1 U8679 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7421) );
  AOI22_X1 U8680 ( .A1(n7001), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n7421), .B2(
        n9633), .ZN(n9625) );
  INV_X1 U8681 ( .A(n6985), .ZN(n6987) );
  INV_X1 U8682 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6988) );
  MUX2_X1 U8683 ( .A(n6988), .B(P1_REG1_REG_8__SCAN_IN), .S(n8880), .Z(n8873)
         );
  NOR2_X1 U8684 ( .A1(n8872), .A2(n8873), .ZN(n8871) );
  NOR2_X1 U8685 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9620), .ZN(n6989) );
  AOI21_X1 U8686 ( .B1(n9620), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6989), .ZN(
        n9611) );
  NAND2_X1 U8687 ( .A1(n9612), .A2(n9611), .ZN(n9610) );
  OAI21_X1 U8688 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9620), .A(n9610), .ZN(
        n9624) );
  NAND2_X1 U8689 ( .A1(n9625), .A2(n9624), .ZN(n9623) );
  OAI21_X1 U8690 ( .B1(n7001), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9623), .ZN(
        n9642) );
  NAND2_X1 U8691 ( .A1(n9643), .A2(n9642), .ZN(n9641) );
  OAI21_X1 U8692 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n9640), .A(n9641), .ZN(
        n6992) );
  INV_X1 U8693 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6990) );
  MUX2_X1 U8694 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6990), .S(n7524), .Z(n6991)
         );
  NAND2_X1 U8695 ( .A1(n6991), .A2(n6992), .ZN(n7523) );
  OAI21_X1 U8696 ( .B1(n6992), .B2(n6991), .A(n7523), .ZN(n7007) );
  NAND2_X1 U8697 ( .A1(n8933), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U8698 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7549) );
  OAI211_X1 U8699 ( .C1(n9634), .C2(n7517), .A(n6993), .B(n7549), .ZN(n7006)
         );
  NOR2_X1 U8700 ( .A1(n9640), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6994) );
  AOI21_X1 U8701 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9640), .A(n6994), .ZN(
        n9646) );
  AOI22_X1 U8702 ( .A1(n8880), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n5023), .B2(
        n6995), .ZN(n8877) );
  OAI21_X1 U8703 ( .B1(n8880), .B2(P1_REG2_REG_8__SCAN_IN), .A(n8876), .ZN(
        n9618) );
  MUX2_X1 U8704 ( .A(n6999), .B(P1_REG2_REG_9__SCAN_IN), .S(n9620), .Z(n9617)
         );
  NOR2_X1 U8705 ( .A1(n9618), .A2(n9617), .ZN(n9616) );
  NAND2_X1 U8706 ( .A1(n7001), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7000) );
  OAI21_X1 U8707 ( .B1(n7001), .B2(P1_REG2_REG_10__SCAN_IN), .A(n7000), .ZN(
        n9628) );
  OAI21_X1 U8708 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9640), .A(n9644), .ZN(
        n7004) );
  NAND2_X1 U8709 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n7524), .ZN(n7002) );
  OAI21_X1 U8710 ( .B1(n7524), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7002), .ZN(
        n7003) );
  NOR2_X1 U8711 ( .A1(n7003), .A2(n7004), .ZN(n7514) );
  AOI211_X1 U8712 ( .C1(n7004), .C2(n7003), .A(n7514), .B(n9626), .ZN(n7005)
         );
  AOI211_X1 U8713 ( .C1(n9661), .C2(n7007), .A(n7006), .B(n7005), .ZN(n7008)
         );
  INV_X1 U8714 ( .A(n7008), .ZN(P1_U3253) );
  OAI21_X1 U8715 ( .B1(n7011), .B2(n7009), .A(n7010), .ZN(n7016) );
  INV_X1 U8716 ( .A(n8831), .ZN(n8848) );
  OAI22_X1 U8717 ( .A1(n8848), .A2(n9699), .B1(n7185), .B2(n8807), .ZN(n7015)
         );
  NAND2_X1 U8718 ( .A1(n8844), .A2(n7187), .ZN(n7013) );
  OAI211_X1 U8719 ( .C1(n9745), .C2(n8837), .A(n7013), .B(n7012), .ZN(n7014)
         );
  AOI211_X1 U8720 ( .C1(n7016), .C2(n8829), .A(n7015), .B(n7014), .ZN(n7017)
         );
  INV_X1 U8721 ( .A(n7017), .ZN(P1_U3225) );
  INV_X1 U8722 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7034) );
  NAND2_X1 U8723 ( .A1(n7103), .A2(n9818), .ZN(n7018) );
  NAND2_X1 U8724 ( .A1(n7019), .A2(n7018), .ZN(n7095) );
  NAND2_X1 U8725 ( .A1(n7095), .A2(n7100), .ZN(n7094) );
  NAND2_X1 U8726 ( .A1(n7020), .A2(n9877), .ZN(n7021) );
  NAND2_X1 U8727 ( .A1(n7022), .A2(n7026), .ZN(n7043) );
  OAI21_X1 U8728 ( .B1(n7022), .B2(n7026), .A(n7043), .ZN(n7023) );
  INV_X1 U8729 ( .A(n7023), .ZN(n7065) );
  NAND2_X1 U8730 ( .A1(n7025), .A2(n7024), .ZN(n7027) );
  XNOR2_X1 U8731 ( .A(n7027), .B(n7026), .ZN(n7028) );
  AOI222_X1 U8732 ( .A1(n9830), .A2(n7028), .B1(n8233), .B2(n8572), .C1(n8235), 
        .C2(n8571), .ZN(n7057) );
  OR2_X1 U8733 ( .A1(n7029), .A2(n7098), .ZN(n7096) );
  OR2_X1 U8734 ( .A1(n7096), .A2(n7031), .ZN(n7047) );
  AOI21_X1 U8735 ( .B1(n7096), .B2(n7031), .A(n9921), .ZN(n7030) );
  AND2_X1 U8736 ( .A1(n7047), .A2(n7030), .ZN(n7062) );
  AOI21_X1 U8737 ( .B1(n9927), .B2(n7031), .A(n7062), .ZN(n7032) );
  OAI211_X1 U8738 ( .C1(n9888), .C2(n7065), .A(n7057), .B(n7032), .ZN(n7035)
         );
  NAND2_X1 U8739 ( .A1(n7035), .A2(n9952), .ZN(n7033) );
  OAI21_X1 U8740 ( .B1(n9952), .B2(n7034), .A(n7033), .ZN(P2_U3525) );
  INV_X1 U8741 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U8742 ( .A1(n7035), .A2(n9937), .ZN(n7036) );
  OAI21_X1 U8743 ( .B1(n9937), .B2(n7037), .A(n7036), .ZN(P2_U3466) );
  INV_X1 U8744 ( .A(n7038), .ZN(n7049) );
  NAND3_X1 U8745 ( .A1(n7050), .A2(n7048), .A3(n7049), .ZN(n7039) );
  INV_X2 U8746 ( .A(n9815), .ZN(n8495) );
  OR2_X1 U8747 ( .A1(n7040), .A2(n8443), .ZN(n7176) );
  AND2_X1 U8748 ( .A1(n7605), .A2(n7176), .ZN(n7041) );
  NAND2_X1 U8749 ( .A1(n8157), .A2(n7060), .ZN(n7042) );
  NAND2_X1 U8750 ( .A1(n7043), .A2(n7042), .ZN(n7110) );
  XNOR2_X1 U8751 ( .A(n7110), .B(n7044), .ZN(n9887) );
  XNOR2_X1 U8752 ( .A(n7045), .B(n7044), .ZN(n7046) );
  AOI222_X1 U8753 ( .A1(n9830), .A2(n7046), .B1(n8232), .B2(n8572), .C1(n8234), 
        .C2(n8571), .ZN(n9886) );
  MUX2_X1 U8754 ( .A(n6906), .B(n9886), .S(n9815), .Z(n7056) );
  AOI21_X1 U8755 ( .B1(n9883), .B2(n7047), .A(n7113), .ZN(n9884) );
  INV_X1 U8756 ( .A(n7048), .ZN(n7052) );
  NAND2_X1 U8757 ( .A1(n7050), .A2(n7049), .ZN(n7051) );
  NOR2_X1 U8758 ( .A1(n9819), .A2(n9921), .ZN(n9845) );
  OR3_X2 U8759 ( .A1(n7052), .A2(n7051), .A3(n8433), .ZN(n9817) );
  OAI22_X1 U8760 ( .A1(n9817), .A2(n7109), .B1(n9814), .B2(n7053), .ZN(n7054)
         );
  AOI21_X1 U8761 ( .B1(n9884), .B2(n9845), .A(n7054), .ZN(n7055) );
  OAI211_X1 U8762 ( .C1(n8604), .C2(n9887), .A(n7056), .B(n7055), .ZN(P2_U3290) );
  MUX2_X1 U8763 ( .A(n6908), .B(n7057), .S(n9815), .Z(n7064) );
  INV_X1 U8764 ( .A(n9819), .ZN(n9811) );
  INV_X1 U8765 ( .A(n7058), .ZN(n7059) );
  OAI22_X1 U8766 ( .A1(n9817), .A2(n7060), .B1(n9814), .B2(n7059), .ZN(n7061)
         );
  AOI21_X1 U8767 ( .B1(n7062), .B2(n9811), .A(n7061), .ZN(n7063) );
  OAI211_X1 U8768 ( .C1(n7065), .C2(n8604), .A(n7064), .B(n7063), .ZN(P2_U3291) );
  MUX2_X1 U8769 ( .A(n6725), .B(n7066), .S(n9815), .Z(n7072) );
  INV_X1 U8770 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7067) );
  OAI22_X1 U8771 ( .A1(n9817), .A2(n7068), .B1(n9814), .B2(n7067), .ZN(n7069)
         );
  AOI21_X1 U8772 ( .B1(n7070), .B2(n9811), .A(n7069), .ZN(n7071) );
  OAI211_X1 U8773 ( .C1(n7073), .C2(n8604), .A(n7072), .B(n7071), .ZN(P2_U3294) );
  INV_X1 U8774 ( .A(n9867), .ZN(n7078) );
  AOI22_X1 U8775 ( .A1(n9867), .A2(n9830), .B1(n8572), .B2(n6830), .ZN(n9869)
         );
  OAI21_X1 U8776 ( .B1(n6831), .B2(n9814), .A(n9869), .ZN(n7075) );
  INV_X1 U8777 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n9785) );
  NOR2_X1 U8778 ( .A1(n9815), .A2(n9785), .ZN(n7074) );
  AOI21_X1 U8779 ( .B1(n9815), .B2(n7075), .A(n7074), .ZN(n7077) );
  INV_X1 U8780 ( .A(n9817), .ZN(n9841) );
  OAI21_X1 U8781 ( .B1(n9845), .B2(n9841), .A(n9865), .ZN(n7076) );
  OAI211_X1 U8782 ( .C1(n7078), .C2(n8604), .A(n7077), .B(n7076), .ZN(P2_U3296) );
  AOI21_X1 U8783 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n9707), .A(n7079), .ZN(
        n7083) );
  NAND2_X1 U8784 ( .A1(n9517), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7082) );
  OAI21_X1 U8785 ( .B1(n9107), .B2(n9692), .A(n7080), .ZN(n7081) );
  OAI211_X1 U8786 ( .C1(n7083), .C2(n9517), .A(n7082), .B(n7081), .ZN(P1_U3291) );
  INV_X1 U8787 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9315) );
  INV_X1 U8788 ( .A(n7084), .ZN(n7085) );
  OAI222_X1 U8789 ( .A1(n8722), .A2(n9315), .B1(n8719), .B2(n7085), .C1(
        P2_U3152), .C2(n8360), .ZN(P2_U3340) );
  INV_X1 U8790 ( .A(n8950), .ZN(n8936) );
  OAI222_X1 U8791 ( .A1(n7086), .A2(n9380), .B1(n6758), .B2(n7085), .C1(
        P1_U3084), .C2(n8936), .ZN(P1_U3335) );
  XOR2_X1 U8792 ( .A(n7088), .B(n7087), .Z(n7093) );
  AOI22_X1 U8793 ( .A1(n7124), .A2(n8844), .B1(n8843), .B2(n8865), .ZN(n7090)
         );
  OAI211_X1 U8794 ( .C1(n7185), .C2(n8848), .A(n7090), .B(n7089), .ZN(n7091)
         );
  AOI21_X1 U8795 ( .B1(n7130), .B2(n8850), .A(n7091), .ZN(n7092) );
  OAI21_X1 U8796 ( .B1(n7093), .B2(n8853), .A(n7092), .ZN(P1_U3211) );
  INV_X1 U8797 ( .A(n8604), .ZN(n9838) );
  OAI21_X1 U8798 ( .B1(n7095), .B2(n7100), .A(n7094), .ZN(n9881) );
  INV_X1 U8799 ( .A(n9845), .ZN(n8387) );
  OAI21_X1 U8800 ( .B1(n7097), .B2(n9877), .A(n7096), .ZN(n9878) );
  AOI22_X1 U8801 ( .A1(n9841), .A2(n7098), .B1(n9839), .B2(n8160), .ZN(n7099)
         );
  OAI21_X1 U8802 ( .B1(n8387), .B2(n9878), .A(n7099), .ZN(n7105) );
  XNOR2_X1 U8803 ( .A(n7101), .B(n7100), .ZN(n7102) );
  OAI222_X1 U8804 ( .A1(n8538), .A2(n8157), .B1(n8536), .B2(n7103), .C1(n7102), 
        .C2(n8533), .ZN(n9879) );
  MUX2_X1 U8805 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n9879), .S(n9815), .Z(n7104)
         );
  AOI211_X1 U8806 ( .C1(n9838), .C2(n9881), .A(n7105), .B(n7104), .ZN(n7106)
         );
  INV_X1 U8807 ( .A(n7106), .ZN(P2_U3292) );
  INV_X1 U8808 ( .A(n7107), .ZN(n7165) );
  AOI22_X1 U8809 ( .A1(n7953), .A2(P1_STATE_REG_SCAN_IN), .B1(n9416), .B2(
        P2_DATAO_REG_19__SCAN_IN), .ZN(n7108) );
  OAI21_X1 U8810 ( .B1(n7165), .B2(n6758), .A(n7108), .ZN(P1_U3334) );
  OAI21_X1 U8811 ( .B1(n7110), .B2(n7109), .A(n7118), .ZN(n7112) );
  NAND2_X1 U8812 ( .A1(n7110), .A2(n7109), .ZN(n7111) );
  NAND2_X1 U8813 ( .A1(n7112), .A2(n7111), .ZN(n7168) );
  XNOR2_X1 U8814 ( .A(n7168), .B(n7167), .ZN(n9895) );
  OAI211_X1 U8815 ( .C1(n7113), .C2(n9893), .A(n7177), .B(n4341), .ZN(n9891)
         );
  AOI22_X1 U8816 ( .A1(n9841), .A2(n8039), .B1(n9839), .B2(n8038), .ZN(n7114)
         );
  OAI21_X1 U8817 ( .B1(n9891), .B2(n9819), .A(n7114), .ZN(n7115) );
  AOI21_X1 U8818 ( .B1(n9895), .B2(n9838), .A(n7115), .ZN(n7121) );
  XNOR2_X1 U8819 ( .A(n7116), .B(n7117), .ZN(n7119) );
  OAI22_X1 U8820 ( .A1(n7262), .A2(n8538), .B1(n7118), .B2(n8536), .ZN(n8037)
         );
  AOI21_X1 U8821 ( .B1(n7119), .B2(n9830), .A(n8037), .ZN(n9892) );
  MUX2_X1 U8822 ( .A(n9892), .B(n6904), .S(n8495), .Z(n7120) );
  NAND2_X1 U8823 ( .A1(n7121), .A2(n7120), .ZN(P2_U3289) );
  XNOR2_X1 U8824 ( .A(n7122), .B(n4674), .ZN(n7123) );
  AOI222_X1 U8825 ( .A1(n9701), .A2(n7123), .B1(n8867), .B2(n9154), .C1(n8865), 
        .C2(n9152), .ZN(n9754) );
  INV_X1 U8826 ( .A(n7124), .ZN(n7125) );
  OAI22_X1 U8827 ( .A1(n9684), .A2(n7126), .B1(n7125), .B2(n9105), .ZN(n7129)
         );
  INV_X1 U8828 ( .A(n9526), .ZN(n9761) );
  AOI21_X1 U8829 ( .B1(n7325), .B2(n7130), .A(n9761), .ZN(n7127) );
  NAND2_X1 U8830 ( .A1(n7127), .A2(n7154), .ZN(n9753) );
  NOR2_X1 U8831 ( .A1(n9753), .A2(n7660), .ZN(n7128) );
  AOI211_X1 U8832 ( .C1(n9107), .C2(n7130), .A(n7129), .B(n7128), .ZN(n7134)
         );
  XNOR2_X1 U8833 ( .A(n7132), .B(n7131), .ZN(n9757) );
  INV_X1 U8834 ( .A(n9176), .ZN(n7307) );
  NAND2_X1 U8835 ( .A1(n9757), .A2(n7307), .ZN(n7133) );
  OAI211_X1 U8836 ( .C1(n9754), .C2(n9708), .A(n7134), .B(n7133), .ZN(P1_U3284) );
  NOR2_X1 U8837 ( .A1(n7141), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7136) );
  NOR2_X1 U8838 ( .A1(n7136), .A2(n7135), .ZN(n7139) );
  INV_X1 U8839 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7137) );
  MUX2_X1 U8840 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7137), .S(n7279), .Z(n7138)
         );
  NAND2_X1 U8841 ( .A1(n7279), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7275) );
  OAI211_X1 U8842 ( .C1(n7279), .C2(P2_REG2_REG_12__SCAN_IN), .A(n7139), .B(
        n7275), .ZN(n7274) );
  OAI211_X1 U8843 ( .C1(n7139), .C2(n7138), .A(n7274), .B(n9784), .ZN(n7151)
         );
  INV_X1 U8844 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7142) );
  MUX2_X1 U8845 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n7142), .S(n7279), .Z(n7143)
         );
  OAI21_X1 U8846 ( .B1(n7144), .B2(n7143), .A(n7278), .ZN(n7149) );
  NOR2_X1 U8847 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7145), .ZN(n7148) );
  INV_X1 U8848 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7146) );
  NOR2_X1 U8849 ( .A1(n9437), .A2(n7146), .ZN(n7147) );
  AOI211_X1 U8850 ( .C1(n9787), .C2(n7149), .A(n7148), .B(n7147), .ZN(n7150)
         );
  OAI211_X1 U8851 ( .C1(n9789), .C2(n7152), .A(n7151), .B(n7150), .ZN(P2_U3257) );
  XNOR2_X1 U8852 ( .A(n7841), .B(n7839), .ZN(n7153) );
  AOI222_X1 U8853 ( .A1(n9701), .A2(n7153), .B1(n8866), .B2(n9154), .C1(n8864), 
        .C2(n9152), .ZN(n7315) );
  AOI211_X1 U8854 ( .C1(n7313), .C2(n7154), .A(n9761), .B(n9669), .ZN(n7312)
         );
  NOR2_X1 U8855 ( .A1(n9710), .A2(n7155), .ZN(n7158) );
  INV_X1 U8856 ( .A(n7156), .ZN(n7293) );
  OAI22_X1 U8857 ( .A1(n9684), .A2(n5023), .B1(n7293), .B2(n9105), .ZN(n7157)
         );
  AOI211_X1 U8858 ( .C1(n7312), .C2(n9170), .A(n7158), .B(n7157), .ZN(n7164)
         );
  NAND2_X1 U8859 ( .A1(n7160), .A2(n7839), .ZN(n7161) );
  NAND2_X1 U8860 ( .A1(n7159), .A2(n7161), .ZN(n7316) );
  INV_X1 U8861 ( .A(n7316), .ZN(n7162) );
  NAND2_X1 U8862 ( .A1(n7162), .A2(n7307), .ZN(n7163) );
  OAI211_X1 U8863 ( .C1(n7315), .C2(n9708), .A(n7164), .B(n7163), .ZN(P1_U3283) );
  OAI222_X1 U8864 ( .A1(n8722), .A2(n7166), .B1(n8719), .B2(n7165), .C1(
        P2_U3152), .C2(n8443), .ZN(P2_U3339) );
  NAND2_X1 U8865 ( .A1(n9893), .A2(n8088), .ZN(n7169) );
  XNOR2_X1 U8866 ( .A(n7250), .B(n7252), .ZN(n9899) );
  NAND2_X1 U8867 ( .A1(n9899), .A2(n7364), .ZN(n7175) );
  OAI21_X1 U8868 ( .B1(n7251), .B2(n7171), .A(n7170), .ZN(n7173) );
  OAI22_X1 U8869 ( .A1(n7359), .A2(n8538), .B1(n8088), .B2(n8536), .ZN(n7172)
         );
  AOI21_X1 U8870 ( .B1(n7173), .B2(n9830), .A(n7172), .ZN(n7174) );
  AND2_X1 U8871 ( .A1(n7175), .A2(n7174), .ZN(n9901) );
  NOR2_X1 U8872 ( .A1(n9840), .A2(n7176), .ZN(n9824) );
  NAND2_X1 U8873 ( .A1(n7177), .A2(n8094), .ZN(n7178) );
  NAND2_X1 U8874 ( .A1(n7267), .A2(n7178), .ZN(n9897) );
  NOR2_X1 U8875 ( .A1(n9897), .A2(n8387), .ZN(n7181) );
  AOI22_X1 U8876 ( .A1(n9840), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n8093), .B2(
        n9839), .ZN(n7179) );
  OAI21_X1 U8877 ( .B1(n4606), .B2(n9817), .A(n7179), .ZN(n7180) );
  AOI211_X1 U8878 ( .C1(n9899), .C2(n9824), .A(n7181), .B(n7180), .ZN(n7182)
         );
  OAI21_X1 U8879 ( .B1(n9901), .B2(n8495), .A(n7182), .ZN(P2_U3288) );
  INV_X1 U8880 ( .A(n9154), .ZN(n9696) );
  INV_X1 U8881 ( .A(n9701), .ZN(n9163) );
  XOR2_X1 U8882 ( .A(n7183), .B(n7770), .Z(n7184) );
  OAI222_X1 U8883 ( .A1(n9696), .A2(n9699), .B1(n9698), .B2(n7185), .C1(n9163), 
        .C2(n7184), .ZN(n9747) );
  INV_X1 U8884 ( .A(n9747), .ZN(n7196) );
  OAI21_X1 U8885 ( .B1(n7204), .B2(n9745), .A(n9526), .ZN(n7186) );
  OR2_X1 U8886 ( .A1(n7186), .A2(n7323), .ZN(n9743) );
  INV_X1 U8887 ( .A(n9743), .ZN(n7190) );
  AOI22_X1 U8888 ( .A1(n9708), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7187), .B2(
        n9707), .ZN(n7188) );
  OAI21_X1 U8889 ( .B1(n9745), .B2(n9710), .A(n7188), .ZN(n7189) );
  AOI21_X1 U8890 ( .B1(n7190), .B2(n9170), .A(n7189), .ZN(n7195) );
  NAND2_X1 U8891 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  NAND2_X1 U8892 ( .A1(n7193), .A2(n7770), .ZN(n9741) );
  NAND3_X1 U8893 ( .A1(n9742), .A2(n9741), .A3(n7307), .ZN(n7194) );
  OAI211_X1 U8894 ( .C1(n7196), .C2(n9517), .A(n7195), .B(n7194), .ZN(P1_U3286) );
  NAND2_X1 U8895 ( .A1(n9695), .A2(n7799), .ZN(n7198) );
  NAND2_X1 U8896 ( .A1(n7198), .A2(n7197), .ZN(n7199) );
  XNOR2_X1 U8897 ( .A(n7199), .B(n7766), .ZN(n7200) );
  NAND2_X1 U8898 ( .A1(n7200), .A2(n9701), .ZN(n7202) );
  AOI22_X1 U8899 ( .A1(n9152), .A2(n8868), .B1(n8870), .B2(n9154), .ZN(n7201)
         );
  NAND2_X1 U8900 ( .A1(n7202), .A2(n7201), .ZN(n9737) );
  INV_X1 U8901 ( .A(n9737), .ZN(n7214) );
  XNOR2_X1 U8902 ( .A(n7203), .B(n7766), .ZN(n9739) );
  INV_X1 U8903 ( .A(n9692), .ZN(n8985) );
  INV_X1 U8904 ( .A(n9689), .ZN(n7206) );
  INV_X1 U8905 ( .A(n7204), .ZN(n7205) );
  OAI21_X1 U8906 ( .B1(n9735), .B2(n7206), .A(n7205), .ZN(n9736) );
  OAI22_X1 U8907 ( .A1(n9684), .A2(n7208), .B1(n7207), .B2(n9105), .ZN(n7209)
         );
  AOI21_X1 U8908 ( .B1(n9107), .B2(n7210), .A(n7209), .ZN(n7211) );
  OAI21_X1 U8909 ( .B1(n8985), .B2(n9736), .A(n7211), .ZN(n7212) );
  AOI21_X1 U8910 ( .B1(n7307), .B2(n9739), .A(n7212), .ZN(n7213) );
  OAI21_X1 U8911 ( .B1(n7214), .B2(n9517), .A(n7213), .ZN(P1_U3287) );
  XNOR2_X1 U8912 ( .A(n7215), .B(n7764), .ZN(n7216) );
  NAND2_X1 U8913 ( .A1(n7216), .A2(n9701), .ZN(n7220) );
  XNOR2_X1 U8914 ( .A(n7217), .B(n7764), .ZN(n9727) );
  INV_X1 U8915 ( .A(n9704), .ZN(n7328) );
  NAND2_X1 U8916 ( .A1(n9727), .A2(n7328), .ZN(n7219) );
  AOI22_X1 U8917 ( .A1(n9154), .A2(n6335), .B1(n8870), .B2(n9152), .ZN(n7218)
         );
  AND3_X1 U8918 ( .A1(n7220), .A2(n7219), .A3(n7218), .ZN(n9729) );
  NOR2_X1 U8919 ( .A1(n9708), .A2(n7221), .ZN(n9693) );
  OR2_X1 U8920 ( .A1(n7222), .A2(n9724), .ZN(n7223) );
  NAND2_X1 U8921 ( .A1(n9688), .A2(n7223), .ZN(n9725) );
  AOI22_X1 U8922 ( .A1(n9708), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9707), .ZN(n7226) );
  NAND2_X1 U8923 ( .A1(n9107), .A2(n6358), .ZN(n7225) );
  OAI211_X1 U8924 ( .C1(n8985), .C2(n9725), .A(n7226), .B(n7225), .ZN(n7227)
         );
  AOI21_X1 U8925 ( .B1(n9693), .B2(n9727), .A(n7227), .ZN(n7228) );
  OAI21_X1 U8926 ( .B1(n9517), .B2(n9729), .A(n7228), .ZN(P1_U3289) );
  INV_X1 U8927 ( .A(n7229), .ZN(n7310) );
  AOI22_X1 U8928 ( .A1(n7957), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n9416), .ZN(n7230) );
  OAI21_X1 U8929 ( .B1(n7310), .B2(n6758), .A(n7230), .ZN(P1_U3333) );
  INV_X1 U8930 ( .A(n7244), .ZN(n7240) );
  INV_X1 U8931 ( .A(n7231), .ZN(n7233) );
  NAND2_X1 U8932 ( .A1(n7233), .A2(n7232), .ZN(n7235) );
  AOI22_X1 U8933 ( .A1(n7240), .A2(n7236), .B1(n7235), .B2(n7234), .ZN(n7243)
         );
  INV_X1 U8934 ( .A(n7269), .ZN(n7237) );
  OAI22_X1 U8935 ( .A1(n8198), .A2(n7237), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5735), .ZN(n7239) );
  OAI22_X1 U8936 ( .A1(n7262), .A2(n8200), .B1(n8199), .B2(n7404), .ZN(n7238)
         );
  AOI211_X1 U8937 ( .C1(n7354), .C2(n8214), .A(n7239), .B(n7238), .ZN(n7242)
         );
  INV_X1 U8938 ( .A(n7359), .ZN(n8230) );
  NAND3_X1 U8939 ( .A1(n7240), .A2(n8180), .A3(n8230), .ZN(n7241) );
  OAI211_X1 U8940 ( .C1(n7243), .C2(n8216), .A(n7242), .B(n7241), .ZN(P2_U3233) );
  INV_X1 U8941 ( .A(n7397), .ZN(n9910) );
  OAI211_X1 U8942 ( .C1(n7245), .C2(n7244), .A(n7339), .B(n8181), .ZN(n7249)
         );
  OAI22_X1 U8943 ( .A1(n7588), .A2(n8199), .B1(n8200), .B2(n7359), .ZN(n7246)
         );
  AOI211_X1 U8944 ( .C1(n7367), .C2(n8209), .A(n7247), .B(n7246), .ZN(n7248)
         );
  OAI211_X1 U8945 ( .C1(n9910), .C2(n8190), .A(n7249), .B(n7248), .ZN(P2_U3219) );
  INV_X1 U8946 ( .A(n7251), .ZN(n7252) );
  INV_X1 U8947 ( .A(n7262), .ZN(n8231) );
  NAND2_X1 U8948 ( .A1(n8094), .A2(n8231), .ZN(n7253) );
  NAND2_X1 U8949 ( .A1(n7254), .A2(n7253), .ZN(n7257) );
  INV_X1 U8950 ( .A(n7257), .ZN(n7255) );
  NAND2_X1 U8951 ( .A1(n7257), .A2(n7258), .ZN(n7259) );
  NAND2_X1 U8952 ( .A1(n7256), .A2(n7259), .ZN(n9906) );
  XNOR2_X1 U8953 ( .A(n7261), .B(n7260), .ZN(n7265) );
  OAI22_X1 U8954 ( .A1(n7262), .A2(n8536), .B1(n7404), .B2(n8538), .ZN(n7263)
         );
  INV_X1 U8955 ( .A(n7263), .ZN(n7264) );
  OAI21_X1 U8956 ( .B1(n7265), .B2(n8533), .A(n7264), .ZN(n7266) );
  AOI21_X1 U8957 ( .B1(n9906), .B2(n7364), .A(n7266), .ZN(n9908) );
  AND2_X1 U8958 ( .A1(n7267), .A2(n7354), .ZN(n7268) );
  OR2_X1 U8959 ( .A1(n7268), .A2(n7365), .ZN(n9904) );
  NOR2_X1 U8960 ( .A1(n9904), .A2(n8387), .ZN(n7272) );
  INV_X1 U8961 ( .A(n7354), .ZN(n9903) );
  AOI22_X1 U8962 ( .A1(n9840), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7269), .B2(
        n9839), .ZN(n7270) );
  OAI21_X1 U8963 ( .B1(n9903), .B2(n9817), .A(n7270), .ZN(n7271) );
  AOI211_X1 U8964 ( .C1(n9906), .C2(n9824), .A(n7272), .B(n7271), .ZN(n7273)
         );
  OAI21_X1 U8965 ( .B1(n9908), .B2(n8495), .A(n7273), .ZN(P2_U3287) );
  NAND2_X1 U8966 ( .A1(n7275), .A2(n7274), .ZN(n7277) );
  INV_X1 U8967 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7376) );
  AOI22_X1 U8968 ( .A1(n7383), .A2(n7376), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7377), .ZN(n7276) );
  NOR2_X1 U8969 ( .A1(n7277), .A2(n7276), .ZN(n7375) );
  AOI21_X1 U8970 ( .B1(n7277), .B2(n7276), .A(n7375), .ZN(n7288) );
  INV_X1 U8971 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9478) );
  AOI22_X1 U8972 ( .A1(n7383), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n9478), .B2(
        n7377), .ZN(n7281) );
  OAI21_X1 U8973 ( .B1(n7279), .B2(P2_REG1_REG_12__SCAN_IN), .A(n7278), .ZN(
        n7280) );
  NAND2_X1 U8974 ( .A1(n7281), .A2(n7280), .ZN(n7382) );
  OAI21_X1 U8975 ( .B1(n7281), .B2(n7280), .A(n7382), .ZN(n7286) );
  INV_X1 U8976 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7283) );
  OAI22_X1 U8977 ( .A1(n9437), .A2(n7283), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7282), .ZN(n7285) );
  NOR2_X1 U8978 ( .A1(n9789), .A2(n7377), .ZN(n7284) );
  AOI211_X1 U8979 ( .C1(n9787), .C2(n7286), .A(n7285), .B(n7284), .ZN(n7287)
         );
  OAI21_X1 U8980 ( .B1(n7288), .B2(n8373), .A(n7287), .ZN(P2_U3258) );
  NAND2_X1 U8981 ( .A1(n4338), .A2(n7289), .ZN(n7291) );
  XNOR2_X1 U8982 ( .A(n7291), .B(n7290), .ZN(n7297) );
  NOR2_X1 U8983 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9321), .ZN(n8875) );
  OAI22_X1 U8984 ( .A1(n8833), .A2(n7293), .B1(n8848), .B2(n7292), .ZN(n7294)
         );
  AOI211_X1 U8985 ( .C1(n8843), .C2(n8864), .A(n8875), .B(n7294), .ZN(n7296)
         );
  NAND2_X1 U8986 ( .A1(n8850), .A2(n7313), .ZN(n7295) );
  OAI211_X1 U8987 ( .C1(n7297), .C2(n8853), .A(n7296), .B(n7295), .ZN(P1_U3219) );
  XNOR2_X1 U8988 ( .A(n7298), .B(n7845), .ZN(n7299) );
  AOI222_X1 U8989 ( .A1(n9701), .A2(n7299), .B1(n8862), .B2(n9152), .C1(n8864), 
        .C2(n9154), .ZN(n7418) );
  OAI21_X1 U8990 ( .B1(n7301), .B2(n7845), .A(n7300), .ZN(n7414) );
  INV_X1 U8991 ( .A(n9671), .ZN(n7303) );
  INV_X1 U8992 ( .A(n7302), .ZN(n9507) );
  AOI211_X1 U8993 ( .C1(n7416), .C2(n7303), .A(n9761), .B(n9507), .ZN(n7415)
         );
  NAND2_X1 U8994 ( .A1(n7415), .A2(n9170), .ZN(n7305) );
  AOI22_X1 U8995 ( .A1(n9708), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7430), .B2(
        n9707), .ZN(n7304) );
  OAI211_X1 U8996 ( .C1(n7435), .C2(n9710), .A(n7305), .B(n7304), .ZN(n7306)
         );
  AOI21_X1 U8997 ( .B1(n7414), .B2(n7307), .A(n7306), .ZN(n7308) );
  OAI21_X1 U8998 ( .B1(n7418), .B2(n9517), .A(n7308), .ZN(P1_U3281) );
  OAI222_X1 U8999 ( .A1(n8722), .A2(n7311), .B1(n8719), .B2(n7310), .C1(n7309), 
        .C2(P2_U3152), .ZN(P2_U3338) );
  AOI21_X1 U9000 ( .B1(n9244), .B2(n7313), .A(n7312), .ZN(n7314) );
  OAI211_X1 U9001 ( .C1(n9529), .C2(n7316), .A(n7315), .B(n7314), .ZN(n7318)
         );
  NAND2_X1 U9002 ( .A1(n7318), .A2(n9783), .ZN(n7317) );
  OAI21_X1 U9003 ( .B1(n9783), .B2(n6988), .A(n7317), .ZN(P1_U3531) );
  NAND2_X1 U9004 ( .A1(n7318), .A2(n9767), .ZN(n7319) );
  OAI21_X1 U9005 ( .B1(n9767), .B2(n5022), .A(n7319), .ZN(P1_U3478) );
  NAND2_X1 U9006 ( .A1(n7321), .A2(n4980), .ZN(n7322) );
  NAND2_X1 U9007 ( .A1(n7320), .A2(n7322), .ZN(n9752) );
  OR2_X1 U9008 ( .A1(n7323), .A2(n9748), .ZN(n7324) );
  NAND2_X1 U9009 ( .A1(n7325), .A2(n7324), .ZN(n9749) );
  AOI22_X1 U9010 ( .A1(n9107), .A2(n8817), .B1(n9707), .B2(n8819), .ZN(n7326)
         );
  OAI21_X1 U9011 ( .B1(n9749), .B2(n8985), .A(n7326), .ZN(n7333) );
  XNOR2_X1 U9012 ( .A(n7829), .B(n4980), .ZN(n7327) );
  NAND2_X1 U9013 ( .A1(n7327), .A2(n9701), .ZN(n7331) );
  NAND2_X1 U9014 ( .A1(n9752), .A2(n7328), .ZN(n7330) );
  AOI22_X1 U9015 ( .A1(n9152), .A2(n8866), .B1(n8868), .B2(n9154), .ZN(n7329)
         );
  NAND3_X1 U9016 ( .A1(n7331), .A2(n7330), .A3(n7329), .ZN(n9750) );
  MUX2_X1 U9017 ( .A(n9750), .B(P1_REG2_REG_6__SCAN_IN), .S(n9708), .Z(n7332)
         );
  AOI211_X1 U9018 ( .C1(n9693), .C2(n9752), .A(n7333), .B(n7332), .ZN(n7334)
         );
  INV_X1 U9019 ( .A(n7334), .ZN(P1_U3285) );
  INV_X1 U9020 ( .A(n7335), .ZN(n7373) );
  AOI22_X1 U9021 ( .A1(n7956), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n9416), .ZN(n7336) );
  OAI21_X1 U9022 ( .B1(n7373), .B2(n6758), .A(n7336), .ZN(P1_U3332) );
  INV_X1 U9023 ( .A(n7589), .ZN(n9920) );
  INV_X1 U9024 ( .A(n7337), .ZN(n7338) );
  AOI21_X1 U9025 ( .B1(n7339), .B2(n7338), .A(n8216), .ZN(n7343) );
  NOR3_X1 U9026 ( .A1(n7340), .A2(n7404), .A3(n8194), .ZN(n7342) );
  OAI21_X1 U9027 ( .B1(n7343), .B2(n7342), .A(n7341), .ZN(n7347) );
  OAI22_X1 U9028 ( .A1(n7404), .A2(n8200), .B1(n8199), .B2(n7600), .ZN(n7344)
         );
  AOI211_X1 U9029 ( .C1(n8209), .C2(n7406), .A(n7345), .B(n7344), .ZN(n7346)
         );
  OAI211_X1 U9030 ( .C1(n9920), .C2(n8190), .A(n7347), .B(n7346), .ZN(P2_U3238) );
  AOI21_X1 U9031 ( .B1(n7349), .B2(n7348), .A(n4337), .ZN(n7353) );
  AOI22_X1 U9032 ( .A1(n9681), .A2(n8844), .B1(n8843), .B2(n8863), .ZN(n7350)
         );
  NAND2_X1 U9033 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9613) );
  OAI211_X1 U9034 ( .C1(n9676), .C2(n8848), .A(n7350), .B(n9613), .ZN(n7351)
         );
  AOI21_X1 U9035 ( .B1(n7705), .B2(n8850), .A(n7351), .ZN(n7352) );
  OAI21_X1 U9036 ( .B1(n7353), .B2(n8853), .A(n7352), .ZN(P1_U3229) );
  OR2_X1 U9037 ( .A1(n7354), .A2(n8230), .ZN(n7355) );
  XNOR2_X1 U9038 ( .A(n7395), .B(n7358), .ZN(n9914) );
  XNOR2_X1 U9039 ( .A(n7357), .B(n7358), .ZN(n7362) );
  OAI22_X1 U9040 ( .A1(n7588), .A2(n8538), .B1(n7359), .B2(n8536), .ZN(n7360)
         );
  INV_X1 U9041 ( .A(n7360), .ZN(n7361) );
  OAI21_X1 U9042 ( .B1(n7362), .B2(n8533), .A(n7361), .ZN(n7363) );
  AOI21_X1 U9043 ( .B1(n9914), .B2(n7364), .A(n7363), .ZN(n9916) );
  NOR2_X1 U9044 ( .A1(n7365), .A2(n9910), .ZN(n7366) );
  OR2_X1 U9045 ( .A1(n7405), .A2(n7366), .ZN(n9911) );
  NOR2_X1 U9046 ( .A1(n9911), .A2(n8387), .ZN(n7370) );
  AOI22_X1 U9047 ( .A1(n9840), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7367), .B2(
        n9839), .ZN(n7368) );
  OAI21_X1 U9048 ( .B1(n9910), .B2(n9817), .A(n7368), .ZN(n7369) );
  AOI211_X1 U9049 ( .C1(n9914), .C2(n9824), .A(n7370), .B(n7369), .ZN(n7371)
         );
  OAI21_X1 U9050 ( .B1(n9916), .B2(n8495), .A(n7371), .ZN(P2_U3286) );
  OAI222_X1 U9051 ( .A1(n8722), .A2(n7374), .B1(n8719), .B2(n7373), .C1(n7372), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  AOI21_X1 U9052 ( .B1(n7377), .B2(n7376), .A(n7375), .ZN(n7380) );
  INV_X1 U9053 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7378) );
  AOI22_X1 U9054 ( .A1(n8312), .A2(n7378), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7381), .ZN(n7379) );
  NOR2_X1 U9055 ( .A1(n7380), .A2(n7379), .ZN(n8306) );
  AOI21_X1 U9056 ( .B1(n7380), .B2(n7379), .A(n8306), .ZN(n7391) );
  INV_X1 U9057 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9472) );
  AOI22_X1 U9058 ( .A1(n8312), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9472), .B2(
        n7381), .ZN(n7385) );
  OAI21_X1 U9059 ( .B1(n7383), .B2(P2_REG1_REG_13__SCAN_IN), .A(n7382), .ZN(
        n7384) );
  OAI21_X1 U9060 ( .B1(n7385), .B2(n7384), .A(n8311), .ZN(n7389) );
  INV_X1 U9061 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7387) );
  NAND2_X1 U9062 ( .A1(n9454), .A2(n8312), .ZN(n7386) );
  NAND2_X1 U9063 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7558) );
  OAI211_X1 U9064 ( .C1(n7387), .C2(n9437), .A(n7386), .B(n7558), .ZN(n7388)
         );
  AOI21_X1 U9065 ( .B1(n7389), .B2(n9787), .A(n7388), .ZN(n7390) );
  OAI21_X1 U9066 ( .B1(n7391), .B2(n8373), .A(n7390), .ZN(P2_U3259) );
  INV_X1 U9067 ( .A(n7392), .ZN(n7412) );
  AOI22_X1 U9068 ( .A1(n7393), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n9416), .ZN(n7394) );
  OAI21_X1 U9069 ( .B1(n7412), .B2(n6758), .A(n7394), .ZN(P1_U3331) );
  INV_X1 U9070 ( .A(n7404), .ZN(n8229) );
  NAND2_X1 U9071 ( .A1(n7397), .A2(n8229), .ZN(n7398) );
  NAND2_X1 U9072 ( .A1(n7400), .A2(n7402), .ZN(n7591) );
  OAI21_X1 U9073 ( .B1(n7400), .B2(n7402), .A(n7591), .ZN(n9918) );
  XNOR2_X1 U9074 ( .A(n7401), .B(n7402), .ZN(n7403) );
  OAI222_X1 U9075 ( .A1(n8538), .A2(n7600), .B1(n8536), .B2(n7404), .C1(n7403), 
        .C2(n8533), .ZN(n9923) );
  NAND2_X1 U9076 ( .A1(n7405), .A2(n9920), .ZN(n9807) );
  OAI21_X1 U9077 ( .B1(n7405), .B2(n9920), .A(n9807), .ZN(n9922) );
  NOR2_X1 U9078 ( .A1(n9922), .A2(n8387), .ZN(n7409) );
  AOI22_X1 U9079 ( .A1(n8495), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7406), .B2(
        n9839), .ZN(n7407) );
  OAI21_X1 U9080 ( .B1(n9920), .B2(n9817), .A(n7407), .ZN(n7408) );
  AOI211_X1 U9081 ( .C1(n9923), .C2(n9815), .A(n7409), .B(n7408), .ZN(n7410)
         );
  OAI21_X1 U9082 ( .B1(n8604), .B2(n9918), .A(n7410), .ZN(P2_U3285) );
  OAI222_X1 U9083 ( .A1(n8722), .A2(n7413), .B1(n8719), .B2(n7412), .C1(
        P2_U3152), .C2(n7411), .ZN(P2_U3336) );
  INV_X1 U9084 ( .A(n7414), .ZN(n7419) );
  AOI21_X1 U9085 ( .B1(n9244), .B2(n7416), .A(n7415), .ZN(n7417) );
  OAI211_X1 U9086 ( .C1(n9529), .C2(n7419), .A(n7418), .B(n7417), .ZN(n7422)
         );
  NAND2_X1 U9087 ( .A1(n7422), .A2(n9783), .ZN(n7420) );
  OAI21_X1 U9088 ( .B1(n9783), .B2(n7421), .A(n7420), .ZN(P1_U3533) );
  NAND2_X1 U9089 ( .A1(n7422), .A2(n9767), .ZN(n7423) );
  OAI21_X1 U9090 ( .B1(n9767), .B2(n5067), .A(n7423), .ZN(P1_U3484) );
  XNOR2_X1 U9091 ( .A(n7426), .B(n7425), .ZN(n7427) );
  XNOR2_X1 U9092 ( .A(n7424), .B(n7427), .ZN(n7428) );
  NAND2_X1 U9093 ( .A1(n7428), .A2(n8829), .ZN(n7434) );
  NOR2_X1 U9094 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7429), .ZN(n9631) );
  INV_X1 U9095 ( .A(n7430), .ZN(n7431) );
  OAI22_X1 U9096 ( .A1(n8833), .A2(n7431), .B1(n7499), .B2(n8807), .ZN(n7432)
         );
  AOI211_X1 U9097 ( .C1(n8831), .C2(n8864), .A(n9631), .B(n7432), .ZN(n7433)
         );
  OAI211_X1 U9098 ( .C1(n7435), .C2(n8837), .A(n7434), .B(n7433), .ZN(P1_U3215) );
  INV_X1 U9099 ( .A(n7341), .ZN(n7438) );
  NOR3_X1 U9100 ( .A1(n7436), .A2(n7588), .A3(n8194), .ZN(n7437) );
  AOI21_X1 U9101 ( .B1(n7438), .B2(n8181), .A(n7437), .ZN(n7448) );
  INV_X1 U9102 ( .A(n9803), .ZN(n7442) );
  OR2_X1 U9103 ( .A1(n7619), .A2(n8538), .ZN(n7440) );
  OR2_X1 U9104 ( .A1(n7588), .A2(n8536), .ZN(n7439) );
  NAND2_X1 U9105 ( .A1(n7440), .A2(n7439), .ZN(n9801) );
  AOI22_X1 U9106 ( .A1(n8129), .A2(n9801), .B1(P2_REG3_REG_12__SCAN_IN), .B2(
        P2_U3152), .ZN(n7441) );
  OAI21_X1 U9107 ( .B1(n7442), .B2(n8198), .A(n7441), .ZN(n7445) );
  NOR2_X1 U9108 ( .A1(n7443), .A2(n8216), .ZN(n7444) );
  AOI211_X1 U9109 ( .C1(n9928), .C2(n8214), .A(n7445), .B(n7444), .ZN(n7446)
         );
  OAI21_X1 U9110 ( .B1(n7448), .B2(n7447), .A(n7446), .ZN(P2_U3226) );
  INV_X1 U9111 ( .A(n7449), .ZN(n7454) );
  AOI21_X1 U9112 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n7450), .A(n6325), .ZN(
        n7451) );
  OAI21_X1 U9113 ( .B1(n7454), .B2(n8719), .A(n7451), .ZN(P2_U3335) );
  NOR2_X1 U9114 ( .A1(n7452), .A2(P1_U3084), .ZN(n7965) );
  AOI21_X1 U9115 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9416), .A(n7965), .ZN(
        n7453) );
  OAI21_X1 U9116 ( .B1(n7454), .B2(n6758), .A(n7453), .ZN(P1_U3330) );
  XNOR2_X1 U9117 ( .A(n7456), .B(n7455), .ZN(n7462) );
  NOR2_X1 U9118 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5081), .ZN(n9639) );
  INV_X1 U9119 ( .A(n9516), .ZN(n7457) );
  OAI22_X1 U9120 ( .A1(n8833), .A2(n7457), .B1(n9511), .B2(n8807), .ZN(n7458)
         );
  AOI211_X1 U9121 ( .C1(n8831), .C2(n8863), .A(n9639), .B(n7458), .ZN(n7461)
         );
  NAND2_X1 U9122 ( .A1(n7459), .A2(n8850), .ZN(n7460) );
  OAI211_X1 U9123 ( .C1(n7462), .C2(n8853), .A(n7461), .B(n7460), .ZN(P1_U3234) );
  INV_X1 U9124 ( .A(n7463), .ZN(n7512) );
  AOI22_X1 U9125 ( .A1(n5474), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n9416), .ZN(n7464) );
  OAI21_X1 U9126 ( .B1(n7512), .B2(n6758), .A(n7464), .ZN(P1_U3329) );
  INV_X1 U9127 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n9988) );
  NOR2_X1 U9128 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7465) );
  AOI21_X1 U9129 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7465), .ZN(n9960) );
  NOR2_X1 U9130 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7466) );
  AOI21_X1 U9131 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7466), .ZN(n9963) );
  NOR2_X1 U9132 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7467) );
  AOI21_X1 U9133 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7467), .ZN(n9966) );
  NOR2_X1 U9134 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7468) );
  AOI21_X1 U9135 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7468), .ZN(n9969) );
  NOR2_X1 U9136 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7469) );
  AOI21_X1 U9137 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7469), .ZN(n9972) );
  NOR2_X1 U9138 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7475) );
  INV_X1 U9139 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9609) );
  XOR2_X1 U9140 ( .A(n9609), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10000) );
  NAND2_X1 U9141 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7473) );
  XOR2_X1 U9142 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n9998) );
  NAND2_X1 U9143 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7471) );
  INV_X1 U9144 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9595) );
  XNOR2_X1 U9145 ( .A(n9595), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(n9996) );
  AOI21_X1 U9146 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9953) );
  INV_X1 U9147 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9957) );
  NAND3_X1 U9148 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9955) );
  OAI21_X1 U9149 ( .B1(n9953), .B2(n9957), .A(n9955), .ZN(n9995) );
  NAND2_X1 U9150 ( .A1(n9996), .A2(n9995), .ZN(n7470) );
  NAND2_X1 U9151 ( .A1(n7471), .A2(n7470), .ZN(n9997) );
  NAND2_X1 U9152 ( .A1(n9998), .A2(n9997), .ZN(n7472) );
  NAND2_X1 U9153 ( .A1(n7473), .A2(n7472), .ZN(n9999) );
  NOR2_X1 U9154 ( .A1(n10000), .A2(n9999), .ZN(n7474) );
  NOR2_X1 U9155 ( .A1(n7475), .A2(n7474), .ZN(n7476) );
  NOR2_X1 U9156 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7476), .ZN(n9984) );
  AND2_X1 U9157 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7476), .ZN(n9983) );
  NOR2_X1 U9158 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9983), .ZN(n7477) );
  NOR2_X1 U9159 ( .A1(n9984), .A2(n7477), .ZN(n7478) );
  NAND2_X1 U9160 ( .A1(n7478), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7480) );
  XOR2_X1 U9161 ( .A(n7478), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n9982) );
  NAND2_X1 U9162 ( .A1(n9982), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U9163 ( .A1(n7480), .A2(n7479), .ZN(n7481) );
  NAND2_X1 U9164 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7481), .ZN(n7483) );
  XOR2_X1 U9165 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7481), .Z(n9994) );
  NAND2_X1 U9166 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n9994), .ZN(n7482) );
  NAND2_X1 U9167 ( .A1(n7483), .A2(n7482), .ZN(n7484) );
  NAND2_X1 U9168 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7484), .ZN(n7486) );
  XOR2_X1 U9169 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7484), .Z(n9993) );
  NAND2_X1 U9170 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n9993), .ZN(n7485) );
  NAND2_X1 U9171 ( .A1(n7486), .A2(n7485), .ZN(n7487) );
  AND2_X1 U9172 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7487), .ZN(n7488) );
  INV_X1 U9173 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n9992) );
  XNOR2_X1 U9174 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7487), .ZN(n9991) );
  NOR2_X1 U9175 ( .A1(n9992), .A2(n9991), .ZN(n9990) );
  NAND2_X1 U9176 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7489) );
  OAI21_X1 U9177 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7489), .ZN(n9980) );
  AOI21_X1 U9178 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9979), .ZN(n9978) );
  NAND2_X1 U9179 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7490) );
  OAI21_X1 U9180 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7490), .ZN(n9977) );
  NOR2_X1 U9181 ( .A1(n9978), .A2(n9977), .ZN(n9976) );
  AOI21_X1 U9182 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9976), .ZN(n9975) );
  NOR2_X1 U9183 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7491) );
  AOI21_X1 U9184 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7491), .ZN(n9974) );
  NAND2_X1 U9185 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  OAI21_X1 U9186 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9973), .ZN(n9971) );
  NAND2_X1 U9187 ( .A1(n9972), .A2(n9971), .ZN(n9970) );
  OAI21_X1 U9188 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9970), .ZN(n9968) );
  NAND2_X1 U9189 ( .A1(n9969), .A2(n9968), .ZN(n9967) );
  OAI21_X1 U9190 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9967), .ZN(n9965) );
  NAND2_X1 U9191 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  OAI21_X1 U9192 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9964), .ZN(n9962) );
  NAND2_X1 U9193 ( .A1(n9963), .A2(n9962), .ZN(n9961) );
  OAI21_X1 U9194 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9961), .ZN(n9959) );
  NAND2_X1 U9195 ( .A1(n9960), .A2(n9959), .ZN(n9958) );
  OAI21_X1 U9196 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9958), .ZN(n9987) );
  NOR2_X1 U9197 ( .A1(n9988), .A2(n9987), .ZN(n7492) );
  NAND2_X1 U9198 ( .A1(n9988), .A2(n9987), .ZN(n9986) );
  OAI21_X1 U9199 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7492), .A(n9986), .ZN(
        n7494) );
  XNOR2_X1 U9200 ( .A(n8959), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7493) );
  XNOR2_X1 U9201 ( .A(n7494), .B(n7493), .ZN(ADD_1071_U4) );
  NAND2_X1 U9202 ( .A1(n7495), .A2(n7774), .ZN(n7496) );
  NAND2_X1 U9203 ( .A1(n7497), .A2(n7496), .ZN(n9546) );
  INV_X1 U9204 ( .A(n9693), .ZN(n7510) );
  XOR2_X1 U9205 ( .A(n7774), .B(n7498), .Z(n7501) );
  OAI22_X1 U9206 ( .A1(n7708), .A2(n9698), .B1(n7499), .B2(n9696), .ZN(n7500)
         );
  AOI21_X1 U9207 ( .B1(n7501), .B2(n9701), .A(n7500), .ZN(n7502) );
  OAI21_X1 U9208 ( .B1(n9704), .B2(n9546), .A(n7502), .ZN(n9549) );
  NAND2_X1 U9209 ( .A1(n9549), .A2(n9684), .ZN(n7509) );
  INV_X1 U9210 ( .A(n7503), .ZN(n7550) );
  OAI22_X1 U9211 ( .A1(n9684), .A2(n7516), .B1(n7550), .B2(n9105), .ZN(n7506)
         );
  INV_X1 U9212 ( .A(n9506), .ZN(n7504) );
  OAI211_X1 U9213 ( .C1(n7504), .C2(n9548), .A(n9526), .B(n9487), .ZN(n9547)
         );
  NOR2_X1 U9214 ( .A1(n9547), .A2(n7660), .ZN(n7505) );
  AOI211_X1 U9215 ( .C1(n9107), .C2(n7507), .A(n7506), .B(n7505), .ZN(n7508)
         );
  OAI211_X1 U9216 ( .C1(n9546), .C2(n7510), .A(n7509), .B(n7508), .ZN(P1_U3279) );
  OAI222_X1 U9217 ( .A1(n7513), .A2(P2_U3152), .B1(n8719), .B2(n7512), .C1(
        n7511), .C2(n8722), .ZN(P2_U3334) );
  MUX2_X1 U9218 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n5129), .S(n8887), .Z(n8894)
         );
  INV_X1 U9219 ( .A(n7514), .ZN(n7515) );
  OAI21_X1 U9220 ( .B1(n7517), .B2(n7516), .A(n7515), .ZN(n8893) );
  NAND2_X1 U9221 ( .A1(n8894), .A2(n8893), .ZN(n8892) );
  NAND2_X1 U9222 ( .A1(n7518), .A2(n7521), .ZN(n7519) );
  NAND2_X1 U9223 ( .A1(n7519), .A2(n9655), .ZN(n8898) );
  XNOR2_X1 U9224 ( .A(n8898), .B(n8905), .ZN(n7520) );
  NOR2_X1 U9225 ( .A1(n5175), .A2(n7520), .ZN(n8899) );
  AOI211_X1 U9226 ( .C1(n7520), .C2(n5175), .A(n8899), .B(n9626), .ZN(n7530)
         );
  INV_X1 U9227 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9540) );
  AOI22_X1 U9228 ( .A1(n9653), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n9540), .B2(
        n7521), .ZN(n9658) );
  INV_X1 U9229 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7522) );
  MUX2_X1 U9230 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n7522), .S(n8887), .Z(n8890)
         );
  OAI21_X1 U9231 ( .B1(n7524), .B2(P1_REG1_REG_12__SCAN_IN), .A(n7523), .ZN(
        n8889) );
  NAND2_X1 U9232 ( .A1(n8890), .A2(n8889), .ZN(n8888) );
  OAI21_X1 U9233 ( .B1(n8887), .B2(P1_REG1_REG_13__SCAN_IN), .A(n8888), .ZN(
        n9659) );
  NAND2_X1 U9234 ( .A1(n9658), .A2(n9659), .ZN(n9657) );
  OAI21_X1 U9235 ( .B1(n9653), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9657), .ZN(
        n8904) );
  XNOR2_X1 U9236 ( .A(n8905), .B(n8904), .ZN(n7526) );
  INV_X1 U9237 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7525) );
  NOR2_X1 U9238 ( .A1(n7525), .A2(n7526), .ZN(n8906) );
  AOI211_X1 U9239 ( .C1(n7526), .C2(n7525), .A(n8906), .B(n9575), .ZN(n7529)
         );
  NAND2_X1 U9240 ( .A1(n8933), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9241 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8846) );
  OAI211_X1 U9242 ( .C1(n8905), .C2(n9634), .A(n7527), .B(n8846), .ZN(n7528)
         );
  OR3_X1 U9243 ( .A1(n7530), .A2(n7529), .A3(n7528), .ZN(P1_U3256) );
  XOR2_X1 U9244 ( .A(n7531), .B(n7776), .Z(n9539) );
  INV_X1 U9245 ( .A(n9539), .ZN(n7544) );
  NAND2_X1 U9246 ( .A1(n7532), .A2(n9701), .ZN(n7536) );
  INV_X1 U9247 ( .A(n7856), .ZN(n7862) );
  INV_X1 U9248 ( .A(n7776), .ZN(n7533) );
  AOI21_X1 U9249 ( .B1(n9492), .B2(n7862), .A(n7533), .ZN(n7535) );
  AOI22_X1 U9250 ( .A1(n9154), .A2(n8860), .B1(n8858), .B2(n9152), .ZN(n7534)
         );
  OAI21_X1 U9251 ( .B1(n7536), .B2(n7535), .A(n7534), .ZN(n9537) );
  INV_X1 U9252 ( .A(n7642), .ZN(n7537) );
  OAI211_X1 U9253 ( .C1(n9536), .C2(n9488), .A(n7537), .B(n9526), .ZN(n9535)
         );
  INV_X1 U9254 ( .A(n7538), .ZN(n7671) );
  OAI22_X1 U9255 ( .A1(n9684), .A2(n7539), .B1(n7671), .B2(n9105), .ZN(n7540)
         );
  AOI21_X1 U9256 ( .B1(n7673), .B2(n9107), .A(n7540), .ZN(n7541) );
  OAI21_X1 U9257 ( .B1(n9535), .B2(n7660), .A(n7541), .ZN(n7542) );
  AOI21_X1 U9258 ( .B1(n9537), .B2(n9684), .A(n7542), .ZN(n7543) );
  OAI21_X1 U9259 ( .B1(n7544), .B2(n9176), .A(n7543), .ZN(P1_U3277) );
  OAI21_X1 U9260 ( .B1(n7547), .B2(n7546), .A(n7545), .ZN(n7548) );
  NAND2_X1 U9261 ( .A1(n7548), .A2(n8829), .ZN(n7554) );
  INV_X1 U9262 ( .A(n7549), .ZN(n7552) );
  OAI22_X1 U9263 ( .A1(n8833), .A2(n7550), .B1(n7708), .B2(n8807), .ZN(n7551)
         );
  AOI211_X1 U9264 ( .C1(n8831), .C2(n8862), .A(n7552), .B(n7551), .ZN(n7553)
         );
  OAI211_X1 U9265 ( .C1(n9548), .C2(n8837), .A(n7554), .B(n7553), .ZN(P1_U3222) );
  NOR3_X1 U9266 ( .A1(n7555), .A2(n7619), .A3(n8194), .ZN(n7556) );
  AOI21_X1 U9267 ( .B1(n7557), .B2(n8181), .A(n7556), .ZN(n7566) );
  INV_X1 U9268 ( .A(n7622), .ZN(n7560) );
  INV_X1 U9269 ( .A(n8200), .ZN(n8174) );
  INV_X1 U9270 ( .A(n7619), .ZN(n8226) );
  AOI22_X1 U9271 ( .A1(n8175), .A2(n4668), .B1(n8174), .B2(n8226), .ZN(n7559)
         );
  OAI211_X1 U9272 ( .C1(n7560), .C2(n8198), .A(n7559), .B(n7558), .ZN(n7563)
         );
  NOR2_X1 U9273 ( .A1(n7561), .A2(n8216), .ZN(n7562) );
  AOI211_X1 U9274 ( .C1(n7620), .C2(n8214), .A(n7563), .B(n7562), .ZN(n7564)
         );
  OAI21_X1 U9275 ( .B1(n7566), .B2(n7565), .A(n7564), .ZN(P2_U3217) );
  INV_X1 U9276 ( .A(n7567), .ZN(n7583) );
  AOI22_X1 U9277 ( .A1(n7568), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n9416), .ZN(n7569) );
  OAI21_X1 U9278 ( .B1(n7583), .B2(n6758), .A(n7569), .ZN(P1_U3328) );
  NAND2_X1 U9279 ( .A1(n4335), .A2(n7570), .ZN(n7571) );
  XNOR2_X1 U9280 ( .A(n7572), .B(n7571), .ZN(n7578) );
  NAND2_X1 U9281 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8884) );
  INV_X1 U9282 ( .A(n8884), .ZN(n7575) );
  INV_X1 U9283 ( .A(n9500), .ZN(n7573) );
  OAI22_X1 U9284 ( .A1(n8833), .A2(n7573), .B1(n9495), .B2(n8807), .ZN(n7574)
         );
  AOI211_X1 U9285 ( .C1(n8831), .C2(n8861), .A(n7575), .B(n7574), .ZN(n7577)
         );
  NAND2_X1 U9286 ( .A1(n9486), .A2(n8850), .ZN(n7576) );
  OAI211_X1 U9287 ( .C1(n7578), .C2(n8853), .A(n7577), .B(n7576), .ZN(P1_U3232) );
  INV_X1 U9288 ( .A(n7579), .ZN(n7586) );
  AOI22_X1 U9289 ( .A1(n7580), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n9416), .ZN(n7581) );
  OAI21_X1 U9290 ( .B1(n7586), .B2(n6758), .A(n7581), .ZN(P1_U3327) );
  OAI222_X1 U9291 ( .A1(n8722), .A2(n7584), .B1(n8719), .B2(n7583), .C1(n7582), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9292 ( .A1(n7587), .A2(P2_U3152), .B1(n8719), .B2(n7586), .C1(
        n7585), .C2(n8722), .ZN(P2_U3332) );
  INV_X1 U9293 ( .A(n7588), .ZN(n8228) );
  NAND2_X1 U9294 ( .A1(n7589), .A2(n8228), .ZN(n7590) );
  AND2_X2 U9295 ( .A1(n7591), .A2(n7590), .ZN(n9806) );
  INV_X1 U9296 ( .A(n7600), .ZN(n8227) );
  OR2_X1 U9297 ( .A1(n9928), .A2(n8227), .ZN(n7593) );
  AND2_X1 U9298 ( .A1(n7594), .A2(n7598), .ZN(n7595) );
  OR2_X1 U9299 ( .A1(n7615), .A2(n7595), .ZN(n7606) );
  INV_X1 U9300 ( .A(n7596), .ZN(n7599) );
  OAI21_X1 U9301 ( .B1(n7599), .B2(n7598), .A(n7597), .ZN(n7603) );
  OAI22_X1 U9302 ( .A1(n7601), .A2(n8538), .B1(n7600), .B2(n8536), .ZN(n7602)
         );
  AOI21_X1 U9303 ( .B1(n7603), .B2(n9830), .A(n7602), .ZN(n7604) );
  OAI21_X1 U9304 ( .B1(n7606), .B2(n7605), .A(n7604), .ZN(n9475) );
  INV_X1 U9305 ( .A(n9475), .ZN(n7613) );
  INV_X1 U9306 ( .A(n7606), .ZN(n9477) );
  AND2_X1 U9307 ( .A1(n9808), .A2(n7614), .ZN(n7607) );
  OR2_X1 U9308 ( .A1(n7607), .A2(n4282), .ZN(n9474) );
  NOR2_X1 U9309 ( .A1(n9474), .A2(n8387), .ZN(n7611) );
  AOI22_X1 U9310 ( .A1(n8495), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7608), .B2(
        n9839), .ZN(n7609) );
  OAI21_X1 U9311 ( .B1(n4598), .B2(n9817), .A(n7609), .ZN(n7610) );
  AOI211_X1 U9312 ( .C1(n9477), .C2(n9824), .A(n7611), .B(n7610), .ZN(n7612)
         );
  OAI21_X1 U9313 ( .B1(n7613), .B2(n9840), .A(n7612), .ZN(P2_U3283) );
  OAI21_X1 U9314 ( .B1(n4333), .B2(n7616), .A(n7990), .ZN(n9471) );
  INV_X1 U9315 ( .A(n9471), .ZN(n7627) );
  XNOR2_X1 U9316 ( .A(n7617), .B(n7616), .ZN(n7618) );
  OAI222_X1 U9317 ( .A1(n8536), .A2(n7619), .B1(n8538), .B2(n8126), .C1(n8533), 
        .C2(n7618), .ZN(n9470) );
  INV_X1 U9318 ( .A(n7620), .ZN(n9467) );
  INV_X1 U9319 ( .A(n8611), .ZN(n7621) );
  OAI21_X1 U9320 ( .B1(n9467), .B2(n4282), .A(n7621), .ZN(n9468) );
  NOR2_X1 U9321 ( .A1(n9468), .A2(n8387), .ZN(n7625) );
  AOI22_X1 U9322 ( .A1(n9840), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7622), .B2(
        n9839), .ZN(n7623) );
  OAI21_X1 U9323 ( .B1(n9467), .B2(n9817), .A(n7623), .ZN(n7624) );
  AOI211_X1 U9324 ( .C1(n9470), .C2(n9815), .A(n7625), .B(n7624), .ZN(n7626)
         );
  OAI21_X1 U9325 ( .B1(n7627), .B2(n8604), .A(n7626), .ZN(P2_U3282) );
  NAND2_X1 U9326 ( .A1(n7628), .A2(n7870), .ZN(n7629) );
  NAND2_X1 U9327 ( .A1(n7630), .A2(n7629), .ZN(n7641) );
  OR2_X1 U9328 ( .A1(n7641), .A2(n9704), .ZN(n7640) );
  NAND2_X1 U9329 ( .A1(n7632), .A2(n7631), .ZN(n7633) );
  NAND2_X1 U9330 ( .A1(n7634), .A2(n7633), .ZN(n7638) );
  NAND2_X1 U9331 ( .A1(n8857), .A2(n9152), .ZN(n7636) );
  NAND2_X1 U9332 ( .A1(n8859), .A2(n9154), .ZN(n7635) );
  NAND2_X1 U9333 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  AOI21_X1 U9334 ( .B1(n7638), .B2(n9701), .A(n7637), .ZN(n7639) );
  INV_X1 U9335 ( .A(n7641), .ZN(n9251) );
  NOR2_X1 U9336 ( .A1(n7642), .A2(n9248), .ZN(n7643) );
  OR2_X1 U9337 ( .A1(n7657), .A2(n7643), .ZN(n9249) );
  AOI22_X1 U9338 ( .A1(n9708), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8845), .B2(
        n9707), .ZN(n7645) );
  NAND2_X1 U9339 ( .A1(n8851), .A2(n9107), .ZN(n7644) );
  OAI211_X1 U9340 ( .C1(n9249), .C2(n8985), .A(n7645), .B(n7644), .ZN(n7646)
         );
  AOI21_X1 U9341 ( .B1(n9251), .B2(n9693), .A(n7646), .ZN(n7647) );
  OAI21_X1 U9342 ( .B1(n9253), .B2(n9708), .A(n7647), .ZN(P1_U3276) );
  INV_X1 U9343 ( .A(n7648), .ZN(n7663) );
  AOI22_X1 U9344 ( .A1(n7649), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n9416), .ZN(n7650) );
  OAI21_X1 U9345 ( .B1(n7663), .B2(n6758), .A(n7650), .ZN(P1_U3326) );
  OAI21_X1 U9346 ( .B1(n7652), .B2(n7872), .A(n7651), .ZN(n9528) );
  INV_X1 U9347 ( .A(n7872), .ZN(n7778) );
  XNOR2_X1 U9348 ( .A(n7653), .B(n7778), .ZN(n7654) );
  NAND2_X1 U9349 ( .A1(n7654), .A2(n9701), .ZN(n7656) );
  AOI22_X1 U9350 ( .A1(n9154), .A2(n8858), .B1(n9155), .B2(n9152), .ZN(n7655)
         );
  NAND2_X1 U9351 ( .A1(n7656), .A2(n7655), .ZN(n9532) );
  OAI211_X1 U9352 ( .C1(n7657), .C2(n9531), .A(n9526), .B(n9169), .ZN(n9530)
         );
  AOI22_X1 U9353 ( .A1(n9708), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8758), .B2(
        n9707), .ZN(n7659) );
  NAND2_X1 U9354 ( .A1(n8762), .A2(n9107), .ZN(n7658) );
  OAI211_X1 U9355 ( .C1(n9530), .C2(n7660), .A(n7659), .B(n7658), .ZN(n7661)
         );
  AOI21_X1 U9356 ( .B1(n9532), .B2(n9684), .A(n7661), .ZN(n7662) );
  OAI21_X1 U9357 ( .B1(n9528), .B2(n9176), .A(n7662), .ZN(P1_U3275) );
  OAI222_X1 U9358 ( .A1(n8722), .A2(n7664), .B1(n8719), .B2(n7663), .C1(n8004), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9359 ( .A(n7665), .ZN(n7667) );
  NAND2_X1 U9360 ( .A1(n7667), .A2(n7666), .ZN(n7669) );
  XNOR2_X1 U9361 ( .A(n7669), .B(n7668), .ZN(n7676) );
  NOR2_X1 U9362 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7670), .ZN(n9652) );
  OAI22_X1 U9363 ( .A1(n8833), .A2(n7671), .B1(n8757), .B2(n8807), .ZN(n7672)
         );
  AOI211_X1 U9364 ( .C1(n8831), .C2(n8860), .A(n9652), .B(n7672), .ZN(n7675)
         );
  NAND2_X1 U9365 ( .A1(n7673), .A2(n8850), .ZN(n7674) );
  OAI211_X1 U9366 ( .C1(n7676), .C2(n8853), .A(n7675), .B(n7674), .ZN(P1_U3213) );
  NAND2_X1 U9367 ( .A1(n9405), .A2(n7684), .ZN(n7678) );
  NAND2_X1 U9368 ( .A1(n5435), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7677) );
  INV_X1 U9369 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U9370 ( .A1(n4267), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n7682) );
  INV_X1 U9371 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n7679) );
  OR2_X1 U9372 ( .A1(n7680), .A2(n7679), .ZN(n7681) );
  OAI211_X1 U9373 ( .C1(n7683), .C2(n8963), .A(n7682), .B(n7681), .ZN(n8962)
         );
  INV_X1 U9374 ( .A(n8962), .ZN(n7756) );
  NAND2_X1 U9375 ( .A1(n5435), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7685) );
  INV_X1 U9376 ( .A(n8855), .ZN(n7687) );
  NAND2_X1 U9377 ( .A1(n8967), .A2(n7687), .ZN(n7686) );
  NAND2_X1 U9378 ( .A1(n7955), .A2(n7686), .ZN(n7793) );
  NAND2_X1 U9379 ( .A1(n7924), .A2(n7688), .ZN(n7689) );
  NAND3_X1 U9380 ( .A1(n7929), .A2(n7925), .A3(n7689), .ZN(n7819) );
  NAND2_X1 U9381 ( .A1(n7924), .A2(n7915), .ZN(n7817) );
  NAND2_X1 U9382 ( .A1(n7747), .A2(n7690), .ZN(n7911) );
  AND2_X1 U9383 ( .A1(n9226), .A2(n9099), .ZN(n7895) );
  NAND2_X1 U9384 ( .A1(n7695), .A2(n7895), .ZN(n7691) );
  NAND2_X1 U9385 ( .A1(n7903), .A2(n7691), .ZN(n7697) );
  OR2_X1 U9386 ( .A1(n7697), .A2(n4550), .ZN(n7811) );
  AND2_X1 U9387 ( .A1(n7885), .A2(n7692), .ZN(n7889) );
  INV_X1 U9388 ( .A(n7889), .ZN(n7693) );
  NAND2_X1 U9389 ( .A1(n7693), .A2(n7892), .ZN(n7694) );
  NOR2_X1 U9390 ( .A1(n7811), .A2(n7694), .ZN(n7699) );
  NAND2_X1 U9391 ( .A1(n7695), .A2(n7900), .ZN(n7901) );
  INV_X1 U9392 ( .A(n7896), .ZN(n7887) );
  NOR2_X1 U9393 ( .A1(n7901), .A2(n7887), .ZN(n7696) );
  OAI21_X1 U9394 ( .B1(n7697), .B2(n7696), .A(n7906), .ZN(n7698) );
  NAND2_X1 U9395 ( .A1(n9243), .A2(n8806), .ZN(n7879) );
  AND2_X1 U9396 ( .A1(n7876), .A2(n7879), .ZN(n7700) );
  NAND2_X1 U9397 ( .A1(n7892), .A2(n7700), .ZN(n7719) );
  INV_X1 U9398 ( .A(n7701), .ZN(n7871) );
  INV_X1 U9399 ( .A(n7863), .ZN(n7702) );
  OR3_X1 U9400 ( .A1(n7719), .A2(n7871), .A3(n7702), .ZN(n7740) );
  INV_X1 U9401 ( .A(n7860), .ZN(n7703) );
  OR2_X1 U9402 ( .A1(n7856), .A2(n7703), .ZN(n7710) );
  NOR2_X1 U9403 ( .A1(n7710), .A2(n7760), .ZN(n7853) );
  INV_X1 U9404 ( .A(n7853), .ZN(n7738) );
  NAND2_X1 U9405 ( .A1(n7705), .A2(n7704), .ZN(n7842) );
  AND2_X1 U9406 ( .A1(n7847), .A2(n7842), .ZN(n7735) );
  AND2_X1 U9407 ( .A1(n7837), .A2(n7706), .ZN(n7840) );
  INV_X1 U9408 ( .A(n7840), .ZN(n7707) );
  AOI21_X1 U9409 ( .B1(n7735), .B2(n7707), .A(n7848), .ZN(n7716) );
  OR2_X1 U9410 ( .A1(n9486), .A2(n7708), .ZN(n7709) );
  AND2_X1 U9411 ( .A1(n7865), .A2(n7709), .ZN(n7866) );
  INV_X1 U9412 ( .A(n7710), .ZN(n7714) );
  INV_X1 U9413 ( .A(n7761), .ZN(n7711) );
  NOR2_X1 U9414 ( .A1(n7712), .A2(n7711), .ZN(n7858) );
  INV_X1 U9415 ( .A(n7858), .ZN(n7713) );
  NAND2_X1 U9416 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  OAI211_X1 U9417 ( .C1(n7738), .C2(n7716), .A(n7866), .B(n7715), .ZN(n7717)
         );
  INV_X1 U9418 ( .A(n7717), .ZN(n7720) );
  AND2_X1 U9419 ( .A1(n7877), .A2(n7718), .ZN(n7874) );
  OAI22_X1 U9420 ( .A1(n7740), .A2(n7720), .B1(n7874), .B2(n7719), .ZN(n7807)
         );
  INV_X1 U9421 ( .A(n7807), .ZN(n7744) );
  INV_X1 U9422 ( .A(n7763), .ZN(n7721) );
  AND2_X1 U9423 ( .A1(n7721), .A2(n7956), .ZN(n7724) );
  OAI211_X1 U9424 ( .C1(n7725), .C2(n7724), .A(n7723), .B(n7722), .ZN(n7727)
         );
  NAND3_X1 U9425 ( .A1(n7727), .A2(n7799), .A3(n7726), .ZN(n7731) );
  AND3_X1 U9426 ( .A1(n7729), .A2(n7831), .A3(n7728), .ZN(n7803) );
  INV_X1 U9427 ( .A(n7803), .ZN(n7730) );
  AOI21_X1 U9428 ( .B1(n7731), .B2(n7798), .A(n7730), .ZN(n7742) );
  INV_X1 U9429 ( .A(n7732), .ZN(n7733) );
  NAND2_X1 U9430 ( .A1(n7831), .A2(n7733), .ZN(n7734) );
  AND3_X1 U9431 ( .A1(n7734), .A2(n7833), .A3(n7828), .ZN(n7805) );
  INV_X1 U9432 ( .A(n7805), .ZN(n7741) );
  INV_X1 U9433 ( .A(n7735), .ZN(n7736) );
  OR4_X1 U9434 ( .A1(n7738), .A2(n7737), .A3(n4531), .A4(n7736), .ZN(n7739) );
  NOR2_X1 U9435 ( .A1(n7740), .A2(n7739), .ZN(n7809) );
  OAI21_X1 U9436 ( .B1(n7742), .B2(n7741), .A(n7809), .ZN(n7743) );
  AND2_X1 U9437 ( .A1(n7744), .A2(n7743), .ZN(n7745) );
  NOR2_X1 U9438 ( .A1(n7811), .A2(n7745), .ZN(n7749) );
  NAND2_X1 U9439 ( .A1(n9211), .A2(n8796), .ZN(n7746) );
  NAND2_X1 U9440 ( .A1(n9015), .A2(n7746), .ZN(n7908) );
  NAND2_X1 U9441 ( .A1(n7908), .A2(n7747), .ZN(n7748) );
  NAND2_X1 U9442 ( .A1(n9016), .A2(n7748), .ZN(n7914) );
  INV_X1 U9443 ( .A(n7914), .ZN(n7812) );
  INV_X1 U9444 ( .A(n7750), .ZN(n7751) );
  NOR2_X1 U9445 ( .A1(n7817), .A2(n7751), .ZN(n7752) );
  NOR2_X1 U9446 ( .A1(n7819), .A2(n7752), .ZN(n7754) );
  NAND2_X1 U9447 ( .A1(n7753), .A2(n7928), .ZN(n7822) );
  OAI21_X1 U9448 ( .B1(n7754), .B2(n7822), .A(n7821), .ZN(n7755) );
  AND2_X1 U9449 ( .A1(n7796), .A2(n7755), .ZN(n7757) );
  OAI21_X1 U9450 ( .B1(n7793), .B2(n7757), .A(n7791), .ZN(n7758) );
  XNOR2_X1 U9451 ( .A(n7758), .B(n7953), .ZN(n7958) );
  INV_X1 U9452 ( .A(n7759), .ZN(n7790) );
  INV_X1 U9453 ( .A(n9042), .ZN(n9052) );
  INV_X1 U9454 ( .A(n7760), .ZN(n7762) );
  AND2_X1 U9455 ( .A1(n7762), .A2(n7761), .ZN(n9509) );
  OR2_X1 U9456 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  NOR2_X1 U9457 ( .A1(n7765), .A2(n9694), .ZN(n7769) );
  INV_X1 U9458 ( .A(n7766), .ZN(n7767) );
  AND4_X1 U9459 ( .A1(n7769), .A2(n4980), .A3(n7768), .A4(n7767), .ZN(n7771)
         );
  NAND4_X1 U9460 ( .A1(n7771), .A2(n4674), .A3(n7839), .A4(n7770), .ZN(n7772)
         );
  NOR2_X1 U9461 ( .A1(n7772), .A2(n7845), .ZN(n7773) );
  NAND4_X1 U9462 ( .A1(n7774), .A2(n9509), .A3(n7773), .A4(n9674), .ZN(n7775)
         );
  NOR3_X1 U9463 ( .A1(n7776), .A2(n4534), .A3(n7775), .ZN(n7777) );
  NAND4_X1 U9464 ( .A1(n9161), .A2(n7870), .A3(n7778), .A4(n7777), .ZN(n7779)
         );
  NOR2_X1 U9465 ( .A1(n9149), .A2(n7779), .ZN(n7780) );
  INV_X1 U9466 ( .A(n9111), .ZN(n9119) );
  NAND4_X1 U9467 ( .A1(n7781), .A2(n9136), .A3(n7780), .A4(n9119), .ZN(n7782)
         );
  NOR2_X1 U9468 ( .A1(n9087), .A2(n7782), .ZN(n7783) );
  NAND4_X1 U9469 ( .A1(n9028), .A2(n9052), .A3(n7783), .A4(n9069), .ZN(n7787)
         );
  INV_X1 U9470 ( .A(n7784), .ZN(n7785) );
  OR3_X1 U9471 ( .A1(n7787), .A2(n8999), .A3(n9019), .ZN(n7788) );
  NOR2_X1 U9472 ( .A1(n8975), .A2(n7788), .ZN(n7789) );
  NAND4_X1 U9473 ( .A1(n7791), .A2(n7790), .A3(n7789), .A4(n7796), .ZN(n7792)
         );
  OR2_X1 U9474 ( .A1(n7793), .A2(n7792), .ZN(n7795) );
  AND2_X1 U9475 ( .A1(n7795), .A2(n7794), .ZN(n7951) );
  INV_X1 U9476 ( .A(n7951), .ZN(n7827) );
  NAND2_X1 U9477 ( .A1(n7796), .A2(n8962), .ZN(n7797) );
  NAND2_X1 U9478 ( .A1(n7797), .A2(n9177), .ZN(n7947) );
  INV_X1 U9479 ( .A(n7798), .ZN(n7804) );
  INV_X1 U9480 ( .A(n7799), .ZN(n7801) );
  NAND2_X1 U9481 ( .A1(n7801), .A2(n7800), .ZN(n7802) );
  OAI211_X1 U9482 ( .C1(n9695), .C2(n7804), .A(n7803), .B(n7802), .ZN(n7806)
         );
  NAND2_X1 U9483 ( .A1(n7806), .A2(n7805), .ZN(n7808) );
  AOI21_X1 U9484 ( .B1(n7809), .B2(n7808), .A(n7807), .ZN(n7810) );
  NOR2_X1 U9485 ( .A1(n7811), .A2(n7810), .ZN(n7813) );
  OAI21_X1 U9486 ( .B1(n7814), .B2(n7813), .A(n7812), .ZN(n7815) );
  INV_X1 U9487 ( .A(n7815), .ZN(n7816) );
  NOR2_X1 U9488 ( .A1(n7817), .A2(n7816), .ZN(n7818) );
  NOR2_X1 U9489 ( .A1(n7819), .A2(n7818), .ZN(n7823) );
  NAND2_X1 U9490 ( .A1(n8962), .A2(n8855), .ZN(n7820) );
  NAND2_X1 U9491 ( .A1(n8967), .A2(n7820), .ZN(n7944) );
  OAI211_X1 U9492 ( .C1(n7823), .C2(n7822), .A(n7944), .B(n7821), .ZN(n7824)
         );
  NAND2_X1 U9493 ( .A1(n7947), .A2(n7824), .ZN(n7825) );
  NAND3_X1 U9494 ( .A1(n7825), .A2(n7956), .A3(n7955), .ZN(n7826) );
  NAND2_X1 U9495 ( .A1(n7827), .A2(n7826), .ZN(n7954) );
  NAND2_X1 U9496 ( .A1(n7829), .A2(n7828), .ZN(n7832) );
  NAND3_X1 U9497 ( .A1(n7832), .A2(n7831), .A3(n7830), .ZN(n7834) );
  NAND3_X1 U9498 ( .A1(n7834), .A2(n7839), .A3(n7833), .ZN(n7836) );
  NAND3_X1 U9499 ( .A1(n7836), .A2(n7842), .A3(n7835), .ZN(n7838) );
  NAND2_X1 U9500 ( .A1(n7838), .A2(n7837), .ZN(n7844) );
  OAI21_X1 U9501 ( .B1(n7841), .B2(n5504), .A(n7840), .ZN(n7843) );
  INV_X1 U9502 ( .A(n7845), .ZN(n7846) );
  INV_X1 U9503 ( .A(n7847), .ZN(n7849) );
  MUX2_X1 U9504 ( .A(n7849), .B(n7848), .S(n7941), .Z(n7850) );
  INV_X1 U9505 ( .A(n7850), .ZN(n7851) );
  NAND2_X1 U9506 ( .A1(n7852), .A2(n9509), .ZN(n7859) );
  NAND2_X1 U9507 ( .A1(n7859), .A2(n7853), .ZN(n7854) );
  OAI211_X1 U9508 ( .C1(n7856), .C2(n7855), .A(n7854), .B(n7866), .ZN(n7857)
         );
  NAND2_X1 U9509 ( .A1(n7857), .A2(n7863), .ZN(n7869) );
  NAND2_X1 U9510 ( .A1(n7859), .A2(n7858), .ZN(n7861) );
  NAND2_X1 U9511 ( .A1(n7861), .A2(n7860), .ZN(n7867) );
  NAND2_X1 U9512 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  AOI22_X1 U9513 ( .A1(n7867), .A2(n7866), .B1(n7865), .B2(n7864), .ZN(n7868)
         );
  NOR2_X1 U9514 ( .A1(n7872), .A2(n7871), .ZN(n7873) );
  MUX2_X1 U9515 ( .A(n7874), .B(n7873), .S(n7943), .Z(n7875) );
  MUX2_X1 U9516 ( .A(n7877), .B(n7876), .S(n7941), .Z(n7878) );
  OAI211_X1 U9517 ( .C1(n7890), .C2(n9155), .A(n7892), .B(n7879), .ZN(n7880)
         );
  NAND2_X1 U9518 ( .A1(n7880), .A2(n7943), .ZN(n7884) );
  INV_X1 U9519 ( .A(n7890), .ZN(n7882) );
  NAND2_X1 U9520 ( .A1(n7882), .A2(n4686), .ZN(n7883) );
  NAND2_X1 U9521 ( .A1(n7884), .A2(n7883), .ZN(n7894) );
  AOI21_X1 U9522 ( .B1(n7894), .B2(n7885), .A(n4550), .ZN(n7888) );
  INV_X1 U9523 ( .A(n7895), .ZN(n7886) );
  OAI21_X1 U9524 ( .B1(n7888), .B2(n7887), .A(n7886), .ZN(n7899) );
  OAI21_X1 U9525 ( .B1(n7890), .B2(n9243), .A(n7889), .ZN(n7893) );
  OAI211_X1 U9526 ( .C1(n7894), .C2(n7893), .A(n7892), .B(n7891), .ZN(n7897)
         );
  AOI21_X1 U9527 ( .B1(n7897), .B2(n7896), .A(n7895), .ZN(n7898) );
  NAND2_X1 U9528 ( .A1(n7901), .A2(n9085), .ZN(n7902) );
  AND2_X1 U9529 ( .A1(n7906), .A2(n7902), .ZN(n7904) );
  MUX2_X1 U9530 ( .A(n7904), .B(n7903), .S(n7941), .Z(n7905) );
  MUX2_X1 U9531 ( .A(n7907), .B(n7906), .S(n7941), .Z(n7910) );
  OR2_X1 U9532 ( .A1(n7911), .A2(n7908), .ZN(n7909) );
  NAND2_X1 U9533 ( .A1(n7911), .A2(n9015), .ZN(n7912) );
  NAND2_X1 U9534 ( .A1(n9017), .A2(n7912), .ZN(n7913) );
  MUX2_X1 U9535 ( .A(n7914), .B(n7913), .S(n7941), .Z(n7917) );
  MUX2_X1 U9536 ( .A(n9016), .B(n7915), .S(n7943), .Z(n7916) );
  OAI21_X1 U9537 ( .B1(n7918), .B2(n7917), .A(n7916), .ZN(n7920) );
  MUX2_X1 U9538 ( .A(n7941), .B(n7920), .S(n7919), .Z(n7923) );
  OR3_X1 U9539 ( .A1(n9196), .A2(n9031), .A3(n7943), .ZN(n7921) );
  NAND3_X1 U9540 ( .A1(n7923), .A2(n7922), .A3(n7921), .ZN(n7927) );
  MUX2_X1 U9541 ( .A(n7925), .B(n7924), .S(n7943), .Z(n7926) );
  NAND3_X1 U9542 ( .A1(n7927), .A2(n8972), .A3(n7926), .ZN(n7931) );
  MUX2_X1 U9543 ( .A(n7929), .B(n7928), .S(n7941), .Z(n7930) );
  AND2_X1 U9544 ( .A1(n7931), .A2(n7930), .ZN(n7937) );
  NAND3_X1 U9545 ( .A1(n7937), .A2(n8979), .A3(n7944), .ZN(n7932) );
  NAND2_X1 U9546 ( .A1(n7932), .A2(n7947), .ZN(n7936) );
  NAND3_X1 U9547 ( .A1(n7947), .A2(n7937), .A3(n9180), .ZN(n7934) );
  AOI21_X1 U9548 ( .B1(n7934), .B2(n7944), .A(n7933), .ZN(n7935) );
  MUX2_X1 U9549 ( .A(n7936), .B(n7935), .S(n7941), .Z(n7949) );
  INV_X1 U9550 ( .A(n7937), .ZN(n7940) );
  NAND3_X1 U9551 ( .A1(n7940), .A2(n7939), .A3(n7938), .ZN(n7946) );
  AND2_X1 U9552 ( .A1(n8979), .A2(n7941), .ZN(n7942) );
  AOI21_X1 U9553 ( .B1(n9180), .B2(n7943), .A(n7942), .ZN(n7945) );
  AND4_X1 U9554 ( .A1(n7947), .A2(n7946), .A3(n7945), .A4(n7944), .ZN(n7948)
         );
  AND2_X1 U9555 ( .A1(n7955), .A2(n7950), .ZN(n7952) );
  NOR4_X1 U9556 ( .A1(n7961), .A2(n7960), .A3(n7959), .A4(n9584), .ZN(n7962)
         );
  AOI211_X1 U9557 ( .C1(n7965), .C2(n6340), .A(n7963), .B(n7962), .ZN(n7964)
         );
  NAND2_X1 U9558 ( .A1(n7966), .A2(n8181), .ZN(n7978) );
  INV_X1 U9559 ( .A(n8612), .ZN(n7970) );
  OR2_X1 U9560 ( .A1(n8137), .A2(n8538), .ZN(n7968) );
  NAND2_X1 U9561 ( .A1(n8225), .A2(n8571), .ZN(n7967) );
  NAND2_X1 U9562 ( .A1(n7968), .A2(n7967), .ZN(n8606) );
  AOI22_X1 U9563 ( .A1(n8129), .A2(n8606), .B1(P2_REG3_REG_15__SCAN_IN), .B2(
        P2_U3152), .ZN(n7969) );
  OAI21_X1 U9564 ( .B1(n7970), .B2(n8198), .A(n7969), .ZN(n7975) );
  INV_X1 U9565 ( .A(n7971), .ZN(n7973) );
  AOI211_X1 U9566 ( .C1(n7973), .C2(n7972), .A(n8126), .B(n8194), .ZN(n7974)
         );
  AOI211_X1 U9567 ( .C1(n7976), .C2(n8214), .A(n7975), .B(n7974), .ZN(n7977)
         );
  OAI21_X1 U9568 ( .B1(n8124), .B2(n7978), .A(n7977), .ZN(P2_U3243) );
  INV_X1 U9569 ( .A(n7979), .ZN(n9412) );
  XOR2_X1 U9570 ( .A(n7983), .B(n7982), .Z(n7984) );
  XNOR2_X1 U9571 ( .A(n4310), .B(n7984), .ZN(n7988) );
  NAND2_X1 U9572 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8957) );
  OAI21_X1 U9573 ( .B1(n8807), .B2(n9099), .A(n8957), .ZN(n7986) );
  OAI22_X1 U9574 ( .A1(n8833), .A2(n9130), .B1(n8848), .B2(n9166), .ZN(n7985)
         );
  AOI211_X1 U9575 ( .C1(n9232), .C2(n8850), .A(n7986), .B(n7985), .ZN(n7987)
         );
  OAI21_X1 U9576 ( .B1(n7988), .B2(n8853), .A(n7987), .ZN(P1_U3217) );
  INV_X1 U9577 ( .A(n8692), .ZN(n8596) );
  INV_X1 U9578 ( .A(n8138), .ZN(n8224) );
  NOR2_X1 U9579 ( .A1(n8677), .A2(n8573), .ZN(n7993) );
  INV_X1 U9580 ( .A(n8677), .ZN(n8553) );
  INV_X1 U9581 ( .A(n8101), .ZN(n8223) );
  INV_X1 U9582 ( .A(n8539), .ZN(n8222) );
  NAND2_X1 U9583 ( .A1(n8524), .A2(n8539), .ZN(n7994) );
  NAND2_X1 U9584 ( .A1(n7995), .A2(n7994), .ZN(n8496) );
  AOI22_X2 U9585 ( .A1(n8496), .A2(n8504), .B1(n8503), .B2(n8106), .ZN(n8483)
         );
  NAND2_X2 U9586 ( .A1(n8447), .A2(n8455), .ZN(n7999) );
  XNOR2_X1 U9587 ( .A(n8000), .B(n8002), .ZN(n8629) );
  INV_X1 U9588 ( .A(P2_B_REG_SCAN_IN), .ZN(n8003) );
  NOR2_X1 U9589 ( .A1(n8004), .A2(n8003), .ZN(n8005) );
  NOR2_X1 U9590 ( .A1(n8538), .A2(n8005), .ZN(n8382) );
  AOI22_X1 U9591 ( .A1(n4471), .A2(n8571), .B1(n8382), .B2(n8218), .ZN(n8006)
         );
  INV_X1 U9592 ( .A(n8628), .ZN(n8010) );
  NOR2_X1 U9593 ( .A1(n8528), .A2(n8668), .ZN(n8497) );
  NAND2_X1 U9594 ( .A1(n8627), .A2(n9811), .ZN(n8009) );
  AOI22_X1 U9595 ( .A1(n8007), .A2(n9839), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8495), .ZN(n8008) );
  OAI211_X1 U9596 ( .C1(n8010), .C2(n9817), .A(n8009), .B(n8008), .ZN(n8011)
         );
  AOI21_X1 U9597 ( .B1(n8626), .B2(n9815), .A(n8011), .ZN(n8012) );
  OAI21_X1 U9598 ( .B1(n8629), .B2(n8604), .A(n8012), .ZN(P2_U3267) );
  NAND2_X1 U9599 ( .A1(n8982), .A2(n4244), .ZN(n8015) );
  NAND2_X1 U9600 ( .A1(n5531), .A2(n8013), .ZN(n8014) );
  NAND2_X1 U9601 ( .A1(n8015), .A2(n8014), .ZN(n8016) );
  XNOR2_X1 U9602 ( .A(n8016), .B(n6362), .ZN(n8020) );
  NOR2_X1 U9603 ( .A1(n9001), .A2(n8017), .ZN(n8018) );
  AOI21_X1 U9604 ( .B1(n8982), .B2(n4247), .A(n8018), .ZN(n8019) );
  XNOR2_X1 U9605 ( .A(n8020), .B(n8019), .ZN(n8027) );
  INV_X1 U9606 ( .A(n8027), .ZN(n8021) );
  NAND2_X1 U9607 ( .A1(n8021), .A2(n8829), .ZN(n8033) );
  NAND4_X1 U9608 ( .A1(n8032), .A2(n8829), .A3(n8026), .A4(n8027), .ZN(n8031)
         );
  OAI22_X1 U9609 ( .A1(n8986), .A2(n8833), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8022), .ZN(n8023) );
  AOI21_X1 U9610 ( .B1(n8843), .B2(n8979), .A(n8023), .ZN(n8024) );
  OAI21_X1 U9611 ( .B1(n8025), .B2(n8848), .A(n8024), .ZN(n8029) );
  NOR3_X1 U9612 ( .A1(n8027), .A2(n8026), .A3(n8853), .ZN(n8028) );
  AOI211_X1 U9613 ( .C1(n8982), .C2(n8850), .A(n8029), .B(n8028), .ZN(n8030)
         );
  OAI211_X1 U9614 ( .C1(n8033), .C2(n8032), .A(n8031), .B(n8030), .ZN(P1_U3218) );
  AOI21_X1 U9615 ( .B1(n8035), .B2(n8034), .A(n8216), .ZN(n8036) );
  NAND2_X1 U9616 ( .A1(n8036), .A2(n8087), .ZN(n8042) );
  AOI22_X1 U9617 ( .A1(n8129), .A2(n8037), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n8041) );
  AOI22_X1 U9618 ( .A1(n8214), .A2(n8039), .B1(n8209), .B2(n8038), .ZN(n8040)
         );
  NAND3_X1 U9619 ( .A1(n8042), .A2(n8041), .A3(n8040), .ZN(P2_U3215) );
  XNOR2_X1 U9620 ( .A(n8044), .B(n8043), .ZN(n8051) );
  OAI22_X1 U9621 ( .A1(n8045), .A2(n8538), .B1(n8111), .B2(n8536), .ZN(n8424)
         );
  INV_X1 U9622 ( .A(n8416), .ZN(n8047) );
  OAI22_X1 U9623 ( .A1(n8047), .A2(n8198), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8046), .ZN(n8048) );
  AOI21_X1 U9624 ( .B1(n8424), .B2(n8129), .A(n8048), .ZN(n8050) );
  NAND2_X1 U9625 ( .A1(n8636), .A2(n8214), .ZN(n8049) );
  OAI211_X1 U9626 ( .C1(n8051), .C2(n8216), .A(n8050), .B(n8049), .ZN(P2_U3216) );
  INV_X1 U9627 ( .A(n8052), .ZN(n8054) );
  NOR2_X1 U9628 ( .A1(n8054), .A2(n8053), .ZN(n8145) );
  INV_X1 U9629 ( .A(n8506), .ZN(n8221) );
  AOI22_X1 U9630 ( .A1(n8052), .A2(n8181), .B1(n8180), .B2(n8221), .ZN(n8059)
         );
  OAI22_X1 U9631 ( .A1(n8198), .A2(n8488), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8055), .ZN(n8057) );
  OAI22_X1 U9632 ( .A1(n8220), .A2(n8199), .B1(n8106), .B2(n8200), .ZN(n8056)
         );
  AOI211_X1 U9633 ( .C1(n8656), .C2(n8214), .A(n8057), .B(n8056), .ZN(n8058)
         );
  OAI21_X1 U9634 ( .B1(n8145), .B2(n8059), .A(n8058), .ZN(P2_U3218) );
  NOR3_X1 U9635 ( .A1(n8194), .A2(n8061), .A3(n8060), .ZN(n8067) );
  INV_X1 U9636 ( .A(n8062), .ZN(n8063) );
  AOI21_X1 U9637 ( .B1(n8064), .B2(n8063), .A(n8216), .ZN(n8066) );
  OAI21_X1 U9638 ( .B1(n8067), .B2(n8066), .A(n8065), .ZN(n8073) );
  INV_X1 U9639 ( .A(n8068), .ZN(n8069) );
  AOI22_X1 U9640 ( .A1(n8214), .A2(n6115), .B1(n8129), .B2(n8069), .ZN(n8072)
         );
  MUX2_X1 U9641 ( .A(P2_STATE_REG_SCAN_IN), .B(n8198), .S(n8070), .Z(n8071) );
  NAND3_X1 U9642 ( .A1(n8073), .A2(n8072), .A3(n8071), .ZN(P2_U3220) );
  INV_X1 U9643 ( .A(n8074), .ZN(n8077) );
  NOR3_X1 U9644 ( .A1(n8075), .A2(n8138), .A3(n8194), .ZN(n8076) );
  AOI21_X1 U9645 ( .B1(n8077), .B2(n8181), .A(n8076), .ZN(n8084) );
  OAI22_X1 U9646 ( .A1(n8101), .A2(n8538), .B1(n8138), .B2(n8536), .ZN(n8557)
         );
  AOI22_X1 U9647 ( .A1(n8129), .A2(n8557), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3152), .ZN(n8078) );
  OAI21_X1 U9648 ( .B1(n8550), .B2(n8198), .A(n8078), .ZN(n8081) );
  NOR2_X1 U9649 ( .A1(n8079), .A2(n8216), .ZN(n8080) );
  AOI211_X1 U9650 ( .C1(n8677), .C2(n8214), .A(n8081), .B(n8080), .ZN(n8082)
         );
  OAI21_X1 U9651 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(P2_U3221) );
  INV_X1 U9652 ( .A(n8085), .ZN(n8086) );
  AOI21_X1 U9653 ( .B1(n8087), .B2(n8086), .A(n8216), .ZN(n8092) );
  NOR3_X1 U9654 ( .A1(n8194), .A2(n8089), .A3(n8088), .ZN(n8091) );
  OAI21_X1 U9655 ( .B1(n8092), .B2(n8091), .A(n8090), .ZN(n8098) );
  AOI22_X1 U9656 ( .A1(n8175), .A2(n8230), .B1(n8174), .B2(n8232), .ZN(n8097)
         );
  AOI22_X1 U9657 ( .A1(n8209), .A2(n8093), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n8096) );
  NAND2_X1 U9658 ( .A1(n8214), .A2(n8094), .ZN(n8095) );
  NAND4_X1 U9659 ( .A1(n8098), .A2(n8097), .A3(n8096), .A4(n8095), .ZN(
        P2_U3223) );
  INV_X1 U9660 ( .A(n8099), .ZN(n8100) );
  AOI21_X1 U9661 ( .B1(n8169), .B2(n8100), .A(n8216), .ZN(n8105) );
  NOR3_X1 U9662 ( .A1(n8102), .A2(n8101), .A3(n8194), .ZN(n8104) );
  OAI21_X1 U9663 ( .B1(n8105), .B2(n8104), .A(n8103), .ZN(n8110) );
  INV_X1 U9664 ( .A(n8106), .ZN(n8480) );
  AOI22_X1 U9665 ( .A1(n8480), .A2(n8572), .B1(n8571), .B2(n8223), .ZN(n8518)
         );
  OAI22_X1 U9666 ( .A1(n8518), .A2(n8212), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8107), .ZN(n8108) );
  AOI21_X1 U9667 ( .B1(n8521), .B2(n8209), .A(n8108), .ZN(n8109) );
  OAI211_X1 U9668 ( .C1(n8524), .C2(n8190), .A(n8110), .B(n8109), .ZN(P2_U3225) );
  INV_X1 U9669 ( .A(n8451), .ZN(n8113) );
  OAI22_X1 U9670 ( .A1(n8111), .A2(n8538), .B1(n8220), .B2(n8536), .ZN(n8457)
         );
  AOI22_X1 U9671 ( .A1(n8457), .A2(n8129), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8112) );
  OAI21_X1 U9672 ( .B1(n8113), .B2(n8198), .A(n8112), .ZN(n8120) );
  NAND3_X1 U9673 ( .A1(n8115), .A2(n8180), .A3(n8472), .ZN(n8116) );
  OAI21_X1 U9674 ( .B1(n8117), .B2(n8216), .A(n8116), .ZN(n8118) );
  AOI211_X1 U9675 ( .C1(n8646), .C2(n8214), .A(n8120), .B(n8119), .ZN(n8121)
         );
  INV_X1 U9676 ( .A(n8121), .ZN(P2_U3227) );
  INV_X1 U9677 ( .A(n8122), .ZN(n8123) );
  AOI21_X1 U9678 ( .B1(n8125), .B2(n8124), .A(n8123), .ZN(n8134) );
  INV_X1 U9679 ( .A(n8594), .ZN(n8131) );
  OR2_X1 U9680 ( .A1(n8126), .A2(n8536), .ZN(n8128) );
  NAND2_X1 U9681 ( .A1(n8570), .A2(n8572), .ZN(n8127) );
  NAND2_X1 U9682 ( .A1(n8128), .A2(n8127), .ZN(n8599) );
  AOI22_X1 U9683 ( .A1(n8129), .A2(n8599), .B1(P2_REG3_REG_16__SCAN_IN), .B2(
        P2_U3152), .ZN(n8130) );
  OAI21_X1 U9684 ( .B1(n8131), .B2(n8198), .A(n8130), .ZN(n8132) );
  AOI21_X1 U9685 ( .B1(n8692), .B2(n8214), .A(n8132), .ZN(n8133) );
  OAI21_X1 U9686 ( .B1(n8134), .B2(n8216), .A(n8133), .ZN(P2_U3228) );
  OAI211_X1 U9687 ( .C1(n4332), .C2(n8136), .A(n8193), .B(n8181), .ZN(n8143)
         );
  OAI22_X1 U9688 ( .A1(n8138), .A2(n8538), .B1(n8137), .B2(n8536), .ZN(n8586)
         );
  INV_X1 U9689 ( .A(n8586), .ZN(n8140) );
  OAI22_X1 U9690 ( .A1(n8212), .A2(n8140), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8139), .ZN(n8141) );
  AOI21_X1 U9691 ( .B1(n8582), .B2(n8209), .A(n8141), .ZN(n8142) );
  OAI211_X1 U9692 ( .C1(n4603), .C2(n8190), .A(n8143), .B(n8142), .ZN(P2_U3230) );
  NOR2_X1 U9693 ( .A1(n8145), .A2(n8144), .ZN(n8147) );
  XNOR2_X1 U9694 ( .A(n8147), .B(n8146), .ZN(n8150) );
  OAI22_X1 U9695 ( .A1(n8150), .A2(n8216), .B1(n8220), .B2(n8194), .ZN(n8148)
         );
  OAI21_X1 U9696 ( .B1(n8150), .B2(n8149), .A(n8148), .ZN(n8156) );
  OAI22_X1 U9697 ( .A1(n8464), .A2(n8198), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8151), .ZN(n8154) );
  OAI22_X1 U9698 ( .A1(n8152), .A2(n8199), .B1(n8506), .B2(n8200), .ZN(n8153)
         );
  AOI211_X1 U9699 ( .C1(n8650), .C2(n8214), .A(n8154), .B(n8153), .ZN(n8155)
         );
  NAND2_X1 U9700 ( .A1(n8156), .A2(n8155), .ZN(P2_U3231) );
  OAI22_X1 U9701 ( .A1(n9877), .A2(n8190), .B1(n8199), .B2(n8157), .ZN(n8158)
         );
  AOI211_X1 U9702 ( .C1(n8160), .C2(n8209), .A(n8159), .B(n8158), .ZN(n8168)
         );
  OAI21_X1 U9703 ( .B1(n8163), .B2(n8065), .A(n8161), .ZN(n8162) );
  NAND2_X1 U9704 ( .A1(n8162), .A2(n8181), .ZN(n8167) );
  NOR3_X1 U9705 ( .A1(n8194), .A2(n8164), .A3(n8163), .ZN(n8165) );
  OAI21_X1 U9706 ( .B1(n8165), .B2(n8174), .A(n8236), .ZN(n8166) );
  NAND3_X1 U9707 ( .A1(n8168), .A2(n8167), .A3(n8166), .ZN(P2_U3232) );
  INV_X1 U9708 ( .A(n8169), .ZN(n8170) );
  AOI211_X1 U9709 ( .C1(n8172), .C2(n8171), .A(n8216), .B(n8170), .ZN(n8179)
         );
  INV_X1 U9710 ( .A(n8671), .ZN(n8532) );
  INV_X1 U9711 ( .A(n8173), .ZN(n8530) );
  AOI22_X1 U9712 ( .A1(n8209), .A2(n8530), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8177) );
  AOI22_X1 U9713 ( .A1(n8175), .A2(n8222), .B1(n8174), .B2(n8573), .ZN(n8176)
         );
  OAI211_X1 U9714 ( .C1(n8532), .C2(n8190), .A(n8177), .B(n8176), .ZN(n8178)
         );
  OR2_X1 U9715 ( .A1(n8179), .A2(n8178), .ZN(P2_U3235) );
  NAND2_X1 U9716 ( .A1(n8480), .A2(n8180), .ZN(n8185) );
  NAND2_X1 U9717 ( .A1(n8182), .A2(n8181), .ZN(n8184) );
  MUX2_X1 U9718 ( .A(n8185), .B(n8184), .S(n8183), .Z(n8189) );
  NOR2_X1 U9719 ( .A1(n8198), .A2(n8500), .ZN(n8187) );
  OAI22_X1 U9720 ( .A1(n8506), .A2(n8199), .B1(n8200), .B2(n8539), .ZN(n8186)
         );
  AOI211_X1 U9721 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8187), 
        .B(n8186), .ZN(n8188) );
  OAI211_X1 U9722 ( .C1(n8503), .C2(n8190), .A(n8189), .B(n8188), .ZN(P2_U3237) );
  INV_X1 U9723 ( .A(n8191), .ZN(n8192) );
  AOI21_X1 U9724 ( .B1(n8193), .B2(n8192), .A(n8216), .ZN(n8197) );
  NOR3_X1 U9725 ( .A1(n8195), .A2(n8201), .A3(n8194), .ZN(n8196) );
  OAI21_X1 U9726 ( .B1(n8197), .B2(n8196), .A(n8074), .ZN(n8205) );
  OAI22_X1 U9727 ( .A1(n8198), .A2(n8564), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8355), .ZN(n8203) );
  OAI22_X1 U9728 ( .A1(n8201), .A2(n8200), .B1(n8199), .B2(n8537), .ZN(n8202)
         );
  AOI211_X1 U9729 ( .C1(n8681), .C2(n8214), .A(n8203), .B(n8202), .ZN(n8204)
         );
  NAND2_X1 U9730 ( .A1(n8205), .A2(n8204), .ZN(P2_U3240) );
  XNOR2_X1 U9731 ( .A(n8207), .B(n8206), .ZN(n8217) );
  AND2_X1 U9732 ( .A1(n8472), .A2(n8571), .ZN(n8208) );
  AOI21_X1 U9733 ( .B1(n8219), .B2(n8572), .A(n8208), .ZN(n8440) );
  INV_X1 U9734 ( .A(n8432), .ZN(n8210) );
  AOI22_X1 U9735 ( .A1(n8210), .A2(n8209), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8211) );
  OAI21_X1 U9736 ( .B1(n8440), .B2(n8212), .A(n8211), .ZN(n8213) );
  AOI21_X1 U9737 ( .B1(n8642), .B2(n8214), .A(n8213), .ZN(n8215) );
  OAI21_X1 U9738 ( .B1(n8217), .B2(n8216), .A(n8215), .ZN(P2_U3242) );
  MUX2_X1 U9739 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8218), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9740 ( .A(n4471), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8238), .Z(
        P2_U3580) );
  MUX2_X1 U9741 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8219), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U9742 ( .A(n8472), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8238), .Z(
        P2_U3577) );
  MUX2_X1 U9743 ( .A(n7996), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8238), .Z(
        P2_U3576) );
  MUX2_X1 U9744 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8221), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U9745 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8480), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U9746 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8222), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U9747 ( .A(n8223), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8238), .Z(
        P2_U3572) );
  MUX2_X1 U9748 ( .A(n8573), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8238), .Z(
        P2_U3571) );
  MUX2_X1 U9749 ( .A(n8224), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8238), .Z(
        P2_U3570) );
  MUX2_X1 U9750 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8570), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U9751 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n4668), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U9752 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8225), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9753 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8226), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9754 ( .A(n8227), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8238), .Z(
        P2_U3564) );
  MUX2_X1 U9755 ( .A(n8228), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8238), .Z(
        P2_U3563) );
  MUX2_X1 U9756 ( .A(n8229), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8238), .Z(
        P2_U3562) );
  MUX2_X1 U9757 ( .A(n8230), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8238), .Z(
        P2_U3561) );
  MUX2_X1 U9758 ( .A(n8231), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8238), .Z(
        P2_U3560) );
  MUX2_X1 U9759 ( .A(n8232), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8238), .Z(
        P2_U3559) );
  MUX2_X1 U9760 ( .A(n8233), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8238), .Z(
        P2_U3558) );
  MUX2_X1 U9761 ( .A(n8234), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8238), .Z(
        P2_U3557) );
  MUX2_X1 U9762 ( .A(n8235), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8238), .Z(
        P2_U3556) );
  MUX2_X1 U9763 ( .A(n8236), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8238), .Z(
        P2_U3555) );
  MUX2_X1 U9764 ( .A(n8237), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8238), .Z(
        P2_U3554) );
  MUX2_X1 U9765 ( .A(n6830), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8238), .Z(
        P2_U3553) );
  OAI211_X1 U9766 ( .C1(n8241), .C2(n8240), .A(n9784), .B(n8239), .ZN(n8252)
         );
  NOR2_X1 U9767 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8242), .ZN(n8243) );
  AOI21_X1 U9768 ( .B1(n9793), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8243), .ZN(
        n8251) );
  NAND2_X1 U9769 ( .A1(n9454), .A2(n8244), .ZN(n8250) );
  AOI21_X1 U9770 ( .B1(n8247), .B2(n8246), .A(n8245), .ZN(n8248) );
  NAND2_X1 U9771 ( .A1(n9787), .A2(n8248), .ZN(n8249) );
  NAND4_X1 U9772 ( .A1(n8252), .A2(n8251), .A3(n8250), .A4(n8249), .ZN(
        P2_U3250) );
  OAI211_X1 U9773 ( .C1(n8255), .C2(n8254), .A(n9784), .B(n8253), .ZN(n8266)
         );
  INV_X1 U9774 ( .A(n8256), .ZN(n8257) );
  AOI21_X1 U9775 ( .B1(n9793), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8257), .ZN(
        n8265) );
  NAND2_X1 U9776 ( .A1(n9454), .A2(n8258), .ZN(n8264) );
  AOI21_X1 U9777 ( .B1(n8261), .B2(n8260), .A(n8259), .ZN(n8262) );
  NAND2_X1 U9778 ( .A1(n9787), .A2(n8262), .ZN(n8263) );
  NAND4_X1 U9779 ( .A1(n8266), .A2(n8265), .A3(n8264), .A4(n8263), .ZN(
        P2_U3251) );
  OAI211_X1 U9780 ( .C1(n8269), .C2(n8268), .A(n9784), .B(n8267), .ZN(n8279)
         );
  AND2_X1 U9781 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8270) );
  AOI21_X1 U9782 ( .B1(n9793), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8270), .ZN(
        n8278) );
  NAND2_X1 U9783 ( .A1(n9454), .A2(n8271), .ZN(n8277) );
  AOI21_X1 U9784 ( .B1(n8274), .B2(n8273), .A(n8272), .ZN(n8275) );
  NAND2_X1 U9785 ( .A1(n9787), .A2(n8275), .ZN(n8276) );
  NAND4_X1 U9786 ( .A1(n8279), .A2(n8278), .A3(n8277), .A4(n8276), .ZN(
        P2_U3252) );
  OAI211_X1 U9787 ( .C1(n8282), .C2(n8281), .A(n9784), .B(n8280), .ZN(n8292)
         );
  NOR2_X1 U9788 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9342), .ZN(n8283) );
  AOI21_X1 U9789 ( .B1(n9793), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8283), .ZN(
        n8291) );
  NAND2_X1 U9790 ( .A1(n9454), .A2(n8284), .ZN(n8290) );
  AOI21_X1 U9791 ( .B1(n8287), .B2(n8286), .A(n8285), .ZN(n8288) );
  NAND2_X1 U9792 ( .A1(n9787), .A2(n8288), .ZN(n8289) );
  NAND4_X1 U9793 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(
        P2_U3253) );
  OAI211_X1 U9794 ( .C1(n8295), .C2(n8294), .A(n9784), .B(n8293), .ZN(n8305)
         );
  NOR2_X1 U9795 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5735), .ZN(n8296) );
  AOI21_X1 U9796 ( .B1(n9793), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8296), .ZN(
        n8304) );
  NAND2_X1 U9797 ( .A1(n9454), .A2(n8297), .ZN(n8303) );
  AOI21_X1 U9798 ( .B1(n8300), .B2(n8299), .A(n8298), .ZN(n8301) );
  NAND2_X1 U9799 ( .A1(n9787), .A2(n8301), .ZN(n8302) );
  NAND4_X1 U9800 ( .A1(n8305), .A2(n8304), .A3(n8303), .A4(n8302), .ZN(
        P2_U3254) );
  NOR2_X1 U9801 ( .A1(n8312), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8307) );
  NOR2_X1 U9802 ( .A1(n8307), .A2(n8306), .ZN(n8325) );
  XNOR2_X1 U9803 ( .A(n8325), .B(n8326), .ZN(n8308) );
  NOR2_X1 U9804 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8308), .ZN(n8327) );
  AOI21_X1 U9805 ( .B1(n8308), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8327), .ZN(
        n8317) );
  INV_X1 U9806 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U9807 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8309) );
  OAI21_X1 U9808 ( .B1(n9437), .B2(n8310), .A(n8309), .ZN(n8315) );
  INV_X1 U9809 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n9466) );
  AOI211_X1 U9810 ( .C1(n8313), .C2(n9466), .A(n8320), .B(n9448), .ZN(n8314)
         );
  AOI211_X1 U9811 ( .C1(n9454), .C2(n8326), .A(n8315), .B(n8314), .ZN(n8316)
         );
  OAI21_X1 U9812 ( .B1(n8317), .B2(n8373), .A(n8316), .ZN(P2_U3260) );
  NOR2_X1 U9813 ( .A1(n8319), .A2(n8318), .ZN(n8321) );
  NOR2_X1 U9814 ( .A1(n8321), .A2(n8320), .ZN(n8334) );
  XNOR2_X1 U9815 ( .A(n8335), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8336) );
  XNOR2_X1 U9816 ( .A(n8334), .B(n8336), .ZN(n8333) );
  NOR2_X1 U9817 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8322), .ZN(n8324) );
  NOR2_X1 U9818 ( .A1(n9789), .A2(n8341), .ZN(n8323) );
  AOI211_X1 U9819 ( .C1(n9793), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8324), .B(
        n8323), .ZN(n8332) );
  NOR2_X1 U9820 ( .A1(n8326), .A2(n8325), .ZN(n8328) );
  NOR2_X1 U9821 ( .A1(n8328), .A2(n8327), .ZN(n8330) );
  INV_X1 U9822 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8342) );
  MUX2_X1 U9823 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n8342), .S(n8335), .Z(n8329)
         );
  NAND2_X1 U9824 ( .A1(n8330), .A2(n8329), .ZN(n8340) );
  OAI211_X1 U9825 ( .C1(n8330), .C2(n8329), .A(n8340), .B(n9784), .ZN(n8331)
         );
  OAI211_X1 U9826 ( .C1(n8333), .C2(n9448), .A(n8332), .B(n8331), .ZN(P2_U3261) );
  XNOR2_X1 U9827 ( .A(n8357), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8339) );
  INV_X1 U9828 ( .A(n8334), .ZN(n8337) );
  OAI22_X1 U9829 ( .A1(n8337), .A2(n8336), .B1(n8335), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n8338) );
  NOR2_X1 U9830 ( .A1(n8338), .A2(n8339), .ZN(n8351) );
  AOI211_X1 U9831 ( .C1(n8339), .C2(n8338), .A(n9448), .B(n8351), .ZN(n8350)
         );
  OAI21_X1 U9832 ( .B1(n8342), .B2(n8341), .A(n8340), .ZN(n8344) );
  XOR2_X1 U9833 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n8357), .Z(n8343) );
  NAND2_X1 U9834 ( .A1(n8343), .A2(n8344), .ZN(n8358) );
  OAI211_X1 U9835 ( .C1(n8344), .C2(n8343), .A(n9784), .B(n8358), .ZN(n8347)
         );
  NOR2_X1 U9836 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8139), .ZN(n8345) );
  AOI21_X1 U9837 ( .B1(n9793), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8345), .ZN(
        n8346) );
  OAI211_X1 U9838 ( .C1(n9789), .C2(n8348), .A(n8347), .B(n8346), .ZN(n8349)
         );
  OR2_X1 U9839 ( .A1(n8350), .A2(n8349), .ZN(P2_U3262) );
  XNOR2_X1 U9840 ( .A(n8360), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8352) );
  OAI21_X1 U9841 ( .B1(n8353), .B2(n8352), .A(n8370), .ZN(n8354) );
  NAND2_X1 U9842 ( .A1(n8354), .A2(n9787), .ZN(n8365) );
  NOR2_X1 U9843 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8355), .ZN(n8356) );
  AOI21_X1 U9844 ( .B1(n9793), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8356), .ZN(
        n8364) );
  NAND2_X1 U9845 ( .A1(n8357), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8359) );
  NAND2_X1 U9846 ( .A1(n8359), .A2(n8358), .ZN(n8366) );
  XNOR2_X1 U9847 ( .A(n8366), .B(n8360), .ZN(n8361) );
  NAND2_X1 U9848 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8361), .ZN(n8368) );
  OAI211_X1 U9849 ( .C1(n8361), .C2(P2_REG2_REG_18__SCAN_IN), .A(n9784), .B(
        n8368), .ZN(n8363) );
  NAND2_X1 U9850 ( .A1(n9454), .A2(n8371), .ZN(n8362) );
  NAND4_X1 U9851 ( .A1(n8365), .A2(n8364), .A3(n8363), .A4(n8362), .ZN(
        P2_U3263) );
  NAND2_X1 U9852 ( .A1(n8371), .A2(n8366), .ZN(n8367) );
  NAND2_X1 U9853 ( .A1(n8368), .A2(n8367), .ZN(n8369) );
  XOR2_X1 U9854 ( .A(n8369), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8374) );
  AOI22_X1 U9855 ( .A1(n8374), .A2(n9784), .B1(n9787), .B2(n8372), .ZN(n8379)
         );
  INV_X1 U9856 ( .A(n8372), .ZN(n8376) );
  NOR2_X1 U9857 ( .A1(n8374), .A2(n8373), .ZN(n8375) );
  AOI211_X1 U9858 ( .C1(n9787), .C2(n8376), .A(n9454), .B(n8375), .ZN(n8378)
         );
  MUX2_X1 U9859 ( .A(n8379), .B(n8378), .S(n8377), .Z(n8381) );
  NAND2_X1 U9860 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8380) );
  OAI211_X1 U9861 ( .C1(n4349), .C2(n9437), .A(n8381), .B(n8380), .ZN(P2_U3264) );
  NAND2_X1 U9862 ( .A1(n8625), .A2(n8388), .ZN(n8621) );
  XNOR2_X1 U9863 ( .A(n8621), .B(n8618), .ZN(n8620) );
  NAND2_X1 U9864 ( .A1(n8383), .A2(n8382), .ZN(n8623) );
  NOR2_X1 U9865 ( .A1(n9840), .A2(n8623), .ZN(n8391) );
  NOR2_X1 U9866 ( .A1(n8384), .A2(n9817), .ZN(n8385) );
  AOI211_X1 U9867 ( .C1(n9840), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8391), .B(
        n8385), .ZN(n8386) );
  OAI21_X1 U9868 ( .B1(n8620), .B2(n8387), .A(n8386), .ZN(P2_U3265) );
  INV_X1 U9869 ( .A(n8388), .ZN(n8389) );
  NAND2_X1 U9870 ( .A1(n8390), .A2(n8389), .ZN(n8622) );
  NAND3_X1 U9871 ( .A1(n8622), .A2(n9845), .A3(n8621), .ZN(n8393) );
  AOI21_X1 U9872 ( .B1(n8495), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8391), .ZN(
        n8392) );
  OAI211_X1 U9873 ( .C1(n8625), .C2(n9817), .A(n8393), .B(n8392), .ZN(P2_U3266) );
  XNOR2_X1 U9874 ( .A(n8395), .B(n8394), .ZN(n8634) );
  INV_X1 U9875 ( .A(n8396), .ZN(n8397) );
  AOI21_X1 U9876 ( .B1(n8630), .B2(n8414), .A(n8397), .ZN(n8631) );
  INV_X1 U9877 ( .A(n8398), .ZN(n8399) );
  AOI22_X1 U9878 ( .A1(n8399), .A2(n9839), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8495), .ZN(n8400) );
  OAI21_X1 U9879 ( .B1(n8401), .B2(n9817), .A(n8400), .ZN(n8411) );
  INV_X1 U9880 ( .A(n8402), .ZN(n8404) );
  AOI21_X1 U9881 ( .B1(n8404), .B2(n8403), .A(n8533), .ZN(n8409) );
  OAI22_X1 U9882 ( .A1(n8406), .A2(n8536), .B1(n8405), .B2(n8538), .ZN(n8407)
         );
  AOI21_X1 U9883 ( .B1(n8409), .B2(n8408), .A(n8407), .ZN(n8633) );
  NOR2_X1 U9884 ( .A1(n8633), .A2(n9840), .ZN(n8410) );
  AOI211_X1 U9885 ( .C1(n8631), .C2(n9845), .A(n8411), .B(n8410), .ZN(n8412)
         );
  OAI21_X1 U9886 ( .B1(n8634), .B2(n8604), .A(n8412), .ZN(P2_U3268) );
  XOR2_X1 U9887 ( .A(n8422), .B(n8413), .Z(n8639) );
  INV_X1 U9888 ( .A(n8414), .ZN(n8415) );
  AOI211_X1 U9889 ( .C1(n8636), .C2(n8430), .A(n9921), .B(n8415), .ZN(n8635)
         );
  INV_X1 U9890 ( .A(n8636), .ZN(n8418) );
  AOI22_X1 U9891 ( .A1(n8416), .A2(n9839), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8495), .ZN(n8417) );
  OAI21_X1 U9892 ( .B1(n8418), .B2(n9817), .A(n8417), .ZN(n8427) );
  INV_X1 U9893 ( .A(n8419), .ZN(n8437) );
  OAI21_X1 U9894 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8423) );
  AOI211_X1 U9895 ( .C1(n8437), .C2(n4751), .A(n8533), .B(n8423), .ZN(n8425)
         );
  NOR2_X1 U9896 ( .A1(n8425), .A2(n8424), .ZN(n8638) );
  NOR2_X1 U9897 ( .A1(n8638), .A2(n8495), .ZN(n8426) );
  AOI211_X1 U9898 ( .C1(n9811), .C2(n8635), .A(n8427), .B(n8426), .ZN(n8428)
         );
  OAI21_X1 U9899 ( .B1(n8639), .B2(n8604), .A(n8428), .ZN(P2_U3269) );
  XOR2_X1 U9900 ( .A(n8439), .B(n8429), .Z(n8644) );
  INV_X1 U9901 ( .A(n8430), .ZN(n8431) );
  AOI211_X1 U9902 ( .C1(n8642), .C2(n4612), .A(n9921), .B(n8431), .ZN(n8641)
         );
  OAI22_X1 U9903 ( .A1(n8434), .A2(n8433), .B1(n9814), .B2(n8432), .ZN(n8442)
         );
  INV_X1 U9904 ( .A(n8435), .ZN(n8436) );
  NAND2_X1 U9905 ( .A1(n8458), .A2(n8436), .ZN(n8438) );
  AOI21_X1 U9906 ( .B1(n8439), .B2(n8438), .A(n8437), .ZN(n8441) );
  OAI21_X1 U9907 ( .B1(n8441), .B2(n8533), .A(n8440), .ZN(n8640) );
  AOI211_X1 U9908 ( .C1(n8641), .C2(n8443), .A(n8442), .B(n8640), .ZN(n8444)
         );
  NOR2_X1 U9909 ( .A1(n8444), .A2(n8495), .ZN(n8445) );
  AOI21_X1 U9910 ( .B1(n8495), .B2(P2_REG2_REG_26__SCAN_IN), .A(n8445), .ZN(
        n8446) );
  OAI21_X1 U9911 ( .B1(n8644), .B2(n8604), .A(n8446), .ZN(P2_U3270) );
  XNOR2_X1 U9912 ( .A(n8448), .B(n8455), .ZN(n8649) );
  AOI211_X1 U9913 ( .C1(n8646), .C2(n8450), .A(n9921), .B(n8449), .ZN(n8645)
         );
  AOI22_X1 U9914 ( .A1(n8451), .A2(n9839), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8495), .ZN(n8452) );
  OAI21_X1 U9915 ( .B1(n8453), .B2(n9817), .A(n8452), .ZN(n8461) );
  INV_X1 U9916 ( .A(n8454), .ZN(n8456) );
  AOI21_X1 U9917 ( .B1(n8456), .B2(n8455), .A(n8533), .ZN(n8459) );
  AOI21_X1 U9918 ( .B1(n8459), .B2(n8458), .A(n8457), .ZN(n8648) );
  NOR2_X1 U9919 ( .A1(n8648), .A2(n8495), .ZN(n8460) );
  AOI211_X1 U9920 ( .C1(n8645), .C2(n9811), .A(n8461), .B(n8460), .ZN(n8462)
         );
  OAI21_X1 U9921 ( .B1(n8649), .B2(n8604), .A(n8462), .ZN(P2_U3271) );
  AOI21_X1 U9922 ( .B1(n8469), .B2(n8463), .A(n4318), .ZN(n8654) );
  XNOR2_X1 U9923 ( .A(n8467), .B(n8485), .ZN(n8651) );
  INV_X1 U9924 ( .A(n8464), .ZN(n8465) );
  AOI22_X1 U9925 ( .A1(n8465), .A2(n9839), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n8495), .ZN(n8466) );
  OAI21_X1 U9926 ( .B1(n8467), .B2(n9817), .A(n8466), .ZN(n8476) );
  OAI211_X1 U9927 ( .C1(n8470), .C2(n8469), .A(n8468), .B(n9830), .ZN(n8474)
         );
  NOR2_X1 U9928 ( .A1(n8506), .A2(n8536), .ZN(n8471) );
  AOI21_X1 U9929 ( .B1(n8472), .B2(n8572), .A(n8471), .ZN(n8473) );
  AND2_X1 U9930 ( .A1(n8474), .A2(n8473), .ZN(n8653) );
  NOR2_X1 U9931 ( .A1(n8653), .A2(n9840), .ZN(n8475) );
  AOI211_X1 U9932 ( .C1(n8651), .C2(n9845), .A(n8476), .B(n8475), .ZN(n8477)
         );
  OAI21_X1 U9933 ( .B1(n8654), .B2(n8604), .A(n8477), .ZN(P2_U3272) );
  OAI21_X1 U9934 ( .B1(n8479), .B2(n4319), .A(n8478), .ZN(n8481) );
  AOI222_X1 U9935 ( .A1(n9830), .A2(n8481), .B1(n8480), .B2(n8571), .C1(n7996), 
        .C2(n8572), .ZN(n8659) );
  OR2_X1 U9936 ( .A1(n8483), .A2(n8482), .ZN(n8655) );
  NAND3_X1 U9937 ( .A1(n8655), .A2(n8484), .A3(n9838), .ZN(n8494) );
  INV_X1 U9938 ( .A(n8498), .ZN(n8487) );
  INV_X1 U9939 ( .A(n8485), .ZN(n8486) );
  AOI21_X1 U9940 ( .B1(n8656), .B2(n8487), .A(n8486), .ZN(n8657) );
  INV_X1 U9941 ( .A(n8488), .ZN(n8489) );
  AOI22_X1 U9942 ( .A1(n8489), .A2(n9839), .B1(P2_REG2_REG_23__SCAN_IN), .B2(
        n8495), .ZN(n8490) );
  OAI21_X1 U9943 ( .B1(n8491), .B2(n9817), .A(n8490), .ZN(n8492) );
  AOI21_X1 U9944 ( .B1(n8657), .B2(n9845), .A(n8492), .ZN(n8493) );
  OAI211_X1 U9945 ( .C1(n8495), .C2(n8659), .A(n8494), .B(n8493), .ZN(P2_U3273) );
  XOR2_X1 U9946 ( .A(n8496), .B(n8504), .Z(n8665) );
  INV_X1 U9947 ( .A(n8497), .ZN(n8499) );
  AOI21_X1 U9948 ( .B1(n8661), .B2(n8499), .A(n8498), .ZN(n8662) );
  INV_X1 U9949 ( .A(n8500), .ZN(n8501) );
  AOI22_X1 U9950 ( .A1(n8501), .A2(n9839), .B1(n8495), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n8502) );
  OAI21_X1 U9951 ( .B1(n8503), .B2(n9817), .A(n8502), .ZN(n8511) );
  AOI21_X1 U9952 ( .B1(n8505), .B2(n8504), .A(n8533), .ZN(n8509) );
  OAI22_X1 U9953 ( .A1(n8506), .A2(n8538), .B1(n8539), .B2(n8536), .ZN(n8507)
         );
  AOI21_X1 U9954 ( .B1(n8509), .B2(n8508), .A(n8507), .ZN(n8664) );
  NOR2_X1 U9955 ( .A1(n8664), .A2(n8495), .ZN(n8510) );
  AOI211_X1 U9956 ( .C1(n8662), .C2(n9845), .A(n8511), .B(n8510), .ZN(n8512)
         );
  OAI21_X1 U9957 ( .B1(n8665), .B2(n8604), .A(n8512), .ZN(P2_U3274) );
  XOR2_X1 U9958 ( .A(n8513), .B(n8517), .Z(n8670) );
  NAND2_X1 U9959 ( .A1(n8514), .A2(n8515), .ZN(n8516) );
  XOR2_X1 U9960 ( .A(n8517), .B(n8516), .Z(n8519) );
  OAI21_X1 U9961 ( .B1(n8519), .B2(n8533), .A(n8518), .ZN(n8666) );
  XNOR2_X1 U9962 ( .A(n8668), .B(n8528), .ZN(n8520) );
  NOR2_X1 U9963 ( .A1(n8520), .A2(n9921), .ZN(n8667) );
  NAND2_X1 U9964 ( .A1(n8667), .A2(n9811), .ZN(n8523) );
  AOI22_X1 U9965 ( .A1(n8495), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8521), .B2(
        n9839), .ZN(n8522) );
  OAI211_X1 U9966 ( .C1(n8524), .C2(n9817), .A(n8523), .B(n8522), .ZN(n8525)
         );
  AOI21_X1 U9967 ( .B1(n8666), .B2(n9815), .A(n8525), .ZN(n8526) );
  OAI21_X1 U9968 ( .B1(n8670), .B2(n8604), .A(n8526), .ZN(P2_U3275) );
  XNOR2_X1 U9969 ( .A(n8527), .B(n8534), .ZN(n8675) );
  INV_X1 U9970 ( .A(n8528), .ZN(n8529) );
  AOI21_X1 U9971 ( .B1(n8671), .B2(n8547), .A(n8529), .ZN(n8672) );
  AOI22_X1 U9972 ( .A1(n9840), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8530), .B2(
        n9839), .ZN(n8531) );
  OAI21_X1 U9973 ( .B1(n8532), .B2(n9817), .A(n8531), .ZN(n8543) );
  AOI21_X1 U9974 ( .B1(n8535), .B2(n8534), .A(n8533), .ZN(n8541) );
  OAI22_X1 U9975 ( .A1(n8539), .A2(n8538), .B1(n8537), .B2(n8536), .ZN(n8540)
         );
  AOI21_X1 U9976 ( .B1(n8541), .B2(n8514), .A(n8540), .ZN(n8674) );
  NOR2_X1 U9977 ( .A1(n8674), .A2(n9840), .ZN(n8542) );
  AOI211_X1 U9978 ( .C1(n8672), .C2(n9845), .A(n8543), .B(n8542), .ZN(n8544)
         );
  OAI21_X1 U9979 ( .B1(n8675), .B2(n8604), .A(n8544), .ZN(P2_U3276) );
  XNOR2_X1 U9980 ( .A(n8545), .B(n8546), .ZN(n8680) );
  INV_X1 U9981 ( .A(n8563), .ZN(n8549) );
  INV_X1 U9982 ( .A(n8547), .ZN(n8548) );
  AOI211_X1 U9983 ( .C1(n8677), .C2(n8549), .A(n9921), .B(n8548), .ZN(n8676)
         );
  INV_X1 U9984 ( .A(n8550), .ZN(n8551) );
  AOI22_X1 U9985 ( .A1(n8495), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8551), .B2(
        n9839), .ZN(n8552) );
  OAI21_X1 U9986 ( .B1(n8553), .B2(n9817), .A(n8552), .ZN(n8560) );
  NAND2_X1 U9987 ( .A1(n8567), .A2(n8554), .ZN(n8556) );
  XNOR2_X1 U9988 ( .A(n8556), .B(n8555), .ZN(n8558) );
  AOI21_X1 U9989 ( .B1(n8558), .B2(n9830), .A(n8557), .ZN(n8679) );
  NOR2_X1 U9990 ( .A1(n8679), .A2(n9840), .ZN(n8559) );
  AOI211_X1 U9991 ( .C1(n8676), .C2(n9811), .A(n8560), .B(n8559), .ZN(n8561)
         );
  OAI21_X1 U9992 ( .B1(n8680), .B2(n8604), .A(n8561), .ZN(P2_U3277) );
  XOR2_X1 U9993 ( .A(n8569), .B(n8562), .Z(n8685) );
  AOI21_X1 U9994 ( .B1(n8681), .B2(n8581), .A(n8563), .ZN(n8682) );
  INV_X1 U9995 ( .A(n8564), .ZN(n8565) );
  AOI22_X1 U9996 ( .A1(n9840), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8565), .B2(
        n9839), .ZN(n8566) );
  OAI21_X1 U9997 ( .B1(n4604), .B2(n9817), .A(n8566), .ZN(n8577) );
  OAI211_X1 U9998 ( .C1(n8569), .C2(n8568), .A(n8567), .B(n9830), .ZN(n8575)
         );
  AOI22_X1 U9999 ( .A1(n8573), .A2(n8572), .B1(n8571), .B2(n8570), .ZN(n8574)
         );
  AND2_X1 U10000 ( .A1(n8575), .A2(n8574), .ZN(n8684) );
  NOR2_X1 U10001 ( .A1(n8684), .A2(n9840), .ZN(n8576) );
  AOI211_X1 U10002 ( .C1(n8682), .C2(n9845), .A(n8577), .B(n8576), .ZN(n8578)
         );
  OAI21_X1 U10003 ( .B1(n8685), .B2(n8604), .A(n8578), .ZN(P2_U3278) );
  AOI21_X1 U10004 ( .B1(n8584), .B2(n8580), .A(n8579), .ZN(n8690) );
  AOI211_X1 U10005 ( .C1(n8687), .C2(n8593), .A(n9921), .B(n4605), .ZN(n8686)
         );
  AOI22_X1 U10006 ( .A1(n9840), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8582), .B2(
        n9839), .ZN(n8583) );
  OAI21_X1 U10007 ( .B1(n4603), .B2(n9817), .A(n8583), .ZN(n8589) );
  XNOR2_X1 U10008 ( .A(n8585), .B(n8584), .ZN(n8587) );
  AOI21_X1 U10009 ( .B1(n8587), .B2(n9830), .A(n8586), .ZN(n8689) );
  NOR2_X1 U10010 ( .A1(n8689), .A2(n9840), .ZN(n8588) );
  AOI211_X1 U10011 ( .C1(n8686), .C2(n9811), .A(n8589), .B(n8588), .ZN(n8590)
         );
  OAI21_X1 U10012 ( .B1(n8690), .B2(n8604), .A(n8590), .ZN(P2_U3279) );
  OAI21_X1 U10013 ( .B1(n8592), .B2(n8597), .A(n8591), .ZN(n8695) );
  AOI211_X1 U10014 ( .C1(n8692), .C2(n8610), .A(n9921), .B(n4600), .ZN(n8691)
         );
  AOI22_X1 U10015 ( .A1(n9840), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8594), .B2(
        n9839), .ZN(n8595) );
  OAI21_X1 U10016 ( .B1(n8596), .B2(n9817), .A(n8595), .ZN(n8602) );
  XOR2_X1 U10017 ( .A(n8598), .B(n8597), .Z(n8600) );
  AOI21_X1 U10018 ( .B1(n8600), .B2(n9830), .A(n8599), .ZN(n8694) );
  NOR2_X1 U10019 ( .A1(n8694), .A2(n9840), .ZN(n8601) );
  AOI211_X1 U10020 ( .C1(n8691), .C2(n9811), .A(n8602), .B(n8601), .ZN(n8603)
         );
  OAI21_X1 U10021 ( .B1(n8695), .B2(n8604), .A(n8603), .ZN(P2_U3280) );
  XNOR2_X1 U10022 ( .A(n8605), .B(n8608), .ZN(n8607) );
  AOI21_X1 U10023 ( .B1(n8607), .B2(n9830), .A(n8606), .ZN(n9462) );
  XNOR2_X1 U10024 ( .A(n8609), .B(n8608), .ZN(n9465) );
  NAND2_X1 U10025 ( .A1(n9465), .A2(n9838), .ZN(n8617) );
  OAI211_X1 U10026 ( .C1(n8611), .C2(n9463), .A(n4341), .B(n8610), .ZN(n9461)
         );
  INV_X1 U10027 ( .A(n9461), .ZN(n8615) );
  AOI22_X1 U10028 ( .A1(n9840), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8612), .B2(
        n9839), .ZN(n8613) );
  OAI21_X1 U10029 ( .B1(n9463), .B2(n9817), .A(n8613), .ZN(n8614) );
  AOI21_X1 U10030 ( .B1(n8615), .B2(n9811), .A(n8614), .ZN(n8616) );
  OAI211_X1 U10031 ( .C1(n8495), .C2(n9462), .A(n8617), .B(n8616), .ZN(
        P2_U3281) );
  NAND2_X1 U10032 ( .A1(n8618), .A2(n9927), .ZN(n8619) );
  OAI211_X1 U10033 ( .C1(n8620), .C2(n9921), .A(n8619), .B(n8623), .ZN(n8696)
         );
  INV_X2 U10034 ( .A(n9950), .ZN(n9952) );
  MUX2_X1 U10035 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8696), .S(n9952), .Z(
        P2_U3551) );
  INV_X1 U10036 ( .A(n9927), .ZN(n9919) );
  NAND3_X1 U10037 ( .A1(n8622), .A2(n4341), .A3(n8621), .ZN(n8624) );
  OAI211_X1 U10038 ( .C1(n8625), .C2(n9919), .A(n8624), .B(n8623), .ZN(n8697)
         );
  MUX2_X1 U10039 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8697), .S(n9952), .Z(
        P2_U3550) );
  MUX2_X1 U10040 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8698), .S(n9952), .Z(
        P2_U3549) );
  AOI22_X1 U10041 ( .A1(n8631), .A2(n4341), .B1(n9927), .B2(n8630), .ZN(n8632)
         );
  OAI211_X1 U10042 ( .C1(n8634), .C2(n9888), .A(n8633), .B(n8632), .ZN(n8699)
         );
  MUX2_X1 U10043 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8699), .S(n9952), .Z(
        P2_U3548) );
  AOI21_X1 U10044 ( .B1(n9927), .B2(n8636), .A(n8635), .ZN(n8637) );
  OAI211_X1 U10045 ( .C1(n8639), .C2(n9888), .A(n8638), .B(n8637), .ZN(n8700)
         );
  MUX2_X1 U10046 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8700), .S(n9952), .Z(
        P2_U3547) );
  AOI211_X1 U10047 ( .C1(n9927), .C2(n8642), .A(n8641), .B(n8640), .ZN(n8643)
         );
  OAI21_X1 U10048 ( .B1(n8644), .B2(n9888), .A(n8643), .ZN(n8701) );
  MUX2_X1 U10049 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8701), .S(n9952), .Z(
        P2_U3546) );
  AOI21_X1 U10050 ( .B1(n9927), .B2(n8646), .A(n8645), .ZN(n8647) );
  OAI211_X1 U10051 ( .C1(n8649), .C2(n9888), .A(n8648), .B(n8647), .ZN(n8702)
         );
  MUX2_X1 U10052 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8702), .S(n9952), .Z(
        P2_U3545) );
  AOI22_X1 U10053 ( .A1(n8651), .A2(n4341), .B1(n9927), .B2(n8650), .ZN(n8652)
         );
  OAI211_X1 U10054 ( .C1(n8654), .C2(n9888), .A(n8653), .B(n8652), .ZN(n8703)
         );
  MUX2_X1 U10055 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8703), .S(n9952), .Z(
        P2_U3544) );
  INV_X1 U10056 ( .A(n9888), .ZN(n9933) );
  NAND3_X1 U10057 ( .A1(n8655), .A2(n8484), .A3(n9933), .ZN(n8660) );
  AOI22_X1 U10058 ( .A1(n8657), .A2(n4341), .B1(n9927), .B2(n8656), .ZN(n8658)
         );
  NAND3_X1 U10059 ( .A1(n8660), .A2(n8659), .A3(n8658), .ZN(n8704) );
  MUX2_X1 U10060 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8704), .S(n9952), .Z(
        P2_U3543) );
  AOI22_X1 U10061 ( .A1(n8662), .A2(n4341), .B1(n9927), .B2(n8661), .ZN(n8663)
         );
  OAI211_X1 U10062 ( .C1(n8665), .C2(n9888), .A(n8664), .B(n8663), .ZN(n8705)
         );
  MUX2_X1 U10063 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8705), .S(n9952), .Z(
        P2_U3542) );
  AOI211_X1 U10064 ( .C1(n9927), .C2(n8668), .A(n8667), .B(n8666), .ZN(n8669)
         );
  OAI21_X1 U10065 ( .B1(n8670), .B2(n9888), .A(n8669), .ZN(n8706) );
  MUX2_X1 U10066 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8706), .S(n9952), .Z(
        P2_U3541) );
  AOI22_X1 U10067 ( .A1(n8672), .A2(n4341), .B1(n9927), .B2(n8671), .ZN(n8673)
         );
  OAI211_X1 U10068 ( .C1(n8675), .C2(n9888), .A(n8674), .B(n8673), .ZN(n8707)
         );
  MUX2_X1 U10069 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8707), .S(n9952), .Z(
        P2_U3540) );
  AOI21_X1 U10070 ( .B1(n9927), .B2(n8677), .A(n8676), .ZN(n8678) );
  OAI211_X1 U10071 ( .C1(n8680), .C2(n9888), .A(n8679), .B(n8678), .ZN(n8708)
         );
  MUX2_X1 U10072 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8708), .S(n9952), .Z(
        P2_U3539) );
  AOI22_X1 U10073 ( .A1(n8682), .A2(n4341), .B1(n9927), .B2(n8681), .ZN(n8683)
         );
  OAI211_X1 U10074 ( .C1(n8685), .C2(n9888), .A(n8684), .B(n8683), .ZN(n8709)
         );
  MUX2_X1 U10075 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8709), .S(n9952), .Z(
        P2_U3538) );
  AOI21_X1 U10076 ( .B1(n9927), .B2(n8687), .A(n8686), .ZN(n8688) );
  OAI211_X1 U10077 ( .C1(n8690), .C2(n9888), .A(n8689), .B(n8688), .ZN(n8710)
         );
  MUX2_X1 U10078 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8710), .S(n9952), .Z(
        P2_U3537) );
  AOI21_X1 U10079 ( .B1(n9927), .B2(n8692), .A(n8691), .ZN(n8693) );
  OAI211_X1 U10080 ( .C1(n8695), .C2(n9888), .A(n8694), .B(n8693), .ZN(n8711)
         );
  MUX2_X1 U10081 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8711), .S(n9952), .Z(
        P2_U3536) );
  INV_X2 U10082 ( .A(n9935), .ZN(n9937) );
  MUX2_X1 U10083 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8696), .S(n9937), .Z(
        P2_U3519) );
  MUX2_X1 U10084 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8697), .S(n9937), .Z(
        P2_U3518) );
  MUX2_X1 U10085 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8698), .S(n9937), .Z(
        P2_U3517) );
  MUX2_X1 U10086 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8699), .S(n9937), .Z(
        P2_U3516) );
  MUX2_X1 U10087 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8700), .S(n9937), .Z(
        P2_U3515) );
  MUX2_X1 U10088 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8701), .S(n9937), .Z(
        P2_U3514) );
  MUX2_X1 U10089 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8702), .S(n9937), .Z(
        P2_U3513) );
  MUX2_X1 U10090 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8703), .S(n9937), .Z(
        P2_U3512) );
  MUX2_X1 U10091 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8704), .S(n9937), .Z(
        P2_U3511) );
  MUX2_X1 U10092 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8705), .S(n9937), .Z(
        P2_U3510) );
  MUX2_X1 U10093 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8706), .S(n9937), .Z(
        P2_U3509) );
  MUX2_X1 U10094 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8707), .S(n9937), .Z(
        P2_U3508) );
  MUX2_X1 U10095 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8708), .S(n9937), .Z(
        P2_U3507) );
  MUX2_X1 U10096 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8709), .S(n9937), .Z(
        P2_U3505) );
  MUX2_X1 U10097 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8710), .S(n9937), .Z(
        P2_U3502) );
  MUX2_X1 U10098 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8711), .S(n9937), .Z(
        P2_U3499) );
  NAND3_X1 U10099 ( .A1(n4494), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8713) );
  OAI22_X1 U10100 ( .A1(n5562), .A2(n8713), .B1(n8712), .B2(n8722), .ZN(n8714)
         );
  AOI21_X1 U10101 ( .B1(n9405), .B2(n8715), .A(n8714), .ZN(n8716) );
  INV_X1 U10102 ( .A(n8716), .ZN(P2_U3327) );
  INV_X1 U10103 ( .A(n8717), .ZN(n9415) );
  OAI222_X1 U10104 ( .A1(n8720), .A2(P2_U3152), .B1(n8719), .B2(n9415), .C1(
        n8718), .C2(n8722), .ZN(P2_U3329) );
  INV_X1 U10105 ( .A(n8721), .ZN(n9418) );
  OAI222_X1 U10106 ( .A1(n6092), .A2(P2_U3152), .B1(n8719), .B2(n9418), .C1(
        n8723), .C2(n8722), .ZN(P2_U3330) );
  MUX2_X1 U10107 ( .A(n8724), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10108 ( .A1(n4798), .A2(n8725), .ZN(n8727) );
  XNOR2_X1 U10109 ( .A(n8727), .B(n8726), .ZN(n8732) );
  OAI22_X1 U10110 ( .A1(n9032), .A2(n8807), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8728), .ZN(n8730) );
  OAI22_X1 U10111 ( .A1(n9100), .A2(n8848), .B1(n8833), .B2(n9064), .ZN(n8729)
         );
  AOI211_X1 U10112 ( .C1(n9211), .C2(n8850), .A(n8730), .B(n8729), .ZN(n8731)
         );
  OAI21_X1 U10113 ( .B1(n8732), .B2(n8853), .A(n8731), .ZN(P1_U3214) );
  INV_X1 U10114 ( .A(n9223), .ZN(n8742) );
  OAI21_X1 U10115 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8736) );
  NAND2_X1 U10116 ( .A1(n8736), .A2(n8829), .ZN(n8741) );
  NOR2_X1 U10117 ( .A1(n8737), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8739) );
  OAI22_X1 U10118 ( .A1(n9100), .A2(n8807), .B1(n8833), .B2(n9104), .ZN(n8738)
         );
  AOI211_X1 U10119 ( .C1(n8831), .C2(n9137), .A(n8739), .B(n8738), .ZN(n8740)
         );
  OAI211_X1 U10120 ( .C1(n8742), .C2(n8837), .A(n8741), .B(n8740), .ZN(
        P1_U3221) );
  INV_X1 U10121 ( .A(n9203), .ZN(n9038) );
  OAI21_X1 U10122 ( .B1(n8744), .B2(n8743), .A(n8824), .ZN(n8745) );
  NAND2_X1 U10123 ( .A1(n8745), .A2(n8829), .ZN(n8751) );
  NOR2_X1 U10124 ( .A1(n8746), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8749) );
  INV_X1 U10125 ( .A(n9035), .ZN(n8747) );
  OAI22_X1 U10126 ( .A1(n9031), .A2(n8807), .B1(n8833), .B2(n8747), .ZN(n8748)
         );
  AOI211_X1 U10127 ( .C1(n8831), .C2(n9072), .A(n8749), .B(n8748), .ZN(n8750)
         );
  OAI211_X1 U10128 ( .C1(n9038), .C2(n8837), .A(n8751), .B(n8750), .ZN(
        P1_U3223) );
  INV_X1 U10129 ( .A(n8753), .ZN(n8754) );
  AOI21_X1 U10130 ( .B1(n8755), .B2(n8752), .A(n8754), .ZN(n8764) );
  OAI22_X1 U10131 ( .A1(n8848), .A2(n8757), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8756), .ZN(n8761) );
  INV_X1 U10132 ( .A(n8758), .ZN(n8759) );
  OAI22_X1 U10133 ( .A1(n8833), .A2(n8759), .B1(n8806), .B2(n8807), .ZN(n8760)
         );
  AOI211_X1 U10134 ( .C1(n8762), .C2(n8850), .A(n8761), .B(n8760), .ZN(n8763)
         );
  OAI21_X1 U10135 ( .B1(n8764), .B2(n8853), .A(n8763), .ZN(P1_U3224) );
  OAI21_X1 U10136 ( .B1(n8767), .B2(n8766), .A(n8765), .ZN(n8768) );
  NAND2_X1 U10137 ( .A1(n8768), .A2(n8829), .ZN(n8772) );
  AOI22_X1 U10138 ( .A1(n8831), .A2(n8857), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3084), .ZN(n8771) );
  AOI22_X1 U10139 ( .A1(n9171), .A2(n8844), .B1(n8843), .B2(n9138), .ZN(n8770)
         );
  NAND2_X1 U10140 ( .A1(n9243), .A2(n8850), .ZN(n8769) );
  NAND4_X1 U10141 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(
        P1_U3226) );
  INV_X1 U10142 ( .A(n8773), .ZN(n8774) );
  AOI21_X1 U10143 ( .B1(n8776), .B2(n8775), .A(n8774), .ZN(n8781) );
  AOI22_X1 U10144 ( .A1(n9054), .A2(n8843), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8778) );
  NAND2_X1 U10145 ( .A1(n9088), .A2(n8831), .ZN(n8777) );
  OAI211_X1 U10146 ( .C1(n8833), .C2(n9046), .A(n8778), .B(n8777), .ZN(n8779)
         );
  AOI21_X1 U10147 ( .B1(n9206), .B2(n8850), .A(n8779), .ZN(n8780) );
  OAI21_X1 U10148 ( .B1(n8781), .B2(n8853), .A(n8780), .ZN(P1_U3227) );
  OAI21_X1 U10149 ( .B1(n8784), .B2(n8783), .A(n8782), .ZN(n8789) );
  AOI22_X1 U10150 ( .A1(n8843), .A2(n9121), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8787) );
  INV_X1 U10151 ( .A(n8785), .ZN(n9116) );
  AOI22_X1 U10152 ( .A1(n9116), .A2(n8844), .B1(n8831), .B2(n9153), .ZN(n8786)
         );
  OAI211_X1 U10153 ( .C1(n9118), .C2(n8837), .A(n8787), .B(n8786), .ZN(n8788)
         );
  AOI21_X1 U10154 ( .B1(n8789), .B2(n8829), .A(n8788), .ZN(n8790) );
  INV_X1 U10155 ( .A(n8790), .ZN(P1_U3231) );
  NAND2_X1 U10156 ( .A1(n8792), .A2(n8791), .ZN(n8793) );
  XOR2_X1 U10157 ( .A(n8794), .B(n8793), .Z(n8800) );
  OAI22_X1 U10158 ( .A1(n8848), .A2(n8795), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9379), .ZN(n8798) );
  OAI22_X1 U10159 ( .A1(n8796), .A2(n8807), .B1(n8833), .B2(n9081), .ZN(n8797)
         );
  AOI211_X1 U10160 ( .C1(n9216), .C2(n8850), .A(n8798), .B(n8797), .ZN(n8799)
         );
  OAI21_X1 U10161 ( .B1(n8800), .B2(n8853), .A(n8799), .ZN(P1_U3233) );
  XNOR2_X1 U10162 ( .A(n8802), .B(n8801), .ZN(n8803) );
  XNOR2_X1 U10163 ( .A(n8804), .B(n8803), .ZN(n8812) );
  OAI22_X1 U10164 ( .A1(n8848), .A2(n8806), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8805), .ZN(n8810) );
  OAI22_X1 U10165 ( .A1(n8833), .A2(n9145), .B1(n8808), .B2(n8807), .ZN(n8809)
         );
  AOI211_X1 U10166 ( .C1(n9236), .C2(n8850), .A(n8810), .B(n8809), .ZN(n8811)
         );
  OAI21_X1 U10167 ( .B1(n8812), .B2(n8853), .A(n8811), .ZN(P1_U3236) );
  OAI21_X1 U10168 ( .B1(n8815), .B2(n8814), .A(n8813), .ZN(n8816) );
  NAND2_X1 U10169 ( .A1(n8816), .A2(n8829), .ZN(n8823) );
  AOI22_X1 U10170 ( .A1(n8817), .A2(n8850), .B1(n8843), .B2(n8866), .ZN(n8822)
         );
  AOI21_X1 U10171 ( .B1(n8831), .B2(n8868), .A(n8818), .ZN(n8821) );
  NAND2_X1 U10172 ( .A1(n8844), .A2(n8819), .ZN(n8820) );
  NAND4_X1 U10173 ( .A1(n8823), .A2(n8822), .A3(n8821), .A4(n8820), .ZN(
        P1_U3237) );
  INV_X1 U10174 ( .A(n9196), .ZN(n9014) );
  INV_X1 U10175 ( .A(n8824), .ZN(n8827) );
  OAI21_X1 U10176 ( .B1(n8827), .B2(n8826), .A(n8825), .ZN(n8830) );
  NAND3_X1 U10177 ( .A1(n8830), .A2(n8829), .A3(n8828), .ZN(n8836) );
  AOI22_X1 U10178 ( .A1(n9054), .A2(n8831), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8832) );
  OAI21_X1 U10179 ( .B1(n8833), .B2(n9011), .A(n8832), .ZN(n8834) );
  AOI21_X1 U10180 ( .B1(n8843), .B2(n9021), .A(n8834), .ZN(n8835) );
  OAI211_X1 U10181 ( .C1(n9014), .C2(n8837), .A(n8836), .B(n8835), .ZN(
        P1_U3238) );
  INV_X1 U10182 ( .A(n8838), .ZN(n8840) );
  NAND2_X1 U10183 ( .A1(n8840), .A2(n8839), .ZN(n8842) );
  XNOR2_X1 U10184 ( .A(n8842), .B(n8841), .ZN(n8854) );
  AOI22_X1 U10185 ( .A1(n8845), .A2(n8844), .B1(n8843), .B2(n8857), .ZN(n8847)
         );
  OAI211_X1 U10186 ( .C1(n9495), .C2(n8848), .A(n8847), .B(n8846), .ZN(n8849)
         );
  AOI21_X1 U10187 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8852) );
  OAI21_X1 U10188 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(P1_U3239) );
  INV_X2 U10189 ( .A(P1_U4006), .ZN(n9587) );
  MUX2_X1 U10190 ( .A(n8962), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9587), .Z(
        P1_U3586) );
  MUX2_X1 U10191 ( .A(n8855), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9587), .Z(
        P1_U3585) );
  MUX2_X1 U10192 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8979), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10193 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n5531), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10194 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9021), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10195 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n8856), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10196 ( .A(n9054), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9587), .Z(
        P1_U3580) );
  MUX2_X1 U10197 ( .A(n9072), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9587), .Z(
        P1_U3579) );
  MUX2_X1 U10198 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9088), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10199 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9071), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10200 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9121), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10201 ( .A(n9137), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9587), .Z(
        P1_U3575) );
  MUX2_X1 U10202 ( .A(n9153), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9587), .Z(
        P1_U3574) );
  MUX2_X1 U10203 ( .A(n9138), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9587), .Z(
        P1_U3573) );
  MUX2_X1 U10204 ( .A(n9155), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9587), .Z(
        P1_U3572) );
  MUX2_X1 U10205 ( .A(n8857), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9587), .Z(
        P1_U3571) );
  MUX2_X1 U10206 ( .A(n8858), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9587), .Z(
        P1_U3570) );
  MUX2_X1 U10207 ( .A(n8859), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9587), .Z(
        P1_U3569) );
  MUX2_X1 U10208 ( .A(n8860), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9587), .Z(
        P1_U3568) );
  MUX2_X1 U10209 ( .A(n8861), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9587), .Z(
        P1_U3567) );
  MUX2_X1 U10210 ( .A(n8862), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9587), .Z(
        P1_U3566) );
  MUX2_X1 U10211 ( .A(n8863), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9587), .Z(
        P1_U3565) );
  MUX2_X1 U10212 ( .A(n8864), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9587), .Z(
        P1_U3564) );
  MUX2_X1 U10213 ( .A(n8865), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9587), .Z(
        P1_U3563) );
  MUX2_X1 U10214 ( .A(n8866), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9587), .Z(
        P1_U3562) );
  MUX2_X1 U10215 ( .A(n8867), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9587), .Z(
        P1_U3561) );
  MUX2_X1 U10216 ( .A(n8868), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9587), .Z(
        P1_U3560) );
  MUX2_X1 U10217 ( .A(n8869), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9587), .Z(
        P1_U3559) );
  MUX2_X1 U10218 ( .A(n8870), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9587), .Z(
        P1_U3558) );
  MUX2_X1 U10219 ( .A(n6363), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9587), .Z(
        P1_U3557) );
  MUX2_X1 U10220 ( .A(n6335), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9587), .Z(
        P1_U3556) );
  MUX2_X1 U10221 ( .A(n6346), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9587), .Z(
        P1_U3555) );
  AOI211_X1 U10222 ( .C1(n8873), .C2(n8872), .A(n9575), .B(n8871), .ZN(n8874)
         );
  INV_X1 U10223 ( .A(n8874), .ZN(n8883) );
  AOI21_X1 U10224 ( .B1(n8933), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n8875), .ZN(
        n8882) );
  OAI21_X1 U10225 ( .B1(n8878), .B2(n8877), .A(n8876), .ZN(n8879) );
  AOI22_X1 U10226 ( .A1(n8880), .A2(n9654), .B1(n9662), .B2(n8879), .ZN(n8881)
         );
  NAND3_X1 U10227 ( .A1(n8883), .A2(n8882), .A3(n8881), .ZN(P1_U3249) );
  INV_X1 U10228 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n8885) );
  OAI21_X1 U10229 ( .B1(n9667), .B2(n8885), .A(n8884), .ZN(n8886) );
  AOI21_X1 U10230 ( .B1(n8887), .B2(n9654), .A(n8886), .ZN(n8897) );
  OAI21_X1 U10231 ( .B1(n8890), .B2(n8889), .A(n8888), .ZN(n8891) );
  NAND2_X1 U10232 ( .A1(n8891), .A2(n9661), .ZN(n8896) );
  OAI211_X1 U10233 ( .C1(n8894), .C2(n8893), .A(n9662), .B(n8892), .ZN(n8895)
         );
  NAND3_X1 U10234 ( .A1(n8897), .A2(n8896), .A3(n8895), .ZN(P1_U3254) );
  NOR2_X1 U10235 ( .A1(n8905), .A2(n8898), .ZN(n8900) );
  NOR2_X1 U10236 ( .A1(n8900), .A2(n8899), .ZN(n8903) );
  NAND2_X1 U10237 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n8921), .ZN(n8901) );
  OAI21_X1 U10238 ( .B1(n8921), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8901), .ZN(
        n8902) );
  NOR2_X1 U10239 ( .A1(n8903), .A2(n8902), .ZN(n8917) );
  AOI211_X1 U10240 ( .C1(n8903), .C2(n8902), .A(n8917), .B(n9626), .ZN(n8916)
         );
  NOR2_X1 U10241 ( .A1(n8905), .A2(n8904), .ZN(n8907) );
  INV_X1 U10242 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8908) );
  MUX2_X1 U10243 ( .A(n8908), .B(P1_REG1_REG_16__SCAN_IN), .S(n8921), .Z(n8909) );
  NOR2_X1 U10244 ( .A1(n8910), .A2(n8909), .ZN(n8920) );
  AOI211_X1 U10245 ( .C1(n8910), .C2(n8909), .A(n8920), .B(n9575), .ZN(n8915)
         );
  NAND2_X1 U10246 ( .A1(n8933), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n8912) );
  NAND2_X1 U10247 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3084), .ZN(n8911) );
  OAI211_X1 U10248 ( .C1(n9634), .C2(n8913), .A(n8912), .B(n8911), .ZN(n8914)
         );
  OR3_X1 U10249 ( .A1(n8916), .A2(n8915), .A3(n8914), .ZN(P1_U3257) );
  XNOR2_X1 U10250 ( .A(n8939), .B(P1_REG2_REG_17__SCAN_IN), .ZN(n8919) );
  AOI21_X1 U10251 ( .B1(n8921), .B2(P1_REG2_REG_16__SCAN_IN), .A(n8917), .ZN(
        n8918) );
  NOR2_X1 U10252 ( .A1(n8918), .A2(n8919), .ZN(n8938) );
  AOI211_X1 U10253 ( .C1(n8919), .C2(n8918), .A(n8938), .B(n9626), .ZN(n8929)
         );
  XNOR2_X1 U10254 ( .A(n8939), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n8923) );
  AOI21_X1 U10255 ( .B1(n8921), .B2(P1_REG1_REG_16__SCAN_IN), .A(n8920), .ZN(
        n8922) );
  NOR2_X1 U10256 ( .A1(n8922), .A2(n8923), .ZN(n8930) );
  AOI211_X1 U10257 ( .C1(n8923), .C2(n8922), .A(n8930), .B(n9575), .ZN(n8928)
         );
  INV_X1 U10258 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n8926) );
  NAND2_X1 U10259 ( .A1(n9654), .A2(n8939), .ZN(n8925) );
  NAND2_X1 U10260 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n8924) );
  OAI211_X1 U10261 ( .C1(n9667), .C2(n8926), .A(n8925), .B(n8924), .ZN(n8927)
         );
  OR3_X1 U10262 ( .A1(n8929), .A2(n8928), .A3(n8927), .ZN(P1_U3258) );
  XNOR2_X1 U10263 ( .A(n8936), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U10264 ( .A1(n8932), .A2(n8931), .ZN(n8949) );
  OAI21_X1 U10265 ( .B1(n8932), .B2(n8931), .A(n8949), .ZN(n8944) );
  NAND2_X1 U10266 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_U3084), .ZN(n8935) );
  NAND2_X1 U10267 ( .A1(n8933), .A2(P1_ADDR_REG_18__SCAN_IN), .ZN(n8934) );
  OAI211_X1 U10268 ( .C1(n8936), .C2(n9634), .A(n8935), .B(n8934), .ZN(n8943)
         );
  NAND2_X1 U10269 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n8950), .ZN(n8937) );
  OAI21_X1 U10270 ( .B1(n8950), .B2(P1_REG2_REG_18__SCAN_IN), .A(n8937), .ZN(
        n8941) );
  AOI211_X1 U10271 ( .C1(n8941), .C2(n8940), .A(n8946), .B(n9626), .ZN(n8942)
         );
  AOI211_X1 U10272 ( .C1(n9661), .C2(n8944), .A(n8943), .B(n8942), .ZN(n8945)
         );
  INV_X1 U10273 ( .A(n8945), .ZN(P1_U3259) );
  INV_X1 U10274 ( .A(n8955), .ZN(n8953) );
  INV_X1 U10275 ( .A(n8948), .ZN(n8952) );
  OAI21_X1 U10276 ( .B1(n8954), .B2(n9575), .A(n9634), .ZN(n8951) );
  AOI22_X1 U10277 ( .A1(n8955), .A2(n9662), .B1(n8954), .B2(n9661), .ZN(n8956)
         );
  OAI211_X1 U10278 ( .C1(n8959), .C2(n9667), .A(n8958), .B(n8957), .ZN(
        P1_U3260) );
  NAND2_X1 U10279 ( .A1(n9523), .A2(n8966), .ZN(n8960) );
  XNOR2_X1 U10280 ( .A(n8960), .B(n9177), .ZN(n9179) );
  NAND2_X1 U10281 ( .A1(n8962), .A2(n8961), .ZN(n9522) );
  NOR2_X1 U10282 ( .A1(n9708), .A2(n9522), .ZN(n8968) );
  NOR2_X1 U10283 ( .A1(n9684), .A2(n8963), .ZN(n8964) );
  AOI211_X1 U10284 ( .C1(n9177), .C2(n9107), .A(n8968), .B(n8964), .ZN(n8965)
         );
  OAI21_X1 U10285 ( .B1(n9179), .B2(n8985), .A(n8965), .ZN(P1_U3261) );
  XNOR2_X1 U10286 ( .A(n8967), .B(n8966), .ZN(n9525) );
  NAND2_X1 U10287 ( .A1(n9525), .A2(n9692), .ZN(n8970) );
  AOI21_X1 U10288 ( .B1(n9517), .B2(P1_REG2_REG_30__SCAN_IN), .A(n8968), .ZN(
        n8969) );
  OAI211_X1 U10289 ( .C1(n9523), .C2(n9710), .A(n8970), .B(n8969), .ZN(
        P1_U3262) );
  NAND2_X1 U10290 ( .A1(n8971), .A2(n8972), .ZN(n8973) );
  NAND2_X1 U10291 ( .A1(n8974), .A2(n8973), .ZN(n9188) );
  AND2_X1 U10292 ( .A1(n8976), .A2(n8975), .ZN(n8977) );
  OAI21_X1 U10293 ( .B1(n8978), .B2(n8977), .A(n9701), .ZN(n8981) );
  AOI22_X1 U10294 ( .A1(n9021), .A2(n9154), .B1(n8979), .B2(n9152), .ZN(n8980)
         );
  NAND2_X1 U10295 ( .A1(n8981), .A2(n8980), .ZN(n9187) );
  NAND2_X1 U10296 ( .A1(n8993), .A2(n8982), .ZN(n8983) );
  NAND2_X1 U10297 ( .A1(n8984), .A2(n8983), .ZN(n9185) );
  NOR2_X1 U10298 ( .A1(n9185), .A2(n8985), .ZN(n8990) );
  INV_X1 U10299 ( .A(n8986), .ZN(n8987) );
  AOI22_X1 U10300 ( .A1(n8987), .A2(n9707), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n9517), .ZN(n8988) );
  OAI21_X1 U10301 ( .B1(n9184), .B2(n9710), .A(n8988), .ZN(n8989) );
  AOI211_X1 U10302 ( .C1(n9187), .C2(n9684), .A(n8990), .B(n8989), .ZN(n8991)
         );
  OAI21_X1 U10303 ( .B1(n9176), .B2(n9188), .A(n8991), .ZN(P1_U3263) );
  XNOR2_X1 U10304 ( .A(n8992), .B(n8999), .ZN(n9195) );
  INV_X1 U10305 ( .A(n9010), .ZN(n8995) );
  INV_X1 U10306 ( .A(n8993), .ZN(n8994) );
  AOI21_X1 U10307 ( .B1(n9191), .B2(n8995), .A(n8994), .ZN(n9192) );
  AOI22_X1 U10308 ( .A1(n8996), .A2(n9707), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n9517), .ZN(n8997) );
  OAI21_X1 U10309 ( .B1(n8998), .B2(n9710), .A(n8997), .ZN(n9006) );
  AOI21_X1 U10310 ( .B1(n9000), .B2(n8999), .A(n9163), .ZN(n9004) );
  OAI22_X1 U10311 ( .A1(n9001), .A2(n9698), .B1(n9031), .B2(n9696), .ZN(n9002)
         );
  AOI21_X1 U10312 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9194) );
  NOR2_X1 U10313 ( .A1(n9194), .A2(n9517), .ZN(n9005) );
  AOI211_X1 U10314 ( .C1(n9692), .C2(n9192), .A(n9006), .B(n9005), .ZN(n9007)
         );
  OAI21_X1 U10315 ( .B1(n9195), .B2(n9176), .A(n9007), .ZN(P1_U3264) );
  XNOR2_X1 U10316 ( .A(n9009), .B(n9008), .ZN(n9200) );
  AOI21_X1 U10317 ( .B1(n9196), .B2(n9033), .A(n9010), .ZN(n9197) );
  INV_X1 U10318 ( .A(n9011), .ZN(n9012) );
  AOI22_X1 U10319 ( .A1(n9012), .A2(n9707), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9517), .ZN(n9013) );
  OAI21_X1 U10320 ( .B1(n9014), .B2(n9710), .A(n9013), .ZN(n9023) );
  NAND2_X1 U10321 ( .A1(n9029), .A2(n9016), .ZN(n9018) );
  NAND2_X1 U10322 ( .A1(n9018), .A2(n9017), .ZN(n9020) );
  NOR2_X1 U10323 ( .A1(n9199), .A2(n9517), .ZN(n9022) );
  AOI211_X1 U10324 ( .C1(n9197), .C2(n9692), .A(n9023), .B(n9022), .ZN(n9024)
         );
  OAI21_X1 U10325 ( .B1(n9176), .B2(n9200), .A(n9024), .ZN(P1_U3265) );
  INV_X1 U10326 ( .A(n9025), .ZN(n9026) );
  AOI21_X1 U10327 ( .B1(n9028), .B2(n9027), .A(n9026), .ZN(n9205) );
  XNOR2_X1 U10328 ( .A(n9029), .B(n9028), .ZN(n9030) );
  OAI222_X1 U10329 ( .A1(n9696), .A2(n9032), .B1(n9698), .B2(n9031), .C1(n9030), .C2(n9163), .ZN(n9201) );
  INV_X1 U10330 ( .A(n9033), .ZN(n9034) );
  AOI211_X1 U10331 ( .C1(n9203), .C2(n9044), .A(n9761), .B(n9034), .ZN(n9202)
         );
  NAND2_X1 U10332 ( .A1(n9202), .A2(n9170), .ZN(n9037) );
  AOI22_X1 U10333 ( .A1(n9035), .A2(n9707), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9517), .ZN(n9036) );
  OAI211_X1 U10334 ( .C1(n9038), .C2(n9710), .A(n9037), .B(n9036), .ZN(n9039)
         );
  AOI21_X1 U10335 ( .B1(n9201), .B2(n9684), .A(n9039), .ZN(n9040) );
  OAI21_X1 U10336 ( .B1(n9205), .B2(n9176), .A(n9040), .ZN(P1_U3266) );
  OAI21_X1 U10337 ( .B1(n9043), .B2(n9042), .A(n9041), .ZN(n9210) );
  INV_X1 U10338 ( .A(n9062), .ZN(n9045) );
  AOI21_X1 U10339 ( .B1(n9206), .B2(n9045), .A(n4505), .ZN(n9207) );
  INV_X1 U10340 ( .A(n9046), .ZN(n9047) );
  AOI22_X1 U10341 ( .A1(n9047), .A2(n9707), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9517), .ZN(n9048) );
  OAI21_X1 U10342 ( .B1(n9049), .B2(n9710), .A(n9048), .ZN(n9057) );
  INV_X1 U10343 ( .A(n9050), .ZN(n9053) );
  OAI21_X1 U10344 ( .B1(n9053), .B2(n9052), .A(n9051), .ZN(n9055) );
  AOI222_X1 U10345 ( .A1(n9701), .A2(n9055), .B1(n9088), .B2(n9154), .C1(n9054), .C2(n9152), .ZN(n9209) );
  NOR2_X1 U10346 ( .A1(n9209), .A2(n9517), .ZN(n9056) );
  AOI211_X1 U10347 ( .C1(n9207), .C2(n9692), .A(n9057), .B(n9056), .ZN(n9058)
         );
  OAI21_X1 U10348 ( .B1(n9176), .B2(n9210), .A(n9058), .ZN(P1_U3267) );
  OAI21_X1 U10349 ( .B1(n9061), .B2(n9060), .A(n9059), .ZN(n9215) );
  INV_X1 U10350 ( .A(n9080), .ZN(n9063) );
  AOI21_X1 U10351 ( .B1(n9211), .B2(n9063), .A(n9062), .ZN(n9212) );
  INV_X1 U10352 ( .A(n9064), .ZN(n9065) );
  AOI22_X1 U10353 ( .A1(n9065), .A2(n9707), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n9517), .ZN(n9066) );
  OAI21_X1 U10354 ( .B1(n9067), .B2(n9710), .A(n9066), .ZN(n9076) );
  OAI211_X1 U10355 ( .C1(n9070), .C2(n9069), .A(n9068), .B(n9701), .ZN(n9074)
         );
  AOI22_X1 U10356 ( .A1(n9072), .A2(n9152), .B1(n9154), .B2(n9071), .ZN(n9073)
         );
  AND2_X1 U10357 ( .A1(n9074), .A2(n9073), .ZN(n9214) );
  NOR2_X1 U10358 ( .A1(n9214), .A2(n9517), .ZN(n9075) );
  AOI211_X1 U10359 ( .C1(n9212), .C2(n9692), .A(n9076), .B(n9075), .ZN(n9077)
         );
  OAI21_X1 U10360 ( .B1(n9176), .B2(n9215), .A(n9077), .ZN(P1_U3268) );
  OAI21_X1 U10361 ( .B1(n9079), .B2(n9087), .A(n9078), .ZN(n9220) );
  AOI21_X1 U10362 ( .B1(n9216), .B2(n9101), .A(n9080), .ZN(n9217) );
  INV_X1 U10363 ( .A(n9216), .ZN(n9084) );
  INV_X1 U10364 ( .A(n9081), .ZN(n9082) );
  AOI22_X1 U10365 ( .A1(n9082), .A2(n9707), .B1(n9708), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9083) );
  OAI21_X1 U10366 ( .B1(n9084), .B2(n9710), .A(n9083), .ZN(n9091) );
  NAND2_X1 U10367 ( .A1(n9094), .A2(n9085), .ZN(n9086) );
  XOR2_X1 U10368 ( .A(n9087), .B(n9086), .Z(n9089) );
  AOI222_X1 U10369 ( .A1(n9701), .A2(n9089), .B1(n9121), .B2(n9154), .C1(n9088), .C2(n9152), .ZN(n9219) );
  NOR2_X1 U10370 ( .A1(n9219), .A2(n9517), .ZN(n9090) );
  AOI211_X1 U10371 ( .C1(n9217), .C2(n9692), .A(n9091), .B(n9090), .ZN(n9092)
         );
  OAI21_X1 U10372 ( .B1(n9176), .B2(n9220), .A(n9092), .ZN(P1_U3269) );
  OAI21_X1 U10373 ( .B1(n4295), .B2(n9097), .A(n9093), .ZN(n9225) );
  INV_X1 U10374 ( .A(n9094), .ZN(n9095) );
  AOI21_X1 U10375 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9098) );
  OAI222_X1 U10376 ( .A1(n9698), .A2(n9100), .B1(n9696), .B2(n9099), .C1(n9163), .C2(n9098), .ZN(n9221) );
  AOI21_X1 U10377 ( .B1(n9113), .B2(n9223), .A(n9761), .ZN(n9102) );
  AND2_X1 U10378 ( .A1(n9102), .A2(n9101), .ZN(n9222) );
  NAND2_X1 U10379 ( .A1(n9222), .A2(n5254), .ZN(n9103) );
  OAI21_X1 U10380 ( .B1(n9105), .B2(n9104), .A(n9103), .ZN(n9106) );
  OAI21_X1 U10381 ( .B1(n9221), .B2(n9106), .A(n9684), .ZN(n9109) );
  AOI22_X1 U10382 ( .A1(n9223), .A2(n9107), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9708), .ZN(n9108) );
  OAI211_X1 U10383 ( .C1(n9225), .C2(n9176), .A(n9109), .B(n9108), .ZN(
        P1_U3270) );
  XNOR2_X1 U10384 ( .A(n9112), .B(n9111), .ZN(n9230) );
  INV_X1 U10385 ( .A(n9128), .ZN(n9115) );
  INV_X1 U10386 ( .A(n9113), .ZN(n9114) );
  AOI21_X1 U10387 ( .B1(n9226), .B2(n9115), .A(n9114), .ZN(n9227) );
  AOI22_X1 U10388 ( .A1(n9708), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9116), .B2(
        n9707), .ZN(n9117) );
  OAI21_X1 U10389 ( .B1(n9118), .B2(n9710), .A(n9117), .ZN(n9124) );
  XNOR2_X1 U10390 ( .A(n9120), .B(n9119), .ZN(n9122) );
  AOI222_X1 U10391 ( .A1(n9701), .A2(n9122), .B1(n9153), .B2(n9154), .C1(n9121), .C2(n9152), .ZN(n9229) );
  NOR2_X1 U10392 ( .A1(n9229), .A2(n9708), .ZN(n9123) );
  AOI211_X1 U10393 ( .C1(n9227), .C2(n9692), .A(n9124), .B(n9123), .ZN(n9125)
         );
  OAI21_X1 U10394 ( .B1(n9230), .B2(n9176), .A(n9125), .ZN(P1_U3271) );
  XNOR2_X1 U10395 ( .A(n9126), .B(n9127), .ZN(n9235) );
  INV_X1 U10396 ( .A(n9144), .ZN(n9129) );
  AOI211_X1 U10397 ( .C1(n9232), .C2(n9129), .A(n9761), .B(n9128), .ZN(n9231)
         );
  INV_X1 U10398 ( .A(n9130), .ZN(n9131) );
  AOI22_X1 U10399 ( .A1(n9708), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9131), .B2(
        n9707), .ZN(n9132) );
  OAI21_X1 U10400 ( .B1(n9133), .B2(n9710), .A(n9132), .ZN(n9141) );
  OAI21_X1 U10401 ( .B1(n9136), .B2(n9135), .A(n9134), .ZN(n9139) );
  AOI222_X1 U10402 ( .A1(n9701), .A2(n9139), .B1(n9138), .B2(n9154), .C1(n9137), .C2(n9152), .ZN(n9234) );
  NOR2_X1 U10403 ( .A1(n9234), .A2(n9708), .ZN(n9140) );
  AOI211_X1 U10404 ( .C1(n9231), .C2(n9170), .A(n9141), .B(n9140), .ZN(n9142)
         );
  OAI21_X1 U10405 ( .B1(n9176), .B2(n9235), .A(n9142), .ZN(P1_U3272) );
  XNOR2_X1 U10406 ( .A(n9143), .B(n9149), .ZN(n9240) );
  AOI21_X1 U10407 ( .B1(n9236), .B2(n9167), .A(n9144), .ZN(n9237) );
  INV_X1 U10408 ( .A(n9236), .ZN(n9148) );
  INV_X1 U10409 ( .A(n9145), .ZN(n9146) );
  AOI22_X1 U10410 ( .A1(n9708), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9146), .B2(
        n9707), .ZN(n9147) );
  OAI21_X1 U10411 ( .B1(n9148), .B2(n9710), .A(n9147), .ZN(n9158) );
  OAI21_X1 U10412 ( .B1(n9151), .B2(n5241), .A(n9150), .ZN(n9156) );
  AOI222_X1 U10413 ( .A1(n9701), .A2(n9156), .B1(n9155), .B2(n9154), .C1(n9153), .C2(n9152), .ZN(n9239) );
  NOR2_X1 U10414 ( .A1(n9239), .A2(n9517), .ZN(n9157) );
  AOI211_X1 U10415 ( .C1(n9237), .C2(n9692), .A(n9158), .B(n9157), .ZN(n9159)
         );
  OAI21_X1 U10416 ( .B1(n9176), .B2(n9240), .A(n9159), .ZN(P1_U3273) );
  XOR2_X1 U10417 ( .A(n9160), .B(n9161), .Z(n9246) );
  XNOR2_X1 U10418 ( .A(n9162), .B(n9161), .ZN(n9164) );
  OAI222_X1 U10419 ( .A1(n9698), .A2(n9166), .B1(n9696), .B2(n9165), .C1(n9164), .C2(n9163), .ZN(n9241) );
  INV_X1 U10420 ( .A(n9167), .ZN(n9168) );
  AOI211_X1 U10421 ( .C1(n9243), .C2(n9169), .A(n9761), .B(n9168), .ZN(n9242)
         );
  NAND2_X1 U10422 ( .A1(n9242), .A2(n9170), .ZN(n9173) );
  AOI22_X1 U10423 ( .A1(n9708), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9171), .B2(
        n9707), .ZN(n9172) );
  OAI211_X1 U10424 ( .C1(n4498), .C2(n9710), .A(n9173), .B(n9172), .ZN(n9174)
         );
  AOI21_X1 U10425 ( .B1(n9241), .B2(n9684), .A(n9174), .ZN(n9175) );
  OAI21_X1 U10426 ( .B1(n9246), .B2(n9176), .A(n9175), .ZN(P1_U3274) );
  NAND2_X1 U10427 ( .A1(n9177), .A2(n9244), .ZN(n9178) );
  OAI211_X1 U10428 ( .C1(n9179), .C2(n9761), .A(n9522), .B(n9178), .ZN(n9254)
         );
  MUX2_X1 U10429 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9254), .S(n9783), .Z(
        P1_U3554) );
  MUX2_X1 U10430 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9255), .S(n9783), .Z(
        P1_U3552) );
  OAI22_X1 U10431 ( .A1(n9185), .A2(n9761), .B1(n9184), .B2(n9759), .ZN(n9186)
         );
  NOR2_X1 U10432 ( .A1(n9187), .A2(n9186), .ZN(n9190) );
  NAND2_X1 U10433 ( .A1(n9190), .A2(n9189), .ZN(n9256) );
  MUX2_X1 U10434 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9256), .S(n9783), .Z(
        P1_U3551) );
  AOI22_X1 U10435 ( .A1(n9192), .A2(n9526), .B1(n9244), .B2(n9191), .ZN(n9193)
         );
  OAI211_X1 U10436 ( .C1(n9195), .C2(n9529), .A(n9194), .B(n9193), .ZN(n9257)
         );
  MUX2_X1 U10437 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9257), .S(n9783), .Z(
        P1_U3550) );
  AOI22_X1 U10438 ( .A1(n9197), .A2(n9526), .B1(n9244), .B2(n9196), .ZN(n9198)
         );
  OAI211_X1 U10439 ( .C1(n9529), .C2(n9200), .A(n9199), .B(n9198), .ZN(n9258)
         );
  MUX2_X1 U10440 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9258), .S(n9783), .Z(
        P1_U3549) );
  OAI21_X1 U10441 ( .B1(n9529), .B2(n9205), .A(n9204), .ZN(n9259) );
  MUX2_X1 U10442 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9259), .S(n9783), .Z(
        P1_U3548) );
  AOI22_X1 U10443 ( .A1(n9207), .A2(n9526), .B1(n9244), .B2(n9206), .ZN(n9208)
         );
  OAI211_X1 U10444 ( .C1(n9529), .C2(n9210), .A(n9209), .B(n9208), .ZN(n9260)
         );
  MUX2_X1 U10445 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9260), .S(n9783), .Z(
        P1_U3547) );
  AOI22_X1 U10446 ( .A1(n9212), .A2(n9526), .B1(n9244), .B2(n9211), .ZN(n9213)
         );
  OAI211_X1 U10447 ( .C1(n9215), .C2(n9529), .A(n9214), .B(n9213), .ZN(n9394)
         );
  MUX2_X1 U10448 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9394), .S(n9783), .Z(
        P1_U3546) );
  AOI22_X1 U10449 ( .A1(n9217), .A2(n9526), .B1(n9244), .B2(n9216), .ZN(n9218)
         );
  OAI211_X1 U10450 ( .C1(n9529), .C2(n9220), .A(n9219), .B(n9218), .ZN(n9395)
         );
  MUX2_X1 U10451 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9395), .S(n9783), .Z(
        P1_U3545) );
  AOI211_X1 U10452 ( .C1(n9244), .C2(n9223), .A(n9222), .B(n9221), .ZN(n9224)
         );
  OAI21_X1 U10453 ( .B1(n9529), .B2(n9225), .A(n9224), .ZN(n9396) );
  MUX2_X1 U10454 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9396), .S(n9783), .Z(
        P1_U3544) );
  AOI22_X1 U10455 ( .A1(n9227), .A2(n9526), .B1(n9244), .B2(n9226), .ZN(n9228)
         );
  OAI211_X1 U10456 ( .C1(n9529), .C2(n9230), .A(n9229), .B(n9228), .ZN(n9397)
         );
  MUX2_X1 U10457 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9397), .S(n9783), .Z(
        P1_U3543) );
  AOI21_X1 U10458 ( .B1(n9244), .B2(n9232), .A(n9231), .ZN(n9233) );
  OAI211_X1 U10459 ( .C1(n9529), .C2(n9235), .A(n9234), .B(n9233), .ZN(n9398)
         );
  MUX2_X1 U10460 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9398), .S(n9783), .Z(
        P1_U3542) );
  AOI22_X1 U10461 ( .A1(n9237), .A2(n9526), .B1(n9244), .B2(n9236), .ZN(n9238)
         );
  OAI211_X1 U10462 ( .C1(n9529), .C2(n9240), .A(n9239), .B(n9238), .ZN(n9399)
         );
  MUX2_X1 U10463 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9399), .S(n9783), .Z(
        P1_U3541) );
  AOI211_X1 U10464 ( .C1(n9244), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9245)
         );
  OAI21_X1 U10465 ( .B1(n9529), .B2(n9246), .A(n9245), .ZN(n9400) );
  MUX2_X1 U10466 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9400), .S(n9783), .Z(
        P1_U3540) );
  INV_X1 U10467 ( .A(n9247), .ZN(n9766) );
  OAI22_X1 U10468 ( .A1(n9249), .A2(n9761), .B1(n9248), .B2(n9759), .ZN(n9250)
         );
  AOI21_X1 U10469 ( .B1(n9251), .B2(n9766), .A(n9250), .ZN(n9252) );
  NAND2_X1 U10470 ( .A1(n9253), .A2(n9252), .ZN(n9401) );
  MUX2_X1 U10471 ( .A(n9401), .B(P1_REG1_REG_15__SCAN_IN), .S(n9780), .Z(
        P1_U3538) );
  MUX2_X1 U10472 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9254), .S(n9767), .Z(
        P1_U3522) );
  MUX2_X1 U10473 ( .A(n9256), .B(P1_REG0_REG_28__SCAN_IN), .S(n4495), .Z(
        P1_U3519) );
  MUX2_X1 U10474 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9257), .S(n9767), .Z(
        P1_U3518) );
  MUX2_X1 U10475 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9258), .S(n9767), .Z(
        P1_U3517) );
  MUX2_X1 U10476 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9259), .S(n9767), .Z(
        P1_U3516) );
  MUX2_X1 U10477 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9260), .S(n9767), .Z(n9393) );
  NOR2_X1 U10478 ( .A1(keyinput53), .A2(keyinput4), .ZN(n9265) );
  NAND2_X1 U10479 ( .A1(keyinput59), .A2(keyinput8), .ZN(n9263) );
  NOR2_X1 U10480 ( .A1(keyinput43), .A2(keyinput10), .ZN(n9261) );
  NAND3_X1 U10481 ( .A1(keyinput23), .A2(keyinput58), .A3(n9261), .ZN(n9262)
         );
  NOR4_X1 U10482 ( .A1(keyinput29), .A2(keyinput14), .A3(n9263), .A4(n9262), 
        .ZN(n9264) );
  NAND4_X1 U10483 ( .A1(keyinput31), .A2(keyinput49), .A3(n9265), .A4(n9264), 
        .ZN(n9285) );
  AND4_X1 U10484 ( .A1(keyinput61), .A2(keyinput21), .A3(keyinput25), .A4(
        keyinput26), .ZN(n9275) );
  NOR4_X1 U10485 ( .A1(keyinput20), .A2(keyinput37), .A3(keyinput36), .A4(
        keyinput60), .ZN(n9274) );
  NAND3_X1 U10486 ( .A1(keyinput24), .A2(keyinput0), .A3(keyinput1), .ZN(n9267) );
  NAND3_X1 U10487 ( .A1(keyinput28), .A2(keyinput48), .A3(keyinput27), .ZN(
        n9266) );
  NOR4_X1 U10488 ( .A1(keyinput54), .A2(keyinput13), .A3(n9267), .A4(n9266), 
        .ZN(n9273) );
  NAND4_X1 U10489 ( .A1(keyinput17), .A2(keyinput45), .A3(keyinput52), .A4(
        keyinput42), .ZN(n9271) );
  NAND4_X1 U10490 ( .A1(keyinput47), .A2(keyinput46), .A3(keyinput35), .A4(
        keyinput50), .ZN(n9270) );
  NAND4_X1 U10491 ( .A1(keyinput62), .A2(keyinput15), .A3(keyinput51), .A4(
        keyinput7), .ZN(n9269) );
  NAND4_X1 U10492 ( .A1(keyinput2), .A2(keyinput6), .A3(keyinput22), .A4(
        keyinput30), .ZN(n9268) );
  NOR4_X1 U10493 ( .A1(n9271), .A2(n9270), .A3(n9269), .A4(n9268), .ZN(n9272)
         );
  NAND4_X1 U10494 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n9284)
         );
  NOR4_X1 U10495 ( .A1(keyinput33), .A2(keyinput41), .A3(keyinput57), .A4(
        keyinput12), .ZN(n9278) );
  NOR4_X1 U10496 ( .A1(keyinput16), .A2(keyinput40), .A3(keyinput32), .A4(
        keyinput38), .ZN(n9277) );
  NOR4_X1 U10497 ( .A1(keyinput39), .A2(keyinput63), .A3(keyinput11), .A4(
        keyinput3), .ZN(n9276) );
  AND3_X1 U10498 ( .A1(n9278), .A2(n9277), .A3(n9276), .ZN(n9282) );
  NOR3_X1 U10499 ( .A1(keyinput19), .A2(keyinput18), .A3(keyinput55), .ZN(
        n9281) );
  AND3_X1 U10500 ( .A1(keyinput44), .A2(keyinput34), .A3(keyinput56), .ZN(
        n9280) );
  AND2_X1 U10501 ( .A1(keyinput9), .A2(keyinput5), .ZN(n9279) );
  NAND4_X1 U10502 ( .A1(n9282), .A2(n9281), .A3(n9280), .A4(n9279), .ZN(n9283)
         );
  NOR3_X1 U10503 ( .A1(n9285), .A2(n9284), .A3(n9283), .ZN(n9352) );
  XNOR2_X1 U10504 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput18), .ZN(n9289) );
  XNOR2_X1 U10505 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput7), .ZN(n9288) );
  XNOR2_X1 U10506 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput40), .ZN(n9287) );
  XNOR2_X1 U10507 ( .A(P1_REG0_REG_21__SCAN_IN), .B(keyinput57), .ZN(n9286) );
  NAND4_X1 U10508 ( .A1(n9289), .A2(n9288), .A3(n9287), .A4(n9286), .ZN(n9295)
         );
  XNOR2_X1 U10509 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput47), .ZN(n9293) );
  XNOR2_X1 U10510 ( .A(P1_REG1_REG_17__SCAN_IN), .B(keyinput32), .ZN(n9292) );
  XNOR2_X1 U10511 ( .A(P1_REG0_REG_25__SCAN_IN), .B(keyinput42), .ZN(n9291) );
  XNOR2_X1 U10512 ( .A(P2_IR_REG_25__SCAN_IN), .B(keyinput38), .ZN(n9290) );
  NAND4_X1 U10513 ( .A1(n9293), .A2(n9292), .A3(n9291), .A4(n9290), .ZN(n9294)
         );
  NOR2_X1 U10514 ( .A1(n9295), .A2(n9294), .ZN(n9311) );
  XNOR2_X1 U10515 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput50), .ZN(n9299) );
  XNOR2_X1 U10516 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput53), .ZN(n9298) );
  XNOR2_X1 U10517 ( .A(SI_11_), .B(keyinput13), .ZN(n9297) );
  XNOR2_X1 U10518 ( .A(P1_REG1_REG_23__SCAN_IN), .B(keyinput60), .ZN(n9296) );
  NAND4_X1 U10519 ( .A1(n9299), .A2(n9298), .A3(n9297), .A4(n9296), .ZN(n9305)
         );
  XNOR2_X1 U10520 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput36), .ZN(n9303) );
  XNOR2_X1 U10521 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput28), .ZN(n9302) );
  XNOR2_X1 U10522 ( .A(P1_REG1_REG_29__SCAN_IN), .B(keyinput31), .ZN(n9301) );
  XNOR2_X1 U10523 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput37), .ZN(n9300) );
  NAND4_X1 U10524 ( .A1(n9303), .A2(n9302), .A3(n9301), .A4(n9300), .ZN(n9304)
         );
  NOR2_X1 U10525 ( .A1(n9305), .A2(n9304), .ZN(n9310) );
  INV_X1 U10526 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n9718) );
  INV_X1 U10527 ( .A(keyinput11), .ZN(n9306) );
  XNOR2_X1 U10528 ( .A(n9718), .B(n9306), .ZN(n9309) );
  INV_X1 U10529 ( .A(keyinput20), .ZN(n9307) );
  XNOR2_X1 U10530 ( .A(n9719), .B(n9307), .ZN(n9308) );
  NAND4_X1 U10531 ( .A1(n9311), .A2(n9310), .A3(n9309), .A4(n9308), .ZN(n9351)
         );
  INV_X1 U10532 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9717) );
  AOI22_X1 U10533 ( .A1(n9717), .A2(keyinput41), .B1(keyinput39), .B2(n9313), 
        .ZN(n9312) );
  OAI221_X1 U10534 ( .B1(n9717), .B2(keyinput41), .C1(n9313), .C2(keyinput39), 
        .A(n9312), .ZN(n9317) );
  INV_X1 U10535 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U10536 ( .A1(n9856), .A2(keyinput45), .B1(n9315), .B2(keyinput6), 
        .ZN(n9314) );
  OAI221_X1 U10537 ( .B1(n9856), .B2(keyinput45), .C1(n9315), .C2(keyinput6), 
        .A(n9314), .ZN(n9316) );
  NOR2_X1 U10538 ( .A1(n9317), .A2(n9316), .ZN(n9325) );
  AOI22_X1 U10539 ( .A1(n6861), .A2(keyinput19), .B1(n9319), .B2(keyinput5), 
        .ZN(n9318) );
  OAI221_X1 U10540 ( .B1(n6861), .B2(keyinput19), .C1(n9319), .C2(keyinput5), 
        .A(n9318), .ZN(n9323) );
  AOI22_X1 U10541 ( .A1(n4878), .A2(keyinput12), .B1(n9321), .B2(keyinput16), 
        .ZN(n9320) );
  OAI221_X1 U10542 ( .B1(n4878), .B2(keyinput12), .C1(n9321), .C2(keyinput16), 
        .A(n9320), .ZN(n9322) );
  NOR2_X1 U10543 ( .A1(n9323), .A2(n9322), .ZN(n9324) );
  AND2_X1 U10544 ( .A1(n9325), .A2(n9324), .ZN(n9349) );
  INV_X1 U10545 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n9716) );
  INV_X1 U10546 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9720) );
  AOI22_X1 U10547 ( .A1(n9716), .A2(keyinput33), .B1(keyinput62), .B2(n9720), 
        .ZN(n9326) );
  OAI221_X1 U10548 ( .B1(n9716), .B2(keyinput33), .C1(n9720), .C2(keyinput62), 
        .A(n9326), .ZN(n9334) );
  INV_X1 U10549 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9328) );
  AOI22_X1 U10550 ( .A1(n4870), .A2(keyinput49), .B1(keyinput4), .B2(n9328), 
        .ZN(n9327) );
  OAI221_X1 U10551 ( .B1(n4870), .B2(keyinput49), .C1(n9328), .C2(keyinput4), 
        .A(n9327), .ZN(n9333) );
  AOI22_X1 U10552 ( .A1(n9331), .A2(keyinput59), .B1(keyinput29), .B2(n9330), 
        .ZN(n9329) );
  OAI221_X1 U10553 ( .B1(n9331), .B2(keyinput59), .C1(n9330), .C2(keyinput29), 
        .A(n9329), .ZN(n9332) );
  NOR3_X1 U10554 ( .A1(n9334), .A2(n9333), .A3(n9332), .ZN(n9348) );
  INV_X1 U10555 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n9854) );
  INV_X1 U10556 ( .A(keyinput63), .ZN(n9336) );
  AOI22_X1 U10557 ( .A1(n9854), .A2(keyinput17), .B1(P1_ADDR_REG_2__SCAN_IN), 
        .B2(n9336), .ZN(n9335) );
  OAI221_X1 U10558 ( .B1(n9854), .B2(keyinput17), .C1(n9336), .C2(
        P1_ADDR_REG_2__SCAN_IN), .A(n9335), .ZN(n9340) );
  INV_X1 U10559 ( .A(keyinput35), .ZN(n9338) );
  AOI22_X1 U10560 ( .A1(n9776), .A2(keyinput2), .B1(P2_ADDR_REG_18__SCAN_IN), 
        .B2(n9338), .ZN(n9337) );
  OAI221_X1 U10561 ( .B1(n9776), .B2(keyinput2), .C1(n9338), .C2(
        P2_ADDR_REG_18__SCAN_IN), .A(n9337), .ZN(n9339) );
  NOR2_X1 U10562 ( .A1(n9340), .A2(n9339), .ZN(n9347) );
  AOI22_X1 U10563 ( .A1(n9342), .A2(keyinput48), .B1(keyinput27), .B2(n6140), 
        .ZN(n9341) );
  OAI221_X1 U10564 ( .B1(n9342), .B2(keyinput48), .C1(n6140), .C2(keyinput27), 
        .A(n9341), .ZN(n9345) );
  AOI22_X1 U10565 ( .A1(n6645), .A2(keyinput14), .B1(n6999), .B2(keyinput8), 
        .ZN(n9343) );
  OAI221_X1 U10566 ( .B1(n6645), .B2(keyinput14), .C1(n6999), .C2(keyinput8), 
        .A(n9343), .ZN(n9344) );
  NOR2_X1 U10567 ( .A1(n9345), .A2(n9344), .ZN(n9346) );
  NAND4_X1 U10568 ( .A1(n9349), .A2(n9348), .A3(n9347), .A4(n9346), .ZN(n9350)
         );
  NOR3_X1 U10569 ( .A1(n9352), .A2(n9351), .A3(n9350), .ZN(n9391) );
  INV_X1 U10570 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n9853) );
  INV_X1 U10571 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9354) );
  AOI22_X1 U10572 ( .A1(n9853), .A2(keyinput23), .B1(n9354), .B2(keyinput10), 
        .ZN(n9353) );
  OAI221_X1 U10573 ( .B1(n9853), .B2(keyinput23), .C1(n9354), .C2(keyinput10), 
        .A(n9353), .ZN(n9366) );
  AOI22_X1 U10574 ( .A1(n9357), .A2(keyinput43), .B1(keyinput58), .B2(n9356), 
        .ZN(n9355) );
  OAI221_X1 U10575 ( .B1(n9357), .B2(keyinput43), .C1(n9356), .C2(keyinput58), 
        .A(n9355), .ZN(n9365) );
  AOI22_X1 U10576 ( .A1(n9360), .A2(keyinput44), .B1(n9359), .B2(keyinput34), 
        .ZN(n9358) );
  OAI221_X1 U10577 ( .B1(n9360), .B2(keyinput44), .C1(n9359), .C2(keyinput34), 
        .A(n9358), .ZN(n9364) );
  AOI22_X1 U10578 ( .A1(n9362), .A2(keyinput56), .B1(keyinput55), .B2(n8139), 
        .ZN(n9361) );
  OAI221_X1 U10579 ( .B1(n9362), .B2(keyinput56), .C1(n8139), .C2(keyinput55), 
        .A(n9361), .ZN(n9363) );
  NOR4_X1 U10580 ( .A1(n9366), .A2(n9365), .A3(n9364), .A4(n9363), .ZN(n9390)
         );
  AOI22_X1 U10581 ( .A1(n5997), .A2(keyinput9), .B1(keyinput46), .B2(n5456), 
        .ZN(n9367) );
  OAI221_X1 U10582 ( .B1(n5997), .B2(keyinput9), .C1(n5456), .C2(keyinput46), 
        .A(n9367), .ZN(n9375) );
  AOI22_X1 U10583 ( .A1(n9369), .A2(keyinput3), .B1(n9714), .B2(keyinput52), 
        .ZN(n9368) );
  OAI221_X1 U10584 ( .B1(n9369), .B2(keyinput3), .C1(n9714), .C2(keyinput52), 
        .A(n9368), .ZN(n9374) );
  AOI22_X1 U10585 ( .A1(P1_U3084), .A2(keyinput15), .B1(keyinput30), .B2(n9436), .ZN(n9370) );
  OAI221_X1 U10586 ( .B1(P1_U3084), .B2(keyinput15), .C1(n9436), .C2(
        keyinput30), .A(n9370), .ZN(n9373) );
  AOI22_X1 U10587 ( .A1(n9472), .A2(keyinput51), .B1(n9721), .B2(keyinput22), 
        .ZN(n9371) );
  OAI221_X1 U10588 ( .B1(n9472), .B2(keyinput51), .C1(n9721), .C2(keyinput22), 
        .A(n9371), .ZN(n9372) );
  NOR4_X1 U10589 ( .A1(n9375), .A2(n9374), .A3(n9373), .A4(n9372), .ZN(n9389)
         );
  AOI22_X1 U10590 ( .A1(n5081), .A2(keyinput61), .B1(n9715), .B2(keyinput21), 
        .ZN(n9376) );
  OAI221_X1 U10591 ( .B1(n5081), .B2(keyinput61), .C1(n9715), .C2(keyinput21), 
        .A(n9376), .ZN(n9387) );
  INV_X1 U10592 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n9855) );
  AOI22_X1 U10593 ( .A1(n6732), .A2(keyinput25), .B1(n9855), .B2(keyinput26), 
        .ZN(n9377) );
  OAI221_X1 U10594 ( .B1(n6732), .B2(keyinput25), .C1(n9855), .C2(keyinput26), 
        .A(n9377), .ZN(n9386) );
  AOI22_X1 U10595 ( .A1(n9380), .A2(keyinput24), .B1(keyinput0), .B2(n9379), 
        .ZN(n9378) );
  OAI221_X1 U10596 ( .B1(n9380), .B2(keyinput24), .C1(n9379), .C2(keyinput0), 
        .A(n9378), .ZN(n9385) );
  AOI22_X1 U10597 ( .A1(n9383), .A2(keyinput1), .B1(keyinput54), .B2(n9382), 
        .ZN(n9381) );
  OAI221_X1 U10598 ( .B1(n9383), .B2(keyinput1), .C1(n9382), .C2(keyinput54), 
        .A(n9381), .ZN(n9384) );
  NOR4_X1 U10599 ( .A1(n9387), .A2(n9386), .A3(n9385), .A4(n9384), .ZN(n9388)
         );
  NAND4_X1 U10600 ( .A1(n9391), .A2(n9390), .A3(n9389), .A4(n9388), .ZN(n9392)
         );
  XNOR2_X1 U10601 ( .A(n9393), .B(n9392), .ZN(P1_U3515) );
  MUX2_X1 U10602 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9394), .S(n9767), .Z(
        P1_U3514) );
  MUX2_X1 U10603 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9395), .S(n9767), .Z(
        P1_U3513) );
  MUX2_X1 U10604 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9396), .S(n9767), .Z(
        P1_U3512) );
  MUX2_X1 U10605 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9397), .S(n9767), .Z(
        P1_U3511) );
  MUX2_X1 U10606 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9398), .S(n9767), .Z(
        P1_U3510) );
  MUX2_X1 U10607 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9399), .S(n9767), .Z(
        P1_U3508) );
  MUX2_X1 U10608 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9400), .S(n9767), .Z(
        P1_U3505) );
  MUX2_X1 U10609 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9401), .S(n9767), .Z(
        P1_U3499) );
  AND2_X1 U10610 ( .A1(n9403), .A2(n9402), .ZN(n9722) );
  MUX2_X1 U10611 ( .A(P1_D_REG_0__SCAN_IN), .B(n9404), .S(n9722), .Z(P1_U3440)
         );
  INV_X1 U10612 ( .A(n9405), .ZN(n9410) );
  NOR4_X1 U10613 ( .A1(n9407), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n9406), .ZN(n9408) );
  AOI21_X1 U10614 ( .B1(n9416), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9408), .ZN(
        n9409) );
  OAI21_X1 U10615 ( .B1(n9410), .B2(n6758), .A(n9409), .ZN(P1_U3322) );
  AOI22_X1 U10616 ( .A1(n4853), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n9416), .ZN(n9411) );
  OAI21_X1 U10617 ( .B1(n9412), .B2(n6758), .A(n9411), .ZN(P1_U3323) );
  AOI22_X1 U10618 ( .A1(n9413), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n9416), .ZN(n9414) );
  OAI21_X1 U10619 ( .B1(n9415), .B2(n6758), .A(n9414), .ZN(P1_U3324) );
  AOI22_X1 U10620 ( .A1(n9589), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n9416), .ZN(n9417) );
  OAI21_X1 U10621 ( .B1(n9418), .B2(n6758), .A(n9417), .ZN(P1_U3325) );
  MUX2_X1 U10622 ( .A(n9419), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI211_X1 U10623 ( .C1(n9422), .C2(n9421), .A(n9420), .B(n9575), .ZN(n9427)
         );
  AOI211_X1 U10624 ( .C1(n9425), .C2(n9424), .A(n9423), .B(n9626), .ZN(n9426)
         );
  AOI211_X1 U10625 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(P1_U3084), .A(n9427), 
        .B(n9426), .ZN(n9432) );
  INV_X1 U10626 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9429) );
  OAI22_X1 U10627 ( .A1(n9667), .A2(n9429), .B1(n9634), .B2(n9428), .ZN(n9430)
         );
  INV_X1 U10628 ( .A(n9430), .ZN(n9431) );
  NAND2_X1 U10629 ( .A1(n9432), .A2(n9431), .ZN(P1_U3244) );
  AOI21_X1 U10630 ( .B1(n9435), .B2(n9434), .A(n9433), .ZN(n9439) );
  OAI22_X1 U10631 ( .A1(n9437), .A2(n9957), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9436), .ZN(n9438) );
  AOI21_X1 U10632 ( .B1(n9787), .B2(n9439), .A(n9438), .ZN(n9442) );
  NAND2_X1 U10633 ( .A1(n9454), .A2(n9440), .ZN(n9441) );
  AND2_X1 U10634 ( .A1(n9442), .A2(n9441), .ZN(n9447) );
  INV_X1 U10635 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9796) );
  NOR2_X1 U10636 ( .A1(n9796), .A2(n9785), .ZN(n9445) );
  OAI211_X1 U10637 ( .C1(n9445), .C2(n9444), .A(n9784), .B(n9443), .ZN(n9446)
         );
  NAND2_X1 U10638 ( .A1(n9447), .A2(n9446), .ZN(P2_U3246) );
  AOI22_X1 U10639 ( .A1(n9793), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9460) );
  AOI211_X1 U10640 ( .C1(n9451), .C2(n9450), .A(n9449), .B(n9448), .ZN(n9452)
         );
  AOI21_X1 U10641 ( .B1(n9454), .B2(n9453), .A(n9452), .ZN(n9459) );
  OAI211_X1 U10642 ( .C1(n9457), .C2(n9456), .A(n9784), .B(n9455), .ZN(n9458)
         );
  NAND3_X1 U10643 ( .A1(n9460), .A2(n9459), .A3(n9458), .ZN(P2_U3247) );
  OAI211_X1 U10644 ( .C1(n9463), .C2(n9919), .A(n9462), .B(n9461), .ZN(n9464)
         );
  AOI21_X1 U10645 ( .B1(n9465), .B2(n9933), .A(n9464), .ZN(n9480) );
  AOI22_X1 U10646 ( .A1(n9952), .A2(n9480), .B1(n9466), .B2(n9950), .ZN(
        P2_U3535) );
  OAI22_X1 U10647 ( .A1(n9468), .A2(n9921), .B1(n9467), .B2(n9919), .ZN(n9469)
         );
  AOI211_X1 U10648 ( .C1(n9471), .C2(n9933), .A(n9470), .B(n9469), .ZN(n9482)
         );
  AOI22_X1 U10649 ( .A1(n9952), .A2(n9482), .B1(n9472), .B2(n9950), .ZN(
        P2_U3534) );
  INV_X1 U10650 ( .A(n9473), .ZN(n9913) );
  OAI22_X1 U10651 ( .A1(n9474), .A2(n9921), .B1(n4598), .B2(n9919), .ZN(n9476)
         );
  AOI211_X1 U10652 ( .C1(n9913), .C2(n9477), .A(n9476), .B(n9475), .ZN(n9484)
         );
  AOI22_X1 U10653 ( .A1(n9952), .A2(n9484), .B1(n9478), .B2(n9950), .ZN(
        P2_U3533) );
  INV_X1 U10654 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9479) );
  AOI22_X1 U10655 ( .A1(n9937), .A2(n9480), .B1(n9479), .B2(n9935), .ZN(
        P2_U3496) );
  INV_X1 U10656 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9481) );
  AOI22_X1 U10657 ( .A1(n9937), .A2(n9482), .B1(n9481), .B2(n9935), .ZN(
        P2_U3493) );
  INV_X1 U10658 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9483) );
  AOI22_X1 U10659 ( .A1(n9937), .A2(n9484), .B1(n9483), .B2(n9935), .ZN(
        P2_U3490) );
  XNOR2_X1 U10660 ( .A(n9485), .B(n4534), .ZN(n9499) );
  INV_X1 U10661 ( .A(n9499), .ZN(n9545) );
  INV_X1 U10662 ( .A(n9486), .ZN(n9541) );
  INV_X1 U10663 ( .A(n9487), .ZN(n9490) );
  INV_X1 U10664 ( .A(n9488), .ZN(n9489) );
  OAI21_X1 U10665 ( .B1(n9541), .B2(n9490), .A(n9489), .ZN(n9542) );
  INV_X1 U10666 ( .A(n9542), .ZN(n9491) );
  AOI22_X1 U10667 ( .A1(n9545), .A2(n9693), .B1(n9692), .B2(n9491), .ZN(n9504)
         );
  OAI21_X1 U10668 ( .B1(n9494), .B2(n9493), .A(n9492), .ZN(n9497) );
  OAI22_X1 U10669 ( .A1(n9511), .A2(n9696), .B1(n9495), .B2(n9698), .ZN(n9496)
         );
  AOI21_X1 U10670 ( .B1(n9497), .B2(n9701), .A(n9496), .ZN(n9498) );
  OAI21_X1 U10671 ( .B1(n9499), .B2(n9704), .A(n9498), .ZN(n9543) );
  AOI22_X1 U10672 ( .A1(n9517), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9500), .B2(
        n9707), .ZN(n9501) );
  OAI21_X1 U10673 ( .B1(n9541), .B2(n9710), .A(n9501), .ZN(n9502) );
  AOI21_X1 U10674 ( .B1(n9543), .B2(n9684), .A(n9502), .ZN(n9503) );
  NAND2_X1 U10675 ( .A1(n9504), .A2(n9503), .ZN(P1_U3278) );
  XNOR2_X1 U10676 ( .A(n9505), .B(n9509), .ZN(n9515) );
  INV_X1 U10677 ( .A(n9515), .ZN(n9556) );
  OAI21_X1 U10678 ( .B1(n9507), .B2(n9552), .A(n9506), .ZN(n9553) );
  INV_X1 U10679 ( .A(n9553), .ZN(n9508) );
  AOI22_X1 U10680 ( .A1(n9556), .A2(n9693), .B1(n9692), .B2(n9508), .ZN(n9521)
         );
  XNOR2_X1 U10681 ( .A(n9510), .B(n9509), .ZN(n9513) );
  OAI22_X1 U10682 ( .A1(n9675), .A2(n9696), .B1(n9511), .B2(n9698), .ZN(n9512)
         );
  AOI21_X1 U10683 ( .B1(n9513), .B2(n9701), .A(n9512), .ZN(n9514) );
  OAI21_X1 U10684 ( .B1(n9515), .B2(n9704), .A(n9514), .ZN(n9554) );
  AOI22_X1 U10685 ( .A1(n9517), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n9516), .B2(
        n9707), .ZN(n9518) );
  OAI21_X1 U10686 ( .B1(n9552), .B2(n9710), .A(n9518), .ZN(n9519) );
  AOI21_X1 U10687 ( .B1(n9554), .B2(n9684), .A(n9519), .ZN(n9520) );
  NAND2_X1 U10688 ( .A1(n9521), .A2(n9520), .ZN(P1_U3280) );
  OAI21_X1 U10689 ( .B1(n9523), .B2(n9759), .A(n9522), .ZN(n9524) );
  AOI21_X1 U10690 ( .B1(n9526), .B2(n9525), .A(n9524), .ZN(n9558) );
  INV_X1 U10691 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9527) );
  AOI22_X1 U10692 ( .A1(n9783), .A2(n9558), .B1(n9527), .B2(n9780), .ZN(
        P1_U3553) );
  INV_X1 U10693 ( .A(n9528), .ZN(n9534) );
  INV_X1 U10694 ( .A(n9529), .ZN(n9758) );
  OAI21_X1 U10695 ( .B1(n9531), .B2(n9759), .A(n9530), .ZN(n9533) );
  AOI211_X1 U10696 ( .C1(n9534), .C2(n9758), .A(n9533), .B(n9532), .ZN(n9559)
         );
  AOI22_X1 U10697 ( .A1(n9783), .A2(n9559), .B1(n8908), .B2(n9780), .ZN(
        P1_U3539) );
  OAI21_X1 U10698 ( .B1(n9536), .B2(n9759), .A(n9535), .ZN(n9538) );
  AOI211_X1 U10699 ( .C1(n9539), .C2(n9758), .A(n9538), .B(n9537), .ZN(n9560)
         );
  AOI22_X1 U10700 ( .A1(n9783), .A2(n9560), .B1(n9540), .B2(n9780), .ZN(
        P1_U3537) );
  OAI22_X1 U10701 ( .A1(n9542), .A2(n9761), .B1(n9541), .B2(n9759), .ZN(n9544)
         );
  AOI211_X1 U10702 ( .C1(n9766), .C2(n9545), .A(n9544), .B(n9543), .ZN(n9561)
         );
  AOI22_X1 U10703 ( .A1(n9783), .A2(n9561), .B1(n7522), .B2(n9780), .ZN(
        P1_U3536) );
  INV_X1 U10704 ( .A(n9546), .ZN(n9551) );
  OAI21_X1 U10705 ( .B1(n9548), .B2(n9759), .A(n9547), .ZN(n9550) );
  AOI211_X1 U10706 ( .C1(n9766), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9562)
         );
  AOI22_X1 U10707 ( .A1(n9783), .A2(n9562), .B1(n6990), .B2(n9780), .ZN(
        P1_U3535) );
  OAI22_X1 U10708 ( .A1(n9553), .A2(n9761), .B1(n9552), .B2(n9759), .ZN(n9555)
         );
  AOI211_X1 U10709 ( .C1(n9766), .C2(n9556), .A(n9555), .B(n9554), .ZN(n9563)
         );
  AOI22_X1 U10710 ( .A1(n9783), .A2(n9563), .B1(n9557), .B2(n9780), .ZN(
        P1_U3534) );
  AOI22_X1 U10711 ( .A1(n9767), .A2(n9558), .B1(n5453), .B2(n4495), .ZN(
        P1_U3521) );
  AOI22_X1 U10712 ( .A1(n9767), .A2(n9559), .B1(n5197), .B2(n4495), .ZN(
        P1_U3502) );
  AOI22_X1 U10713 ( .A1(n9767), .A2(n9560), .B1(n5148), .B2(n4495), .ZN(
        P1_U3496) );
  AOI22_X1 U10714 ( .A1(n9767), .A2(n9561), .B1(n5128), .B2(n4495), .ZN(
        P1_U3493) );
  AOI22_X1 U10715 ( .A1(n9767), .A2(n9562), .B1(n5107), .B2(n4495), .ZN(
        P1_U3490) );
  AOI22_X1 U10716 ( .A1(n9767), .A2(n9563), .B1(n5084), .B2(n4495), .ZN(
        P1_U3487) );
  XNOR2_X1 U10717 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10718 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10719 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9564) );
  OAI22_X1 U10720 ( .A1(n9667), .A2(n9564), .B1(n9634), .B2(n4502), .ZN(n9565)
         );
  INV_X1 U10721 ( .A(n9565), .ZN(n9574) );
  NAND2_X1 U10722 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9568) );
  AOI211_X1 U10723 ( .C1(n9568), .C2(n9567), .A(n9566), .B(n9575), .ZN(n9572)
         );
  AOI211_X1 U10724 ( .C1(n9583), .C2(n9570), .A(n9569), .B(n9626), .ZN(n9571)
         );
  AOI211_X1 U10725 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9572), 
        .B(n9571), .ZN(n9573) );
  NAND2_X1 U10726 ( .A1(n9574), .A2(n9573), .ZN(P1_U3242) );
  AOI211_X1 U10727 ( .C1(n9578), .C2(n9577), .A(n9576), .B(n9575), .ZN(n9579)
         );
  AOI21_X1 U10728 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n9579), 
        .ZN(n9594) );
  AOI211_X1 U10729 ( .C1(n9582), .C2(n9581), .A(n9580), .B(n9626), .ZN(n9591)
         );
  INV_X1 U10730 ( .A(n9583), .ZN(n9586) );
  MUX2_X1 U10731 ( .A(n9586), .B(n9585), .S(n9584), .Z(n9590) );
  AOI211_X1 U10732 ( .C1(n9590), .C2(n9589), .A(n9588), .B(n9587), .ZN(n9604)
         );
  AOI211_X1 U10733 ( .C1(n9654), .C2(n9592), .A(n9591), .B(n9604), .ZN(n9593)
         );
  OAI211_X1 U10734 ( .C1(n9595), .C2(n9667), .A(n9594), .B(n9593), .ZN(
        P1_U3243) );
  OAI21_X1 U10735 ( .B1(n9598), .B2(n9597), .A(n9596), .ZN(n9599) );
  AOI22_X1 U10736 ( .A1(n9600), .A2(n9654), .B1(n9662), .B2(n9599), .ZN(n9608)
         );
  OAI21_X1 U10737 ( .B1(n9603), .B2(n9602), .A(n9601), .ZN(n9606) );
  NOR2_X1 U10738 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6861), .ZN(n9605) );
  AOI211_X1 U10739 ( .C1(n9661), .C2(n9606), .A(n9605), .B(n9604), .ZN(n9607)
         );
  OAI211_X1 U10740 ( .C1(n9667), .C2(n9609), .A(n9608), .B(n9607), .ZN(
        P1_U3245) );
  OAI21_X1 U10741 ( .B1(n9612), .B2(n9611), .A(n9610), .ZN(n9615) );
  INV_X1 U10742 ( .A(n9613), .ZN(n9614) );
  AOI21_X1 U10743 ( .B1(n9615), .B2(n9661), .A(n9614), .ZN(n9622) );
  AOI211_X1 U10744 ( .C1(n9618), .C2(n9617), .A(n9616), .B(n9626), .ZN(n9619)
         );
  AOI21_X1 U10745 ( .B1(n9654), .B2(n9620), .A(n9619), .ZN(n9621) );
  OAI211_X1 U10746 ( .C1(n9667), .C2(n9992), .A(n9622), .B(n9621), .ZN(
        P1_U3250) );
  OAI21_X1 U10747 ( .B1(n9625), .B2(n9624), .A(n9623), .ZN(n9632) );
  AOI211_X1 U10748 ( .C1(n9629), .C2(n9628), .A(n9627), .B(n9626), .ZN(n9630)
         );
  AOI211_X1 U10749 ( .C1(n9632), .C2(n9661), .A(n9631), .B(n9630), .ZN(n9638)
         );
  INV_X1 U10750 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9635) );
  OAI22_X1 U10751 ( .A1(n9667), .A2(n9635), .B1(n9634), .B2(n9633), .ZN(n9636)
         );
  INV_X1 U10752 ( .A(n9636), .ZN(n9637) );
  NAND2_X1 U10753 ( .A1(n9638), .A2(n9637), .ZN(P1_U3251) );
  INV_X1 U10754 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9651) );
  AOI21_X1 U10755 ( .B1(n9654), .B2(n9640), .A(n9639), .ZN(n9650) );
  OAI21_X1 U10756 ( .B1(n9643), .B2(n9642), .A(n9641), .ZN(n9648) );
  OAI21_X1 U10757 ( .B1(n9646), .B2(n9645), .A(n9644), .ZN(n9647) );
  AOI22_X1 U10758 ( .A1(n9648), .A2(n9661), .B1(n9647), .B2(n9662), .ZN(n9649)
         );
  OAI211_X1 U10759 ( .C1(n9667), .C2(n9651), .A(n9650), .B(n9649), .ZN(
        P1_U3252) );
  INV_X1 U10760 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9666) );
  AOI21_X1 U10761 ( .B1(n9654), .B2(n9653), .A(n9652), .ZN(n9665) );
  OAI21_X1 U10762 ( .B1(n9656), .B2(n7539), .A(n9655), .ZN(n9663) );
  OAI21_X1 U10763 ( .B1(n9659), .B2(n9658), .A(n9657), .ZN(n9660) );
  AOI22_X1 U10764 ( .A1(n9663), .A2(n9662), .B1(n9661), .B2(n9660), .ZN(n9664)
         );
  OAI211_X1 U10765 ( .C1(n9667), .C2(n9666), .A(n9665), .B(n9664), .ZN(
        P1_U3255) );
  XOR2_X1 U10766 ( .A(n9668), .B(n9674), .Z(n9680) );
  INV_X1 U10767 ( .A(n9680), .ZN(n9765) );
  NOR2_X1 U10768 ( .A1(n9669), .A2(n9760), .ZN(n9670) );
  OR2_X1 U10769 ( .A1(n9671), .A2(n9670), .ZN(n9762) );
  INV_X1 U10770 ( .A(n9762), .ZN(n9672) );
  AOI22_X1 U10771 ( .A1(n9765), .A2(n9693), .B1(n9692), .B2(n9672), .ZN(n9686)
         );
  XOR2_X1 U10772 ( .A(n9674), .B(n9673), .Z(n9678) );
  OAI22_X1 U10773 ( .A1(n9676), .A2(n9696), .B1(n9675), .B2(n9698), .ZN(n9677)
         );
  AOI21_X1 U10774 ( .B1(n9678), .B2(n9701), .A(n9677), .ZN(n9679) );
  OAI21_X1 U10775 ( .B1(n9680), .B2(n9704), .A(n9679), .ZN(n9763) );
  AOI22_X1 U10776 ( .A1(n9708), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n9681), .B2(
        n9707), .ZN(n9682) );
  OAI21_X1 U10777 ( .B1(n9760), .B2(n9710), .A(n9682), .ZN(n9683) );
  AOI21_X1 U10778 ( .B1(n9763), .B2(n9684), .A(n9683), .ZN(n9685) );
  NAND2_X1 U10779 ( .A1(n9686), .A2(n9685), .ZN(P1_U3282) );
  XOR2_X1 U10780 ( .A(n9694), .B(n9687), .Z(n9705) );
  INV_X1 U10781 ( .A(n9705), .ZN(n9734) );
  INV_X1 U10782 ( .A(n9688), .ZN(n9690) );
  OAI21_X1 U10783 ( .B1(n9690), .B2(n9730), .A(n9689), .ZN(n9731) );
  INV_X1 U10784 ( .A(n9731), .ZN(n9691) );
  AOI22_X1 U10785 ( .A1(n9734), .A2(n9693), .B1(n9692), .B2(n9691), .ZN(n9713)
         );
  XNOR2_X1 U10786 ( .A(n9695), .B(n9694), .ZN(n9702) );
  OAI22_X1 U10787 ( .A1(n9699), .A2(n9698), .B1(n9697), .B2(n9696), .ZN(n9700)
         );
  AOI21_X1 U10788 ( .B1(n9702), .B2(n9701), .A(n9700), .ZN(n9703) );
  OAI21_X1 U10789 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9732) );
  AOI22_X1 U10790 ( .A1(n9708), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9707), .B2(
        n9706), .ZN(n9709) );
  OAI21_X1 U10791 ( .B1(n9730), .B2(n9710), .A(n9709), .ZN(n9711) );
  AOI21_X1 U10792 ( .B1(n9732), .B2(n9684), .A(n9711), .ZN(n9712) );
  NAND2_X1 U10793 ( .A1(n9713), .A2(n9712), .ZN(P1_U3288) );
  AND2_X1 U10794 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9723), .ZN(P1_U3292) );
  AND2_X1 U10795 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9723), .ZN(P1_U3293) );
  AND2_X1 U10796 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9723), .ZN(P1_U3294) );
  AND2_X1 U10797 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9723), .ZN(P1_U3295) );
  AND2_X1 U10798 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9723), .ZN(P1_U3296) );
  NOR2_X1 U10799 ( .A1(n9722), .A2(n9714), .ZN(P1_U3297) );
  AND2_X1 U10800 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9723), .ZN(P1_U3298) );
  NOR2_X1 U10801 ( .A1(n9722), .A2(n9715), .ZN(P1_U3299) );
  AND2_X1 U10802 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9723), .ZN(P1_U3300) );
  NOR2_X1 U10803 ( .A1(n9722), .A2(n9716), .ZN(P1_U3301) );
  AND2_X1 U10804 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9723), .ZN(P1_U3302) );
  NOR2_X1 U10805 ( .A1(n9722), .A2(n9717), .ZN(P1_U3303) );
  AND2_X1 U10806 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9723), .ZN(P1_U3304) );
  AND2_X1 U10807 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9723), .ZN(P1_U3305) );
  NOR2_X1 U10808 ( .A1(n9722), .A2(n9718), .ZN(P1_U3306) );
  AND2_X1 U10809 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9723), .ZN(P1_U3307) );
  AND2_X1 U10810 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9723), .ZN(P1_U3308) );
  AND2_X1 U10811 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9723), .ZN(P1_U3309) );
  NOR2_X1 U10812 ( .A1(n9722), .A2(n9719), .ZN(P1_U3310) );
  AND2_X1 U10813 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9723), .ZN(P1_U3311) );
  NOR2_X1 U10814 ( .A1(n9722), .A2(n9720), .ZN(P1_U3312) );
  AND2_X1 U10815 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9723), .ZN(P1_U3313) );
  NOR2_X1 U10816 ( .A1(n9722), .A2(n9721), .ZN(P1_U3314) );
  AND2_X1 U10817 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9723), .ZN(P1_U3315) );
  AND2_X1 U10818 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9723), .ZN(P1_U3316) );
  AND2_X1 U10819 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9723), .ZN(P1_U3317) );
  AND2_X1 U10820 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9723), .ZN(P1_U3318) );
  AND2_X1 U10821 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9723), .ZN(P1_U3319) );
  AND2_X1 U10822 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9723), .ZN(P1_U3320) );
  AND2_X1 U10823 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9723), .ZN(P1_U3321) );
  OAI22_X1 U10824 ( .A1(n9725), .A2(n9761), .B1(n9724), .B2(n9759), .ZN(n9726)
         );
  AOI21_X1 U10825 ( .B1(n9727), .B2(n9766), .A(n9726), .ZN(n9728) );
  AND2_X1 U10826 ( .A1(n9729), .A2(n9728), .ZN(n9769) );
  AOI22_X1 U10827 ( .A1(n9767), .A2(n9769), .B1(n4855), .B2(n4495), .ZN(
        P1_U3460) );
  OAI22_X1 U10828 ( .A1(n9731), .A2(n9761), .B1(n9730), .B2(n9759), .ZN(n9733)
         );
  AOI211_X1 U10829 ( .C1(n9766), .C2(n9734), .A(n9733), .B(n9732), .ZN(n9771)
         );
  AOI22_X1 U10830 ( .A1(n9767), .A2(n9771), .B1(n4900), .B2(n4495), .ZN(
        P1_U3463) );
  OAI22_X1 U10831 ( .A1(n9736), .A2(n9761), .B1(n9735), .B2(n9759), .ZN(n9738)
         );
  AOI211_X1 U10832 ( .C1(n9758), .C2(n9739), .A(n9738), .B(n9737), .ZN(n9773)
         );
  INV_X1 U10833 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9740) );
  AOI22_X1 U10834 ( .A1(n9767), .A2(n9773), .B1(n9740), .B2(n4495), .ZN(
        P1_U3466) );
  NAND3_X1 U10835 ( .A1(n9742), .A2(n9741), .A3(n9758), .ZN(n9744) );
  OAI211_X1 U10836 ( .C1(n9745), .C2(n9759), .A(n9744), .B(n9743), .ZN(n9746)
         );
  NOR2_X1 U10837 ( .A1(n9747), .A2(n9746), .ZN(n9775) );
  AOI22_X1 U10838 ( .A1(n9767), .A2(n9775), .B1(n4941), .B2(n4495), .ZN(
        P1_U3469) );
  OAI22_X1 U10839 ( .A1(n9749), .A2(n9761), .B1(n9748), .B2(n9759), .ZN(n9751)
         );
  AOI211_X1 U10840 ( .C1(n9766), .C2(n9752), .A(n9751), .B(n9750), .ZN(n9777)
         );
  AOI22_X1 U10841 ( .A1(n9767), .A2(n9777), .B1(n4962), .B2(n4495), .ZN(
        P1_U3472) );
  OAI211_X1 U10842 ( .C1(n9755), .C2(n9759), .A(n9754), .B(n9753), .ZN(n9756)
         );
  AOI21_X1 U10843 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9779) );
  AOI22_X1 U10844 ( .A1(n9767), .A2(n9779), .B1(n5000), .B2(n4495), .ZN(
        P1_U3475) );
  OAI22_X1 U10845 ( .A1(n9762), .A2(n9761), .B1(n9760), .B2(n9759), .ZN(n9764)
         );
  AOI211_X1 U10846 ( .C1(n9766), .C2(n9765), .A(n9764), .B(n9763), .ZN(n9782)
         );
  AOI22_X1 U10847 ( .A1(n9767), .A2(n9782), .B1(n5044), .B2(n4495), .ZN(
        P1_U3481) );
  INV_X1 U10848 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U10849 ( .A1(n9783), .A2(n9769), .B1(n9768), .B2(n9780), .ZN(
        P1_U3525) );
  INV_X1 U10850 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9770) );
  AOI22_X1 U10851 ( .A1(n9783), .A2(n9771), .B1(n9770), .B2(n9780), .ZN(
        P1_U3526) );
  INV_X1 U10852 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9772) );
  AOI22_X1 U10853 ( .A1(n9783), .A2(n9773), .B1(n9772), .B2(n9780), .ZN(
        P1_U3527) );
  INV_X1 U10854 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9774) );
  AOI22_X1 U10855 ( .A1(n9783), .A2(n9775), .B1(n9774), .B2(n9780), .ZN(
        P1_U3528) );
  AOI22_X1 U10856 ( .A1(n9783), .A2(n9777), .B1(n9776), .B2(n9780), .ZN(
        P1_U3529) );
  INV_X1 U10857 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9778) );
  AOI22_X1 U10858 ( .A1(n9783), .A2(n9779), .B1(n9778), .B2(n9780), .ZN(
        P1_U3530) );
  INV_X1 U10859 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9781) );
  AOI22_X1 U10860 ( .A1(n9783), .A2(n9782), .B1(n9781), .B2(n9780), .ZN(
        P1_U3532) );
  AOI22_X1 U10861 ( .A1(n9784), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9787), .ZN(n9797) );
  INV_X1 U10862 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9786) );
  NAND2_X1 U10863 ( .A1(n9787), .A2(n9786), .ZN(n9788) );
  OAI211_X1 U10864 ( .C1(n9790), .C2(P2_REG2_REG_0__SCAN_IN), .A(n9789), .B(
        n9788), .ZN(n9791) );
  INV_X1 U10865 ( .A(n9791), .ZN(n9795) );
  AOI22_X1 U10866 ( .A1(n9793), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n9794) );
  OAI221_X1 U10867 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n9797), .C1(n9796), .C2(
        n9795), .A(n9794), .ZN(P2_U3245) );
  NAND2_X1 U10868 ( .A1(n9799), .A2(n9798), .ZN(n9800) );
  XNOR2_X1 U10869 ( .A(n9800), .B(n9804), .ZN(n9802) );
  AOI21_X1 U10870 ( .B1(n9802), .B2(n9830), .A(n9801), .ZN(n9931) );
  AOI222_X1 U10871 ( .A1(n9928), .A2(n9841), .B1(P2_REG2_REG_12__SCAN_IN), 
        .B2(n9840), .C1(n9839), .C2(n9803), .ZN(n9813) );
  OAI21_X1 U10872 ( .B1(n9806), .B2(n7592), .A(n9805), .ZN(n9934) );
  AOI21_X1 U10873 ( .B1(n9807), .B2(n9928), .A(n9921), .ZN(n9809) );
  NAND2_X1 U10874 ( .A1(n9809), .A2(n9808), .ZN(n9929) );
  INV_X1 U10875 ( .A(n9929), .ZN(n9810) );
  AOI22_X1 U10876 ( .A1(n9934), .A2(n9838), .B1(n9811), .B2(n9810), .ZN(n9812)
         );
  OAI211_X1 U10877 ( .C1(n9840), .C2(n9931), .A(n9813), .B(n9812), .ZN(
        P2_U3284) );
  OAI22_X1 U10878 ( .A1(n9815), .A2(n6724), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9814), .ZN(n9822) );
  INV_X1 U10879 ( .A(n9816), .ZN(n9820) );
  OAI22_X1 U10880 ( .A1(n9820), .A2(n9819), .B1(n9818), .B2(n9817), .ZN(n9821)
         );
  AOI211_X1 U10881 ( .C1(n9824), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9825)
         );
  OAI21_X1 U10882 ( .B1(n9840), .B2(n9826), .A(n9825), .ZN(P2_U3293) );
  INV_X1 U10883 ( .A(n6297), .ZN(n9831) );
  INV_X1 U10884 ( .A(n9827), .ZN(n9828) );
  NAND2_X1 U10885 ( .A1(n6801), .A2(n9828), .ZN(n9829) );
  OAI211_X1 U10886 ( .C1(n9832), .C2(n9831), .A(n9830), .B(n9829), .ZN(n9834)
         );
  AND2_X1 U10887 ( .A1(n9834), .A2(n9833), .ZN(n9875) );
  OR2_X1 U10888 ( .A1(n6801), .A2(n9835), .ZN(n9836) );
  NAND2_X1 U10889 ( .A1(n9837), .A2(n9836), .ZN(n9873) );
  NAND2_X1 U10890 ( .A1(n9838), .A2(n9873), .ZN(n9849) );
  AOI22_X1 U10891 ( .A1(n9840), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n9839), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n9848) );
  NAND2_X1 U10892 ( .A1(n9841), .A2(n6114), .ZN(n9847) );
  NAND2_X1 U10893 ( .A1(n6114), .A2(n9865), .ZN(n9842) );
  NAND2_X1 U10894 ( .A1(n9843), .A2(n9842), .ZN(n9871) );
  INV_X1 U10895 ( .A(n9871), .ZN(n9844) );
  NAND2_X1 U10896 ( .A1(n9845), .A2(n9844), .ZN(n9846) );
  AND4_X1 U10897 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(n9850)
         );
  OAI21_X1 U10898 ( .B1(n8495), .B2(n9875), .A(n9850), .ZN(P2_U3295) );
  NAND2_X1 U10899 ( .A1(n9852), .A2(n9851), .ZN(n9861) );
  AND2_X1 U10900 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n9861), .ZN(P2_U3297) );
  INV_X1 U10901 ( .A(n9861), .ZN(n9859) );
  NOR2_X1 U10902 ( .A1(n9859), .A2(n9853), .ZN(P2_U3298) );
  AND2_X1 U10903 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n9861), .ZN(P2_U3299) );
  AND2_X1 U10904 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n9861), .ZN(P2_U3300) );
  AND2_X1 U10905 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n9861), .ZN(P2_U3301) );
  AND2_X1 U10906 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n9861), .ZN(P2_U3302) );
  AND2_X1 U10907 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n9861), .ZN(P2_U3303) );
  AND2_X1 U10908 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n9861), .ZN(P2_U3304) );
  AND2_X1 U10909 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n9861), .ZN(P2_U3305) );
  AND2_X1 U10910 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n9861), .ZN(P2_U3306) );
  AND2_X1 U10911 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n9861), .ZN(P2_U3307) );
  AND2_X1 U10912 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n9861), .ZN(P2_U3308) );
  AND2_X1 U10913 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n9861), .ZN(P2_U3309) );
  AND2_X1 U10914 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n9861), .ZN(P2_U3310) );
  AND2_X1 U10915 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n9861), .ZN(P2_U3311) );
  NOR2_X1 U10916 ( .A1(n9859), .A2(n9854), .ZN(P2_U3312) );
  AND2_X1 U10917 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n9861), .ZN(P2_U3313) );
  AND2_X1 U10918 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n9861), .ZN(P2_U3314) );
  NOR2_X1 U10919 ( .A1(n9859), .A2(n9855), .ZN(P2_U3315) );
  AND2_X1 U10920 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n9861), .ZN(P2_U3316) );
  AND2_X1 U10921 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n9861), .ZN(P2_U3317) );
  AND2_X1 U10922 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n9861), .ZN(P2_U3318) );
  AND2_X1 U10923 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n9861), .ZN(P2_U3319) );
  AND2_X1 U10924 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n9861), .ZN(P2_U3320) );
  AND2_X1 U10925 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n9861), .ZN(P2_U3321) );
  AND2_X1 U10926 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n9861), .ZN(P2_U3322) );
  AND2_X1 U10927 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n9861), .ZN(P2_U3323) );
  AND2_X1 U10928 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n9861), .ZN(P2_U3324) );
  AND2_X1 U10929 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n9861), .ZN(P2_U3325) );
  NOR2_X1 U10930 ( .A1(n9859), .A2(n9856), .ZN(P2_U3326) );
  OAI22_X1 U10931 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n9859), .B1(n9858), .B2(
        n9857), .ZN(n9860) );
  INV_X1 U10932 ( .A(n9860), .ZN(P2_U3437) );
  INV_X1 U10933 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9862) );
  AOI22_X1 U10934 ( .A1(n9864), .A2(n9863), .B1(n9862), .B2(n9861), .ZN(
        P2_U3438) );
  AOI22_X1 U10935 ( .A1(n9867), .A2(n9933), .B1(n9866), .B2(n9865), .ZN(n9868)
         );
  AND2_X1 U10936 ( .A1(n9869), .A2(n9868), .ZN(n9938) );
  INV_X1 U10937 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9870) );
  AOI22_X1 U10938 ( .A1(n9937), .A2(n9938), .B1(n9870), .B2(n9935), .ZN(
        P2_U3451) );
  OAI22_X1 U10939 ( .A1(n9871), .A2(n9921), .B1(n6759), .B2(n9919), .ZN(n9872)
         );
  AOI21_X1 U10940 ( .B1(n9873), .B2(n9933), .A(n9872), .ZN(n9874) );
  AND2_X1 U10941 ( .A1(n9875), .A2(n9874), .ZN(n9939) );
  INV_X1 U10942 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9876) );
  AOI22_X1 U10943 ( .A1(n9937), .A2(n9939), .B1(n9876), .B2(n9935), .ZN(
        P2_U3454) );
  OAI22_X1 U10944 ( .A1(n9878), .A2(n9921), .B1(n9877), .B2(n9919), .ZN(n9880)
         );
  AOI211_X1 U10945 ( .C1(n9933), .C2(n9881), .A(n9880), .B(n9879), .ZN(n9941)
         );
  INV_X1 U10946 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9882) );
  AOI22_X1 U10947 ( .A1(n9937), .A2(n9941), .B1(n9882), .B2(n9935), .ZN(
        P2_U3463) );
  AOI22_X1 U10948 ( .A1(n9884), .A2(n4341), .B1(n9927), .B2(n9883), .ZN(n9885)
         );
  OAI211_X1 U10949 ( .C1(n9888), .C2(n9887), .A(n9886), .B(n9885), .ZN(n9889)
         );
  INV_X1 U10950 ( .A(n9889), .ZN(n9943) );
  INV_X1 U10951 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9890) );
  AOI22_X1 U10952 ( .A1(n9937), .A2(n9943), .B1(n9890), .B2(n9935), .ZN(
        P2_U3469) );
  OAI211_X1 U10953 ( .C1(n9893), .C2(n9919), .A(n9892), .B(n9891), .ZN(n9894)
         );
  AOI21_X1 U10954 ( .B1(n9895), .B2(n9933), .A(n9894), .ZN(n9945) );
  INV_X1 U10955 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9896) );
  AOI22_X1 U10956 ( .A1(n9937), .A2(n9945), .B1(n9896), .B2(n9935), .ZN(
        P2_U3472) );
  OAI22_X1 U10957 ( .A1(n9897), .A2(n9921), .B1(n4606), .B2(n9919), .ZN(n9898)
         );
  AOI21_X1 U10958 ( .B1(n9899), .B2(n9913), .A(n9898), .ZN(n9900) );
  AND2_X1 U10959 ( .A1(n9901), .A2(n9900), .ZN(n9946) );
  INV_X1 U10960 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9902) );
  AOI22_X1 U10961 ( .A1(n9937), .A2(n9946), .B1(n9902), .B2(n9935), .ZN(
        P2_U3475) );
  OAI22_X1 U10962 ( .A1(n9904), .A2(n9921), .B1(n9903), .B2(n9919), .ZN(n9905)
         );
  AOI21_X1 U10963 ( .B1(n9906), .B2(n9913), .A(n9905), .ZN(n9907) );
  AND2_X1 U10964 ( .A1(n9908), .A2(n9907), .ZN(n9947) );
  INV_X1 U10965 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9909) );
  AOI22_X1 U10966 ( .A1(n9937), .A2(n9947), .B1(n9909), .B2(n9935), .ZN(
        P2_U3478) );
  OAI22_X1 U10967 ( .A1(n9911), .A2(n9921), .B1(n9910), .B2(n9919), .ZN(n9912)
         );
  AOI21_X1 U10968 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(n9915) );
  AND2_X1 U10969 ( .A1(n9916), .A2(n9915), .ZN(n9948) );
  INV_X1 U10970 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9917) );
  AOI22_X1 U10971 ( .A1(n9937), .A2(n9948), .B1(n9917), .B2(n9935), .ZN(
        P2_U3481) );
  INV_X1 U10972 ( .A(n9918), .ZN(n9925) );
  OAI22_X1 U10973 ( .A1(n9922), .A2(n9921), .B1(n9920), .B2(n9919), .ZN(n9924)
         );
  AOI211_X1 U10974 ( .C1(n9925), .C2(n9933), .A(n9924), .B(n9923), .ZN(n9949)
         );
  INV_X1 U10975 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9926) );
  AOI22_X1 U10976 ( .A1(n9937), .A2(n9949), .B1(n9926), .B2(n9935), .ZN(
        P2_U3484) );
  NAND2_X1 U10977 ( .A1(n9928), .A2(n9927), .ZN(n9930) );
  NAND3_X1 U10978 ( .A1(n9931), .A2(n9930), .A3(n9929), .ZN(n9932) );
  AOI21_X1 U10979 ( .B1(n9934), .B2(n9933), .A(n9932), .ZN(n9951) );
  INV_X1 U10980 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n9936) );
  AOI22_X1 U10981 ( .A1(n9937), .A2(n9951), .B1(n9936), .B2(n9935), .ZN(
        P2_U3487) );
  AOI22_X1 U10982 ( .A1(n9952), .A2(n9938), .B1(n9786), .B2(n9950), .ZN(
        P2_U3520) );
  AOI22_X1 U10983 ( .A1(n9952), .A2(n9939), .B1(n6712), .B2(n9950), .ZN(
        P2_U3521) );
  INV_X1 U10984 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n9940) );
  AOI22_X1 U10985 ( .A1(n9952), .A2(n9941), .B1(n9940), .B2(n9950), .ZN(
        P2_U3524) );
  INV_X1 U10986 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9942) );
  AOI22_X1 U10987 ( .A1(n9952), .A2(n9943), .B1(n9942), .B2(n9950), .ZN(
        P2_U3526) );
  INV_X1 U10988 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9944) );
  AOI22_X1 U10989 ( .A1(n9952), .A2(n9945), .B1(n9944), .B2(n9950), .ZN(
        P2_U3527) );
  AOI22_X1 U10990 ( .A1(n9952), .A2(n9946), .B1(n6896), .B2(n9950), .ZN(
        P2_U3528) );
  AOI22_X1 U10991 ( .A1(n9952), .A2(n9947), .B1(n6897), .B2(n9950), .ZN(
        P2_U3529) );
  AOI22_X1 U10992 ( .A1(n9952), .A2(n9948), .B1(n6898), .B2(n9950), .ZN(
        P2_U3530) );
  AOI22_X1 U10993 ( .A1(n9952), .A2(n9949), .B1(n6972), .B2(n9950), .ZN(
        P2_U3531) );
  AOI22_X1 U10994 ( .A1(n9952), .A2(n9951), .B1(n7142), .B2(n9950), .ZN(
        P2_U3532) );
  INV_X1 U10995 ( .A(n9953), .ZN(n9954) );
  NAND2_X1 U10996 ( .A1(n9955), .A2(n9954), .ZN(n9956) );
  XOR2_X1 U10997 ( .A(n9957), .B(n9956), .Z(ADD_1071_U5) );
  XOR2_X1 U10998 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U10999 ( .B1(n9960), .B2(n9959), .A(n9958), .ZN(ADD_1071_U56) );
  OAI21_X1 U11000 ( .B1(n9963), .B2(n9962), .A(n9961), .ZN(ADD_1071_U57) );
  OAI21_X1 U11001 ( .B1(n9966), .B2(n9965), .A(n9964), .ZN(ADD_1071_U58) );
  OAI21_X1 U11002 ( .B1(n9969), .B2(n9968), .A(n9967), .ZN(ADD_1071_U59) );
  OAI21_X1 U11003 ( .B1(n9972), .B2(n9971), .A(n9970), .ZN(ADD_1071_U60) );
  OAI21_X1 U11004 ( .B1(n9975), .B2(n9974), .A(n9973), .ZN(ADD_1071_U61) );
  AOI21_X1 U11005 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(ADD_1071_U62) );
  AOI21_X1 U11006 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(ADD_1071_U63) );
  XOR2_X1 U11007 ( .A(n9982), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11008 ( .A1(n9984), .A2(n9983), .ZN(n9985) );
  XOR2_X1 U11009 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n9985), .Z(ADD_1071_U51) );
  OAI21_X1 U11010 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n9989) );
  XNOR2_X1 U11011 ( .A(n9989), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11012 ( .B1(n9992), .B2(n9991), .A(n9990), .ZN(ADD_1071_U47) );
  XOR2_X1 U11013 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n9993), .Z(ADD_1071_U48) );
  XOR2_X1 U11014 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n9994), .Z(ADD_1071_U49) );
  XOR2_X1 U11015 ( .A(n9996), .B(n9995), .Z(ADD_1071_U54) );
  XOR2_X1 U11016 ( .A(n9998), .B(n9997), .Z(ADD_1071_U53) );
  XNOR2_X1 U11017 ( .A(n10000), .B(n9999), .ZN(ADD_1071_U52) );
  CLKBUF_X2 U4754 ( .A(n4672), .Z(n7684) );
  CLKBUF_X1 U4755 ( .A(n5623), .Z(n6151) );
  CLKBUF_X3 U4767 ( .A(n4934), .Z(n4267) );
endmodule

