

module b21_C_SARLock_k_128_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, ADD_1071_U4, ADD_1071_U55, 
        ADD_1071_U56, ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, 
        ADD_1071_U61, ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, 
        ADD_1071_U49, ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, 
        ADD_1071_U54, ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, 
        P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, 
        P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, 
        P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, 
        P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, 
        P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, 
        P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, 
        P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, 
        P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, 
        P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, 
        P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, 
        P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, 
        P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, 
        P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, 
        P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, 
        P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, 
        P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, 
        P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, 
        P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, 
        P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, 
        P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, 
        P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, 
        P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, 
        P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, 
        P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, 
        P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, 
        P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, 
        P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366;

  INV_X2 U4890 ( .A(n10222), .ZN(n10224) );
  NAND2_X1 U4891 ( .A1(n8695), .A2(n4401), .ZN(n8631) );
  NAND2_X2 U4892 ( .A1(n6062), .A2(n6061), .ZN(n8789) );
  INV_X1 U4893 ( .A(n8250), .ZN(n6013) );
  INV_X1 U4894 ( .A(n6286), .ZN(n6111) );
  CLKBUF_X2 U4896 ( .A(n5817), .Z(n8250) );
  INV_X2 U4897 ( .A(n6501), .ZN(n7634) );
  BUF_X1 U4898 ( .A(n5823), .Z(n4390) );
  NOR3_X1 U4899 ( .A1(n8724), .A2(n8704), .A3(n8703), .ZN(n8702) );
  OR2_X1 U4900 ( .A1(n6401), .A2(n6415), .ZN(n5041) );
  INV_X1 U4901 ( .A(n8138), .ZN(n6201) );
  OR2_X1 U4902 ( .A1(n8752), .A2(n8836), .ZN(n8754) );
  AND2_X1 U4903 ( .A1(n6969), .A2(n10275), .ZN(n6971) );
  OAI211_X1 U4904 ( .C1(n6401), .C2(n6414), .A(n5804), .B(n5803), .ZN(n6200)
         );
  OAI21_X1 U4905 ( .B1(n9161), .B2(n9162), .A(n5589), .ZN(n9139) );
  AOI21_X1 U4906 ( .B1(n8718), .B2(n8716), .A(n8717), .ZN(n8724) );
  INV_X1 U4907 ( .A(n5179), .ZN(n5136) );
  INV_X1 U4908 ( .A(n5485), .ZN(n5177) );
  CLKBUF_X2 U4909 ( .A(n5178), .Z(n6478) );
  NOR2_X1 U4910 ( .A1(n9408), .A2(n9168), .ZN(n9155) );
  NAND2_X1 U4911 ( .A1(n9225), .A2(n4777), .ZN(n9227) );
  MUX2_X1 U4912 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8889), .S(n6401), .Z(n10214)
         );
  NAND2_X1 U4913 ( .A1(n5814), .A2(n4428), .ZN(n8468) );
  XOR2_X1 U4914 ( .A(n6119), .B(n8385), .Z(n4384) );
  CLKBUF_X3 U4915 ( .A(n7679), .Z(n4386) );
  INV_X1 U4916 ( .A(n6501), .ZN(n4385) );
  NOR2_X2 U4917 ( .A1(n9266), .A2(n9439), .ZN(n9252) );
  AND2_X2 U4918 ( .A1(n5798), .A2(n5724), .ZN(n5828) );
  AND2_X1 U4919 ( .A1(n7501), .A2(n9810), .ZN(n7556) );
  NOR2_X2 U4920 ( .A1(n7499), .A2(n8850), .ZN(n7501) );
  AOI22_X2 U4921 ( .A1(n9215), .A2(n5715), .B1(n8924), .B2(n5714), .ZN(n9197)
         );
  NAND2_X2 U4922 ( .A1(n6023), .A2(n5040), .ZN(n8664) );
  OAI222_X1 U4923 ( .A1(n8883), .A2(n8107), .B1(P2_U3152), .B2(n5754), .C1(
        n7734), .C2(n8888), .ZN(P2_U3329) );
  AOI21_X4 U4924 ( .B1(n9227), .B2(n5522), .A(n7891), .ZN(n9202) );
  XNOR2_X2 U4925 ( .A(n8789), .B(n8608), .ZN(n8259) );
  NAND2_X2 U4926 ( .A1(n5542), .A2(n5541), .ZN(n9419) );
  OAI22_X2 U4927 ( .A1(n7476), .A2(n8419), .B1(n7484), .B2(n8458), .ZN(n7555)
         );
  XNOR2_X2 U4928 ( .A(n8468), .B(n8290), .ZN(n10187) );
  OAI22_X2 U4929 ( .A1(n9276), .A2(n9283), .B1(n8915), .B2(n9281), .ZN(n9272)
         );
  AOI21_X2 U4930 ( .B1(n9290), .B2(n5713), .A(n5712), .ZN(n9276) );
  AND3_X1 U4931 ( .A1(n7695), .A2(n8979), .A3(n7701), .ZN(n8904) );
  NAND2_X2 U4932 ( .A1(n8276), .A2(n8277), .ZN(n8401) );
  CLKBUF_X2 U4933 ( .A(n7679), .Z(n4391) );
  INV_X1 U4934 ( .A(n10182), .ZN(n10262) );
  CLKBUF_X3 U4935 ( .A(n7679), .Z(n4388) );
  INV_X1 U4936 ( .A(n6562), .ZN(n10087) );
  INV_X1 U4937 ( .A(n9998), .ZN(n10093) );
  NAND2_X1 U4938 ( .A1(n6088), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5776) );
  CLKBUF_X2 U4940 ( .A(n5791), .Z(n6077) );
  INV_X1 U4941 ( .A(n10023), .ZN(n10028) );
  CLKBUF_X2 U4943 ( .A(n5452), .Z(n5582) );
  INV_X1 U4944 ( .A(n5754), .ZN(n5752) );
  INV_X2 U4945 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4946 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5761) );
  AOI21_X1 U4947 ( .B1(n4384), .B2(n10302), .A(n4733), .ZN(n4732) );
  NOR2_X1 U4948 ( .A1(n8961), .A2(n8960), .ZN(n8959) );
  AOI21_X1 U4949 ( .B1(n4751), .B2(n4750), .A(n8441), .ZN(n8452) );
  OAI21_X1 U4950 ( .B1(n8570), .B2(n8573), .A(n4990), .ZN(n8557) );
  NAND2_X1 U4951 ( .A1(n7694), .A2(n7693), .ZN(n8979) );
  AOI211_X1 U4952 ( .C1(n9987), .C2(n9143), .A(n9142), .B(n9141), .ZN(n9404)
         );
  NAND2_X1 U4953 ( .A1(n4631), .A2(n4630), .ZN(n8914) );
  NAND2_X1 U4954 ( .A1(n5002), .A2(n5003), .ZN(n8693) );
  NAND2_X1 U4955 ( .A1(n4620), .A2(n4415), .ZN(n9012) );
  NAND2_X1 U4956 ( .A1(n7633), .A2(n7632), .ZN(n8891) );
  OR2_X1 U4957 ( .A1(n7537), .A2(n7538), .ZN(n7565) );
  OAI211_X1 U4958 ( .C1(n4944), .C2(n4645), .A(n7623), .B(n4642), .ZN(n7630)
         );
  OAI21_X1 U4959 ( .B1(n5577), .B2(n5576), .A(n5591), .ZN(n7571) );
  OR2_X1 U4960 ( .A1(n8689), .A2(n8218), .ZN(n5040) );
  NAND2_X1 U4961 ( .A1(n5483), .A2(n5482), .ZN(n9439) );
  NAND2_X1 U4962 ( .A1(n6025), .A2(n6024), .ZN(n8814) );
  NAND2_X1 U4963 ( .A1(n5360), .A2(n5359), .ZN(n9457) );
  NAND2_X1 U4964 ( .A1(n5339), .A2(n5338), .ZN(n9464) );
  OAI21_X1 U4965 ( .B1(n5382), .B2(n5381), .A(n5380), .ZN(n5404) );
  NAND2_X1 U4966 ( .A1(n5319), .A2(n5318), .ZN(n9468) );
  NAND2_X1 U4967 ( .A1(n5301), .A2(n5300), .ZN(n7326) );
  NAND2_X1 U4968 ( .A1(n5906), .A2(n5905), .ZN(n7264) );
  OR3_X2 U4969 ( .A1(n6220), .A2(n8851), .A3(n6400), .ZN(n8233) );
  NAND2_X1 U4970 ( .A1(n5292), .A2(n5291), .ZN(n5312) );
  INV_X2 U4971 ( .A(n10134), .ZN(n4387) );
  AND2_X2 U4972 ( .A1(n6734), .A2(n6383), .ZN(n7770) );
  NAND2_X2 U4973 ( .A1(n4810), .A2(n8445), .ZN(n8138) );
  OAI211_X1 U4974 ( .C1(n6190), .C2(n6320), .A(n5212), .B(n5211), .ZN(n7102)
         );
  AND2_X1 U4975 ( .A1(n7934), .A2(n6861), .ZN(n6732) );
  AND2_X2 U4976 ( .A1(n9873), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U4006) );
  NAND4_X1 U4977 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n10206)
         );
  XNOR2_X1 U4978 ( .A(n5106), .B(n5105), .ZN(n7934) );
  OAI211_X1 U4979 ( .C1(n6190), .C2(n6264), .A(n5176), .B(n5175), .ZN(n6562)
         );
  NAND4_X1 U4980 ( .A1(n5167), .A2(n5166), .A3(n5165), .A4(n5164), .ZN(n10009)
         );
  INV_X4 U4981 ( .A(n5177), .ZN(n6484) );
  NAND2_X1 U4982 ( .A1(n5104), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5106) );
  OR2_X1 U4983 ( .A1(n7806), .A2(n6260), .ZN(n5160) );
  NAND2_X2 U4984 ( .A1(n7596), .A2(n5119), .ZN(n5485) );
  OAI21_X1 U4985 ( .B1(n4562), .B2(n4514), .A(n4512), .ZN(n5206) );
  INV_X1 U4986 ( .A(n5120), .ZN(n5119) );
  NAND2_X1 U4987 ( .A1(n5143), .A2(n6259), .ZN(n5219) );
  AOI21_X1 U4988 ( .B1(n5189), .B2(n4513), .A(n4460), .ZN(n4512) );
  OAI21_X1 U4989 ( .B1(n5241), .B2(n4883), .A(n5250), .ZN(n4882) );
  NAND4_X1 U4990 ( .A1(n4590), .A2(n4589), .A3(n4588), .A4(n4587), .ZN(n5753)
         );
  NAND2_X1 U4991 ( .A1(n4729), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4728) );
  NAND2_X1 U4992 ( .A1(n5736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5737) );
  CLKBUF_X1 U4993 ( .A(n5640), .Z(n9874) );
  XNOR2_X1 U4994 ( .A(n5128), .B(n5127), .ZN(n5640) );
  NAND2_X1 U4995 ( .A1(n5116), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5118) );
  NAND2_X1 U4996 ( .A1(n9772), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5115) );
  NAND2_X2 U4997 ( .A1(n7800), .A2(P1_U3084), .ZN(n9782) );
  OR2_X1 U4998 ( .A1(n5126), .A2(n5280), .ZN(n5128) );
  INV_X2 U4999 ( .A(n9777), .ZN(n4389) );
  NOR2_X1 U5000 ( .A1(n4417), .A2(n4958), .ZN(n4957) );
  AND2_X1 U5002 ( .A1(n5087), .A2(n5079), .ZN(n5037) );
  BUF_X4 U5003 ( .A(n5134), .Z(n6259) );
  AND2_X1 U5004 ( .A1(n5245), .A2(n5065), .ZN(n5257) );
  AND2_X1 U5005 ( .A1(n4821), .A2(n4818), .ZN(n5044) );
  NOR2_X1 U5006 ( .A1(n5220), .A2(n5078), .ZN(n5336) );
  AND2_X1 U5007 ( .A1(n5828), .A2(n4424), .ZN(n4814) );
  AND4_X1 U5008 ( .A1(n4472), .A2(n4942), .A3(n5063), .A4(n5062), .ZN(n5245)
         );
  NAND2_X2 U5009 ( .A1(n4508), .A2(n4506), .ZN(n5134) );
  INV_X1 U5010 ( .A(n4959), .ZN(n4958) );
  NAND3_X1 U5011 ( .A1(n4511), .A2(n4510), .A3(n4509), .ZN(n4508) );
  NAND3_X1 U5012 ( .A1(n4507), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4506) );
  AND2_X1 U5013 ( .A1(n5066), .A2(n5075), .ZN(n4959) );
  AND2_X1 U5014 ( .A1(n4816), .A2(n4815), .ZN(n4821) );
  AND3_X1 U5015 ( .A1(n5726), .A2(n4820), .A3(n4819), .ZN(n4818) );
  NOR2_X2 U5016 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5062) );
  INV_X1 U5017 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6121) );
  NOR2_X1 U5018 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n4815) );
  NOR2_X2 U5019 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5063) );
  INV_X1 U5020 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6009) );
  NOR2_X1 U5021 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4816) );
  INV_X1 U5022 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5079) );
  NOR2_X1 U5023 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5724) );
  NOR2_X2 U5024 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5798) );
  NOR2_X1 U5025 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n5084) );
  INV_X1 U5026 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5725) );
  INV_X2 U5027 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  INV_X1 U5028 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5075) );
  INV_X1 U5029 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5102) );
  INV_X1 U5030 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4507) );
  NAND4_X4 U5031 ( .A1(n5776), .A2(n5775), .A3(n5774), .A4(n5773), .ZN(n5787)
         );
  OAI21_X2 U5032 ( .B1(n6957), .B2(n5848), .A(n5847), .ZN(n6968) );
  NAND2_X1 U5033 ( .A1(n5833), .A2(n5832), .ZN(n6957) );
  OR2_X2 U5034 ( .A1(n7489), .A2(n8328), .ZN(n7491) );
  OAI22_X2 U5035 ( .A1(n7311), .A2(n7312), .B1(n10295), .B2(n8460), .ZN(n7489)
         );
  AOI21_X2 U5036 ( .B1(n8693), .B2(n6006), .A(n6005), .ZN(n8678) );
  OAI22_X2 U5037 ( .A1(n9167), .A2(n8048), .B1(n9029), .B2(n9412), .ZN(n9154)
         );
  INV_X1 U5038 ( .A(n4794), .ZN(n9167) );
  NAND2_X1 U5039 ( .A1(n5753), .A2(n5754), .ZN(n5823) );
  AND2_X1 U5040 ( .A1(n6384), .A2(n6733), .ZN(n7679) );
  AOI21_X1 U5041 ( .B1(n4790), .B2(n4788), .A(n4441), .ZN(n4787) );
  INV_X1 U5042 ( .A(n4413), .ZN(n4788) );
  AOI21_X1 U5043 ( .B1(n4462), .B2(n8371), .A(n4559), .ZN(n4558) );
  INV_X1 U5044 ( .A(n8375), .ZN(n4559) );
  INV_X1 U5045 ( .A(n8369), .ZN(n4561) );
  NAND2_X1 U5046 ( .A1(n7938), .A2(n4858), .ZN(n8024) );
  NAND2_X1 U5047 ( .A1(n6401), .A2(n6259), .ZN(n5817) );
  AOI21_X1 U5048 ( .B1(n4888), .B2(n4890), .A(n4885), .ZN(n4884) );
  INV_X1 U5049 ( .A(n5590), .ZN(n4885) );
  INV_X1 U5050 ( .A(n5552), .ZN(n4895) );
  INV_X2 U5051 ( .A(n5845), .ZN(n8249) );
  NAND2_X2 U5052 ( .A1(n6401), .A2(n7800), .ZN(n5845) );
  INV_X1 U5053 ( .A(n4787), .ZN(n4786) );
  AOI21_X1 U5054 ( .B1(n4787), .B2(n4789), .A(n4785), .ZN(n4784) );
  AND2_X1 U5055 ( .A1(n5113), .A2(n5112), .ZN(n9989) );
  AOI21_X1 U5056 ( .B1(n4558), .B2(n4560), .A(n8374), .ZN(n4557) );
  INV_X1 U5057 ( .A(n8371), .ZN(n4560) );
  NAND2_X1 U5058 ( .A1(n5254), .A2(n5253), .ZN(n5272) );
  NAND3_X1 U5059 ( .A1(n8433), .A2(n10243), .A3(n8436), .ZN(n4810) );
  INV_X1 U5060 ( .A(n4983), .ZN(n4981) );
  NAND2_X1 U5061 ( .A1(n8583), .A2(n8259), .ZN(n4975) );
  NOR2_X1 U5062 ( .A1(n8637), .A2(n5000), .ZN(n4999) );
  NOR2_X1 U5063 ( .A1(n4394), .A2(n6038), .ZN(n5000) );
  NAND2_X1 U5064 ( .A1(n4599), .A2(n8656), .ZN(n4598) );
  INV_X1 U5065 ( .A(n4601), .ZN(n4599) );
  AND2_X1 U5066 ( .A1(n8716), .A2(n8340), .ZN(n8744) );
  OR2_X1 U5067 ( .A1(n7367), .A2(n5931), .ZN(n8317) );
  OR2_X1 U5068 ( .A1(n10275), .A2(n8466), .ZN(n8298) );
  NAND2_X1 U5069 ( .A1(n8836), .A2(n8720), .ZN(n5004) );
  OR2_X1 U5070 ( .A1(n6160), .A2(n4591), .ZN(n4590) );
  INV_X1 U5071 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5748) );
  AND2_X1 U5072 ( .A1(n5761), .A2(n5982), .ZN(n4812) );
  OAI21_X1 U5073 ( .B1(n7926), .B2(n4927), .A(n4926), .ZN(n7932) );
  NAND2_X1 U5074 ( .A1(n7931), .A2(n7930), .ZN(n4926) );
  NAND2_X1 U5075 ( .A1(n5195), .A2(n5011), .ZN(n7818) );
  NAND2_X1 U5076 ( .A1(n5135), .A2(n6747), .ZN(n5680) );
  NAND2_X1 U5077 ( .A1(n5025), .A2(n5023), .ZN(n9172) );
  NAND2_X1 U5078 ( .A1(n5024), .A2(n8048), .ZN(n5023) );
  INV_X1 U5079 ( .A(n5027), .ZN(n5024) );
  AOI21_X1 U5080 ( .B1(n4876), .B2(n4874), .A(n4491), .ZN(n4873) );
  INV_X1 U5081 ( .A(n5607), .ZN(n4874) );
  AOI21_X1 U5082 ( .B1(n5553), .B2(n4894), .A(n4892), .ZN(n4891) );
  INV_X1 U5083 ( .A(n5570), .ZN(n4892) );
  AND2_X1 U5084 ( .A1(n5590), .A2(n5575), .ZN(n5576) );
  NAND2_X1 U5085 ( .A1(n5540), .A2(n5539), .ZN(n5554) );
  NAND2_X1 U5086 ( .A1(n4900), .A2(n4898), .ZN(n5540) );
  AOI21_X1 U5087 ( .B1(n4901), .B2(n4475), .A(n4899), .ZN(n4898) );
  OAI21_X1 U5088 ( .B1(n5477), .B2(n5476), .A(n5475), .ZN(n5495) );
  AND2_X1 U5089 ( .A1(n5496), .A2(n5481), .ZN(n5494) );
  OAI21_X1 U5090 ( .B1(n5404), .B2(n5403), .A(n5402), .ZN(n5421) );
  XNOR2_X1 U5091 ( .A(n5378), .B(SI_14_), .ZN(n5377) );
  NAND2_X1 U5092 ( .A1(n4909), .A2(n4907), .ZN(n5382) );
  AOI21_X1 U5093 ( .B1(n4911), .B2(n4914), .A(n4908), .ZN(n4907) );
  NAND2_X1 U5094 ( .A1(n5331), .A2(n4911), .ZN(n4909) );
  INV_X1 U5095 ( .A(n5368), .ZN(n4908) );
  NOR2_X1 U5096 ( .A1(n5350), .A2(n4918), .ZN(n4917) );
  INV_X1 U5097 ( .A(n5330), .ZN(n4918) );
  NAND2_X1 U5098 ( .A1(n4581), .A2(n5313), .ZN(n5331) );
  NAND2_X1 U5099 ( .A1(n5312), .A2(n5039), .ZN(n4581) );
  NAND2_X1 U5100 ( .A1(n4879), .A2(n4878), .ZN(n5274) );
  AOI21_X1 U5101 ( .B1(n4881), .B2(n4883), .A(n4453), .ZN(n4878) );
  INV_X1 U5102 ( .A(n4882), .ZN(n4881) );
  NAND2_X1 U5103 ( .A1(n8180), .A2(n4571), .ZN(n4569) );
  AOI21_X1 U5104 ( .B1(n4691), .B2(n8166), .A(n4459), .ZN(n4689) );
  INV_X1 U5105 ( .A(n8167), .ZN(n8119) );
  INV_X1 U5106 ( .A(n6218), .ZN(n4842) );
  NAND2_X1 U5107 ( .A1(n4811), .A2(n8680), .ZN(n8433) );
  NAND2_X2 U5108 ( .A1(n8881), .A2(n5754), .ZN(n6286) );
  NAND2_X1 U5109 ( .A1(n4975), .A2(n4974), .ZN(n4984) );
  AND2_X1 U5110 ( .A1(n4988), .A2(n4393), .ZN(n4974) );
  NAND2_X1 U5111 ( .A1(n8648), .A2(n4999), .ZN(n4997) );
  NAND2_X1 U5112 ( .A1(n4596), .A2(n4595), .ZN(n8655) );
  AOI21_X1 U5113 ( .B1(n4601), .B2(n4603), .A(n4600), .ZN(n4595) );
  NAND2_X1 U5114 ( .A1(n4602), .A2(n4601), .ZN(n4596) );
  NOR2_X1 U5115 ( .A1(n8721), .A2(n8826), .ZN(n6005) );
  NAND2_X1 U5116 ( .A1(n7248), .A2(n5875), .ZN(n4970) );
  NAND2_X1 U5117 ( .A1(n5859), .A2(n4971), .ZN(n4969) );
  NOR2_X1 U5118 ( .A1(n8297), .A2(n4972), .ZN(n4971) );
  NAND2_X1 U5119 ( .A1(n6097), .A2(n6096), .ZN(n8771) );
  AND2_X1 U5120 ( .A1(n6695), .A2(n4936), .ZN(n4935) );
  NAND2_X1 U5122 ( .A1(n5121), .A2(n5120), .ZN(n5179) );
  AND2_X1 U5123 ( .A1(n7596), .A2(n5120), .ZN(n5178) );
  NOR2_X1 U5124 ( .A1(n4717), .A2(n9401), .ZN(n4713) );
  OAI21_X1 U5125 ( .B1(n4778), .B2(n4777), .A(n4452), .ZN(n4776) );
  OR2_X1 U5126 ( .A1(n9826), .A2(n9016), .ZN(n5038) );
  INV_X1 U5127 ( .A(n5710), .ZN(n4791) );
  NAND2_X1 U5128 ( .A1(n4793), .A2(n4413), .ZN(n4792) );
  INV_X1 U5129 ( .A(n9344), .ZN(n4793) );
  INV_X1 U5130 ( .A(n7806), .ZN(n5466) );
  INV_X1 U5131 ( .A(n6190), .ZN(n5465) );
  AND2_X1 U5132 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  INV_X1 U5133 ( .A(n10116), .ZN(n9822) );
  AND2_X1 U5134 ( .A1(n5539), .A2(n5529), .ZN(n5537) );
  NAND2_X1 U5135 ( .A1(n5495), .A2(n5494), .ZN(n5497) );
  AOI21_X1 U5136 ( .B1(n7766), .B2(n8711), .A(n7765), .ZN(n4617) );
  NAND2_X1 U5137 ( .A1(n4799), .A2(n4798), .ZN(n5718) );
  AOI21_X1 U5138 ( .B1(n4396), .B2(n4801), .A(n4451), .ZN(n4798) );
  OAI21_X1 U5139 ( .B1(n8289), .B2(n8269), .A(n4445), .ZN(n8270) );
  INV_X1 U5140 ( .A(n8294), .ZN(n4520) );
  NAND2_X1 U5141 ( .A1(n4518), .A2(n8380), .ZN(n4517) );
  INV_X1 U5142 ( .A(n8298), .ZN(n4518) );
  NOR2_X1 U5143 ( .A1(n4532), .A2(n4759), .ZN(n4531) );
  INV_X1 U5144 ( .A(n8331), .ZN(n4532) );
  NAND2_X1 U5145 ( .A1(n8417), .A2(n8334), .ZN(n4530) );
  NOR2_X1 U5146 ( .A1(n4530), .A2(n8416), .ZN(n4527) );
  AND2_X1 U5147 ( .A1(n8744), .A2(n8339), .ZN(n4533) );
  INV_X1 U5148 ( .A(n7903), .ZN(n4505) );
  NAND2_X1 U5149 ( .A1(n4458), .A2(n4549), .ZN(n4548) );
  NAND2_X1 U5150 ( .A1(n8357), .A2(n4550), .ZN(n4549) );
  INV_X1 U5151 ( .A(n8355), .ZN(n4550) );
  NOR2_X1 U5152 ( .A1(n9027), .A2(n7933), .ZN(n4930) );
  NAND2_X1 U5153 ( .A1(n4503), .A2(n7918), .ZN(n7919) );
  INV_X1 U5154 ( .A(n4873), .ZN(n4871) );
  AOI21_X1 U5155 ( .B1(n4554), .B2(n4556), .A(n4463), .ZN(n4553) );
  INV_X1 U5156 ( .A(n4557), .ZN(n4556) );
  NAND2_X1 U5157 ( .A1(n9412), .A2(n9186), .ZN(n7904) );
  OR2_X1 U5158 ( .A1(n9412), .A2(n9186), .ZN(n7939) );
  INV_X1 U5159 ( .A(n8003), .ZN(n5021) );
  OAI21_X1 U5160 ( .B1(n9261), .B2(n5021), .A(n7960), .ZN(n5020) );
  INV_X1 U5161 ( .A(n4864), .ZN(n4863) );
  OAI21_X1 U5162 ( .B1(n4866), .B2(n4865), .A(n5458), .ZN(n4864) );
  INV_X1 U5163 ( .A(n5440), .ZN(n4865) );
  NAND2_X1 U5164 ( .A1(n5333), .A2(n5332), .ZN(n5349) );
  NAND2_X1 U5165 ( .A1(n5277), .A2(n5276), .ZN(n5291) );
  INV_X1 U5166 ( .A(n8155), .ZN(n4578) );
  INV_X1 U5167 ( .A(n7446), .ZN(n4686) );
  OR2_X1 U5168 ( .A1(n8762), .A2(n8253), .ZN(n8392) );
  INV_X1 U5169 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4960) );
  INV_X1 U5170 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5726) );
  NOR2_X1 U5171 ( .A1(n8426), .A2(n4985), .ZN(n4983) );
  NAND2_X1 U5172 ( .A1(n8561), .A2(n6095), .ZN(n4989) );
  AND2_X1 U5173 ( .A1(n4989), .A2(n4990), .ZN(n4988) );
  OR2_X1 U5174 ( .A1(n8777), .A2(n6095), .ZN(n8377) );
  OR2_X1 U5175 ( .A1(n8783), .A2(n8151), .ZN(n8375) );
  NOR2_X1 U5176 ( .A1(n4770), .A2(n8372), .ZN(n4769) );
  INV_X1 U5177 ( .A(n4999), .ZN(n4994) );
  OR2_X1 U5178 ( .A1(n8792), .A2(n8159), .ZN(n8365) );
  INV_X1 U5179 ( .A(n8656), .ZN(n4600) );
  INV_X1 U5180 ( .A(n8681), .ZN(n4772) );
  OR2_X1 U5181 ( .A1(n8831), .A2(n7581), .ZN(n8261) );
  AND2_X1 U5182 ( .A1(n4604), .A2(n4758), .ZN(n8746) );
  NAND2_X1 U5183 ( .A1(n4605), .A2(n4761), .ZN(n4604) );
  OR2_X1 U5184 ( .A1(n7484), .A2(n7450), .ZN(n8333) );
  NAND2_X1 U5185 ( .A1(n4737), .A2(n4736), .ZN(n7188) );
  INV_X1 U5186 ( .A(n8300), .ZN(n4748) );
  AND2_X1 U5187 ( .A1(n8280), .A2(n8276), .ZN(n4757) );
  OR2_X2 U5188 ( .A1(n5787), .A2(n10246), .ZN(n8277) );
  NAND2_X1 U5189 ( .A1(n8610), .A2(n8365), .ZN(n8588) );
  OR2_X1 U5190 ( .A1(n8738), .A2(n8744), .ZN(n5005) );
  INV_X1 U5191 ( .A(n4943), .ZN(n4643) );
  NOR2_X1 U5192 ( .A1(n4947), .A2(n4946), .ZN(n4945) );
  INV_X1 U5193 ( .A(n4949), .ZN(n4946) );
  INV_X1 U5194 ( .A(n4484), .ZN(n4947) );
  AND2_X1 U5195 ( .A1(n7403), .A2(n7402), .ZN(n4943) );
  INV_X1 U5196 ( .A(n7406), .ZN(n7403) );
  AOI21_X1 U5197 ( .B1(n4639), .B2(n4641), .A(n4446), .ZN(n4638) );
  OR2_X1 U5198 ( .A1(n7387), .A2(n7386), .ZN(n7396) );
  XNOR2_X1 U5199 ( .A(n4621), .B(n7716), .ZN(n6753) );
  NAND2_X1 U5200 ( .A1(n6685), .A2(n4622), .ZN(n4621) );
  NAND2_X1 U5201 ( .A1(n9986), .A2(n4386), .ZN(n4622) );
  INV_X1 U5202 ( .A(n7735), .ZN(n4629) );
  OR2_X1 U5203 ( .A1(n7710), .A2(n7709), .ZN(n4956) );
  NOR2_X1 U5204 ( .A1(n9401), .A2(n9164), .ZN(n7810) );
  OR2_X1 U5205 ( .A1(n9396), .A2(n7727), .ZN(n8019) );
  AND2_X1 U5206 ( .A1(n9401), .A2(n9164), .ZN(n8011) );
  NOR2_X1 U5207 ( .A1(n9241), .A2(n9427), .ZN(n4711) );
  OR2_X1 U5208 ( .A1(n9427), .A2(n8924), .ZN(n8028) );
  NOR2_X1 U5209 ( .A1(n9318), .A2(n9340), .ZN(n4724) );
  OR2_X1 U5210 ( .A1(n9318), .A2(n9016), .ZN(n7859) );
  NAND2_X1 U5211 ( .A1(n9366), .A2(n9365), .ZN(n5036) );
  OR2_X1 U5212 ( .A1(n7326), .A2(n5311), .ZN(n7973) );
  NAND2_X1 U5213 ( .A1(n6800), .A2(n5031), .ZN(n7014) );
  NOR2_X1 U5214 ( .A1(n5033), .A2(n5032), .ZN(n5031) );
  INV_X1 U5215 ( .A(n7996), .ZN(n5033) );
  AND2_X1 U5216 ( .A1(n7013), .A2(n7996), .ZN(n8036) );
  NAND2_X1 U5217 ( .A1(n10007), .A2(n4434), .ZN(n9982) );
  NAND2_X1 U5218 ( .A1(n5680), .A2(n6740), .ZN(n8060) );
  NAND2_X1 U5219 ( .A1(n10074), .A2(n6492), .ZN(n4809) );
  INV_X1 U5220 ( .A(n9143), .ZN(n9176) );
  AOI21_X1 U5221 ( .B1(n5028), .B2(n9203), .A(n5548), .ZN(n5027) );
  XNOR2_X1 U5222 ( .A(n7797), .B(n7796), .ZN(n7794) );
  INV_X1 U5223 ( .A(n5623), .ZN(n4877) );
  NOR2_X1 U5224 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4808) );
  AOI21_X1 U5225 ( .B1(n4891), .B2(n4893), .A(n4889), .ZN(n4888) );
  INV_X1 U5226 ( .A(n5576), .ZN(n4889) );
  INV_X1 U5227 ( .A(n4891), .ZN(n4890) );
  INV_X1 U5228 ( .A(n5377), .ZN(n5381) );
  NAND2_X1 U5229 ( .A1(n5402), .A2(n5386), .ZN(n5403) );
  NAND2_X1 U5230 ( .A1(n5272), .A2(n5256), .ZN(n5273) );
  INV_X1 U5231 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n4941) );
  XNOR2_X1 U5232 ( .A(n5252), .B(SI_7_), .ZN(n5249) );
  INV_X1 U5233 ( .A(n5240), .ZN(n5241) );
  NAND2_X1 U5234 ( .A1(n5218), .A2(n5217), .ZN(n5242) );
  AND2_X1 U5235 ( .A1(n8174), .A2(n8143), .ZN(n8148) );
  INV_X1 U5236 ( .A(n8120), .ZN(n4692) );
  OAI211_X1 U5237 ( .C1(n6401), .C2(n6465), .A(n5846), .B(n4515), .ZN(n6192)
         );
  OR2_X1 U5238 ( .A1(n6266), .A2(n5845), .ZN(n4515) );
  NAND2_X1 U5239 ( .A1(n5745), .A2(n5744), .ZN(n6034) );
  INV_X1 U5240 ( .A(n6027), .ZN(n5745) );
  OR2_X1 U5241 ( .A1(n6034), .A2(n8189), .ZN(n6041) );
  NOR2_X1 U5242 ( .A1(n10298), .A2(n8680), .ZN(n6725) );
  NAND2_X1 U5243 ( .A1(n4584), .A2(n7149), .ZN(n4583) );
  INV_X1 U5244 ( .A(n7261), .ZN(n4584) );
  AND2_X1 U5245 ( .A1(n7031), .A2(n7074), .ZN(n7030) );
  OR2_X1 U5246 ( .A1(n7037), .A2(n7036), .ZN(n7031) );
  OAI21_X1 U5247 ( .B1(n6819), .B2(n4824), .A(n4822), .ZN(n7075) );
  INV_X1 U5248 ( .A(n4823), .ZN(n4822) );
  OAI21_X1 U5249 ( .B1(n4825), .B2(n4824), .A(n6837), .ZN(n4823) );
  INV_X1 U5250 ( .A(n6836), .ZN(n4824) );
  XNOR2_X1 U5251 ( .A(n7043), .B(n4421), .ZN(n7037) );
  NAND2_X1 U5252 ( .A1(n10139), .A2(n10140), .ZN(n10138) );
  AND2_X1 U5253 ( .A1(n4836), .A2(n4835), .ZN(n4834) );
  INV_X1 U5254 ( .A(n8236), .ZN(n4835) );
  NAND3_X1 U5255 ( .A1(n4696), .A2(n4694), .A3(n4693), .ZN(n4837) );
  OR2_X1 U5256 ( .A1(n8156), .A2(n4695), .ZN(n4694) );
  INV_X1 U5257 ( .A(n4697), .ZN(n4696) );
  NAND2_X1 U5258 ( .A1(n4698), .A2(n4397), .ZN(n4693) );
  NOR2_X1 U5259 ( .A1(n7534), .A2(n4686), .ZN(n4684) );
  NAND2_X1 U5260 ( .A1(n4684), .A2(n7303), .ZN(n4680) );
  NAND2_X1 U5261 ( .A1(n7534), .A2(n4686), .ZN(n4685) );
  INV_X1 U5262 ( .A(n7303), .ZN(n4683) );
  AND2_X1 U5263 ( .A1(n8392), .A2(n8390), .ZN(n8399) );
  AND2_X1 U5264 ( .A1(n8762), .A2(n8253), .ZN(n8395) );
  OR2_X1 U5265 ( .A1(n8553), .A2(n6146), .ZN(n8391) );
  INV_X1 U5266 ( .A(n6290), .ZN(n5921) );
  OAI21_X1 U5267 ( .B1(n8533), .B2(n8732), .A(n8522), .ZN(n7743) );
  NAND2_X1 U5268 ( .A1(n6109), .A2(n6108), .ZN(n7759) );
  NAND2_X1 U5269 ( .A1(n8558), .A2(n8181), .ZN(n7599) );
  NAND2_X1 U5270 ( .A1(n8783), .A2(n8151), .ZN(n8562) );
  NAND2_X1 U5271 ( .A1(n4735), .A2(n4991), .ZN(n8576) );
  NAND2_X1 U5272 ( .A1(n8588), .A2(n8587), .ZN(n4771) );
  NAND2_X1 U5273 ( .A1(n4771), .A2(n4769), .ZN(n8571) );
  OR2_X1 U5274 ( .A1(n6052), .A2(n6051), .ZN(n6065) );
  AOI21_X1 U5275 ( .B1(n4999), .B2(n4394), .A(n4457), .ZN(n4998) );
  OR2_X1 U5276 ( .A1(n8804), .A2(n8190), .ZN(n8615) );
  NAND3_X1 U5277 ( .A1(n8636), .A2(n8625), .A3(n8615), .ZN(n8616) );
  AND2_X1 U5278 ( .A1(n8615), .A2(n8349), .ZN(n8637) );
  NAND2_X1 U5279 ( .A1(n8356), .A2(n4772), .ZN(n4603) );
  NAND2_X1 U5280 ( .A1(n4406), .A2(n8356), .ZN(n4601) );
  AND2_X1 U5281 ( .A1(n8814), .A2(n8658), .ZN(n6031) );
  AND2_X1 U5282 ( .A1(n8360), .A2(n8638), .ZN(n8656) );
  AOI21_X1 U5283 ( .B1(n4395), .B2(n8744), .A(n4455), .ZN(n5003) );
  NAND2_X1 U5284 ( .A1(n8261), .A2(n8262), .ZN(n8717) );
  OR2_X1 U5285 ( .A1(n8836), .A2(n7566), .ZN(n8716) );
  NAND2_X1 U5286 ( .A1(n7556), .A2(n8335), .ZN(n8752) );
  INV_X1 U5287 ( .A(n8333), .ZN(n4762) );
  INV_X1 U5288 ( .A(n7477), .ZN(n4760) );
  INV_X1 U5289 ( .A(n4605), .ZN(n7478) );
  NAND2_X1 U5290 ( .A1(n7478), .A2(n8419), .ZN(n7477) );
  INV_X1 U5291 ( .A(n4610), .ZN(n4609) );
  AOI21_X1 U5292 ( .B1(n4964), .B2(n4966), .A(n4442), .ZN(n4963) );
  NAND2_X1 U5293 ( .A1(n7189), .A2(n7225), .ZN(n7317) );
  AND2_X1 U5294 ( .A1(n8312), .A2(n8304), .ZN(n8411) );
  NAND2_X1 U5295 ( .A1(n5915), .A2(n5914), .ZN(n7178) );
  NAND2_X1 U5296 ( .A1(n4612), .A2(n8411), .ZN(n7184) );
  INV_X1 U5297 ( .A(n7181), .ZN(n4612) );
  NOR2_X1 U5298 ( .A1(n8307), .A2(n4968), .ZN(n4967) );
  INV_X1 U5299 ( .A(n4970), .ZN(n4968) );
  AND2_X1 U5300 ( .A1(n6133), .A2(n8298), .ZN(n6134) );
  NAND2_X1 U5301 ( .A1(n6134), .A2(n8297), .ZN(n6981) );
  OR2_X1 U5302 ( .A1(n5845), .A2(n6263), .ZN(n5819) );
  NAND2_X1 U5303 ( .A1(n6159), .A2(P2_IR_REG_30__SCAN_IN), .ZN(n4587) );
  OR2_X1 U5304 ( .A1(n4593), .A2(n4591), .ZN(n4588) );
  NAND2_X1 U5305 ( .A1(n6160), .A2(n5008), .ZN(n4729) );
  NOR2_X1 U5306 ( .A1(n4404), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n4857) );
  NAND2_X1 U5307 ( .A1(n5760), .A2(n5761), .ZN(n4813) );
  XNOR2_X1 U5308 ( .A(n5777), .B(P2_IR_REG_1__SCAN_IN), .ZN(n9791) );
  NAND2_X1 U5309 ( .A1(n7695), .A2(n8979), .ZN(n4649) );
  NOR2_X1 U5310 ( .A1(n7664), .A2(n9004), .ZN(n4635) );
  INV_X1 U5311 ( .A(n7657), .ZN(n4633) );
  INV_X1 U5312 ( .A(n6702), .ZN(n6700) );
  INV_X1 U5313 ( .A(n8901), .ZN(n4647) );
  NAND2_X1 U5314 ( .A1(n8914), .A2(n4950), .ZN(n4948) );
  OR2_X1 U5315 ( .A1(n8911), .A2(n8912), .ZN(n4950) );
  NOR2_X1 U5316 ( .A1(n7735), .A2(n4954), .ZN(n4953) );
  INV_X1 U5317 ( .A(n4956), .ZN(n4954) );
  OR2_X1 U5318 ( .A1(n7937), .A2(n4925), .ZN(n4924) );
  NOR2_X1 U5319 ( .A1(n8058), .A2(n8093), .ZN(n4922) );
  NAND2_X1 U5320 ( .A1(n5201), .A2(n5202), .ZN(n4624) );
  OR2_X1 U5321 ( .A1(n5452), .A2(n6557), .ZN(n5145) );
  OR2_X1 U5322 ( .A1(n9917), .A2(n4477), .ZN(n4672) );
  NAND2_X1 U5323 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  INV_X1 U5324 ( .A(n6369), .ZN(n4671) );
  NAND2_X1 U5325 ( .A1(n6361), .A2(n6362), .ZN(n6599) );
  NAND2_X1 U5326 ( .A1(n6636), .A2(n6637), .ZN(n6999) );
  OR2_X1 U5327 ( .A1(n9044), .A2(n9335), .ZN(n4676) );
  NOR2_X1 U5328 ( .A1(n9821), .A2(n4715), .ZN(n4714) );
  NAND2_X1 U5329 ( .A1(n4716), .A2(n9150), .ZN(n4715) );
  INV_X1 U5330 ( .A(n4717), .ZN(n4716) );
  OR3_X1 U5331 ( .A1(n5614), .A2(n5613), .A3(n5612), .ZN(n5655) );
  NAND2_X1 U5332 ( .A1(n9140), .A2(n4802), .ZN(n4801) );
  INV_X1 U5333 ( .A(n4804), .ZN(n4802) );
  NAND2_X1 U5334 ( .A1(n9150), .A2(n9164), .ZN(n4803) );
  NOR2_X1 U5335 ( .A1(n9138), .A2(n7810), .ZN(n9122) );
  NAND2_X1 U5336 ( .A1(n8019), .A2(n8014), .ZN(n9128) );
  INV_X1 U5337 ( .A(n9136), .ZN(n9140) );
  INV_X1 U5338 ( .A(n9028), .ZN(n9164) );
  OR2_X1 U5339 ( .A1(n9188), .A2(n9412), .ZN(n9168) );
  NOR2_X1 U5340 ( .A1(n9184), .A2(n7815), .ZN(n5028) );
  OR2_X1 U5341 ( .A1(n9202), .A2(n9203), .ZN(n5029) );
  INV_X1 U5342 ( .A(n8046), .ZN(n9184) );
  NAND2_X1 U5343 ( .A1(n5059), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5518) );
  INV_X1 U5344 ( .A(n5500), .ZN(n5059) );
  INV_X1 U5345 ( .A(n4779), .ZN(n4778) );
  OAI21_X1 U5346 ( .B1(n9245), .B2(n4782), .A(n4405), .ZN(n4779) );
  NOR2_X1 U5347 ( .A1(n9245), .A2(n9261), .ZN(n4780) );
  INV_X1 U5348 ( .A(n5450), .ZN(n5057) );
  NAND2_X1 U5349 ( .A1(n9295), .A2(n5034), .ZN(n9282) );
  NOR2_X1 U5350 ( .A1(n8043), .A2(n7957), .ZN(n5034) );
  NAND2_X1 U5351 ( .A1(n9297), .A2(n9296), .ZN(n9295) );
  OR2_X1 U5352 ( .A1(n9340), .A2(n9357), .ZN(n9307) );
  INV_X1 U5353 ( .A(n7851), .ZN(n9331) );
  NAND2_X1 U5354 ( .A1(n5036), .A2(n5035), .ZN(n9359) );
  AND2_X1 U5355 ( .A1(n9343), .A2(n7978), .ZN(n5035) );
  OR2_X1 U5356 ( .A1(n5707), .A2(n5706), .ZN(n5708) );
  NAND2_X1 U5357 ( .A1(n5289), .A2(n5013), .ZN(n7209) );
  NOR2_X1 U5358 ( .A1(n8039), .A2(n5014), .ZN(n5013) );
  NAND2_X1 U5359 ( .A1(n7014), .A2(n7972), .ZN(n5289) );
  INV_X1 U5360 ( .A(n8036), .ZN(n9963) );
  AND2_X1 U5361 ( .A1(n7828), .A2(n7995), .ZN(n8034) );
  OAI21_X1 U5362 ( .B1(n7819), .B2(n5230), .A(n8074), .ZN(n6801) );
  NAND2_X1 U5363 ( .A1(n6801), .A2(n8034), .ZN(n6800) );
  OR2_X1 U5364 ( .A1(n7936), .A2(n6380), .ZN(n10010) );
  OR2_X1 U5365 ( .A1(n7936), .A2(n9874), .ZN(n10012) );
  OR2_X1 U5366 ( .A1(n6388), .A2(n6529), .ZN(n6740) );
  NAND2_X1 U5367 ( .A1(n5579), .A2(n5578), .ZN(n9408) );
  XNOR2_X1 U5368 ( .A(n7803), .B(n7802), .ZN(n8876) );
  NAND2_X1 U5369 ( .A1(n7799), .A2(n7798), .ZN(n7803) );
  XNOR2_X1 U5370 ( .A(n5572), .B(n5571), .ZN(n7544) );
  NAND2_X1 U5371 ( .A1(n4896), .A2(n5552), .ZN(n5572) );
  NAND2_X1 U5372 ( .A1(n4897), .A2(n5549), .ZN(n4896) );
  INV_X1 U5373 ( .A(n5554), .ZN(n4897) );
  XNOR2_X1 U5374 ( .A(n5074), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U5375 ( .A1(n5098), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5074) );
  INV_X1 U5376 ( .A(n5509), .ZN(n4903) );
  INV_X1 U5377 ( .A(n4902), .ZN(n4901) );
  OAI21_X1 U5378 ( .B1(n4905), .B2(n4475), .A(n5523), .ZN(n4902) );
  NAND2_X1 U5379 ( .A1(n4904), .A2(n5509), .ZN(n5525) );
  NAND2_X1 U5380 ( .A1(n5497), .A2(n4905), .ZN(n4904) );
  NAND2_X1 U5381 ( .A1(n4862), .A2(n5440), .ZN(n5459) );
  NAND2_X1 U5382 ( .A1(n5423), .A2(n4866), .ZN(n4862) );
  NAND2_X1 U5383 ( .A1(n5423), .A2(n5422), .ZN(n5442) );
  NAND2_X1 U5384 ( .A1(n4910), .A2(n4915), .ZN(n5367) );
  XNOR2_X1 U5385 ( .A(n5331), .B(n5327), .ZN(n6315) );
  XNOR2_X1 U5386 ( .A(n5172), .B(SI_2_), .ZN(n5170) );
  AND2_X1 U5387 ( .A1(n7300), .A2(n7299), .ZN(n7302) );
  NAND2_X1 U5388 ( .A1(n5739), .A2(n5738), .ZN(n8798) );
  NAND2_X1 U5389 ( .A1(n4848), .A2(n4849), .ZN(n8167) );
  AOI21_X1 U5390 ( .B1(n4851), .B2(n4853), .A(n4433), .ZN(n4849) );
  NOR2_X1 U5391 ( .A1(n4568), .A2(n4570), .ZN(n4564) );
  NOR2_X1 U5392 ( .A1(n8183), .A2(n4571), .ZN(n4570) );
  INV_X1 U5393 ( .A(n8180), .ZN(n4567) );
  NAND2_X1 U5394 ( .A1(n4829), .A2(n4827), .ZN(n8175) );
  AOI21_X1 U5395 ( .B1(n4830), .B2(n4833), .A(n4828), .ZN(n4827) );
  NAND2_X1 U5396 ( .A1(n8198), .A2(n4830), .ZN(n4829) );
  INV_X1 U5397 ( .A(n8148), .ZN(n4828) );
  NAND2_X1 U5398 ( .A1(n5935), .A2(n5934), .ZN(n10295) );
  NAND2_X1 U5399 ( .A1(n7535), .A2(n4585), .ZN(n7537) );
  NAND2_X1 U5400 ( .A1(n7533), .A2(n7532), .ZN(n7535) );
  NAND2_X1 U5401 ( .A1(n7447), .A2(n4586), .ZN(n4585) );
  AND2_X1 U5402 ( .A1(n7534), .A2(n7446), .ZN(n4586) );
  NAND2_X1 U5403 ( .A1(n6860), .A2(n6213), .ZN(n6217) );
  NAND2_X1 U5404 ( .A1(n4847), .A2(n4846), .ZN(n4845) );
  NAND2_X1 U5405 ( .A1(n4843), .A2(n4845), .ZN(n6915) );
  INV_X1 U5406 ( .A(n4844), .ZN(n4843) );
  AND2_X1 U5407 ( .A1(n6223), .A2(n6222), .ZN(n8242) );
  NAND2_X1 U5408 ( .A1(n4837), .A2(n4834), .ZN(n4841) );
  NAND2_X1 U5409 ( .A1(n8235), .A2(n8236), .ZN(n4706) );
  NAND2_X1 U5410 ( .A1(n4837), .A2(n4836), .ZN(n8235) );
  NAND2_X1 U5411 ( .A1(n8783), .A2(n8228), .ZN(n4704) );
  NAND2_X1 U5412 ( .A1(n6461), .A2(n6462), .ZN(n6460) );
  NAND2_X1 U5413 ( .A1(n6519), .A2(n6520), .ZN(n6654) );
  XOR2_X1 U5414 ( .A(n8538), .B(n7743), .Z(n8535) );
  INV_X1 U5415 ( .A(n4977), .ZN(n4976) );
  INV_X1 U5416 ( .A(n8771), .ZN(n8181) );
  INV_X1 U5417 ( .A(n8426), .ZN(n7597) );
  NAND2_X1 U5418 ( .A1(n4984), .A2(n4982), .ZN(n7598) );
  INV_X1 U5419 ( .A(n4985), .ZN(n4982) );
  AOI21_X1 U5420 ( .B1(n7608), .B2(n10193), .A(n7607), .ZN(n8774) );
  NAND2_X1 U5421 ( .A1(n10222), .A2(n6903), .ZN(n10200) );
  NAND2_X1 U5422 ( .A1(n7764), .A2(n4497), .ZN(n6185) );
  INV_X1 U5423 ( .A(n6149), .ZN(n7764) );
  AND2_X1 U5424 ( .A1(n4732), .A2(n4734), .ZN(n4497) );
  NAND2_X1 U5425 ( .A1(n7766), .A2(n8852), .ZN(n4734) );
  NAND2_X1 U5426 ( .A1(n5371), .A2(n5370), .ZN(n9351) );
  NAND2_X1 U5427 ( .A1(n5468), .A2(n5467), .ZN(n9442) );
  NAND4_X1 U5428 ( .A1(n5326), .A2(n5325), .A3(n5324), .A4(n5323), .ZN(n9032)
         );
  AND2_X1 U5429 ( .A1(n5153), .A2(n5168), .ZN(n9860) );
  OAI21_X1 U5430 ( .B1(n9104), .B2(n9944), .A(n4656), .ZN(n4655) );
  OR2_X1 U5431 ( .A1(n9106), .A2(n9907), .ZN(n4656) );
  OAI21_X1 U5432 ( .B1(n9109), .B2(n9108), .A(n9107), .ZN(n4651) );
  OAI21_X1 U5433 ( .B1(n9942), .B2(n4511), .A(n9110), .ZN(n4653) );
  INV_X1 U5434 ( .A(n9321), .ZN(n9387) );
  OAI21_X1 U5435 ( .B1(n4727), .B2(n4398), .A(n5143), .ZN(n4726) );
  NOR2_X1 U5436 ( .A1(n6269), .A2(n7800), .ZN(n4727) );
  NAND2_X1 U5437 ( .A1(n5111), .A2(n10099), .ZN(n9994) );
  INV_X1 U5438 ( .A(n10029), .ZN(n9350) );
  INV_X1 U5439 ( .A(n4501), .ZN(n4500) );
  OAI21_X1 U5440 ( .B1(n9395), .B2(n9823), .A(n9393), .ZN(n4501) );
  XNOR2_X1 U5441 ( .A(n5108), .B(n5071), .ZN(n8092) );
  NAND2_X1 U5442 ( .A1(n4523), .A2(n4521), .ZN(n8289) );
  NAND2_X1 U5443 ( .A1(n8403), .A2(n8380), .ZN(n4523) );
  OAI21_X1 U5444 ( .B1(n7836), .B2(n8039), .A(n7835), .ZN(n7838) );
  MUX2_X1 U5445 ( .A(n7834), .B(n7833), .S(n7920), .Z(n7836) );
  OAI21_X1 U5446 ( .B1(n4431), .B2(n4519), .A(n4516), .ZN(n8308) );
  AND2_X1 U5447 ( .A1(n8297), .A2(n4517), .ZN(n4516) );
  AOI21_X1 U5448 ( .B1(n8287), .B2(n8286), .A(n4520), .ZN(n4519) );
  OR2_X1 U5449 ( .A1(n4538), .A2(n4471), .ZN(n4534) );
  OR2_X1 U5450 ( .A1(n4540), .A2(n4468), .ZN(n4535) );
  OAI21_X1 U5451 ( .B1(n8316), .B2(n8305), .A(n8380), .ZN(n4540) );
  OAI21_X1 U5452 ( .B1(n8316), .B2(n8313), .A(n8393), .ZN(n4538) );
  OR2_X1 U5453 ( .A1(n7875), .A2(n7862), .ZN(n7877) );
  INV_X1 U5454 ( .A(n4547), .ZN(n4546) );
  OAI21_X1 U5455 ( .B1(n4548), .B2(n4551), .A(n4448), .ZN(n4547) );
  NOR2_X1 U5456 ( .A1(n8348), .A2(n4482), .ZN(n4551) );
  AND2_X1 U5457 ( .A1(n4533), .A2(n4529), .ZN(n4528) );
  OR2_X1 U5458 ( .A1(n4531), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U5459 ( .A1(n7902), .A2(n4504), .ZN(n7914) );
  NOR2_X1 U5460 ( .A1(n4505), .A2(n4422), .ZN(n4504) );
  AOI21_X1 U5461 ( .B1(n4546), .B2(n4548), .A(n4545), .ZN(n4544) );
  INV_X1 U5462 ( .A(n8615), .ZN(n4545) );
  NAND2_X1 U5463 ( .A1(n8135), .A2(n8206), .ZN(n4699) );
  AOI21_X1 U5464 ( .B1(n4557), .B2(n4555), .A(n8379), .ZN(n4554) );
  INV_X1 U5465 ( .A(n4558), .ZN(n4555) );
  OR2_X1 U5466 ( .A1(n7759), .A2(n6118), .ZN(n8387) );
  INV_X1 U5467 ( .A(n8455), .ZN(n6095) );
  AND2_X1 U5468 ( .A1(n5834), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5851) );
  NAND2_X1 U5469 ( .A1(n8288), .A2(n6950), .ZN(n4522) );
  INV_X1 U5470 ( .A(n4640), .ZN(n4639) );
  OAI21_X1 U5471 ( .B1(n4945), .B2(n4641), .A(n8921), .ZN(n4640) );
  INV_X1 U5472 ( .A(n8971), .ZN(n4641) );
  NAND2_X1 U5473 ( .A1(n7793), .A2(n4410), .ZN(n8026) );
  NAND2_X1 U5474 ( .A1(n4931), .A2(n4929), .ZN(n4928) );
  NAND2_X1 U5475 ( .A1(n7809), .A2(n7933), .ZN(n4931) );
  NOR2_X1 U5476 ( .A1(n7919), .A2(n4930), .ZN(n4929) );
  AND2_X1 U5477 ( .A1(n9408), .A2(n9176), .ZN(n8013) );
  OR2_X1 U5478 ( .A1(n5702), .A2(n9372), .ZN(n5704) );
  AND2_X1 U5479 ( .A1(n8048), .A2(n5028), .ZN(n5026) );
  NAND2_X1 U5480 ( .A1(n4868), .A2(n4869), .ZN(n7797) );
  AOI21_X1 U5481 ( .B1(n4875), .B2(n4870), .A(n4411), .ZN(n4869) );
  INV_X1 U5482 ( .A(n5537), .ZN(n4899) );
  AOI21_X1 U5483 ( .B1(n4915), .B2(n4913), .A(n4912), .ZN(n4911) );
  INV_X1 U5484 ( .A(n5047), .ZN(n4912) );
  INV_X1 U5485 ( .A(n4917), .ZN(n4913) );
  INV_X1 U5486 ( .A(n4915), .ZN(n4914) );
  NAND2_X1 U5487 ( .A1(n5296), .A2(n5295), .ZN(n5313) );
  INV_X1 U5488 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n4942) );
  NAND2_X1 U5489 ( .A1(n4840), .A2(n4839), .ZN(n4838) );
  INV_X1 U5490 ( .A(n8195), .ZN(n4839) );
  INV_X1 U5491 ( .A(n8196), .ZN(n4840) );
  INV_X1 U5492 ( .A(n8187), .ZN(n4688) );
  INV_X1 U5493 ( .A(n8206), .ZN(n4700) );
  OAI21_X1 U5494 ( .B1(n4702), .B2(n4419), .A(n4838), .ZN(n4697) );
  OR2_X1 U5495 ( .A1(n4419), .A2(n8155), .ZN(n4695) );
  NAND2_X1 U5496 ( .A1(n8387), .A2(n8386), .ZN(n8428) );
  NAND2_X1 U5497 ( .A1(n4769), .A2(n8259), .ZN(n4766) );
  INV_X1 U5498 ( .A(n4769), .ZN(n4767) );
  OR2_X1 U5499 ( .A1(n8771), .A2(n6147), .ZN(n8382) );
  NOR2_X1 U5500 ( .A1(n8809), .A2(n4741), .ZN(n4740) );
  INV_X1 U5501 ( .A(n4742), .ZN(n4741) );
  NOR2_X1 U5502 ( .A1(n8814), .A2(n8823), .ZN(n4742) );
  OR2_X1 U5503 ( .A1(n5960), .A2(n9683), .ZN(n5974) );
  NAND2_X1 U5504 ( .A1(n4606), .A2(n8330), .ZN(n4605) );
  NAND2_X1 U5505 ( .A1(n7492), .A2(n8328), .ZN(n4606) );
  NAND2_X1 U5506 ( .A1(n5741), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5960) );
  INV_X1 U5507 ( .A(n5951), .ZN(n5741) );
  NAND2_X1 U5508 ( .A1(n5740), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5951) );
  INV_X1 U5509 ( .A(n5937), .ZN(n5740) );
  OAI21_X1 U5510 ( .B1(n8411), .B2(n4611), .A(n8321), .ZN(n4610) );
  INV_X1 U5511 ( .A(n4965), .ZN(n4964) );
  OAI21_X1 U5512 ( .B1(n5914), .B2(n4966), .A(n8414), .ZN(n4965) );
  INV_X1 U5513 ( .A(n5916), .ZN(n4966) );
  INV_X1 U5514 ( .A(n4522), .ZN(n8405) );
  NOR2_X1 U5515 ( .A1(n10217), .A2(n6200), .ZN(n10197) );
  NAND2_X1 U5516 ( .A1(n4592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4591) );
  NOR2_X1 U5517 ( .A1(n5009), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n5008) );
  NAND2_X1 U5518 ( .A1(n6161), .A2(n5010), .ZN(n5009) );
  NAND2_X1 U5519 ( .A1(n4938), .A2(n6688), .ZN(n4936) );
  INV_X1 U5520 ( .A(n6683), .ZN(n4938) );
  NOR2_X1 U5521 ( .A1(n7936), .A2(n8092), .ZN(n4925) );
  NAND2_X1 U5522 ( .A1(n4719), .A2(n4718), .ZN(n4717) );
  OR2_X1 U5523 ( .A1(n9392), .A2(n9123), .ZN(n8020) );
  INV_X1 U5524 ( .A(n8013), .ZN(n5589) );
  OR2_X1 U5525 ( .A1(n9408), .A2(n9176), .ZN(n7940) );
  AOI21_X1 U5526 ( .B1(n5019), .B2(n5021), .A(n5017), .ZN(n5016) );
  INV_X1 U5527 ( .A(n5020), .ZN(n5019) );
  AND2_X1 U5528 ( .A1(n4723), .A2(n4724), .ZN(n4722) );
  NOR2_X1 U5529 ( .A1(n9973), .A2(n9968), .ZN(n4708) );
  INV_X1 U5530 ( .A(n4809), .ZN(n6738) );
  NAND2_X1 U5531 ( .A1(n9252), .A2(n9237), .ZN(n9236) );
  INV_X1 U5532 ( .A(n4708), .ZN(n9974) );
  INV_X1 U5533 ( .A(n7095), .ZN(n6786) );
  NAND2_X1 U5534 ( .A1(n10022), .A2(n10087), .ZN(n9999) );
  INV_X1 U5535 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5095) );
  NOR2_X1 U5536 ( .A1(n5510), .A2(n4906), .ZN(n4905) );
  INV_X1 U5537 ( .A(n5496), .ZN(n4906) );
  NAND2_X1 U5538 ( .A1(n4861), .A2(n4860), .ZN(n5477) );
  AOI21_X1 U5539 ( .B1(n4863), .B2(n4865), .A(n4485), .ZN(n4860) );
  NOR2_X1 U5540 ( .A1(n5441), .A2(n4867), .ZN(n4866) );
  INV_X1 U5541 ( .A(n5422), .ZN(n4867) );
  AOI21_X1 U5542 ( .B1(n4919), .B2(n4917), .A(n4916), .ZN(n4915) );
  INV_X1 U5543 ( .A(n5349), .ZN(n4916) );
  NAND2_X1 U5544 ( .A1(n5329), .A2(SI_11_), .ZN(n5330) );
  NAND2_X1 U5545 ( .A1(n5349), .A2(n5335), .ZN(n5350) );
  INV_X1 U5546 ( .A(n5327), .ZN(n4919) );
  NAND2_X1 U5547 ( .A1(n5290), .A2(n5046), .ZN(n5292) );
  INV_X1 U5548 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5064) );
  INV_X1 U5549 ( .A(n5174), .ZN(n4513) );
  NAND2_X1 U5550 ( .A1(n5134), .A2(n5132), .ZN(n5133) );
  AND2_X1 U5551 ( .A1(n4826), .A2(n6770), .ZN(n4825) );
  INV_X1 U5552 ( .A(n6776), .ZN(n4826) );
  NAND2_X1 U5553 ( .A1(n4580), .A2(n4576), .ZN(n4575) );
  OR2_X1 U5554 ( .A1(n8230), .A2(n4572), .ZN(n4574) );
  NAND2_X1 U5555 ( .A1(n4577), .A2(n4573), .ZN(n4572) );
  INV_X1 U5556 ( .A(n8128), .ZN(n4573) );
  INV_X1 U5557 ( .A(n4852), .ZN(n4851) );
  OAI21_X1 U5558 ( .B1(n4854), .B2(n4853), .A(n8108), .ZN(n4852) );
  INV_X1 U5559 ( .A(n4856), .ZN(n4853) );
  INV_X1 U5560 ( .A(n8174), .ZN(n4571) );
  AOI21_X1 U5561 ( .B1(n4832), .B2(n4834), .A(n4831), .ZN(n4830) );
  INV_X1 U5562 ( .A(n8147), .ZN(n4831) );
  INV_X1 U5563 ( .A(n4838), .ZN(n4832) );
  INV_X1 U5564 ( .A(n4834), .ZN(n4833) );
  AND2_X1 U5565 ( .A1(n6724), .A2(n6195), .ZN(n10140) );
  NAND2_X1 U5566 ( .A1(n5742), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5976) );
  INV_X1 U5567 ( .A(n5974), .ZN(n5742) );
  NAND2_X1 U5568 ( .A1(n8119), .A2(n8118), .ZN(n8164) );
  AND2_X1 U5569 ( .A1(n8659), .A2(n6204), .ZN(n8128) );
  NAND2_X1 U5570 ( .A1(n5746), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6043) );
  NAND3_X1 U5571 ( .A1(n10138), .A2(n6203), .A3(n6199), .ZN(n4844) );
  NOR2_X1 U5572 ( .A1(n7579), .A2(n4855), .ZN(n4854) );
  INV_X1 U5573 ( .A(n7564), .ZN(n4855) );
  OR2_X1 U5574 ( .A1(n7578), .A2(n7577), .ZN(n4856) );
  NAND2_X1 U5575 ( .A1(n8196), .A2(n8195), .ZN(n4836) );
  CLKBUF_X1 U5576 ( .A(n6290), .Z(n6114) );
  OR2_X1 U5577 ( .A1(n5888), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5903) );
  AND2_X1 U5578 ( .A1(n7136), .A2(n7135), .ZN(n8505) );
  INV_X1 U5579 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5727) );
  AND2_X1 U5580 ( .A1(n5725), .A2(n4960), .ZN(n4817) );
  OAI21_X1 U5581 ( .B1(n7521), .B2(n7520), .A(n7519), .ZN(n8512) );
  AND2_X1 U5582 ( .A1(n8516), .A2(n7508), .ZN(n7511) );
  OAI21_X1 U5583 ( .B1(n4981), .B2(n4393), .A(n4979), .ZN(n4977) );
  AOI21_X1 U5584 ( .B1(n4983), .B2(n4980), .A(n4456), .ZN(n4979) );
  INV_X1 U5585 ( .A(n4988), .ZN(n4980) );
  NOR2_X1 U5586 ( .A1(n4981), .A2(n8587), .ZN(n4978) );
  NAND2_X1 U5587 ( .A1(n4987), .A2(n4986), .ZN(n4985) );
  NAND2_X1 U5588 ( .A1(n4988), .A2(n8573), .ZN(n4987) );
  NAND2_X1 U5589 ( .A1(n4461), .A2(n4989), .ZN(n4986) );
  NAND2_X1 U5590 ( .A1(n4613), .A2(n4763), .ZN(n7604) );
  AOI21_X1 U5591 ( .B1(n4765), .B2(n4767), .A(n4764), .ZN(n4763) );
  NAND2_X1 U5592 ( .A1(n8588), .A2(n4765), .ZN(n4613) );
  INV_X1 U5593 ( .A(n8377), .ZN(n4764) );
  AND2_X1 U5594 ( .A1(n8382), .A2(n8381), .ZN(n8426) );
  NAND2_X1 U5595 ( .A1(n4991), .A2(n8151), .ZN(n4990) );
  NAND2_X1 U5596 ( .A1(n6063), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6075) );
  NAND2_X1 U5597 ( .A1(n8616), .A2(n4614), .ZN(n8610) );
  AND2_X1 U5598 ( .A1(n8605), .A2(n8606), .ZN(n4614) );
  AOI21_X1 U5599 ( .B1(n4995), .B2(n4994), .A(n5001), .ZN(n4993) );
  AND2_X1 U5600 ( .A1(n8798), .A2(n8457), .ZN(n5001) );
  NAND2_X1 U5601 ( .A1(n8365), .A2(n8369), .ZN(n8596) );
  AND2_X1 U5602 ( .A1(n6139), .A2(n4598), .ZN(n4597) );
  AND2_X1 U5603 ( .A1(n8637), .A2(n8638), .ZN(n6139) );
  NAND2_X1 U5604 ( .A1(n8695), .A2(n4740), .ZN(n8649) );
  NAND2_X1 U5605 ( .A1(n8695), .A2(n8689), .ZN(n8679) );
  OR2_X1 U5606 ( .A1(n5976), .A2(n5765), .ZN(n5986) );
  NAND2_X1 U5607 ( .A1(n5743), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6000) );
  INV_X1 U5608 ( .A(n5986), .ZN(n5743) );
  NAND2_X1 U5609 ( .A1(n8746), .A2(n8340), .ZN(n8718) );
  OR2_X1 U5610 ( .A1(n5923), .A2(n5922), .ZN(n5937) );
  INV_X1 U5611 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8487) );
  OR2_X1 U5612 ( .A1(n5907), .A2(n8487), .ZN(n5923) );
  NAND2_X1 U5613 ( .A1(n6134), .A2(n4443), .ZN(n4607) );
  INV_X1 U5614 ( .A(n8410), .ZN(n5900) );
  AND2_X1 U5615 ( .A1(n8310), .A2(n8314), .ZN(n8410) );
  OAI21_X1 U5616 ( .B1(n6134), .B2(n4745), .A(n4744), .ZN(n7230) );
  NAND2_X1 U5617 ( .A1(n5879), .A2(n4494), .ZN(n6992) );
  NAND2_X1 U5618 ( .A1(n6279), .A2(n8249), .ZN(n4494) );
  INV_X1 U5619 ( .A(n4737), .ZN(n7240) );
  NAND2_X1 U5620 ( .A1(n5850), .A2(n5849), .ZN(n6975) );
  NAND2_X1 U5621 ( .A1(n8298), .A2(n8294), .ZN(n8407) );
  NAND2_X1 U5622 ( .A1(n4738), .A2(n10262), .ZN(n6947) );
  INV_X1 U5623 ( .A(n10196), .ZN(n4738) );
  NAND2_X1 U5624 ( .A1(n4755), .A2(n8266), .ZN(n10174) );
  NAND2_X1 U5625 ( .A1(n4753), .A2(n10187), .ZN(n4755) );
  NAND2_X1 U5626 ( .A1(n10197), .A2(n10256), .ZN(n10196) );
  AND2_X1 U5627 ( .A1(n7759), .A2(n8851), .ZN(n4733) );
  NAND2_X1 U5628 ( .A1(n6084), .A2(n6083), .ZN(n8777) );
  AND2_X1 U5629 ( .A1(n4997), .A2(n4995), .ZN(n8803) );
  NAND2_X1 U5630 ( .A1(n5005), .A2(n4395), .ZN(n8714) );
  AND2_X1 U5631 ( .A1(n5005), .A2(n5004), .ZN(n8715) );
  AND2_X1 U5632 ( .A1(n5006), .A2(n5750), .ZN(n4593) );
  AND2_X1 U5633 ( .A1(n5008), .A2(n5748), .ZN(n5006) );
  INV_X1 U5634 ( .A(n5009), .ZN(n5007) );
  OAI21_X1 U5635 ( .B1(n6127), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6164) );
  OR2_X1 U5636 ( .A1(n5903), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n5917) );
  NAND2_X1 U5637 ( .A1(n5060), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5638 ( .A1(n6878), .A2(n4403), .ZN(n6886) );
  INV_X1 U5639 ( .A(n6883), .ZN(n4940) );
  NOR2_X1 U5640 ( .A1(n5048), .A2(n5042), .ZN(n7402) );
  NAND2_X1 U5641 ( .A1(n7395), .A2(n7394), .ZN(n4944) );
  NAND2_X1 U5642 ( .A1(n9012), .A2(n9015), .ZN(n4939) );
  NAND2_X1 U5643 ( .A1(n5056), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5429) );
  INV_X1 U5644 ( .A(n5414), .ZN(n5056) );
  NAND2_X1 U5645 ( .A1(n6590), .A2(n6591), .ZN(n6684) );
  NAND2_X1 U5646 ( .A1(n8911), .A2(n8912), .ZN(n4949) );
  OR2_X1 U5647 ( .A1(n5341), .A2(n5340), .ZN(n5361) );
  NAND2_X1 U5648 ( .A1(n4944), .A2(n4943), .ZN(n7468) );
  OR2_X1 U5649 ( .A1(n5429), .A2(n8953), .ZN(n5450) );
  OR3_X1 U5650 ( .A1(n6577), .A2(n8099), .A3(n10072), .ZN(n6503) );
  OR2_X1 U5651 ( .A1(n8931), .A2(n4629), .ZN(n4628) );
  NOR2_X1 U5652 ( .A1(n4447), .A2(n9025), .ZN(n4627) );
  NAND2_X1 U5653 ( .A1(n8101), .A2(n8092), .ZN(n6734) );
  NAND2_X1 U5654 ( .A1(n5114), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5130) );
  INV_X1 U5655 ( .A(n5582), .ZN(n5630) );
  NAND4_X1 U5656 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n6492)
         );
  NAND2_X1 U5657 ( .A1(n5178), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5122) );
  NOR3_X1 U5658 ( .A1(n6311), .A2(n6389), .A3(n9852), .ZN(n9851) );
  AOI22_X1 U5659 ( .A1(n9879), .A2(n9878), .B1(n6330), .B2(n6329), .ZN(n9895)
         );
  AND2_X1 U5660 ( .A1(n9895), .A2(n9894), .ZN(n9897) );
  NAND2_X1 U5661 ( .A1(n6343), .A2(n6342), .ZN(n6341) );
  NOR2_X1 U5662 ( .A1(n9909), .A2(n9910), .ZN(n9908) );
  NAND2_X1 U5663 ( .A1(n6599), .A2(n4476), .ZN(n9931) );
  AND2_X1 U5664 ( .A1(n4670), .A2(n4669), .ZN(n9934) );
  NAND2_X1 U5665 ( .A1(n6607), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5666 ( .A1(n9934), .A2(n9935), .ZN(n9933) );
  OR2_X1 U5667 ( .A1(n6647), .A2(n6646), .ZN(n4663) );
  NAND2_X1 U5668 ( .A1(n6999), .A2(n4489), .ZN(n7000) );
  AND2_X1 U5669 ( .A1(n4663), .A2(n4662), .ZN(n9041) );
  NAND2_X1 U5670 ( .A1(n7006), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4662) );
  NAND2_X1 U5671 ( .A1(n7808), .A2(n7807), .ZN(n7938) );
  NAND2_X1 U5672 ( .A1(n5622), .A2(n7917), .ZN(n9125) );
  AND2_X1 U5673 ( .A1(n8012), .A2(n5604), .ZN(n9136) );
  NAND2_X1 U5674 ( .A1(n7940), .A2(n5589), .ZN(n9162) );
  NAND2_X1 U5675 ( .A1(n9252), .A2(n4709), .ZN(n9188) );
  AND2_X1 U5676 ( .A1(n4400), .A2(n5716), .ZN(n4709) );
  OAI21_X1 U5677 ( .B1(n9182), .B2(n4796), .A(n4795), .ZN(n4794) );
  AND2_X1 U5678 ( .A1(n9419), .A2(n9204), .ZN(n4796) );
  NAND2_X1 U5679 ( .A1(n5716), .A2(n9175), .ZN(n4795) );
  NAND2_X1 U5680 ( .A1(n9252), .A2(n4711), .ZN(n9220) );
  OR2_X1 U5681 ( .A1(n5488), .A2(n5058), .ZN(n5500) );
  AND2_X1 U5682 ( .A1(n9346), .A2(n4720), .ZN(n9277) );
  NOR2_X1 U5683 ( .A1(n9447), .A2(n4721), .ZN(n4720) );
  INV_X1 U5684 ( .A(n4722), .ZN(n4721) );
  NAND2_X1 U5685 ( .A1(n9346), .A2(n9832), .ZN(n9337) );
  NAND2_X1 U5686 ( .A1(n9346), .A2(n4724), .ZN(n9314) );
  NAND2_X1 U5687 ( .A1(n5420), .A2(n4785), .ZN(n9309) );
  NAND2_X1 U5688 ( .A1(n5055), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5396) );
  INV_X1 U5689 ( .A(n5361), .ZN(n5055) );
  OR3_X1 U5690 ( .A1(n5396), .A2(n5395), .A3(n8894), .ZN(n5414) );
  NAND2_X1 U5691 ( .A1(n9330), .A2(n9331), .ZN(n9329) );
  NAND2_X1 U5692 ( .A1(n5036), .A2(n7978), .ZN(n9355) );
  AND2_X1 U5693 ( .A1(n9379), .A2(n9840), .ZN(n9346) );
  INV_X1 U5694 ( .A(n9365), .ZN(n9372) );
  NOR2_X1 U5695 ( .A1(n9377), .A2(n9457), .ZN(n9379) );
  NAND2_X1 U5696 ( .A1(n5348), .A2(n7976), .ZN(n9366) );
  AND2_X1 U5697 ( .A1(n7847), .A2(n7978), .ZN(n9365) );
  OR2_X1 U5698 ( .A1(n7436), .A2(n9464), .ZN(n9377) );
  NAND2_X1 U5699 ( .A1(n5054), .A2(n5053), .ZN(n5321) );
  INV_X1 U5700 ( .A(n7837), .ZN(n8040) );
  NAND2_X1 U5701 ( .A1(n7272), .A2(n7275), .ZN(n7436) );
  AND2_X1 U5702 ( .A1(n7431), .A2(n7839), .ZN(n7837) );
  NAND2_X1 U5703 ( .A1(n4708), .A2(n4707), .ZN(n7211) );
  NOR2_X1 U5704 ( .A1(n7211), .A2(n7326), .ZN(n7272) );
  NOR2_X1 U5705 ( .A1(n4807), .A2(n4806), .ZN(n4805) );
  INV_X1 U5706 ( .A(n5697), .ZN(n4806) );
  AND2_X1 U5707 ( .A1(n7104), .A2(n6786), .ZN(n6803) );
  OR2_X1 U5708 ( .A1(n9999), .A2(n9998), .ZN(n10001) );
  NOR2_X1 U5709 ( .A1(n10001), .A2(n7102), .ZN(n7104) );
  NAND2_X1 U5710 ( .A1(n8067), .A2(n5195), .ZN(n5012) );
  NOR2_X1 U5711 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  INV_X1 U5712 ( .A(n10012), .ZN(n9987) );
  AND2_X1 U5713 ( .A1(n4425), .A2(n9129), .ZN(n9397) );
  NAND2_X1 U5714 ( .A1(n9202), .A2(n5028), .ZN(n5022) );
  OR2_X1 U5715 ( .A1(n7933), .A2(n5653), .ZN(n9473) );
  AND2_X1 U5716 ( .A1(n10070), .A2(n5676), .ZN(n6525) );
  INV_X1 U5717 ( .A(n6863), .ZN(n6529) );
  OR3_X1 U5718 ( .A1(n5661), .A2(n5660), .A3(n7573), .ZN(n10036) );
  XNOR2_X1 U5719 ( .A(n7595), .B(n5627), .ZN(n7733) );
  NAND2_X1 U5720 ( .A1(n4872), .A2(n4873), .ZN(n7595) );
  NAND2_X1 U5721 ( .A1(n5605), .A2(n4876), .ZN(n4872) );
  XNOR2_X1 U5722 ( .A(n5605), .B(n5606), .ZN(n7586) );
  NAND2_X1 U5723 ( .A1(n4887), .A2(n4891), .ZN(n5577) );
  OAI21_X1 U5724 ( .B1(n5554), .B2(n4890), .A(n4888), .ZN(n5591) );
  NAND2_X1 U5725 ( .A1(n5554), .A2(n4894), .ZN(n4887) );
  NAND2_X1 U5726 ( .A1(n5101), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5727 ( .A1(n5497), .A2(n5496), .ZN(n5511) );
  NAND2_X1 U5728 ( .A1(n5257), .A2(n4959), .ZN(n5299) );
  XNOR2_X1 U5729 ( .A(n5312), .B(n5039), .ZN(n6300) );
  NAND2_X1 U5730 ( .A1(n4880), .A2(n5244), .ZN(n5251) );
  XNOR2_X1 U5731 ( .A(n5215), .B(SI_5_), .ZN(n5213) );
  AND2_X1 U5732 ( .A1(n5063), .A2(n5062), .ZN(n5184) );
  NAND2_X1 U5733 ( .A1(n6819), .A2(n6770), .ZN(n6777) );
  INV_X1 U5734 ( .A(n4841), .ZN(n8234) );
  NAND2_X1 U5735 ( .A1(n5959), .A2(n5958), .ZN(n7484) );
  OAI21_X1 U5736 ( .B1(n8119), .B2(n4690), .A(n4689), .ZN(n8188) );
  INV_X1 U5737 ( .A(n6192), .ZN(n10270) );
  NAND2_X1 U5738 ( .A1(n7565), .A2(n7564), .ZN(n7580) );
  NAND2_X1 U5739 ( .A1(n6050), .A2(n6049), .ZN(n8792) );
  AND2_X1 U5740 ( .A1(n8242), .A2(n10189), .ZN(n10137) );
  AND2_X1 U5741 ( .A1(n6230), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8210) );
  NAND2_X1 U5742 ( .A1(n6916), .A2(n6209), .ZN(n6860) );
  AND2_X1 U5743 ( .A1(n8242), .A2(n10190), .ZN(n10136) );
  NAND2_X1 U5744 ( .A1(n8164), .A2(n8120), .ZN(n8216) );
  INV_X1 U5745 ( .A(n8210), .ZN(n8240) );
  NAND2_X1 U5746 ( .A1(n7031), .A2(n4582), .ZN(n7041) );
  OR2_X1 U5747 ( .A1(n7037), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U5748 ( .A1(n5920), .A2(n5919), .ZN(n7367) );
  NAND2_X1 U5749 ( .A1(n4850), .A2(n4856), .ZN(n8109) );
  NAND2_X1 U5750 ( .A1(n7565), .A2(n4854), .ZN(n4850) );
  NAND2_X1 U5751 ( .A1(n5997), .A2(n5996), .ZN(n8826) );
  INV_X1 U5752 ( .A(n6975), .ZN(n10275) );
  INV_X1 U5753 ( .A(n10136), .ZN(n8225) );
  INV_X1 U5754 ( .A(n10137), .ZN(n8224) );
  OAI211_X1 U5755 ( .C1(n4682), .C2(n7302), .A(n4681), .B(n4679), .ZN(n7533)
         );
  NAND2_X1 U5756 ( .A1(n4683), .A2(n7534), .ZN(n4682) );
  AND2_X1 U5757 ( .A1(n4680), .A2(n4685), .ZN(n4679) );
  NAND2_X1 U5758 ( .A1(n5971), .A2(n5970), .ZN(n8844) );
  XNOR2_X1 U5759 ( .A(n4752), .B(n8730), .ZN(n4751) );
  AOI21_X1 U5760 ( .B1(n8254), .B2(n8399), .A(n8395), .ZN(n4752) );
  NAND2_X1 U5761 ( .A1(n6204), .A2(n8255), .ZN(n4750) );
  NAND2_X1 U5762 ( .A1(n5921), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5797) );
  INV_X1 U5763 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5132) );
  NAND2_X1 U5764 ( .A1(n9794), .A2(n4438), .ZN(n9805) );
  NAND2_X1 U5765 ( .A1(n6460), .A2(n4435), .ZN(n6450) );
  NAND2_X1 U5766 ( .A1(n6654), .A2(n4481), .ZN(n8472) );
  NAND2_X1 U5767 ( .A1(n8484), .A2(n6657), .ZN(n6658) );
  AOI21_X1 U5768 ( .B1(n7128), .B2(n5925), .A(n7127), .ZN(n8499) );
  NAND2_X1 U5769 ( .A1(n4961), .A2(n5044), .ZN(n5932) );
  INV_X1 U5770 ( .A(n5843), .ZN(n4961) );
  AOI21_X1 U5771 ( .B1(n7133), .B2(n7497), .A(n10159), .ZN(n7132) );
  XNOR2_X1 U5772 ( .A(n4495), .B(n6016), .ZN(n7753) );
  NAND2_X1 U5773 ( .A1(n8534), .A2(n7744), .ZN(n4495) );
  AND2_X1 U5774 ( .A1(n6419), .A2(n6418), .ZN(n10151) );
  NAND2_X1 U5775 ( .A1(n8252), .A2(n8251), .ZN(n8762) );
  AOI21_X1 U5776 ( .B1(n7790), .B2(n8249), .A(n8244), .ZN(n8769) );
  NOR2_X1 U5777 ( .A1(n4768), .A2(n8372), .ZN(n8572) );
  INV_X1 U5778 ( .A(n4771), .ZN(n4768) );
  NAND2_X1 U5779 ( .A1(n7544), .A2(n8249), .ZN(n6062) );
  INV_X1 U5780 ( .A(n8792), .ZN(n6059) );
  NAND2_X1 U5781 ( .A1(n4997), .A2(n4998), .ZN(n8626) );
  AOI21_X1 U5782 ( .B1(n8648), .B2(n6038), .A(n4394), .ZN(n8630) );
  NAND2_X1 U5783 ( .A1(n4594), .A2(n4601), .ZN(n8657) );
  OR2_X1 U5784 ( .A1(n4602), .A2(n4603), .ZN(n4594) );
  NAND2_X1 U5785 ( .A1(n5985), .A2(n5984), .ZN(n8831) );
  NAND2_X1 U5786 ( .A1(n5764), .A2(n5763), .ZN(n8836) );
  NAND2_X1 U5787 ( .A1(n7477), .A2(n4761), .ZN(n7550) );
  NOR2_X1 U5788 ( .A1(n4760), .A2(n4762), .ZN(n7551) );
  NAND2_X1 U5789 ( .A1(n5948), .A2(n5947), .ZN(n8850) );
  NAND2_X1 U5790 ( .A1(n7178), .A2(n5916), .ZN(n7219) );
  NAND2_X1 U5791 ( .A1(n7184), .A2(n8312), .ZN(n7220) );
  OR2_X1 U5792 ( .A1(n8446), .A2(n6226), .ZN(n10218) );
  NAND2_X1 U5793 ( .A1(n4969), .A2(n4970), .ZN(n6987) );
  INV_X1 U5794 ( .A(n6134), .ZN(n6713) );
  NAND2_X1 U5795 ( .A1(n8272), .A2(n8276), .ZN(n6936) );
  INV_X1 U5796 ( .A(n10200), .ZN(n10183) );
  AND2_X1 U5797 ( .A1(n6295), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10240) );
  XNOR2_X1 U5798 ( .A(n6167), .B(P2_IR_REG_24__SCAN_IN), .ZN(n7455) );
  XNOR2_X1 U5799 ( .A(n6126), .B(n6125), .ZN(n8436) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9744) );
  OR2_X1 U5801 ( .A1(n4953), .A2(n4480), .ZN(n4951) );
  AND2_X1 U5802 ( .A1(n4649), .A2(n4648), .ZN(n8902) );
  NAND2_X1 U5803 ( .A1(n6568), .A2(n6569), .ZN(n6589) );
  NAND2_X1 U5804 ( .A1(n7664), .A2(n9004), .ZN(n4630) );
  NOR2_X1 U5805 ( .A1(n4635), .A2(n4633), .ZN(n4632) );
  NAND2_X1 U5806 ( .A1(n7776), .A2(n7775), .ZN(n7788) );
  NAND2_X1 U5807 ( .A1(n8968), .A2(n8971), .ZN(n8922) );
  NAND2_X1 U5808 ( .A1(n4944), .A2(n7402), .ZN(n7405) );
  NAND2_X2 U5809 ( .A1(n5560), .A2(n5559), .ZN(n9412) );
  NAND2_X1 U5810 ( .A1(n7544), .A2(n7804), .ZN(n5560) );
  NAND2_X1 U5811 ( .A1(n4939), .A2(n9013), .ZN(n8939) );
  INV_X1 U5812 ( .A(n9019), .ZN(n9005) );
  NAND2_X1 U5813 ( .A1(n4948), .A2(n4949), .ZN(n8970) );
  AND2_X1 U5814 ( .A1(n6382), .A2(n6381), .ZN(n8951) );
  NAND2_X1 U5815 ( .A1(n4636), .A2(n7663), .ZN(n9001) );
  NAND2_X1 U5816 ( .A1(n4634), .A2(n7664), .ZN(n9002) );
  INV_X1 U5817 ( .A(n4636), .ZN(n4634) );
  INV_X1 U5818 ( .A(n8951), .ZN(n9025) );
  AND2_X1 U5819 ( .A1(n6580), .A2(n6579), .ZN(n9021) );
  CLKBUF_X1 U5820 ( .A(n5641), .Z(n9869) );
  INV_X1 U5821 ( .A(n7934), .ZN(n8101) );
  NAND2_X1 U5822 ( .A1(n8094), .A2(n8093), .ZN(n4920) );
  NAND2_X1 U5823 ( .A1(n5203), .A2(n4623), .ZN(n9986) );
  NOR2_X1 U5824 ( .A1(n4429), .A2(n4624), .ZN(n4623) );
  OR2_X1 U5825 ( .A1(n5582), .A2(n9993), .ZN(n5181) );
  OR2_X1 U5826 ( .A1(n5179), .A2(n5144), .ZN(n5146) );
  NAND2_X1 U5827 ( .A1(n5178), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5148) );
  OR2_X1 U5828 ( .A1(n5452), .A2(n6865), .ZN(n5139) );
  NOR2_X1 U5829 ( .A1(n9863), .A2(n9862), .ZN(n9861) );
  NOR2_X1 U5830 ( .A1(n9866), .A2(n9865), .ZN(n9864) );
  NOR2_X1 U5831 ( .A1(n9849), .A2(n4659), .ZN(n9866) );
  INV_X1 U5832 ( .A(n6245), .ZN(n4659) );
  AND2_X1 U5833 ( .A1(n4661), .A2(n4660), .ZN(n6322) );
  NAND2_X1 U5834 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  NOR2_X1 U5835 ( .A1(n6348), .A2(n6349), .ZN(n6347) );
  NAND2_X1 U5836 ( .A1(n9891), .A2(n4668), .ZN(n6348) );
  OR2_X1 U5837 ( .A1(n9901), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n4668) );
  NOR2_X1 U5838 ( .A1(n6347), .A2(n4665), .ZN(n6323) );
  NOR2_X1 U5839 ( .A1(n4667), .A2(n4666), .ZN(n4665) );
  AND2_X1 U5840 ( .A1(n5262), .A2(n5261), .ZN(n9914) );
  INV_X1 U5841 ( .A(n4672), .ZN(n6370) );
  INV_X1 U5842 ( .A(n4670), .ZN(n6606) );
  NOR2_X1 U5843 ( .A1(n6642), .A2(n4664), .ZN(n6647) );
  AND2_X1 U5844 ( .A1(n6643), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4664) );
  INV_X1 U5845 ( .A(n4663), .ZN(n7005) );
  XNOR2_X1 U5846 ( .A(n9041), .B(n9040), .ZN(n7007) );
  INV_X1 U5847 ( .A(n4676), .ZN(n9056) );
  NOR2_X1 U5848 ( .A1(n9065), .A2(n9064), .ZN(n9070) );
  OAI21_X1 U5849 ( .B1(n9044), .B2(n4674), .A(n4673), .ZN(n9078) );
  NAND2_X1 U5850 ( .A1(n4677), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n4674) );
  NAND2_X1 U5851 ( .A1(n9057), .A2(n4677), .ZN(n4673) );
  INV_X1 U5852 ( .A(n9061), .ZN(n4677) );
  INV_X1 U5853 ( .A(n9057), .ZN(n4675) );
  AOI21_X1 U5854 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n9102), .A(n9101), .ZN(
        n9953) );
  INV_X1 U5855 ( .A(n7938), .ZN(n9390) );
  OAI21_X1 U5856 ( .B1(n4418), .B2(n9128), .A(n9127), .ZN(n9400) );
  NAND2_X1 U5857 ( .A1(n4800), .A2(n4396), .ZN(n9127) );
  INV_X1 U5858 ( .A(n9408), .ZN(n9159) );
  NAND2_X1 U5859 ( .A1(n5029), .A2(n7897), .ZN(n9183) );
  NAND2_X1 U5860 ( .A1(n5517), .A2(n5516), .ZN(n9427) );
  NAND2_X1 U5861 ( .A1(n4775), .A2(n4778), .ZN(n9233) );
  NAND2_X1 U5862 ( .A1(n4774), .A2(n4780), .ZN(n4775) );
  NAND2_X1 U5863 ( .A1(n5018), .A2(n8003), .ZN(n9246) );
  NAND2_X1 U5864 ( .A1(n9262), .A2(n9261), .ZN(n5018) );
  AOI21_X1 U5865 ( .B1(n4774), .B2(n9271), .A(n4781), .ZN(n9244) );
  NAND2_X1 U5866 ( .A1(n4783), .A2(n4787), .ZN(n9305) );
  NAND2_X1 U5867 ( .A1(n9344), .A2(n4790), .ZN(n4783) );
  NAND2_X1 U5868 ( .A1(n5412), .A2(n5411), .ZN(n9318) );
  NAND2_X1 U5869 ( .A1(n4792), .A2(n4790), .ZN(n9326) );
  NAND2_X1 U5870 ( .A1(n4792), .A2(n5710), .ZN(n9324) );
  NAND2_X1 U5871 ( .A1(n5289), .A2(n7967), .ZN(n7207) );
  NAND2_X1 U5872 ( .A1(n6800), .A2(n7995), .ZN(n9964) );
  OR3_X1 U5873 ( .A1(n9387), .A2(n6862), .A3(n8097), .ZN(n10032) );
  MUX2_X1 U5874 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9783), .S(n5143), .Z(n6863) );
  INV_X1 U5875 ( .A(n10032), .ZN(n10003) );
  AOI211_X1 U5876 ( .C1(n9822), .C2(n9821), .A(n9820), .B(n9819), .ZN(n9844)
         );
  NOR2_X1 U5877 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n5030) );
  XNOR2_X1 U5878 ( .A(n5624), .B(n5623), .ZN(n9778) );
  OAI21_X1 U5879 ( .B1(n5497), .B2(n4475), .A(n4901), .ZN(n5538) );
  INV_X1 U5880 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9730) );
  NAND2_X1 U5881 ( .A1(n4562), .A2(n5174), .ZN(n5190) );
  INV_X1 U5882 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9547) );
  XNOR2_X1 U5883 ( .A(n4678), .B(n5131), .ZN(n9856) );
  NAND2_X1 U5884 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4678) );
  NOR2_X1 U5885 ( .A1(n7360), .A2(n10356), .ZN(n10347) );
  NOR2_X1 U5886 ( .A1(n6398), .A2(n10234), .ZN(P2_U3966) );
  OAI211_X1 U5887 ( .C1(n8175), .C2(n4565), .A(n4563), .B(n4483), .ZN(P2_U3222) );
  NAND2_X1 U5888 ( .A1(n4566), .A2(n4567), .ZN(n4565) );
  NAND2_X1 U5889 ( .A1(n8175), .A2(n4564), .ZN(n4563) );
  AND2_X1 U5890 ( .A1(n4845), .A2(n6203), .ZN(n6622) );
  NAND2_X1 U5891 ( .A1(n4705), .A2(n4703), .ZN(P2_U3242) );
  AND2_X1 U5892 ( .A1(n8243), .A2(n4704), .ZN(n4703) );
  AOI21_X1 U5893 ( .B1(n4384), .B2(n10202), .A(n4616), .ZN(n4615) );
  INV_X1 U5894 ( .A(n4617), .ZN(n4616) );
  NOR2_X1 U5895 ( .A1(n8774), .A2(n10224), .ZN(n7609) );
  NAND2_X1 U5896 ( .A1(n10317), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U5897 ( .A1(n6185), .A2(n10319), .ZN(n4731) );
  INV_X1 U5898 ( .A(n4653), .ZN(n4652) );
  NAND2_X1 U5899 ( .A1(n4655), .A2(n8092), .ZN(n4654) );
  OAI21_X1 U5900 ( .B1(n9395), .B2(n9323), .A(n5720), .ZN(n5721) );
  NAND2_X1 U5901 ( .A1(n4499), .A2(n4498), .ZN(P1_U3552) );
  NAND2_X1 U5902 ( .A1(n10134), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U5903 ( .A1(n4408), .A2(n8134), .ZN(n4702) );
  OR2_X1 U5904 ( .A1(n8789), .A2(n8456), .ZN(n4393) );
  INV_X1 U5905 ( .A(n4773), .ZN(n4602) );
  AND2_X1 U5906 ( .A1(n8654), .A2(n8641), .ZN(n4394) );
  AND2_X1 U5907 ( .A1(n8717), .A2(n5004), .ZN(n4395) );
  AND2_X1 U5908 ( .A1(n9128), .A2(n4803), .ZN(n4396) );
  AND2_X1 U5909 ( .A1(n4702), .A2(n4444), .ZN(n4397) );
  INV_X1 U5910 ( .A(n7967), .ZN(n5014) );
  INV_X1 U5911 ( .A(n8419), .ZN(n4759) );
  INV_X1 U5912 ( .A(n7995), .ZN(n5032) );
  AND2_X1 U5913 ( .A1(n7800), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4398) );
  AND2_X1 U5914 ( .A1(n4691), .A2(n8187), .ZN(n4399) );
  NAND2_X1 U5915 ( .A1(n5629), .A2(n5628), .ZN(n9392) );
  INV_X1 U5916 ( .A(n9392), .ZN(n4718) );
  INV_X1 U5917 ( .A(n7885), .ZN(n4777) );
  AND2_X1 U5918 ( .A1(n4711), .A2(n4710), .ZN(n4400) );
  AND2_X1 U5919 ( .A1(n4740), .A2(n4739), .ZN(n4401) );
  OR2_X1 U5920 ( .A1(n7267), .A2(n7275), .ZN(n4402) );
  AND2_X1 U5921 ( .A1(n6877), .A2(n4940), .ZN(n4403) );
  OR2_X1 U5922 ( .A1(n6124), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n4404) );
  OR2_X1 U5923 ( .A1(n9255), .A2(n9230), .ZN(n4405) );
  OR2_X1 U5924 ( .A1(n8671), .A2(n8670), .ZN(n4406) );
  INV_X1 U5925 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5091) );
  OR2_X1 U5926 ( .A1(n4600), .A2(n4603), .ZN(n4407) );
  AND2_X1 U5927 ( .A1(n4580), .A2(n4579), .ZN(n4408) );
  AND3_X1 U5928 ( .A1(n4535), .A2(n4534), .A3(n4473), .ZN(n4409) );
  INV_X1 U5929 ( .A(n8039), .ZN(n4807) );
  AND2_X1 U5930 ( .A1(n4859), .A2(n7792), .ZN(n4410) );
  AND2_X1 U5931 ( .A1(n7593), .A2(SI_29_), .ZN(n4411) );
  INV_X2 U5932 ( .A(n6725), .ZN(n6204) );
  INV_X1 U5933 ( .A(n8136), .ZN(n8135) );
  OR2_X1 U5934 ( .A1(n4579), .A2(n8134), .ZN(n4412) );
  NAND2_X1 U5935 ( .A1(n9351), .A2(n9327), .ZN(n4413) );
  AND2_X1 U5936 ( .A1(n6700), .A2(n7089), .ZN(n4414) );
  AND2_X1 U5937 ( .A1(n8890), .A2(n7639), .ZN(n4415) );
  AND3_X1 U5938 ( .A1(n5796), .A2(n5795), .A3(n5794), .ZN(n4416) );
  OR2_X1 U5939 ( .A1(n5070), .A2(n5069), .ZN(n4417) );
  AND2_X1 U5940 ( .A1(n4800), .A2(n4803), .ZN(n4418) );
  NAND2_X1 U5941 ( .A1(n9282), .A2(n7987), .ZN(n9262) );
  AND2_X1 U5942 ( .A1(n6980), .A2(n8306), .ZN(n8297) );
  INV_X1 U5943 ( .A(n8297), .ZN(n4749) );
  INV_X1 U5944 ( .A(n8048), .ZN(n9173) );
  AND2_X1 U5945 ( .A1(n7939), .A2(n7904), .ZN(n8048) );
  AND2_X1 U5946 ( .A1(n4699), .A2(n8135), .ZN(n4419) );
  INV_X1 U5947 ( .A(n8290), .ZN(n10256) );
  OAI211_X1 U5948 ( .C1(n6401), .C2(n6476), .A(n5819), .B(n5818), .ZN(n8290)
         );
  XNOR2_X1 U5949 ( .A(n5328), .B(SI_11_), .ZN(n5327) );
  NOR2_X1 U5950 ( .A1(n5717), .A2(n4804), .ZN(n4420) );
  NAND2_X1 U5951 ( .A1(n5597), .A2(n5596), .ZN(n9401) );
  AND2_X1 U5952 ( .A1(n8461), .A2(n6204), .ZN(n4421) );
  AND2_X1 U5953 ( .A1(n7817), .A2(n7933), .ZN(n4422) );
  INV_X1 U5954 ( .A(n9306), .ZN(n4785) );
  INV_X1 U5955 ( .A(n8259), .ZN(n8587) );
  NAND2_X1 U5956 ( .A1(n5531), .A2(n5530), .ZN(n9422) );
  INV_X1 U5957 ( .A(n9422), .ZN(n4710) );
  INV_X1 U5958 ( .A(n7951), .ZN(n5017) );
  NAND2_X1 U5959 ( .A1(n4502), .A2(n5037), .ZN(n4423) );
  AND3_X1 U5960 ( .A1(n5725), .A2(n4960), .A3(n5727), .ZN(n4424) );
  OR2_X1 U5961 ( .A1(n9144), .A2(n9396), .ZN(n4425) );
  AND2_X1 U5962 ( .A1(n4773), .A2(n4772), .ZN(n4426) );
  AND2_X1 U5963 ( .A1(n4780), .A2(n7885), .ZN(n4427) );
  NAND2_X1 U5964 ( .A1(n5448), .A2(n5447), .ZN(n9447) );
  NAND2_X1 U5965 ( .A1(n6082), .A2(n6081), .ZN(n8565) );
  AND3_X1 U5966 ( .A1(n5813), .A2(n5811), .A3(n5812), .ZN(n4428) );
  NAND2_X1 U5967 ( .A1(n6033), .A2(n6032), .ZN(n8809) );
  NOR2_X1 U5968 ( .A1(n6480), .A2(n5200), .ZN(n4429) );
  AND2_X1 U5969 ( .A1(n4701), .A2(n8136), .ZN(n4430) );
  AND2_X1 U5970 ( .A1(n8296), .A2(n8380), .ZN(n4431) );
  AND2_X1 U5971 ( .A1(n4461), .A2(n8562), .ZN(n4432) );
  AND2_X1 U5972 ( .A1(n8112), .A2(n8111), .ZN(n4433) );
  NAND2_X1 U5973 ( .A1(n5499), .A2(n5498), .ZN(n9241) );
  AND2_X1 U5974 ( .A1(n8063), .A2(n8064), .ZN(n4434) );
  NAND2_X1 U5975 ( .A1(n5428), .A2(n5427), .ZN(n9452) );
  INV_X1 U5976 ( .A(n9452), .ZN(n4723) );
  OR2_X1 U5977 ( .A1(n6465), .A2(n6959), .ZN(n4435) );
  NOR2_X1 U5978 ( .A1(n4762), .A2(n7554), .ZN(n4761) );
  NAND2_X1 U5979 ( .A1(n5393), .A2(n5392), .ZN(n9340) );
  AND2_X1 U5980 ( .A1(n8375), .A2(n8562), .ZN(n8573) );
  INV_X1 U5981 ( .A(n8573), .ZN(n4770) );
  INV_X1 U5982 ( .A(n4735), .ZN(n8586) );
  NOR2_X1 U5983 ( .A1(n8600), .A2(n8789), .ZN(n4735) );
  INV_X1 U5984 ( .A(n6259), .ZN(n7800) );
  AND2_X1 U5985 ( .A1(n8364), .A2(n8606), .ZN(n8625) );
  AND2_X1 U5986 ( .A1(n5022), .A2(n5027), .ZN(n4436) );
  NAND2_X1 U5987 ( .A1(n7646), .A2(n7647), .ZN(n4437) );
  OR2_X1 U5988 ( .A1(n6415), .A2(n5771), .ZN(n4438) );
  INV_X1 U5989 ( .A(n8823), .ZN(n8689) );
  NAND2_X1 U5990 ( .A1(n6015), .A2(n6014), .ZN(n8823) );
  AND2_X1 U5991 ( .A1(n4676), .A2(n4675), .ZN(n4439) );
  INV_X1 U5992 ( .A(n9821), .ZN(n9117) );
  NAND2_X1 U5993 ( .A1(n7793), .A2(n7792), .ZN(n9821) );
  AND2_X1 U5994 ( .A1(n5257), .A2(n5066), .ZN(n5260) );
  OR2_X1 U5995 ( .A1(n9422), .A2(n9211), .ZN(n4440) );
  INV_X1 U5996 ( .A(n9261), .ZN(n9271) );
  AND2_X1 U5997 ( .A1(n7959), .A2(n8003), .ZN(n9261) );
  AND2_X1 U5998 ( .A1(n9340), .A2(n9311), .ZN(n4441) );
  AND2_X1 U5999 ( .A1(n7367), .A2(n8461), .ZN(n4442) );
  NOR2_X1 U6000 ( .A1(n4749), .A2(n4748), .ZN(n4443) );
  NOR2_X1 U6001 ( .A1(n8135), .A2(n4700), .ZN(n4444) );
  AND2_X1 U6002 ( .A1(n8268), .A2(n8298), .ZN(n4445) );
  AND2_X1 U6003 ( .A1(n7686), .A2(n7685), .ZN(n4446) );
  NOR2_X1 U6004 ( .A1(n4629), .A2(n4956), .ZN(n4447) );
  AND2_X1 U6005 ( .A1(n8349), .A2(n8638), .ZN(n4448) );
  AND2_X1 U6006 ( .A1(n8844), .A2(n8336), .ZN(n4449) );
  INV_X1 U6007 ( .A(n8408), .ZN(n8307) );
  NAND2_X1 U6008 ( .A1(n8309), .A2(n8300), .ZN(n8408) );
  INV_X1 U6009 ( .A(n4568), .ZN(n4566) );
  NAND2_X1 U6010 ( .A1(n4569), .A2(n8182), .ZN(n4568) );
  AND2_X1 U6011 ( .A1(n4432), .A2(n4766), .ZN(n4765) );
  AND2_X1 U6012 ( .A1(n8245), .A2(n4496), .ZN(n4450) );
  AND2_X1 U6013 ( .A1(n9396), .A2(n9137), .ZN(n4451) );
  NAND2_X1 U6014 ( .A1(n9241), .A2(n9212), .ZN(n4452) );
  AND2_X1 U6015 ( .A1(n5252), .A2(SI_7_), .ZN(n4453) );
  NAND2_X1 U6016 ( .A1(n8127), .A2(n8126), .ZN(n4454) );
  AND2_X1 U6017 ( .A1(n8835), .A2(n7581), .ZN(n4455) );
  INV_X1 U6018 ( .A(n4782), .ZN(n4781) );
  NAND2_X1 U6019 ( .A1(n9442), .A2(n9284), .ZN(n4782) );
  NOR2_X1 U6020 ( .A1(n8771), .A2(n8564), .ZN(n4456) );
  NOR2_X1 U6021 ( .A1(n8804), .A2(n8659), .ZN(n4457) );
  INV_X1 U6022 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5994) );
  INV_X1 U6023 ( .A(n8305), .ZN(n4541) );
  INV_X1 U6024 ( .A(n8313), .ZN(n4542) );
  INV_X1 U6025 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5735) );
  INV_X1 U6026 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5117) );
  AND2_X1 U6027 ( .A1(n8360), .A2(n8356), .ZN(n4458) );
  INV_X1 U6028 ( .A(n4691), .ZN(n4690) );
  NOR2_X1 U6029 ( .A1(n8215), .A2(n4692), .ZN(n4691) );
  AND2_X1 U6030 ( .A1(n8124), .A2(n8123), .ZN(n4459) );
  AND2_X1 U6031 ( .A1(n5192), .A2(SI_3_), .ZN(n4460) );
  OAI21_X1 U6032 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5290) );
  AND2_X1 U6033 ( .A1(n8377), .A2(n8376), .ZN(n4461) );
  OAI21_X1 U6034 ( .B1(n4689), .B2(n4688), .A(n4454), .ZN(n4687) );
  NAND2_X1 U6035 ( .A1(n4886), .A2(n4884), .ZN(n5605) );
  OR2_X1 U6036 ( .A1(n4561), .A2(n8259), .ZN(n4462) );
  OR2_X1 U6037 ( .A1(n8814), .A2(n8684), .ZN(n8356) );
  NAND2_X1 U6038 ( .A1(n8426), .A2(n8378), .ZN(n4463) );
  INV_X1 U6039 ( .A(n4645), .ZN(n4644) );
  NAND2_X1 U6040 ( .A1(n7621), .A2(n7467), .ZN(n4645) );
  AND2_X1 U6041 ( .A1(n6688), .A2(n6591), .ZN(n4464) );
  OR2_X1 U6042 ( .A1(n8702), .A2(n6138), .ZN(n4773) );
  AND2_X1 U6043 ( .A1(n5029), .A2(n5028), .ZN(n4465) );
  OR2_X1 U6044 ( .A1(n4710), .A2(n9187), .ZN(n4466) );
  AND2_X1 U6045 ( .A1(n4808), .A2(n5129), .ZN(n4467) );
  AND2_X1 U6046 ( .A1(n4541), .A2(n8300), .ZN(n4468) );
  OR2_X1 U6047 ( .A1(n4648), .A2(n8901), .ZN(n4469) );
  AND2_X1 U6048 ( .A1(n4955), .A2(n4953), .ZN(n4470) );
  AOI21_X1 U6049 ( .B1(n4761), .B2(n4759), .A(n4449), .ZN(n4758) );
  INV_X1 U6050 ( .A(n8312), .ZN(n4611) );
  OR2_X1 U6051 ( .A1(n7264), .A2(n7231), .ZN(n8312) );
  AND2_X1 U6052 ( .A1(n4542), .A2(n4539), .ZN(n4471) );
  INV_X1 U6053 ( .A(n9419), .ZN(n5716) );
  AND2_X1 U6054 ( .A1(n5064), .A2(n4941), .ZN(n4472) );
  INV_X1 U6055 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U6056 ( .A1(n8316), .A2(n8315), .ZN(n4473) );
  NAND2_X1 U6057 ( .A1(n9860), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4474) );
  INV_X1 U6058 ( .A(n4996), .ZN(n4995) );
  NAND2_X1 U6059 ( .A1(n4998), .A2(n8424), .ZN(n4996) );
  INV_X1 U6060 ( .A(n6128), .ZN(n8432) );
  NAND2_X1 U6061 ( .A1(n8948), .A2(n7657), .ZN(n4636) );
  INV_X1 U6062 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n4666) );
  OR2_X1 U6063 ( .A1(n5524), .A2(n4903), .ZN(n4475) );
  OR2_X1 U6064 ( .A1(n6607), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4476) );
  AND2_X1 U6065 ( .A1(n4502), .A2(n5079), .ZN(n5357) );
  AND2_X1 U6066 ( .A1(n9924), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4477) );
  AND4_X1 U6067 ( .A1(n5828), .A2(n4821), .A3(n4818), .A4(n4817), .ZN(n4478)
         );
  NAND2_X1 U6068 ( .A1(n6073), .A2(n6072), .ZN(n8783) );
  INV_X1 U6069 ( .A(n8783), .ZN(n4991) );
  NAND2_X1 U6070 ( .A1(n5611), .A2(n5610), .ZN(n9396) );
  INV_X1 U6071 ( .A(n9396), .ZN(n4719) );
  INV_X1 U6072 ( .A(n9027), .ZN(n9123) );
  NAND2_X1 U6073 ( .A1(n9252), .A2(n4400), .ZN(n4712) );
  NAND2_X1 U6074 ( .A1(n4948), .A2(n4945), .ZN(n8968) );
  AND2_X1 U6075 ( .A1(n9295), .A2(n5436), .ZN(n4479) );
  AND2_X1 U6076 ( .A1(n7712), .A2(n7713), .ZN(n4480) );
  NAND2_X1 U6077 ( .A1(n8695), .A2(n4742), .ZN(n4743) );
  NAND2_X1 U6078 ( .A1(n9346), .A2(n4722), .ZN(n4725) );
  OR2_X1 U6079 ( .A1(n6655), .A2(n6990), .ZN(n4481) );
  NAND2_X1 U6080 ( .A1(n8347), .A2(n8346), .ZN(n4482) );
  AND2_X1 U6081 ( .A1(n8185), .A2(n8186), .ZN(n4483) );
  NAND2_X1 U6082 ( .A1(n7675), .A2(n7676), .ZN(n4484) );
  AND2_X1 U6083 ( .A1(n8329), .A2(n8330), .ZN(n8328) );
  OR2_X1 U6084 ( .A1(n8230), .A2(n8128), .ZN(n4580) );
  AND2_X1 U6085 ( .A1(n5460), .A2(SI_18_), .ZN(n4485) );
  NAND2_X1 U6086 ( .A1(n5828), .A2(n5725), .ZN(n5843) );
  NAND2_X1 U6087 ( .A1(n7395), .A2(n8991), .ZN(n4486) );
  AND2_X1 U6088 ( .A1(n9390), .A2(n9111), .ZN(n8052) );
  AND2_X1 U6089 ( .A1(n6684), .A2(n6683), .ZN(n4487) );
  AND2_X1 U6090 ( .A1(n6819), .A2(n4825), .ZN(n4488) );
  OR2_X1 U6091 ( .A1(n7006), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4489) );
  AND2_X1 U6092 ( .A1(n7468), .A2(n7467), .ZN(n7622) );
  NAND2_X1 U6093 ( .A1(n6040), .A2(n6039), .ZN(n8804) );
  INV_X1 U6094 ( .A(n8804), .ZN(n4739) );
  NAND2_X1 U6095 ( .A1(n6698), .A2(n7089), .ZN(n6699) );
  NAND2_X1 U6096 ( .A1(n5698), .A2(n5697), .ZN(n7204) );
  AND2_X1 U6097 ( .A1(n6981), .A2(n8299), .ZN(n4490) );
  INV_X1 U6098 ( .A(n4790), .ZN(n4789) );
  NOR2_X1 U6099 ( .A1(n9331), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U6100 ( .A1(n6160), .A2(n6161), .ZN(n6169) );
  INV_X1 U6101 ( .A(n4894), .ZN(n4893) );
  NOR2_X1 U6102 ( .A1(n5571), .A2(n4895), .ZN(n4894) );
  AND2_X1 U6103 ( .A1(n5626), .A2(n5625), .ZN(n4491) );
  INV_X1 U6104 ( .A(n4876), .ZN(n4875) );
  AND3_X1 U6105 ( .A1(n8280), .A2(n8278), .A3(n8276), .ZN(n4492) );
  INV_X1 U6106 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6159) );
  NOR2_X1 U6107 ( .A1(n4871), .A2(n7594), .ZN(n4870) );
  INV_X1 U6108 ( .A(n10211), .ZN(n10190) );
  NAND2_X1 U6109 ( .A1(n5283), .A2(n5282), .ZN(n7195) );
  INV_X1 U6110 ( .A(n7195), .ZN(n4707) );
  CLKBUF_X1 U6111 ( .A(n6492), .Z(n9039) );
  XNOR2_X1 U6112 ( .A(n6164), .B(n6163), .ZN(n8257) );
  NOR2_X2 U6113 ( .A1(n8686), .A2(n10293), .ZN(n8848) );
  INV_X1 U6114 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5010) );
  NAND2_X1 U6115 ( .A1(n5891), .A2(n5890), .ZN(n7421) );
  INV_X1 U6116 ( .A(n7421), .ZN(n4736) );
  AND2_X1 U6117 ( .A1(n10138), .A2(n6199), .ZN(n4493) );
  INV_X1 U6118 ( .A(n6331), .ZN(n4667) );
  INV_X1 U6119 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4509) );
  AND2_X1 U6120 ( .A1(n6011), .A2(n6120), .ZN(n8680) );
  INV_X1 U6121 ( .A(n8680), .ZN(n8730) );
  INV_X1 U6122 ( .A(n5121), .ZN(n7596) );
  NOR2_X1 U6123 ( .A1(n9850), .A2(n9871), .ZN(n9849) );
  INV_X1 U6124 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4511) );
  INV_X1 U6125 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4592) );
  INV_X1 U6126 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U6127 ( .A1(n4522), .A2(n8393), .ZN(n4521) );
  BUF_X2 U6128 ( .A(n5143), .Z(n6190) );
  NOR2_X1 U6129 ( .A1(n5690), .A2(n8069), .ZN(n5011) );
  NAND2_X1 U6130 ( .A1(n9476), .A2(n4387), .ZN(n4499) );
  NAND2_X1 U6131 ( .A1(n9394), .A2(n4500), .ZN(n9476) );
  NAND2_X1 U6132 ( .A1(n8486), .A2(n8485), .ZN(n8484) );
  NAND2_X1 U6133 ( .A1(n4731), .A2(n4730), .ZN(P2_U3549) );
  NAND2_X1 U6134 ( .A1(n9805), .A2(n9806), .ZN(n9804) );
  OR2_X1 U6135 ( .A1(n6141), .A2(n8385), .ZN(n4496) );
  NAND2_X1 U6136 ( .A1(n6141), .A2(n8385), .ZN(n8245) );
  NAND2_X1 U6137 ( .A1(n4746), .A2(n4607), .ZN(n6136) );
  NAND2_X1 U6138 ( .A1(n10008), .A2(n10014), .ZN(n10007) );
  NAND2_X1 U6139 ( .A1(n7209), .A2(n7973), .ZN(n7268) );
  NAND2_X1 U6140 ( .A1(n4651), .A2(n9192), .ZN(n4650) );
  NAND2_X1 U6141 ( .A1(n4928), .A2(n8021), .ZN(n4927) );
  XNOR2_X1 U6142 ( .A(n5214), .B(n5213), .ZN(n6266) );
  NAND2_X1 U6143 ( .A1(n4923), .A2(n4922), .ZN(n4921) );
  NAND2_X1 U6144 ( .A1(n4921), .A2(n4920), .ZN(n8105) );
  NAND4_X1 U6145 ( .A1(n7916), .A2(n7915), .A3(n9136), .A4(n7917), .ZN(n4503)
         );
  NAND4_X1 U6146 ( .A1(n4942), .A2(n5062), .A3(n5064), .A4(n5063), .ZN(n5220)
         );
  NAND2_X1 U6147 ( .A1(n7205), .A2(n5699), .ZN(n7267) );
  NAND2_X1 U6148 ( .A1(n5685), .A2(n5684), .ZN(n6921) );
  NAND2_X2 U6149 ( .A1(n5709), .A2(n5708), .ZN(n9344) );
  OAI21_X1 U6150 ( .B1(n6784), .B2(n7820), .A(n5693), .ZN(n6811) );
  NAND2_X1 U6151 ( .A1(n9197), .A2(n4440), .ZN(n4797) );
  NAND2_X1 U6152 ( .A1(n4797), .A2(n4466), .ZN(n9182) );
  NAND2_X1 U6153 ( .A1(n5698), .A2(n4805), .ZN(n7205) );
  INV_X1 U6154 ( .A(n5189), .ZN(n4514) );
  NAND2_X1 U6155 ( .A1(n5206), .A2(n5205), .ZN(n5210) );
  NAND2_X1 U6156 ( .A1(n8327), .A2(n8380), .ZN(n4526) );
  NAND2_X1 U6157 ( .A1(n8326), .A2(n8393), .ZN(n4525) );
  NAND2_X1 U6158 ( .A1(n4524), .A2(n4528), .ZN(n8343) );
  NAND3_X1 U6159 ( .A1(n4526), .A2(n4525), .A3(n4527), .ZN(n4524) );
  OR2_X1 U6160 ( .A1(n8311), .A2(n4538), .ZN(n4537) );
  OR2_X1 U6161 ( .A1(n8301), .A2(n4540), .ZN(n4536) );
  NAND3_X1 U6162 ( .A1(n4537), .A2(n4536), .A3(n4409), .ZN(n8325) );
  AND2_X1 U6163 ( .A1(n8310), .A2(n8309), .ZN(n4539) );
  NAND2_X1 U6164 ( .A1(n8354), .A2(n4546), .ZN(n4543) );
  NAND2_X1 U6165 ( .A1(n4543), .A2(n4544), .ZN(n8351) );
  NAND2_X1 U6166 ( .A1(n4552), .A2(n4553), .ZN(n8384) );
  NAND2_X1 U6167 ( .A1(n8370), .A2(n4554), .ZN(n4552) );
  NAND2_X1 U6168 ( .A1(n5171), .A2(n5170), .ZN(n4562) );
  NAND3_X1 U6169 ( .A1(n4575), .A2(n4412), .A3(n4574), .ZN(n8156) );
  NAND4_X1 U6170 ( .A1(n4575), .A2(n4412), .A3(n4578), .A4(n4574), .ZN(n4698)
         );
  INV_X1 U6171 ( .A(n8133), .ZN(n4579) );
  NOR2_X1 U6172 ( .A1(n8133), .A2(n4577), .ZN(n4576) );
  INV_X1 U6173 ( .A(n8134), .ZN(n4577) );
  AOI21_X2 U6174 ( .B1(n8167), .B2(n4399), .A(n4687), .ZN(n8129) );
  AOI21_X2 U6175 ( .B1(n8207), .B2(n8206), .A(n4430), .ZN(n8198) );
  AND2_X1 U6176 ( .A1(n6160), .A2(n5006), .ZN(n5751) );
  NAND2_X1 U6177 ( .A1(n4593), .A2(n6160), .ZN(n8878) );
  NAND3_X1 U6178 ( .A1(n4593), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6160), .ZN(
        n4589) );
  OAI21_X2 U6179 ( .B1(n4602), .B2(n4407), .A(n4597), .ZN(n8636) );
  NAND2_X1 U6180 ( .A1(n7181), .A2(n8312), .ZN(n4608) );
  NAND2_X1 U6181 ( .A1(n4608), .A2(n4609), .ZN(n6137) );
  INV_X1 U6182 ( .A(n10187), .ZN(n10195) );
  NAND2_X1 U6183 ( .A1(n4618), .A2(n4615), .ZN(P2_U3267) );
  NAND2_X1 U6184 ( .A1(n6149), .A2(n10222), .ZN(n4618) );
  NAND3_X1 U6185 ( .A1(n4939), .A2(n4437), .A3(n9013), .ZN(n8937) );
  NAND2_X1 U6186 ( .A1(n4619), .A2(n7640), .ZN(n9013) );
  NAND2_X1 U6187 ( .A1(n4620), .A2(n8890), .ZN(n4619) );
  NAND2_X1 U6188 ( .A1(n8891), .A2(n8893), .ZN(n4620) );
  NAND2_X1 U6189 ( .A1(n6698), .A2(n4414), .ZN(n6878) );
  NAND2_X1 U6190 ( .A1(n6878), .A2(n6877), .ZN(n6884) );
  NOR2_X1 U6191 ( .A1(n4470), .A2(n4625), .ZN(n7736) );
  NAND2_X1 U6192 ( .A1(n4626), .A2(n4627), .ZN(n4625) );
  OR2_X1 U6193 ( .A1(n8930), .A2(n4628), .ZN(n4626) );
  OR2_X1 U6194 ( .A1(n8930), .A2(n8931), .ZN(n4955) );
  NAND2_X1 U6195 ( .A1(n8948), .A2(n4632), .ZN(n4631) );
  NAND2_X1 U6196 ( .A1(n4948), .A2(n4639), .ZN(n4637) );
  NAND2_X1 U6197 ( .A1(n4637), .A2(n4638), .ZN(n7691) );
  NAND2_X1 U6198 ( .A1(n4643), .A2(n4644), .ZN(n4642) );
  NAND2_X1 U6199 ( .A1(n4646), .A2(n4469), .ZN(n8900) );
  NAND3_X1 U6200 ( .A1(n7695), .A2(n4647), .A3(n8979), .ZN(n4646) );
  NOR2_X2 U6201 ( .A1(n8900), .A2(n8904), .ZN(n8961) );
  INV_X1 U6202 ( .A(n7701), .ZN(n4648) );
  NAND3_X1 U6203 ( .A1(n4654), .A2(n4652), .A3(n4650), .ZN(P1_U3260) );
  INV_X1 U6204 ( .A(n4657), .ZN(n4658) );
  OAI21_X1 U6205 ( .B1(n9865), .B2(n6245), .A(n4474), .ZN(n4657) );
  OAI21_X1 U6206 ( .B1(n6244), .B2(n9865), .A(n4658), .ZN(n4661) );
  INV_X1 U6207 ( .A(n4661), .ZN(n6250) );
  INV_X1 U6208 ( .A(n6249), .ZN(n4660) );
  XNOR2_X1 U6209 ( .A(n9055), .B(n9063), .ZN(n9044) );
  MUX2_X1 U6210 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6243), .S(n9856), .Z(n9850)
         );
  OR2_X1 U6211 ( .A1(n7302), .A2(n7303), .ZN(n7447) );
  NAND2_X1 U6212 ( .A1(n7302), .A2(n4684), .ZN(n4681) );
  NAND2_X1 U6213 ( .A1(n4698), .A2(n4702), .ZN(n4701) );
  XNOR2_X1 U6214 ( .A(n4701), .B(n8135), .ZN(n8207) );
  NAND3_X1 U6215 ( .A1(n4706), .A2(n4841), .A3(n10141), .ZN(n4705) );
  INV_X1 U6216 ( .A(n4712), .ZN(n9198) );
  NAND2_X1 U6217 ( .A1(n9155), .A2(n9150), .ZN(n9144) );
  NAND2_X1 U6218 ( .A1(n9155), .A2(n4714), .ZN(n9115) );
  AND2_X1 U6219 ( .A1(n9155), .A2(n4713), .ZN(n9116) );
  INV_X1 U6220 ( .A(n4725), .ZN(n9291) );
  OAI21_X2 U6221 ( .B1(n6190), .B2(n9856), .A(n4726), .ZN(n6747) );
  NAND2_X2 U6222 ( .A1(n5640), .A2(n5641), .ZN(n5143) );
  NAND2_X2 U6223 ( .A1(n5143), .A2(n7800), .ZN(n7806) );
  NOR2_X2 U6224 ( .A1(n8754), .A2(n8831), .ZN(n8694) );
  XNOR2_X2 U6225 ( .A(n4728), .B(n5748), .ZN(n6417) );
  AND2_X2 U6226 ( .A1(n5760), .A2(n5734), .ZN(n6160) );
  NOR2_X2 U6227 ( .A1(n8576), .A2(n8777), .ZN(n8558) );
  NOR2_X2 U6228 ( .A1(n7188), .A2(n7264), .ZN(n7189) );
  NOR2_X2 U6229 ( .A1(n6717), .A2(n6992), .ZN(n4737) );
  NOR2_X2 U6230 ( .A1(n6947), .A2(n6192), .ZN(n6969) );
  INV_X1 U6231 ( .A(n4743), .ZN(n8665) );
  AOI21_X1 U6232 ( .B1(n8299), .B2(n4749), .A(n4748), .ZN(n4744) );
  INV_X1 U6233 ( .A(n8299), .ZN(n4745) );
  INV_X1 U6234 ( .A(n4747), .ZN(n4746) );
  OAI21_X1 U6235 ( .B1(n8299), .B2(n4748), .A(n8410), .ZN(n4747) );
  NAND2_X1 U6236 ( .A1(n4754), .A2(n8278), .ZN(n4753) );
  NAND2_X1 U6237 ( .A1(n4757), .A2(n8272), .ZN(n4754) );
  NAND2_X1 U6238 ( .A1(n4756), .A2(n8278), .ZN(n10188) );
  NAND2_X1 U6239 ( .A1(n8272), .A2(n4492), .ZN(n4756) );
  NAND2_X1 U6240 ( .A1(n8280), .A2(n8278), .ZN(n8402) );
  NAND2_X1 U6241 ( .A1(n6160), .A2(n5007), .ZN(n5736) );
  NAND2_X1 U6242 ( .A1(n6131), .A2(n6130), .ZN(n10176) );
  AOI21_X1 U6243 ( .B1(n7604), .B2(n8426), .A(n6140), .ZN(n6141) );
  OAI21_X2 U6244 ( .B1(n7313), .B2(n8323), .A(n8322), .ZN(n7492) );
  NAND2_X1 U6245 ( .A1(n8277), .A2(n10207), .ZN(n8272) );
  NAND2_X1 U6246 ( .A1(n6137), .A2(n8317), .ZN(n7313) );
  OR2_X1 U6247 ( .A1(n5845), .A2(n6269), .ZN(n5779) );
  OR2_X1 U6248 ( .A1(n5845), .A2(n6261), .ZN(n5804) );
  NAND2_X4 U6249 ( .A1(n6417), .A2(n7589), .ZN(n6401) );
  NAND2_X1 U6250 ( .A1(n5806), .A2(n10251), .ZN(n8280) );
  AOI21_X2 U6251 ( .B1(n9272), .B2(n4427), .A(n4776), .ZN(n9215) );
  CLKBUF_X1 U6252 ( .A(n9272), .Z(n4774) );
  OAI21_X2 U6253 ( .B1(n9344), .B2(n4786), .A(n4784), .ZN(n9304) );
  OR2_X1 U6254 ( .A1(n5717), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U6255 ( .A1(n5717), .A2(n4396), .ZN(n4799) );
  AND2_X1 U6256 ( .A1(n9408), .A2(n9143), .ZN(n4804) );
  NAND3_X1 U6257 ( .A1(n5037), .A2(n5336), .A3(n4808), .ZN(n5114) );
  AND3_X2 U6258 ( .A1(n5037), .A2(n5336), .A3(n4467), .ZN(n5126) );
  NAND3_X1 U6259 ( .A1(n5037), .A2(n4502), .A3(n5091), .ZN(n5089) );
  NAND2_X1 U6260 ( .A1(n4809), .A2(n5680), .ZN(n6737) );
  NAND2_X1 U6261 ( .A1(n4809), .A2(n8062), .ZN(n8065) );
  AND2_X1 U6262 ( .A1(n8060), .A2(n4809), .ZN(n10008) );
  INV_X1 U6263 ( .A(n8257), .ZN(n4811) );
  NAND2_X1 U6264 ( .A1(n5760), .A2(n4812), .ZN(n5993) );
  NAND2_X1 U6265 ( .A1(n4813), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5762) );
  INV_X1 U6266 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n4820) );
  INV_X1 U6267 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n4819) );
  AND2_X2 U6268 ( .A1(n4814), .A2(n5044), .ZN(n5760) );
  NAND3_X1 U6269 ( .A1(n6860), .A2(n4842), .A3(n6213), .ZN(n6766) );
  NAND2_X1 U6270 ( .A1(n4844), .A2(n4845), .ZN(n6207) );
  INV_X1 U6271 ( .A(n6912), .ZN(n4846) );
  INV_X1 U6272 ( .A(n6202), .ZN(n4847) );
  NAND2_X1 U6273 ( .A1(n7565), .A2(n4851), .ZN(n4848) );
  NAND2_X1 U6274 ( .A1(n5995), .A2(n5994), .ZN(n6123) );
  NAND2_X1 U6275 ( .A1(n5995), .A2(n4857), .ZN(n6127) );
  NAND2_X1 U6276 ( .A1(n8026), .A2(n9111), .ZN(n4858) );
  INV_X1 U6277 ( .A(n7928), .ZN(n4859) );
  NAND2_X1 U6278 ( .A1(n5423), .A2(n4863), .ZN(n4861) );
  NAND2_X1 U6279 ( .A1(n5609), .A2(n4870), .ZN(n4868) );
  OAI21_X1 U6280 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5624) );
  AOI21_X1 U6281 ( .B1(n5608), .B2(n5607), .A(n4877), .ZN(n4876) );
  NAND2_X1 U6282 ( .A1(n5242), .A2(n4881), .ZN(n4879) );
  NAND2_X1 U6283 ( .A1(n5242), .A2(n5241), .ZN(n4880) );
  INV_X1 U6284 ( .A(n5244), .ZN(n4883) );
  NAND2_X1 U6285 ( .A1(n5554), .A2(n4888), .ZN(n4886) );
  NAND2_X1 U6286 ( .A1(n5497), .A2(n4901), .ZN(n4900) );
  NAND2_X1 U6287 ( .A1(n5331), .A2(n4917), .ZN(n4910) );
  OAI21_X1 U6288 ( .B1(n5331), .B2(n4919), .A(n5330), .ZN(n5351) );
  NAND3_X1 U6289 ( .A1(n8059), .A2(n8053), .A3(n4924), .ZN(n4923) );
  NAND2_X1 U6290 ( .A1(n6393), .A2(n4934), .ZN(n4933) );
  NAND2_X1 U6291 ( .A1(n6391), .A2(n6392), .ZN(n4934) );
  NAND2_X1 U6292 ( .A1(n4933), .A2(n4932), .ZN(n6500) );
  OR2_X1 U6293 ( .A1(n4934), .A2(n7770), .ZN(n4932) );
  OAI21_X1 U6294 ( .B1(n6393), .B2(n4934), .A(n4933), .ZN(n9870) );
  NAND2_X1 U6295 ( .A1(n6590), .A2(n4464), .ZN(n4937) );
  NAND2_X1 U6296 ( .A1(n4937), .A2(n4935), .ZN(n6698) );
  NAND3_X1 U6297 ( .A1(n5063), .A2(n5062), .A3(n5064), .ZN(n5187) );
  OAI21_X1 U6298 ( .B1(n8930), .B2(n4952), .A(n4951), .ZN(n7776) );
  OR2_X1 U6299 ( .A1(n8931), .A2(n4480), .ZN(n4952) );
  NAND2_X1 U6300 ( .A1(n5257), .A2(n4957), .ZN(n5107) );
  NAND2_X1 U6301 ( .A1(n5915), .A2(n4964), .ZN(n4962) );
  NAND2_X1 U6302 ( .A1(n4962), .A2(n4963), .ZN(n7311) );
  NAND2_X1 U6303 ( .A1(n4969), .A2(n4967), .ZN(n6985) );
  NAND2_X1 U6304 ( .A1(n5859), .A2(n5858), .ZN(n6712) );
  INV_X1 U6305 ( .A(n5858), .ZN(n4972) );
  NAND2_X1 U6306 ( .A1(n4973), .A2(n4976), .ZN(n6119) );
  NAND2_X1 U6307 ( .A1(n8583), .A2(n4978), .ZN(n4973) );
  AND2_X2 U6308 ( .A1(n4975), .A2(n4393), .ZN(n8570) );
  OR2_X1 U6309 ( .A1(n8648), .A2(n4996), .ZN(n4992) );
  AND2_X2 U6310 ( .A1(n4992), .A2(n4993), .ZN(n8597) );
  NAND2_X1 U6311 ( .A1(n8738), .A2(n4395), .ZN(n5002) );
  INV_X1 U6312 ( .A(n5005), .ZN(n8740) );
  XNOR2_X1 U6313 ( .A(n5012), .B(n7109), .ZN(n7099) );
  NAND2_X1 U6314 ( .A1(n9262), .A2(n5019), .ZN(n5015) );
  NAND2_X1 U6315 ( .A1(n5015), .A2(n5016), .ZN(n9225) );
  NAND2_X1 U6316 ( .A1(n9202), .A2(n5026), .ZN(n5025) );
  NAND2_X1 U6317 ( .A1(n5126), .A2(n5127), .ZN(n5116) );
  NAND2_X1 U6318 ( .A1(n5126), .A2(n5030), .ZN(n9772) );
  AND2_X1 U6319 ( .A1(n10007), .A2(n8064), .ZN(n7944) );
  AND2_X2 U6320 ( .A1(n8064), .A2(n8062), .ZN(n10014) );
  INV_X1 U6321 ( .A(n5806), .ZN(n5805) );
  OR2_X1 U6322 ( .A1(n8770), .A2(n8848), .ZN(n8776) );
  OAI211_X1 U6323 ( .C1(n5134), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5133), .ZN(n5156) );
  INV_X1 U6324 ( .A(n5721), .ZN(n5722) );
  NAND2_X1 U6325 ( .A1(n7937), .A2(n7935), .ZN(n8059) );
  XNOR2_X1 U6326 ( .A(n5103), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5719) );
  INV_X1 U6327 ( .A(n5753), .ZN(n8881) );
  NAND2_X1 U6328 ( .A1(n5752), .A2(n5753), .ZN(n5791) );
  INV_X1 U6329 ( .A(n8129), .ZN(n8132) );
  INV_X1 U6330 ( .A(n7691), .ZN(n7694) );
  XNOR2_X1 U6331 ( .A(n8783), .B(n8138), .ZN(n8144) );
  NAND2_X1 U6332 ( .A1(n5100), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5110) );
  OAI21_X1 U6333 ( .B1(n5100), .B2(n5073), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5096) );
  OR2_X1 U6334 ( .A1(n5485), .A2(n10128), .ZN(n5147) );
  OR2_X1 U6335 ( .A1(n5485), .A2(n6389), .ZN(n5140) );
  OR2_X1 U6336 ( .A1(n5485), .A2(n6235), .ZN(n5125) );
  AOI21_X2 U6337 ( .B1(n8664), .B2(n8671), .A(n6031), .ZN(n8648) );
  AND2_X1 U6338 ( .A1(n5313), .A2(n5298), .ZN(n5039) );
  AND2_X1 U6339 ( .A1(n7401), .A2(n7400), .ZN(n5042) );
  AND2_X1 U6340 ( .A1(n5094), .A2(n5093), .ZN(n5043) );
  INV_X1 U6341 ( .A(n8411), .ZN(n5914) );
  AND2_X1 U6342 ( .A1(n5422), .A2(n5407), .ZN(n5045) );
  AND2_X1 U6343 ( .A1(n5291), .A2(n5279), .ZN(n5046) );
  AND2_X1 U6344 ( .A1(n5368), .A2(n5356), .ZN(n5047) );
  NOR2_X1 U6345 ( .A1(n7399), .A2(n8992), .ZN(n5048) );
  INV_X1 U6346 ( .A(n10021), .ZN(n9321) );
  INV_X1 U6347 ( .A(n8456), .ZN(n8608) );
  NOR2_X1 U6348 ( .A1(n7293), .A2(n7292), .ZN(n5049) );
  NOR2_X1 U6349 ( .A1(n7925), .A2(n7924), .ZN(n7926) );
  INV_X1 U6350 ( .A(n8428), .ZN(n8385) );
  INV_X1 U6351 ( .A(n7385), .ZN(n7386) );
  INV_X1 U6352 ( .A(n8130), .ZN(n8131) );
  INV_X1 U6353 ( .A(n6041), .ZN(n5746) );
  NOR2_X1 U6354 ( .A1(n5881), .A2(n6509), .ZN(n5880) );
  INV_X1 U6355 ( .A(n6065), .ZN(n6063) );
  INV_X1 U6356 ( .A(n5993), .ZN(n5995) );
  OR2_X1 U6357 ( .A1(n6493), .A2(n6732), .ZN(n6501) );
  INV_X1 U6358 ( .A(n5532), .ZN(n5060) );
  INV_X1 U6359 ( .A(n5305), .ZN(n5054) );
  INV_X1 U6360 ( .A(n5580), .ZN(n5061) );
  INV_X1 U6361 ( .A(n5457), .ZN(n5458) );
  INV_X1 U6362 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5314) );
  INV_X1 U6363 ( .A(n5249), .ZN(n5250) );
  NOR2_X1 U6364 ( .A1(n8132), .A2(n8131), .ZN(n8133) );
  AND3_X1 U6365 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n5834) );
  INV_X1 U6366 ( .A(n8166), .ZN(n8118) );
  NAND2_X1 U6367 ( .A1(n5787), .A2(n6204), .ZN(n6198) );
  OR2_X1 U6368 ( .A1(n6086), .A2(n6085), .ZN(n6100) );
  OR2_X1 U6369 ( .A1(n6043), .A2(n9715), .ZN(n6052) );
  OR2_X1 U6370 ( .A1(n6000), .A2(n8536), .ZN(n6027) );
  NAND2_X1 U6371 ( .A1(n5851), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5881) );
  INV_X1 U6372 ( .A(n6401), .ZN(n6012) );
  NAND2_X1 U6373 ( .A1(n7606), .A2(n7605), .ZN(n7607) );
  AOI21_X1 U6374 ( .B1(n6007), .B2(n9648), .A(n6159), .ZN(n6008) );
  INV_X1 U6375 ( .A(n7631), .ZN(n7632) );
  INV_X1 U6376 ( .A(n7692), .ZN(n7693) );
  INV_X1 U6377 ( .A(n7663), .ZN(n7664) );
  OR3_X1 U6378 ( .A1(n5563), .A2(n5562), .A3(n5561), .ZN(n5580) );
  NAND2_X1 U6379 ( .A1(n5057), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6380 ( .A1(n5052), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5305) );
  NAND2_X1 U6381 ( .A1(n5061), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5614) );
  INV_X1 U6382 ( .A(n9310), .ZN(n5711) );
  OR2_X1 U6383 ( .A1(n5321), .A2(n9622), .ZN(n5341) );
  OR2_X1 U6384 ( .A1(n10036), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5678) );
  INV_X1 U6385 ( .A(n5606), .ZN(n5608) );
  NAND2_X1 U6386 ( .A1(n5384), .A2(n5383), .ZN(n5402) );
  INV_X1 U6387 ( .A(n8565), .ZN(n8151) );
  AND2_X1 U6388 ( .A1(n6100), .A2(n6087), .ZN(n8559) );
  INV_X1 U6389 ( .A(n5791), .ZN(n6088) );
  INV_X1 U6390 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n6509) );
  INV_X1 U6391 ( .A(n10179), .ZN(n6130) );
  AND2_X1 U6392 ( .A1(n8333), .A2(n8332), .ZN(n8419) );
  AND2_X1 U6393 ( .A1(n8318), .A2(n8322), .ZN(n7312) );
  AND2_X1 U6394 ( .A1(n7545), .A2(n6168), .ZN(n6171) );
  INV_X1 U6395 ( .A(n9137), .ZN(n7727) );
  XNOR2_X1 U6396 ( .A(n7164), .B(n7716), .ZN(n7387) );
  AND2_X1 U6397 ( .A1(n7782), .A2(n8951), .ZN(n7777) );
  XNOR2_X1 U6398 ( .A(n7617), .B(n7716), .ZN(n7712) );
  AND2_X1 U6399 ( .A1(n6547), .A2(n6566), .ZN(n6553) );
  INV_X1 U6400 ( .A(n9007), .ZN(n9017) );
  XNOR2_X1 U6401 ( .A(n5130), .B(n5129), .ZN(n5641) );
  AND2_X1 U6402 ( .A1(n5615), .A2(n5655), .ZN(n9130) );
  OR2_X1 U6403 ( .A1(n5518), .A2(n8982), .ZN(n5532) );
  OR2_X1 U6404 ( .A1(n5179), .A2(n6243), .ZN(n5123) );
  INV_X1 U6405 ( .A(n9401), .ZN(n9150) );
  INV_X1 U6406 ( .A(n8092), .ZN(n9192) );
  NAND2_X1 U6407 ( .A1(n8020), .A2(n8088), .ZN(n8050) );
  INV_X1 U6408 ( .A(n10118), .ZN(n9469) );
  INV_X1 U6409 ( .A(n6747), .ZN(n10074) );
  AND2_X1 U6410 ( .A1(n6221), .A2(n6150), .ZN(n8851) );
  INV_X1 U6411 ( .A(n10143), .ZN(n8228) );
  INV_X1 U6412 ( .A(n6414), .ZN(n9803) );
  AND2_X1 U6413 ( .A1(n6408), .A2(n7589), .ZN(n10168) );
  NAND2_X1 U6414 ( .A1(n8356), .A2(n8357), .ZN(n8671) );
  INV_X1 U6415 ( .A(n10210), .ZN(n10189) );
  INV_X1 U6416 ( .A(n10219), .ZN(n8711) );
  AND2_X1 U6417 ( .A1(n8774), .A2(n8773), .ZN(n8775) );
  INV_X1 U6418 ( .A(n8851), .ZN(n10296) );
  AND2_X1 U6419 ( .A1(n6129), .A2(n6128), .ZN(n10293) );
  INV_X1 U6420 ( .A(n8848), .ZN(n10302) );
  NOR2_X1 U6421 ( .A1(n6171), .A2(n7574), .ZN(n10225) );
  INV_X1 U6422 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6161) );
  AND2_X1 U6423 ( .A1(n6709), .A2(n9822), .ZN(n9023) );
  NAND4_X2 U6424 ( .A1(n5148), .A2(n5147), .A3(n5146), .A4(n5145), .ZN(n6542)
         );
  AND2_X1 U6425 ( .A1(n9105), .A2(n9874), .ZN(n9950) );
  AND2_X1 U6426 ( .A1(n7960), .A2(n7951), .ZN(n9245) );
  INV_X1 U6427 ( .A(n8043), .ZN(n9283) );
  INV_X1 U6428 ( .A(n10010), .ZN(n9985) );
  INV_X1 U6429 ( .A(n9989), .ZN(n10019) );
  OR2_X1 U6430 ( .A1(n6862), .A2(n6861), .ZN(n10116) );
  XNOR2_X1 U6431 ( .A(n5718), .B(n8050), .ZN(n9395) );
  AND2_X1 U6432 ( .A1(n10015), .A2(n9473), .ZN(n9823) );
  AND2_X1 U6433 ( .A1(n6524), .A2(n6523), .ZN(n6533) );
  INV_X1 U6434 ( .A(n9473), .ZN(n10099) );
  INV_X1 U6435 ( .A(n5657), .ZN(n5658) );
  INV_X1 U6436 ( .A(n10240), .ZN(n10234) );
  AND2_X1 U6437 ( .A1(n6219), .A2(n10218), .ZN(n10143) );
  NAND2_X1 U6438 ( .A1(n6107), .A2(n6106), .ZN(n8564) );
  INV_X1 U6439 ( .A(n10166), .ZN(n10152) );
  OR2_X1 U6440 ( .A1(n6904), .A2(n6204), .ZN(n10219) );
  AND3_X1 U6441 ( .A1(n8750), .A2(n8749), .A3(n8748), .ZN(n8842) );
  INV_X1 U6442 ( .A(n10319), .ZN(n10317) );
  INV_X1 U6443 ( .A(n10306), .ZN(n10304) );
  INV_X1 U6444 ( .A(n10235), .ZN(n10237) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n9678) );
  INV_X1 U6446 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6265) );
  NAND2_X1 U6447 ( .A1(n5588), .A2(n5587), .ZN(n9143) );
  OR2_X1 U6448 ( .A1(n10021), .A2(n6377), .ZN(n10029) );
  OR3_X1 U6449 ( .A1(n9387), .A2(n6527), .A3(n7770), .ZN(n9323) );
  AND2_X1 U6450 ( .A1(n9830), .A2(n9829), .ZN(n9845) );
  NAND2_X1 U6451 ( .A1(n6525), .A2(n6533), .ZN(n10124) );
  CLKBUF_X1 U6452 ( .A(n10062), .Z(n10069) );
  NAND2_X1 U6453 ( .A1(n6384), .A2(n5099), .ZN(n10072) );
  NOR2_X1 U6454 ( .A1(n10347), .A2(n10346), .ZN(n10345) );
  NAND3_X1 U6455 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5224) );
  INV_X1 U6456 ( .A(n5224), .ZN(n5050) );
  NAND2_X1 U6457 ( .A1(n5050), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5234) );
  INV_X1 U6458 ( .A(n5234), .ZN(n5051) );
  NAND2_X1 U6459 ( .A1(n5051), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5265) );
  INV_X1 U6460 ( .A(n5265), .ZN(n5052) );
  AND2_X1 U6461 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n5053) );
  INV_X1 U6462 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9622) );
  INV_X1 U6463 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5340) );
  INV_X1 U6464 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5395) );
  INV_X1 U6465 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8894) );
  INV_X1 U6466 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8953) );
  NAND2_X1 U6467 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5058) );
  INV_X1 U6468 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8982) );
  INV_X1 U6469 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5562) );
  INV_X1 U6470 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5561) );
  INV_X1 U6471 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5613) );
  INV_X1 U6472 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5612) );
  INV_X1 U6473 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5065) );
  INV_X1 U6474 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5066) );
  NOR2_X1 U6475 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5083) );
  NAND3_X1 U6476 ( .A1(n5084), .A2(n5083), .A3(n5314), .ZN(n5070) );
  INV_X1 U6477 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5443) );
  INV_X1 U6478 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5068) );
  INV_X1 U6479 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5067) );
  NAND4_X1 U6480 ( .A1(n5443), .A2(n5068), .A3(n5067), .A4(n5079), .ZN(n5069)
         );
  INV_X1 U6481 ( .A(n5107), .ZN(n5072) );
  INV_X1 U6482 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5071) );
  NAND2_X1 U6483 ( .A1(n5072), .A2(n5071), .ZN(n5100) );
  INV_X1 U6484 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5109) );
  INV_X1 U6485 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5105) );
  NAND3_X1 U6486 ( .A1(n5102), .A2(n5109), .A3(n5105), .ZN(n5073) );
  NAND2_X1 U6487 ( .A1(n5096), .A2(n5095), .ZN(n5098) );
  NOR2_X1 U6488 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5077) );
  NOR2_X1 U6489 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5076) );
  NAND4_X1 U6490 ( .A1(n5077), .A2(n5076), .A3(n5075), .A4(n5314), .ZN(n5078)
         );
  NOR2_X1 U6491 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5082) );
  NOR2_X1 U6492 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5081) );
  NOR2_X1 U6493 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5080) );
  NAND4_X1 U6494 ( .A1(n5083), .A2(n5082), .A3(n5081), .A4(n5080), .ZN(n5086)
         );
  NAND3_X1 U6495 ( .A1(n5084), .A2(n5102), .A3(n5095), .ZN(n5085) );
  NOR2_X1 U6496 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  NAND2_X1 U6497 ( .A1(n5089), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5088) );
  MUX2_X1 U6498 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5088), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n5090) );
  NAND2_X1 U6499 ( .A1(n5090), .A2(n5114), .ZN(n7573) );
  INV_X1 U6500 ( .A(n7573), .ZN(n5094) );
  NAND2_X1 U6501 ( .A1(n4423), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5092) );
  XNOR2_X1 U6502 ( .A(n5092), .B(n5091), .ZN(n7549) );
  INV_X1 U6503 ( .A(n7549), .ZN(n5093) );
  NAND2_X2 U6504 ( .A1(n5657), .A2(n5043), .ZN(n6384) );
  OR2_X1 U6505 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  NAND2_X1 U6506 ( .A1(n5098), .A2(n5097), .ZN(n7418) );
  AND2_X1 U6507 ( .A1(n7418), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5099) );
  NAND2_X1 U6508 ( .A1(n5110), .A2(n5109), .ZN(n5101) );
  NOR2_X1 U6509 ( .A1(n10072), .A2(n4392), .ZN(n5111) );
  NAND2_X1 U6510 ( .A1(n5103), .A2(n5102), .ZN(n5104) );
  NAND2_X1 U6511 ( .A1(n5107), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5108) );
  NAND2_X2 U6512 ( .A1(n7934), .A2(n9192), .ZN(n7933) );
  XNOR2_X1 U6513 ( .A(n5110), .B(n5109), .ZN(n8093) );
  INV_X1 U6514 ( .A(n8093), .ZN(n5653) );
  OR2_X1 U6515 ( .A1(n7934), .A2(n8092), .ZN(n5113) );
  NAND2_X1 U6516 ( .A1(n4392), .A2(n5653), .ZN(n5112) );
  INV_X1 U6517 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5127) );
  XNOR2_X2 U6518 ( .A(n5115), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5121) );
  XNOR2_X2 U6519 ( .A(n5118), .B(n5117), .ZN(n5120) );
  INV_X1 U6520 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6235) );
  NAND2_X2 U6521 ( .A1(n5121), .A2(n5119), .ZN(n5452) );
  INV_X1 U6522 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6505) );
  OR2_X1 U6523 ( .A1(n5452), .A2(n6505), .ZN(n5124) );
  INV_X1 U6524 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6243) );
  INV_X1 U6525 ( .A(n6492), .ZN(n5135) );
  INV_X1 U6526 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5129) );
  INV_X1 U6527 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5131) );
  INV_X1 U6528 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9621) );
  XNOR2_X1 U6529 ( .A(n5156), .B(SI_1_), .ZN(n5155) );
  MUX2_X1 U6530 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5134), .Z(n5154) );
  XNOR2_X1 U6531 ( .A(n5155), .B(n5154), .ZN(n6269) );
  INV_X1 U6532 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6389) );
  INV_X1 U6533 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6865) );
  NAND2_X1 U6534 ( .A1(n5178), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U6535 ( .A1(n5136), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5137) );
  NAND4_X2 U6536 ( .A1(n5140), .A2(n5139), .A3(n5138), .A4(n5137), .ZN(n6388)
         );
  INV_X1 U6537 ( .A(SI_0_), .ZN(n5141) );
  NOR2_X1 U6538 ( .A1(n7800), .A2(n5141), .ZN(n5142) );
  XNOR2_X1 U6539 ( .A(n5142), .B(n5132), .ZN(n9783) );
  INV_X1 U6540 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10128) );
  INV_X1 U6541 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5144) );
  INV_X1 U6542 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6557) );
  NOR2_X1 U6543 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5151) );
  INV_X1 U6544 ( .A(n5151), .ZN(n5149) );
  NAND2_X1 U6545 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n5149), .ZN(n5150) );
  INV_X1 U6546 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5152) );
  MUX2_X1 U6547 ( .A(n5150), .B(P1_IR_REG_31__SCAN_IN), .S(n5152), .Z(n5153)
         );
  NAND2_X1 U6548 ( .A1(n5152), .A2(n5151), .ZN(n5168) );
  INV_X1 U6549 ( .A(n9860), .ZN(n6262) );
  NAND2_X1 U6550 ( .A1(n5155), .A2(n5154), .ZN(n5159) );
  INV_X1 U6551 ( .A(n5156), .ZN(n5157) );
  NAND2_X1 U6552 ( .A1(n5157), .A2(SI_1_), .ZN(n5158) );
  NAND2_X1 U6553 ( .A1(n5159), .A2(n5158), .ZN(n5171) );
  INV_X1 U6554 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6257) );
  INV_X1 U6555 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6260) );
  MUX2_X1 U6556 ( .A(n6257), .B(n6260), .S(n5134), .Z(n5172) );
  XNOR2_X1 U6557 ( .A(n5171), .B(n5170), .ZN(n6261) );
  OR2_X1 U6558 ( .A1(n5219), .A2(n6261), .ZN(n5161) );
  OAI211_X2 U6559 ( .C1(n6190), .C2(n6262), .A(n5161), .B(n5160), .ZN(n10023)
         );
  OR2_X2 U6560 ( .A1(n6542), .A2(n10028), .ZN(n8064) );
  NAND2_X1 U6561 ( .A1(n6542), .A2(n10028), .ZN(n8062) );
  NAND2_X1 U6562 ( .A1(n5178), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5167) );
  INV_X1 U6563 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5162) );
  OR2_X1 U6564 ( .A1(n5485), .A2(n5162), .ZN(n5166) );
  OR2_X1 U6565 ( .A1(n5452), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5165) );
  INV_X1 U6566 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5163) );
  OR2_X1 U6567 ( .A1(n5179), .A2(n5163), .ZN(n5164) );
  NAND2_X1 U6568 ( .A1(n5168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5169) );
  XNOR2_X1 U6569 ( .A(n5169), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6328) );
  INV_X1 U6570 ( .A(n6328), .ZN(n6264) );
  INV_X1 U6571 ( .A(n5172), .ZN(n5173) );
  NAND2_X1 U6572 ( .A1(n5173), .A2(SI_2_), .ZN(n5174) );
  INV_X1 U6573 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6258) );
  MUX2_X1 U6574 ( .A(n6258), .B(n9547), .S(n5134), .Z(n5191) );
  XNOR2_X1 U6575 ( .A(n5191), .B(SI_3_), .ZN(n5189) );
  XNOR2_X1 U6576 ( .A(n5190), .B(n5189), .ZN(n6263) );
  OR2_X1 U6577 ( .A1(n5219), .A2(n6263), .ZN(n5176) );
  OR2_X1 U6578 ( .A1(n7806), .A2(n9547), .ZN(n5175) );
  OR2_X1 U6579 ( .A1(n10009), .A2(n10087), .ZN(n8063) );
  INV_X1 U6580 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6330) );
  OR2_X1 U6581 ( .A1(n6484), .A2(n6330), .ZN(n5183) );
  NAND2_X1 U6582 ( .A1(n6478), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5182) );
  XNOR2_X1 U6583 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n9993) );
  INV_X1 U6584 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6321) );
  OR2_X1 U6585 ( .A1(n6480), .A2(n6321), .ZN(n5180) );
  NAND4_X2 U6586 ( .A1(n5183), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n9038)
         );
  INV_X1 U6587 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5280) );
  NOR2_X1 U6588 ( .A1(n5184), .A2(n5280), .ZN(n5185) );
  MUX2_X1 U6589 ( .A(n5280), .B(n5185), .S(P1_IR_REG_4__SCAN_IN), .Z(n5186) );
  INV_X1 U6590 ( .A(n5186), .ZN(n5188) );
  NAND2_X1 U6591 ( .A1(n5188), .A2(n5187), .ZN(n6329) );
  INV_X1 U6592 ( .A(n5191), .ZN(n5192) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6267) );
  MUX2_X1 U6594 ( .A(n9744), .B(n6267), .S(n6259), .Z(n5207) );
  XNOR2_X1 U6595 ( .A(n5207), .B(SI_4_), .ZN(n5205) );
  XNOR2_X1 U6596 ( .A(n5206), .B(n5205), .ZN(n6268) );
  OR2_X1 U6597 ( .A1(n5219), .A2(n6268), .ZN(n5194) );
  OR2_X1 U6598 ( .A1(n7806), .A2(n6267), .ZN(n5193) );
  OAI211_X1 U6599 ( .C1(n6190), .C2(n6329), .A(n5194), .B(n5193), .ZN(n9998)
         );
  NAND2_X1 U6600 ( .A1(n9038), .A2(n10093), .ZN(n7945) );
  NAND2_X1 U6601 ( .A1(n10009), .A2(n10087), .ZN(n9981) );
  AND2_X1 U6602 ( .A1(n7945), .A2(n9981), .ZN(n8070) );
  NAND2_X1 U6603 ( .A1(n9982), .A2(n8070), .ZN(n5195) );
  OR2_X1 U6604 ( .A1(n9038), .A2(n10093), .ZN(n8067) );
  NAND2_X1 U6605 ( .A1(n6478), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5203) );
  INV_X1 U6606 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5196) );
  OR2_X1 U6607 ( .A1(n5485), .A2(n5196), .ZN(n5202) );
  INV_X1 U6608 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5198) );
  NAND2_X1 U6609 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5197) );
  NAND2_X1 U6610 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  NAND2_X1 U6611 ( .A1(n5224), .A2(n5199), .ZN(n7106) );
  OR2_X1 U6612 ( .A1(n5452), .A2(n7106), .ZN(n5201) );
  INV_X1 U6613 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5200) );
  NAND2_X1 U6614 ( .A1(n5187), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5204) );
  XNOR2_X1 U6615 ( .A(n5204), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9901) );
  INV_X1 U6616 ( .A(n9901), .ZN(n6320) );
  INV_X1 U6617 ( .A(n5207), .ZN(n5208) );
  NAND2_X1 U6618 ( .A1(n5208), .A2(SI_4_), .ZN(n5209) );
  NAND2_X1 U6619 ( .A1(n5210), .A2(n5209), .ZN(n5214) );
  MUX2_X1 U6620 ( .A(n6265), .B(n9730), .S(n6259), .Z(n5215) );
  OR2_X1 U6621 ( .A1(n6266), .A2(n5219), .ZN(n5212) );
  OR2_X1 U6622 ( .A1(n7806), .A2(n9730), .ZN(n5211) );
  INV_X1 U6623 ( .A(n7102), .ZN(n10105) );
  NOR2_X1 U6624 ( .A1(n9986), .A2(n10105), .ZN(n5690) );
  NAND2_X1 U6625 ( .A1(n9986), .A2(n10105), .ZN(n7822) );
  NAND2_X1 U6626 ( .A1(n7818), .A2(n7822), .ZN(n7819) );
  NAND2_X1 U6627 ( .A1(n5214), .A2(n5213), .ZN(n5218) );
  INV_X1 U6628 ( .A(n5215), .ZN(n5216) );
  NAND2_X1 U6629 ( .A1(n5216), .A2(SI_5_), .ZN(n5217) );
  MUX2_X1 U6630 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n6259), .Z(n5243) );
  XNOR2_X2 U6631 ( .A(n5243), .B(SI_6_), .ZN(n5240) );
  XNOR2_X1 U6632 ( .A(n5242), .B(n5240), .ZN(n6270) );
  INV_X2 U6633 ( .A(n5219), .ZN(n7804) );
  NAND2_X1 U6634 ( .A1(n6270), .A2(n7804), .ZN(n5223) );
  NAND2_X1 U6635 ( .A1(n5220), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6636 ( .A(n5221), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6331) );
  AOI22_X1 U6637 ( .A1(n5466), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5465), .B2(
        n6331), .ZN(n5222) );
  NAND2_X1 U6638 ( .A1(n5223), .A2(n5222), .ZN(n7095) );
  NAND2_X1 U6639 ( .A1(n6478), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5229) );
  INV_X1 U6640 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6326) );
  OR2_X1 U6641 ( .A1(n6484), .A2(n6326), .ZN(n5228) );
  INV_X1 U6642 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6344) );
  NAND2_X1 U6643 ( .A1(n5224), .A2(n6344), .ZN(n5225) );
  NAND2_X1 U6644 ( .A1(n5234), .A2(n5225), .ZN(n7084) );
  OR2_X1 U6645 ( .A1(n5582), .A2(n7084), .ZN(n5227) );
  OR2_X1 U6646 ( .A1(n6480), .A2(n4666), .ZN(n5226) );
  NAND4_X1 U6647 ( .A1(n5229), .A2(n5228), .A3(n5227), .A4(n5226), .ZN(n9037)
         );
  NAND2_X1 U6648 ( .A1(n6786), .A2(n9037), .ZN(n7827) );
  INV_X1 U6649 ( .A(n7827), .ZN(n5230) );
  OR2_X1 U6650 ( .A1(n9037), .A2(n6786), .ZN(n8074) );
  NAND2_X1 U6651 ( .A1(n6478), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5239) );
  INV_X1 U6652 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5231) );
  OR2_X1 U6653 ( .A1(n6484), .A2(n5231), .ZN(n5238) );
  INV_X1 U6654 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5232) );
  OR2_X1 U6655 ( .A1(n6480), .A2(n5232), .ZN(n5237) );
  INV_X1 U6656 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5233) );
  NAND2_X1 U6657 ( .A1(n5234), .A2(n5233), .ZN(n5235) );
  NAND2_X1 U6658 ( .A1(n5265), .A2(n5235), .ZN(n6805) );
  OR2_X1 U6659 ( .A1(n5582), .A2(n6805), .ZN(n5236) );
  NAND4_X1 U6660 ( .A1(n5239), .A2(n5238), .A3(n5237), .A4(n5236), .ZN(n9036)
         );
  INV_X1 U6661 ( .A(n9036), .ZN(n9967) );
  NAND2_X1 U6662 ( .A1(n5243), .A2(SI_6_), .ZN(n5244) );
  MUX2_X1 U6663 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6259), .Z(n5252) );
  XNOR2_X1 U6664 ( .A(n5251), .B(n5249), .ZN(n6273) );
  NAND2_X1 U6665 ( .A1(n6273), .A2(n7804), .ZN(n5248) );
  OR2_X1 U6666 ( .A1(n5245), .A2(n5280), .ZN(n5246) );
  XNOR2_X1 U6667 ( .A(n5246), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6366) );
  AOI22_X1 U6668 ( .A1(n5466), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5465), .B2(
        n6366), .ZN(n5247) );
  NAND2_X1 U6669 ( .A1(n5248), .A2(n5247), .ZN(n6703) );
  OR2_X1 U6670 ( .A1(n9967), .A2(n6703), .ZN(n7828) );
  NAND2_X1 U6671 ( .A1(n9967), .A2(n6703), .ZN(n7995) );
  INV_X1 U6672 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6282) );
  INV_X1 U6673 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6280) );
  MUX2_X1 U6674 ( .A(n6282), .B(n6280), .S(n6259), .Z(n5254) );
  INV_X1 U6675 ( .A(SI_8_), .ZN(n5253) );
  INV_X1 U6676 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6677 ( .A1(n5255), .A2(SI_8_), .ZN(n5256) );
  XNOR2_X1 U6678 ( .A(n5274), .B(n5273), .ZN(n6279) );
  NAND2_X1 U6679 ( .A1(n6279), .A2(n7804), .ZN(n5264) );
  NOR2_X1 U6680 ( .A1(n5257), .A2(n5280), .ZN(n5258) );
  MUX2_X1 U6681 ( .A(n5280), .B(n5258), .S(P1_IR_REG_8__SCAN_IN), .Z(n5259) );
  INV_X1 U6682 ( .A(n5259), .ZN(n5262) );
  INV_X1 U6683 ( .A(n5260), .ZN(n5261) );
  AOI22_X1 U6684 ( .A1(n5466), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5465), .B2(
        n9914), .ZN(n5263) );
  NAND2_X1 U6685 ( .A1(n5264), .A2(n5263), .ZN(n9968) );
  NAND2_X1 U6686 ( .A1(n6478), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5271) );
  INV_X1 U6687 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6358) );
  OR2_X1 U6688 ( .A1(n6484), .A2(n6358), .ZN(n5270) );
  INV_X1 U6689 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6889) );
  NAND2_X1 U6690 ( .A1(n5265), .A2(n6889), .ZN(n5266) );
  NAND2_X1 U6691 ( .A1(n5305), .A2(n5266), .ZN(n9969) );
  OR2_X1 U6692 ( .A1(n5582), .A2(n9969), .ZN(n5269) );
  INV_X1 U6693 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5267) );
  OR2_X1 U6694 ( .A1(n6480), .A2(n5267), .ZN(n5268) );
  NAND4_X1 U6695 ( .A1(n5271), .A2(n5270), .A3(n5269), .A4(n5268), .ZN(n9035)
         );
  INV_X1 U6696 ( .A(n9035), .ZN(n6704) );
  NAND2_X1 U6697 ( .A1(n9968), .A2(n6704), .ZN(n7996) );
  INV_X1 U6698 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6299) );
  INV_X1 U6699 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5275) );
  MUX2_X1 U6700 ( .A(n6299), .B(n5275), .S(n6259), .Z(n5277) );
  INV_X1 U6701 ( .A(SI_9_), .ZN(n5276) );
  INV_X1 U6702 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6703 ( .A1(n5278), .A2(SI_9_), .ZN(n5279) );
  XNOR2_X1 U6704 ( .A(n5290), .B(n5046), .ZN(n6292) );
  NAND2_X1 U6705 ( .A1(n6292), .A2(n7804), .ZN(n5283) );
  OR2_X1 U6706 ( .A1(n5260), .A2(n5280), .ZN(n5281) );
  XNOR2_X1 U6707 ( .A(n5281), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9924) );
  AOI22_X1 U6708 ( .A1(n5466), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5465), .B2(
        n9924), .ZN(n5282) );
  NAND2_X1 U6709 ( .A1(n6478), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5288) );
  INV_X1 U6710 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5284) );
  OR2_X1 U6711 ( .A1(n6484), .A2(n5284), .ZN(n5287) );
  INV_X1 U6712 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7061) );
  XNOR2_X1 U6713 ( .A(n5305), .B(n7061), .ZN(n7062) );
  OR2_X1 U6714 ( .A1(n5582), .A2(n7062), .ZN(n5286) );
  INV_X1 U6715 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6367) );
  OR2_X1 U6716 ( .A1(n6480), .A2(n6367), .ZN(n5285) );
  NAND4_X1 U6717 ( .A1(n5288), .A2(n5287), .A3(n5286), .A4(n5285), .ZN(n9034)
         );
  INV_X1 U6718 ( .A(n9034), .ZN(n9966) );
  NOR2_X1 U6719 ( .A1(n7195), .A2(n9966), .ZN(n7824) );
  INV_X1 U6720 ( .A(n7824), .ZN(n7011) );
  OR2_X1 U6721 ( .A1(n9968), .A2(n6704), .ZN(n7013) );
  AND2_X1 U6722 ( .A1(n7011), .A2(n7013), .ZN(n7972) );
  NAND2_X1 U6723 ( .A1(n7195), .A2(n9966), .ZN(n7967) );
  INV_X1 U6724 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5294) );
  INV_X1 U6725 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n5293) );
  MUX2_X1 U6726 ( .A(n5294), .B(n5293), .S(n6259), .Z(n5296) );
  INV_X1 U6727 ( .A(SI_10_), .ZN(n5295) );
  INV_X1 U6728 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6729 ( .A1(n5297), .A2(SI_10_), .ZN(n5298) );
  NAND2_X1 U6730 ( .A1(n6300), .A2(n7804), .ZN(n5301) );
  NAND2_X1 U6731 ( .A1(n5299), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5315) );
  XNOR2_X1 U6732 ( .A(n5315), .B(P1_IR_REG_10__SCAN_IN), .ZN(n6607) );
  AOI22_X1 U6733 ( .A1(n5466), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5465), .B2(
        n6607), .ZN(n5300) );
  NAND2_X1 U6734 ( .A1(n6478), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5310) );
  INV_X1 U6735 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n5302) );
  OR2_X1 U6736 ( .A1(n6484), .A2(n5302), .ZN(n5309) );
  INV_X1 U6737 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n5303) );
  OR2_X1 U6738 ( .A1(n6480), .A2(n5303), .ZN(n5308) );
  INV_X1 U6739 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5304) );
  OAI21_X1 U6740 ( .B1(n5305), .B2(n7061), .A(n5304), .ZN(n5306) );
  NAND2_X1 U6741 ( .A1(n5306), .A2(n5321), .ZN(n7327) );
  OR2_X1 U6742 ( .A1(n5582), .A2(n7327), .ZN(n5307) );
  NAND4_X1 U6743 ( .A1(n5310), .A2(n5309), .A3(n5308), .A4(n5307), .ZN(n9033)
         );
  INV_X1 U6744 ( .A(n9033), .ZN(n5311) );
  NAND2_X1 U6745 ( .A1(n7326), .A2(n5311), .ZN(n7968) );
  NAND2_X1 U6746 ( .A1(n7973), .A2(n7968), .ZN(n8039) );
  INV_X1 U6747 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6316) );
  INV_X1 U6748 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6317) );
  MUX2_X1 U6749 ( .A(n6316), .B(n6317), .S(n6259), .Z(n5328) );
  NAND2_X1 U6750 ( .A1(n6315), .A2(n7804), .ZN(n5319) );
  NAND2_X1 U6751 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  NAND2_X1 U6752 ( .A1(n5316), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  XNOR2_X1 U6753 ( .A(n5317), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9929) );
  AOI22_X1 U6754 ( .A1(n5466), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5465), .B2(
        n9929), .ZN(n5318) );
  NAND2_X1 U6755 ( .A1(n6478), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5326) );
  INV_X1 U6756 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5320) );
  OR2_X1 U6757 ( .A1(n6484), .A2(n5320), .ZN(n5325) );
  NAND2_X1 U6758 ( .A1(n5321), .A2(n9622), .ZN(n5322) );
  NAND2_X1 U6759 ( .A1(n5341), .A2(n5322), .ZN(n8990) );
  OR2_X1 U6760 ( .A1(n5582), .A2(n8990), .ZN(n5324) );
  INV_X1 U6761 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7276) );
  OR2_X1 U6762 ( .A1(n6480), .A2(n7276), .ZN(n5323) );
  INV_X1 U6763 ( .A(n9032), .ZN(n7435) );
  NAND2_X1 U6764 ( .A1(n9468), .A2(n7435), .ZN(n7839) );
  NAND2_X1 U6765 ( .A1(n7268), .A2(n7839), .ZN(n7432) );
  INV_X1 U6766 ( .A(n5328), .ZN(n5329) );
  INV_X1 U6767 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6356) );
  INV_X1 U6768 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6354) );
  MUX2_X1 U6769 ( .A(n6356), .B(n6354), .S(n6259), .Z(n5333) );
  INV_X1 U6770 ( .A(SI_12_), .ZN(n5332) );
  INV_X1 U6771 ( .A(n5333), .ZN(n5334) );
  NAND2_X1 U6772 ( .A1(n5334), .A2(SI_12_), .ZN(n5335) );
  XNOR2_X1 U6773 ( .A(n5351), .B(n5350), .ZN(n6353) );
  NAND2_X1 U6774 ( .A1(n6353), .A2(n7804), .ZN(n5339) );
  OR2_X1 U6775 ( .A1(n4502), .A2(n5280), .ZN(n5337) );
  XNOR2_X1 U6776 ( .A(n5337), .B(P1_IR_REG_12__SCAN_IN), .ZN(n6643) );
  AOI22_X1 U6777 ( .A1(n5466), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5465), .B2(
        n6643), .ZN(n5338) );
  NAND2_X1 U6778 ( .A1(n6478), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5347) );
  INV_X1 U6779 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6600) );
  OR2_X1 U6780 ( .A1(n6484), .A2(n6600), .ZN(n5346) );
  NAND2_X1 U6781 ( .A1(n5341), .A2(n5340), .ZN(n5342) );
  NAND2_X1 U6782 ( .A1(n5361), .A2(n5342), .ZN(n7440) );
  OR2_X1 U6783 ( .A1(n5582), .A2(n7440), .ZN(n5345) );
  INV_X1 U6784 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n5343) );
  OR2_X1 U6785 ( .A1(n6480), .A2(n5343), .ZN(n5344) );
  NAND4_X1 U6786 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n9031)
         );
  INV_X1 U6787 ( .A(n9031), .ZN(n9367) );
  NOR2_X1 U6788 ( .A1(n9464), .A2(n9367), .ZN(n7841) );
  INV_X1 U6789 ( .A(n7841), .ZN(n5701) );
  OR2_X1 U6790 ( .A1(n9468), .A2(n7435), .ZN(n7431) );
  AND2_X1 U6791 ( .A1(n5701), .A2(n7431), .ZN(n7974) );
  NAND2_X1 U6792 ( .A1(n7432), .A2(n7974), .ZN(n5348) );
  NAND2_X1 U6793 ( .A1(n9464), .A2(n9367), .ZN(n7976) );
  INV_X1 U6794 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n5352) );
  MUX2_X1 U6795 ( .A(n9678), .B(n5352), .S(n6259), .Z(n5354) );
  INV_X1 U6796 ( .A(SI_13_), .ZN(n5353) );
  NAND2_X1 U6797 ( .A1(n5354), .A2(n5353), .ZN(n5368) );
  INV_X1 U6798 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6799 ( .A1(n5355), .A2(SI_13_), .ZN(n5356) );
  XNOR2_X1 U6800 ( .A(n5367), .B(n5047), .ZN(n6396) );
  NAND2_X1 U6801 ( .A1(n6396), .A2(n7804), .ZN(n5360) );
  OR2_X1 U6802 ( .A1(n5357), .A2(n5280), .ZN(n5358) );
  XNOR2_X1 U6803 ( .A(n5358), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7006) );
  AOI22_X1 U6804 ( .A1(n5466), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5465), .B2(
        n7006), .ZN(n5359) );
  NAND2_X1 U6805 ( .A1(n6478), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5366) );
  INV_X1 U6806 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6634) );
  OR2_X1 U6807 ( .A1(n6484), .A2(n6634), .ZN(n5365) );
  INV_X1 U6808 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U6809 ( .A1(n5361), .A2(n6633), .ZN(n5362) );
  NAND2_X1 U6810 ( .A1(n5396), .A2(n5362), .ZN(n9380) );
  OR2_X1 U6811 ( .A1(n5452), .A2(n9380), .ZN(n5364) );
  INV_X1 U6812 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6644) );
  OR2_X1 U6813 ( .A1(n6480), .A2(n6644), .ZN(n5363) );
  NAND4_X1 U6814 ( .A1(n5366), .A2(n5365), .A3(n5364), .A4(n5363), .ZN(n9030)
         );
  INV_X1 U6815 ( .A(n9030), .ZN(n9356) );
  OR2_X1 U6816 ( .A1(n9457), .A2(n9356), .ZN(n7847) );
  NAND2_X1 U6817 ( .A1(n9457), .A2(n9356), .ZN(n7978) );
  INV_X1 U6818 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6489) );
  INV_X1 U6819 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6490) );
  MUX2_X1 U6820 ( .A(n6489), .B(n6490), .S(n6259), .Z(n5378) );
  XNOR2_X1 U6821 ( .A(n5382), .B(n5377), .ZN(n6488) );
  NAND2_X1 U6822 ( .A1(n6488), .A2(n7804), .ZN(n5371) );
  INV_X1 U6823 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5369) );
  AND2_X1 U6824 ( .A1(n5357), .A2(n5369), .ZN(n5409) );
  OR2_X1 U6825 ( .A1(n5409), .A2(n5280), .ZN(n5388) );
  XNOR2_X1 U6826 ( .A(n5388), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9047) );
  AOI22_X1 U6827 ( .A1(n5466), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5465), .B2(
        n9047), .ZN(n5370) );
  NAND2_X1 U6828 ( .A1(n6478), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5376) );
  INV_X1 U6829 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6997) );
  OR2_X1 U6830 ( .A1(n6484), .A2(n6997), .ZN(n5375) );
  INV_X1 U6831 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5372) );
  OR2_X1 U6832 ( .A1(n6480), .A2(n5372), .ZN(n5374) );
  XNOR2_X1 U6833 ( .A(n5396), .B(n8894), .ZN(n9348) );
  OR2_X1 U6834 ( .A1(n5582), .A2(n9348), .ZN(n5373) );
  NAND4_X1 U6835 ( .A1(n5376), .A2(n5375), .A3(n5374), .A4(n5373), .ZN(n9327)
         );
  XNOR2_X1 U6836 ( .A(n9351), .B(n9327), .ZN(n9343) );
  INV_X1 U6837 ( .A(n9343), .ZN(n9354) );
  INV_X1 U6838 ( .A(n9327), .ZN(n9368) );
  OR2_X1 U6839 ( .A1(n9351), .A2(n9368), .ZN(n7850) );
  NAND2_X1 U6840 ( .A1(n9359), .A2(n7850), .ZN(n9330) );
  INV_X1 U6841 ( .A(n5378), .ZN(n5379) );
  NAND2_X1 U6842 ( .A1(n5379), .A2(SI_14_), .ZN(n5380) );
  INV_X1 U6843 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6616) );
  INV_X1 U6844 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6617) );
  MUX2_X1 U6845 ( .A(n6616), .B(n6617), .S(n6259), .Z(n5384) );
  INV_X1 U6846 ( .A(SI_15_), .ZN(n5383) );
  INV_X1 U6847 ( .A(n5384), .ZN(n5385) );
  NAND2_X1 U6848 ( .A1(n5385), .A2(SI_15_), .ZN(n5386) );
  XNOR2_X1 U6849 ( .A(n5404), .B(n5403), .ZN(n6615) );
  NAND2_X1 U6850 ( .A1(n6615), .A2(n7804), .ZN(n5393) );
  INV_X1 U6851 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5387) );
  NAND2_X1 U6852 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  NAND2_X1 U6853 ( .A1(n5389), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5391) );
  INV_X1 U6854 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5390) );
  XNOR2_X1 U6855 ( .A(n5391), .B(n5390), .ZN(n9063) );
  INV_X1 U6856 ( .A(n9063), .ZN(n9051) );
  AOI22_X1 U6857 ( .A1(n5466), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5465), .B2(
        n9051), .ZN(n5392) );
  NAND2_X1 U6858 ( .A1(n5177), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5401) );
  INV_X1 U6859 ( .A(n6478), .ZN(n5616) );
  INV_X1 U6860 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5394) );
  OR2_X1 U6861 ( .A1(n5616), .A2(n5394), .ZN(n5400) );
  OAI21_X1 U6862 ( .B1(n5396), .B2(n8894), .A(n5395), .ZN(n5397) );
  NAND2_X1 U6863 ( .A1(n5397), .A2(n5414), .ZN(n9334) );
  OR2_X1 U6864 ( .A1(n5452), .A2(n9334), .ZN(n5399) );
  INV_X1 U6865 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9335) );
  OR2_X1 U6866 ( .A1(n6480), .A2(n9335), .ZN(n5398) );
  NAND4_X1 U6867 ( .A1(n5401), .A2(n5400), .A3(n5399), .A4(n5398), .ZN(n9311)
         );
  INV_X1 U6868 ( .A(n9311), .ZN(n9357) );
  NAND2_X1 U6869 ( .A1(n9340), .A2(n9357), .ZN(n7993) );
  NAND2_X1 U6870 ( .A1(n9307), .A2(n7993), .ZN(n7851) );
  NAND2_X1 U6871 ( .A1(n9329), .A2(n9307), .ZN(n5420) );
  INV_X1 U6872 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6626) );
  INV_X1 U6873 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9709) );
  MUX2_X1 U6874 ( .A(n6626), .B(n9709), .S(n6259), .Z(n5405) );
  INV_X1 U6875 ( .A(SI_16_), .ZN(n9584) );
  NAND2_X1 U6876 ( .A1(n5405), .A2(n9584), .ZN(n5422) );
  INV_X1 U6877 ( .A(n5405), .ZN(n5406) );
  NAND2_X1 U6878 ( .A1(n5406), .A2(SI_16_), .ZN(n5407) );
  XNOR2_X1 U6879 ( .A(n5421), .B(n5045), .ZN(n6625) );
  NAND2_X1 U6880 ( .A1(n6625), .A2(n7804), .ZN(n5412) );
  NOR2_X1 U6881 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5408) );
  NAND2_X1 U6882 ( .A1(n5409), .A2(n5408), .ZN(n5425) );
  NAND2_X1 U6883 ( .A1(n5425), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5410) );
  XNOR2_X1 U6884 ( .A(n5410), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9083) );
  AOI22_X1 U6885 ( .A1(n5466), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5465), .B2(
        n9083), .ZN(n5411) );
  NAND2_X1 U6886 ( .A1(n5177), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5419) );
  INV_X1 U6887 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n5413) );
  OR2_X1 U6888 ( .A1(n5616), .A2(n5413), .ZN(n5418) );
  INV_X1 U6889 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n8942) );
  NAND2_X1 U6890 ( .A1(n5414), .A2(n8942), .ZN(n5415) );
  NAND2_X1 U6891 ( .A1(n5429), .A2(n5415), .ZN(n9316) );
  OR2_X1 U6892 ( .A1(n5452), .A2(n9316), .ZN(n5417) );
  INV_X1 U6893 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9058) );
  OR2_X1 U6894 ( .A1(n6480), .A2(n9058), .ZN(n5416) );
  NAND4_X1 U6895 ( .A1(n5419), .A2(n5418), .A3(n5417), .A4(n5416), .ZN(n9328)
         );
  INV_X1 U6896 ( .A(n9328), .ZN(n9016) );
  NAND2_X1 U6897 ( .A1(n9318), .A2(n9016), .ZN(n7986) );
  NAND2_X1 U6898 ( .A1(n7859), .A2(n7986), .ZN(n9306) );
  NAND2_X1 U6899 ( .A1(n9309), .A2(n7859), .ZN(n9297) );
  NAND2_X1 U6900 ( .A1(n5421), .A2(n5045), .ZN(n5423) );
  INV_X1 U6901 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6632) );
  INV_X1 U6902 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5424) );
  MUX2_X1 U6903 ( .A(n6632), .B(n5424), .S(n6259), .Z(n5438) );
  XNOR2_X1 U6904 ( .A(n5438), .B(SI_17_), .ZN(n5437) );
  XNOR2_X1 U6905 ( .A(n5442), .B(n5437), .ZN(n6629) );
  NAND2_X1 U6906 ( .A1(n6629), .A2(n7804), .ZN(n5428) );
  OR2_X1 U6907 ( .A1(n5425), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6908 ( .A1(n5426), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5444) );
  XNOR2_X1 U6909 ( .A(n5444), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9102) );
  AOI22_X1 U6910 ( .A1(n5466), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5465), .B2(
        n9102), .ZN(n5427) );
  NAND2_X1 U6911 ( .A1(n6478), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5435) );
  INV_X1 U6912 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9084) );
  OR2_X1 U6913 ( .A1(n6484), .A2(n9084), .ZN(n5434) );
  NAND2_X1 U6914 ( .A1(n5429), .A2(n8953), .ZN(n5430) );
  NAND2_X1 U6915 ( .A1(n5450), .A2(n5430), .ZN(n9292) );
  OR2_X1 U6916 ( .A1(n5582), .A2(n9292), .ZN(n5433) );
  INV_X1 U6917 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5431) );
  OR2_X1 U6918 ( .A1(n6480), .A2(n5431), .ZN(n5432) );
  NAND4_X1 U6919 ( .A1(n5435), .A2(n5434), .A3(n5433), .A4(n5432), .ZN(n9310)
         );
  NOR2_X1 U6920 ( .A1(n9452), .A2(n5711), .ZN(n7957) );
  INV_X1 U6921 ( .A(n7957), .ZN(n5436) );
  NAND2_X1 U6922 ( .A1(n9452), .A2(n5711), .ZN(n7985) );
  NAND2_X1 U6923 ( .A1(n5436), .A2(n7985), .ZN(n9289) );
  INV_X1 U6924 ( .A(n9289), .ZN(n9296) );
  INV_X1 U6925 ( .A(n5437), .ZN(n5441) );
  INV_X1 U6926 ( .A(n5438), .ZN(n5439) );
  NAND2_X1 U6927 ( .A1(n5439), .A2(SI_17_), .ZN(n5440) );
  MUX2_X1 U6928 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6259), .Z(n5460) );
  XNOR2_X1 U6929 ( .A(n5460), .B(SI_18_), .ZN(n5457) );
  XNOR2_X1 U6930 ( .A(n5459), .B(n5457), .ZN(n6750) );
  NAND2_X1 U6931 ( .A1(n6750), .A2(n7804), .ZN(n5448) );
  NAND2_X1 U6932 ( .A1(n5444), .A2(n5443), .ZN(n5445) );
  NAND2_X1 U6933 ( .A1(n5445), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5446) );
  XNOR2_X1 U6934 ( .A(n5446), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9951) );
  AOI22_X1 U6935 ( .A1(n5466), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5465), .B2(
        n9951), .ZN(n5447) );
  NAND2_X1 U6936 ( .A1(n6478), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5456) );
  INV_X1 U6937 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9100) );
  OR2_X1 U6938 ( .A1(n5485), .A2(n9100), .ZN(n5455) );
  INV_X1 U6939 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6940 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NAND2_X1 U6941 ( .A1(n5488), .A2(n5451), .ZN(n9278) );
  OR2_X1 U6942 ( .A1(n5452), .A2(n9278), .ZN(n5454) );
  INV_X1 U6943 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9096) );
  OR2_X1 U6944 ( .A1(n6480), .A2(n9096), .ZN(n5453) );
  NAND4_X1 U6945 ( .A1(n5456), .A2(n5455), .A3(n5454), .A4(n5453), .ZN(n9298)
         );
  INV_X1 U6946 ( .A(n9298), .ZN(n8915) );
  OR2_X1 U6947 ( .A1(n9447), .A2(n8915), .ZN(n7954) );
  NAND2_X1 U6948 ( .A1(n9447), .A2(n8915), .ZN(n7987) );
  NAND2_X1 U6949 ( .A1(n7954), .A2(n7987), .ZN(n8043) );
  INV_X1 U6950 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6870) );
  INV_X1 U6951 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n6871) );
  MUX2_X1 U6952 ( .A(n6870), .B(n6871), .S(n6259), .Z(n5462) );
  INV_X1 U6953 ( .A(SI_19_), .ZN(n5461) );
  NAND2_X1 U6954 ( .A1(n5462), .A2(n5461), .ZN(n5475) );
  INV_X1 U6955 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U6956 ( .A1(n5463), .A2(SI_19_), .ZN(n5464) );
  NAND2_X1 U6957 ( .A1(n5475), .A2(n5464), .ZN(n5476) );
  XNOR2_X1 U6958 ( .A(n5477), .B(n5476), .ZN(n6869) );
  NAND2_X1 U6959 ( .A1(n6869), .A2(n7804), .ZN(n5468) );
  AOI22_X1 U6960 ( .A1(n5466), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9192), .B2(
        n5465), .ZN(n5467) );
  NAND2_X1 U6961 ( .A1(n6478), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5474) );
  INV_X1 U6962 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5469) );
  OR2_X1 U6963 ( .A1(n6484), .A2(n5469), .ZN(n5473) );
  INV_X1 U6964 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5487) );
  XNOR2_X1 U6965 ( .A(n5488), .B(n5487), .ZN(n9267) );
  OR2_X1 U6966 ( .A1(n5582), .A2(n9267), .ZN(n5472) );
  INV_X1 U6967 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5470) );
  OR2_X1 U6968 ( .A1(n6480), .A2(n5470), .ZN(n5471) );
  NAND4_X1 U6969 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n9284)
         );
  INV_X1 U6970 ( .A(n9284), .ZN(n9248) );
  OR2_X1 U6971 ( .A1(n9442), .A2(n9248), .ZN(n7959) );
  NAND2_X1 U6972 ( .A1(n9442), .A2(n9248), .ZN(n8003) );
  INV_X1 U6973 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n9717) );
  INV_X1 U6974 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7098) );
  MUX2_X1 U6975 ( .A(n9717), .B(n7098), .S(n6259), .Z(n5479) );
  INV_X1 U6976 ( .A(SI_20_), .ZN(n5478) );
  NAND2_X1 U6977 ( .A1(n5479), .A2(n5478), .ZN(n5496) );
  INV_X1 U6978 ( .A(n5479), .ZN(n5480) );
  NAND2_X1 U6979 ( .A1(n5480), .A2(SI_20_), .ZN(n5481) );
  XNOR2_X1 U6980 ( .A(n5495), .B(n5494), .ZN(n7097) );
  NAND2_X1 U6981 ( .A1(n7097), .A2(n7804), .ZN(n5483) );
  OR2_X1 U6982 ( .A1(n7806), .A2(n7098), .ZN(n5482) );
  NAND2_X1 U6983 ( .A1(n6478), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5493) );
  INV_X1 U6984 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5484) );
  OR2_X1 U6985 ( .A1(n5485), .A2(n5484), .ZN(n5492) );
  INV_X1 U6986 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5486) );
  OAI21_X1 U6987 ( .B1(n5488), .B2(n5487), .A(n5486), .ZN(n5489) );
  NAND2_X1 U6988 ( .A1(n5489), .A2(n5500), .ZN(n9253) );
  OR2_X1 U6989 ( .A1(n5582), .A2(n9253), .ZN(n5491) );
  INV_X1 U6990 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9254) );
  OR2_X1 U6991 ( .A1(n6480), .A2(n9254), .ZN(n5490) );
  NAND4_X1 U6992 ( .A1(n5493), .A2(n5492), .A3(n5491), .A4(n5490), .ZN(n9263)
         );
  INV_X1 U6993 ( .A(n9263), .ZN(n9230) );
  NOR2_X1 U6994 ( .A1(n9439), .A2(n9230), .ZN(n7884) );
  INV_X1 U6995 ( .A(n7884), .ZN(n7960) );
  NAND2_X1 U6996 ( .A1(n9439), .A2(n9230), .ZN(n7951) );
  INV_X1 U6997 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7161) );
  INV_X1 U6998 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7125) );
  MUX2_X1 U6999 ( .A(n7161), .B(n7125), .S(n6259), .Z(n5507) );
  XNOR2_X1 U7000 ( .A(n5507), .B(SI_21_), .ZN(n5506) );
  XNOR2_X1 U7001 ( .A(n5511), .B(n5506), .ZN(n7124) );
  NAND2_X1 U7002 ( .A1(n7124), .A2(n7804), .ZN(n5499) );
  OR2_X1 U7003 ( .A1(n7806), .A2(n7125), .ZN(n5498) );
  INV_X1 U7004 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U7005 ( .A1(n5500), .A2(n9746), .ZN(n5501) );
  NAND2_X1 U7006 ( .A1(n5518), .A2(n5501), .ZN(n9234) );
  OR2_X1 U7007 ( .A1(n9234), .A2(n5582), .ZN(n5505) );
  NAND2_X1 U7008 ( .A1(n5177), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7009 ( .A1(n5136), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5503) );
  NAND2_X1 U7010 ( .A1(n6478), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5502) );
  NAND4_X1 U7011 ( .A1(n5505), .A2(n5504), .A3(n5503), .A4(n5502), .ZN(n9212)
         );
  INV_X1 U7012 ( .A(n9212), .ZN(n9249) );
  OR2_X1 U7013 ( .A1(n9241), .A2(n9249), .ZN(n7962) );
  NAND2_X1 U7014 ( .A1(n9241), .A2(n9249), .ZN(n9209) );
  NAND2_X1 U7015 ( .A1(n7962), .A2(n9209), .ZN(n7885) );
  INV_X1 U7016 ( .A(n5506), .ZN(n5510) );
  INV_X1 U7017 ( .A(n5507), .ZN(n5508) );
  NAND2_X1 U7018 ( .A1(n5508), .A2(SI_21_), .ZN(n5509) );
  INV_X1 U7019 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7613) );
  INV_X1 U7020 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9583) );
  MUX2_X1 U7021 ( .A(n7613), .B(n9583), .S(n6259), .Z(n5513) );
  INV_X1 U7022 ( .A(SI_22_), .ZN(n5512) );
  NAND2_X1 U7023 ( .A1(n5513), .A2(n5512), .ZN(n5523) );
  INV_X1 U7024 ( .A(n5513), .ZN(n5514) );
  NAND2_X1 U7025 ( .A1(n5514), .A2(SI_22_), .ZN(n5515) );
  NAND2_X1 U7026 ( .A1(n5523), .A2(n5515), .ZN(n5524) );
  XNOR2_X1 U7027 ( .A(n5525), .B(n5524), .ZN(n7414) );
  NAND2_X1 U7028 ( .A1(n7414), .A2(n7804), .ZN(n5517) );
  OR2_X1 U7029 ( .A1(n7806), .A2(n9583), .ZN(n5516) );
  NAND2_X1 U7030 ( .A1(n5518), .A2(n8982), .ZN(n5519) );
  NAND2_X1 U7031 ( .A1(n5532), .A2(n5519), .ZN(n9217) );
  AOI22_X1 U7032 ( .A1(n5177), .A2(P1_REG1_REG_22__SCAN_IN), .B1(n6478), .B2(
        P1_REG0_REG_22__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7033 ( .A1(n5136), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5520) );
  OAI211_X1 U7034 ( .C1(n9217), .C2(n5582), .A(n5521), .B(n5520), .ZN(n9228)
         );
  INV_X1 U7035 ( .A(n9228), .ZN(n8924) );
  NAND2_X1 U7036 ( .A1(n9427), .A2(n8924), .ZN(n8027) );
  NAND2_X1 U7037 ( .A1(n8027), .A2(n9209), .ZN(n7953) );
  INV_X1 U7038 ( .A(n7953), .ZN(n5522) );
  INV_X1 U7039 ( .A(n8028), .ZN(n7891) );
  INV_X1 U7040 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7416) );
  INV_X1 U7041 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7420) );
  MUX2_X1 U7042 ( .A(n7416), .B(n7420), .S(n6259), .Z(n5527) );
  INV_X1 U7043 ( .A(SI_23_), .ZN(n5526) );
  NAND2_X1 U7044 ( .A1(n5527), .A2(n5526), .ZN(n5539) );
  INV_X1 U7045 ( .A(n5527), .ZN(n5528) );
  NAND2_X1 U7046 ( .A1(n5528), .A2(SI_23_), .ZN(n5529) );
  XNOR2_X1 U7047 ( .A(n5538), .B(n5537), .ZN(n7417) );
  NAND2_X1 U7048 ( .A1(n7417), .A2(n7804), .ZN(n5531) );
  OR2_X1 U7049 ( .A1(n7806), .A2(n7420), .ZN(n5530) );
  INV_X1 U7050 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n5536) );
  INV_X1 U7051 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U7052 ( .A1(n5532), .A2(n9668), .ZN(n5533) );
  NAND2_X1 U7053 ( .A1(n5563), .A2(n5533), .ZN(n9199) );
  OR2_X1 U7054 ( .A1(n9199), .A2(n5582), .ZN(n5535) );
  AOI22_X1 U7055 ( .A1(n5177), .A2(P1_REG1_REG_23__SCAN_IN), .B1(n6478), .B2(
        P1_REG0_REG_23__SCAN_IN), .ZN(n5534) );
  OAI211_X1 U7056 ( .C1(n6480), .C2(n5536), .A(n5535), .B(n5534), .ZN(n9211)
         );
  INV_X1 U7057 ( .A(n9211), .ZN(n9187) );
  NOR2_X1 U7058 ( .A1(n9422), .A2(n9187), .ZN(n7815) );
  INV_X1 U7059 ( .A(n7815), .ZN(n7897) );
  AND2_X1 U7060 ( .A1(n9422), .A2(n9187), .ZN(n8006) );
  INV_X1 U7061 ( .A(n8006), .ZN(n7900) );
  NAND2_X1 U7062 ( .A1(n7897), .A2(n7900), .ZN(n9203) );
  INV_X1 U7063 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7457) );
  INV_X1 U7064 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7731) );
  MUX2_X1 U7065 ( .A(n7457), .B(n7731), .S(n6259), .Z(n5550) );
  XNOR2_X1 U7066 ( .A(n5550), .B(SI_24_), .ZN(n5549) );
  XNOR2_X1 U7067 ( .A(n5554), .B(n5549), .ZN(n7456) );
  NAND2_X1 U7068 ( .A1(n7456), .A2(n7804), .ZN(n5542) );
  OR2_X1 U7069 ( .A1(n7806), .A2(n7731), .ZN(n5541) );
  XNOR2_X1 U7070 ( .A(n5563), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9190) );
  NAND2_X1 U7071 ( .A1(n9190), .A2(n5630), .ZN(n5547) );
  INV_X1 U7072 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9554) );
  NAND2_X1 U7073 ( .A1(n6478), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U7074 ( .A1(n5136), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5543) );
  OAI211_X1 U7075 ( .C1(n6484), .C2(n9554), .A(n5544), .B(n5543), .ZN(n5545)
         );
  INV_X1 U7076 ( .A(n5545), .ZN(n5546) );
  NAND2_X1 U7077 ( .A1(n5547), .A2(n5546), .ZN(n9204) );
  XNOR2_X1 U7078 ( .A(n9419), .B(n9204), .ZN(n8046) );
  INV_X1 U7079 ( .A(n9204), .ZN(n9175) );
  NAND2_X1 U7080 ( .A1(n9419), .A2(n9175), .ZN(n7899) );
  INV_X1 U7081 ( .A(n7899), .ZN(n5548) );
  INV_X1 U7082 ( .A(n5549), .ZN(n5553) );
  INV_X1 U7083 ( .A(n5550), .ZN(n5551) );
  NAND2_X1 U7084 ( .A1(n5551), .A2(SI_24_), .ZN(n5552) );
  INV_X1 U7085 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7546) );
  INV_X1 U7086 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7547) );
  MUX2_X1 U7087 ( .A(n7546), .B(n7547), .S(n6259), .Z(n5556) );
  INV_X1 U7088 ( .A(SI_25_), .ZN(n5555) );
  NAND2_X1 U7089 ( .A1(n5556), .A2(n5555), .ZN(n5570) );
  INV_X1 U7090 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U7091 ( .A1(n5557), .A2(SI_25_), .ZN(n5558) );
  NAND2_X1 U7092 ( .A1(n5570), .A2(n5558), .ZN(n5571) );
  OR2_X1 U7093 ( .A1(n7806), .A2(n7547), .ZN(n5559) );
  OAI21_X1 U7094 ( .B1(n5563), .B2(n5562), .A(n5561), .ZN(n5564) );
  AND2_X1 U7095 ( .A1(n5564), .A2(n5580), .ZN(n9177) );
  NAND2_X1 U7096 ( .A1(n9177), .A2(n5630), .ZN(n5569) );
  INV_X1 U7097 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9567) );
  NAND2_X1 U7098 ( .A1(n5177), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7099 ( .A1(n5136), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5565) );
  OAI211_X1 U7100 ( .C1(n5616), .C2(n9567), .A(n5566), .B(n5565), .ZN(n5567)
         );
  INV_X1 U7101 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U7102 ( .A1(n5569), .A2(n5568), .ZN(n9029) );
  INV_X1 U7103 ( .A(n9029), .ZN(n9186) );
  INV_X1 U7104 ( .A(n7904), .ZN(n7906) );
  NOR2_X1 U7105 ( .A1(n9172), .A2(n7906), .ZN(n9161) );
  INV_X1 U7106 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7576) );
  INV_X1 U7107 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7572) );
  MUX2_X1 U7108 ( .A(n7576), .B(n7572), .S(n6259), .Z(n5573) );
  INV_X1 U7109 ( .A(SI_26_), .ZN(n9635) );
  NAND2_X1 U7110 ( .A1(n5573), .A2(n9635), .ZN(n5590) );
  INV_X1 U7111 ( .A(n5573), .ZN(n5574) );
  NAND2_X1 U7112 ( .A1(n5574), .A2(SI_26_), .ZN(n5575) );
  NAND2_X1 U7113 ( .A1(n7571), .A2(n7804), .ZN(n5579) );
  OR2_X1 U7114 ( .A1(n7806), .A2(n7572), .ZN(n5578) );
  INV_X1 U7115 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9733) );
  NAND2_X1 U7116 ( .A1(n5580), .A2(n9733), .ZN(n5581) );
  NAND2_X1 U7117 ( .A1(n5614), .A2(n5581), .ZN(n9156) );
  OR2_X1 U7118 ( .A1(n9156), .A2(n5582), .ZN(n5588) );
  INV_X1 U7119 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5585) );
  NAND2_X1 U7120 ( .A1(n6478), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5584) );
  NAND2_X1 U7121 ( .A1(n5136), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5583) );
  OAI211_X1 U7122 ( .C1(n6484), .C2(n5585), .A(n5584), .B(n5583), .ZN(n5586)
         );
  INV_X1 U7123 ( .A(n5586), .ZN(n5587) );
  INV_X1 U7124 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7591) );
  INV_X1 U7125 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5595) );
  MUX2_X1 U7126 ( .A(n7591), .B(n5595), .S(n6259), .Z(n5592) );
  INV_X1 U7127 ( .A(SI_27_), .ZN(n9747) );
  NAND2_X1 U7128 ( .A1(n5592), .A2(n9747), .ZN(n5607) );
  INV_X1 U7129 ( .A(n5592), .ZN(n5593) );
  NAND2_X1 U7130 ( .A1(n5593), .A2(SI_27_), .ZN(n5594) );
  AND2_X1 U7131 ( .A1(n5607), .A2(n5594), .ZN(n5606) );
  NAND2_X1 U7132 ( .A1(n7586), .A2(n7804), .ZN(n5597) );
  OR2_X1 U7133 ( .A1(n7806), .A2(n5595), .ZN(n5596) );
  XNOR2_X1 U7134 ( .A(n5614), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U7135 ( .A1(n9147), .A2(n5630), .ZN(n5603) );
  INV_X1 U7136 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U7137 ( .A1(n5136), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5599) );
  NAND2_X1 U7138 ( .A1(n6478), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5598) );
  OAI211_X1 U7139 ( .C1(n6484), .C2(n5600), .A(n5599), .B(n5598), .ZN(n5601)
         );
  INV_X1 U7140 ( .A(n5601), .ZN(n5602) );
  NAND2_X1 U7141 ( .A1(n5603), .A2(n5602), .ZN(n9028) );
  INV_X1 U7142 ( .A(n7810), .ZN(n8012) );
  INV_X1 U7143 ( .A(n8011), .ZN(n5604) );
  NOR2_X1 U7144 ( .A1(n9139), .A2(n9140), .ZN(n9138) );
  INV_X1 U7145 ( .A(n9122), .ZN(n5622) );
  INV_X1 U7146 ( .A(n5605), .ZN(n5609) );
  INV_X1 U7147 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8887) );
  INV_X1 U7148 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9781) );
  MUX2_X1 U7149 ( .A(n8887), .B(n9781), .S(n6259), .Z(n5626) );
  XNOR2_X1 U7150 ( .A(n5626), .B(SI_28_), .ZN(n5623) );
  NAND2_X1 U7151 ( .A1(n9778), .A2(n7804), .ZN(n5611) );
  OR2_X1 U7152 ( .A1(n7806), .A2(n9781), .ZN(n5610) );
  OAI21_X1 U7153 ( .B1(n5614), .B2(n5613), .A(n5612), .ZN(n5615) );
  NAND2_X1 U7154 ( .A1(n9130), .A2(n5630), .ZN(n5621) );
  INV_X1 U7155 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U7156 ( .A1(n5136), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5618) );
  INV_X1 U7157 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9628) );
  OR2_X1 U7158 ( .A1(n5616), .A2(n9628), .ZN(n5617) );
  OAI211_X1 U7159 ( .C1(n6484), .C2(n9545), .A(n5618), .B(n5617), .ZN(n5619)
         );
  INV_X1 U7160 ( .A(n5619), .ZN(n5620) );
  NAND2_X1 U7161 ( .A1(n5621), .A2(n5620), .ZN(n9137) );
  NAND2_X1 U7162 ( .A1(n9396), .A2(n7727), .ZN(n8014) );
  INV_X1 U7163 ( .A(n9128), .ZN(n7917) );
  NAND2_X1 U7164 ( .A1(n9125), .A2(n8019), .ZN(n5639) );
  INV_X1 U7165 ( .A(SI_28_), .ZN(n5625) );
  INV_X1 U7166 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8106) );
  INV_X1 U7167 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7734) );
  MUX2_X1 U7168 ( .A(n8106), .B(n7734), .S(n7800), .Z(n7592) );
  XNOR2_X1 U7169 ( .A(n7592), .B(SI_29_), .ZN(n5627) );
  NAND2_X1 U7170 ( .A1(n7733), .A2(n7804), .ZN(n5629) );
  OR2_X1 U7171 ( .A1(n7806), .A2(n8106), .ZN(n5628) );
  INV_X1 U7172 ( .A(n5655), .ZN(n5631) );
  NAND2_X1 U7173 ( .A1(n5631), .A2(n5630), .ZN(n5637) );
  INV_X1 U7174 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7175 ( .A1(n6478), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7176 ( .A1(n5136), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5632) );
  OAI211_X1 U7177 ( .C1(n6484), .C2(n5634), .A(n5633), .B(n5632), .ZN(n5635)
         );
  INV_X1 U7178 ( .A(n5635), .ZN(n5636) );
  NAND2_X1 U7179 ( .A1(n5637), .A2(n5636), .ZN(n9027) );
  NAND2_X1 U7180 ( .A1(n9392), .A2(n9123), .ZN(n8088) );
  INV_X1 U7181 ( .A(n8050), .ZN(n5638) );
  XNOR2_X1 U7182 ( .A(n5639), .B(n5638), .ZN(n5651) );
  NAND2_X1 U7183 ( .A1(n8101), .A2(n4392), .ZN(n7936) );
  OR2_X1 U7184 ( .A1(n7727), .A2(n10012), .ZN(n5649) );
  INV_X1 U7185 ( .A(n9874), .ZN(n6380) );
  INV_X1 U7186 ( .A(P1_B_REG_SCAN_IN), .ZN(n5656) );
  NOR2_X1 U7187 ( .A1(n9869), .A2(n5656), .ZN(n5642) );
  NOR2_X1 U7188 ( .A1(n10010), .A2(n5642), .ZN(n9112) );
  INV_X1 U7189 ( .A(n9112), .ZN(n5647) );
  NAND2_X1 U7190 ( .A1(n6478), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5646) );
  INV_X1 U7191 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5643) );
  OR2_X1 U7192 ( .A1(n6484), .A2(n5643), .ZN(n5645) );
  INV_X1 U7193 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9118) );
  OR2_X1 U7194 ( .A1(n6480), .A2(n9118), .ZN(n5644) );
  AND3_X1 U7195 ( .A1(n5646), .A2(n5645), .A3(n5644), .ZN(n7928) );
  OR2_X1 U7196 ( .A1(n5647), .A2(n7928), .ZN(n5648) );
  OAI21_X1 U7197 ( .B1(n9989), .B2(n5651), .A(n5650), .ZN(n5652) );
  INV_X1 U7198 ( .A(n5652), .ZN(n9394) );
  INV_X1 U7199 ( .A(n9241), .ZN(n9237) );
  OR2_X1 U7200 ( .A1(n6747), .A2(n6863), .ZN(n10024) );
  INV_X1 U7201 ( .A(n6703), .ZN(n6808) );
  NAND2_X1 U7202 ( .A1(n6803), .A2(n6808), .ZN(n9973) );
  INV_X1 U7203 ( .A(n9468), .ZN(n7275) );
  INV_X1 U7204 ( .A(n9351), .ZN(n9840) );
  INV_X1 U7205 ( .A(n9340), .ZN(n9832) );
  INV_X1 U7206 ( .A(n9447), .ZN(n9281) );
  INV_X1 U7207 ( .A(n9442), .ZN(n9270) );
  NAND2_X1 U7208 ( .A1(n9277), .A2(n9270), .ZN(n9266) );
  INV_X1 U7209 ( .A(n4392), .ZN(n8054) );
  NAND2_X1 U7210 ( .A1(n7934), .A2(n8054), .ZN(n6862) );
  OR2_X1 U7211 ( .A1(n6862), .A2(n5653), .ZN(n10118) );
  AOI211_X1 U7212 ( .C1(n9392), .C2(n4425), .A(n10118), .B(n9116), .ZN(n9391)
         );
  NAND2_X1 U7213 ( .A1(n9391), .A2(n8092), .ZN(n5654) );
  OAI211_X1 U7214 ( .C1(n5655), .C2(n9994), .A(n9394), .B(n5654), .ZN(n5679)
         );
  AND2_X1 U7215 ( .A1(n5657), .A2(n5656), .ZN(n5661) );
  AND2_X1 U7216 ( .A1(n7549), .A2(P1_B_REG_SCAN_IN), .ZN(n5659) );
  AND2_X1 U7217 ( .A1(n5658), .A2(n5659), .ZN(n5660) );
  OR2_X1 U7218 ( .A1(n10036), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7219 ( .A1(n5658), .A2(n7573), .ZN(n5662) );
  NAND2_X1 U7220 ( .A1(n5663), .A2(n5662), .ZN(n6375) );
  INV_X1 U7221 ( .A(n10072), .ZN(n6379) );
  AND2_X1 U7222 ( .A1(n6375), .A2(n6379), .ZN(n10070) );
  NOR4_X1 U7223 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5667) );
  NOR4_X1 U7224 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5666) );
  NOR4_X1 U7225 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n5665) );
  NOR4_X1 U7226 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n5664) );
  NAND4_X1 U7227 ( .A1(n5667), .A2(n5666), .A3(n5665), .A4(n5664), .ZN(n5673)
         );
  NOR2_X1 U7228 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .ZN(
        n5671) );
  NOR4_X1 U7229 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n5670) );
  NOR4_X1 U7230 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5669) );
  NOR4_X1 U7231 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5668) );
  NAND4_X1 U7232 ( .A1(n5671), .A2(n5670), .A3(n5669), .A4(n5668), .ZN(n5672)
         );
  NOR2_X1 U7233 ( .A1(n5673), .A2(n5672), .ZN(n5674) );
  NOR2_X1 U7234 ( .A1(n10036), .A2(n5674), .ZN(n6376) );
  AND2_X1 U7235 ( .A1(n8093), .A2(n8092), .ZN(n6861) );
  OR2_X1 U7236 ( .A1(n7936), .A2(n6861), .ZN(n6574) );
  INV_X1 U7237 ( .A(n6574), .ZN(n5675) );
  NOR2_X1 U7238 ( .A1(n6376), .A2(n5675), .ZN(n5676) );
  NAND2_X1 U7239 ( .A1(n7573), .A2(n7549), .ZN(n5677) );
  NAND2_X1 U7240 ( .A1(n5678), .A2(n5677), .ZN(n6524) );
  INV_X1 U7241 ( .A(n6524), .ZN(n6276) );
  NAND2_X1 U7242 ( .A1(n6525), .A2(n6276), .ZN(n6804) );
  AND2_X2 U7243 ( .A1(n6804), .A2(n9994), .ZN(n10021) );
  NAND2_X1 U7244 ( .A1(n5679), .A2(n9321), .ZN(n5723) );
  NAND2_X1 U7245 ( .A1(n6388), .A2(n6863), .ZN(n6730) );
  NAND2_X1 U7246 ( .A1(n6737), .A2(n6730), .ZN(n5682) );
  OR2_X1 U7247 ( .A1(n9039), .A2(n6747), .ZN(n5681) );
  NAND2_X1 U7248 ( .A1(n5682), .A2(n5681), .ZN(n10013) );
  INV_X1 U7249 ( .A(n10014), .ZN(n5683) );
  NAND2_X1 U7250 ( .A1(n10013), .A2(n5683), .ZN(n5685) );
  OR2_X1 U7251 ( .A1(n6542), .A2(n10023), .ZN(n5684) );
  AND2_X1 U7252 ( .A1(n8063), .A2(n9981), .ZN(n8030) );
  INV_X1 U7253 ( .A(n8030), .ZN(n6922) );
  NAND2_X1 U7254 ( .A1(n6921), .A2(n6922), .ZN(n5687) );
  OR2_X1 U7255 ( .A1(n10009), .A2(n6562), .ZN(n5686) );
  NAND2_X1 U7256 ( .A1(n5687), .A2(n5686), .ZN(n9980) );
  NAND2_X1 U7257 ( .A1(n8067), .A2(n7945), .ZN(n9984) );
  NAND2_X1 U7258 ( .A1(n9980), .A2(n9984), .ZN(n5689) );
  OR2_X1 U7259 ( .A1(n9038), .A2(n9998), .ZN(n5688) );
  NAND2_X1 U7260 ( .A1(n5689), .A2(n5688), .ZN(n7110) );
  INV_X1 U7261 ( .A(n7110), .ZN(n5691) );
  INV_X1 U7262 ( .A(n5690), .ZN(n7950) );
  NAND2_X1 U7263 ( .A1(n7950), .A2(n7822), .ZN(n8031) );
  INV_X1 U7264 ( .A(n8031), .ZN(n7109) );
  NAND2_X1 U7265 ( .A1(n5691), .A2(n8031), .ZN(n10102) );
  NAND2_X1 U7266 ( .A1(n9986), .A2(n7102), .ZN(n5692) );
  NAND2_X1 U7267 ( .A1(n10102), .A2(n5692), .ZN(n6784) );
  AND2_X1 U7268 ( .A1(n8074), .A2(n7827), .ZN(n7820) );
  OR2_X1 U7269 ( .A1(n9037), .A2(n7095), .ZN(n5693) );
  INV_X1 U7270 ( .A(n8034), .ZN(n6812) );
  NOR2_X1 U7271 ( .A1(n6703), .A2(n9036), .ZN(n5694) );
  AOI21_X1 U7272 ( .B1(n6811), .B2(n6812), .A(n5694), .ZN(n9961) );
  NAND2_X1 U7273 ( .A1(n9961), .A2(n9963), .ZN(n9960) );
  NAND2_X1 U7274 ( .A1(n9968), .A2(n9035), .ZN(n5695) );
  NAND2_X1 U7275 ( .A1(n9960), .A2(n5695), .ZN(n7012) );
  OR2_X1 U7276 ( .A1(n7195), .A2(n9034), .ZN(n5696) );
  NAND2_X1 U7277 ( .A1(n7012), .A2(n5696), .ZN(n5698) );
  NAND2_X1 U7278 ( .A1(n7195), .A2(n9034), .ZN(n5697) );
  OR2_X1 U7279 ( .A1(n7326), .A2(n9033), .ZN(n5699) );
  NAND2_X1 U7280 ( .A1(n7267), .A2(n8040), .ZN(n7266) );
  NAND2_X1 U7281 ( .A1(n7266), .A2(n9032), .ZN(n5700) );
  NAND2_X1 U7282 ( .A1(n5700), .A2(n4402), .ZN(n7430) );
  NAND2_X1 U7283 ( .A1(n5701), .A2(n7976), .ZN(n9369) );
  NAND2_X1 U7284 ( .A1(n9457), .A2(n9030), .ZN(n5705) );
  INV_X1 U7285 ( .A(n5705), .ZN(n5702) );
  AND2_X1 U7286 ( .A1(n9369), .A2(n5704), .ZN(n5703) );
  NAND2_X1 U7287 ( .A1(n7430), .A2(n5703), .ZN(n5709) );
  INV_X1 U7288 ( .A(n5704), .ZN(n5707) );
  NAND2_X1 U7289 ( .A1(n9464), .A2(n9031), .ZN(n9370) );
  AND2_X1 U7290 ( .A1(n9370), .A2(n5705), .ZN(n5706) );
  OR2_X1 U7291 ( .A1(n9351), .A2(n9327), .ZN(n5710) );
  INV_X1 U7292 ( .A(n9318), .ZN(n9826) );
  NAND2_X1 U7293 ( .A1(n9304), .A2(n5038), .ZN(n9290) );
  NAND2_X1 U7294 ( .A1(n4723), .A2(n5711), .ZN(n5713) );
  NAND2_X1 U7295 ( .A1(n9452), .A2(n9310), .ZN(n7862) );
  INV_X1 U7296 ( .A(n7862), .ZN(n5712) );
  INV_X1 U7297 ( .A(n9439), .ZN(n9255) );
  NAND2_X1 U7298 ( .A1(n9427), .A2(n9228), .ZN(n5715) );
  INV_X1 U7299 ( .A(n9427), .ZN(n5714) );
  AOI21_X1 U7300 ( .B1(n9176), .B2(n9159), .A(n9154), .ZN(n5717) );
  NAND2_X1 U7301 ( .A1(n5719), .A2(n8093), .ZN(n6383) );
  OR2_X1 U7302 ( .A1(n6734), .A2(n6383), .ZN(n8099) );
  INV_X1 U7303 ( .A(n8099), .ZN(n6527) );
  OR2_X1 U7304 ( .A1(n6862), .A2(n8093), .ZN(n6377) );
  AOI22_X1 U7305 ( .A1(n9392), .A2(n9350), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n9387), .ZN(n5720) );
  NAND2_X1 U7306 ( .A1(n5723), .A2(n5722), .ZN(P1_U3355) );
  NOR2_X1 U7307 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5730) );
  NOR2_X1 U7308 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5729) );
  INV_X1 U7309 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5728) );
  NAND4_X1 U7310 ( .A1(n5761), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n5733)
         );
  NAND2_X1 U7311 ( .A1(n6009), .A2(n6121), .ZN(n6124) );
  INV_X1 U7312 ( .A(n6124), .ZN(n5731) );
  NAND3_X1 U7313 ( .A1(n5731), .A2(n5994), .A3(n5982), .ZN(n5732) );
  NOR2_X1 U7314 ( .A1(n5733), .A2(n5732), .ZN(n5734) );
  XNOR2_X2 U7315 ( .A(n5737), .B(n5735), .ZN(n7589) );
  NAND2_X1 U7316 ( .A1(n7417), .A2(n8249), .ZN(n5739) );
  OR2_X1 U7317 ( .A1(n8250), .A2(n7416), .ZN(n5738) );
  NAND2_X1 U7318 ( .A1(n5880), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5907) );
  INV_X1 U7319 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5922) );
  INV_X1 U7320 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n9683) );
  INV_X1 U7321 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5765) );
  INV_X1 U7322 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8536) );
  AND2_X1 U7323 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5744) );
  INV_X1 U7324 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8189) );
  INV_X1 U7325 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9715) );
  NAND2_X1 U7326 ( .A1(n6043), .A2(n9715), .ZN(n5747) );
  NAND2_X1 U7327 ( .A1(n6052), .A2(n5747), .ZN(n8620) );
  OR2_X2 U7328 ( .A1(n5751), .A2(n6159), .ZN(n5749) );
  INV_X1 U7329 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5750) );
  XNOR2_X2 U7330 ( .A(n5749), .B(n5750), .ZN(n5754) );
  OR2_X1 U7331 ( .A1(n8620), .A2(n6110), .ZN(n5759) );
  NAND2_X4 U7332 ( .A1(n8881), .A2(n5752), .ZN(n6290) );
  INV_X1 U7333 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9569) );
  INV_X2 U7334 ( .A(n5823), .ZN(n6284) );
  NAND2_X1 U7335 ( .A1(n6284), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5756) );
  INV_X1 U7336 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9728) );
  OR2_X1 U7337 ( .A1(n6286), .A2(n9728), .ZN(n5755) );
  OAI211_X1 U7338 ( .C1(n6290), .C2(n9569), .A(n5756), .B(n5755), .ZN(n5757)
         );
  INV_X1 U7339 ( .A(n5757), .ZN(n5758) );
  NAND2_X1 U7340 ( .A1(n5759), .A2(n5758), .ZN(n8457) );
  NAND2_X1 U7341 ( .A1(n6625), .A2(n8249), .ZN(n5764) );
  XNOR2_X1 U7342 ( .A(n5762), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7747) );
  AOI22_X1 U7343 ( .A1(n6013), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6012), .B2(
        n7747), .ZN(n5763) );
  INV_X1 U7344 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9719) );
  OR2_X1 U7345 ( .A1(n6286), .A2(n9719), .ZN(n5770) );
  INV_X1 U7346 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8756) );
  OR2_X1 U7347 ( .A1(n4390), .A2(n8756), .ZN(n5769) );
  NAND2_X1 U7348 ( .A1(n5976), .A2(n5765), .ZN(n5766) );
  NAND2_X1 U7349 ( .A1(n5986), .A2(n5766), .ZN(n8755) );
  OR2_X1 U7350 ( .A1(n6077), .A2(n8755), .ZN(n5768) );
  INV_X1 U7351 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7509) );
  OR2_X1 U7352 ( .A1(n6114), .A2(n7509), .ZN(n5767) );
  NAND4_X1 U7353 ( .A1(n5770), .A2(n5769), .A3(n5768), .A4(n5767), .ZN(n8720)
         );
  INV_X1 U7354 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6403) );
  OR2_X2 U7355 ( .A1(n6290), .A2(n6403), .ZN(n5775) );
  INV_X1 U7356 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5771) );
  OR2_X1 U7357 ( .A1(n5823), .A2(n5771), .ZN(n5774) );
  INV_X1 U7358 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5772) );
  OR2_X1 U7359 ( .A1(n6286), .A2(n5772), .ZN(n5773) );
  INV_X1 U7360 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6256) );
  OR2_X1 U7361 ( .A1(n5817), .A2(n6256), .ZN(n5778) );
  NAND2_X1 U7362 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5777) );
  INV_X1 U7363 ( .A(n9791), .ZN(n6415) );
  NAND3_X2 U7364 ( .A1(n5779), .A2(n5778), .A3(n5041), .ZN(n10215) );
  INV_X2 U7365 ( .A(n10215), .ZN(n10246) );
  NAND2_X1 U7366 ( .A1(n5787), .A2(n10246), .ZN(n8276) );
  NAND2_X1 U7367 ( .A1(n6284), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5785) );
  INV_X1 U7368 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n6901) );
  OR2_X1 U7369 ( .A1(n5791), .A2(n6901), .ZN(n5784) );
  INV_X1 U7370 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5780) );
  OR2_X1 U7371 ( .A1(n6290), .A2(n5780), .ZN(n5783) );
  INV_X1 U7372 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5781) );
  OR2_X1 U7373 ( .A1(n6286), .A2(n5781), .ZN(n5782) );
  NAND2_X1 U7374 ( .A1(n7800), .A2(SI_0_), .ZN(n5786) );
  XNOR2_X1 U7375 ( .A(n5786), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n8889) );
  NAND2_X1 U7376 ( .A1(n10206), .A2(n10214), .ZN(n10204) );
  NAND2_X1 U7377 ( .A1(n8401), .A2(n10204), .ZN(n5789) );
  OR2_X1 U7378 ( .A1(n5787), .A2(n10215), .ZN(n5788) );
  NAND2_X1 U7379 ( .A1(n5789), .A2(n5788), .ZN(n6935) );
  INV_X1 U7380 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n5790) );
  INV_X1 U7381 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6941) );
  OR2_X1 U7382 ( .A1(n5791), .A2(n6941), .ZN(n5796) );
  INV_X1 U7383 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5792) );
  OR2_X1 U7384 ( .A1(n6286), .A2(n5792), .ZN(n5795) );
  INV_X1 U7385 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n5793) );
  OR2_X1 U7386 ( .A1(n5823), .A2(n5793), .ZN(n5794) );
  NAND2_X2 U7387 ( .A1(n5797), .A2(n4416), .ZN(n5806) );
  INV_X1 U7388 ( .A(n5798), .ZN(n5799) );
  NAND2_X1 U7389 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n5799), .ZN(n5800) );
  MUX2_X1 U7390 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5800), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n5802) );
  INV_X1 U7391 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5801) );
  NAND2_X1 U7392 ( .A1(n5801), .A2(n5798), .ZN(n5815) );
  NAND2_X1 U7393 ( .A1(n5802), .A2(n5815), .ZN(n6414) );
  OR2_X1 U7394 ( .A1(n5817), .A2(n6257), .ZN(n5803) );
  INV_X1 U7395 ( .A(n6200), .ZN(n10251) );
  NAND2_X1 U7396 ( .A1(n5805), .A2(n6200), .ZN(n8278) );
  NAND2_X1 U7397 ( .A1(n6935), .A2(n8402), .ZN(n5808) );
  OR2_X1 U7398 ( .A1(n5806), .A2(n6200), .ZN(n5807) );
  NAND2_X1 U7399 ( .A1(n5808), .A2(n5807), .ZN(n10194) );
  NAND2_X1 U7400 ( .A1(n5921), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5814) );
  OR2_X1 U7401 ( .A1(n6077), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5813) );
  INV_X1 U7402 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5809) );
  OR2_X1 U7403 ( .A1(n4390), .A2(n5809), .ZN(n5812) );
  INV_X1 U7404 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5810) );
  OR2_X1 U7405 ( .A1(n6286), .A2(n5810), .ZN(n5811) );
  NAND2_X1 U7406 ( .A1(n5815), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5816) );
  XNOR2_X1 U7407 ( .A(n5816), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6413) );
  INV_X1 U7408 ( .A(n6413), .ZN(n6476) );
  OR2_X1 U7409 ( .A1(n5817), .A2(n6258), .ZN(n5818) );
  NAND2_X1 U7410 ( .A1(n10194), .A2(n10195), .ZN(n5821) );
  OR2_X1 U7411 ( .A1(n8468), .A2(n8290), .ZN(n5820) );
  NAND2_X1 U7412 ( .A1(n5821), .A2(n5820), .ZN(n10178) );
  NAND2_X1 U7413 ( .A1(n6111), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5827) );
  INV_X1 U7414 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5822) );
  OR2_X1 U7415 ( .A1(n4390), .A2(n5822), .ZN(n5826) );
  XNOR2_X1 U7416 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n10180) );
  OR2_X1 U7417 ( .A1(n6110), .A2(n10180), .ZN(n5825) );
  INV_X1 U7418 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6406) );
  OR2_X1 U7419 ( .A1(n6290), .A2(n6406), .ZN(n5824) );
  NAND4_X1 U7420 ( .A1(n5827), .A2(n5826), .A3(n5825), .A4(n5824), .ZN(n10191)
         );
  OR2_X1 U7421 ( .A1(n5828), .A2(n6159), .ZN(n5829) );
  XNOR2_X1 U7422 ( .A(n5829), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6435) );
  INV_X1 U7423 ( .A(n6435), .ZN(n6424) );
  OR2_X1 U7424 ( .A1(n5845), .A2(n6268), .ZN(n5831) );
  OR2_X1 U7425 ( .A1(n8250), .A2(n9744), .ZN(n5830) );
  OAI211_X1 U7426 ( .C1(n6401), .C2(n6424), .A(n5831), .B(n5830), .ZN(n10182)
         );
  OR2_X1 U7427 ( .A1(n10191), .A2(n10262), .ZN(n8267) );
  NAND2_X1 U7428 ( .A1(n10191), .A2(n10262), .ZN(n6950) );
  NAND2_X1 U7429 ( .A1(n8267), .A2(n6950), .ZN(n10179) );
  NAND2_X1 U7430 ( .A1(n10178), .A2(n10179), .ZN(n5833) );
  OR2_X1 U7431 ( .A1(n10191), .A2(n10182), .ZN(n5832) );
  NAND2_X1 U7432 ( .A1(n6111), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5842) );
  INV_X1 U7433 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6959) );
  OR2_X1 U7434 ( .A1(n4390), .A2(n6959), .ZN(n5841) );
  INV_X1 U7435 ( .A(n5834), .ZN(n5852) );
  INV_X1 U7436 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U7437 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5835) );
  NAND2_X1 U7438 ( .A1(n5836), .A2(n5835), .ZN(n5837) );
  NAND2_X1 U7439 ( .A1(n5852), .A2(n5837), .ZN(n6958) );
  OR2_X1 U7440 ( .A1(n6110), .A2(n6958), .ZN(n5840) );
  INV_X1 U7441 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5838) );
  OR2_X1 U7442 ( .A1(n6290), .A2(n5838), .ZN(n5839) );
  NAND4_X1 U7443 ( .A1(n5842), .A2(n5841), .A3(n5840), .A4(n5839), .ZN(n8467)
         );
  NAND2_X1 U7444 ( .A1(n5843), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5844) );
  XNOR2_X1 U7445 ( .A(n5844), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6434) );
  INV_X1 U7446 ( .A(n6434), .ZN(n6465) );
  OR2_X1 U7447 ( .A1(n8250), .A2(n6265), .ZN(n5846) );
  NOR2_X1 U7448 ( .A1(n8467), .A2(n6192), .ZN(n5848) );
  NAND2_X1 U7449 ( .A1(n8467), .A2(n6192), .ZN(n5847) );
  NAND2_X1 U7450 ( .A1(n6270), .A2(n8249), .ZN(n5850) );
  NOR2_X1 U7451 ( .A1(n5843), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7452 ( .A1(n5877), .A2(n6159), .ZN(n5870) );
  XNOR2_X1 U7453 ( .A(n5870), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6433) );
  AOI22_X1 U7454 ( .A1(n6013), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6012), .B2(
        n6433), .ZN(n5849) );
  NAND2_X1 U7455 ( .A1(n6111), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5857) );
  INV_X1 U7456 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6973) );
  OR2_X1 U7457 ( .A1(n4390), .A2(n6973), .ZN(n5856) );
  INV_X1 U7458 ( .A(n5851), .ZN(n5862) );
  INV_X1 U7459 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U7460 ( .A1(n5852), .A2(n6443), .ZN(n5853) );
  NAND2_X1 U7461 ( .A1(n5862), .A2(n5853), .ZN(n6972) );
  OR2_X1 U7462 ( .A1(n6077), .A2(n6972), .ZN(n5855) );
  INV_X1 U7463 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6427) );
  OR2_X1 U7464 ( .A1(n6114), .A2(n6427), .ZN(n5854) );
  NAND4_X1 U7465 ( .A1(n5857), .A2(n5856), .A3(n5855), .A4(n5854), .ZN(n8466)
         );
  NAND2_X1 U7466 ( .A1(n10275), .A2(n8466), .ZN(n8294) );
  NAND2_X1 U7467 ( .A1(n6968), .A2(n8407), .ZN(n5859) );
  NAND2_X1 U7468 ( .A1(n8466), .A2(n6975), .ZN(n5858) );
  NAND2_X1 U7469 ( .A1(n6111), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5868) );
  INV_X1 U7470 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5860) );
  OR2_X1 U7471 ( .A1(n4390), .A2(n5860), .ZN(n5867) );
  INV_X1 U7472 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U7473 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  NAND2_X1 U7474 ( .A1(n5881), .A2(n5863), .ZN(n6779) );
  OR2_X1 U7475 ( .A1(n6077), .A2(n6779), .ZN(n5866) );
  INV_X1 U7476 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n5864) );
  OR2_X1 U7477 ( .A1(n6290), .A2(n5864), .ZN(n5865) );
  NAND4_X1 U7478 ( .A1(n5868), .A2(n5867), .A3(n5866), .A4(n5865), .ZN(n8465)
         );
  INV_X1 U7479 ( .A(n8465), .ZN(n5875) );
  NAND2_X1 U7480 ( .A1(n6273), .A2(n8249), .ZN(n5874) );
  INV_X1 U7481 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U7482 ( .A1(n5870), .A2(n5869), .ZN(n5871) );
  NAND2_X1 U7483 ( .A1(n5871), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5872) );
  XNOR2_X1 U7484 ( .A(n5872), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6516) );
  AOI22_X1 U7485 ( .A1(n6013), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6012), .B2(
        n6516), .ZN(n5873) );
  NAND2_X1 U7486 ( .A1(n5874), .A2(n5873), .ZN(n6771) );
  OR2_X1 U7487 ( .A1(n5875), .A2(n6771), .ZN(n6980) );
  NAND2_X1 U7488 ( .A1(n5875), .A2(n6771), .ZN(n8306) );
  NOR2_X1 U7489 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5876) );
  NAND2_X1 U7490 ( .A1(n5877), .A2(n5876), .ZN(n5888) );
  NAND2_X1 U7491 ( .A1(n5888), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5878) );
  XNOR2_X1 U7492 ( .A(n5878), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6662) );
  AOI22_X1 U7493 ( .A1(n6013), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6012), .B2(
        n6662), .ZN(n5879) );
  NAND2_X1 U7494 ( .A1(n6111), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5886) );
  INV_X1 U7495 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6990) );
  OR2_X1 U7496 ( .A1(n4390), .A2(n6990), .ZN(n5885) );
  INV_X1 U7497 ( .A(n5880), .ZN(n5893) );
  NAND2_X1 U7498 ( .A1(n5881), .A2(n6509), .ZN(n5882) );
  NAND2_X1 U7499 ( .A1(n5893), .A2(n5882), .ZN(n6989) );
  OR2_X1 U7500 ( .A1(n6110), .A2(n6989), .ZN(n5884) );
  INV_X1 U7501 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6511) );
  OR2_X1 U7502 ( .A1(n6290), .A2(n6511), .ZN(n5883) );
  NAND4_X1 U7503 ( .A1(n5886), .A2(n5885), .A3(n5884), .A4(n5883), .ZN(n8464)
         );
  INV_X1 U7504 ( .A(n8464), .ZN(n7232) );
  OR2_X1 U7505 ( .A1(n6992), .A2(n7232), .ZN(n8309) );
  NAND2_X1 U7506 ( .A1(n6992), .A2(n7232), .ZN(n8300) );
  NAND2_X1 U7507 ( .A1(n6992), .A2(n8464), .ZN(n5887) );
  NAND2_X1 U7508 ( .A1(n6985), .A2(n5887), .ZN(n7235) );
  INV_X1 U7509 ( .A(n7235), .ZN(n5901) );
  NAND2_X1 U7510 ( .A1(n6292), .A2(n8249), .ZN(n5891) );
  NAND2_X1 U7511 ( .A1(n5903), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5889) );
  XNOR2_X1 U7512 ( .A(n5889), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8475) );
  AOI22_X1 U7513 ( .A1(n6013), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6012), .B2(
        n8475), .ZN(n5890) );
  NAND2_X1 U7514 ( .A1(n6111), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5898) );
  OR2_X1 U7515 ( .A1(n4390), .A2(n6653), .ZN(n5897) );
  INV_X1 U7516 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7517 ( .A1(n5893), .A2(n5892), .ZN(n5894) );
  NAND2_X1 U7518 ( .A1(n5907), .A2(n5894), .ZN(n7070) );
  OR2_X1 U7519 ( .A1(n6077), .A2(n7070), .ZN(n5896) );
  INV_X1 U7520 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6663) );
  OR2_X1 U7521 ( .A1(n6114), .A2(n6663), .ZN(n5895) );
  NAND4_X1 U7522 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n8463)
         );
  INV_X1 U7523 ( .A(n8463), .ZN(n5899) );
  OR2_X1 U7524 ( .A1(n7421), .A2(n5899), .ZN(n8310) );
  NAND2_X1 U7525 ( .A1(n7421), .A2(n5899), .ZN(n8314) );
  NAND2_X1 U7526 ( .A1(n5901), .A2(n5900), .ZN(n7233) );
  OR2_X1 U7527 ( .A1(n7421), .A2(n8463), .ZN(n5902) );
  NAND2_X1 U7528 ( .A1(n7233), .A2(n5902), .ZN(n7176) );
  INV_X1 U7529 ( .A(n7176), .ZN(n5915) );
  NAND2_X1 U7530 ( .A1(n6300), .A2(n8249), .ZN(n5906) );
  NAND2_X1 U7531 ( .A1(n5917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5904) );
  XNOR2_X1 U7532 ( .A(n5904), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8489) );
  AOI22_X1 U7533 ( .A1(n6013), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6012), .B2(
        n8489), .ZN(n5905) );
  NAND2_X1 U7534 ( .A1(n6111), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5913) );
  INV_X1 U7535 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7187) );
  OR2_X1 U7536 ( .A1(n4390), .A2(n7187), .ZN(n5912) );
  NAND2_X1 U7537 ( .A1(n5907), .A2(n8487), .ZN(n5908) );
  NAND2_X1 U7538 ( .A1(n5923), .A2(n5908), .ZN(n7257) );
  OR2_X1 U7539 ( .A1(n6077), .A2(n7257), .ZN(n5911) );
  INV_X1 U7540 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n5909) );
  OR2_X1 U7541 ( .A1(n6290), .A2(n5909), .ZN(n5910) );
  NAND4_X1 U7542 ( .A1(n5913), .A2(n5912), .A3(n5911), .A4(n5910), .ZN(n8462)
         );
  INV_X1 U7543 ( .A(n8462), .ZN(n7231) );
  NAND2_X1 U7544 ( .A1(n7264), .A2(n7231), .ZN(n8304) );
  NAND2_X1 U7545 ( .A1(n7264), .A2(n8462), .ZN(n5916) );
  NAND2_X1 U7546 ( .A1(n6315), .A2(n8249), .ZN(n5920) );
  OAI21_X1 U7547 ( .B1(n5917), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5918) );
  XNOR2_X1 U7548 ( .A(n5918), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7134) );
  AOI22_X1 U7549 ( .A1(n6013), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6012), .B2(
        n7134), .ZN(n5919) );
  NAND2_X1 U7550 ( .A1(n5921), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5930) );
  NAND2_X1 U7551 ( .A1(n5923), .A2(n5922), .ZN(n5924) );
  NAND2_X1 U7552 ( .A1(n5937), .A2(n5924), .ZN(n7224) );
  OR2_X1 U7553 ( .A1(n6110), .A2(n7224), .ZN(n5929) );
  INV_X1 U7554 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5925) );
  OR2_X1 U7555 ( .A1(n4390), .A2(n5925), .ZN(n5928) );
  INV_X1 U7556 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5926) );
  OR2_X1 U7557 ( .A1(n6286), .A2(n5926), .ZN(n5927) );
  NAND4_X1 U7558 ( .A1(n5930), .A2(n5929), .A3(n5928), .A4(n5927), .ZN(n8461)
         );
  INV_X1 U7559 ( .A(n8461), .ZN(n5931) );
  NAND2_X1 U7560 ( .A1(n7367), .A2(n5931), .ZN(n8321) );
  NAND2_X1 U7561 ( .A1(n8317), .A2(n8321), .ZN(n8414) );
  NAND2_X1 U7562 ( .A1(n6353), .A2(n8249), .ZN(n5935) );
  NAND2_X1 U7563 ( .A1(n5932), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5933) );
  XNOR2_X1 U7564 ( .A(n5933), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8502) );
  AOI22_X1 U7565 ( .A1(n6013), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6012), .B2(
        n8502), .ZN(n5934) );
  NAND2_X1 U7566 ( .A1(n6111), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5942) );
  INV_X1 U7567 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7320) );
  OR2_X1 U7568 ( .A1(n4390), .A2(n7320), .ZN(n5941) );
  INV_X1 U7569 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n5936) );
  OR2_X1 U7570 ( .A1(n6290), .A2(n5936), .ZN(n5940) );
  INV_X1 U7571 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8500) );
  NAND2_X1 U7572 ( .A1(n5937), .A2(n8500), .ZN(n5938) );
  NAND2_X1 U7573 ( .A1(n5951), .A2(n5938), .ZN(n7319) );
  OR2_X1 U7574 ( .A1(n6077), .A2(n7319), .ZN(n5939) );
  NAND4_X1 U7575 ( .A1(n5942), .A2(n5941), .A3(n5940), .A4(n5939), .ZN(n8460)
         );
  INV_X1 U7576 ( .A(n8460), .ZN(n7155) );
  OR2_X1 U7577 ( .A1(n10295), .A2(n7155), .ZN(n8318) );
  NAND2_X1 U7578 ( .A1(n10295), .A2(n7155), .ZN(n8322) );
  NAND2_X1 U7579 ( .A1(n6396), .A2(n8249), .ZN(n5948) );
  NOR2_X1 U7580 ( .A1(n4478), .A2(n6159), .ZN(n5943) );
  MUX2_X1 U7581 ( .A(n6159), .B(n5943), .S(P2_IR_REG_13__SCAN_IN), .Z(n5944)
         );
  INV_X1 U7582 ( .A(n5944), .ZN(n5946) );
  INV_X1 U7583 ( .A(n5760), .ZN(n5945) );
  AND2_X1 U7584 ( .A1(n5946), .A2(n5945), .ZN(n10167) );
  AOI22_X1 U7585 ( .A1(n6013), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6012), .B2(
        n10167), .ZN(n5947) );
  NAND2_X1 U7586 ( .A1(n6111), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5956) );
  INV_X1 U7587 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7497) );
  OR2_X1 U7588 ( .A1(n4390), .A2(n7497), .ZN(n5955) );
  INV_X1 U7589 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5949) );
  OR2_X1 U7590 ( .A1(n6114), .A2(n5949), .ZN(n5954) );
  INV_X1 U7591 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7592 ( .A1(n5951), .A2(n5950), .ZN(n5952) );
  NAND2_X1 U7593 ( .A1(n5960), .A2(n5952), .ZN(n7496) );
  OR2_X1 U7594 ( .A1(n6110), .A2(n7496), .ZN(n5953) );
  NAND4_X1 U7595 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n8459)
         );
  INV_X1 U7596 ( .A(n8459), .ZN(n7304) );
  OR2_X1 U7597 ( .A1(n8850), .A2(n7304), .ZN(n8329) );
  NAND2_X1 U7598 ( .A1(n8850), .A2(n7304), .ZN(n8330) );
  NAND2_X1 U7599 ( .A1(n8850), .A2(n8459), .ZN(n5957) );
  NAND2_X1 U7600 ( .A1(n7491), .A2(n5957), .ZN(n7476) );
  NAND2_X1 U7601 ( .A1(n6488), .A2(n8249), .ZN(n5959) );
  OR2_X1 U7602 ( .A1(n5760), .A2(n6159), .ZN(n5967) );
  XNOR2_X1 U7603 ( .A(n5967), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7515) );
  AOI22_X1 U7604 ( .A1(n6013), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6012), .B2(
        n7515), .ZN(n5958) );
  NAND2_X1 U7605 ( .A1(n6111), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5965) );
  NAND2_X1 U7606 ( .A1(n5960), .A2(n9683), .ZN(n5961) );
  NAND2_X1 U7607 ( .A1(n5974), .A2(n5961), .ZN(n7482) );
  OR2_X1 U7608 ( .A1(n6110), .A2(n7482), .ZN(n5964) );
  OR2_X1 U7609 ( .A1(n4390), .A2(n7130), .ZN(n5963) );
  INV_X1 U7610 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7139) );
  OR2_X1 U7611 ( .A1(n6290), .A2(n7139), .ZN(n5962) );
  NAND4_X1 U7612 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(n8458)
         );
  INV_X1 U7613 ( .A(n8458), .ZN(n7450) );
  NAND2_X1 U7614 ( .A1(n7484), .A2(n7450), .ZN(n8332) );
  NAND2_X1 U7615 ( .A1(n6615), .A2(n8249), .ZN(n5971) );
  INV_X1 U7616 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5966) );
  NAND2_X1 U7617 ( .A1(n5967), .A2(n5966), .ZN(n5968) );
  NAND2_X1 U7618 ( .A1(n5968), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5969) );
  XNOR2_X1 U7619 ( .A(n5969), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8515) );
  AOI22_X1 U7620 ( .A1(n6013), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6012), .B2(
        n8515), .ZN(n5970) );
  NAND2_X1 U7621 ( .A1(n6284), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5981) );
  INV_X1 U7622 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5972) );
  OR2_X1 U7623 ( .A1(n6286), .A2(n5972), .ZN(n5980) );
  INV_X1 U7624 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7625 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U7626 ( .A1(n5976), .A2(n5975), .ZN(n7558) );
  OR2_X1 U7627 ( .A1(n6077), .A2(n7558), .ZN(n5979) );
  INV_X1 U7628 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5977) );
  OR2_X1 U7629 ( .A1(n6290), .A2(n5977), .ZN(n5978) );
  NAND4_X1 U7630 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n8743)
         );
  INV_X1 U7631 ( .A(n8743), .ZN(n8336) );
  XNOR2_X1 U7632 ( .A(n8844), .B(n8336), .ZN(n7554) );
  NAND2_X1 U7633 ( .A1(n7555), .A2(n7554), .ZN(n7553) );
  OR2_X1 U7634 ( .A1(n8844), .A2(n8743), .ZN(n8337) );
  NAND2_X1 U7635 ( .A1(n7553), .A2(n8337), .ZN(n8738) );
  INV_X1 U7636 ( .A(n8720), .ZN(n7566) );
  NAND2_X1 U7637 ( .A1(n8836), .A2(n7566), .ZN(n8340) );
  NAND2_X1 U7638 ( .A1(n6629), .A2(n8249), .ZN(n5985) );
  NAND2_X1 U7639 ( .A1(n5993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5983) );
  XNOR2_X1 U7640 ( .A(n5983), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7748) );
  AOI22_X1 U7641 ( .A1(n6013), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6012), .B2(
        n7748), .ZN(n5984) );
  NAND2_X1 U7642 ( .A1(n6111), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5992) );
  INV_X1 U7643 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8732) );
  OR2_X1 U7644 ( .A1(n4390), .A2(n8732), .ZN(n5991) );
  INV_X1 U7645 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8525) );
  NAND2_X1 U7646 ( .A1(n5986), .A2(n8525), .ZN(n5987) );
  NAND2_X1 U7647 ( .A1(n6000), .A2(n5987), .ZN(n8731) );
  OR2_X1 U7648 ( .A1(n6110), .A2(n8731), .ZN(n5990) );
  INV_X1 U7649 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n5988) );
  OR2_X1 U7650 ( .A1(n6290), .A2(n5988), .ZN(n5989) );
  NAND4_X1 U7651 ( .A1(n5992), .A2(n5991), .A3(n5990), .A4(n5989), .ZN(n8742)
         );
  INV_X1 U7652 ( .A(n8742), .ZN(n7581) );
  NAND2_X1 U7653 ( .A1(n8831), .A2(n7581), .ZN(n8262) );
  NAND2_X1 U7654 ( .A1(n6750), .A2(n8249), .ZN(n5997) );
  NAND2_X1 U7655 ( .A1(n6123), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7656 ( .A(n6007), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8538) );
  AOI22_X1 U7657 ( .A1(n6013), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6012), .B2(
        n8538), .ZN(n5996) );
  INV_X1 U7658 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U7659 ( .A1(n6111), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5998) );
  OAI21_X1 U7660 ( .B1(n4390), .B2(n5999), .A(n5998), .ZN(n6004) );
  NAND2_X1 U7661 ( .A1(n6000), .A2(n8536), .ZN(n6001) );
  NAND2_X1 U7662 ( .A1(n6027), .A2(n6001), .ZN(n8697) );
  INV_X1 U7663 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n7745) );
  OR2_X1 U7664 ( .A1(n6290), .A2(n7745), .ZN(n6002) );
  OAI21_X1 U7665 ( .B1(n8697), .B2(n6077), .A(n6002), .ZN(n6003) );
  OR2_X1 U7666 ( .A1(n6004), .A2(n6003), .ZN(n8721) );
  NAND2_X1 U7667 ( .A1(n8826), .A2(n8721), .ZN(n6006) );
  INV_X1 U7668 ( .A(n8721), .ZN(n8683) );
  INV_X1 U7669 ( .A(n8826), .ZN(n8701) );
  NAND2_X1 U7670 ( .A1(n6869), .A2(n8249), .ZN(n6015) );
  NAND2_X1 U7671 ( .A1(n6008), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n6011) );
  INV_X1 U7672 ( .A(n6008), .ZN(n6010) );
  NAND2_X1 U7673 ( .A1(n6010), .A2(n6009), .ZN(n6120) );
  AOI22_X1 U7674 ( .A1(n6013), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8680), .B2(
        n6012), .ZN(n6014) );
  INV_X1 U7675 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n6021) );
  XNOR2_X1 U7676 ( .A(n6027), .B(P2_REG3_REG_19__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U7677 ( .A1(n8687), .A2(n6088), .ZN(n6020) );
  INV_X1 U7678 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7679 ( .A1(n4390), .A2(n6016), .ZN(n6018) );
  INV_X1 U7680 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n7750) );
  OR2_X1 U7681 ( .A1(n6114), .A2(n7750), .ZN(n6017) );
  AND2_X1 U7682 ( .A1(n6018), .A2(n6017), .ZN(n6019) );
  OAI211_X1 U7683 ( .C1(n6286), .C2(n6021), .A(n6020), .B(n6019), .ZN(n8707)
         );
  OR2_X1 U7684 ( .A1(n8823), .A2(n8707), .ZN(n6022) );
  NAND2_X1 U7685 ( .A1(n8678), .A2(n6022), .ZN(n6023) );
  INV_X1 U7686 ( .A(n8707), .ZN(n8218) );
  NAND2_X1 U7687 ( .A1(n7097), .A2(n8249), .ZN(n6025) );
  OR2_X1 U7688 ( .A1(n8250), .A2(n9717), .ZN(n6024) );
  INV_X1 U7689 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9681) );
  INV_X1 U7690 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6026) );
  INV_X1 U7691 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8217) );
  OAI21_X1 U7692 ( .B1(n6027), .B2(n6026), .A(n8217), .ZN(n6028) );
  NAND2_X1 U7693 ( .A1(n6034), .A2(n6028), .ZN(n8666) );
  OR2_X1 U7694 ( .A1(n8666), .A2(n6110), .ZN(n6030) );
  AOI22_X1 U7695 ( .A1(n5921), .A2(P2_REG1_REG_20__SCAN_IN), .B1(n6284), .B2(
        P2_REG2_REG_20__SCAN_IN), .ZN(n6029) );
  OAI211_X1 U7696 ( .C1(n6286), .C2(n9681), .A(n6030), .B(n6029), .ZN(n8658)
         );
  INV_X1 U7697 ( .A(n8658), .ZN(n8684) );
  NAND2_X1 U7698 ( .A1(n8814), .A2(n8684), .ZN(n8357) );
  NAND2_X1 U7699 ( .A1(n7124), .A2(n8249), .ZN(n6033) );
  OR2_X1 U7700 ( .A1(n8250), .A2(n7161), .ZN(n6032) );
  NAND2_X1 U7701 ( .A1(n6034), .A2(n8189), .ZN(n6035) );
  NAND2_X1 U7702 ( .A1(n6041), .A2(n6035), .ZN(n8651) );
  AOI22_X1 U7703 ( .A1(n5921), .A2(P2_REG1_REG_21__SCAN_IN), .B1(n6284), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n6037) );
  NAND2_X1 U7704 ( .A1(n6111), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6036) );
  OAI211_X1 U7705 ( .C1(n8651), .C2(n6077), .A(n6037), .B(n6036), .ZN(n8673)
         );
  NAND2_X1 U7706 ( .A1(n8809), .A2(n8673), .ZN(n6038) );
  INV_X1 U7707 ( .A(n8809), .ZN(n8654) );
  INV_X1 U7708 ( .A(n8673), .ZN(n8641) );
  NAND2_X1 U7709 ( .A1(n7414), .A2(n8249), .ZN(n6040) );
  OR2_X1 U7710 ( .A1(n8250), .A2(n7613), .ZN(n6039) );
  INV_X1 U7711 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U7712 ( .A1(n6041), .A2(n8223), .ZN(n6042) );
  NAND2_X1 U7713 ( .A1(n6043), .A2(n6042), .ZN(n8633) );
  OR2_X1 U7714 ( .A1(n8633), .A2(n6110), .ZN(n6048) );
  INV_X1 U7715 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9571) );
  NAND2_X1 U7716 ( .A1(n6284), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6045) );
  NAND2_X1 U7717 ( .A1(n6111), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6044) );
  OAI211_X1 U7718 ( .C1(n9571), .C2(n6114), .A(n6045), .B(n6044), .ZN(n6046)
         );
  INV_X1 U7719 ( .A(n6046), .ZN(n6047) );
  NAND2_X1 U7720 ( .A1(n6048), .A2(n6047), .ZN(n8659) );
  INV_X1 U7721 ( .A(n8659), .ZN(n8190) );
  NAND2_X1 U7722 ( .A1(n8804), .A2(n8190), .ZN(n8349) );
  INV_X1 U7723 ( .A(n8457), .ZN(n8642) );
  OR2_X1 U7724 ( .A1(n8798), .A2(n8642), .ZN(n8364) );
  NAND2_X1 U7725 ( .A1(n8798), .A2(n8642), .ZN(n8606) );
  NAND2_X1 U7726 ( .A1(n7456), .A2(n8249), .ZN(n6050) );
  OR2_X1 U7727 ( .A1(n8250), .A2(n7457), .ZN(n6049) );
  INV_X1 U7728 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7729 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  AND2_X1 U7730 ( .A1(n6065), .A2(n6053), .ZN(n8603) );
  NAND2_X1 U7731 ( .A1(n8603), .A2(n6088), .ZN(n6058) );
  INV_X1 U7732 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9735) );
  NAND2_X1 U7733 ( .A1(n6284), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6055) );
  INV_X1 U7734 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9721) );
  OR2_X1 U7735 ( .A1(n6286), .A2(n9721), .ZN(n6054) );
  OAI211_X1 U7736 ( .C1(n6290), .C2(n9735), .A(n6055), .B(n6054), .ZN(n6056)
         );
  INV_X1 U7737 ( .A(n6056), .ZN(n6057) );
  NAND2_X1 U7738 ( .A1(n6058), .A2(n6057), .ZN(n8618) );
  INV_X1 U7739 ( .A(n8618), .ZN(n8159) );
  NAND2_X1 U7740 ( .A1(n8792), .A2(n8159), .ZN(n8369) );
  NAND2_X1 U7741 ( .A1(n8597), .A2(n8596), .ZN(n8595) );
  NAND2_X1 U7742 ( .A1(n6059), .A2(n8159), .ZN(n6060) );
  NAND2_X1 U7743 ( .A1(n8595), .A2(n6060), .ZN(n8583) );
  OR2_X1 U7744 ( .A1(n8250), .A2(n7546), .ZN(n6061) );
  INV_X1 U7745 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U7746 ( .A1(n6065), .A2(n6064), .ZN(n6066) );
  NAND2_X1 U7747 ( .A1(n6075), .A2(n6066), .ZN(n8585) );
  OR2_X1 U7748 ( .A1(n8585), .A2(n6077), .ZN(n6071) );
  INV_X1 U7749 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U7750 ( .A1(n6111), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7751 ( .A1(n6284), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6067) );
  OAI211_X1 U7752 ( .C1(n9580), .C2(n6290), .A(n6068), .B(n6067), .ZN(n6069)
         );
  INV_X1 U7753 ( .A(n6069), .ZN(n6070) );
  NAND2_X1 U7754 ( .A1(n6071), .A2(n6070), .ZN(n8456) );
  NAND2_X1 U7755 ( .A1(n7571), .A2(n8249), .ZN(n6073) );
  OR2_X1 U7756 ( .A1(n8250), .A2(n7576), .ZN(n6072) );
  INV_X1 U7757 ( .A(n6075), .ZN(n6074) );
  NAND2_X1 U7758 ( .A1(n6074), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6086) );
  INV_X1 U7759 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8239) );
  NAND2_X1 U7760 ( .A1(n6075), .A2(n8239), .ZN(n6076) );
  NAND2_X1 U7761 ( .A1(n6086), .A2(n6076), .ZN(n8579) );
  OR2_X1 U7762 ( .A1(n8579), .A2(n6077), .ZN(n6082) );
  INV_X1 U7763 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9684) );
  NAND2_X1 U7764 ( .A1(n6111), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7765 ( .A1(n5921), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6078) );
  OAI211_X1 U7766 ( .C1(n4390), .C2(n9684), .A(n6079), .B(n6078), .ZN(n6080)
         );
  INV_X1 U7767 ( .A(n6080), .ZN(n6081) );
  NAND2_X1 U7768 ( .A1(n7586), .A2(n8249), .ZN(n6084) );
  OR2_X1 U7769 ( .A1(n8250), .A2(n7591), .ZN(n6083) );
  INV_X1 U7770 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U7771 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  NAND2_X1 U7772 ( .A1(n8559), .A2(n6088), .ZN(n6094) );
  INV_X1 U7773 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6091) );
  NAND2_X1 U7774 ( .A1(n6284), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6090) );
  NAND2_X1 U7775 ( .A1(n6111), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6089) );
  OAI211_X1 U7776 ( .C1(n6091), .C2(n6290), .A(n6090), .B(n6089), .ZN(n6092)
         );
  INV_X1 U7777 ( .A(n6092), .ZN(n6093) );
  NAND2_X1 U7778 ( .A1(n6094), .A2(n6093), .ZN(n8455) );
  NAND2_X1 U7779 ( .A1(n8777), .A2(n6095), .ZN(n8376) );
  INV_X1 U7780 ( .A(n8777), .ZN(n8561) );
  NAND2_X1 U7781 ( .A1(n9778), .A2(n8249), .ZN(n6097) );
  OR2_X1 U7782 ( .A1(n8250), .A2(n8887), .ZN(n6096) );
  INV_X1 U7783 ( .A(n6100), .ZN(n6098) );
  NAND2_X1 U7784 ( .A1(n6098), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7760) );
  INV_X1 U7785 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U7786 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  NAND2_X1 U7787 ( .A1(n7760), .A2(n6101), .ZN(n7602) );
  OR2_X1 U7788 ( .A1(n7602), .A2(n6110), .ZN(n6107) );
  INV_X1 U7789 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6104) );
  NAND2_X1 U7790 ( .A1(n6111), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7791 ( .A1(n6284), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6102) );
  OAI211_X1 U7792 ( .C1(n6104), .C2(n6114), .A(n6103), .B(n6102), .ZN(n6105)
         );
  INV_X1 U7793 ( .A(n6105), .ZN(n6106) );
  NAND2_X1 U7794 ( .A1(n8771), .A2(n6147), .ZN(n8381) );
  NAND2_X1 U7795 ( .A1(n7733), .A2(n8249), .ZN(n6109) );
  OR2_X1 U7796 ( .A1(n8250), .A2(n7734), .ZN(n6108) );
  OR2_X1 U7797 ( .A1(n7760), .A2(n6110), .ZN(n6117) );
  INV_X1 U7798 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9742) );
  NAND2_X1 U7799 ( .A1(n6284), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7800 ( .A1(n6111), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7801 ( .C1(n6114), .C2(n9742), .A(n6113), .B(n6112), .ZN(n6115)
         );
  INV_X1 U7802 ( .A(n6115), .ZN(n6116) );
  NAND2_X1 U7803 ( .A1(n6117), .A2(n6116), .ZN(n8454) );
  INV_X1 U7804 ( .A(n8454), .ZN(n6118) );
  NAND2_X1 U7805 ( .A1(n7759), .A2(n6118), .ZN(n8386) );
  NAND2_X1 U7806 ( .A1(n6120), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6122) );
  XNOR2_X1 U7807 ( .A(n6122), .B(n6121), .ZN(n6128) );
  NAND2_X1 U7808 ( .A1(n6127), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6126) );
  INV_X1 U7809 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6125) );
  INV_X1 U7810 ( .A(n8436), .ZN(n8271) );
  NAND2_X1 U7811 ( .A1(n6128), .A2(n8271), .ZN(n8445) );
  INV_X1 U7812 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6163) );
  XNOR2_X1 U7813 ( .A(n8445), .B(n4811), .ZN(n8725) );
  AND2_X1 U7814 ( .A1(n8725), .A2(n8730), .ZN(n8686) );
  AND2_X1 U7815 ( .A1(n8257), .A2(n8680), .ZN(n6129) );
  OR2_X1 U7816 ( .A1(n6128), .A2(n8436), .ZN(n8255) );
  NAND2_X1 U7817 ( .A1(n8255), .A2(n8433), .ZN(n10193) );
  INV_X1 U7818 ( .A(n10193), .ZN(n6148) );
  INV_X1 U7819 ( .A(n10214), .ZN(n10242) );
  OR2_X1 U7820 ( .A1(n10206), .A2(n10242), .ZN(n10207) );
  OR2_X1 U7821 ( .A1(n8468), .A2(n10256), .ZN(n8266) );
  INV_X1 U7822 ( .A(n10174), .ZN(n6131) );
  NAND2_X1 U7823 ( .A1(n8467), .A2(n10270), .ZN(n8288) );
  NAND2_X1 U7824 ( .A1(n10176), .A2(n8405), .ZN(n6132) );
  OR2_X1 U7825 ( .A1(n8467), .A2(n10270), .ZN(n8268) );
  NAND2_X1 U7826 ( .A1(n6132), .A2(n8268), .ZN(n6964) );
  INV_X1 U7827 ( .A(n8407), .ZN(n6967) );
  NAND2_X1 U7828 ( .A1(n6964), .A2(n6967), .ZN(n6133) );
  INV_X1 U7829 ( .A(n6980), .ZN(n6135) );
  NOR2_X1 U7830 ( .A1(n8408), .A2(n6135), .ZN(n8299) );
  NAND2_X1 U7831 ( .A1(n6136), .A2(n8314), .ZN(n7181) );
  INV_X1 U7832 ( .A(n8318), .ZN(n8323) );
  INV_X1 U7833 ( .A(n7554), .ZN(n8417) );
  INV_X1 U7834 ( .A(n8261), .ZN(n8704) );
  OR2_X1 U7835 ( .A1(n8826), .A2(n8683), .ZN(n8353) );
  NAND2_X1 U7836 ( .A1(n8826), .A2(n8683), .ZN(n8346) );
  NAND2_X1 U7837 ( .A1(n8353), .A2(n8346), .ZN(n8703) );
  INV_X1 U7838 ( .A(n8346), .ZN(n6138) );
  OR2_X1 U7839 ( .A1(n8823), .A2(n8218), .ZN(n8355) );
  NAND2_X1 U7840 ( .A1(n8823), .A2(n8218), .ZN(n8347) );
  NAND2_X1 U7841 ( .A1(n8355), .A2(n8347), .ZN(n8681) );
  INV_X1 U7842 ( .A(n8347), .ZN(n8670) );
  OR2_X1 U7843 ( .A1(n8809), .A2(n8641), .ZN(n8360) );
  NAND2_X1 U7844 ( .A1(n8809), .A2(n8641), .ZN(n8638) );
  INV_X1 U7845 ( .A(n8596), .ZN(n8605) );
  NOR2_X1 U7846 ( .A1(n8789), .A2(n8608), .ZN(n8372) );
  INV_X1 U7847 ( .A(n8382), .ZN(n6140) );
  INV_X1 U7848 ( .A(n8564), .ZN(n6147) );
  OR2_X1 U7849 ( .A1(n8257), .A2(n8436), .ZN(n6294) );
  OR2_X1 U7850 ( .A1(n6294), .A2(n6417), .ZN(n10210) );
  INV_X1 U7851 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U7852 ( .A1(n6284), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6144) );
  INV_X1 U7853 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6142) );
  OR2_X1 U7854 ( .A1(n6286), .A2(n6142), .ZN(n6143) );
  OAI211_X1 U7855 ( .C1(n6290), .C2(n9581), .A(n6144), .B(n6143), .ZN(n8453)
         );
  INV_X1 U7856 ( .A(n8453), .ZN(n6146) );
  INV_X1 U7857 ( .A(n7589), .ZN(n8443) );
  INV_X1 U7858 ( .A(n6417), .ZN(n8442) );
  OR2_X1 U7859 ( .A1(n6294), .A2(n8442), .ZN(n10211) );
  AOI21_X1 U7860 ( .B1(n8443), .B2(P2_B_REG_SCAN_IN), .A(n10211), .ZN(n8548)
         );
  INV_X1 U7861 ( .A(n8548), .ZN(n6145) );
  OAI222_X1 U7862 ( .A1(n6148), .A2(n4450), .B1(n6147), .B2(n10210), .C1(n6146), .C2(n6145), .ZN(n6149) );
  OR2_X1 U7863 ( .A1(n10215), .A2(n10214), .ZN(n10217) );
  INV_X1 U7864 ( .A(n6771), .ZN(n7248) );
  NAND2_X1 U7865 ( .A1(n6971), .A2(n7248), .ZN(n6717) );
  INV_X1 U7866 ( .A(n7367), .ZN(n7225) );
  OR2_X2 U7867 ( .A1(n7317), .A2(n10295), .ZN(n7499) );
  INV_X1 U7868 ( .A(n7484), .ZN(n9810) );
  INV_X1 U7869 ( .A(n8844), .ZN(n8335) );
  AND2_X2 U7870 ( .A1(n8694), .A2(n8701), .ZN(n8695) );
  NOR2_X1 U7871 ( .A1(n8798), .A2(n8631), .ZN(n8599) );
  NAND2_X1 U7872 ( .A1(n6059), .A2(n8599), .ZN(n8600) );
  NOR2_X2 U7873 ( .A1(n7599), .A2(n7759), .ZN(n8551) );
  AOI21_X1 U7874 ( .B1(n7759), .B2(n7599), .A(n8551), .ZN(n7766) );
  NAND2_X1 U7875 ( .A1(n8257), .A2(n8436), .ZN(n10243) );
  OR2_X2 U7876 ( .A1(n10243), .A2(n8432), .ZN(n10298) );
  INV_X1 U7877 ( .A(n10298), .ZN(n8852) );
  NAND2_X1 U7878 ( .A1(n6128), .A2(n8730), .ZN(n6221) );
  INV_X1 U7879 ( .A(n10243), .ZN(n6150) );
  NOR4_X1 U7880 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n6154) );
  NOR4_X1 U7881 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6153) );
  NOR4_X1 U7882 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6152) );
  NOR4_X1 U7883 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6151) );
  NAND4_X1 U7884 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n6173)
         );
  NOR2_X1 U7885 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .ZN(
        n6158) );
  NOR4_X1 U7886 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6157) );
  NOR4_X1 U7887 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6156) );
  NOR4_X1 U7888 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n6155) );
  NAND4_X1 U7889 ( .A1(n6158), .A2(n6157), .A3(n6156), .A4(n6155), .ZN(n6172)
         );
  OR2_X1 U7890 ( .A1(n6160), .A2(n6159), .ZN(n6162) );
  XNOR2_X1 U7891 ( .A(n6162), .B(n6161), .ZN(n7545) );
  NAND2_X1 U7892 ( .A1(n6164), .A2(n6163), .ZN(n6165) );
  NAND2_X1 U7893 ( .A1(n6165), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  INV_X1 U7894 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6175) );
  NAND2_X1 U7895 ( .A1(n6176), .A2(n6175), .ZN(n6166) );
  NAND2_X1 U7896 ( .A1(n6166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6167) );
  XOR2_X1 U7897 ( .A(n7455), .B(P2_B_REG_SCAN_IN), .Z(n6168) );
  NAND2_X1 U7898 ( .A1(n6169), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6170) );
  XNOR2_X1 U7899 ( .A(n6170), .B(n5010), .ZN(n7574) );
  OAI21_X1 U7900 ( .B1(n6173), .B2(n6172), .A(n10225), .ZN(n6214) );
  NOR2_X1 U7901 ( .A1(n7574), .A2(n7545), .ZN(n6174) );
  NAND2_X1 U7902 ( .A1(n7455), .A2(n6174), .ZN(n6398) );
  XNOR2_X1 U7903 ( .A(n6176), .B(n6175), .ZN(n6295) );
  NAND2_X1 U7904 ( .A1(n6398), .A2(n10240), .ZN(n8446) );
  INV_X1 U7905 ( .A(n6294), .ZN(n6400) );
  NAND2_X1 U7906 ( .A1(n6400), .A2(n6221), .ZN(n6228) );
  INV_X1 U7907 ( .A(n6228), .ZN(n6177) );
  NOR2_X1 U7908 ( .A1(n8446), .A2(n6177), .ZN(n6899) );
  NAND2_X1 U7909 ( .A1(n10293), .A2(n8436), .ZN(n6226) );
  NAND3_X1 U7910 ( .A1(n6214), .A2(n6899), .A3(n6226), .ZN(n6179) );
  INV_X1 U7911 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10238) );
  INV_X1 U7912 ( .A(n7574), .ZN(n6180) );
  INV_X1 U7913 ( .A(n7545), .ZN(n6178) );
  NOR2_X1 U7914 ( .A1(n6180), .A2(n6178), .ZN(n10239) );
  AOI21_X1 U7915 ( .B1(n10225), .B2(n10238), .A(n10239), .ZN(n6215) );
  NOR2_X1 U7916 ( .A1(n6179), .A2(n6215), .ZN(n6184) );
  OR2_X1 U7917 ( .A1(n7455), .A2(n6180), .ZN(n10233) );
  INV_X1 U7918 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7919 ( .A1(n10225), .A2(n6181), .ZN(n6182) );
  NAND2_X1 U7920 ( .A1(n10233), .A2(n6182), .ZN(n6897) );
  INV_X1 U7921 ( .A(n6897), .ZN(n6183) );
  AND2_X2 U7922 ( .A1(n6184), .A2(n6183), .ZN(n10319) );
  AND2_X2 U7923 ( .A1(n6184), .A2(n6897), .ZN(n10306) );
  NAND2_X1 U7924 ( .A1(n6185), .A2(n10306), .ZN(n6188) );
  INV_X1 U7925 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6186) );
  OR2_X1 U7926 ( .A1(n10306), .A2(n6186), .ZN(n6187) );
  NAND2_X1 U7927 ( .A1(n6188), .A2(n6187), .ZN(P2_U3517) );
  NAND2_X1 U7928 ( .A1(n7936), .A2(n6384), .ZN(n6189) );
  NAND2_X1 U7929 ( .A1(n6189), .A2(n7418), .ZN(n6248) );
  NAND2_X1 U7930 ( .A1(n6248), .A2(n6190), .ZN(n6310) );
  NAND2_X1 U7931 ( .A1(n6310), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X1 U7932 ( .A(n7418), .ZN(n6191) );
  NOR2_X1 U7933 ( .A1(n6384), .A2(n6191), .ZN(n9873) );
  XNOR2_X1 U7934 ( .A(n6192), .B(n6201), .ZN(n6816) );
  NAND2_X1 U7935 ( .A1(n8467), .A2(n6204), .ZN(n6193) );
  OR2_X1 U7936 ( .A1(n6816), .A2(n6193), .ZN(n6764) );
  NAND2_X1 U7937 ( .A1(n6193), .A2(n6816), .ZN(n6194) );
  NAND2_X1 U7938 ( .A1(n6764), .A2(n6194), .ZN(n6218) );
  OR2_X1 U7939 ( .A1(n10204), .A2(n6725), .ZN(n6724) );
  OR2_X1 U7940 ( .A1(n8138), .A2(n10214), .ZN(n6195) );
  XNOR2_X1 U7941 ( .A(n10215), .B(n8138), .ZN(n6196) );
  XNOR2_X1 U7942 ( .A(n6198), .B(n6196), .ZN(n10139) );
  INV_X1 U7943 ( .A(n6196), .ZN(n6197) );
  NAND2_X1 U7944 ( .A1(n6198), .A2(n6197), .ZN(n6199) );
  NAND2_X1 U7945 ( .A1(n5806), .A2(n6204), .ZN(n6202) );
  XNOR2_X1 U7946 ( .A(n6201), .B(n6200), .ZN(n6912) );
  NAND2_X1 U7947 ( .A1(n6202), .A2(n6912), .ZN(n6203) );
  NAND2_X1 U7948 ( .A1(n8468), .A2(n6204), .ZN(n6205) );
  XNOR2_X1 U7949 ( .A(n6201), .B(n8290), .ZN(n6849) );
  OR2_X1 U7950 ( .A1(n6205), .A2(n6849), .ZN(n6208) );
  NAND2_X1 U7951 ( .A1(n6205), .A2(n6849), .ZN(n6206) );
  AND2_X1 U7952 ( .A1(n6208), .A2(n6206), .ZN(n6913) );
  NAND2_X1 U7953 ( .A1(n6207), .A2(n6913), .ZN(n6916) );
  NAND2_X1 U7954 ( .A1(n10191), .A2(n6204), .ZN(n6212) );
  XNOR2_X1 U7955 ( .A(n10182), .B(n8138), .ZN(n6210) );
  XNOR2_X1 U7956 ( .A(n6212), .B(n6210), .ZN(n6850) );
  AND2_X1 U7957 ( .A1(n6850), .A2(n6208), .ZN(n6209) );
  INV_X1 U7958 ( .A(n6210), .ZN(n6211) );
  NAND2_X1 U7959 ( .A1(n6212), .A2(n6211), .ZN(n6213) );
  NAND2_X1 U7960 ( .A1(n6215), .A2(n6214), .ZN(n6895) );
  NOR2_X1 U7961 ( .A1(n6897), .A2(n6895), .ZN(n6225) );
  INV_X1 U7962 ( .A(n8446), .ZN(n6216) );
  NAND2_X1 U7963 ( .A1(n6225), .A2(n6216), .ZN(n6220) );
  INV_X1 U7964 ( .A(n6766), .ZN(n6818) );
  AOI211_X1 U7965 ( .C1(n6218), .C2(n6217), .A(n8233), .B(n6818), .ZN(n6234)
         );
  OR2_X1 U7966 ( .A1(n10243), .A2(n6128), .ZN(n10205) );
  OR2_X1 U7967 ( .A1(n6220), .A2(n10205), .ZN(n6219) );
  NOR2_X1 U7968 ( .A1(n10143), .A2(n10270), .ZN(n6233) );
  INV_X1 U7969 ( .A(n10191), .ZN(n6909) );
  INV_X1 U7970 ( .A(n6220), .ZN(n6223) );
  INV_X1 U7971 ( .A(n6221), .ZN(n6222) );
  INV_X1 U7972 ( .A(n8466), .ZN(n6224) );
  OAI22_X1 U7973 ( .A1(n6909), .A2(n8224), .B1(n8225), .B2(n6224), .ZN(n6232)
         );
  INV_X1 U7974 ( .A(n6225), .ZN(n6227) );
  NAND2_X1 U7975 ( .A1(n6227), .A2(n6226), .ZN(n6619) );
  AND3_X1 U7976 ( .A1(n6398), .A2(n6295), .A3(n6228), .ZN(n6229) );
  NAND2_X1 U7977 ( .A1(n6619), .A2(n6229), .ZN(n6230) );
  OAI22_X1 U7978 ( .A1(n8240), .A2(n6958), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5836), .ZN(n6231) );
  OR4_X1 U7979 ( .A1(n6234), .A2(n6233), .A3(n6232), .A4(n6231), .ZN(P2_U3229)
         );
  INV_X1 U7980 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6929) );
  NOR2_X1 U7981 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6929), .ZN(n6570) );
  OR2_X1 U7982 ( .A1(n9856), .A2(n6235), .ZN(n6237) );
  INV_X1 U7983 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6311) );
  MUX2_X1 U7984 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6235), .S(n9856), .Z(n9852)
         );
  INV_X1 U7985 ( .A(n9851), .ZN(n6236) );
  AND2_X1 U7986 ( .A1(n6237), .A2(n6236), .ZN(n9863) );
  XNOR2_X1 U7987 ( .A(n9860), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n9862) );
  AOI21_X1 U7988 ( .B1(n9860), .B2(P1_REG1_REG_2__SCAN_IN), .A(n9861), .ZN(
        n6242) );
  NAND2_X1 U7989 ( .A1(P1_REG1_REG_3__SCAN_IN), .A2(n6328), .ZN(n6238) );
  OAI21_X1 U7990 ( .B1(n6328), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6238), .ZN(
        n6241) );
  NOR2_X1 U7991 ( .A1(n6242), .A2(n6241), .ZN(n6327) );
  OR2_X1 U7992 ( .A1(n9874), .A2(P1_U3084), .ZN(n9779) );
  INV_X1 U7993 ( .A(n9869), .ZN(n6239) );
  NOR2_X1 U7994 ( .A1(n9779), .A2(n6239), .ZN(n6240) );
  NAND2_X1 U7995 ( .A1(n6248), .A2(n6240), .ZN(n9907) );
  AOI211_X1 U7996 ( .C1(n6242), .C2(n6241), .A(n6327), .B(n9907), .ZN(n6254)
         );
  OR2_X1 U7997 ( .A1(n9856), .A2(n6243), .ZN(n6245) );
  NAND2_X1 U7998 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n9871) );
  INV_X1 U7999 ( .A(n9849), .ZN(n6244) );
  NAND2_X1 U8000 ( .A1(n9860), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6246) );
  OAI21_X1 U8001 ( .B1(n9860), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6246), .ZN(
        n9865) );
  NAND2_X1 U8002 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(n6328), .ZN(n6247) );
  OAI21_X1 U8003 ( .B1(n6328), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6247), .ZN(
        n6249) );
  NOR2_X1 U8004 ( .A1(n9869), .A2(P1_U3084), .ZN(n7587) );
  AND2_X1 U8005 ( .A1(n6248), .A2(n7587), .ZN(n9105) );
  NAND2_X1 U8006 ( .A1(n9105), .A2(n6380), .ZN(n9944) );
  AOI211_X1 U8007 ( .C1(n6250), .C2(n6249), .A(n6322), .B(n9944), .ZN(n6253)
         );
  INV_X1 U8008 ( .A(n9950), .ZN(n9091) );
  OR2_X1 U8009 ( .A1(P1_U3083), .A2(n9873), .ZN(n9942) );
  INV_X1 U8010 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6251) );
  OAI22_X1 U8011 ( .A1(n9091), .A2(n6264), .B1(n9942), .B2(n6251), .ZN(n6252)
         );
  OR4_X1 U8012 ( .A1(n6570), .A2(n6254), .A3(n6253), .A4(n6252), .ZN(P1_U3244)
         );
  AND2_X1 U8013 ( .A1(n6259), .A2(P2_U3152), .ZN(n6751) );
  INV_X2 U8014 ( .A(n6751), .ZN(n8888) );
  AND2_X1 U8015 ( .A1(n7800), .A2(P2_U3152), .ZN(n8884) );
  INV_X2 U8016 ( .A(n8884), .ZN(n8883) );
  OAI222_X1 U8017 ( .A1(n8888), .A2(n6256), .B1(n8883), .B2(n6269), .C1(n6415), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U8018 ( .A1(n8888), .A2(n6257), .B1(n8883), .B2(n6261), .C1(
        P2_U3152), .C2(n6414), .ZN(P2_U3356) );
  OAI222_X1 U8019 ( .A1(n8888), .A2(n6258), .B1(n8883), .B2(n6263), .C1(
        P2_U3152), .C2(n6476), .ZN(P2_U3355) );
  AND2_X1 U8020 ( .A1(n6259), .A2(P1_U3084), .ZN(n9777) );
  OAI222_X1 U8021 ( .A1(n6262), .A2(P1_U3084), .B1(n4389), .B2(n6261), .C1(
        n6260), .C2(n9782), .ZN(P1_U3351) );
  OAI222_X1 U8022 ( .A1(n6264), .A2(P1_U3084), .B1(n4389), .B2(n6263), .C1(
        n9547), .C2(n9782), .ZN(P1_U3350) );
  OAI222_X1 U8023 ( .A1(n8888), .A2(n9744), .B1(n8883), .B2(n6268), .C1(
        P2_U3152), .C2(n6424), .ZN(P2_U3354) );
  OAI222_X1 U8024 ( .A1(n8888), .A2(n6265), .B1(n8883), .B2(n6266), .C1(
        P2_U3152), .C2(n6465), .ZN(P2_U3353) );
  OAI222_X1 U8025 ( .A1(n9782), .A2(n9730), .B1(n4389), .B2(n6266), .C1(n6320), 
        .C2(P1_U3084), .ZN(P1_U3348) );
  OAI222_X1 U8026 ( .A1(n6329), .A2(P1_U3084), .B1(n4389), .B2(n6268), .C1(
        n6267), .C2(n9782), .ZN(P1_U3349) );
  OAI222_X1 U8027 ( .A1(P1_U3084), .A2(n9856), .B1(n4389), .B2(n6269), .C1(
        n9621), .C2(n9782), .ZN(P1_U3352) );
  INV_X1 U8028 ( .A(n6270), .ZN(n6272) );
  INV_X1 U8029 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6271) );
  OAI222_X1 U8030 ( .A1(n4667), .A2(P1_U3084), .B1(n4389), .B2(n6272), .C1(
        n6271), .C2(n9782), .ZN(P1_U3347) );
  INV_X1 U8031 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9731) );
  INV_X1 U8032 ( .A(n6433), .ZN(n6454) );
  OAI222_X1 U8033 ( .A1(n8888), .A2(n9731), .B1(n8883), .B2(n6272), .C1(
        P2_U3152), .C2(n6454), .ZN(P2_U3352) );
  INV_X1 U8034 ( .A(n6366), .ZN(n6336) );
  INV_X1 U8035 ( .A(n6273), .ZN(n6274) );
  INV_X1 U8036 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9659) );
  OAI222_X1 U8037 ( .A1(n6336), .A2(P1_U3084), .B1(n4389), .B2(n6274), .C1(
        n9659), .C2(n9782), .ZN(P1_U3346) );
  INV_X1 U8038 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6275) );
  INV_X1 U8039 ( .A(n6516), .ZN(n6442) );
  OAI222_X1 U8040 ( .A1(n8888), .A2(n6275), .B1(n8883), .B2(n6274), .C1(
        P2_U3152), .C2(n6442), .ZN(P2_U3351) );
  INV_X1 U8041 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U8042 ( .A1(n6276), .A2(n6379), .ZN(n6277) );
  OAI21_X1 U8043 ( .B1(n6379), .B2(n6278), .A(n6277), .ZN(P1_U3441) );
  INV_X1 U8044 ( .A(n9914), .ZN(n6364) );
  INV_X1 U8045 ( .A(n6279), .ZN(n6281) );
  OAI222_X1 U8046 ( .A1(n6364), .A2(P1_U3084), .B1(n4389), .B2(n6281), .C1(
        n6280), .C2(n9782), .ZN(P1_U3345) );
  INV_X1 U8047 ( .A(n6662), .ZN(n6655) );
  OAI222_X1 U8048 ( .A1(n8888), .A2(n6282), .B1(n8883), .B2(n6281), .C1(
        P2_U3152), .C2(n6655), .ZN(P2_U3350) );
  NAND2_X1 U8049 ( .A1(n10206), .A2(P2_U3966), .ZN(n6283) );
  OAI21_X1 U8050 ( .B1(P2_U3966), .B2(n5132), .A(n6283), .ZN(P2_U3552) );
  INV_X1 U8051 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U8052 ( .A1(n6284), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6288) );
  INV_X1 U8053 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6285) );
  OR2_X1 U8054 ( .A1(n6286), .A2(n6285), .ZN(n6287) );
  OAI211_X1 U8055 ( .C1(n6290), .C2(n6289), .A(n6288), .B(n6287), .ZN(n8547)
         );
  NAND2_X1 U8056 ( .A1(n8547), .A2(P2_U3966), .ZN(n6291) );
  OAI21_X1 U8057 ( .B1(P2_U3966), .B2(n7805), .A(n6291), .ZN(P2_U3583) );
  INV_X1 U8058 ( .A(n6292), .ZN(n6298) );
  INV_X1 U8059 ( .A(n9782), .ZN(n9774) );
  AOI22_X1 U8060 ( .A1(n9924), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n9774), .ZN(n6293) );
  OAI21_X1 U8061 ( .B1(n6298), .B2(n4389), .A(n6293), .ZN(P1_U3344) );
  OAI21_X1 U8062 ( .B1(n8446), .B2(n6294), .A(n6401), .ZN(n6297) );
  OR2_X1 U8063 ( .A1(n6295), .A2(P2_U3152), .ZN(n8451) );
  NAND2_X1 U8064 ( .A1(n8446), .A2(n8451), .ZN(n6296) );
  NAND2_X1 U8065 ( .A1(n6297), .A2(n6296), .ZN(n9788) );
  INV_X1 U8066 ( .A(n9788), .ZN(n10162) );
  NOR2_X1 U8067 ( .A1(n10162), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8068 ( .A(n8475), .ZN(n6652) );
  OAI222_X1 U8069 ( .A1(n8888), .A2(n6299), .B1(n8883), .B2(n6298), .C1(n6652), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  INV_X1 U8070 ( .A(n6300), .ZN(n6303) );
  AOI22_X1 U8071 ( .A1(n6607), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9774), .ZN(n6301) );
  OAI21_X1 U8072 ( .B1(n6303), .B2(n4389), .A(n6301), .ZN(P1_U3343) );
  AOI22_X1 U8073 ( .A1(n8489), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n6751), .ZN(n6302) );
  OAI21_X1 U8074 ( .B1(n6303), .B2(n8883), .A(n6302), .ZN(P2_U3348) );
  INV_X1 U8075 ( .A(n9942), .ZN(n9955) );
  AND2_X1 U8076 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6304) );
  OAI22_X1 U8077 ( .A1(n9869), .A2(n6304), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n6389), .ZN(n6308) );
  NOR2_X1 U8078 ( .A1(n9869), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6305) );
  OR2_X1 U8079 ( .A1(n9779), .A2(n6305), .ZN(n6307) );
  NAND2_X1 U8080 ( .A1(P1_STATE_REG_SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6306) );
  NAND2_X1 U8081 ( .A1(n6307), .A2(n6306), .ZN(n9872) );
  OAI21_X1 U8082 ( .B1(n9874), .B2(n6308), .A(n9872), .ZN(n6309) );
  OAI22_X1 U8083 ( .A1(n6310), .A2(n6309), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6865), .ZN(n6313) );
  NOR3_X1 U8084 ( .A1(n9907), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6311), .ZN(
        n6312) );
  AOI211_X1 U8085 ( .C1(P1_ADDR_REG_0__SCAN_IN), .C2(n9955), .A(n6313), .B(
        n6312), .ZN(n6314) );
  INV_X1 U8086 ( .A(n6314), .ZN(P1_U3241) );
  INV_X1 U8087 ( .A(n6315), .ZN(n6318) );
  INV_X1 U8088 ( .A(n7134), .ZN(n7128) );
  OAI222_X1 U8089 ( .A1(n8888), .A2(n6316), .B1(n8883), .B2(n6318), .C1(n7128), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  INV_X1 U8090 ( .A(n9929), .ZN(n6598) );
  OAI222_X1 U8091 ( .A1(P1_U3084), .A2(n6598), .B1(n4389), .B2(n6318), .C1(
        n6317), .C2(n9782), .ZN(P1_U3342) );
  INV_X1 U8092 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n6340) );
  INV_X1 U8093 ( .A(n9944), .ZN(n9937) );
  NOR2_X1 U8094 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6366), .ZN(n6319) );
  AOI21_X1 U8095 ( .B1(n6366), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6319), .ZN(
        n6324) );
  MUX2_X1 U8096 ( .A(n4666), .B(P1_REG2_REG_6__SCAN_IN), .S(n6331), .Z(n6349)
         );
  AOI22_X1 U8097 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n9901), .B1(n6320), .B2(
        n5200), .ZN(n9892) );
  INV_X1 U8098 ( .A(n6329), .ZN(n9881) );
  MUX2_X1 U8099 ( .A(n6321), .B(P1_REG2_REG_4__SCAN_IN), .S(n6329), .Z(n9883)
         );
  AOI21_X1 U8100 ( .B1(n6328), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6322), .ZN(
        n9884) );
  NAND2_X1 U8101 ( .A1(n9883), .A2(n9884), .ZN(n9882) );
  OAI21_X1 U8102 ( .B1(P1_REG2_REG_4__SCAN_IN), .B2(n9881), .A(n9882), .ZN(
        n9893) );
  NAND2_X1 U8103 ( .A1(n6324), .A2(n6323), .ZN(n6365) );
  OAI21_X1 U8104 ( .B1(n6324), .B2(n6323), .A(n6365), .ZN(n6338) );
  INV_X1 U8105 ( .A(n9907), .ZN(n9956) );
  NOR2_X1 U8106 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6366), .ZN(n6325) );
  AOI21_X1 U8107 ( .B1(n6366), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6325), .ZN(
        n6333) );
  MUX2_X1 U8108 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6326), .S(n6331), .Z(n6342)
         );
  XNOR2_X1 U8109 ( .A(n6329), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9879) );
  AOI21_X1 U8110 ( .B1(n6328), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6327), .ZN(
        n9878) );
  MUX2_X1 U8111 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5196), .S(n9901), .Z(n9894)
         );
  AOI21_X1 U8112 ( .B1(n9901), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9897), .ZN(
        n6343) );
  OAI21_X1 U8113 ( .B1(n6331), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6341), .ZN(
        n6332) );
  NAND2_X1 U8114 ( .A1(n6333), .A2(n6332), .ZN(n6359) );
  OAI21_X1 U8115 ( .B1(n6333), .B2(n6332), .A(n6359), .ZN(n6334) );
  AND2_X1 U8116 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6706) );
  AOI21_X1 U8117 ( .B1(n9956), .B2(n6334), .A(n6706), .ZN(n6335) );
  OAI21_X1 U8118 ( .B1(n9091), .B2(n6336), .A(n6335), .ZN(n6337) );
  AOI21_X1 U8119 ( .B1(n9937), .B2(n6338), .A(n6337), .ZN(n6339) );
  OAI21_X1 U8120 ( .B1(n9942), .B2(n6340), .A(n6339), .ZN(P1_U3248) );
  OAI21_X1 U8121 ( .B1(n6343), .B2(n6342), .A(n6341), .ZN(n6345) );
  NOR2_X1 U8122 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6344), .ZN(n7081) );
  AOI21_X1 U8123 ( .B1(n9956), .B2(n6345), .A(n7081), .ZN(n6346) );
  OAI21_X1 U8124 ( .B1(n9091), .B2(n4667), .A(n6346), .ZN(n6351) );
  AOI211_X1 U8125 ( .C1(n6349), .C2(n6348), .A(n6347), .B(n9944), .ZN(n6350)
         );
  AOI211_X1 U8126 ( .C1(P1_ADDR_REG_6__SCAN_IN), .C2(n9955), .A(n6351), .B(
        n6350), .ZN(n6352) );
  INV_X1 U8127 ( .A(n6352), .ZN(P1_U3247) );
  INV_X1 U8128 ( .A(n6643), .ZN(n6604) );
  INV_X1 U8129 ( .A(n6353), .ZN(n6355) );
  OAI222_X1 U8130 ( .A1(n6604), .A2(P1_U3084), .B1(n4389), .B2(n6355), .C1(
        n6354), .C2(n9782), .ZN(P1_U3341) );
  INV_X1 U8131 ( .A(n8502), .ZN(n7126) );
  OAI222_X1 U8132 ( .A1(n8888), .A2(n6356), .B1(n8883), .B2(n6355), .C1(
        P2_U3152), .C2(n7126), .ZN(P2_U3346) );
  INV_X1 U8133 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6374) );
  NOR2_X1 U8134 ( .A1(P1_REG1_REG_10__SCAN_IN), .A2(n6607), .ZN(n6357) );
  AOI21_X1 U8135 ( .B1(n6607), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6357), .ZN(
        n6362) );
  MUX2_X1 U8136 ( .A(n6358), .B(P1_REG1_REG_8__SCAN_IN), .S(n9914), .Z(n9909)
         );
  OAI21_X1 U8137 ( .B1(n6366), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6359), .ZN(
        n9910) );
  AOI21_X1 U8138 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9914), .A(n9908), .ZN(
        n9923) );
  NOR2_X1 U8139 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n9924), .ZN(n6360) );
  AOI21_X1 U8140 ( .B1(n9924), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6360), .ZN(
        n9922) );
  NAND2_X1 U8141 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  OAI21_X1 U8142 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9924), .A(n9921), .ZN(
        n6361) );
  OAI21_X1 U8143 ( .B1(n6362), .B2(n6361), .A(n6599), .ZN(n6363) );
  NAND2_X1 U8144 ( .A1(n6363), .A2(n9956), .ZN(n6373) );
  AND2_X1 U8145 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7170) );
  AOI22_X1 U8146 ( .A1(n9914), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n5267), .B2(
        n6364), .ZN(n9906) );
  OAI21_X1 U8147 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n6366), .A(n6365), .ZN(
        n9905) );
  NAND2_X1 U8148 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  OAI21_X1 U8149 ( .B1(n9914), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9904), .ZN(
        n9919) );
  MUX2_X1 U8150 ( .A(n6367), .B(P1_REG2_REG_9__SCAN_IN), .S(n9924), .Z(n9918)
         );
  NOR2_X1 U8151 ( .A1(n9919), .A2(n9918), .ZN(n9917) );
  NAND2_X1 U8152 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n6607), .ZN(n6368) );
  OAI21_X1 U8153 ( .B1(n6607), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6368), .ZN(
        n6369) );
  AOI211_X1 U8154 ( .C1(n6370), .C2(n6369), .A(n6606), .B(n9944), .ZN(n6371)
         );
  AOI211_X1 U8155 ( .C1(n9950), .C2(n6607), .A(n7170), .B(n6371), .ZN(n6372)
         );
  OAI211_X1 U8156 ( .C1(n9942), .C2(n6374), .A(n6373), .B(n6372), .ZN(P1_U3251) );
  OR2_X1 U8157 ( .A1(n6376), .A2(n6375), .ZN(n6532) );
  NOR2_X1 U8158 ( .A1(n6532), .A2(n6524), .ZN(n6382) );
  INV_X1 U8159 ( .A(n6382), .ZN(n6577) );
  AOI21_X1 U8160 ( .B1(n8099), .B2(n6377), .A(n10072), .ZN(n6378) );
  NAND2_X1 U8161 ( .A1(n6577), .A2(n6378), .ZN(n6579) );
  AND2_X1 U8162 ( .A1(n6379), .A2(n6574), .ZN(n6534) );
  AND2_X1 U8163 ( .A1(n6579), .A2(n6534), .ZN(n6709) );
  INV_X1 U8164 ( .A(n6709), .ZN(n8929) );
  AOI21_X1 U8165 ( .B1(n6577), .B2(n10116), .A(n8929), .ZN(n6558) );
  NOR2_X2 U8166 ( .A1(n6503), .A2(n6380), .ZN(n9007) );
  NAND2_X1 U8167 ( .A1(n10116), .A2(n7936), .ZN(n6573) );
  NOR2_X1 U8168 ( .A1(n6573), .A2(n10072), .ZN(n6381) );
  NAND2_X1 U8169 ( .A1(n6384), .A2(n6383), .ZN(n6493) );
  NAND2_X1 U8170 ( .A1(n4385), .A2(n6388), .ZN(n6387) );
  INV_X1 U8171 ( .A(n6383), .ZN(n6733) );
  INV_X1 U8172 ( .A(n6384), .ZN(n6385) );
  AOI22_X1 U8173 ( .A1(n4386), .A2(n6863), .B1(n6385), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6386) );
  AND2_X1 U8174 ( .A1(n6387), .A2(n6386), .ZN(n6393) );
  NAND2_X1 U8175 ( .A1(n6388), .A2(n4391), .ZN(n6392) );
  OAI22_X1 U8176 ( .A1(n6493), .A2(n6529), .B1(n6384), .B2(n6389), .ZN(n6390)
         );
  INV_X1 U8177 ( .A(n6390), .ZN(n6391) );
  AOI22_X1 U8178 ( .A1(n9007), .A2(n9039), .B1(n8951), .B2(n9870), .ZN(n6395)
         );
  NAND2_X1 U8179 ( .A1(n9023), .A2(n6863), .ZN(n6394) );
  OAI211_X1 U8180 ( .C1(n6558), .C2(n6865), .A(n6395), .B(n6394), .ZN(P1_U3230) );
  INV_X1 U8181 ( .A(n6396), .ZN(n6477) );
  AOI22_X1 U8182 ( .A1(n7006), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9774), .ZN(n6397) );
  OAI21_X1 U8183 ( .B1(n6477), .B2(n4389), .A(n6397), .ZN(P1_U3340) );
  OR2_X1 U8184 ( .A1(n6417), .A2(P2_U3152), .ZN(n8885) );
  OR2_X1 U8185 ( .A1(n6398), .A2(n8885), .ZN(n6399) );
  OAI211_X1 U8186 ( .C1(n8446), .C2(n6400), .A(n8451), .B(n6399), .ZN(n6402)
         );
  NAND2_X1 U8187 ( .A1(n6402), .A2(n6401), .ZN(n6407) );
  INV_X2 U8188 ( .A(P2_U3966), .ZN(n8469) );
  NAND2_X1 U8189 ( .A1(n6407), .A2(n8469), .ZN(n6419) );
  AND2_X1 U8190 ( .A1(n6419), .A2(n6417), .ZN(n10166) );
  AND2_X1 U8191 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6412) );
  NAND2_X1 U8192 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9785) );
  MUX2_X1 U8193 ( .A(n6403), .B(P2_REG1_REG_1__SCAN_IN), .S(n9791), .Z(n9786)
         );
  NOR2_X1 U8194 ( .A1(n9785), .A2(n9786), .ZN(n9784) );
  AOI21_X1 U8195 ( .B1(n9791), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9784), .ZN(
        n9801) );
  NAND2_X1 U8196 ( .A1(n9803), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6404) );
  OAI21_X1 U8197 ( .B1(n9803), .B2(P2_REG1_REG_2__SCAN_IN), .A(n6404), .ZN(
        n9800) );
  NOR2_X1 U8198 ( .A1(n9801), .A2(n9800), .ZN(n9799) );
  AOI21_X1 U8199 ( .B1(n9803), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9799), .ZN(
        n6468) );
  NAND2_X1 U8200 ( .A1(n6413), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6405) );
  OAI21_X1 U8201 ( .B1(n6413), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6405), .ZN(
        n6467) );
  NOR2_X1 U8202 ( .A1(n6468), .A2(n6467), .ZN(n6466) );
  AOI21_X1 U8203 ( .B1(n6413), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6466), .ZN(
        n6410) );
  MUX2_X1 U8204 ( .A(n6406), .B(P2_REG1_REG_4__SCAN_IN), .S(n6435), .Z(n6409)
         );
  NOR2_X1 U8205 ( .A1(n6410), .A2(n6409), .ZN(n6425) );
  INV_X1 U8206 ( .A(n6407), .ZN(n6408) );
  INV_X1 U8207 ( .A(n10168), .ZN(n10153) );
  AOI211_X1 U8208 ( .C1(n6410), .C2(n6409), .A(n6425), .B(n10153), .ZN(n6411)
         );
  AOI211_X1 U8209 ( .C1(n10162), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6412), .B(
        n6411), .ZN(n6423) );
  AOI22_X1 U8210 ( .A1(n6435), .A2(P2_REG2_REG_4__SCAN_IN), .B1(n5822), .B2(
        n6424), .ZN(n6421) );
  AOI22_X1 U8211 ( .A1(n6413), .A2(P2_REG2_REG_3__SCAN_IN), .B1(n5809), .B2(
        n6476), .ZN(n6473) );
  NAND2_X1 U8212 ( .A1(n9803), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6416) );
  AOI22_X1 U8213 ( .A1(n9803), .A2(P2_REG2_REG_2__SCAN_IN), .B1(n5793), .B2(
        n6414), .ZN(n9806) );
  AOI22_X1 U8214 ( .A1(n9791), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n5771), .B2(
        n6415), .ZN(n9796) );
  NAND3_X1 U8215 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n9796), .ZN(n9794) );
  NAND2_X1 U8216 ( .A1(n6416), .A2(n9804), .ZN(n6472) );
  NAND2_X1 U8217 ( .A1(n6473), .A2(n6472), .ZN(n6471) );
  OAI21_X1 U8218 ( .B1(n5809), .B2(n6476), .A(n6471), .ZN(n6420) );
  NOR2_X1 U8219 ( .A1(n6417), .A2(n7589), .ZN(n6418) );
  NAND2_X1 U8220 ( .A1(n6421), .A2(n6420), .ZN(n6436) );
  OAI211_X1 U8221 ( .C1(n6421), .C2(n6420), .A(n10151), .B(n6436), .ZN(n6422)
         );
  OAI211_X1 U8222 ( .C1(n10152), .C2(n6424), .A(n6423), .B(n6422), .ZN(
        P2_U3249) );
  AND2_X1 U8223 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6432) );
  AOI21_X1 U8224 ( .B1(n6435), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6425), .ZN(
        n6457) );
  NAND2_X1 U8225 ( .A1(n6434), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6426) );
  OAI21_X1 U8226 ( .B1(n6434), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6426), .ZN(
        n6456) );
  NOR2_X1 U8227 ( .A1(n6457), .A2(n6456), .ZN(n6455) );
  AOI21_X1 U8228 ( .B1(n6434), .B2(P2_REG1_REG_5__SCAN_IN), .A(n6455), .ZN(
        n6446) );
  MUX2_X1 U8229 ( .A(n6427), .B(P2_REG1_REG_6__SCAN_IN), .S(n6433), .Z(n6445)
         );
  NOR2_X1 U8230 ( .A1(n6446), .A2(n6445), .ZN(n6444) );
  AOI21_X1 U8231 ( .B1(n6433), .B2(P2_REG1_REG_6__SCAN_IN), .A(n6444), .ZN(
        n6430) );
  NAND2_X1 U8232 ( .A1(n6516), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6428) );
  OAI21_X1 U8233 ( .B1(n6516), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6428), .ZN(
        n6429) );
  NOR2_X1 U8234 ( .A1(n6430), .A2(n6429), .ZN(n6510) );
  AOI211_X1 U8235 ( .C1(n6430), .C2(n6429), .A(n6510), .B(n10153), .ZN(n6431)
         );
  AOI211_X1 U8236 ( .C1(n10162), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6432), .B(
        n6431), .ZN(n6441) );
  AOI22_X1 U8237 ( .A1(n6516), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n5860), .B2(
        n6442), .ZN(n6439) );
  AOI22_X1 U8238 ( .A1(n6433), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n6973), .B2(
        n6454), .ZN(n6451) );
  AOI22_X1 U8239 ( .A1(n6434), .A2(P2_REG2_REG_5__SCAN_IN), .B1(n6959), .B2(
        n6465), .ZN(n6462) );
  NAND2_X1 U8240 ( .A1(n6435), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6437) );
  NAND2_X1 U8241 ( .A1(n6437), .A2(n6436), .ZN(n6461) );
  NAND2_X1 U8242 ( .A1(n6451), .A2(n6450), .ZN(n6449) );
  OAI21_X1 U8243 ( .B1(n6973), .B2(n6454), .A(n6449), .ZN(n6438) );
  NAND2_X1 U8244 ( .A1(n6439), .A2(n6438), .ZN(n6517) );
  OAI211_X1 U8245 ( .C1(n6439), .C2(n6438), .A(n10151), .B(n6517), .ZN(n6440)
         );
  OAI211_X1 U8246 ( .C1(n10152), .C2(n6442), .A(n6441), .B(n6440), .ZN(
        P2_U3252) );
  NOR2_X1 U8247 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6443), .ZN(n6448) );
  AOI211_X1 U8248 ( .C1(n6446), .C2(n6445), .A(n6444), .B(n10153), .ZN(n6447)
         );
  AOI211_X1 U8249 ( .C1(n10162), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6448), .B(
        n6447), .ZN(n6453) );
  OAI211_X1 U8250 ( .C1(n6451), .C2(n6450), .A(n10151), .B(n6449), .ZN(n6452)
         );
  OAI211_X1 U8251 ( .C1(n10152), .C2(n6454), .A(n6453), .B(n6452), .ZN(
        P2_U3251) );
  NOR2_X1 U8252 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5836), .ZN(n6459) );
  AOI211_X1 U8253 ( .C1(n6457), .C2(n6456), .A(n6455), .B(n10153), .ZN(n6458)
         );
  AOI211_X1 U8254 ( .C1(n10162), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6459), .B(
        n6458), .ZN(n6464) );
  OAI211_X1 U8255 ( .C1(n6462), .C2(n6461), .A(n10151), .B(n6460), .ZN(n6463)
         );
  OAI211_X1 U8256 ( .C1(n10152), .C2(n6465), .A(n6464), .B(n6463), .ZN(
        P2_U3250) );
  INV_X1 U8257 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6908) );
  NOR2_X1 U8258 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6908), .ZN(n6470) );
  AOI211_X1 U8259 ( .C1(n6468), .C2(n6467), .A(n6466), .B(n10153), .ZN(n6469)
         );
  AOI211_X1 U8260 ( .C1(n10162), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6470), .B(
        n6469), .ZN(n6475) );
  OAI211_X1 U8261 ( .C1(n6473), .C2(n6472), .A(n10151), .B(n6471), .ZN(n6474)
         );
  OAI211_X1 U8262 ( .C1(n10152), .C2(n6476), .A(n6475), .B(n6474), .ZN(
        P2_U3248) );
  INV_X1 U8263 ( .A(n10167), .ZN(n7133) );
  OAI222_X1 U8264 ( .A1(n8888), .A2(n9678), .B1(n8883), .B2(n6477), .C1(n7133), 
        .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8265 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9647) );
  INV_X1 U8266 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6483) );
  NAND2_X1 U8267 ( .A1(n6478), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6482) );
  INV_X1 U8268 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6479) );
  OR2_X1 U8269 ( .A1(n6480), .A2(n6479), .ZN(n6481) );
  OAI211_X1 U8270 ( .C1(n6484), .C2(n6483), .A(n6482), .B(n6481), .ZN(n9111)
         );
  NAND2_X1 U8271 ( .A1(P1_U4006), .A2(n9111), .ZN(n6485) );
  OAI21_X1 U8272 ( .B1(P1_U4006), .B2(n9647), .A(n6485), .ZN(P1_U3586) );
  INV_X1 U8273 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6487) );
  NAND2_X1 U8274 ( .A1(P1_U4006), .A2(n6388), .ZN(n6486) );
  OAI21_X1 U8275 ( .B1(P1_U4006), .B2(n6487), .A(n6486), .ZN(P1_U3555) );
  INV_X1 U8276 ( .A(n6488), .ZN(n6491) );
  INV_X1 U8277 ( .A(n7515), .ZN(n7144) );
  OAI222_X1 U8278 ( .A1(n8888), .A2(n6489), .B1(n8883), .B2(n6491), .C1(n7144), 
        .C2(P2_U3152), .ZN(P2_U3344) );
  INV_X1 U8279 ( .A(n9047), .ZN(n9040) );
  OAI222_X1 U8280 ( .A1(P1_U3084), .A2(n9040), .B1(n4389), .B2(n6491), .C1(
        n6490), .C2(n9782), .ZN(P1_U3339) );
  INV_X1 U8281 ( .A(n6500), .ZN(n6498) );
  NAND2_X1 U8282 ( .A1(n6492), .A2(n4391), .ZN(n6495) );
  NAND2_X1 U8284 ( .A1(n6674), .A2(n6747), .ZN(n6494) );
  NAND2_X1 U8285 ( .A1(n6495), .A2(n6494), .ZN(n6496) );
  XNOR2_X1 U8286 ( .A(n6496), .B(n7770), .ZN(n6499) );
  INV_X1 U8287 ( .A(n6499), .ZN(n6497) );
  NAND2_X1 U8288 ( .A1(n6498), .A2(n6497), .ZN(n6549) );
  NAND2_X1 U8289 ( .A1(n6500), .A2(n6499), .ZN(n6550) );
  NAND2_X1 U8290 ( .A1(n6549), .A2(n6550), .ZN(n6502) );
  AOI22_X1 U8291 ( .A1(n7634), .A2(n9039), .B1(n4388), .B2(n6747), .ZN(n6548)
         );
  XNOR2_X1 U8292 ( .A(n6502), .B(n6548), .ZN(n6508) );
  NOR2_X2 U8293 ( .A1(n6503), .A2(n9874), .ZN(n9019) );
  AOI22_X1 U8294 ( .A1(n9007), .A2(n6542), .B1(n9019), .B2(n6388), .ZN(n6504)
         );
  OAI21_X1 U8295 ( .B1(n6558), .B2(n6505), .A(n6504), .ZN(n6506) );
  AOI21_X1 U8296 ( .B1(n9023), .B2(n6747), .A(n6506), .ZN(n6507) );
  OAI21_X1 U8297 ( .B1(n6508), .B2(n9025), .A(n6507), .ZN(P1_U3220) );
  NOR2_X1 U8298 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6509), .ZN(n6515) );
  AOI21_X1 U8299 ( .B1(n6516), .B2(P2_REG1_REG_7__SCAN_IN), .A(n6510), .ZN(
        n6513) );
  MUX2_X1 U8300 ( .A(n6511), .B(P2_REG1_REG_8__SCAN_IN), .S(n6662), .Z(n6512)
         );
  NOR2_X1 U8301 ( .A1(n6513), .A2(n6512), .ZN(n6661) );
  AOI211_X1 U8302 ( .C1(n6513), .C2(n6512), .A(n6661), .B(n10153), .ZN(n6514)
         );
  AOI211_X1 U8303 ( .C1(n10162), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6515), .B(
        n6514), .ZN(n6522) );
  AOI22_X1 U8304 ( .A1(n6662), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n6990), .B2(
        n6655), .ZN(n6520) );
  NAND2_X1 U8305 ( .A1(n6516), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8306 ( .A1(n6518), .A2(n6517), .ZN(n6519) );
  OAI211_X1 U8307 ( .C1(n6520), .C2(n6519), .A(n10151), .B(n6654), .ZN(n6521)
         );
  OAI211_X1 U8308 ( .C1(n10152), .C2(n6655), .A(n6522), .B(n6521), .ZN(
        P2_U3253) );
  OR2_X1 U8309 ( .A1(n9473), .A2(n4392), .ZN(n6523) );
  INV_X2 U8310 ( .A(n10124), .ZN(n10126) );
  INV_X1 U8311 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8312 ( .A1(n6388), .A2(n6529), .ZN(n8061) );
  INV_X1 U8313 ( .A(n6862), .ZN(n6526) );
  AOI211_X1 U8314 ( .C1(n6740), .C2(n8061), .A(n6527), .B(n6526), .ZN(n6528)
         );
  AOI21_X1 U8315 ( .B1(n9985), .B2(n9039), .A(n6528), .ZN(n6864) );
  OAI21_X1 U8316 ( .B1(n6529), .B2(n6862), .A(n6864), .ZN(n6536) );
  NAND2_X1 U8317 ( .A1(n6536), .A2(n10126), .ZN(n6530) );
  OAI21_X1 U8318 ( .B1(n10126), .B2(n6531), .A(n6530), .ZN(P1_U3454) );
  INV_X1 U8319 ( .A(n6532), .ZN(n6535) );
  NAND3_X1 U8320 ( .A1(n6535), .A2(n6534), .A3(n6533), .ZN(n10134) );
  NAND2_X1 U8321 ( .A1(n6536), .A2(n4387), .ZN(n6537) );
  OAI21_X1 U8322 ( .B1(n4387), .B2(n6389), .A(n6537), .ZN(P1_U3523) );
  OR2_X1 U8323 ( .A1(n10028), .A2(n10116), .ZN(n10080) );
  OAI22_X1 U8324 ( .A1(n9005), .A2(n5135), .B1(n8929), .B2(n10080), .ZN(n6538)
         );
  AOI21_X1 U8325 ( .B1(n9007), .B2(n10009), .A(n6538), .ZN(n6556) );
  NAND2_X1 U8326 ( .A1(n6542), .A2(n4388), .ZN(n6540) );
  NAND2_X1 U8327 ( .A1(n6674), .A2(n10023), .ZN(n6539) );
  NAND2_X1 U8328 ( .A1(n6540), .A2(n6539), .ZN(n6541) );
  XNOR2_X1 U8329 ( .A(n6541), .B(n7770), .ZN(n6546) );
  INV_X1 U8330 ( .A(n6546), .ZN(n6544) );
  AOI22_X1 U8331 ( .A1(n7634), .A2(n6542), .B1(n4388), .B2(n10023), .ZN(n6545)
         );
  INV_X1 U8332 ( .A(n6545), .ZN(n6543) );
  NAND2_X1 U8333 ( .A1(n6544), .A2(n6543), .ZN(n6547) );
  NAND2_X1 U8334 ( .A1(n6546), .A2(n6545), .ZN(n6566) );
  NAND2_X1 U8335 ( .A1(n6549), .A2(n6548), .ZN(n6551) );
  NAND2_X1 U8336 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  NAND2_X1 U8337 ( .A1(n6552), .A2(n6553), .ZN(n6567) );
  OAI21_X1 U8338 ( .B1(n6553), .B2(n6552), .A(n6567), .ZN(n6554) );
  NAND2_X1 U8339 ( .A1(n6554), .A2(n8951), .ZN(n6555) );
  OAI211_X1 U8340 ( .C1(n6558), .C2(n6557), .A(n6556), .B(n6555), .ZN(P1_U3235) );
  NAND2_X1 U8341 ( .A1(n10009), .A2(n4386), .ZN(n6560) );
  NAND2_X1 U8342 ( .A1(n6674), .A2(n6562), .ZN(n6559) );
  NAND2_X1 U8343 ( .A1(n6560), .A2(n6559), .ZN(n6561) );
  XNOR2_X1 U8344 ( .A(n6561), .B(n7770), .ZN(n6564) );
  AOI22_X1 U8345 ( .A1(n7634), .A2(n10009), .B1(n4388), .B2(n6562), .ZN(n6563)
         );
  NAND2_X1 U8346 ( .A1(n6564), .A2(n6563), .ZN(n6588) );
  OR2_X1 U8347 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  AND2_X1 U8348 ( .A1(n6588), .A2(n6565), .ZN(n6569) );
  NAND2_X1 U8349 ( .A1(n6567), .A2(n6566), .ZN(n6568) );
  OAI21_X1 U8350 ( .B1(n6569), .B2(n6568), .A(n6589), .ZN(n6583) );
  INV_X1 U8351 ( .A(n9038), .ZN(n6572) );
  AOI21_X1 U8352 ( .B1(n9019), .B2(n6542), .A(n6570), .ZN(n6571) );
  OAI21_X1 U8353 ( .B1(n9017), .B2(n6572), .A(n6571), .ZN(n6582) );
  INV_X1 U8354 ( .A(n9023), .ZN(n8958) );
  INV_X1 U8355 ( .A(n6573), .ZN(n6576) );
  NAND3_X1 U8356 ( .A1(n6574), .A2(n6384), .A3(n7418), .ZN(n6575) );
  AOI21_X1 U8357 ( .B1(n6577), .B2(n6576), .A(n6575), .ZN(n6578) );
  OR2_X1 U8358 ( .A1(n6578), .A2(P1_U3084), .ZN(n6580) );
  OAI22_X1 U8359 ( .A1(n8958), .A2(n10087), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9021), .ZN(n6581) );
  AOI211_X1 U8360 ( .C1(n8951), .C2(n6583), .A(n6582), .B(n6581), .ZN(n6584)
         );
  INV_X1 U8361 ( .A(n6584), .ZN(P1_U3216) );
  NAND2_X1 U8362 ( .A1(n9038), .A2(n4391), .ZN(n6586) );
  NAND2_X1 U8363 ( .A1(n6674), .A2(n9998), .ZN(n6585) );
  NAND2_X1 U8364 ( .A1(n6586), .A2(n6585), .ZN(n6587) );
  INV_X2 U8365 ( .A(n7770), .ZN(n7716) );
  XNOR2_X1 U8366 ( .A(n6587), .B(n7716), .ZN(n6680) );
  AOI22_X1 U8367 ( .A1(n7634), .A2(n9038), .B1(n4386), .B2(n9998), .ZN(n6681)
         );
  XNOR2_X1 U8368 ( .A(n6680), .B(n6681), .ZN(n6591) );
  NAND2_X1 U8369 ( .A1(n6589), .A2(n6588), .ZN(n6590) );
  OAI21_X1 U8370 ( .B1(n6591), .B2(n6590), .A(n6684), .ZN(n6596) );
  INV_X1 U8371 ( .A(n9986), .ZN(n6593) );
  AND2_X1 U8372 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9887) );
  AOI21_X1 U8373 ( .B1(n9019), .B2(n10009), .A(n9887), .ZN(n6592) );
  OAI21_X1 U8374 ( .B1(n9017), .B2(n6593), .A(n6592), .ZN(n6595) );
  OAI22_X1 U8375 ( .A1(n8958), .A2(n10093), .B1(n9021), .B2(n9993), .ZN(n6594)
         );
  AOI211_X1 U8376 ( .C1(n6596), .C2(n8951), .A(n6595), .B(n6594), .ZN(n6597)
         );
  INV_X1 U8377 ( .A(n6597), .ZN(P1_U3228) );
  AOI22_X1 U8378 ( .A1(n9929), .A2(P1_REG1_REG_11__SCAN_IN), .B1(n5320), .B2(
        n6598), .ZN(n9932) );
  NAND2_X1 U8379 ( .A1(n9932), .A2(n9931), .ZN(n9930) );
  OAI21_X1 U8380 ( .B1(n9929), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9930), .ZN(
        n6602) );
  MUX2_X1 U8381 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n6600), .S(n6643), .Z(n6601)
         );
  NAND2_X1 U8382 ( .A1(n6601), .A2(n6602), .ZN(n6635) );
  OAI21_X1 U8383 ( .B1(n6602), .B2(n6601), .A(n6635), .ZN(n6613) );
  NAND2_X1 U8384 ( .A1(n9955), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U8385 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7407) );
  OAI211_X1 U8386 ( .C1(n9091), .C2(n6604), .A(n6603), .B(n7407), .ZN(n6612)
         );
  NOR2_X1 U8387 ( .A1(n9929), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6605) );
  AOI21_X1 U8388 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9929), .A(n6605), .ZN(
        n9935) );
  OAI21_X1 U8389 ( .B1(n9929), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9933), .ZN(
        n6610) );
  NAND2_X1 U8390 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n6643), .ZN(n6608) );
  OAI21_X1 U8391 ( .B1(n6643), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6608), .ZN(
        n6609) );
  NOR2_X1 U8392 ( .A1(n6609), .A2(n6610), .ZN(n6642) );
  AOI211_X1 U8393 ( .C1(n6610), .C2(n6609), .A(n6642), .B(n9944), .ZN(n6611)
         );
  AOI211_X1 U8394 ( .C1(n6613), .C2(n9956), .A(n6612), .B(n6611), .ZN(n6614)
         );
  INV_X1 U8395 ( .A(n6614), .ZN(P1_U3253) );
  INV_X1 U8396 ( .A(n6615), .ZN(n6618) );
  INV_X1 U8397 ( .A(n8515), .ZN(n7520) );
  OAI222_X1 U8398 ( .A1(n8888), .A2(n6616), .B1(n8883), .B2(n6618), .C1(
        P2_U3152), .C2(n7520), .ZN(P2_U3343) );
  OAI222_X1 U8399 ( .A1(n9063), .A2(P1_U3084), .B1(n4389), .B2(n6618), .C1(
        n6617), .C2(n9782), .ZN(P1_U3338) );
  INV_X1 U8400 ( .A(n8468), .ZN(n8291) );
  INV_X1 U8401 ( .A(n5787), .ZN(n6938) );
  OAI22_X1 U8402 ( .A1(n8291), .A2(n8225), .B1(n8224), .B2(n6938), .ZN(n6621)
         );
  AND2_X1 U8403 ( .A1(n6619), .A2(n6899), .ZN(n10150) );
  OAI22_X1 U8404 ( .A1(n10143), .A2(n10251), .B1(n10150), .B2(n6941), .ZN(
        n6620) );
  NOR2_X1 U8405 ( .A1(n6621), .A2(n6620), .ZN(n6624) );
  INV_X1 U8406 ( .A(n8233), .ZN(n10141) );
  OAI211_X1 U8407 ( .C1(n4493), .C2(n6622), .A(n6915), .B(n10141), .ZN(n6623)
         );
  NAND2_X1 U8408 ( .A1(n6624), .A2(n6623), .ZN(P2_U3239) );
  INV_X1 U8409 ( .A(n6625), .ZN(n6628) );
  INV_X1 U8410 ( .A(n7747), .ZN(n7742) );
  OAI222_X1 U8411 ( .A1(n8888), .A2(n6626), .B1(n8883), .B2(n6628), .C1(n7742), 
        .C2(P2_U3152), .ZN(P2_U3342) );
  INV_X1 U8412 ( .A(n9083), .ZN(n6627) );
  OAI222_X1 U8413 ( .A1(n9782), .A2(n9709), .B1(n4389), .B2(n6628), .C1(
        P1_U3084), .C2(n6627), .ZN(P1_U3337) );
  INV_X1 U8414 ( .A(n6629), .ZN(n6631) );
  AOI22_X1 U8415 ( .A1(n9102), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9774), .ZN(n6630) );
  OAI21_X1 U8416 ( .B1(n6631), .B2(n4389), .A(n6630), .ZN(P1_U3336) );
  INV_X1 U8417 ( .A(n7748), .ZN(n8533) );
  OAI222_X1 U8418 ( .A1(n8888), .A2(n6632), .B1(n8883), .B2(n6631), .C1(n8533), 
        .C2(P2_U3152), .ZN(P2_U3341) );
  INV_X1 U8419 ( .A(n7006), .ZN(n6641) );
  NOR2_X1 U8420 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6633), .ZN(n7471) );
  INV_X1 U8421 ( .A(n7471), .ZN(n6640) );
  MUX2_X1 U8422 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n6634), .S(n7006), .Z(n6637)
         );
  OAI21_X1 U8423 ( .B1(n6643), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6635), .ZN(
        n6636) );
  OAI21_X1 U8424 ( .B1(n6637), .B2(n6636), .A(n6999), .ZN(n6638) );
  NAND2_X1 U8425 ( .A1(n9956), .A2(n6638), .ZN(n6639) );
  OAI211_X1 U8426 ( .C1(n9091), .C2(n6641), .A(n6640), .B(n6639), .ZN(n6649)
         );
  NOR2_X1 U8427 ( .A1(n7006), .A2(n6644), .ZN(n6645) );
  AOI21_X1 U8428 ( .B1(n7006), .B2(n6644), .A(n6645), .ZN(n6646) );
  AOI211_X1 U8429 ( .C1(n6647), .C2(n6646), .A(n7005), .B(n9944), .ZN(n6648)
         );
  AOI211_X1 U8430 ( .C1(P1_ADDR_REG_13__SCAN_IN), .C2(n9955), .A(n6649), .B(
        n6648), .ZN(n6650) );
  INV_X1 U8431 ( .A(n6650), .ZN(P1_U3254) );
  AOI22_X1 U8432 ( .A1(n7134), .A2(n5925), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n7128), .ZN(n6659) );
  NAND2_X1 U8433 ( .A1(n8489), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6657) );
  MUX2_X1 U8434 ( .A(n7187), .B(P2_REG2_REG_10__SCAN_IN), .S(n8489), .Z(n6651)
         );
  INV_X1 U8435 ( .A(n6651), .ZN(n8485) );
  NAND2_X1 U8436 ( .A1(n8475), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6656) );
  INV_X1 U8437 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6653) );
  AOI22_X1 U8438 ( .A1(n8475), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n6653), .B2(
        n6652), .ZN(n8471) );
  NAND2_X1 U8439 ( .A1(n8471), .A2(n8472), .ZN(n8470) );
  NAND2_X1 U8440 ( .A1(n6656), .A2(n8470), .ZN(n8486) );
  NOR2_X1 U8441 ( .A1(n6659), .A2(n6658), .ZN(n7127) );
  AOI21_X1 U8442 ( .B1(n6659), .B2(n6658), .A(n7127), .ZN(n6673) );
  INV_X1 U8443 ( .A(n10151), .ZN(n10172) );
  NOR2_X1 U8444 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5922), .ZN(n6660) );
  AOI21_X1 U8445 ( .B1(n10162), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6660), .ZN(
        n6670) );
  INV_X1 U8446 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7373) );
  MUX2_X1 U8447 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7373), .S(n7134), .Z(n6668)
         );
  MUX2_X1 U8448 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n5909), .S(n8489), .Z(n8492)
         );
  NAND2_X1 U8449 ( .A1(n8475), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6665) );
  AOI21_X1 U8450 ( .B1(n6662), .B2(P2_REG1_REG_8__SCAN_IN), .A(n6661), .ZN(
        n8477) );
  MUX2_X1 U8451 ( .A(n6663), .B(P2_REG1_REG_9__SCAN_IN), .S(n8475), .Z(n8478)
         );
  NOR2_X1 U8452 ( .A1(n8477), .A2(n8478), .ZN(n8476) );
  INV_X1 U8453 ( .A(n8476), .ZN(n6664) );
  NAND2_X1 U8454 ( .A1(n6665), .A2(n6664), .ZN(n8491) );
  NAND2_X1 U8455 ( .A1(n8492), .A2(n8491), .ZN(n8490) );
  NAND2_X1 U8456 ( .A1(n8489), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6666) );
  NAND2_X1 U8457 ( .A1(n8490), .A2(n6666), .ZN(n6667) );
  NAND2_X1 U8458 ( .A1(n6667), .A2(n6668), .ZN(n7136) );
  OAI211_X1 U8459 ( .C1(n6668), .C2(n6667), .A(n10168), .B(n7136), .ZN(n6669)
         );
  OAI211_X1 U8460 ( .C1(n10152), .C2(n7128), .A(n6670), .B(n6669), .ZN(n6671)
         );
  INV_X1 U8461 ( .A(n6671), .ZN(n6672) );
  OAI21_X1 U8462 ( .B1(n6673), .B2(n10172), .A(n6672), .ZN(P2_U3256) );
  NAND2_X1 U8463 ( .A1(n6703), .A2(n6674), .ZN(n6676) );
  NAND2_X1 U8464 ( .A1(n9036), .A2(n4388), .ZN(n6675) );
  NAND2_X1 U8465 ( .A1(n6676), .A2(n6675), .ZN(n6677) );
  XNOR2_X1 U8466 ( .A(n6677), .B(n7716), .ZN(n6873) );
  NAND2_X1 U8467 ( .A1(n6703), .A2(n4391), .ZN(n6679) );
  NAND2_X1 U8468 ( .A1(n7634), .A2(n9036), .ZN(n6678) );
  NAND2_X1 U8469 ( .A1(n6679), .A2(n6678), .ZN(n6874) );
  XNOR2_X1 U8470 ( .A(n6873), .B(n6874), .ZN(n6702) );
  INV_X1 U8471 ( .A(n6680), .ZN(n6682) );
  NAND2_X1 U8472 ( .A1(n6682), .A2(n6681), .ZN(n6683) );
  NAND2_X1 U8473 ( .A1(n6674), .A2(n7102), .ZN(n6685) );
  NAND2_X1 U8474 ( .A1(n7634), .A2(n9986), .ZN(n6687) );
  NAND2_X1 U8475 ( .A1(n4386), .A2(n7102), .ZN(n6686) );
  NAND2_X1 U8476 ( .A1(n6687), .A2(n6686), .ZN(n6692) );
  NAND2_X1 U8477 ( .A1(n6753), .A2(n6692), .ZN(n6688) );
  NAND2_X1 U8478 ( .A1(n9037), .A2(n4391), .ZN(n6690) );
  NAND2_X1 U8479 ( .A1(n7095), .A2(n6674), .ZN(n6689) );
  NAND2_X1 U8480 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  XNOR2_X1 U8481 ( .A(n6691), .B(n7770), .ZN(n6697) );
  AOI22_X1 U8482 ( .A1(n7634), .A2(n9037), .B1(n4388), .B2(n7095), .ZN(n6696)
         );
  NAND2_X1 U8483 ( .A1(n6697), .A2(n6696), .ZN(n7088) );
  INV_X1 U8484 ( .A(n6753), .ZN(n6693) );
  INV_X1 U8485 ( .A(n6692), .ZN(n6755) );
  NAND2_X1 U8486 ( .A1(n6693), .A2(n6755), .ZN(n6694) );
  AND2_X1 U8487 ( .A1(n7088), .A2(n6694), .ZN(n6695) );
  OR2_X1 U8488 ( .A1(n6697), .A2(n6696), .ZN(n7089) );
  INV_X1 U8489 ( .A(n6878), .ZN(n6701) );
  AOI21_X1 U8490 ( .B1(n6702), .B2(n6699), .A(n6701), .ZN(n6711) );
  AND2_X1 U8491 ( .A1(n6703), .A2(n9822), .ZN(n10109) );
  NOR2_X1 U8492 ( .A1(n9017), .A2(n6704), .ZN(n6705) );
  AOI211_X1 U8493 ( .C1(n9019), .C2(n9037), .A(n6706), .B(n6705), .ZN(n6707)
         );
  OAI21_X1 U8494 ( .B1(n9021), .B2(n6805), .A(n6707), .ZN(n6708) );
  AOI21_X1 U8495 ( .B1(n6709), .B2(n10109), .A(n6708), .ZN(n6710) );
  OAI21_X1 U8496 ( .B1(n6711), .B2(n9025), .A(n6710), .ZN(P1_U3211) );
  XNOR2_X1 U8497 ( .A(n6712), .B(n4749), .ZN(n7254) );
  AOI21_X1 U8498 ( .B1(n6713), .B2(n4749), .A(n6148), .ZN(n6716) );
  NAND2_X1 U8499 ( .A1(n8466), .A2(n10189), .ZN(n6715) );
  NAND2_X1 U8500 ( .A1(n8464), .A2(n10190), .ZN(n6714) );
  NAND2_X1 U8501 ( .A1(n6715), .A2(n6714), .ZN(n6778) );
  AOI21_X1 U8502 ( .B1(n6716), .B2(n6981), .A(n6778), .ZN(n7249) );
  INV_X1 U8503 ( .A(n6971), .ZN(n6718) );
  INV_X1 U8504 ( .A(n6717), .ZN(n6988) );
  AOI21_X1 U8505 ( .B1(n6771), .B2(n6718), .A(n6988), .ZN(n7252) );
  AOI22_X1 U8506 ( .A1(n7252), .A2(n8852), .B1(n8851), .B2(n6771), .ZN(n6719)
         );
  OAI211_X1 U8507 ( .C1(n7254), .C2(n8848), .A(n7249), .B(n6719), .ZN(n6721)
         );
  NAND2_X1 U8508 ( .A1(n6721), .A2(n10319), .ZN(n6720) );
  OAI21_X1 U8509 ( .B1(n10319), .B2(n5864), .A(n6720), .ZN(P2_U3527) );
  INV_X1 U8510 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6723) );
  NAND2_X1 U8511 ( .A1(n6721), .A2(n10306), .ZN(n6722) );
  OAI21_X1 U8512 ( .B1(n10306), .B2(n6723), .A(n6722), .ZN(P2_U3472) );
  INV_X1 U8513 ( .A(n6724), .ZN(n6729) );
  NOR2_X1 U8514 ( .A1(n8233), .A2(n6725), .ZN(n8229) );
  AOI22_X1 U8515 ( .A1(n8229), .A2(n10206), .B1(n10214), .B2(n10141), .ZN(
        n6728) );
  OAI22_X1 U8516 ( .A1(n10143), .A2(n10242), .B1(n10150), .B2(n6901), .ZN(
        n6726) );
  AOI21_X1 U8517 ( .B1(n10136), .B2(n5787), .A(n6726), .ZN(n6727) );
  OAI21_X1 U8518 ( .B1(n6729), .B2(n6728), .A(n6727), .ZN(P2_U3234) );
  OR2_X1 U8519 ( .A1(n6383), .A2(n8092), .ZN(n6926) );
  INV_X1 U8520 ( .A(n6926), .ZN(n6746) );
  XOR2_X1 U8521 ( .A(n6737), .B(n6730), .Z(n6744) );
  INV_X1 U8522 ( .A(n6744), .ZN(n10077) );
  NAND2_X1 U8523 ( .A1(n6747), .A2(n6863), .ZN(n6731) );
  NAND3_X1 U8524 ( .A1(n9469), .A2(n10024), .A3(n6731), .ZN(n10073) );
  OAI22_X1 U8525 ( .A1(n9192), .A2(n10073), .B1(n9994), .B2(n6505), .ZN(n6745)
         );
  NAND2_X1 U8526 ( .A1(n6732), .A2(n4392), .ZN(n6736) );
  OR2_X1 U8527 ( .A1(n6734), .A2(n6733), .ZN(n6735) );
  AND2_X1 U8528 ( .A1(n6736), .A2(n6735), .ZN(n10015) );
  AOI22_X1 U8529 ( .A1(n9985), .A2(n6542), .B1(n6388), .B2(n9987), .ZN(n6743)
         );
  INV_X1 U8530 ( .A(n6737), .ZN(n6741) );
  NOR2_X1 U8531 ( .A1(n8060), .A2(n6738), .ZN(n8029) );
  INV_X1 U8532 ( .A(n8029), .ZN(n6739) );
  OAI211_X1 U8533 ( .C1(n6741), .C2(n6740), .A(n6739), .B(n10019), .ZN(n6742)
         );
  OAI211_X1 U8534 ( .C1(n6744), .C2(n10015), .A(n6743), .B(n6742), .ZN(n10075)
         );
  AOI211_X1 U8535 ( .C1(n6746), .C2(n10077), .A(n6745), .B(n10075), .ZN(n6749)
         );
  AOI22_X1 U8536 ( .A1(n9350), .A2(n6747), .B1(n10021), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6748) );
  OAI21_X1 U8537 ( .B1(n6749), .B2(n9387), .A(n6748), .ZN(P1_U3290) );
  INV_X1 U8538 ( .A(n6750), .ZN(n6763) );
  AOI22_X1 U8539 ( .A1(n8538), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n6751), .ZN(n6752) );
  OAI21_X1 U8540 ( .B1(n6763), .B2(n8883), .A(n6752), .ZN(P2_U3340) );
  NOR2_X1 U8541 ( .A1(n4487), .A2(n6753), .ZN(n7085) );
  AOI21_X1 U8542 ( .B1(n4487), .B2(n6753), .A(n7085), .ZN(n6754) );
  NAND2_X1 U8543 ( .A1(n6754), .A2(n6755), .ZN(n7087) );
  OAI21_X1 U8544 ( .B1(n6755), .B2(n6754), .A(n7087), .ZN(n6760) );
  INV_X1 U8545 ( .A(n9037), .ZN(n6757) );
  NOR2_X1 U8546 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5198), .ZN(n9899) );
  AOI21_X1 U8547 ( .B1(n9019), .B2(n9038), .A(n9899), .ZN(n6756) );
  OAI21_X1 U8548 ( .B1(n9017), .B2(n6757), .A(n6756), .ZN(n6759) );
  OAI22_X1 U8549 ( .A1(n8958), .A2(n10105), .B1(n9021), .B2(n7106), .ZN(n6758)
         );
  AOI211_X1 U8550 ( .C1(n6760), .C2(n8951), .A(n6759), .B(n6758), .ZN(n6761)
         );
  INV_X1 U8551 ( .A(n6761), .ZN(P1_U3225) );
  INV_X1 U8552 ( .A(n9951), .ZN(n9099) );
  INV_X1 U8553 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6762) );
  OAI222_X1 U8554 ( .A1(n9099), .A2(P1_U3084), .B1(n4389), .B2(n6763), .C1(
        n6762), .C2(n9782), .ZN(P1_U3335) );
  XNOR2_X1 U8555 ( .A(n6975), .B(n8138), .ZN(n6767) );
  NAND2_X1 U8556 ( .A1(n8466), .A2(n6204), .ZN(n6768) );
  XNOR2_X1 U8557 ( .A(n6767), .B(n6768), .ZN(n6829) );
  AND2_X1 U8558 ( .A1(n6829), .A2(n6764), .ZN(n6765) );
  NAND2_X1 U8559 ( .A1(n6766), .A2(n6765), .ZN(n6819) );
  INV_X1 U8560 ( .A(n6767), .ZN(n6769) );
  NAND2_X1 U8561 ( .A1(n6769), .A2(n6768), .ZN(n6770) );
  XNOR2_X1 U8562 ( .A(n6771), .B(n8138), .ZN(n6831) );
  AND2_X1 U8563 ( .A1(n8465), .A2(n6204), .ZN(n6772) );
  NAND2_X1 U8564 ( .A1(n6831), .A2(n6772), .ZN(n6836) );
  INV_X1 U8565 ( .A(n6831), .ZN(n6774) );
  INV_X1 U8566 ( .A(n6772), .ZN(n6773) );
  NAND2_X1 U8567 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  NAND2_X1 U8568 ( .A1(n6836), .A2(n6775), .ZN(n6776) );
  AOI211_X1 U8569 ( .C1(n6777), .C2(n6776), .A(n8233), .B(n4488), .ZN(n6783)
         );
  AOI22_X1 U8570 ( .A1(n8242), .A2(n6778), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n6781) );
  INV_X1 U8571 ( .A(n6779), .ZN(n7246) );
  NAND2_X1 U8572 ( .A1(n8210), .A2(n7246), .ZN(n6780) );
  OAI211_X1 U8573 ( .C1(n7248), .C2(n10143), .A(n6781), .B(n6780), .ZN(n6782)
         );
  OR2_X1 U8574 ( .A1(n6783), .A2(n6782), .ZN(P2_U3215) );
  INV_X1 U8575 ( .A(n7820), .ZN(n8032) );
  XNOR2_X1 U8576 ( .A(n6784), .B(n8032), .ZN(n6795) );
  XNOR2_X1 U8577 ( .A(n7819), .B(n8032), .ZN(n6785) );
  AOI222_X1 U8578 ( .A1(n10019), .A2(n6785), .B1(n9036), .B2(n9985), .C1(n9986), .C2(n9987), .ZN(n6794) );
  OAI21_X1 U8579 ( .B1(n7104), .B2(n6786), .A(n9469), .ZN(n6787) );
  NOR2_X1 U8580 ( .A1(n6787), .A2(n6803), .ZN(n6792) );
  NAND2_X1 U8581 ( .A1(n6792), .A2(n8092), .ZN(n6788) );
  OAI211_X1 U8582 ( .C1(n9994), .C2(n7084), .A(n6794), .B(n6788), .ZN(n6789)
         );
  NAND2_X1 U8583 ( .A1(n6789), .A2(n9321), .ZN(n6791) );
  AOI22_X1 U8584 ( .A1(n9350), .A2(n7095), .B1(n10021), .B2(
        P1_REG2_REG_6__SCAN_IN), .ZN(n6790) );
  OAI211_X1 U8585 ( .C1(n9323), .C2(n6795), .A(n6791), .B(n6790), .ZN(P1_U3285) );
  INV_X1 U8586 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n6797) );
  AOI21_X1 U8587 ( .B1(n9822), .B2(n7095), .A(n6792), .ZN(n6793) );
  OAI211_X1 U8588 ( .C1(n9823), .C2(n6795), .A(n6794), .B(n6793), .ZN(n6798)
         );
  NAND2_X1 U8589 ( .A1(n6798), .A2(n10126), .ZN(n6796) );
  OAI21_X1 U8590 ( .B1(n10126), .B2(n6797), .A(n6796), .ZN(P1_U3472) );
  NAND2_X1 U8591 ( .A1(n6798), .A2(n4387), .ZN(n6799) );
  OAI21_X1 U8592 ( .B1(n4387), .B2(n6326), .A(n6799), .ZN(P1_U3529) );
  OAI21_X1 U8593 ( .B1(n8034), .B2(n6801), .A(n6800), .ZN(n6802) );
  AOI222_X1 U8594 ( .A1(n10019), .A2(n6802), .B1(n9037), .B2(n9987), .C1(n9035), .C2(n9985), .ZN(n10112) );
  OAI211_X1 U8595 ( .C1(n6803), .C2(n6808), .A(n9469), .B(n9973), .ZN(n10110)
         );
  INV_X1 U8596 ( .A(n10110), .ZN(n6810) );
  OR2_X1 U8597 ( .A1(n6804), .A2(n9192), .ZN(n9353) );
  INV_X1 U8598 ( .A(n9353), .ZN(n7438) );
  NOR2_X1 U8599 ( .A1(n9994), .A2(n6805), .ZN(n6806) );
  AOI21_X1 U8600 ( .B1(n10021), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6806), .ZN(
        n6807) );
  OAI21_X1 U8601 ( .B1(n10029), .B2(n6808), .A(n6807), .ZN(n6809) );
  AOI21_X1 U8602 ( .B1(n6810), .B2(n7438), .A(n6809), .ZN(n6814) );
  XNOR2_X1 U8603 ( .A(n6811), .B(n6812), .ZN(n10114) );
  INV_X1 U8604 ( .A(n9323), .ZN(n9363) );
  NAND2_X1 U8605 ( .A1(n10114), .A2(n9363), .ZN(n6813) );
  OAI211_X1 U8606 ( .C1(n10112), .C2(n9387), .A(n6814), .B(n6813), .ZN(
        P1_U3284) );
  INV_X1 U8607 ( .A(n8229), .ZN(n7151) );
  INV_X1 U8608 ( .A(n8467), .ZN(n6815) );
  NOR3_X1 U8609 ( .A1(n7151), .A2(n6816), .A3(n6815), .ZN(n6817) );
  AOI21_X1 U8610 ( .B1(n6818), .B2(n10141), .A(n6817), .ZN(n6830) );
  INV_X1 U8611 ( .A(n6819), .ZN(n6827) );
  NAND2_X1 U8612 ( .A1(n8467), .A2(n10189), .ZN(n6821) );
  NAND2_X1 U8613 ( .A1(n8465), .A2(n10190), .ZN(n6820) );
  AND2_X1 U8614 ( .A1(n6821), .A2(n6820), .ZN(n6965) );
  INV_X1 U8615 ( .A(n6965), .ZN(n6822) );
  AOI22_X1 U8616 ( .A1(n8242), .A2(n6822), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n6825) );
  INV_X1 U8617 ( .A(n6972), .ZN(n6823) );
  NAND2_X1 U8618 ( .A1(n8210), .A2(n6823), .ZN(n6824) );
  OAI211_X1 U8619 ( .C1(n10275), .C2(n10143), .A(n6825), .B(n6824), .ZN(n6826)
         );
  AOI21_X1 U8620 ( .B1(n6827), .B2(n10141), .A(n6826), .ZN(n6828) );
  OAI21_X1 U8621 ( .B1(n6830), .B2(n6829), .A(n6828), .ZN(P2_U3241) );
  NAND3_X1 U8622 ( .A1(n8229), .A2(n6831), .A3(n8465), .ZN(n6839) );
  XNOR2_X1 U8623 ( .A(n6992), .B(n8138), .ZN(n6832) );
  AND2_X1 U8624 ( .A1(n8464), .A2(n6204), .ZN(n6833) );
  NAND2_X1 U8625 ( .A1(n6832), .A2(n6833), .ZN(n7029) );
  INV_X1 U8626 ( .A(n6832), .ZN(n7067) );
  INV_X1 U8627 ( .A(n6833), .ZN(n6834) );
  NAND2_X1 U8628 ( .A1(n7067), .A2(n6834), .ZN(n6835) );
  AND2_X1 U8629 ( .A1(n7029), .A2(n6835), .ZN(n6837) );
  OAI21_X1 U8630 ( .B1(n4488), .B2(n6837), .A(n10141), .ZN(n6838) );
  INV_X1 U8631 ( .A(n7075), .ZN(n7069) );
  AOI21_X1 U8632 ( .B1(n6839), .B2(n6838), .A(n7069), .ZN(n6847) );
  INV_X1 U8633 ( .A(n6992), .ZN(n10281) );
  NAND2_X1 U8634 ( .A1(n8465), .A2(n10189), .ZN(n6841) );
  NAND2_X1 U8635 ( .A1(n8463), .A2(n10190), .ZN(n6840) );
  AND2_X1 U8636 ( .A1(n6841), .A2(n6840), .ZN(n6983) );
  INV_X1 U8637 ( .A(n6983), .ZN(n6842) );
  AOI22_X1 U8638 ( .A1(n8242), .A2(n6842), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n6845) );
  INV_X1 U8639 ( .A(n6989), .ZN(n6843) );
  NAND2_X1 U8640 ( .A1(n8210), .A2(n6843), .ZN(n6844) );
  OAI211_X1 U8641 ( .C1(n10281), .C2(n10143), .A(n6845), .B(n6844), .ZN(n6846)
         );
  OR2_X1 U8642 ( .A1(n6847), .A2(n6846), .ZN(P2_U3223) );
  NAND2_X1 U8643 ( .A1(n8229), .A2(n8468), .ZN(n6848) );
  OAI22_X1 U8644 ( .A1(n6916), .A2(n8233), .B1(n6849), .B2(n6848), .ZN(n6858)
         );
  INV_X1 U8645 ( .A(n6850), .ZN(n6857) );
  INV_X1 U8646 ( .A(n8242), .ZN(n8202) );
  NAND2_X1 U8647 ( .A1(n8468), .A2(n10189), .ZN(n6852) );
  NAND2_X1 U8648 ( .A1(n8467), .A2(n10190), .ZN(n6851) );
  NAND2_X1 U8649 ( .A1(n6852), .A2(n6851), .ZN(n10175) );
  INV_X1 U8650 ( .A(n10175), .ZN(n6854) );
  INV_X1 U8651 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6853) );
  OAI22_X1 U8652 ( .A1(n8202), .A2(n6854), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6853), .ZN(n6856) );
  OAI22_X1 U8653 ( .A1(n10262), .A2(n10143), .B1(n8240), .B2(n10180), .ZN(
        n6855) );
  AOI211_X1 U8654 ( .C1(n6858), .C2(n6857), .A(n6856), .B(n6855), .ZN(n6859)
         );
  OAI21_X1 U8655 ( .B1(n6860), .B2(n8233), .A(n6859), .ZN(P2_U3232) );
  INV_X1 U8656 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9550) );
  INV_X1 U8657 ( .A(n6861), .ZN(n8097) );
  OAI21_X1 U8658 ( .B1(n9350), .B2(n10003), .A(n6863), .ZN(n6868) );
  OAI21_X1 U8659 ( .B1(n6865), .B2(n9994), .A(n6864), .ZN(n6866) );
  NAND2_X1 U8660 ( .A1(n6866), .A2(n9321), .ZN(n6867) );
  OAI211_X1 U8661 ( .C1(n9550), .C2(n9321), .A(n6868), .B(n6867), .ZN(P1_U3291) );
  INV_X1 U8662 ( .A(n6869), .ZN(n6872) );
  OAI222_X1 U8663 ( .A1(n8888), .A2(n6870), .B1(n8883), .B2(n6872), .C1(n8730), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U8664 ( .A1(P1_U3084), .A2(n8092), .B1(n4389), .B2(n6872), .C1(
        n6871), .C2(n9782), .ZN(P1_U3334) );
  INV_X1 U8665 ( .A(n6873), .ZN(n6876) );
  INV_X1 U8666 ( .A(n6874), .ZN(n6875) );
  NAND2_X1 U8667 ( .A1(n6876), .A2(n6875), .ZN(n6877) );
  AND2_X1 U8668 ( .A1(n7634), .A2(n9035), .ZN(n6879) );
  AOI21_X1 U8669 ( .B1(n9968), .B2(n4391), .A(n6879), .ZN(n6883) );
  NAND2_X1 U8670 ( .A1(n9968), .A2(n6674), .ZN(n6881) );
  NAND2_X1 U8671 ( .A1(n9035), .A2(n4386), .ZN(n6880) );
  NAND2_X1 U8672 ( .A1(n6881), .A2(n6880), .ZN(n6882) );
  XNOR2_X1 U8673 ( .A(n6882), .B(n7770), .ZN(n6885) );
  NAND2_X1 U8674 ( .A1(n6886), .A2(n6885), .ZN(n7056) );
  INV_X1 U8675 ( .A(n7056), .ZN(n6888) );
  NAND2_X1 U8676 ( .A1(n6884), .A2(n6883), .ZN(n7055) );
  AOI21_X1 U8677 ( .B1(n6886), .B2(n7055), .A(n6885), .ZN(n6887) );
  AOI21_X1 U8678 ( .B1(n6888), .B2(n7055), .A(n6887), .ZN(n6894) );
  NOR2_X1 U8679 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6889), .ZN(n9912) );
  AOI21_X1 U8680 ( .B1(n9019), .B2(n9036), .A(n9912), .ZN(n6891) );
  NAND2_X1 U8681 ( .A1(n9007), .A2(n9034), .ZN(n6890) );
  OAI211_X1 U8682 ( .C1(n9021), .C2(n9969), .A(n6891), .B(n6890), .ZN(n6892)
         );
  AOI21_X1 U8683 ( .B1(n9023), .B2(n9968), .A(n6892), .ZN(n6893) );
  OAI21_X1 U8684 ( .B1(n6894), .B2(n9025), .A(n6893), .ZN(P1_U3219) );
  NAND2_X1 U8685 ( .A1(n10206), .A2(n10242), .ZN(n8275) );
  NAND2_X1 U8686 ( .A1(n10207), .A2(n8275), .ZN(n10245) );
  INV_X1 U8687 ( .A(n10245), .ZN(n6907) );
  INV_X1 U8688 ( .A(n6895), .ZN(n6896) );
  AND2_X1 U8689 ( .A1(n6897), .A2(n6896), .ZN(n6898) );
  NAND2_X1 U8690 ( .A1(n6899), .A2(n6898), .ZN(n6904) );
  NAND2_X2 U8691 ( .A1(n6904), .A2(n10218), .ZN(n10222) );
  INV_X1 U8692 ( .A(n8686), .ZN(n8741) );
  OR2_X1 U8693 ( .A1(n8445), .A2(n8730), .ZN(n7179) );
  NAND2_X1 U8694 ( .A1(n8741), .A2(n7179), .ZN(n10213) );
  NAND2_X1 U8695 ( .A1(n10222), .A2(n10213), .ZN(n8713) );
  AND2_X1 U8696 ( .A1(n5787), .A2(n10190), .ZN(n6900) );
  AOI21_X1 U8697 ( .B1(n10245), .B2(n10193), .A(n6900), .ZN(n10241) );
  OAI22_X1 U8698 ( .A1(n10224), .A2(n10241), .B1(n6901), .B2(n10218), .ZN(
        n6902) );
  AOI21_X1 U8699 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n10224), .A(n6902), .ZN(
        n6906) );
  INV_X1 U8700 ( .A(n10205), .ZN(n6903) );
  OAI21_X1 U8701 ( .B1(n10183), .B2(n8711), .A(n10214), .ZN(n6905) );
  OAI211_X1 U8702 ( .C1(n6907), .C2(n8713), .A(n6906), .B(n6905), .ZN(P2_U3296) );
  OAI22_X1 U8703 ( .A1(n8240), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n6908), .ZN(n6911) );
  OAI22_X1 U8704 ( .A1(n8225), .A2(n6909), .B1(n10256), .B2(n10143), .ZN(n6910) );
  AOI211_X1 U8705 ( .C1(n10137), .C2(n5806), .A(n6911), .B(n6910), .ZN(n6920)
         );
  NOR3_X1 U8706 ( .A1(n7151), .A2(n6912), .A3(n5805), .ZN(n6918) );
  INV_X1 U8707 ( .A(n6913), .ZN(n6914) );
  AOI21_X1 U8708 ( .B1(n6915), .B2(n6914), .A(n8233), .ZN(n6917) );
  OAI21_X1 U8709 ( .B1(n6918), .B2(n6917), .A(n6916), .ZN(n6919) );
  NAND2_X1 U8710 ( .A1(n6920), .A2(n6919), .ZN(P2_U3220) );
  XNOR2_X1 U8711 ( .A(n6921), .B(n8030), .ZN(n6927) );
  AOI22_X1 U8712 ( .A1(n9987), .A2(n6542), .B1(n9038), .B2(n9985), .ZN(n6925)
         );
  XNOR2_X1 U8713 ( .A(n7944), .B(n6922), .ZN(n6923) );
  NAND2_X1 U8714 ( .A1(n6923), .A2(n10019), .ZN(n6924) );
  OAI211_X1 U8715 ( .C1(n6927), .C2(n10015), .A(n6925), .B(n6924), .ZN(n10089)
         );
  INV_X1 U8716 ( .A(n10089), .ZN(n6934) );
  OR2_X1 U8717 ( .A1(n10021), .A2(n6926), .ZN(n10027) );
  INV_X1 U8718 ( .A(n10027), .ZN(n10004) );
  INV_X1 U8719 ( .A(n6927), .ZN(n10091) );
  OR2_X1 U8720 ( .A1(n10022), .A2(n10087), .ZN(n6928) );
  NAND2_X1 U8721 ( .A1(n9999), .A2(n6928), .ZN(n10088) );
  NOR2_X1 U8722 ( .A1(n10032), .A2(n10088), .ZN(n6932) );
  INV_X1 U8723 ( .A(n9994), .ZN(n10020) );
  AOI22_X1 U8724 ( .A1(n10021), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n10020), .B2(
        n6929), .ZN(n6930) );
  OAI21_X1 U8725 ( .B1(n10029), .B2(n10087), .A(n6930), .ZN(n6931) );
  AOI211_X1 U8726 ( .C1(n10004), .C2(n10091), .A(n6932), .B(n6931), .ZN(n6933)
         );
  OAI21_X1 U8727 ( .B1(n10021), .B2(n6934), .A(n6933), .ZN(P1_U3288) );
  XNOR2_X1 U8728 ( .A(n6935), .B(n8402), .ZN(n10255) );
  INV_X1 U8729 ( .A(n10255), .ZN(n6946) );
  XOR2_X1 U8730 ( .A(n8402), .B(n6936), .Z(n6937) );
  OAI222_X1 U8731 ( .A1(n10210), .A2(n6938), .B1(n10211), .B2(n8291), .C1(
        n6148), .C2(n6937), .ZN(n10253) );
  INV_X1 U8732 ( .A(n10217), .ZN(n6940) );
  INV_X1 U8733 ( .A(n10197), .ZN(n6939) );
  OAI21_X1 U8734 ( .B1(n10251), .B2(n6940), .A(n6939), .ZN(n10252) );
  OAI22_X1 U8735 ( .A1(n10219), .A2(n10252), .B1(n6941), .B2(n10218), .ZN(
        n6942) );
  AOI21_X1 U8736 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10224), .A(n6942), .ZN(
        n6943) );
  OAI21_X1 U8737 ( .B1(n10251), .B2(n10200), .A(n6943), .ZN(n6944) );
  AOI21_X1 U8738 ( .B1(n10253), .B2(n10222), .A(n6944), .ZN(n6945) );
  OAI21_X1 U8739 ( .B1(n6946), .B2(n8713), .A(n6945), .ZN(P2_U3294) );
  INV_X1 U8740 ( .A(n6947), .ZN(n6949) );
  INV_X1 U8741 ( .A(n6969), .ZN(n6948) );
  OAI211_X1 U8742 ( .C1(n10270), .C2(n6949), .A(n6948), .B(n8852), .ZN(n10269)
         );
  INV_X1 U8743 ( .A(n10269), .ZN(n6955) );
  NAND2_X1 U8744 ( .A1(n10176), .A2(n6950), .ZN(n6951) );
  NAND2_X1 U8745 ( .A1(n8268), .A2(n8288), .ZN(n6956) );
  XNOR2_X1 U8746 ( .A(n6951), .B(n6956), .ZN(n6952) );
  NAND2_X1 U8747 ( .A1(n6952), .A2(n10193), .ZN(n6954) );
  AOI22_X1 U8748 ( .A1(n10189), .A2(n10191), .B1(n8466), .B2(n10190), .ZN(
        n6953) );
  NAND2_X1 U8749 ( .A1(n6954), .A2(n6953), .ZN(n10271) );
  AOI21_X1 U8750 ( .B1(n6955), .B2(n8730), .A(n10271), .ZN(n6963) );
  XNOR2_X1 U8751 ( .A(n6957), .B(n6956), .ZN(n10273) );
  INV_X1 U8752 ( .A(n8713), .ZN(n10202) );
  NOR2_X1 U8753 ( .A1(n10200), .A2(n10270), .ZN(n6961) );
  OAI22_X1 U8754 ( .A1(n10222), .A2(n6959), .B1(n6958), .B2(n10218), .ZN(n6960) );
  AOI211_X1 U8755 ( .C1(n10273), .C2(n10202), .A(n6961), .B(n6960), .ZN(n6962)
         );
  OAI21_X1 U8756 ( .B1(n6963), .B2(n10224), .A(n6962), .ZN(P2_U3291) );
  XNOR2_X1 U8757 ( .A(n6964), .B(n8407), .ZN(n6966) );
  OAI21_X1 U8758 ( .B1(n6966), .B2(n6148), .A(n6965), .ZN(n10277) );
  INV_X1 U8759 ( .A(n10277), .ZN(n6979) );
  XNOR2_X1 U8760 ( .A(n6968), .B(n6967), .ZN(n10279) );
  NOR2_X1 U8761 ( .A1(n6969), .A2(n10275), .ZN(n6970) );
  OR2_X1 U8762 ( .A1(n6971), .A2(n6970), .ZN(n10276) );
  OAI22_X1 U8763 ( .A1(n10222), .A2(n6973), .B1(n6972), .B2(n10218), .ZN(n6974) );
  AOI21_X1 U8764 ( .B1(n10183), .B2(n6975), .A(n6974), .ZN(n6976) );
  OAI21_X1 U8765 ( .B1(n10276), .B2(n10219), .A(n6976), .ZN(n6977) );
  AOI21_X1 U8766 ( .B1(n10279), .B2(n10202), .A(n6977), .ZN(n6978) );
  OAI21_X1 U8767 ( .B1(n6979), .B2(n10224), .A(n6978), .ZN(P2_U3290) );
  AOI21_X1 U8768 ( .B1(n6981), .B2(n6980), .A(n8307), .ZN(n6982) );
  OAI21_X1 U8769 ( .B1(n4490), .B2(n6982), .A(n10193), .ZN(n6984) );
  NAND2_X1 U8770 ( .A1(n6984), .A2(n6983), .ZN(n10284) );
  INV_X1 U8771 ( .A(n10284), .ZN(n6996) );
  INV_X1 U8772 ( .A(n6985), .ZN(n6986) );
  AOI21_X1 U8773 ( .B1(n8307), .B2(n6987), .A(n6986), .ZN(n10285) );
  OAI21_X1 U8774 ( .B1(n6988), .B2(n10281), .A(n7240), .ZN(n10282) );
  OAI22_X1 U8775 ( .A1(n10222), .A2(n6990), .B1(n6989), .B2(n10218), .ZN(n6991) );
  AOI21_X1 U8776 ( .B1(n10183), .B2(n6992), .A(n6991), .ZN(n6993) );
  OAI21_X1 U8777 ( .B1(n10282), .B2(n10219), .A(n6993), .ZN(n6994) );
  AOI21_X1 U8778 ( .B1(n10285), .B2(n10202), .A(n6994), .ZN(n6995) );
  OAI21_X1 U8779 ( .B1(n10224), .B2(n6996), .A(n6995), .ZN(P2_U3288) );
  NAND2_X1 U8780 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3084), .ZN(n7004) );
  NOR2_X1 U8781 ( .A1(n9040), .A2(n6997), .ZN(n6998) );
  AOI21_X1 U8782 ( .B1(n6997), .B2(n9040), .A(n6998), .ZN(n7001) );
  NAND2_X1 U8783 ( .A1(n7001), .A2(n7000), .ZN(n9046) );
  OAI21_X1 U8784 ( .B1(n7001), .B2(n7000), .A(n9046), .ZN(n7002) );
  NAND2_X1 U8785 ( .A1(n9956), .A2(n7002), .ZN(n7003) );
  OAI211_X1 U8786 ( .C1(n9091), .C2(n9040), .A(n7004), .B(n7003), .ZN(n7009)
         );
  NOR2_X1 U8787 ( .A1(n5372), .A2(n7007), .ZN(n9042) );
  AOI211_X1 U8788 ( .C1(n7007), .C2(n5372), .A(n9042), .B(n9944), .ZN(n7008)
         );
  AOI211_X1 U8789 ( .C1(P1_ADDR_REG_14__SCAN_IN), .C2(n9955), .A(n7009), .B(
        n7008), .ZN(n7010) );
  INV_X1 U8790 ( .A(n7010), .ZN(P1_U3255) );
  AND2_X1 U8791 ( .A1(n7011), .A2(n7967), .ZN(n8035) );
  XNOR2_X1 U8792 ( .A(n7012), .B(n8035), .ZN(n7194) );
  INV_X1 U8793 ( .A(n10015), .ZN(n9992) );
  NAND2_X1 U8794 ( .A1(n7014), .A2(n7013), .ZN(n7015) );
  XNOR2_X1 U8795 ( .A(n7015), .B(n8035), .ZN(n7017) );
  AOI22_X1 U8796 ( .A1(n9987), .A2(n9035), .B1(n9033), .B2(n9985), .ZN(n7016)
         );
  OAI21_X1 U8797 ( .B1(n7017), .B2(n9989), .A(n7016), .ZN(n7018) );
  AOI21_X1 U8798 ( .B1(n7194), .B2(n9992), .A(n7018), .ZN(n7198) );
  INV_X1 U8799 ( .A(n7211), .ZN(n7019) );
  AOI21_X1 U8800 ( .B1(n7195), .B2(n9974), .A(n7019), .ZN(n7196) );
  NAND2_X1 U8801 ( .A1(n7196), .A2(n10003), .ZN(n7022) );
  NOR2_X1 U8802 ( .A1(n9994), .A2(n7062), .ZN(n7020) );
  AOI21_X1 U8803 ( .B1(n10021), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7020), .ZN(
        n7021) );
  OAI211_X1 U8804 ( .C1(n4707), .C2(n10029), .A(n7022), .B(n7021), .ZN(n7023)
         );
  AOI21_X1 U8805 ( .B1(n7194), .B2(n10004), .A(n7023), .ZN(n7024) );
  OAI21_X1 U8806 ( .B1(n7198), .B2(n9387), .A(n7024), .ZN(P1_U3282) );
  XNOR2_X1 U8807 ( .A(n10295), .B(n6201), .ZN(n7025) );
  NAND2_X1 U8808 ( .A1(n8460), .A2(n6204), .ZN(n7026) );
  NAND2_X1 U8809 ( .A1(n7025), .A2(n7026), .ZN(n7292) );
  INV_X1 U8810 ( .A(n7025), .ZN(n7028) );
  INV_X1 U8811 ( .A(n7026), .ZN(n7027) );
  NAND2_X1 U8812 ( .A1(n7028), .A2(n7027), .ZN(n7289) );
  NAND2_X1 U8813 ( .A1(n7292), .A2(n7289), .ZN(n7044) );
  XNOR2_X1 U8814 ( .A(n7421), .B(n8138), .ZN(n7038) );
  NAND2_X1 U8815 ( .A1(n8463), .A2(n6204), .ZN(n7039) );
  XNOR2_X1 U8816 ( .A(n7038), .B(n7039), .ZN(n7079) );
  AND2_X1 U8817 ( .A1(n7079), .A2(n7029), .ZN(n7074) );
  XNOR2_X1 U8818 ( .A(n7367), .B(n8138), .ZN(n7043) );
  XNOR2_X1 U8819 ( .A(n7264), .B(n8138), .ZN(n7032) );
  AND2_X1 U8820 ( .A1(n8462), .A2(n6204), .ZN(n7033) );
  NAND2_X1 U8821 ( .A1(n7032), .A2(n7033), .ZN(n7036) );
  NAND2_X1 U8822 ( .A1(n7075), .A2(n7030), .ZN(n7042) );
  INV_X1 U8823 ( .A(n7032), .ZN(n7152) );
  INV_X1 U8824 ( .A(n7033), .ZN(n7034) );
  NAND2_X1 U8825 ( .A1(n7152), .A2(n7034), .ZN(n7035) );
  NAND2_X1 U8826 ( .A1(n7036), .A2(n7035), .ZN(n7261) );
  INV_X1 U8827 ( .A(n7038), .ZN(n7040) );
  NAND2_X1 U8828 ( .A1(n7040), .A2(n7039), .ZN(n7149) );
  NAND2_X1 U8829 ( .A1(n7042), .A2(n7041), .ZN(n7295) );
  NAND2_X1 U8830 ( .A1(n7043), .A2(n4421), .ZN(n7290) );
  NAND2_X1 U8831 ( .A1(n7295), .A2(n7290), .ZN(n7117) );
  XOR2_X1 U8832 ( .A(n7044), .B(n7117), .Z(n7050) );
  NOR2_X1 U8833 ( .A1(n8240), .A2(n7319), .ZN(n7048) );
  NAND2_X1 U8834 ( .A1(n8461), .A2(n10189), .ZN(n7046) );
  NAND2_X1 U8835 ( .A1(n8459), .A2(n10190), .ZN(n7045) );
  AND2_X1 U8836 ( .A1(n7046), .A2(n7045), .ZN(n7315) );
  OAI22_X1 U8837 ( .A1(n8202), .A2(n7315), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8500), .ZN(n7047) );
  AOI211_X1 U8838 ( .C1(n10295), .C2(n8228), .A(n7048), .B(n7047), .ZN(n7049)
         );
  OAI21_X1 U8839 ( .B1(n7050), .B2(n8233), .A(n7049), .ZN(P2_U3226) );
  NAND2_X1 U8840 ( .A1(n7195), .A2(n6674), .ZN(n7052) );
  NAND2_X1 U8841 ( .A1(n9034), .A2(n4386), .ZN(n7051) );
  NAND2_X1 U8842 ( .A1(n7052), .A2(n7051), .ZN(n7053) );
  XNOR2_X1 U8843 ( .A(n7053), .B(n7716), .ZN(n7166) );
  AND2_X1 U8844 ( .A1(n7634), .A2(n9034), .ZN(n7054) );
  AOI21_X1 U8845 ( .B1(n7195), .B2(n4388), .A(n7054), .ZN(n7167) );
  XNOR2_X1 U8846 ( .A(n7166), .B(n7167), .ZN(n7058) );
  NAND2_X1 U8847 ( .A1(n7056), .A2(n7055), .ZN(n7057) );
  NAND2_X1 U8848 ( .A1(n7057), .A2(n7058), .ZN(n7395) );
  OAI21_X1 U8849 ( .B1(n7058), .B2(n7057), .A(n7395), .ZN(n7059) );
  NAND2_X1 U8850 ( .A1(n7059), .A2(n8951), .ZN(n7066) );
  NAND2_X1 U8851 ( .A1(n9019), .A2(n9035), .ZN(n7060) );
  OAI21_X1 U8852 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7061), .A(n7060), .ZN(n7064) );
  NOR2_X1 U8853 ( .A1(n9021), .A2(n7062), .ZN(n7063) );
  AOI211_X1 U8854 ( .C1(n9007), .C2(n9033), .A(n7064), .B(n7063), .ZN(n7065)
         );
  OAI211_X1 U8855 ( .C1(n4707), .C2(n8958), .A(n7066), .B(n7065), .ZN(P1_U3229) );
  NOR3_X1 U8856 ( .A1(n7151), .A2(n7067), .A3(n7232), .ZN(n7068) );
  AOI21_X1 U8857 ( .B1(n7069), .B2(n10141), .A(n7068), .ZN(n7080) );
  NAND2_X1 U8858 ( .A1(n10137), .A2(n8464), .ZN(n7073) );
  NAND2_X1 U8859 ( .A1(n10136), .A2(n8462), .ZN(n7072) );
  NAND2_X1 U8860 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n8473) );
  INV_X1 U8861 ( .A(n7070), .ZN(n7241) );
  NAND2_X1 U8862 ( .A1(n8210), .A2(n7241), .ZN(n7071) );
  NAND4_X1 U8863 ( .A1(n7073), .A2(n7072), .A3(n8473), .A4(n7071), .ZN(n7077)
         );
  NAND2_X1 U8864 ( .A1(n7075), .A2(n7074), .ZN(n7150) );
  NOR2_X1 U8865 ( .A1(n7150), .A2(n8233), .ZN(n7076) );
  AOI211_X1 U8866 ( .C1(n7421), .C2(n8228), .A(n7077), .B(n7076), .ZN(n7078)
         );
  OAI21_X1 U8867 ( .B1(n7080), .B2(n7079), .A(n7078), .ZN(P2_U3233) );
  AOI21_X1 U8868 ( .B1(n9007), .B2(n9036), .A(n7081), .ZN(n7083) );
  NAND2_X1 U8869 ( .A1(n9019), .A2(n9986), .ZN(n7082) );
  OAI211_X1 U8870 ( .C1(n9021), .C2(n7084), .A(n7083), .B(n7082), .ZN(n7094)
         );
  INV_X1 U8871 ( .A(n7085), .ZN(n7086) );
  NAND2_X1 U8872 ( .A1(n7087), .A2(n7086), .ZN(n7091) );
  NAND2_X1 U8873 ( .A1(n7089), .A2(n7088), .ZN(n7090) );
  XNOR2_X1 U8874 ( .A(n7091), .B(n7090), .ZN(n7092) );
  NOR2_X1 U8875 ( .A1(n7092), .A2(n9025), .ZN(n7093) );
  AOI211_X1 U8876 ( .C1(n9023), .C2(n7095), .A(n7094), .B(n7093), .ZN(n7096)
         );
  INV_X1 U8877 ( .A(n7096), .ZN(P1_U3237) );
  INV_X1 U8878 ( .A(n7097), .ZN(n7116) );
  OAI222_X1 U8879 ( .A1(n8093), .A2(P1_U3084), .B1(n4389), .B2(n7116), .C1(
        n7098), .C2(n9782), .ZN(P1_U3333) );
  NAND2_X1 U8880 ( .A1(n7099), .A2(n10019), .ZN(n7101) );
  AOI22_X1 U8881 ( .A1(n9987), .A2(n9038), .B1(n9037), .B2(n9985), .ZN(n7100)
         );
  NAND2_X1 U8882 ( .A1(n7101), .A2(n7100), .ZN(n10107) );
  INV_X1 U8883 ( .A(n10107), .ZN(n7115) );
  NOR2_X1 U8884 ( .A1(n9387), .A2(n9192), .ZN(n9258) );
  NAND2_X1 U8885 ( .A1(n10001), .A2(n7102), .ZN(n7103) );
  NAND2_X1 U8886 ( .A1(n7103), .A2(n9469), .ZN(n7105) );
  OR2_X1 U8887 ( .A1(n7105), .A2(n7104), .ZN(n10103) );
  INV_X1 U8888 ( .A(n10103), .ZN(n7113) );
  NOR2_X1 U8889 ( .A1(n9994), .A2(n7106), .ZN(n7107) );
  AOI21_X1 U8890 ( .B1(n10021), .B2(P1_REG2_REG_5__SCAN_IN), .A(n7107), .ZN(
        n7108) );
  OAI21_X1 U8891 ( .B1(n10029), .B2(n10105), .A(n7108), .ZN(n7112) );
  NAND2_X1 U8892 ( .A1(n7110), .A2(n7109), .ZN(n10101) );
  AND3_X1 U8893 ( .A1(n10102), .A2(n9363), .A3(n10101), .ZN(n7111) );
  AOI211_X1 U8894 ( .C1(n9258), .C2(n7113), .A(n7112), .B(n7111), .ZN(n7114)
         );
  OAI21_X1 U8895 ( .B1(n10021), .B2(n7115), .A(n7114), .ZN(P1_U3286) );
  OAI222_X1 U8896 ( .A1(n8888), .A2(n9717), .B1(P2_U3152), .B2(n6128), .C1(
        n8883), .C2(n7116), .ZN(P2_U3338) );
  NAND2_X1 U8897 ( .A1(n7117), .A2(n7292), .ZN(n7118) );
  NAND2_X1 U8898 ( .A1(n7118), .A2(n7289), .ZN(n7119) );
  XNOR2_X1 U8899 ( .A(n8850), .B(n8138), .ZN(n7288) );
  NAND2_X1 U8900 ( .A1(n8459), .A2(n6204), .ZN(n7286) );
  XNOR2_X1 U8901 ( .A(n7288), .B(n7286), .ZN(n7297) );
  XNOR2_X1 U8902 ( .A(n7119), .B(n7297), .ZN(n7123) );
  OAI22_X1 U8903 ( .A1(n8240), .A2(n7496), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5950), .ZN(n7121) );
  OAI22_X1 U8904 ( .A1(n7155), .A2(n8224), .B1(n8225), .B2(n7450), .ZN(n7120)
         );
  AOI211_X1 U8905 ( .C1(n8850), .C2(n8228), .A(n7121), .B(n7120), .ZN(n7122)
         );
  OAI21_X1 U8906 ( .B1(n7123), .B2(n8233), .A(n7122), .ZN(P2_U3236) );
  INV_X1 U8907 ( .A(n7124), .ZN(n7160) );
  OAI222_X1 U8908 ( .A1(n8054), .A2(P1_U3084), .B1(n4389), .B2(n7160), .C1(
        n7125), .C2(n9782), .ZN(P1_U3332) );
  NAND2_X1 U8909 ( .A1(n8502), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7129) );
  AOI22_X1 U8910 ( .A1(n8502), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7320), .B2(
        n7126), .ZN(n8498) );
  NAND2_X1 U8911 ( .A1(n8498), .A2(n8499), .ZN(n8497) );
  NAND2_X1 U8912 ( .A1(n7129), .A2(n8497), .ZN(n10161) );
  AOI22_X1 U8913 ( .A1(n10167), .A2(n7497), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7133), .ZN(n10160) );
  NOR2_X1 U8914 ( .A1(n10161), .A2(n10160), .ZN(n10159) );
  INV_X1 U8915 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7130) );
  AOI22_X1 U8916 ( .A1(n7515), .A2(n7130), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7144), .ZN(n7131) );
  NOR2_X1 U8917 ( .A1(n7132), .A2(n7131), .ZN(n7516) );
  AOI21_X1 U8918 ( .B1(n7132), .B2(n7131), .A(n7516), .ZN(n7148) );
  AOI22_X1 U8919 ( .A1(n10167), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n5949), .B2(
        n7133), .ZN(n10165) );
  NAND2_X1 U8920 ( .A1(n7134), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7135) );
  OR2_X1 U8921 ( .A1(n8502), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8922 ( .A1(n8502), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7137) );
  AND2_X1 U8923 ( .A1(n7138), .A2(n7137), .ZN(n8504) );
  NAND2_X1 U8924 ( .A1(n8505), .A2(n8504), .ZN(n8503) );
  OAI21_X1 U8925 ( .B1(n8502), .B2(P2_REG1_REG_12__SCAN_IN), .A(n8503), .ZN(
        n10164) );
  NAND2_X1 U8926 ( .A1(n10165), .A2(n10164), .ZN(n10163) );
  OAI21_X1 U8927 ( .B1(n10167), .B2(P2_REG1_REG_13__SCAN_IN), .A(n10163), .ZN(
        n7142) );
  NOR2_X1 U8928 ( .A1(n7144), .A2(n7139), .ZN(n7140) );
  AOI21_X1 U8929 ( .B1(n7139), .B2(n7144), .A(n7140), .ZN(n7141) );
  NAND2_X1 U8930 ( .A1(n7141), .A2(n7142), .ZN(n7506) );
  OAI21_X1 U8931 ( .B1(n7142), .B2(n7141), .A(n7506), .ZN(n7146) );
  NOR2_X1 U8932 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9683), .ZN(n7306) );
  AOI21_X1 U8933 ( .B1(n10162), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n7306), .ZN(
        n7143) );
  OAI21_X1 U8934 ( .B1(n10152), .B2(n7144), .A(n7143), .ZN(n7145) );
  AOI21_X1 U8935 ( .B1(n7146), .B2(n10168), .A(n7145), .ZN(n7147) );
  OAI21_X1 U8936 ( .B1(n7148), .B2(n10172), .A(n7147), .ZN(P2_U3259) );
  NAND2_X1 U8937 ( .A1(n7150), .A2(n7149), .ZN(n7260) );
  OR2_X1 U8938 ( .A1(n7260), .A2(n7261), .ZN(n7258) );
  AOI21_X1 U8939 ( .B1(n7258), .B2(n7037), .A(n8233), .ZN(n7154) );
  NOR3_X1 U8940 ( .A1(n7152), .A2(n7231), .A3(n7151), .ZN(n7153) );
  OAI21_X1 U8941 ( .B1(n7154), .B2(n7153), .A(n7295), .ZN(n7159) );
  OAI22_X1 U8942 ( .A1(n8240), .A2(n7224), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5922), .ZN(n7157) );
  OAI22_X1 U8943 ( .A1(n7155), .A2(n8225), .B1(n8224), .B2(n7231), .ZN(n7156)
         );
  AOI211_X1 U8944 ( .C1(n7367), .C2(n8228), .A(n7157), .B(n7156), .ZN(n7158)
         );
  NAND2_X1 U8945 ( .A1(n7159), .A2(n7158), .ZN(P2_U3238) );
  OAI222_X1 U8946 ( .A1(n8888), .A2(n7161), .B1(P2_U3152), .B2(n8436), .C1(
        n8883), .C2(n7160), .ZN(P2_U3337) );
  NAND2_X1 U8947 ( .A1(n7326), .A2(n6674), .ZN(n7163) );
  NAND2_X1 U8948 ( .A1(n9033), .A2(n4388), .ZN(n7162) );
  NAND2_X1 U8949 ( .A1(n7163), .A2(n7162), .ZN(n7164) );
  AND2_X1 U8950 ( .A1(n7634), .A2(n9033), .ZN(n7165) );
  AOI21_X1 U8951 ( .B1(n7326), .B2(n4386), .A(n7165), .ZN(n7385) );
  XNOR2_X1 U8952 ( .A(n7387), .B(n7385), .ZN(n7397) );
  INV_X1 U8953 ( .A(n7166), .ZN(n7168) );
  NAND2_X1 U8954 ( .A1(n7168), .A2(n7167), .ZN(n7388) );
  NAND2_X1 U8955 ( .A1(n7395), .A2(n7388), .ZN(n7169) );
  XOR2_X1 U8956 ( .A(n7397), .B(n7169), .Z(n7175) );
  AOI21_X1 U8957 ( .B1(n9019), .B2(n9034), .A(n7170), .ZN(n7172) );
  NAND2_X1 U8958 ( .A1(n9007), .A2(n9032), .ZN(n7171) );
  OAI211_X1 U8959 ( .C1(n9021), .C2(n7327), .A(n7172), .B(n7171), .ZN(n7173)
         );
  AOI21_X1 U8960 ( .B1(n9023), .B2(n7326), .A(n7173), .ZN(n7174) );
  OAI21_X1 U8961 ( .B1(n7175), .B2(n9025), .A(n7174), .ZN(P1_U3215) );
  NAND2_X1 U8962 ( .A1(n7176), .A2(n8411), .ZN(n7177) );
  NAND2_X1 U8963 ( .A1(n7178), .A2(n7177), .ZN(n10287) );
  INV_X1 U8964 ( .A(n7179), .ZN(n7180) );
  AND2_X1 U8965 ( .A1(n10222), .A2(n7180), .ZN(n8760) );
  INV_X1 U8966 ( .A(n8760), .ZN(n8736) );
  AOI21_X1 U8967 ( .B1(n7181), .B2(n5914), .A(n6148), .ZN(n7185) );
  NAND2_X1 U8968 ( .A1(n8463), .A2(n10189), .ZN(n7183) );
  NAND2_X1 U8969 ( .A1(n8461), .A2(n10190), .ZN(n7182) );
  NAND2_X1 U8970 ( .A1(n7183), .A2(n7182), .ZN(n7255) );
  AOI21_X1 U8971 ( .B1(n7185), .B2(n7184), .A(n7255), .ZN(n7186) );
  OAI21_X1 U8972 ( .B1(n10287), .B2(n8741), .A(n7186), .ZN(n10290) );
  NAND2_X1 U8973 ( .A1(n10290), .A2(n10222), .ZN(n7193) );
  OAI22_X1 U8974 ( .A1(n10222), .A2(n7187), .B1(n7257), .B2(n10218), .ZN(n7191) );
  INV_X1 U8975 ( .A(n7264), .ZN(n10288) );
  INV_X1 U8976 ( .A(n7188), .ZN(n7239) );
  INV_X1 U8977 ( .A(n7189), .ZN(n7223) );
  OAI21_X1 U8978 ( .B1(n10288), .B2(n7239), .A(n7223), .ZN(n10289) );
  NOR2_X1 U8979 ( .A1(n10289), .A2(n10219), .ZN(n7190) );
  AOI211_X1 U8980 ( .C1(n10183), .C2(n7264), .A(n7191), .B(n7190), .ZN(n7192)
         );
  OAI211_X1 U8981 ( .C1(n10287), .C2(n8736), .A(n7193), .B(n7192), .ZN(
        P2_U3286) );
  INV_X1 U8982 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7201) );
  INV_X1 U8983 ( .A(n7194), .ZN(n7199) );
  AOI22_X1 U8984 ( .A1(n7196), .A2(n9469), .B1(n9822), .B2(n7195), .ZN(n7197)
         );
  OAI211_X1 U8985 ( .C1(n9473), .C2(n7199), .A(n7198), .B(n7197), .ZN(n7202)
         );
  NAND2_X1 U8986 ( .A1(n7202), .A2(n10126), .ZN(n7200) );
  OAI21_X1 U8987 ( .B1(n10126), .B2(n7201), .A(n7200), .ZN(P1_U3481) );
  NAND2_X1 U8988 ( .A1(n7202), .A2(n4387), .ZN(n7203) );
  OAI21_X1 U8989 ( .B1(n4387), .B2(n5284), .A(n7203), .ZN(P1_U3532) );
  INV_X1 U8990 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7216) );
  INV_X1 U8991 ( .A(n7205), .ZN(n7206) );
  AOI21_X1 U8992 ( .B1(n4807), .B2(n7204), .A(n7206), .ZN(n7336) );
  AOI21_X1 U8993 ( .B1(n7207), .B2(n8039), .A(n9989), .ZN(n7210) );
  OAI22_X1 U8994 ( .A1(n7435), .A2(n10010), .B1(n9966), .B2(n10012), .ZN(n7208) );
  AOI21_X1 U8995 ( .B1(n7210), .B2(n7209), .A(n7208), .ZN(n7331) );
  NAND2_X1 U8996 ( .A1(n7211), .A2(n7326), .ZN(n7212) );
  NAND2_X1 U8997 ( .A1(n7212), .A2(n9469), .ZN(n7213) );
  NOR2_X1 U8998 ( .A1(n7272), .A2(n7213), .ZN(n7334) );
  AOI21_X1 U8999 ( .B1(n9822), .B2(n7326), .A(n7334), .ZN(n7214) );
  OAI211_X1 U9000 ( .C1(n7336), .C2(n9823), .A(n7331), .B(n7214), .ZN(n7217)
         );
  NAND2_X1 U9001 ( .A1(n7217), .A2(n10126), .ZN(n7215) );
  OAI21_X1 U9002 ( .B1(n10126), .B2(n7216), .A(n7215), .ZN(P1_U3484) );
  NAND2_X1 U9003 ( .A1(n7217), .A2(n4387), .ZN(n7218) );
  OAI21_X1 U9004 ( .B1(n4387), .B2(n5302), .A(n7218), .ZN(P1_U3533) );
  XNOR2_X1 U9005 ( .A(n7219), .B(n8414), .ZN(n7371) );
  XNOR2_X1 U9006 ( .A(n7220), .B(n8414), .ZN(n7221) );
  AOI222_X1 U9007 ( .A1(n10193), .A2(n7221), .B1(n8462), .B2(n10189), .C1(
        n8460), .C2(n10190), .ZN(n7370) );
  OR2_X1 U9008 ( .A1(n7370), .A2(n10224), .ZN(n7229) );
  INV_X1 U9009 ( .A(n7317), .ZN(n7222) );
  AOI21_X1 U9010 ( .B1(n7367), .B2(n7223), .A(n7222), .ZN(n7368) );
  OAI22_X1 U9011 ( .A1(n10218), .A2(n7224), .B1(n5925), .B2(n10222), .ZN(n7227) );
  NOR2_X1 U9012 ( .A1(n7225), .A2(n10200), .ZN(n7226) );
  AOI211_X1 U9013 ( .C1(n7368), .C2(n8711), .A(n7227), .B(n7226), .ZN(n7228)
         );
  OAI211_X1 U9014 ( .C1(n7371), .C2(n8713), .A(n7229), .B(n7228), .ZN(P2_U3285) );
  XNOR2_X1 U9015 ( .A(n7230), .B(n8410), .ZN(n7238) );
  OAI22_X1 U9016 ( .A1(n7232), .A2(n10210), .B1(n7231), .B2(n10211), .ZN(n7237) );
  INV_X1 U9017 ( .A(n7233), .ZN(n7234) );
  AOI21_X1 U9018 ( .B1(n8410), .B2(n7235), .A(n7234), .ZN(n7425) );
  NOR2_X1 U9019 ( .A1(n7425), .A2(n8741), .ZN(n7236) );
  AOI211_X1 U9020 ( .C1(n7238), .C2(n10193), .A(n7237), .B(n7236), .ZN(n7424)
         );
  AOI21_X1 U9021 ( .B1(n7421), .B2(n7240), .A(n7239), .ZN(n7422) );
  INV_X1 U9022 ( .A(n10218), .ZN(n8698) );
  AOI22_X1 U9023 ( .A1(n10224), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n7241), .B2(
        n8698), .ZN(n7242) );
  OAI21_X1 U9024 ( .B1(n4736), .B2(n10200), .A(n7242), .ZN(n7244) );
  NOR2_X1 U9025 ( .A1(n7425), .A2(n8736), .ZN(n7243) );
  AOI211_X1 U9026 ( .C1(n7422), .C2(n8711), .A(n7244), .B(n7243), .ZN(n7245)
         );
  OAI21_X1 U9027 ( .B1(n7424), .B2(n10224), .A(n7245), .ZN(P2_U3287) );
  AOI22_X1 U9028 ( .A1(n10224), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7246), .B2(
        n8698), .ZN(n7247) );
  OAI21_X1 U9029 ( .B1(n7248), .B2(n10200), .A(n7247), .ZN(n7251) );
  NOR2_X1 U9030 ( .A1(n7249), .A2(n10224), .ZN(n7250) );
  AOI211_X1 U9031 ( .C1(n7252), .C2(n8711), .A(n7251), .B(n7250), .ZN(n7253)
         );
  OAI21_X1 U9032 ( .B1(n8713), .B2(n7254), .A(n7253), .ZN(P2_U3289) );
  AOI22_X1 U9033 ( .A1(n8242), .A2(n7255), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7256) );
  OAI21_X1 U9034 ( .B1(n7257), .B2(n8240), .A(n7256), .ZN(n7263) );
  INV_X1 U9035 ( .A(n7258), .ZN(n7259) );
  AOI211_X1 U9036 ( .C1(n7261), .C2(n7260), .A(n8233), .B(n7259), .ZN(n7262)
         );
  AOI211_X1 U9037 ( .C1(n7264), .C2(n8228), .A(n7263), .B(n7262), .ZN(n7265)
         );
  INV_X1 U9038 ( .A(n7265), .ZN(P2_U3219) );
  OAI21_X1 U9039 ( .B1(n7267), .B2(n8040), .A(n7266), .ZN(n9467) );
  XNOR2_X1 U9040 ( .A(n7268), .B(n7837), .ZN(n7270) );
  AOI22_X1 U9041 ( .A1(n9985), .A2(n9031), .B1(n9033), .B2(n9987), .ZN(n7269)
         );
  OAI21_X1 U9042 ( .B1(n7270), .B2(n9989), .A(n7269), .ZN(n7271) );
  AOI21_X1 U9043 ( .B1(n9992), .B2(n9467), .A(n7271), .ZN(n9472) );
  INV_X1 U9044 ( .A(n7272), .ZN(n7274) );
  INV_X1 U9045 ( .A(n7436), .ZN(n7273) );
  AOI21_X1 U9046 ( .B1(n9468), .B2(n7274), .A(n7273), .ZN(n9470) );
  NOR2_X1 U9047 ( .A1(n7275), .A2(n10029), .ZN(n7278) );
  OAI22_X1 U9048 ( .A1(n9321), .A2(n7276), .B1(n8990), .B2(n9994), .ZN(n7277)
         );
  AOI211_X1 U9049 ( .C1(n9470), .C2(n10003), .A(n7278), .B(n7277), .ZN(n7280)
         );
  NAND2_X1 U9050 ( .A1(n9467), .A2(n10004), .ZN(n7279) );
  OAI211_X1 U9051 ( .C1(n9472), .C2(n9387), .A(n7280), .B(n7279), .ZN(P1_U3280) );
  XNOR2_X1 U9052 ( .A(n7484), .B(n6201), .ZN(n7281) );
  NAND2_X1 U9053 ( .A1(n8458), .A2(n6204), .ZN(n7282) );
  NAND2_X1 U9054 ( .A1(n7281), .A2(n7282), .ZN(n7446) );
  INV_X1 U9055 ( .A(n7281), .ZN(n7284) );
  INV_X1 U9056 ( .A(n7282), .ZN(n7283) );
  NAND2_X1 U9057 ( .A1(n7284), .A2(n7283), .ZN(n7285) );
  NAND2_X1 U9058 ( .A1(n7446), .A2(n7285), .ZN(n7303) );
  INV_X1 U9059 ( .A(n7286), .ZN(n7287) );
  NAND2_X1 U9060 ( .A1(n7288), .A2(n7287), .ZN(n7296) );
  AND2_X1 U9061 ( .A1(n7289), .A2(n7296), .ZN(n7291) );
  AND2_X1 U9062 ( .A1(n7290), .A2(n7291), .ZN(n7294) );
  INV_X1 U9063 ( .A(n7291), .ZN(n7293) );
  AOI21_X1 U9064 ( .B1(n7295), .B2(n7294), .A(n5049), .ZN(n7300) );
  INV_X1 U9065 ( .A(n7296), .ZN(n7298) );
  OR2_X1 U9066 ( .A1(n7298), .A2(n7297), .ZN(n7299) );
  INV_X1 U9067 ( .A(n7447), .ZN(n7301) );
  AOI21_X1 U9068 ( .B1(n7303), .B2(n7302), .A(n7301), .ZN(n7310) );
  INV_X1 U9069 ( .A(n7482), .ZN(n7307) );
  OAI22_X1 U9070 ( .A1(n8336), .A2(n8225), .B1(n8224), .B2(n7304), .ZN(n7305)
         );
  AOI211_X1 U9071 ( .C1(n8210), .C2(n7307), .A(n7306), .B(n7305), .ZN(n7309)
         );
  NAND2_X1 U9072 ( .A1(n7484), .A2(n8228), .ZN(n7308) );
  OAI211_X1 U9073 ( .C1(n7310), .C2(n8233), .A(n7309), .B(n7308), .ZN(P2_U3217) );
  XNOR2_X1 U9074 ( .A(n7311), .B(n7312), .ZN(n10303) );
  INV_X1 U9075 ( .A(n10303), .ZN(n7325) );
  INV_X1 U9076 ( .A(n7312), .ZN(n8415) );
  XNOR2_X1 U9077 ( .A(n7313), .B(n8415), .ZN(n7314) );
  NAND2_X1 U9078 ( .A1(n7314), .A2(n10193), .ZN(n7316) );
  NAND2_X1 U9079 ( .A1(n7316), .A2(n7315), .ZN(n10300) );
  NAND2_X1 U9080 ( .A1(n7317), .A2(n10295), .ZN(n7318) );
  NAND2_X1 U9081 ( .A1(n7499), .A2(n7318), .ZN(n10299) );
  OAI22_X1 U9082 ( .A1(n10222), .A2(n7320), .B1(n7319), .B2(n10218), .ZN(n7321) );
  AOI21_X1 U9083 ( .B1(n10295), .B2(n10183), .A(n7321), .ZN(n7322) );
  OAI21_X1 U9084 ( .B1(n10299), .B2(n10219), .A(n7322), .ZN(n7323) );
  AOI21_X1 U9085 ( .B1(n10300), .B2(n10222), .A(n7323), .ZN(n7324) );
  OAI21_X1 U9086 ( .B1(n7325), .B2(n8713), .A(n7324), .ZN(P2_U3284) );
  INV_X1 U9087 ( .A(n7326), .ZN(n7330) );
  INV_X1 U9088 ( .A(n7327), .ZN(n7328) );
  AOI22_X1 U9089 ( .A1(n9387), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7328), .B2(
        n10020), .ZN(n7329) );
  OAI21_X1 U9090 ( .B1(n10029), .B2(n7330), .A(n7329), .ZN(n7333) );
  NOR2_X1 U9091 ( .A1(n7331), .A2(n9387), .ZN(n7332) );
  AOI211_X1 U9092 ( .C1(n7334), .C2(n7438), .A(n7333), .B(n7332), .ZN(n7335)
         );
  OAI21_X1 U9093 ( .B1(n9323), .B2(n7336), .A(n7335), .ZN(P1_U3281) );
  INV_X1 U9094 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10354) );
  NOR2_X1 U9095 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7337) );
  AOI21_X1 U9096 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7337), .ZN(n10326) );
  NOR2_X1 U9097 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7338) );
  AOI21_X1 U9098 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7338), .ZN(n10329) );
  NOR2_X1 U9099 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n7339) );
  AOI21_X1 U9100 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n7339), .ZN(n10332) );
  NOR2_X1 U9101 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7340) );
  AOI21_X1 U9102 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7340), .ZN(n10335) );
  NOR2_X1 U9103 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .ZN(n7341) );
  AOI21_X1 U9104 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n7341), .ZN(n10338) );
  NOR2_X1 U9105 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7347) );
  XNOR2_X1 U9106 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10366) );
  NAND2_X1 U9107 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7345) );
  XOR2_X1 U9108 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10364) );
  NAND2_X1 U9109 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7343) );
  XOR2_X1 U9110 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10362) );
  AOI21_X1 U9111 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10320) );
  INV_X1 U9112 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9787) );
  NAND3_X1 U9113 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10322) );
  OAI21_X1 U9114 ( .B1(n10320), .B2(n9787), .A(n10322), .ZN(n10361) );
  NAND2_X1 U9115 ( .A1(n10362), .A2(n10361), .ZN(n7342) );
  NAND2_X1 U9116 ( .A1(n7343), .A2(n7342), .ZN(n10363) );
  NAND2_X1 U9117 ( .A1(n10364), .A2(n10363), .ZN(n7344) );
  NAND2_X1 U9118 ( .A1(n7345), .A2(n7344), .ZN(n10365) );
  NOR2_X1 U9119 ( .A1(n10366), .A2(n10365), .ZN(n7346) );
  NOR2_X1 U9120 ( .A1(n7347), .A2(n7346), .ZN(n7348) );
  NOR2_X1 U9121 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7348), .ZN(n10350) );
  AND2_X1 U9122 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7348), .ZN(n10349) );
  NOR2_X1 U9123 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10349), .ZN(n7349) );
  NOR2_X1 U9124 ( .A1(n10350), .A2(n7349), .ZN(n7350) );
  NAND2_X1 U9125 ( .A1(n7350), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7352) );
  XOR2_X1 U9126 ( .A(n7350), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10348) );
  NAND2_X1 U9127 ( .A1(n10348), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7351) );
  NAND2_X1 U9128 ( .A1(n7352), .A2(n7351), .ZN(n7353) );
  NAND2_X1 U9129 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7353), .ZN(n7355) );
  XOR2_X1 U9130 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n7353), .Z(n10360) );
  NAND2_X1 U9131 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10360), .ZN(n7354) );
  NAND2_X1 U9132 ( .A1(n7355), .A2(n7354), .ZN(n7356) );
  NAND2_X1 U9133 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7356), .ZN(n7358) );
  XOR2_X1 U9134 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7356), .Z(n10359) );
  NAND2_X1 U9135 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10359), .ZN(n7357) );
  NAND2_X1 U9136 ( .A1(n7358), .A2(n7357), .ZN(n7359) );
  AND2_X1 U9137 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7359), .ZN(n7360) );
  INV_X1 U9138 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10358) );
  XNOR2_X1 U9139 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7359), .ZN(n10357) );
  NOR2_X1 U9140 ( .A1(n10358), .A2(n10357), .ZN(n10356) );
  NAND2_X1 U9141 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7361) );
  OAI21_X1 U9142 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7361), .ZN(n10346) );
  AOI21_X1 U9143 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10345), .ZN(n10344) );
  NAND2_X1 U9144 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7362) );
  OAI21_X1 U9145 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7362), .ZN(n10343) );
  NOR2_X1 U9146 ( .A1(n10344), .A2(n10343), .ZN(n10342) );
  AOI21_X1 U9147 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10342), .ZN(n10341) );
  NOR2_X1 U9148 ( .A1(P1_ADDR_REG_12__SCAN_IN), .A2(P2_ADDR_REG_12__SCAN_IN), 
        .ZN(n7363) );
  AOI21_X1 U9149 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n7363), .ZN(n10340) );
  NAND2_X1 U9150 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  OAI21_X1 U9151 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n10339), .ZN(n10337) );
  NAND2_X1 U9152 ( .A1(n10338), .A2(n10337), .ZN(n10336) );
  OAI21_X1 U9153 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10336), .ZN(n10334) );
  NAND2_X1 U9154 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  OAI21_X1 U9155 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10333), .ZN(n10331) );
  NAND2_X1 U9156 ( .A1(n10332), .A2(n10331), .ZN(n10330) );
  OAI21_X1 U9157 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10330), .ZN(n10328) );
  NAND2_X1 U9158 ( .A1(n10329), .A2(n10328), .ZN(n10327) );
  OAI21_X1 U9159 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10327), .ZN(n10325) );
  NAND2_X1 U9160 ( .A1(n10326), .A2(n10325), .ZN(n10324) );
  OAI21_X1 U9161 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10324), .ZN(n10353) );
  NOR2_X1 U9162 ( .A1(n10354), .A2(n10353), .ZN(n7364) );
  NAND2_X1 U9163 ( .A1(n10354), .A2(n10353), .ZN(n10352) );
  OAI21_X1 U9164 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7364), .A(n10352), .ZN(
        n7366) );
  XNOR2_X1 U9165 ( .A(n4511), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7365) );
  XNOR2_X1 U9166 ( .A(n7366), .B(n7365), .ZN(ADD_1071_U4) );
  AOI22_X1 U9167 ( .A1(n7368), .A2(n8852), .B1(n8851), .B2(n7367), .ZN(n7369)
         );
  OAI211_X1 U9168 ( .C1(n8848), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7374)
         );
  NAND2_X1 U9169 ( .A1(n7374), .A2(n10319), .ZN(n7372) );
  OAI21_X1 U9170 ( .B1(n10319), .B2(n7373), .A(n7372), .ZN(P2_U3531) );
  NAND2_X1 U9171 ( .A1(n7374), .A2(n10306), .ZN(n7375) );
  OAI21_X1 U9172 ( .B1(n10306), .B2(n5926), .A(n7375), .ZN(P2_U3484) );
  NAND2_X1 U9173 ( .A1(n9464), .A2(n6674), .ZN(n7377) );
  NAND2_X1 U9174 ( .A1(n9031), .A2(n4388), .ZN(n7376) );
  NAND2_X1 U9175 ( .A1(n7377), .A2(n7376), .ZN(n7378) );
  XNOR2_X1 U9176 ( .A(n7378), .B(n7770), .ZN(n7380) );
  AND2_X1 U9177 ( .A1(n7634), .A2(n9031), .ZN(n7379) );
  AOI21_X1 U9178 ( .B1(n9464), .B2(n4386), .A(n7379), .ZN(n7381) );
  NAND2_X1 U9179 ( .A1(n7380), .A2(n7381), .ZN(n7467) );
  INV_X1 U9180 ( .A(n7380), .ZN(n7383) );
  INV_X1 U9181 ( .A(n7381), .ZN(n7382) );
  NAND2_X1 U9182 ( .A1(n7383), .A2(n7382), .ZN(n7384) );
  NAND2_X1 U9183 ( .A1(n7467), .A2(n7384), .ZN(n7406) );
  AND2_X1 U9184 ( .A1(n7388), .A2(n7396), .ZN(n8991) );
  NAND2_X1 U9185 ( .A1(n9468), .A2(n6674), .ZN(n7390) );
  NAND2_X1 U9186 ( .A1(n9032), .A2(n4388), .ZN(n7389) );
  NAND2_X1 U9187 ( .A1(n7390), .A2(n7389), .ZN(n7391) );
  XNOR2_X1 U9188 ( .A(n7391), .B(n7770), .ZN(n8994) );
  AND2_X1 U9189 ( .A1(n7634), .A2(n9032), .ZN(n7392) );
  AOI21_X1 U9190 ( .B1(n9468), .B2(n4388), .A(n7392), .ZN(n8993) );
  AND2_X1 U9191 ( .A1(n8994), .A2(n8993), .ZN(n7399) );
  INV_X1 U9192 ( .A(n7399), .ZN(n7393) );
  AND2_X1 U9193 ( .A1(n8991), .A2(n7393), .ZN(n7394) );
  INV_X1 U9194 ( .A(n7396), .ZN(n7398) );
  OR2_X1 U9195 ( .A1(n7398), .A2(n7397), .ZN(n8992) );
  INV_X1 U9196 ( .A(n8994), .ZN(n7401) );
  INV_X1 U9197 ( .A(n8993), .ZN(n7400) );
  INV_X1 U9198 ( .A(n7468), .ZN(n7404) );
  AOI21_X1 U9199 ( .B1(n7406), .B2(n7405), .A(n7404), .ZN(n7413) );
  INV_X1 U9200 ( .A(n7407), .ZN(n7409) );
  NOR2_X1 U9201 ( .A1(n9005), .A2(n7435), .ZN(n7408) );
  AOI211_X1 U9202 ( .C1(n9007), .C2(n9030), .A(n7409), .B(n7408), .ZN(n7410)
         );
  OAI21_X1 U9203 ( .B1(n9021), .B2(n7440), .A(n7410), .ZN(n7411) );
  AOI21_X1 U9204 ( .B1(n9023), .B2(n9464), .A(n7411), .ZN(n7412) );
  OAI21_X1 U9205 ( .B1(n7413), .B2(n9025), .A(n7412), .ZN(P1_U3222) );
  INV_X1 U9206 ( .A(n7414), .ZN(n7612) );
  OAI222_X1 U9207 ( .A1(P1_U3084), .A2(n7934), .B1(n4389), .B2(n7612), .C1(
        n9583), .C2(n9782), .ZN(P1_U3331) );
  NAND2_X1 U9208 ( .A1(n7417), .A2(n8884), .ZN(n7415) );
  OAI211_X1 U9209 ( .C1(n7416), .C2(n8888), .A(n7415), .B(n8451), .ZN(P2_U3335) );
  NAND2_X1 U9210 ( .A1(n7417), .A2(n9777), .ZN(n7419) );
  NOR2_X1 U9211 ( .A1(n7418), .A2(P1_U3084), .ZN(n8096) );
  INV_X1 U9212 ( .A(n8096), .ZN(n8100) );
  OAI211_X1 U9213 ( .C1(n7420), .C2(n9782), .A(n7419), .B(n8100), .ZN(P1_U3330) );
  INV_X1 U9214 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7427) );
  INV_X1 U9215 ( .A(n10293), .ZN(n8855) );
  AOI22_X1 U9216 ( .A1(n7422), .A2(n8852), .B1(n8851), .B2(n7421), .ZN(n7423)
         );
  OAI211_X1 U9217 ( .C1(n7425), .C2(n8855), .A(n7424), .B(n7423), .ZN(n7428)
         );
  NAND2_X1 U9218 ( .A1(n7428), .A2(n10306), .ZN(n7426) );
  OAI21_X1 U9219 ( .B1(n10306), .B2(n7427), .A(n7426), .ZN(P2_U3478) );
  NAND2_X1 U9220 ( .A1(n7428), .A2(n10319), .ZN(n7429) );
  OAI21_X1 U9221 ( .B1(n10319), .B2(n6663), .A(n7429), .ZN(P2_U3529) );
  XNOR2_X1 U9222 ( .A(n7430), .B(n9369), .ZN(n9466) );
  NAND2_X1 U9223 ( .A1(n7432), .A2(n7431), .ZN(n7433) );
  XOR2_X1 U9224 ( .A(n9369), .B(n7433), .Z(n7434) );
  OAI222_X1 U9225 ( .A1(n10010), .A2(n9356), .B1(n10012), .B2(n7435), .C1(
        n9989), .C2(n7434), .ZN(n9462) );
  AOI21_X1 U9226 ( .B1(n7436), .B2(n9464), .A(n10118), .ZN(n7437) );
  AND2_X1 U9227 ( .A1(n7437), .A2(n9377), .ZN(n9463) );
  NAND2_X1 U9228 ( .A1(n9463), .A2(n7438), .ZN(n7443) );
  NAND2_X1 U9229 ( .A1(n10021), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7439) );
  OAI21_X1 U9230 ( .B1(n9994), .B2(n7440), .A(n7439), .ZN(n7441) );
  AOI21_X1 U9231 ( .B1(n9464), .B2(n9350), .A(n7441), .ZN(n7442) );
  NAND2_X1 U9232 ( .A1(n7443), .A2(n7442), .ZN(n7444) );
  AOI21_X1 U9233 ( .B1(n9462), .B2(n9321), .A(n7444), .ZN(n7445) );
  OAI21_X1 U9234 ( .B1(n9323), .B2(n9466), .A(n7445), .ZN(P1_U3279) );
  NAND2_X1 U9235 ( .A1(n8229), .A2(n8743), .ZN(n7449) );
  AND2_X1 U9236 ( .A1(n8743), .A2(n6204), .ZN(n7532) );
  OR2_X1 U9237 ( .A1(n8233), .A2(n7532), .ZN(n7448) );
  XNOR2_X1 U9238 ( .A(n8844), .B(n8138), .ZN(n7534) );
  MUX2_X1 U9239 ( .A(n7449), .B(n7448), .S(n7533), .Z(n7454) );
  OAI22_X1 U9240 ( .A1(n8240), .A2(n7558), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5973), .ZN(n7452) );
  OAI22_X1 U9241 ( .A1(n7450), .A2(n8224), .B1(n8225), .B2(n7566), .ZN(n7451)
         );
  AOI211_X1 U9242 ( .C1(n8844), .C2(n8228), .A(n7452), .B(n7451), .ZN(n7453)
         );
  NAND2_X1 U9243 ( .A1(n7454), .A2(n7453), .ZN(P2_U3243) );
  INV_X1 U9244 ( .A(n7455), .ZN(n7458) );
  INV_X1 U9245 ( .A(n7456), .ZN(n7732) );
  OAI222_X1 U9246 ( .A1(n7458), .A2(P2_U3152), .B1(n8883), .B2(n7732), .C1(
        n7457), .C2(n8888), .ZN(P2_U3334) );
  NAND2_X1 U9247 ( .A1(n9457), .A2(n6674), .ZN(n7460) );
  NAND2_X1 U9248 ( .A1(n9030), .A2(n4386), .ZN(n7459) );
  NAND2_X1 U9249 ( .A1(n7460), .A2(n7459), .ZN(n7461) );
  XNOR2_X1 U9250 ( .A(n7461), .B(n7770), .ZN(n7463) );
  AND2_X1 U9251 ( .A1(n7634), .A2(n9030), .ZN(n7462) );
  AOI21_X1 U9252 ( .B1(n9457), .B2(n4391), .A(n7462), .ZN(n7464) );
  NAND2_X1 U9253 ( .A1(n7463), .A2(n7464), .ZN(n7621) );
  INV_X1 U9254 ( .A(n7463), .ZN(n7466) );
  INV_X1 U9255 ( .A(n7464), .ZN(n7465) );
  NAND2_X1 U9256 ( .A1(n7466), .A2(n7465), .ZN(n7623) );
  NAND2_X1 U9257 ( .A1(n7621), .A2(n7623), .ZN(n7469) );
  XOR2_X1 U9258 ( .A(n7469), .B(n7622), .Z(n7475) );
  NOR2_X1 U9259 ( .A1(n9017), .A2(n9368), .ZN(n7470) );
  AOI211_X1 U9260 ( .C1(n9019), .C2(n9031), .A(n7471), .B(n7470), .ZN(n7472)
         );
  OAI21_X1 U9261 ( .B1(n9021), .B2(n9380), .A(n7472), .ZN(n7473) );
  AOI21_X1 U9262 ( .B1(n9023), .B2(n9457), .A(n7473), .ZN(n7474) );
  OAI21_X1 U9263 ( .B1(n7475), .B2(n9025), .A(n7474), .ZN(P1_U3232) );
  XNOR2_X1 U9264 ( .A(n7476), .B(n8419), .ZN(n9814) );
  INV_X1 U9265 ( .A(n9814), .ZN(n7488) );
  OAI211_X1 U9266 ( .C1(n7478), .C2(n8419), .A(n7477), .B(n10193), .ZN(n7480)
         );
  AOI22_X1 U9267 ( .A1(n10190), .A2(n8743), .B1(n8459), .B2(n10189), .ZN(n7479) );
  NAND2_X1 U9268 ( .A1(n7480), .A2(n7479), .ZN(n9812) );
  INV_X1 U9269 ( .A(n7556), .ZN(n7481) );
  OAI21_X1 U9270 ( .B1(n9810), .B2(n7501), .A(n7481), .ZN(n9811) );
  OAI22_X1 U9271 ( .A1(n10222), .A2(n7130), .B1(n7482), .B2(n10218), .ZN(n7483) );
  AOI21_X1 U9272 ( .B1(n7484), .B2(n10183), .A(n7483), .ZN(n7485) );
  OAI21_X1 U9273 ( .B1(n9811), .B2(n10219), .A(n7485), .ZN(n7486) );
  AOI21_X1 U9274 ( .B1(n9812), .B2(n10222), .A(n7486), .ZN(n7487) );
  OAI21_X1 U9275 ( .B1(n7488), .B2(n8713), .A(n7487), .ZN(P2_U3282) );
  NAND2_X1 U9276 ( .A1(n7489), .A2(n8328), .ZN(n7490) );
  NAND2_X1 U9277 ( .A1(n7491), .A2(n7490), .ZN(n8856) );
  AOI22_X1 U9278 ( .A1(n10189), .A2(n8460), .B1(n8458), .B2(n10190), .ZN(n7495) );
  XNOR2_X1 U9279 ( .A(n7492), .B(n8328), .ZN(n7493) );
  NAND2_X1 U9280 ( .A1(n7493), .A2(n10193), .ZN(n7494) );
  OAI211_X1 U9281 ( .C1(n8856), .C2(n8741), .A(n7495), .B(n7494), .ZN(n8858)
         );
  OAI22_X1 U9282 ( .A1(n10222), .A2(n7497), .B1(n7496), .B2(n10218), .ZN(n7498) );
  AOI21_X1 U9283 ( .B1(n8850), .B2(n10183), .A(n7498), .ZN(n7503) );
  AND2_X1 U9284 ( .A1(n7499), .A2(n8850), .ZN(n7500) );
  NOR2_X1 U9285 ( .A1(n7501), .A2(n7500), .ZN(n8853) );
  NAND2_X1 U9286 ( .A1(n8853), .A2(n8711), .ZN(n7502) );
  OAI211_X1 U9287 ( .C1(n8856), .C2(n8736), .A(n7503), .B(n7502), .ZN(n7504)
         );
  AOI21_X1 U9288 ( .B1(n8858), .B2(n10222), .A(n7504), .ZN(n7505) );
  INV_X1 U9289 ( .A(n7505), .ZN(P2_U3283) );
  OAI21_X1 U9290 ( .B1(n7515), .B2(P2_REG1_REG_14__SCAN_IN), .A(n7506), .ZN(
        n7507) );
  XNOR2_X1 U9291 ( .A(n7507), .B(n8515), .ZN(n8517) );
  NAND2_X1 U9292 ( .A1(n8517), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8516) );
  OR2_X1 U9293 ( .A1(n7520), .A2(n7507), .ZN(n7508) );
  XNOR2_X1 U9294 ( .A(n7747), .B(n7509), .ZN(n7510) );
  NAND2_X1 U9295 ( .A1(n7510), .A2(n7511), .ZN(n7746) );
  OAI21_X1 U9296 ( .B1(n7511), .B2(n7510), .A(n7746), .ZN(n7514) );
  INV_X1 U9297 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U9298 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7539) );
  OAI21_X1 U9299 ( .B1(n9788), .B2(n7512), .A(n7539), .ZN(n7513) );
  AOI21_X1 U9300 ( .B1(n10168), .B2(n7514), .A(n7513), .ZN(n7526) );
  AOI22_X1 U9301 ( .A1(n7747), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8756), .B2(
        n7742), .ZN(n7524) );
  NOR2_X1 U9302 ( .A1(n7515), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n7517) );
  NOR2_X1 U9303 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  OR2_X1 U9304 ( .A1(n7518), .A2(n8515), .ZN(n7519) );
  INV_X1 U9305 ( .A(n7519), .ZN(n7522) );
  INV_X1 U9306 ( .A(n7518), .ZN(n7521) );
  NOR2_X1 U9307 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n8512), .ZN(n8511) );
  NOR2_X1 U9308 ( .A1(n7522), .A2(n8511), .ZN(n7523) );
  NAND2_X1 U9309 ( .A1(n7524), .A2(n7523), .ZN(n7741) );
  OAI211_X1 U9310 ( .C1(n7524), .C2(n7523), .A(n10151), .B(n7741), .ZN(n7525)
         );
  OAI211_X1 U9311 ( .C1(n10152), .C2(n7742), .A(n7526), .B(n7525), .ZN(
        P2_U3261) );
  XNOR2_X1 U9312 ( .A(n8836), .B(n6201), .ZN(n7527) );
  NAND2_X1 U9313 ( .A1(n8720), .A2(n6204), .ZN(n7528) );
  NAND2_X1 U9314 ( .A1(n7527), .A2(n7528), .ZN(n7564) );
  INV_X1 U9315 ( .A(n7527), .ZN(n7530) );
  INV_X1 U9316 ( .A(n7528), .ZN(n7529) );
  NAND2_X1 U9317 ( .A1(n7530), .A2(n7529), .ZN(n7531) );
  NAND2_X1 U9318 ( .A1(n7564), .A2(n7531), .ZN(n7538) );
  INV_X1 U9319 ( .A(n7565), .ZN(n7536) );
  AOI21_X1 U9320 ( .B1(n7538), .B2(n7537), .A(n7536), .ZN(n7543) );
  AOI22_X1 U9321 ( .A1(n10137), .A2(n8743), .B1(n10136), .B2(n8742), .ZN(n7540) );
  OAI211_X1 U9322 ( .C1(n8240), .C2(n8755), .A(n7540), .B(n7539), .ZN(n7541)
         );
  AOI21_X1 U9323 ( .B1(n8836), .B2(n8228), .A(n7541), .ZN(n7542) );
  OAI21_X1 U9324 ( .B1(n7543), .B2(n8233), .A(n7542), .ZN(P2_U3228) );
  INV_X1 U9325 ( .A(n7544), .ZN(n7548) );
  OAI222_X1 U9326 ( .A1(n8888), .A2(n7546), .B1(n8883), .B2(n7548), .C1(n7545), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9327 ( .A1(P1_U3084), .A2(n7549), .B1(n4389), .B2(n7548), .C1(
        n7547), .C2(n9782), .ZN(P1_U3328) );
  OAI21_X1 U9328 ( .B1(n7551), .B2(n8417), .A(n7550), .ZN(n7552) );
  AOI222_X1 U9329 ( .A1(n10193), .A2(n7552), .B1(n8720), .B2(n10190), .C1(
        n8458), .C2(n10189), .ZN(n8847) );
  OAI21_X1 U9330 ( .B1(n7555), .B2(n7554), .A(n7553), .ZN(n8843) );
  OR2_X1 U9331 ( .A1(n7556), .A2(n8335), .ZN(n7557) );
  AND2_X1 U9332 ( .A1(n8752), .A2(n7557), .ZN(n8845) );
  NAND2_X1 U9333 ( .A1(n8845), .A2(n8711), .ZN(n7561) );
  INV_X1 U9334 ( .A(n7558), .ZN(n7559) );
  AOI22_X1 U9335 ( .A1(n10224), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n7559), .B2(
        n8698), .ZN(n7560) );
  OAI211_X1 U9336 ( .C1(n8335), .C2(n10200), .A(n7561), .B(n7560), .ZN(n7562)
         );
  AOI21_X1 U9337 ( .B1(n8843), .B2(n10202), .A(n7562), .ZN(n7563) );
  OAI21_X1 U9338 ( .B1(n8847), .B2(n10224), .A(n7563), .ZN(P2_U3281) );
  XNOR2_X1 U9339 ( .A(n8831), .B(n6201), .ZN(n7578) );
  NAND2_X1 U9340 ( .A1(n8742), .A2(n6204), .ZN(n7577) );
  XNOR2_X1 U9341 ( .A(n7578), .B(n7577), .ZN(n7579) );
  XNOR2_X1 U9342 ( .A(n7580), .B(n7579), .ZN(n7570) );
  OAI22_X1 U9343 ( .A1(n8240), .A2(n8731), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8525), .ZN(n7568) );
  OAI22_X1 U9344 ( .A1(n7566), .A2(n8224), .B1(n8225), .B2(n8683), .ZN(n7567)
         );
  AOI211_X1 U9345 ( .C1(n8831), .C2(n8228), .A(n7568), .B(n7567), .ZN(n7569)
         );
  OAI21_X1 U9346 ( .B1(n7570), .B2(n8233), .A(n7569), .ZN(P2_U3230) );
  INV_X1 U9347 ( .A(n7571), .ZN(n7575) );
  OAI222_X1 U9348 ( .A1(P1_U3084), .A2(n7573), .B1(n4389), .B2(n7575), .C1(
        n7572), .C2(n9782), .ZN(P1_U3327) );
  OAI222_X1 U9349 ( .A1(n8888), .A2(n7576), .B1(n8883), .B2(n7575), .C1(n7574), 
        .C2(P2_U3152), .ZN(P2_U3332) );
  XNOR2_X1 U9350 ( .A(n8826), .B(n8138), .ZN(n8112) );
  NAND2_X1 U9351 ( .A1(n8721), .A2(n6204), .ZN(n8110) );
  XNOR2_X1 U9352 ( .A(n8112), .B(n8110), .ZN(n8108) );
  XNOR2_X1 U9353 ( .A(n8109), .B(n8108), .ZN(n7585) );
  OAI22_X1 U9354 ( .A1(n8240), .A2(n8697), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8536), .ZN(n7583) );
  OAI22_X1 U9355 ( .A1(n7581), .A2(n8224), .B1(n8225), .B2(n8218), .ZN(n7582)
         );
  AOI211_X1 U9356 ( .C1(n8826), .C2(n8228), .A(n7583), .B(n7582), .ZN(n7584)
         );
  OAI21_X1 U9357 ( .B1(n7585), .B2(n8233), .A(n7584), .ZN(P2_U3240) );
  INV_X1 U9358 ( .A(n7586), .ZN(n7590) );
  AOI21_X1 U9359 ( .B1(n9774), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n7587), .ZN(
        n7588) );
  OAI21_X1 U9360 ( .B1(n7590), .B2(n4389), .A(n7588), .ZN(P1_U3326) );
  OAI222_X1 U9361 ( .A1(n8888), .A2(n7591), .B1(n8883), .B2(n7590), .C1(n7589), 
        .C2(P2_U3152), .ZN(P2_U3331) );
  INV_X1 U9362 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7791) );
  INV_X1 U9363 ( .A(n7592), .ZN(n7593) );
  NOR2_X1 U9364 ( .A1(n7593), .A2(SI_29_), .ZN(n7594) );
  MUX2_X1 U9365 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7800), .Z(n7796) );
  XNOR2_X1 U9366 ( .A(n7794), .B(SI_30_), .ZN(n7790) );
  INV_X1 U9367 ( .A(n7790), .ZN(n8882) );
  OAI222_X1 U9368 ( .A1(n9782), .A2(n7791), .B1(n4389), .B2(n8882), .C1(
        P1_U3084), .C2(n7596), .ZN(P1_U3323) );
  XNOR2_X1 U9369 ( .A(n7598), .B(n7597), .ZN(n8770) );
  INV_X1 U9370 ( .A(n8558), .ZN(n7601) );
  INV_X1 U9371 ( .A(n7599), .ZN(n7600) );
  AOI21_X1 U9372 ( .B1(n8771), .B2(n7601), .A(n7600), .ZN(n8772) );
  INV_X1 U9373 ( .A(n7602), .ZN(n8184) );
  AOI22_X1 U9374 ( .A1(n8184), .A2(n8698), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n10224), .ZN(n7603) );
  OAI21_X1 U9375 ( .B1(n8181), .B2(n10200), .A(n7603), .ZN(n7610) );
  XOR2_X1 U9376 ( .A(n8426), .B(n7604), .Z(n7608) );
  NAND2_X1 U9377 ( .A1(n8454), .A2(n10190), .ZN(n7606) );
  NAND2_X1 U9378 ( .A1(n8455), .A2(n10189), .ZN(n7605) );
  AOI211_X1 U9379 ( .C1(n8711), .C2(n8772), .A(n7610), .B(n7609), .ZN(n7611)
         );
  OAI21_X1 U9380 ( .B1(n8770), .B2(n8713), .A(n7611), .ZN(P2_U3268) );
  OAI222_X1 U9381 ( .A1(n8888), .A2(n7613), .B1(n8883), .B2(n7612), .C1(n8257), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  AND2_X1 U9382 ( .A1(n9143), .A2(n7634), .ZN(n7614) );
  AOI21_X1 U9383 ( .B1(n9408), .B2(n4388), .A(n7614), .ZN(n7711) );
  INV_X1 U9384 ( .A(n7711), .ZN(n7713) );
  NAND2_X1 U9385 ( .A1(n9408), .A2(n6674), .ZN(n7616) );
  NAND2_X1 U9386 ( .A1(n9143), .A2(n4388), .ZN(n7615) );
  NAND2_X1 U9387 ( .A1(n7616), .A2(n7615), .ZN(n7617) );
  AOI22_X1 U9388 ( .A1(n9419), .A2(n4386), .B1(n7634), .B2(n9204), .ZN(n7704)
         );
  NAND2_X1 U9389 ( .A1(n9419), .A2(n6674), .ZN(n7619) );
  NAND2_X1 U9390 ( .A1(n9204), .A2(n4388), .ZN(n7618) );
  NAND2_X1 U9391 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  XNOR2_X1 U9392 ( .A(n7620), .B(n7716), .ZN(n7702) );
  INV_X1 U9393 ( .A(n7702), .ZN(n7703) );
  NAND2_X1 U9394 ( .A1(n9351), .A2(n6674), .ZN(n7625) );
  NAND2_X1 U9395 ( .A1(n9327), .A2(n4388), .ZN(n7624) );
  NAND2_X1 U9396 ( .A1(n7625), .A2(n7624), .ZN(n7626) );
  XNOR2_X1 U9397 ( .A(n7626), .B(n7716), .ZN(n7631) );
  NAND2_X1 U9398 ( .A1(n7630), .A2(n7631), .ZN(n8890) );
  NAND2_X1 U9399 ( .A1(n9340), .A2(n6674), .ZN(n7628) );
  NAND2_X1 U9400 ( .A1(n9311), .A2(n4386), .ZN(n7627) );
  NAND2_X1 U9401 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  XNOR2_X1 U9402 ( .A(n7629), .B(n7770), .ZN(n7639) );
  INV_X1 U9403 ( .A(n7630), .ZN(n7633) );
  NAND2_X1 U9404 ( .A1(n9351), .A2(n4386), .ZN(n7636) );
  NAND2_X1 U9405 ( .A1(n7634), .A2(n9327), .ZN(n7635) );
  NAND2_X1 U9406 ( .A1(n7636), .A2(n7635), .ZN(n8893) );
  NAND2_X1 U9407 ( .A1(n9340), .A2(n4386), .ZN(n7638) );
  NAND2_X1 U9408 ( .A1(n7634), .A2(n9311), .ZN(n7637) );
  NAND2_X1 U9409 ( .A1(n7638), .A2(n7637), .ZN(n9015) );
  INV_X1 U9410 ( .A(n7639), .ZN(n7640) );
  NAND2_X1 U9411 ( .A1(n9318), .A2(n6674), .ZN(n7642) );
  NAND2_X1 U9412 ( .A1(n9328), .A2(n4388), .ZN(n7641) );
  NAND2_X1 U9413 ( .A1(n7642), .A2(n7641), .ZN(n7643) );
  XNOR2_X1 U9414 ( .A(n7643), .B(n7716), .ZN(n7646) );
  NAND2_X1 U9415 ( .A1(n9318), .A2(n4386), .ZN(n7645) );
  NAND2_X1 U9416 ( .A1(n7634), .A2(n9328), .ZN(n7644) );
  NAND2_X1 U9417 ( .A1(n7645), .A2(n7644), .ZN(n7647) );
  INV_X1 U9418 ( .A(n7646), .ZN(n7649) );
  INV_X1 U9419 ( .A(n7647), .ZN(n7648) );
  NAND2_X1 U9420 ( .A1(n7649), .A2(n7648), .ZN(n8940) );
  NAND2_X1 U9421 ( .A1(n8937), .A2(n8940), .ZN(n8949) );
  NAND2_X1 U9422 ( .A1(n9452), .A2(n6674), .ZN(n7651) );
  NAND2_X1 U9423 ( .A1(n9310), .A2(n4388), .ZN(n7650) );
  NAND2_X1 U9424 ( .A1(n7651), .A2(n7650), .ZN(n7652) );
  XNOR2_X1 U9425 ( .A(n7652), .B(n7716), .ZN(n7654) );
  AND2_X1 U9426 ( .A1(n7634), .A2(n9310), .ZN(n7653) );
  AOI21_X1 U9427 ( .B1(n9452), .B2(n4391), .A(n7653), .ZN(n7655) );
  XNOR2_X1 U9428 ( .A(n7654), .B(n7655), .ZN(n8950) );
  NAND2_X1 U9429 ( .A1(n8949), .A2(n8950), .ZN(n8948) );
  INV_X1 U9430 ( .A(n7654), .ZN(n7656) );
  NAND2_X1 U9431 ( .A1(n7656), .A2(n7655), .ZN(n7657) );
  NAND2_X1 U9432 ( .A1(n9447), .A2(n6674), .ZN(n7659) );
  NAND2_X1 U9433 ( .A1(n9298), .A2(n4386), .ZN(n7658) );
  NAND2_X1 U9434 ( .A1(n7659), .A2(n7658), .ZN(n7660) );
  XNOR2_X1 U9435 ( .A(n7660), .B(n7770), .ZN(n7663) );
  NAND2_X1 U9436 ( .A1(n9447), .A2(n4391), .ZN(n7662) );
  NAND2_X1 U9437 ( .A1(n7634), .A2(n9298), .ZN(n7661) );
  NAND2_X1 U9438 ( .A1(n7662), .A2(n7661), .ZN(n9004) );
  NAND2_X1 U9439 ( .A1(n9442), .A2(n6674), .ZN(n7666) );
  NAND2_X1 U9440 ( .A1(n9284), .A2(n4391), .ZN(n7665) );
  NAND2_X1 U9441 ( .A1(n7666), .A2(n7665), .ZN(n7667) );
  XNOR2_X1 U9442 ( .A(n7667), .B(n7716), .ZN(n8911) );
  NAND2_X1 U9443 ( .A1(n9442), .A2(n4386), .ZN(n7669) );
  NAND2_X1 U9444 ( .A1(n7634), .A2(n9284), .ZN(n7668) );
  NAND2_X1 U9445 ( .A1(n7669), .A2(n7668), .ZN(n8912) );
  NAND2_X1 U9446 ( .A1(n9439), .A2(n6674), .ZN(n7671) );
  NAND2_X1 U9447 ( .A1(n9263), .A2(n4388), .ZN(n7670) );
  NAND2_X1 U9448 ( .A1(n7671), .A2(n7670), .ZN(n7672) );
  XNOR2_X1 U9449 ( .A(n7672), .B(n7716), .ZN(n7675) );
  NAND2_X1 U9450 ( .A1(n9439), .A2(n4388), .ZN(n7674) );
  NAND2_X1 U9451 ( .A1(n7634), .A2(n9263), .ZN(n7673) );
  NAND2_X1 U9452 ( .A1(n7674), .A2(n7673), .ZN(n7676) );
  INV_X1 U9453 ( .A(n7675), .ZN(n7678) );
  INV_X1 U9454 ( .A(n7676), .ZN(n7677) );
  NAND2_X1 U9455 ( .A1(n7678), .A2(n7677), .ZN(n8971) );
  NAND2_X1 U9456 ( .A1(n9241), .A2(n6674), .ZN(n7681) );
  NAND2_X1 U9457 ( .A1(n9212), .A2(n4388), .ZN(n7680) );
  NAND2_X1 U9458 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  XNOR2_X1 U9459 ( .A(n7682), .B(n7716), .ZN(n7684) );
  AND2_X1 U9460 ( .A1(n7634), .A2(n9212), .ZN(n7683) );
  AOI21_X1 U9461 ( .B1(n9241), .B2(n4386), .A(n7683), .ZN(n7685) );
  XNOR2_X1 U9462 ( .A(n7684), .B(n7685), .ZN(n8921) );
  INV_X1 U9463 ( .A(n7684), .ZN(n7686) );
  AND2_X1 U9464 ( .A1(n9228), .A2(n7634), .ZN(n7687) );
  AOI21_X1 U9465 ( .B1(n9427), .B2(n4386), .A(n7687), .ZN(n7692) );
  NAND2_X1 U9466 ( .A1(n7691), .A2(n7692), .ZN(n8978) );
  NAND2_X1 U9467 ( .A1(n9427), .A2(n6674), .ZN(n7689) );
  NAND2_X1 U9468 ( .A1(n9228), .A2(n4388), .ZN(n7688) );
  NAND2_X1 U9469 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  XNOR2_X1 U9470 ( .A(n7690), .B(n7716), .ZN(n8981) );
  NAND2_X1 U9471 ( .A1(n8978), .A2(n8981), .ZN(n7695) );
  NAND2_X1 U9472 ( .A1(n9422), .A2(n6674), .ZN(n7697) );
  NAND2_X1 U9473 ( .A1(n9211), .A2(n4391), .ZN(n7696) );
  NAND2_X1 U9474 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  XNOR2_X1 U9475 ( .A(n7698), .B(n7770), .ZN(n7701) );
  NAND2_X1 U9476 ( .A1(n9422), .A2(n4386), .ZN(n7700) );
  NAND2_X1 U9477 ( .A1(n9211), .A2(n4385), .ZN(n7699) );
  NAND2_X1 U9478 ( .A1(n7700), .A2(n7699), .ZN(n8901) );
  XOR2_X1 U9479 ( .A(n7704), .B(n7702), .Z(n8960) );
  AOI21_X1 U9480 ( .B1(n7704), .B2(n7703), .A(n8959), .ZN(n8930) );
  AOI22_X1 U9481 ( .A1(n9412), .A2(n4386), .B1(n7634), .B2(n9029), .ZN(n7708)
         );
  NAND2_X1 U9482 ( .A1(n9412), .A2(n6674), .ZN(n7706) );
  NAND2_X1 U9483 ( .A1(n9029), .A2(n4391), .ZN(n7705) );
  NAND2_X1 U9484 ( .A1(n7706), .A2(n7705), .ZN(n7707) );
  XNOR2_X1 U9485 ( .A(n7707), .B(n7716), .ZN(n7710) );
  XOR2_X1 U9486 ( .A(n7708), .B(n7710), .Z(n8931) );
  INV_X1 U9487 ( .A(n7708), .ZN(n7709) );
  XOR2_X1 U9488 ( .A(n7711), .B(n7712), .Z(n7735) );
  NAND2_X1 U9489 ( .A1(n9401), .A2(n6674), .ZN(n7715) );
  NAND2_X1 U9490 ( .A1(n9028), .A2(n4386), .ZN(n7714) );
  NAND2_X1 U9491 ( .A1(n7715), .A2(n7714), .ZN(n7717) );
  XNOR2_X1 U9492 ( .A(n7717), .B(n7716), .ZN(n7723) );
  INV_X1 U9493 ( .A(n7723), .ZN(n7721) );
  NAND2_X1 U9494 ( .A1(n9401), .A2(n4391), .ZN(n7719) );
  NAND2_X1 U9495 ( .A1(n9028), .A2(n7634), .ZN(n7718) );
  NAND2_X1 U9496 ( .A1(n7719), .A2(n7718), .ZN(n7722) );
  INV_X1 U9497 ( .A(n7722), .ZN(n7720) );
  NAND2_X1 U9498 ( .A1(n7721), .A2(n7720), .ZN(n7782) );
  NAND2_X1 U9499 ( .A1(n7723), .A2(n7722), .ZN(n7775) );
  NAND2_X1 U9500 ( .A1(n7782), .A2(n7775), .ZN(n7724) );
  XNOR2_X1 U9501 ( .A(n7776), .B(n7724), .ZN(n7730) );
  AOI22_X1 U9502 ( .A1(n9019), .A2(n9143), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n7726) );
  INV_X1 U9503 ( .A(n9021), .ZN(n8962) );
  NAND2_X1 U9504 ( .A1(n8962), .A2(n9147), .ZN(n7725) );
  OAI211_X1 U9505 ( .C1(n7727), .C2(n9017), .A(n7726), .B(n7725), .ZN(n7728)
         );
  AOI21_X1 U9506 ( .B1(n9401), .B2(n9023), .A(n7728), .ZN(n7729) );
  OAI21_X1 U9507 ( .B1(n7730), .B2(n9025), .A(n7729), .ZN(P1_U3212) );
  OAI222_X1 U9508 ( .A1(n5658), .A2(P1_U3084), .B1(n4389), .B2(n7732), .C1(
        n7731), .C2(n9782), .ZN(P1_U3329) );
  INV_X1 U9509 ( .A(n7733), .ZN(n8107) );
  INV_X1 U9510 ( .A(n7736), .ZN(n7740) );
  NOR2_X1 U9511 ( .A1(n9021), .A2(n9156), .ZN(n7738) );
  OAI22_X1 U9512 ( .A1(n9164), .A2(n9017), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9733), .ZN(n7737) );
  AOI211_X1 U9513 ( .C1(n9019), .C2(n9029), .A(n7738), .B(n7737), .ZN(n7739)
         );
  OAI211_X1 U9514 ( .C1(n9159), .C2(n8958), .A(n7740), .B(n7739), .ZN(P1_U3238) );
  AOI22_X1 U9515 ( .A1(n7748), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n8732), .B2(
        n8533), .ZN(n8523) );
  OAI21_X1 U9516 ( .B1(n8756), .B2(n7742), .A(n7741), .ZN(n8524) );
  NAND2_X1 U9517 ( .A1(n8523), .A2(n8524), .ZN(n8522) );
  NAND2_X1 U9518 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8535), .ZN(n8534) );
  NAND2_X1 U9519 ( .A1(n7743), .A2(n8538), .ZN(n7744) );
  XNOR2_X1 U9520 ( .A(n8538), .B(n7745), .ZN(n8541) );
  XNOR2_X1 U9521 ( .A(n7748), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n8527) );
  OAI21_X1 U9522 ( .B1(n7747), .B2(P2_REG1_REG_16__SCAN_IN), .A(n7746), .ZN(
        n8528) );
  NOR2_X1 U9523 ( .A1(n8527), .A2(n8528), .ZN(n8526) );
  AOI21_X1 U9524 ( .B1(n7748), .B2(P2_REG1_REG_17__SCAN_IN), .A(n8526), .ZN(
        n8540) );
  NAND2_X1 U9525 ( .A1(n8541), .A2(n8540), .ZN(n8539) );
  OR2_X1 U9526 ( .A1(n8538), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n7749) );
  NAND2_X1 U9527 ( .A1(n8539), .A2(n7749), .ZN(n7751) );
  XNOR2_X1 U9528 ( .A(n7751), .B(n7750), .ZN(n7755) );
  INV_X1 U9529 ( .A(n7755), .ZN(n7752) );
  AOI22_X1 U9530 ( .A1(n7753), .A2(n10151), .B1(n7752), .B2(n10168), .ZN(n7757) );
  NOR2_X1 U9531 ( .A1(n7753), .A2(n10172), .ZN(n7754) );
  AOI211_X1 U9532 ( .C1(n10168), .C2(n7755), .A(n10166), .B(n7754), .ZN(n7756)
         );
  MUX2_X1 U9533 ( .A(n7757), .B(n7756), .S(n8680), .Z(n7758) );
  NAND2_X1 U9534 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8168) );
  OAI211_X1 U9535 ( .C1(n4510), .C2(n9788), .A(n7758), .B(n8168), .ZN(P2_U3264) );
  INV_X1 U9536 ( .A(n7759), .ZN(n7763) );
  INV_X1 U9537 ( .A(n7760), .ZN(n7761) );
  AOI22_X1 U9538 ( .A1(n7761), .A2(n8698), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n10224), .ZN(n7762) );
  OAI21_X1 U9539 ( .B1(n7763), .B2(n10200), .A(n7762), .ZN(n7765) );
  NAND2_X1 U9540 ( .A1(n9396), .A2(n6674), .ZN(n7769) );
  NAND2_X1 U9541 ( .A1(n9137), .A2(n4388), .ZN(n7768) );
  NAND2_X1 U9542 ( .A1(n7769), .A2(n7768), .ZN(n7771) );
  XNOR2_X1 U9543 ( .A(n7771), .B(n7770), .ZN(n7773) );
  AOI22_X1 U9544 ( .A1(n9396), .A2(n4388), .B1(n7634), .B2(n9137), .ZN(n7772)
         );
  XNOR2_X1 U9545 ( .A(n7773), .B(n7772), .ZN(n7783) );
  INV_X1 U9546 ( .A(n7783), .ZN(n7774) );
  NAND2_X1 U9547 ( .A1(n7774), .A2(n8951), .ZN(n7789) );
  AND2_X1 U9548 ( .A1(n7783), .A2(n7777), .ZN(n7778) );
  NAND2_X1 U9549 ( .A1(n7788), .A2(n7778), .ZN(n7787) );
  INV_X1 U9550 ( .A(n9130), .ZN(n7781) );
  AOI22_X1 U9551 ( .A1(n9007), .A2(n9027), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7780) );
  NAND2_X1 U9552 ( .A1(n9028), .A2(n9019), .ZN(n7779) );
  OAI211_X1 U9553 ( .C1(n9021), .C2(n7781), .A(n7780), .B(n7779), .ZN(n7785)
         );
  NOR3_X1 U9554 ( .A1(n7783), .A2(n9025), .A3(n7782), .ZN(n7784) );
  AOI211_X1 U9555 ( .C1(n9023), .C2(n9396), .A(n7785), .B(n7784), .ZN(n7786)
         );
  OAI211_X1 U9556 ( .C1(n7789), .C2(n7788), .A(n7787), .B(n7786), .ZN(P1_U3218) );
  NAND2_X1 U9557 ( .A1(n7790), .A2(n7804), .ZN(n7793) );
  OR2_X1 U9558 ( .A1(n7806), .A2(n7791), .ZN(n7792) );
  INV_X1 U9559 ( .A(n7794), .ZN(n7795) );
  NAND2_X1 U9560 ( .A1(n7795), .A2(SI_30_), .ZN(n7799) );
  NAND2_X1 U9561 ( .A1(n7797), .A2(n7796), .ZN(n7798) );
  MUX2_X1 U9562 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7800), .Z(n7801) );
  XNOR2_X1 U9563 ( .A(n7801), .B(SI_31_), .ZN(n7802) );
  NAND2_X1 U9564 ( .A1(n8876), .A2(n7804), .ZN(n7808) );
  INV_X1 U9565 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7805) );
  OR2_X1 U9566 ( .A1(n7806), .A2(n7805), .ZN(n7807) );
  NAND2_X1 U9567 ( .A1(n8024), .A2(n9392), .ZN(n7809) );
  MUX2_X1 U9568 ( .A(n8011), .B(n7810), .S(n7933), .Z(n7812) );
  MUX2_X1 U9569 ( .A(n8019), .B(n8014), .S(n7933), .Z(n7811) );
  OAI21_X1 U9570 ( .B1(n7812), .B2(n9128), .A(n7811), .ZN(n7918) );
  OR2_X1 U9571 ( .A1(n9419), .A2(n9175), .ZN(n7898) );
  NAND2_X1 U9572 ( .A1(n7904), .A2(n7899), .ZN(n8010) );
  AND2_X1 U9573 ( .A1(n7898), .A2(n8006), .ZN(n7813) );
  NOR2_X1 U9574 ( .A1(n8010), .A2(n7813), .ZN(n7814) );
  INV_X1 U9575 ( .A(n7933), .ZN(n7920) );
  MUX2_X1 U9576 ( .A(n7898), .B(n7814), .S(n7920), .Z(n7903) );
  NAND2_X1 U9577 ( .A1(n7899), .A2(n7815), .ZN(n7816) );
  NAND2_X1 U9578 ( .A1(n7939), .A2(n7816), .ZN(n7817) );
  MUX2_X1 U9579 ( .A(n7819), .B(n7818), .S(n7933), .Z(n7821) );
  NAND2_X1 U9580 ( .A1(n7821), .A2(n7820), .ZN(n7829) );
  INV_X1 U9581 ( .A(n7822), .ZN(n8075) );
  OAI211_X1 U9582 ( .C1(n7829), .C2(n8075), .A(n8074), .B(n7995), .ZN(n7823)
         );
  NAND3_X1 U9583 ( .A1(n7823), .A2(n8036), .A3(n7828), .ZN(n7826) );
  AND2_X1 U9584 ( .A1(n7967), .A2(n7996), .ZN(n7825) );
  AOI21_X1 U9585 ( .B1(n7826), .B2(n7825), .A(n7824), .ZN(n7834) );
  AND2_X1 U9586 ( .A1(n7828), .A2(n7827), .ZN(n7964) );
  NAND2_X1 U9587 ( .A1(n7829), .A2(n7964), .ZN(n7831) );
  NOR2_X1 U9588 ( .A1(n9963), .A2(n5032), .ZN(n7830) );
  NAND2_X1 U9589 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  AOI21_X1 U9590 ( .B1(n7832), .B2(n7972), .A(n5014), .ZN(n7833) );
  MUX2_X1 U9591 ( .A(n7968), .B(n7973), .S(n7933), .Z(n7835) );
  NAND2_X1 U9592 ( .A1(n7838), .A2(n7837), .ZN(n7848) );
  AND2_X1 U9593 ( .A1(n7976), .A2(n7839), .ZN(n7966) );
  AND2_X1 U9594 ( .A1(n7978), .A2(n7966), .ZN(n7840) );
  NAND2_X1 U9595 ( .A1(n7850), .A2(n7847), .ZN(n7979) );
  AOI21_X1 U9596 ( .B1(n7848), .B2(n7840), .A(n7979), .ZN(n7845) );
  INV_X1 U9597 ( .A(n7976), .ZN(n7842) );
  MUX2_X1 U9598 ( .A(n7842), .B(n7841), .S(n7920), .Z(n7843) );
  NAND3_X1 U9599 ( .A1(n7850), .A2(n9365), .A3(n7843), .ZN(n7844) );
  OAI21_X1 U9600 ( .B1(n7845), .B2(n7933), .A(n7844), .ZN(n7846) );
  NAND2_X1 U9601 ( .A1(n9351), .A2(n9368), .ZN(n7983) );
  NAND2_X1 U9602 ( .A1(n7846), .A2(n7983), .ZN(n7855) );
  NAND3_X1 U9603 ( .A1(n7848), .A2(n7974), .A3(n7847), .ZN(n7849) );
  AND2_X1 U9604 ( .A1(n7983), .A2(n7978), .ZN(n7994) );
  NAND2_X1 U9605 ( .A1(n7849), .A2(n7994), .ZN(n7853) );
  AND2_X1 U9606 ( .A1(n7850), .A2(n7933), .ZN(n7852) );
  AOI21_X1 U9607 ( .B1(n7853), .B2(n7852), .A(n7851), .ZN(n7854) );
  NAND2_X1 U9608 ( .A1(n7855), .A2(n7854), .ZN(n7858) );
  AND2_X1 U9609 ( .A1(n7986), .A2(n7993), .ZN(n7856) );
  AND2_X1 U9610 ( .A1(n7859), .A2(n9307), .ZN(n7989) );
  MUX2_X1 U9611 ( .A(n7856), .B(n7989), .S(n7933), .Z(n7857) );
  NAND2_X1 U9612 ( .A1(n7858), .A2(n7857), .ZN(n7861) );
  MUX2_X1 U9613 ( .A(n7859), .B(n7986), .S(n7933), .Z(n7860) );
  NAND2_X1 U9614 ( .A1(n7861), .A2(n7860), .ZN(n7875) );
  NAND4_X1 U9615 ( .A1(n7877), .A2(n7954), .A3(n7959), .A4(n7933), .ZN(n7883)
         );
  AOI21_X1 U9616 ( .B1(n7875), .B2(n5711), .A(n9452), .ZN(n7882) );
  NAND2_X1 U9617 ( .A1(n9298), .A2(n7920), .ZN(n7864) );
  OAI22_X1 U9618 ( .A1(n9447), .A2(n7864), .B1(n9248), .B2(n7933), .ZN(n7863)
         );
  INV_X1 U9619 ( .A(n7863), .ZN(n7866) );
  OR3_X1 U9620 ( .A1(n9447), .A2(n9248), .A3(n7864), .ZN(n7865) );
  OAI21_X1 U9621 ( .B1(n7866), .B2(n9442), .A(n7865), .ZN(n7867) );
  NAND2_X1 U9622 ( .A1(n7951), .A2(n7867), .ZN(n7873) );
  NOR2_X1 U9623 ( .A1(n9298), .A2(n7920), .ZN(n7868) );
  NAND2_X1 U9624 ( .A1(n9447), .A2(n7868), .ZN(n7869) );
  OAI21_X1 U9625 ( .B1(n7920), .B2(n9284), .A(n7869), .ZN(n7871) );
  INV_X1 U9626 ( .A(n7869), .ZN(n7870) );
  AOI22_X1 U9627 ( .A1(n7871), .A2(n9442), .B1(n7870), .B2(n9248), .ZN(n7872)
         );
  OAI211_X1 U9628 ( .C1(n7951), .C2(n7920), .A(n7873), .B(n7872), .ZN(n7874)
         );
  INV_X1 U9629 ( .A(n7874), .ZN(n7881) );
  NAND2_X1 U9630 ( .A1(n7875), .A2(n4723), .ZN(n7876) );
  NAND2_X1 U9631 ( .A1(n7876), .A2(n5711), .ZN(n7879) );
  NAND2_X1 U9632 ( .A1(n8003), .A2(n7987), .ZN(n7955) );
  NOR2_X1 U9633 ( .A1(n7955), .A2(n7933), .ZN(n7878) );
  NAND4_X1 U9634 ( .A1(n7879), .A2(n7878), .A3(n7877), .A4(n7951), .ZN(n7880)
         );
  OAI211_X1 U9635 ( .C1(n7883), .C2(n7882), .A(n7881), .B(n7880), .ZN(n7887)
         );
  OR2_X1 U9636 ( .A1(n7885), .A2(n7884), .ZN(n7888) );
  INV_X1 U9637 ( .A(n7888), .ZN(n7886) );
  AND2_X1 U9638 ( .A1(n7887), .A2(n7886), .ZN(n7896) );
  NAND2_X1 U9639 ( .A1(n7888), .A2(n9209), .ZN(n7889) );
  NAND2_X1 U9640 ( .A1(n7889), .A2(n8028), .ZN(n7890) );
  MUX2_X1 U9641 ( .A(n7890), .B(n7953), .S(n7933), .Z(n7895) );
  INV_X1 U9642 ( .A(n8027), .ZN(n7892) );
  MUX2_X1 U9643 ( .A(n7892), .B(n7891), .S(n7933), .Z(n7893) );
  INV_X1 U9644 ( .A(n7893), .ZN(n7894) );
  OAI21_X1 U9645 ( .B1(n7896), .B2(n7895), .A(n7894), .ZN(n7901) );
  AND2_X1 U9646 ( .A1(n7898), .A2(n7897), .ZN(n7942) );
  NAND4_X1 U9647 ( .A1(n7901), .A2(n7942), .A3(n7900), .A4(n7899), .ZN(n7902)
         );
  MUX2_X1 U9648 ( .A(n9408), .B(n9143), .S(n7933), .Z(n7913) );
  MUX2_X1 U9649 ( .A(n7939), .B(n7904), .S(n7933), .Z(n7905) );
  NAND3_X1 U9650 ( .A1(n7914), .A2(n7913), .A3(n7905), .ZN(n7912) );
  AOI21_X1 U9651 ( .B1(n9176), .B2(n7906), .A(n9408), .ZN(n7909) );
  INV_X1 U9652 ( .A(n7939), .ZN(n7907) );
  AOI21_X1 U9653 ( .B1(n9159), .B2(n7907), .A(n9143), .ZN(n7908) );
  MUX2_X1 U9654 ( .A(n7909), .B(n7908), .S(n7920), .Z(n7910) );
  INV_X1 U9655 ( .A(n7910), .ZN(n7911) );
  NAND2_X1 U9656 ( .A1(n7912), .A2(n7911), .ZN(n7916) );
  OR2_X1 U9657 ( .A1(n7914), .A2(n7913), .ZN(n7915) );
  INV_X1 U9658 ( .A(n8024), .ZN(n7925) );
  NAND3_X1 U9659 ( .A1(n7919), .A2(n4718), .A3(n9123), .ZN(n7923) );
  NAND2_X1 U9660 ( .A1(n9027), .A2(n7933), .ZN(n7922) );
  NAND2_X1 U9661 ( .A1(n9392), .A2(n7920), .ZN(n7921) );
  NAND3_X1 U9662 ( .A1(n7923), .A2(n7922), .A3(n7921), .ZN(n7924) );
  INV_X1 U9663 ( .A(n9111), .ZN(n7927) );
  NAND2_X1 U9664 ( .A1(n7938), .A2(n7927), .ZN(n8089) );
  NAND2_X1 U9665 ( .A1(n8089), .A2(n7933), .ZN(n7931) );
  NAND2_X1 U9666 ( .A1(n9111), .A2(n4859), .ZN(n7929) );
  NAND2_X1 U9667 ( .A1(n9821), .A2(n7929), .ZN(n8021) );
  INV_X1 U9668 ( .A(n8021), .ZN(n7930) );
  OAI21_X1 U9669 ( .B1(n8024), .B2(n7933), .A(n7932), .ZN(n7937) );
  NAND2_X1 U9670 ( .A1(n7934), .A2(n4392), .ZN(n7935) );
  AND2_X1 U9671 ( .A1(n7940), .A2(n7939), .ZN(n7941) );
  NAND2_X1 U9672 ( .A1(n8012), .A2(n7941), .ZN(n8016) );
  INV_X1 U9673 ( .A(n7942), .ZN(n7943) );
  NOR2_X1 U9674 ( .A1(n8016), .A2(n7943), .ZN(n8078) );
  INV_X1 U9675 ( .A(n7944), .ZN(n7948) );
  INV_X1 U9676 ( .A(n7945), .ZN(n7946) );
  OAI21_X1 U9677 ( .B1(n7946), .B2(n8063), .A(n8067), .ZN(n7947) );
  AOI21_X1 U9678 ( .B1(n7948), .B2(n8070), .A(n7947), .ZN(n7949) );
  NOR2_X1 U9679 ( .A1(n7949), .A2(n8075), .ZN(n7991) );
  NAND2_X1 U9680 ( .A1(n8074), .A2(n7950), .ZN(n8068) );
  AND2_X1 U9681 ( .A1(n7962), .A2(n5017), .ZN(n7952) );
  OR2_X1 U9682 ( .A1(n7953), .A2(n7952), .ZN(n8002) );
  INV_X1 U9683 ( .A(n7954), .ZN(n7958) );
  INV_X1 U9684 ( .A(n7955), .ZN(n7956) );
  OAI21_X1 U9685 ( .B1(n7958), .B2(n7957), .A(n7956), .ZN(n7961) );
  AND4_X1 U9686 ( .A1(n7962), .A2(n7961), .A3(n7960), .A4(n7959), .ZN(n7963)
         );
  OAI21_X1 U9687 ( .B1(n8002), .B2(n7963), .A(n8028), .ZN(n7992) );
  INV_X1 U9688 ( .A(n7964), .ZN(n7965) );
  NOR2_X1 U9689 ( .A1(n7992), .A2(n7965), .ZN(n8077) );
  INV_X1 U9690 ( .A(n7966), .ZN(n7971) );
  NAND2_X1 U9691 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  AND2_X1 U9692 ( .A1(n7969), .A2(n7973), .ZN(n7970) );
  NOR2_X1 U9693 ( .A1(n7971), .A2(n7970), .ZN(n7997) );
  NAND2_X1 U9694 ( .A1(n7973), .A2(n7972), .ZN(n7977) );
  INV_X1 U9695 ( .A(n7974), .ZN(n7975) );
  AOI22_X1 U9696 ( .A1(n7997), .A2(n7977), .B1(n7976), .B2(n7975), .ZN(n7982)
         );
  INV_X1 U9697 ( .A(n7978), .ZN(n7981) );
  INV_X1 U9698 ( .A(n7979), .ZN(n7980) );
  OAI21_X1 U9699 ( .B1(n7982), .B2(n7981), .A(n7980), .ZN(n7984) );
  NAND3_X1 U9700 ( .A1(n7984), .A2(n7993), .A3(n7983), .ZN(n7988) );
  NAND3_X1 U9701 ( .A1(n7987), .A2(n7986), .A3(n7985), .ZN(n8001) );
  AOI21_X1 U9702 ( .B1(n7989), .B2(n7988), .A(n8001), .ZN(n8072) );
  INV_X1 U9703 ( .A(n8072), .ZN(n7990) );
  OAI211_X1 U9704 ( .C1(n7991), .C2(n8068), .A(n8077), .B(n7990), .ZN(n8009)
         );
  INV_X1 U9705 ( .A(n7992), .ZN(n8008) );
  INV_X1 U9706 ( .A(n7993), .ZN(n8000) );
  INV_X1 U9707 ( .A(n7994), .ZN(n7999) );
  NAND3_X1 U9708 ( .A1(n7997), .A2(n7996), .A3(n7995), .ZN(n7998) );
  NOR4_X1 U9709 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n8005)
         );
  INV_X1 U9710 ( .A(n8002), .ZN(n8004) );
  OAI211_X1 U9711 ( .C1(n8072), .C2(n8005), .A(n8004), .B(n8003), .ZN(n8007)
         );
  AOI21_X1 U9712 ( .B1(n8008), .B2(n8007), .A(n8006), .ZN(n8081) );
  NAND2_X1 U9713 ( .A1(n8009), .A2(n8081), .ZN(n8018) );
  INV_X1 U9714 ( .A(n8010), .ZN(n8017) );
  AOI21_X1 U9715 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8015) );
  OAI211_X1 U9716 ( .C1(n8017), .C2(n8016), .A(n8015), .B(n8014), .ZN(n8084)
         );
  AOI21_X1 U9717 ( .B1(n8078), .B2(n8018), .A(n8084), .ZN(n8022) );
  NAND2_X1 U9718 ( .A1(n8020), .A2(n8019), .ZN(n8082) );
  OAI211_X1 U9719 ( .C1(n8022), .C2(n8082), .A(n8021), .B(n8088), .ZN(n8023)
         );
  AOI211_X1 U9720 ( .C1(n8024), .C2(n8023), .A(n8054), .B(n8052), .ZN(n8025)
         );
  NOR2_X1 U9721 ( .A1(n8025), .A2(n9192), .ZN(n8057) );
  INV_X1 U9722 ( .A(n8026), .ZN(n8086) );
  NAND2_X1 U9723 ( .A1(n8028), .A2(n8027), .ZN(n9214) );
  NAND4_X1 U9724 ( .A1(n8030), .A2(n10014), .A3(n8029), .A4(n8061), .ZN(n8033)
         );
  NOR4_X1 U9725 ( .A1(n8033), .A2(n8032), .A3(n8031), .A4(n9984), .ZN(n8037)
         );
  NAND4_X1 U9726 ( .A1(n8037), .A2(n8036), .A3(n8035), .A4(n8034), .ZN(n8038)
         );
  NOR4_X1 U9727 ( .A1(n9369), .A2(n8040), .A3(n8039), .A4(n8038), .ZN(n8041)
         );
  NAND4_X1 U9728 ( .A1(n9331), .A2(n9365), .A3(n8041), .A4(n9343), .ZN(n8042)
         );
  NOR4_X1 U9729 ( .A1(n8043), .A2(n9289), .A3(n9306), .A4(n8042), .ZN(n8044)
         );
  NAND4_X1 U9730 ( .A1(n4777), .A2(n9245), .A3(n9261), .A4(n8044), .ZN(n8045)
         );
  NOR4_X1 U9731 ( .A1(n9162), .A2(n9203), .A3(n9214), .A4(n8045), .ZN(n8047)
         );
  NAND4_X1 U9732 ( .A1(n9136), .A2(n8048), .A3(n8047), .A4(n8046), .ZN(n8049)
         );
  NOR4_X1 U9733 ( .A1(n8086), .A2(n9128), .A3(n8050), .A4(n8049), .ZN(n8051)
         );
  NAND2_X1 U9734 ( .A1(n8051), .A2(n8089), .ZN(n8055) );
  INV_X1 U9735 ( .A(n8052), .ZN(n8053) );
  OAI21_X1 U9736 ( .B1(n9117), .B2(n4859), .A(n8053), .ZN(n8090) );
  OAI21_X1 U9737 ( .B1(n8055), .B2(n8090), .A(n8054), .ZN(n8056) );
  MUX2_X1 U9738 ( .A(n9192), .B(n8057), .S(n8056), .Z(n8058) );
  AOI21_X1 U9739 ( .B1(n4392), .B2(n8061), .A(n8060), .ZN(n8066) );
  OAI211_X1 U9740 ( .C1(n8066), .C2(n8065), .A(n8064), .B(n8063), .ZN(n8071)
         );
  INV_X1 U9741 ( .A(n8067), .ZN(n8069) );
  AOI211_X1 U9742 ( .C1(n8071), .C2(n8070), .A(n8069), .B(n8068), .ZN(n8073)
         );
  AOI211_X1 U9743 ( .C1(n8075), .C2(n8074), .A(n8073), .B(n8072), .ZN(n8076)
         );
  NAND2_X1 U9744 ( .A1(n8077), .A2(n8076), .ZN(n8080) );
  INV_X1 U9745 ( .A(n8078), .ZN(n8079) );
  AOI21_X1 U9746 ( .B1(n8081), .B2(n8080), .A(n8079), .ZN(n8085) );
  INV_X1 U9747 ( .A(n8082), .ZN(n8083) );
  OAI21_X1 U9748 ( .B1(n8085), .B2(n8084), .A(n8083), .ZN(n8087) );
  AOI21_X1 U9749 ( .B1(n8088), .B2(n8087), .A(n8086), .ZN(n8091) );
  OAI21_X1 U9750 ( .B1(n8091), .B2(n8090), .A(n8089), .ZN(n8095) );
  NOR2_X1 U9751 ( .A1(n8095), .A2(n8092), .ZN(n8094) );
  INV_X1 U9752 ( .A(n8095), .ZN(n8098) );
  OAI21_X1 U9753 ( .B1(n8098), .B2(n8097), .A(n8096), .ZN(n8104) );
  NOR4_X1 U9754 ( .A1(n8099), .A2(n10072), .A3(n9874), .A4(n9869), .ZN(n8103)
         );
  OAI21_X1 U9755 ( .B1(n8101), .B2(n8100), .A(P1_B_REG_SCAN_IN), .ZN(n8102) );
  OAI22_X1 U9756 ( .A1(n8105), .A2(n8104), .B1(n8103), .B2(n8102), .ZN(
        P1_U3240) );
  OAI222_X1 U9757 ( .A1(n4389), .A2(n8107), .B1(n5120), .B2(P1_U3084), .C1(
        n8106), .C2(n9782), .ZN(P1_U3324) );
  INV_X1 U9758 ( .A(n8110), .ZN(n8111) );
  XNOR2_X1 U9759 ( .A(n8823), .B(n6201), .ZN(n8113) );
  NAND2_X1 U9760 ( .A1(n8707), .A2(n6204), .ZN(n8114) );
  NAND2_X1 U9761 ( .A1(n8113), .A2(n8114), .ZN(n8120) );
  INV_X1 U9762 ( .A(n8113), .ZN(n8116) );
  INV_X1 U9763 ( .A(n8114), .ZN(n8115) );
  NAND2_X1 U9764 ( .A1(n8116), .A2(n8115), .ZN(n8117) );
  NAND2_X1 U9765 ( .A1(n8120), .A2(n8117), .ZN(n8166) );
  XNOR2_X1 U9766 ( .A(n8814), .B(n6201), .ZN(n8121) );
  NAND2_X1 U9767 ( .A1(n8658), .A2(n6204), .ZN(n8122) );
  XNOR2_X1 U9768 ( .A(n8121), .B(n8122), .ZN(n8215) );
  INV_X1 U9769 ( .A(n8121), .ZN(n8124) );
  INV_X1 U9770 ( .A(n8122), .ZN(n8123) );
  XNOR2_X1 U9771 ( .A(n8809), .B(n8138), .ZN(n8127) );
  NAND2_X1 U9772 ( .A1(n8673), .A2(n6204), .ZN(n8125) );
  XNOR2_X1 U9773 ( .A(n8127), .B(n8125), .ZN(n8187) );
  INV_X1 U9774 ( .A(n8125), .ZN(n8126) );
  XOR2_X1 U9775 ( .A(n8138), .B(n8804), .Z(n8130) );
  XNOR2_X1 U9776 ( .A(n8129), .B(n8130), .ZN(n8230) );
  XNOR2_X1 U9777 ( .A(n8798), .B(n8138), .ZN(n8134) );
  NAND2_X1 U9778 ( .A1(n8457), .A2(n6204), .ZN(n8155) );
  XNOR2_X1 U9779 ( .A(n8792), .B(n8138), .ZN(n8136) );
  AND2_X1 U9780 ( .A1(n8618), .A2(n6204), .ZN(n8206) );
  XOR2_X1 U9781 ( .A(n8138), .B(n8789), .Z(n8196) );
  NAND2_X1 U9782 ( .A1(n8456), .A2(n6204), .ZN(n8195) );
  AND2_X1 U9783 ( .A1(n8565), .A2(n6204), .ZN(n8137) );
  NAND2_X1 U9784 ( .A1(n8144), .A2(n8137), .ZN(n8147) );
  OAI21_X1 U9785 ( .B1(n8144), .B2(n8137), .A(n8147), .ZN(n8236) );
  XNOR2_X1 U9786 ( .A(n8777), .B(n8138), .ZN(n8139) );
  AND2_X1 U9787 ( .A1(n8455), .A2(n6204), .ZN(n8140) );
  NAND2_X1 U9788 ( .A1(n8139), .A2(n8140), .ZN(n8174) );
  INV_X1 U9789 ( .A(n8139), .ZN(n8142) );
  INV_X1 U9790 ( .A(n8140), .ZN(n8141) );
  NAND2_X1 U9791 ( .A1(n8142), .A2(n8141), .ZN(n8143) );
  NOR2_X1 U9792 ( .A1(n8234), .A2(n8148), .ZN(n8146) );
  NAND3_X1 U9793 ( .A1(n8144), .A2(n8229), .A3(n8565), .ZN(n8145) );
  OAI21_X1 U9794 ( .B1(n8146), .B2(n8233), .A(n8145), .ZN(n8149) );
  NAND2_X1 U9795 ( .A1(n8149), .A2(n8175), .ZN(n8154) );
  AOI22_X1 U9796 ( .A1(n8559), .A2(n8210), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8150) );
  OAI21_X1 U9797 ( .B1(n8151), .B2(n8224), .A(n8150), .ZN(n8152) );
  AOI21_X1 U9798 ( .B1(n10136), .B2(n8564), .A(n8152), .ZN(n8153) );
  OAI211_X1 U9799 ( .C1(n8561), .C2(n10143), .A(n8154), .B(n8153), .ZN(
        P2_U3216) );
  NAND2_X1 U9800 ( .A1(n8155), .A2(n10141), .ZN(n8158) );
  NAND2_X1 U9801 ( .A1(n8457), .A2(n8229), .ZN(n8157) );
  MUX2_X1 U9802 ( .A(n8158), .B(n8157), .S(n8156), .Z(n8163) );
  OAI22_X1 U9803 ( .A1(n8240), .A2(n8620), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9715), .ZN(n8161) );
  OAI22_X1 U9804 ( .A1(n8159), .A2(n8225), .B1(n8224), .B2(n8190), .ZN(n8160)
         );
  AOI211_X1 U9805 ( .C1(n8798), .C2(n8228), .A(n8161), .B(n8160), .ZN(n8162)
         );
  NAND2_X1 U9806 ( .A1(n8163), .A2(n8162), .ZN(P2_U3218) );
  INV_X1 U9807 ( .A(n8164), .ZN(n8165) );
  AOI21_X1 U9808 ( .B1(n8167), .B2(n8166), .A(n8165), .ZN(n8173) );
  INV_X1 U9809 ( .A(n8687), .ZN(n8170) );
  AOI22_X1 U9810 ( .A1(n10137), .A2(n8721), .B1(n10136), .B2(n8658), .ZN(n8169) );
  OAI211_X1 U9811 ( .C1(n8240), .C2(n8170), .A(n8169), .B(n8168), .ZN(n8171)
         );
  AOI21_X1 U9812 ( .B1(n8823), .B2(n8228), .A(n8171), .ZN(n8172) );
  OAI21_X1 U9813 ( .B1(n8173), .B2(n8233), .A(n8172), .ZN(P2_U3221) );
  NAND2_X1 U9814 ( .A1(n8564), .A2(n6204), .ZN(n8176) );
  XNOR2_X1 U9815 ( .A(n8176), .B(n8138), .ZN(n8179) );
  NOR3_X1 U9816 ( .A1(n8181), .A2(n8228), .A3(n8179), .ZN(n8177) );
  AOI21_X1 U9817 ( .B1(n8181), .B2(n8179), .A(n8177), .ZN(n8183) );
  NAND3_X1 U9818 ( .A1(n8771), .A2(n10143), .A3(n8179), .ZN(n8178) );
  OAI21_X1 U9819 ( .B1(n8771), .B2(n8179), .A(n8178), .ZN(n8180) );
  OAI21_X1 U9820 ( .B1(n8181), .B2(n10143), .A(n8233), .ZN(n8182) );
  AOI22_X1 U9821 ( .A1(n8184), .A2(n8210), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n8186) );
  AOI22_X1 U9822 ( .A1(n8454), .A2(n10136), .B1(n8455), .B2(n10137), .ZN(n8185) );
  XNOR2_X1 U9823 ( .A(n8188), .B(n8187), .ZN(n8194) );
  OAI22_X1 U9824 ( .A1(n8240), .A2(n8651), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8189), .ZN(n8192) );
  OAI22_X1 U9825 ( .A1(n8684), .A2(n8224), .B1(n8225), .B2(n8190), .ZN(n8191)
         );
  AOI211_X1 U9826 ( .C1(n8809), .C2(n8228), .A(n8192), .B(n8191), .ZN(n8193)
         );
  OAI21_X1 U9827 ( .B1(n8194), .B2(n8233), .A(n8193), .ZN(P2_U3225) );
  XNOR2_X1 U9828 ( .A(n8196), .B(n8195), .ZN(n8197) );
  XNOR2_X1 U9829 ( .A(n8198), .B(n8197), .ZN(n8205) );
  AND2_X1 U9830 ( .A1(n8618), .A2(n10189), .ZN(n8199) );
  AOI21_X1 U9831 ( .B1(n8565), .B2(n10190), .A(n8199), .ZN(n8589) );
  INV_X1 U9832 ( .A(n8585), .ZN(n8200) );
  AOI22_X1 U9833 ( .A1(n8200), .A2(n8210), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8201) );
  OAI21_X1 U9834 ( .B1(n8589), .B2(n8202), .A(n8201), .ZN(n8203) );
  AOI21_X1 U9835 ( .B1(n8789), .B2(n8228), .A(n8203), .ZN(n8204) );
  OAI21_X1 U9836 ( .B1(n8205), .B2(n8233), .A(n8204), .ZN(P2_U3227) );
  NAND2_X1 U9837 ( .A1(n8618), .A2(n8229), .ZN(n8209) );
  OR2_X1 U9838 ( .A1(n8206), .A2(n8233), .ZN(n8208) );
  MUX2_X1 U9839 ( .A(n8209), .B(n8208), .S(n8207), .Z(n8214) );
  AOI22_X1 U9840 ( .A1(n8603), .A2(n8210), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8213) );
  AOI22_X1 U9841 ( .A1(n8456), .A2(n10136), .B1(n10137), .B2(n8457), .ZN(n8212) );
  NAND2_X1 U9842 ( .A1(n8792), .A2(n8228), .ZN(n8211) );
  NAND4_X1 U9843 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(
        P2_U3231) );
  XNOR2_X1 U9844 ( .A(n8216), .B(n8215), .ZN(n8222) );
  OAI22_X1 U9845 ( .A1(n8240), .A2(n8666), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8217), .ZN(n8220) );
  OAI22_X1 U9846 ( .A1(n8218), .A2(n8224), .B1(n8225), .B2(n8641), .ZN(n8219)
         );
  AOI211_X1 U9847 ( .C1(n8814), .C2(n8228), .A(n8220), .B(n8219), .ZN(n8221)
         );
  OAI21_X1 U9848 ( .B1(n8222), .B2(n8233), .A(n8221), .ZN(P2_U3235) );
  OAI22_X1 U9849 ( .A1(n8240), .A2(n8633), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8223), .ZN(n8227) );
  OAI22_X1 U9850 ( .A1(n8642), .A2(n8225), .B1(n8224), .B2(n8641), .ZN(n8226)
         );
  AOI211_X1 U9851 ( .C1(n8804), .C2(n8228), .A(n8227), .B(n8226), .ZN(n8232)
         );
  NAND3_X1 U9852 ( .A1(n8230), .A2(n8229), .A3(n8659), .ZN(n8231) );
  OAI211_X1 U9853 ( .C1(n4580), .C2(n8233), .A(n8232), .B(n8231), .ZN(P2_U3237) );
  NAND2_X1 U9854 ( .A1(n8455), .A2(n10190), .ZN(n8238) );
  NAND2_X1 U9855 ( .A1(n8456), .A2(n10189), .ZN(n8237) );
  NAND2_X1 U9856 ( .A1(n8238), .A2(n8237), .ZN(n8574) );
  OAI22_X1 U9857 ( .A1(n8579), .A2(n8240), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8239), .ZN(n8241) );
  AOI21_X1 U9858 ( .B1(n8574), .B2(n8242), .A(n8241), .ZN(n8243) );
  OR2_X1 U9859 ( .A1(n8547), .A2(n8436), .ZN(n8246) );
  INV_X1 U9860 ( .A(n8246), .ZN(n8248) );
  INV_X1 U9861 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9722) );
  NOR2_X1 U9862 ( .A1(n8250), .A2(n9722), .ZN(n8244) );
  INV_X1 U9863 ( .A(n8769), .ZN(n8553) );
  OAI211_X1 U9864 ( .C1(n8769), .C2(n8246), .A(n8245), .B(n8386), .ZN(n8247)
         );
  OAI21_X1 U9865 ( .B1(n8248), .B2(n8391), .A(n8247), .ZN(n8254) );
  NAND2_X1 U9866 ( .A1(n8876), .A2(n8249), .ZN(n8252) );
  OR2_X1 U9867 ( .A1(n8250), .A2(n9647), .ZN(n8251) );
  INV_X1 U9868 ( .A(n8547), .ZN(n8253) );
  NAND2_X1 U9869 ( .A1(n8553), .A2(n6146), .ZN(n8390) );
  INV_X1 U9870 ( .A(n8395), .ZN(n8256) );
  AND2_X1 U9871 ( .A1(n8256), .A2(n8391), .ZN(n8400) );
  NAND3_X1 U9872 ( .A1(n8257), .A2(n8271), .A3(n8680), .ZN(n8393) );
  MUX2_X1 U9873 ( .A(n8399), .B(n8400), .S(n8393), .Z(n8398) );
  NAND2_X1 U9874 ( .A1(n8789), .A2(n8608), .ZN(n8258) );
  OAI211_X1 U9875 ( .C1(n8259), .C2(n8369), .A(n8573), .B(n8258), .ZN(n8260)
         );
  NAND2_X1 U9876 ( .A1(n8260), .A2(n8393), .ZN(n8371) );
  INV_X1 U9877 ( .A(n8625), .ZN(n8424) );
  NAND2_X1 U9878 ( .A1(n8353), .A2(n8261), .ZN(n8264) );
  INV_X1 U9879 ( .A(n8262), .ZN(n8263) );
  INV_X1 U9880 ( .A(n8393), .ZN(n8380) );
  MUX2_X1 U9881 ( .A(n8264), .B(n8263), .S(n8380), .Z(n8265) );
  INV_X1 U9882 ( .A(n8265), .ZN(n8345) );
  NAND2_X1 U9883 ( .A1(n8268), .A2(n8267), .ZN(n8403) );
  AND2_X1 U9884 ( .A1(n8267), .A2(n8266), .ZN(n8269) );
  NAND2_X1 U9885 ( .A1(n8270), .A2(n8393), .ZN(n8287) );
  INV_X1 U9886 ( .A(n8289), .ZN(n8285) );
  AND2_X1 U9887 ( .A1(n8275), .A2(n8271), .ZN(n8273) );
  OAI211_X1 U9888 ( .C1(n8273), .C2(n8272), .A(n8280), .B(n8276), .ZN(n8274)
         );
  NAND2_X1 U9889 ( .A1(n8274), .A2(n8278), .ZN(n8283) );
  NAND2_X1 U9890 ( .A1(n8276), .A2(n8275), .ZN(n8279) );
  NAND3_X1 U9891 ( .A1(n8279), .A2(n8278), .A3(n8277), .ZN(n8281) );
  NAND2_X1 U9892 ( .A1(n8281), .A2(n8280), .ZN(n8282) );
  MUX2_X1 U9893 ( .A(n8283), .B(n8282), .S(n8380), .Z(n8284) );
  NAND3_X1 U9894 ( .A1(n8285), .A2(n8284), .A3(n10187), .ZN(n8286) );
  NAND2_X1 U9895 ( .A1(n8289), .A2(n8288), .ZN(n8293) );
  OAI21_X1 U9896 ( .B1(n8291), .B2(n8290), .A(n8405), .ZN(n8292) );
  NAND2_X1 U9897 ( .A1(n8293), .A2(n8292), .ZN(n8295) );
  NAND2_X1 U9898 ( .A1(n8295), .A2(n8294), .ZN(n8296) );
  NAND2_X1 U9899 ( .A1(n8308), .A2(n8299), .ZN(n8301) );
  AND2_X1 U9900 ( .A1(n8304), .A2(n8314), .ZN(n8302) );
  MUX2_X1 U9901 ( .A(n8310), .B(n8302), .S(n8393), .Z(n8303) );
  AND2_X1 U9902 ( .A1(n8303), .A2(n8312), .ZN(n8316) );
  NAND2_X1 U9903 ( .A1(n8321), .A2(n8304), .ZN(n8305) );
  NAND3_X1 U9904 ( .A1(n8308), .A2(n8307), .A3(n8306), .ZN(n8311) );
  NAND2_X1 U9905 ( .A1(n8317), .A2(n8312), .ZN(n8313) );
  INV_X1 U9906 ( .A(n8314), .ZN(n8315) );
  AND2_X1 U9907 ( .A1(n8318), .A2(n8317), .ZN(n8320) );
  INV_X1 U9908 ( .A(n8322), .ZN(n8319) );
  AOI21_X1 U9909 ( .B1(n8325), .B2(n8320), .A(n8319), .ZN(n8327) );
  AND2_X1 U9910 ( .A1(n8322), .A2(n8321), .ZN(n8324) );
  AOI21_X1 U9911 ( .B1(n8325), .B2(n8324), .A(n8323), .ZN(n8326) );
  INV_X1 U9912 ( .A(n8328), .ZN(n8416) );
  MUX2_X1 U9913 ( .A(n8330), .B(n8329), .S(n8393), .Z(n8331) );
  MUX2_X1 U9914 ( .A(n8333), .B(n8332), .S(n8393), .Z(n8334) );
  MUX2_X1 U9915 ( .A(n8336), .B(n8335), .S(n8393), .Z(n8338) );
  NAND2_X1 U9916 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  INV_X1 U9917 ( .A(n8717), .ZN(n8342) );
  MUX2_X1 U9918 ( .A(n8716), .B(n8340), .S(n8393), .Z(n8341) );
  NAND3_X1 U9919 ( .A1(n8343), .A2(n8342), .A3(n8341), .ZN(n8344) );
  NAND2_X1 U9920 ( .A1(n8345), .A2(n8344), .ZN(n8354) );
  INV_X1 U9921 ( .A(n8357), .ZN(n8348) );
  INV_X1 U9922 ( .A(n8349), .ZN(n8350) );
  MUX2_X1 U9923 ( .A(n8351), .B(n8350), .S(n8380), .Z(n8352) );
  OAI22_X1 U9924 ( .A1(n8424), .A2(n8352), .B1(n8380), .B2(n8606), .ZN(n8363)
         );
  AOI21_X1 U9925 ( .B1(n8354), .B2(n8353), .A(n4482), .ZN(n8359) );
  NAND2_X1 U9926 ( .A1(n8356), .A2(n8355), .ZN(n8358) );
  OAI211_X1 U9927 ( .C1(n8359), .C2(n8358), .A(n8357), .B(n8638), .ZN(n8361)
         );
  NAND4_X1 U9928 ( .A1(n8615), .A2(n8361), .A3(n8380), .A4(n8360), .ZN(n8362)
         );
  NAND3_X1 U9929 ( .A1(n8363), .A2(n8365), .A3(n8362), .ZN(n8368) );
  NAND2_X1 U9930 ( .A1(n8365), .A2(n8364), .ZN(n8366) );
  NAND2_X1 U9931 ( .A1(n8366), .A2(n8380), .ZN(n8367) );
  NAND2_X1 U9932 ( .A1(n8368), .A2(n8367), .ZN(n8370) );
  INV_X1 U9933 ( .A(n8372), .ZN(n8373) );
  AOI21_X1 U9934 ( .B1(n8375), .B2(n8373), .A(n8393), .ZN(n8374) );
  OAI21_X1 U9935 ( .B1(n8562), .B2(n8393), .A(n4461), .ZN(n8379) );
  MUX2_X1 U9936 ( .A(n8377), .B(n8376), .S(n8393), .Z(n8378) );
  MUX2_X1 U9937 ( .A(n8382), .B(n8381), .S(n8380), .Z(n8383) );
  NAND3_X1 U9938 ( .A1(n8385), .A2(n8384), .A3(n8383), .ZN(n8389) );
  MUX2_X1 U9939 ( .A(n8387), .B(n8386), .S(n8393), .Z(n8388) );
  NAND4_X1 U9940 ( .A1(n8391), .A2(n8390), .A3(n8389), .A4(n8388), .ZN(n8397)
         );
  INV_X1 U9941 ( .A(n8392), .ZN(n8394) );
  MUX2_X1 U9942 ( .A(n8395), .B(n8394), .S(n8393), .Z(n8396) );
  AOI21_X1 U9943 ( .B1(n8398), .B2(n8397), .A(n8396), .ZN(n8434) );
  INV_X1 U9944 ( .A(n8434), .ZN(n8440) );
  OAI21_X1 U9945 ( .B1(n8432), .B2(n8433), .A(n10298), .ZN(n8439) );
  INV_X1 U9946 ( .A(n8399), .ZN(n8430) );
  INV_X1 U9947 ( .A(n8400), .ZN(n8429) );
  INV_X1 U9948 ( .A(n8671), .ZN(n8422) );
  NOR4_X1 U9949 ( .A1(n8402), .A2(n8401), .A3(n10245), .A4(n6128), .ZN(n8406)
         );
  INV_X1 U9950 ( .A(n8403), .ZN(n8404) );
  NAND4_X1 U9951 ( .A1(n8406), .A2(n8405), .A3(n8404), .A4(n10187), .ZN(n8409)
         );
  NOR4_X1 U9952 ( .A1(n8409), .A2(n8408), .A3(n4749), .A4(n8407), .ZN(n8412)
         );
  NAND3_X1 U9953 ( .A1(n8412), .A2(n8411), .A3(n8410), .ZN(n8413) );
  NOR4_X1 U9954 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), .ZN(n8418)
         );
  NAND4_X1 U9955 ( .A1(n8744), .A2(n8419), .A3(n8418), .A4(n8417), .ZN(n8420)
         );
  NOR4_X1 U9956 ( .A1(n8681), .A2(n8703), .A3(n8717), .A4(n8420), .ZN(n8421)
         );
  NAND4_X1 U9957 ( .A1(n8637), .A2(n8422), .A3(n8656), .A4(n8421), .ZN(n8423)
         );
  NOR4_X1 U9958 ( .A1(n4770), .A2(n8424), .A3(n8596), .A4(n8423), .ZN(n8425)
         );
  NAND4_X1 U9959 ( .A1(n8426), .A2(n4461), .A3(n8425), .A4(n8587), .ZN(n8427)
         );
  NOR4_X1 U9960 ( .A1(n8430), .A2(n8429), .A3(n8428), .A4(n8427), .ZN(n8431)
         );
  XNOR2_X1 U9961 ( .A(n8431), .B(n8730), .ZN(n8437) );
  AOI21_X1 U9962 ( .B1(n8434), .B2(n8433), .A(n8432), .ZN(n8435) );
  AOI21_X1 U9963 ( .B1(n8437), .B2(n8436), .A(n8435), .ZN(n8438) );
  AOI21_X1 U9964 ( .B1(n8440), .B2(n8439), .A(n8438), .ZN(n8441) );
  INV_X1 U9965 ( .A(n8451), .ZN(n8448) );
  NAND3_X1 U9966 ( .A1(n8730), .A2(n8443), .A3(n8442), .ZN(n8444) );
  NOR3_X1 U9967 ( .A1(n8446), .A2(n8445), .A3(n8444), .ZN(n8447) );
  MUX2_X1 U9968 ( .A(n8448), .B(n8447), .S(n4811), .Z(n8450) );
  INV_X1 U9969 ( .A(P2_B_REG_SCAN_IN), .ZN(n8449) );
  OAI22_X1 U9970 ( .A1(n8452), .A2(n8451), .B1(n8450), .B2(n8449), .ZN(
        P2_U3244) );
  MUX2_X1 U9971 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8453), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9972 ( .A(n8454), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8469), .Z(
        P2_U3581) );
  MUX2_X1 U9973 ( .A(n8564), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8469), .Z(
        P2_U3580) );
  MUX2_X1 U9974 ( .A(n8455), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8469), .Z(
        P2_U3579) );
  MUX2_X1 U9975 ( .A(n8565), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8469), .Z(
        P2_U3578) );
  MUX2_X1 U9976 ( .A(n8456), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8469), .Z(
        P2_U3577) );
  MUX2_X1 U9977 ( .A(n8618), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8469), .Z(
        P2_U3576) );
  MUX2_X1 U9978 ( .A(n8457), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8469), .Z(
        P2_U3575) );
  MUX2_X1 U9979 ( .A(n8659), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8469), .Z(
        P2_U3574) );
  MUX2_X1 U9980 ( .A(n8673), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8469), .Z(
        P2_U3573) );
  MUX2_X1 U9981 ( .A(n8658), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8469), .Z(
        P2_U3572) );
  MUX2_X1 U9982 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8707), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U9983 ( .A(n8721), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8469), .Z(
        P2_U3570) );
  MUX2_X1 U9984 ( .A(n8742), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8469), .Z(
        P2_U3569) );
  MUX2_X1 U9985 ( .A(n8720), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8469), .Z(
        P2_U3568) );
  MUX2_X1 U9986 ( .A(n8743), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8469), .Z(
        P2_U3567) );
  MUX2_X1 U9987 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8458), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U9988 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8459), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U9989 ( .A(n8460), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8469), .Z(
        P2_U3564) );
  MUX2_X1 U9990 ( .A(n8461), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8469), .Z(
        P2_U3563) );
  MUX2_X1 U9991 ( .A(n8462), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8469), .Z(
        P2_U3562) );
  MUX2_X1 U9992 ( .A(n8463), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8469), .Z(
        P2_U3561) );
  MUX2_X1 U9993 ( .A(n8464), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8469), .Z(
        P2_U3560) );
  MUX2_X1 U9994 ( .A(n8465), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8469), .Z(
        P2_U3559) );
  MUX2_X1 U9995 ( .A(n8466), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8469), .Z(
        P2_U3558) );
  MUX2_X1 U9996 ( .A(n8467), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8469), .Z(
        P2_U3557) );
  MUX2_X1 U9997 ( .A(n10191), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8469), .Z(
        P2_U3556) );
  MUX2_X1 U9998 ( .A(n8468), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8469), .Z(
        P2_U3555) );
  MUX2_X1 U9999 ( .A(n5806), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8469), .Z(
        P2_U3554) );
  MUX2_X1 U10000 ( .A(n5787), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8469), .Z(
        P2_U3553) );
  OAI211_X1 U10001 ( .C1(n8472), .C2(n8471), .A(n10151), .B(n8470), .ZN(n8483)
         );
  INV_X1 U10002 ( .A(n8473), .ZN(n8474) );
  AOI21_X1 U10003 ( .B1(n10162), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n8474), .ZN(
        n8482) );
  NAND2_X1 U10004 ( .A1(n10166), .A2(n8475), .ZN(n8481) );
  AOI21_X1 U10005 ( .B1(n8478), .B2(n8477), .A(n8476), .ZN(n8479) );
  NAND2_X1 U10006 ( .A1(n10168), .A2(n8479), .ZN(n8480) );
  NAND4_X1 U10007 ( .A1(n8483), .A2(n8482), .A3(n8481), .A4(n8480), .ZN(
        P2_U3254) );
  OAI211_X1 U10008 ( .C1(n8486), .C2(n8485), .A(n10151), .B(n8484), .ZN(n8496)
         );
  NOR2_X1 U10009 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8487), .ZN(n8488) );
  AOI21_X1 U10010 ( .B1(n10162), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n8488), .ZN(
        n8495) );
  NAND2_X1 U10011 ( .A1(n10166), .A2(n8489), .ZN(n8494) );
  OAI211_X1 U10012 ( .C1(n8492), .C2(n8491), .A(n10168), .B(n8490), .ZN(n8493)
         );
  NAND4_X1 U10013 ( .A1(n8496), .A2(n8495), .A3(n8494), .A4(n8493), .ZN(
        P2_U3255) );
  OAI211_X1 U10014 ( .C1(n8499), .C2(n8498), .A(n10151), .B(n8497), .ZN(n8510)
         );
  NOR2_X1 U10015 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8500), .ZN(n8501) );
  AOI21_X1 U10016 ( .B1(n10162), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8501), .ZN(
        n8509) );
  NAND2_X1 U10017 ( .A1(n10166), .A2(n8502), .ZN(n8508) );
  OAI21_X1 U10018 ( .B1(n8505), .B2(n8504), .A(n8503), .ZN(n8506) );
  NAND2_X1 U10019 ( .A1(n10168), .A2(n8506), .ZN(n8507) );
  NAND4_X1 U10020 ( .A1(n8510), .A2(n8509), .A3(n8508), .A4(n8507), .ZN(
        P2_U3257) );
  AOI21_X1 U10021 ( .B1(n8512), .B2(P2_REG2_REG_15__SCAN_IN), .A(n8511), .ZN(
        n8513) );
  OR2_X1 U10022 ( .A1(n8513), .A2(n10172), .ZN(n8521) );
  NOR2_X1 U10023 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5973), .ZN(n8514) );
  AOI21_X1 U10024 ( .B1(n10162), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8514), .ZN(
        n8520) );
  NAND2_X1 U10025 ( .A1(n10166), .A2(n8515), .ZN(n8519) );
  OAI211_X1 U10026 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n8517), .A(n10168), .B(
        n8516), .ZN(n8518) );
  NAND4_X1 U10027 ( .A1(n8521), .A2(n8520), .A3(n8519), .A4(n8518), .ZN(
        P2_U3260) );
  OAI211_X1 U10028 ( .C1(n8524), .C2(n8523), .A(n10151), .B(n8522), .ZN(n8532)
         );
  NOR2_X1 U10029 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8525), .ZN(n8530) );
  AOI211_X1 U10030 ( .C1(n8528), .C2(n8527), .A(n8526), .B(n10153), .ZN(n8529)
         );
  AOI211_X1 U10031 ( .C1(n10162), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n8530), .B(
        n8529), .ZN(n8531) );
  OAI211_X1 U10032 ( .C1(n10152), .C2(n8533), .A(n8532), .B(n8531), .ZN(
        P2_U3262) );
  OAI211_X1 U10033 ( .C1(P2_REG2_REG_18__SCAN_IN), .C2(n8535), .A(n10151), .B(
        n8534), .ZN(n8546) );
  NOR2_X1 U10034 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8536), .ZN(n8537) );
  AOI21_X1 U10035 ( .B1(n10162), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8537), .ZN(
        n8545) );
  NAND2_X1 U10036 ( .A1(n10166), .A2(n8538), .ZN(n8544) );
  OAI21_X1 U10037 ( .B1(n8541), .B2(n8540), .A(n8539), .ZN(n8542) );
  NAND2_X1 U10038 ( .A1(n10168), .A2(n8542), .ZN(n8543) );
  NAND4_X1 U10039 ( .A1(n8546), .A2(n8545), .A3(n8544), .A4(n8543), .ZN(
        P2_U3263) );
  NAND2_X1 U10040 ( .A1(n8769), .A2(n8551), .ZN(n8765) );
  XNOR2_X1 U10041 ( .A(n8765), .B(n8762), .ZN(n8764) );
  NAND2_X1 U10042 ( .A1(n8548), .A2(n8547), .ZN(n8767) );
  NOR2_X1 U10043 ( .A1(n10224), .A2(n8767), .ZN(n8554) );
  AOI21_X1 U10044 ( .B1(n10224), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8554), .ZN(
        n8550) );
  NAND2_X1 U10045 ( .A1(n8762), .A2(n10183), .ZN(n8549) );
  OAI211_X1 U10046 ( .C1(n8764), .C2(n10219), .A(n8550), .B(n8549), .ZN(
        P2_U3265) );
  INV_X1 U10047 ( .A(n8551), .ZN(n8552) );
  NAND2_X1 U10048 ( .A1(n8553), .A2(n8552), .ZN(n8766) );
  NAND3_X1 U10049 ( .A1(n8766), .A2(n8711), .A3(n8765), .ZN(n8556) );
  AOI21_X1 U10050 ( .B1(n10224), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8554), .ZN(
        n8555) );
  OAI211_X1 U10051 ( .C1(n8769), .C2(n10200), .A(n8556), .B(n8555), .ZN(
        P2_U3266) );
  XNOR2_X1 U10052 ( .A(n8557), .B(n4461), .ZN(n8781) );
  AOI21_X1 U10053 ( .B1(n8777), .B2(n8576), .A(n8558), .ZN(n8778) );
  AOI22_X1 U10054 ( .A1(n8559), .A2(n8698), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n10224), .ZN(n8560) );
  OAI21_X1 U10055 ( .B1(n8561), .B2(n10200), .A(n8560), .ZN(n8568) );
  NAND2_X1 U10056 ( .A1(n8571), .A2(n8562), .ZN(n8563) );
  XNOR2_X1 U10057 ( .A(n8563), .B(n4461), .ZN(n8566) );
  AOI222_X1 U10058 ( .A1(n10193), .A2(n8566), .B1(n8565), .B2(n10189), .C1(
        n8564), .C2(n10190), .ZN(n8780) );
  NOR2_X1 U10059 ( .A1(n8780), .A2(n10224), .ZN(n8567) );
  AOI211_X1 U10060 ( .C1(n8778), .C2(n8711), .A(n8568), .B(n8567), .ZN(n8569)
         );
  OAI21_X1 U10061 ( .B1(n8781), .B2(n8713), .A(n8569), .ZN(P2_U3269) );
  XNOR2_X1 U10062 ( .A(n8570), .B(n4770), .ZN(n8786) );
  AOI22_X1 U10063 ( .A1(n8783), .A2(n10183), .B1(n10224), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8582) );
  OAI21_X1 U10064 ( .B1(n8573), .B2(n8572), .A(n8571), .ZN(n8575) );
  AOI21_X1 U10065 ( .B1(n8575), .B2(n10193), .A(n8574), .ZN(n8785) );
  INV_X1 U10066 ( .A(n8576), .ZN(n8577) );
  AOI211_X1 U10067 ( .C1(n8783), .C2(n8586), .A(n10298), .B(n8577), .ZN(n8782)
         );
  NAND2_X1 U10068 ( .A1(n8782), .A2(n8730), .ZN(n8578) );
  OAI211_X1 U10069 ( .C1(n10218), .C2(n8579), .A(n8785), .B(n8578), .ZN(n8580)
         );
  NAND2_X1 U10070 ( .A1(n8580), .A2(n10222), .ZN(n8581) );
  OAI211_X1 U10071 ( .C1(n8786), .C2(n8713), .A(n8582), .B(n8581), .ZN(
        P2_U3270) );
  XNOR2_X1 U10072 ( .A(n8583), .B(n8587), .ZN(n8791) );
  INV_X1 U10073 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n8584) );
  OAI22_X1 U10074 ( .A1(n8585), .A2(n10218), .B1(n8584), .B2(n10222), .ZN(
        n8593) );
  AOI211_X1 U10075 ( .C1(n8789), .C2(n8600), .A(n10298), .B(n4735), .ZN(n8788)
         );
  XNOR2_X1 U10076 ( .A(n8588), .B(n8587), .ZN(n8590) );
  OAI21_X1 U10077 ( .B1(n8590), .B2(n6148), .A(n8589), .ZN(n8787) );
  AOI21_X1 U10078 ( .B1(n8788), .B2(n8730), .A(n8787), .ZN(n8591) );
  NOR2_X1 U10079 ( .A1(n8591), .A2(n10224), .ZN(n8592) );
  AOI211_X1 U10080 ( .C1(n10183), .C2(n8789), .A(n8593), .B(n8592), .ZN(n8594)
         );
  OAI21_X1 U10081 ( .B1(n8713), .B2(n8791), .A(n8594), .ZN(P2_U3271) );
  OAI21_X1 U10082 ( .B1(n8597), .B2(n8596), .A(n8595), .ZN(n8598) );
  INV_X1 U10083 ( .A(n8598), .ZN(n8796) );
  INV_X1 U10084 ( .A(n8599), .ZN(n8602) );
  INV_X1 U10085 ( .A(n8600), .ZN(n8601) );
  AOI21_X1 U10086 ( .B1(n8792), .B2(n8602), .A(n8601), .ZN(n8793) );
  AOI22_X1 U10087 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(n10224), .B1(n8603), 
        .B2(n8698), .ZN(n8604) );
  OAI21_X1 U10088 ( .B1(n6059), .B2(n10200), .A(n8604), .ZN(n8613) );
  AOI21_X1 U10089 ( .B1(n8616), .B2(n8606), .A(n8605), .ZN(n8607) );
  NOR2_X1 U10090 ( .A1(n8607), .A2(n6148), .ZN(n8611) );
  OAI22_X1 U10091 ( .A1(n8608), .A2(n10211), .B1(n8642), .B2(n10210), .ZN(
        n8609) );
  AOI21_X1 U10092 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8795) );
  NOR2_X1 U10093 ( .A1(n8795), .A2(n10224), .ZN(n8612) );
  AOI211_X1 U10094 ( .C1(n8793), .C2(n8711), .A(n8613), .B(n8612), .ZN(n8614)
         );
  OAI21_X1 U10095 ( .B1(n8796), .B2(n8713), .A(n8614), .ZN(P2_U3272) );
  AND2_X1 U10096 ( .A1(n8636), .A2(n8615), .ZN(n8617) );
  OAI21_X1 U10097 ( .B1(n8617), .B2(n8625), .A(n8616), .ZN(n8619) );
  AOI222_X1 U10098 ( .A1(n10193), .A2(n8619), .B1(n8659), .B2(n10189), .C1(
        n8618), .C2(n10190), .ZN(n8801) );
  XOR2_X1 U10099 ( .A(n8631), .B(n8798), .Z(n8799) );
  INV_X1 U10100 ( .A(n8798), .ZN(n8623) );
  INV_X1 U10101 ( .A(n8620), .ZN(n8621) );
  AOI22_X1 U10102 ( .A1(n10224), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8621), 
        .B2(n8698), .ZN(n8622) );
  OAI21_X1 U10103 ( .B1(n8623), .B2(n10200), .A(n8622), .ZN(n8624) );
  AOI21_X1 U10104 ( .B1(n8799), .B2(n8711), .A(n8624), .ZN(n8629) );
  INV_X1 U10105 ( .A(n8803), .ZN(n8627) );
  NAND2_X1 U10106 ( .A1(n8626), .A2(n8625), .ZN(n8797) );
  NAND3_X1 U10107 ( .A1(n8627), .A2(n10202), .A3(n8797), .ZN(n8628) );
  OAI211_X1 U10108 ( .C1(n8801), .C2(n10224), .A(n8629), .B(n8628), .ZN(
        P2_U3273) );
  XOR2_X1 U10109 ( .A(n8637), .B(n8630), .Z(n8808) );
  INV_X1 U10110 ( .A(n8631), .ZN(n8632) );
  AOI21_X1 U10111 ( .B1(n8804), .B2(n8649), .A(n8632), .ZN(n8805) );
  INV_X1 U10112 ( .A(n8633), .ZN(n8634) );
  AOI22_X1 U10113 ( .A1(n10224), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8634), 
        .B2(n8698), .ZN(n8635) );
  OAI21_X1 U10114 ( .B1(n4739), .B2(n10200), .A(n8635), .ZN(n8646) );
  INV_X1 U10115 ( .A(n8636), .ZN(n8640) );
  AOI21_X1 U10116 ( .B1(n8655), .B2(n8638), .A(n8637), .ZN(n8639) );
  NOR3_X1 U10117 ( .A1(n8640), .A2(n8639), .A3(n6148), .ZN(n8644) );
  OAI22_X1 U10118 ( .A1(n8642), .A2(n10211), .B1(n8641), .B2(n10210), .ZN(
        n8643) );
  NOR2_X1 U10119 ( .A1(n8644), .A2(n8643), .ZN(n8807) );
  NOR2_X1 U10120 ( .A1(n8807), .A2(n10224), .ZN(n8645) );
  AOI211_X1 U10121 ( .C1(n8805), .C2(n8711), .A(n8646), .B(n8645), .ZN(n8647)
         );
  OAI21_X1 U10122 ( .B1(n8808), .B2(n8713), .A(n8647), .ZN(P2_U3274) );
  XNOR2_X1 U10123 ( .A(n8648), .B(n8656), .ZN(n8813) );
  INV_X1 U10124 ( .A(n8649), .ZN(n8650) );
  AOI21_X1 U10125 ( .B1(n8809), .B2(n4743), .A(n8650), .ZN(n8810) );
  INV_X1 U10126 ( .A(n8651), .ZN(n8652) );
  AOI22_X1 U10127 ( .A1(n10224), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8652), 
        .B2(n8698), .ZN(n8653) );
  OAI21_X1 U10128 ( .B1(n8654), .B2(n10200), .A(n8653), .ZN(n8662) );
  OAI21_X1 U10129 ( .B1(n8657), .B2(n8656), .A(n8655), .ZN(n8660) );
  AOI222_X1 U10130 ( .A1(n10193), .A2(n8660), .B1(n8659), .B2(n10190), .C1(
        n8658), .C2(n10189), .ZN(n8812) );
  NOR2_X1 U10131 ( .A1(n8812), .A2(n10224), .ZN(n8661) );
  AOI211_X1 U10132 ( .C1(n8810), .C2(n8711), .A(n8662), .B(n8661), .ZN(n8663)
         );
  OAI21_X1 U10133 ( .B1(n8713), .B2(n8813), .A(n8663), .ZN(P2_U3275) );
  XNOR2_X1 U10134 ( .A(n8664), .B(n8671), .ZN(n8818) );
  AOI21_X1 U10135 ( .B1(n8814), .B2(n8679), .A(n8665), .ZN(n8815) );
  INV_X1 U10136 ( .A(n8814), .ZN(n8669) );
  INV_X1 U10137 ( .A(n8666), .ZN(n8667) );
  AOI22_X1 U10138 ( .A1(n10224), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8667), 
        .B2(n8698), .ZN(n8668) );
  OAI21_X1 U10139 ( .B1(n8669), .B2(n10200), .A(n8668), .ZN(n8676) );
  NOR2_X1 U10140 ( .A1(n4426), .A2(n8670), .ZN(n8672) );
  XNOR2_X1 U10141 ( .A(n8672), .B(n8671), .ZN(n8674) );
  AOI222_X1 U10142 ( .A1(n10193), .A2(n8674), .B1(n8673), .B2(n10190), .C1(
        n8707), .C2(n10189), .ZN(n8817) );
  NOR2_X1 U10143 ( .A1(n8817), .A2(n10224), .ZN(n8675) );
  AOI211_X1 U10144 ( .C1(n8815), .C2(n8711), .A(n8676), .B(n8675), .ZN(n8677)
         );
  OAI21_X1 U10145 ( .B1(n8713), .B2(n8818), .A(n8677), .ZN(P2_U3276) );
  XOR2_X1 U10146 ( .A(n8678), .B(n8681), .Z(n8819) );
  OAI211_X1 U10147 ( .C1(n8689), .C2(n8695), .A(n8852), .B(n8679), .ZN(n8820)
         );
  NOR2_X1 U10148 ( .A1(n8820), .A2(n8680), .ZN(n8685) );
  AOI21_X1 U10149 ( .B1(n4602), .B2(n8681), .A(n4426), .ZN(n8682) );
  OAI222_X1 U10150 ( .A1(n10211), .A2(n8684), .B1(n10210), .B2(n8683), .C1(
        n6148), .C2(n8682), .ZN(n8821) );
  AOI211_X1 U10151 ( .C1(n8686), .C2(n8819), .A(n8685), .B(n8821), .ZN(n8692)
         );
  AOI22_X1 U10152 ( .A1(n10224), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n8687), 
        .B2(n8698), .ZN(n8688) );
  OAI21_X1 U10153 ( .B1(n8689), .B2(n10200), .A(n8688), .ZN(n8690) );
  AOI21_X1 U10154 ( .B1(n8819), .B2(n8760), .A(n8690), .ZN(n8691) );
  OAI21_X1 U10155 ( .B1(n8692), .B2(n10224), .A(n8691), .ZN(P2_U3277) );
  XOR2_X1 U10156 ( .A(n8693), .B(n8703), .Z(n8830) );
  INV_X1 U10157 ( .A(n8694), .ZN(n8696) );
  AOI21_X1 U10158 ( .B1(n8826), .B2(n8696), .A(n8695), .ZN(n8827) );
  INV_X1 U10159 ( .A(n8697), .ZN(n8699) );
  AOI22_X1 U10160 ( .A1(n10224), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8699), 
        .B2(n8698), .ZN(n8700) );
  OAI21_X1 U10161 ( .B1(n8701), .B2(n10200), .A(n8700), .ZN(n8710) );
  INV_X1 U10162 ( .A(n8702), .ZN(n8706) );
  OAI21_X1 U10163 ( .B1(n8724), .B2(n8704), .A(n8703), .ZN(n8705) );
  NAND2_X1 U10164 ( .A1(n8706), .A2(n8705), .ZN(n8708) );
  AOI222_X1 U10165 ( .A1(n10193), .A2(n8708), .B1(n8707), .B2(n10190), .C1(
        n8742), .C2(n10189), .ZN(n8829) );
  NOR2_X1 U10166 ( .A1(n8829), .A2(n10224), .ZN(n8709) );
  AOI211_X1 U10167 ( .C1(n8827), .C2(n8711), .A(n8710), .B(n8709), .ZN(n8712)
         );
  OAI21_X1 U10168 ( .B1(n8830), .B2(n8713), .A(n8712), .ZN(P2_U3278) );
  OAI21_X1 U10169 ( .B1(n8715), .B2(n8717), .A(n8714), .ZN(n8832) );
  INV_X1 U10170 ( .A(n8832), .ZN(n8737) );
  NAND3_X1 U10171 ( .A1(n8718), .A2(n8717), .A3(n8716), .ZN(n8719) );
  NAND2_X1 U10172 ( .A1(n8719), .A2(n10193), .ZN(n8723) );
  AOI22_X1 U10173 ( .A1(n10190), .A2(n8721), .B1(n8720), .B2(n10189), .ZN(
        n8722) );
  OAI21_X1 U10174 ( .B1(n8724), .B2(n8723), .A(n8722), .ZN(n8729) );
  INV_X1 U10175 ( .A(n8725), .ZN(n8727) );
  XOR2_X1 U10176 ( .A(n8754), .B(n8831), .Z(n8726) );
  AOI21_X1 U10177 ( .B1(n8852), .B2(n8726), .A(n8729), .ZN(n8833) );
  OAI21_X1 U10178 ( .B1(n8737), .B2(n8727), .A(n8833), .ZN(n8728) );
  OAI211_X1 U10179 ( .C1(n8730), .C2(n8729), .A(n8728), .B(n10222), .ZN(n8735)
         );
  OAI22_X1 U10180 ( .A1(n10222), .A2(n8732), .B1(n8731), .B2(n10218), .ZN(
        n8733) );
  AOI21_X1 U10181 ( .B1(n8831), .B2(n10183), .A(n8733), .ZN(n8734) );
  OAI211_X1 U10182 ( .C1(n8737), .C2(n8736), .A(n8735), .B(n8734), .ZN(
        P2_U3279) );
  AND2_X1 U10183 ( .A1(n8738), .A2(n8744), .ZN(n8739) );
  OR2_X1 U10184 ( .A1(n8740), .A2(n8739), .ZN(n8751) );
  OR2_X1 U10185 ( .A1(n8751), .A2(n8741), .ZN(n8750) );
  AOI22_X1 U10186 ( .A1(n10189), .A2(n8743), .B1(n8742), .B2(n10190), .ZN(
        n8749) );
  INV_X1 U10187 ( .A(n8744), .ZN(n8745) );
  XNOR2_X1 U10188 ( .A(n8746), .B(n8745), .ZN(n8747) );
  NAND2_X1 U10189 ( .A1(n8747), .A2(n10193), .ZN(n8748) );
  INV_X1 U10190 ( .A(n8751), .ZN(n8840) );
  NAND2_X1 U10191 ( .A1(n8752), .A2(n8836), .ZN(n8753) );
  NAND2_X1 U10192 ( .A1(n8754), .A2(n8753), .ZN(n8838) );
  OAI22_X1 U10193 ( .A1(n10222), .A2(n8756), .B1(n8755), .B2(n10218), .ZN(
        n8757) );
  AOI21_X1 U10194 ( .B1(n8836), .B2(n10183), .A(n8757), .ZN(n8758) );
  OAI21_X1 U10195 ( .B1(n8838), .B2(n10219), .A(n8758), .ZN(n8759) );
  AOI21_X1 U10196 ( .B1(n8840), .B2(n8760), .A(n8759), .ZN(n8761) );
  OAI21_X1 U10197 ( .B1(n8842), .B2(n10224), .A(n8761), .ZN(P2_U3280) );
  NAND2_X1 U10198 ( .A1(n8762), .A2(n8851), .ZN(n8763) );
  OAI211_X1 U10199 ( .C1(n8764), .C2(n10298), .A(n8763), .B(n8767), .ZN(n8859)
         );
  MUX2_X1 U10200 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8859), .S(n10319), .Z(
        P2_U3551) );
  NAND3_X1 U10201 ( .A1(n8766), .A2(n8852), .A3(n8765), .ZN(n8768) );
  OAI211_X1 U10202 ( .C1(n8769), .C2(n10296), .A(n8768), .B(n8767), .ZN(n8860)
         );
  MUX2_X1 U10203 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8860), .S(n10319), .Z(
        P2_U3550) );
  AOI22_X1 U10204 ( .A1(n8772), .A2(n8852), .B1(n8851), .B2(n8771), .ZN(n8773)
         );
  NAND2_X1 U10205 ( .A1(n8776), .A2(n8775), .ZN(n8861) );
  MUX2_X1 U10206 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8861), .S(n10319), .Z(
        P2_U3548) );
  AOI22_X1 U10207 ( .A1(n8778), .A2(n8852), .B1(n8851), .B2(n8777), .ZN(n8779)
         );
  OAI211_X1 U10208 ( .C1(n8781), .C2(n8848), .A(n8780), .B(n8779), .ZN(n8862)
         );
  MUX2_X1 U10209 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8862), .S(n10319), .Z(
        P2_U3547) );
  AOI21_X1 U10210 ( .B1(n8851), .B2(n8783), .A(n8782), .ZN(n8784) );
  OAI211_X1 U10211 ( .C1(n8786), .C2(n8848), .A(n8785), .B(n8784), .ZN(n8863)
         );
  MUX2_X1 U10212 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8863), .S(n10319), .Z(
        P2_U3546) );
  AOI211_X1 U10213 ( .C1(n8851), .C2(n8789), .A(n8788), .B(n8787), .ZN(n8790)
         );
  OAI21_X1 U10214 ( .B1(n8791), .B2(n8848), .A(n8790), .ZN(n8864) );
  MUX2_X1 U10215 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8864), .S(n10319), .Z(
        P2_U3545) );
  AOI22_X1 U10216 ( .A1(n8793), .A2(n8852), .B1(n8851), .B2(n8792), .ZN(n8794)
         );
  OAI211_X1 U10217 ( .C1(n8796), .C2(n8848), .A(n8795), .B(n8794), .ZN(n8865)
         );
  MUX2_X1 U10218 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8865), .S(n10319), .Z(
        P2_U3544) );
  NAND2_X1 U10219 ( .A1(n8797), .A2(n10302), .ZN(n8802) );
  AOI22_X1 U10220 ( .A1(n8799), .A2(n8852), .B1(n8851), .B2(n8798), .ZN(n8800)
         );
  OAI211_X1 U10221 ( .C1(n8803), .C2(n8802), .A(n8801), .B(n8800), .ZN(n8866)
         );
  MUX2_X1 U10222 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8866), .S(n10319), .Z(
        P2_U3543) );
  AOI22_X1 U10223 ( .A1(n8805), .A2(n8852), .B1(n8851), .B2(n8804), .ZN(n8806)
         );
  OAI211_X1 U10224 ( .C1(n8808), .C2(n8848), .A(n8807), .B(n8806), .ZN(n8867)
         );
  MUX2_X1 U10225 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8867), .S(n10319), .Z(
        P2_U3542) );
  AOI22_X1 U10226 ( .A1(n8810), .A2(n8852), .B1(n8851), .B2(n8809), .ZN(n8811)
         );
  OAI211_X1 U10227 ( .C1(n8848), .C2(n8813), .A(n8812), .B(n8811), .ZN(n8868)
         );
  MUX2_X1 U10228 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8868), .S(n10319), .Z(
        P2_U3541) );
  AOI22_X1 U10229 ( .A1(n8815), .A2(n8852), .B1(n8851), .B2(n8814), .ZN(n8816)
         );
  OAI211_X1 U10230 ( .C1(n8848), .C2(n8818), .A(n8817), .B(n8816), .ZN(n8869)
         );
  MUX2_X1 U10231 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8869), .S(n10319), .Z(
        P2_U3540) );
  INV_X1 U10232 ( .A(n8819), .ZN(n8825) );
  INV_X1 U10233 ( .A(n8820), .ZN(n8822) );
  AOI211_X1 U10234 ( .C1(n8851), .C2(n8823), .A(n8822), .B(n8821), .ZN(n8824)
         );
  OAI21_X1 U10235 ( .B1(n8848), .B2(n8825), .A(n8824), .ZN(n8870) );
  MUX2_X1 U10236 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n8870), .S(n10319), .Z(
        P2_U3539) );
  AOI22_X1 U10237 ( .A1(n8827), .A2(n8852), .B1(n8851), .B2(n8826), .ZN(n8828)
         );
  OAI211_X1 U10238 ( .C1(n8830), .C2(n8848), .A(n8829), .B(n8828), .ZN(n8871)
         );
  MUX2_X1 U10239 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8871), .S(n10319), .Z(
        P2_U3538) );
  INV_X1 U10240 ( .A(n8831), .ZN(n8835) );
  NAND2_X1 U10241 ( .A1(n8832), .A2(n10302), .ZN(n8834) );
  OAI211_X1 U10242 ( .C1(n8835), .C2(n10296), .A(n8834), .B(n8833), .ZN(n8872)
         );
  MUX2_X1 U10243 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8872), .S(n10319), .Z(
        P2_U3537) );
  INV_X1 U10244 ( .A(n8836), .ZN(n8837) );
  OAI22_X1 U10245 ( .A1(n8838), .A2(n10298), .B1(n8837), .B2(n10296), .ZN(
        n8839) );
  AOI21_X1 U10246 ( .B1(n8840), .B2(n10293), .A(n8839), .ZN(n8841) );
  NAND2_X1 U10247 ( .A1(n8842), .A2(n8841), .ZN(n8873) );
  MUX2_X1 U10248 ( .A(n8873), .B(P2_REG1_REG_16__SCAN_IN), .S(n10317), .Z(
        P2_U3536) );
  INV_X1 U10249 ( .A(n8843), .ZN(n8849) );
  AOI22_X1 U10250 ( .A1(n8845), .A2(n8852), .B1(n8851), .B2(n8844), .ZN(n8846)
         );
  OAI211_X1 U10251 ( .C1(n8849), .C2(n8848), .A(n8847), .B(n8846), .ZN(n8874)
         );
  MUX2_X1 U10252 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8874), .S(n10319), .Z(
        P2_U3535) );
  AOI22_X1 U10253 ( .A1(n8853), .A2(n8852), .B1(n8851), .B2(n8850), .ZN(n8854)
         );
  OAI21_X1 U10254 ( .B1(n8856), .B2(n8855), .A(n8854), .ZN(n8857) );
  OR2_X1 U10255 ( .A1(n8858), .A2(n8857), .ZN(n8875) );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8875), .S(n10319), .Z(
        P2_U3533) );
  MUX2_X1 U10257 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8859), .S(n10306), .Z(
        P2_U3519) );
  MUX2_X1 U10258 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8860), .S(n10306), .Z(
        P2_U3518) );
  MUX2_X1 U10259 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8861), .S(n10306), .Z(
        P2_U3516) );
  MUX2_X1 U10260 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8862), .S(n10306), .Z(
        P2_U3515) );
  MUX2_X1 U10261 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8863), .S(n10306), .Z(
        P2_U3514) );
  MUX2_X1 U10262 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8864), .S(n10306), .Z(
        P2_U3513) );
  MUX2_X1 U10263 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8865), .S(n10306), .Z(
        P2_U3512) );
  MUX2_X1 U10264 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8866), .S(n10306), .Z(
        P2_U3511) );
  MUX2_X1 U10265 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8867), .S(n10306), .Z(
        P2_U3510) );
  MUX2_X1 U10266 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8868), .S(n10306), .Z(
        P2_U3509) );
  MUX2_X1 U10267 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8869), .S(n10306), .Z(
        P2_U3508) );
  MUX2_X1 U10268 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n8870), .S(n10306), .Z(
        P2_U3507) );
  MUX2_X1 U10269 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8871), .S(n10306), .Z(
        P2_U3505) );
  MUX2_X1 U10270 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8872), .S(n10306), .Z(
        P2_U3502) );
  MUX2_X1 U10271 ( .A(n8873), .B(P2_REG0_REG_16__SCAN_IN), .S(n10304), .Z(
        P2_U3499) );
  MUX2_X1 U10272 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8874), .S(n10306), .Z(
        P2_U3496) );
  MUX2_X1 U10273 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n8875), .S(n10306), .Z(
        P2_U3490) );
  INV_X1 U10274 ( .A(n8876), .ZN(n9776) );
  NAND3_X1 U10275 ( .A1(n4592), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n8877) );
  OAI22_X1 U10276 ( .A1(n8878), .A2(n8877), .B1(n9647), .B2(n8888), .ZN(n8879)
         );
  INV_X1 U10277 ( .A(n8879), .ZN(n8880) );
  OAI21_X1 U10278 ( .B1(n9776), .B2(n8883), .A(n8880), .ZN(P2_U3327) );
  OAI222_X1 U10279 ( .A1(n8888), .A2(n9722), .B1(n8883), .B2(n8882), .C1(n8881), .C2(P2_U3152), .ZN(P2_U3328) );
  NAND2_X1 U10280 ( .A1(n9778), .A2(n8884), .ZN(n8886) );
  OAI211_X1 U10281 ( .C1(n8888), .C2(n8887), .A(n8886), .B(n8885), .ZN(
        P2_U3330) );
  MUX2_X1 U10282 ( .A(n8889), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10283 ( .A1(n8891), .A2(n8890), .ZN(n8892) );
  XOR2_X1 U10284 ( .A(n8893), .B(n8892), .Z(n8899) );
  OAI22_X1 U10285 ( .A1(n9005), .A2(n9356), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8894), .ZN(n8895) );
  AOI21_X1 U10286 ( .B1(n9007), .B2(n9311), .A(n8895), .ZN(n8896) );
  OAI21_X1 U10287 ( .B1(n9021), .B2(n9348), .A(n8896), .ZN(n8897) );
  AOI21_X1 U10288 ( .B1(n9351), .B2(n9023), .A(n8897), .ZN(n8898) );
  OAI21_X1 U10289 ( .B1(n8899), .B2(n9025), .A(n8898), .ZN(P1_U3213) );
  INV_X1 U10290 ( .A(n8900), .ZN(n8905) );
  OAI21_X1 U10291 ( .B1(n8902), .B2(n8904), .A(n8901), .ZN(n8903) );
  OAI21_X1 U10292 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8906) );
  NAND2_X1 U10293 ( .A1(n8906), .A2(n8951), .ZN(n8910) );
  NOR2_X1 U10294 ( .A1(n9021), .A2(n9199), .ZN(n8908) );
  OAI22_X1 U10295 ( .A1(n9017), .A2(n9175), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9668), .ZN(n8907) );
  AOI211_X1 U10296 ( .C1(n9019), .C2(n9228), .A(n8908), .B(n8907), .ZN(n8909)
         );
  OAI211_X1 U10297 ( .C1(n4710), .C2(n8958), .A(n8910), .B(n8909), .ZN(
        P1_U3214) );
  XOR2_X1 U10298 ( .A(n8912), .B(n8911), .Z(n8913) );
  XNOR2_X1 U10299 ( .A(n8914), .B(n8913), .ZN(n8920) );
  NAND2_X1 U10300 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9110) );
  OAI21_X1 U10301 ( .B1(n9005), .B2(n8915), .A(n9110), .ZN(n8916) );
  AOI21_X1 U10302 ( .B1(n9007), .B2(n9263), .A(n8916), .ZN(n8917) );
  OAI21_X1 U10303 ( .B1(n9021), .B2(n9267), .A(n8917), .ZN(n8918) );
  AOI21_X1 U10304 ( .B1(n9442), .B2(n9023), .A(n8918), .ZN(n8919) );
  OAI21_X1 U10305 ( .B1(n8920), .B2(n9025), .A(n8919), .ZN(P1_U3217) );
  NAND2_X1 U10306 ( .A1(n9241), .A2(n9822), .ZN(n9434) );
  XNOR2_X1 U10307 ( .A(n8922), .B(n8921), .ZN(n8923) );
  NAND2_X1 U10308 ( .A1(n8923), .A2(n8951), .ZN(n8928) );
  NOR2_X1 U10309 ( .A1(n9021), .A2(n9234), .ZN(n8926) );
  OAI22_X1 U10310 ( .A1(n9017), .A2(n8924), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9746), .ZN(n8925) );
  AOI211_X1 U10311 ( .C1(n9019), .C2(n9263), .A(n8926), .B(n8925), .ZN(n8927)
         );
  OAI211_X1 U10312 ( .C1(n8929), .C2(n9434), .A(n8928), .B(n8927), .ZN(
        P1_U3221) );
  XOR2_X1 U10313 ( .A(n8931), .B(n8930), .Z(n8936) );
  NAND2_X1 U10314 ( .A1(n8962), .A2(n9177), .ZN(n8933) );
  AOI22_X1 U10315 ( .A1(n9007), .A2(n9143), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8932) );
  OAI211_X1 U10316 ( .C1(n9175), .C2(n9005), .A(n8933), .B(n8932), .ZN(n8934)
         );
  AOI21_X1 U10317 ( .B1(n9412), .B2(n9023), .A(n8934), .ZN(n8935) );
  OAI21_X1 U10318 ( .B1(n8936), .B2(n9025), .A(n8935), .ZN(P1_U3223) );
  INV_X1 U10319 ( .A(n8937), .ZN(n8941) );
  NAND2_X1 U10320 ( .A1(n4437), .A2(n8940), .ZN(n8938) );
  AOI22_X1 U10321 ( .A1(n8941), .A2(n8940), .B1(n8939), .B2(n8938), .ZN(n8947)
         );
  NOR2_X1 U10322 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8942), .ZN(n9071) );
  NOR2_X1 U10323 ( .A1(n9005), .A2(n9357), .ZN(n8943) );
  AOI211_X1 U10324 ( .C1(n9007), .C2(n9310), .A(n9071), .B(n8943), .ZN(n8944)
         );
  OAI21_X1 U10325 ( .B1(n9021), .B2(n9316), .A(n8944), .ZN(n8945) );
  AOI21_X1 U10326 ( .B1(n9318), .B2(n9023), .A(n8945), .ZN(n8946) );
  OAI21_X1 U10327 ( .B1(n8947), .B2(n9025), .A(n8946), .ZN(P1_U3224) );
  OAI21_X1 U10328 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8952) );
  NAND2_X1 U10329 ( .A1(n8952), .A2(n8951), .ZN(n8957) );
  NOR2_X1 U10330 ( .A1(n9021), .A2(n9292), .ZN(n8955) );
  OAI22_X1 U10331 ( .A1(n9005), .A2(n9016), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8953), .ZN(n8954) );
  AOI211_X1 U10332 ( .C1(n9007), .C2(n9298), .A(n8955), .B(n8954), .ZN(n8956)
         );
  OAI211_X1 U10333 ( .C1(n4723), .C2(n8958), .A(n8957), .B(n8956), .ZN(
        P1_U3226) );
  AOI21_X1 U10334 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(n8967) );
  NAND2_X1 U10335 ( .A1(n8962), .A2(n9190), .ZN(n8964) );
  AOI22_X1 U10336 ( .A1(n9007), .A2(n9029), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n8963) );
  OAI211_X1 U10337 ( .C1(n9187), .C2(n9005), .A(n8964), .B(n8963), .ZN(n8965)
         );
  AOI21_X1 U10338 ( .B1(n9419), .B2(n9023), .A(n8965), .ZN(n8966) );
  OAI21_X1 U10339 ( .B1(n8967), .B2(n9025), .A(n8966), .ZN(P1_U3227) );
  INV_X1 U10340 ( .A(n8968), .ZN(n8972) );
  NAND2_X1 U10341 ( .A1(n4484), .A2(n8971), .ZN(n8969) );
  AOI22_X1 U10342 ( .A1(n8972), .A2(n8971), .B1(n8970), .B2(n8969), .ZN(n8977)
         );
  AOI22_X1 U10343 ( .A1(n9007), .A2(n9212), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8974) );
  NAND2_X1 U10344 ( .A1(n9019), .A2(n9284), .ZN(n8973) );
  OAI211_X1 U10345 ( .C1(n9021), .C2(n9253), .A(n8974), .B(n8973), .ZN(n8975)
         );
  AOI21_X1 U10346 ( .B1(n9439), .B2(n9023), .A(n8975), .ZN(n8976) );
  OAI21_X1 U10347 ( .B1(n8977), .B2(n9025), .A(n8976), .ZN(P1_U3231) );
  NAND2_X1 U10348 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  XOR2_X1 U10349 ( .A(n8981), .B(n8980), .Z(n8987) );
  OAI22_X1 U10350 ( .A1(n9017), .A2(n9187), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8982), .ZN(n8983) );
  AOI21_X1 U10351 ( .B1(n9019), .B2(n9212), .A(n8983), .ZN(n8984) );
  OAI21_X1 U10352 ( .B1(n9021), .B2(n9217), .A(n8984), .ZN(n8985) );
  AOI21_X1 U10353 ( .B1(n9427), .B2(n9023), .A(n8985), .ZN(n8986) );
  OAI21_X1 U10354 ( .B1(n8987), .B2(n9025), .A(n8986), .ZN(P1_U3233) );
  NOR2_X1 U10355 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9622), .ZN(n9928) );
  AOI21_X1 U10356 ( .B1(n9019), .B2(n9033), .A(n9928), .ZN(n8989) );
  NAND2_X1 U10357 ( .A1(n9007), .A2(n9031), .ZN(n8988) );
  OAI211_X1 U10358 ( .C1(n9021), .C2(n8990), .A(n8989), .B(n8988), .ZN(n8999)
         );
  AND2_X1 U10359 ( .A1(n4486), .A2(n8992), .ZN(n8996) );
  XNOR2_X1 U10360 ( .A(n8994), .B(n8993), .ZN(n8995) );
  XNOR2_X1 U10361 ( .A(n8996), .B(n8995), .ZN(n8997) );
  NOR2_X1 U10362 ( .A1(n8997), .A2(n9025), .ZN(n8998) );
  AOI211_X1 U10363 ( .C1(n9023), .C2(n9468), .A(n8999), .B(n8998), .ZN(n9000)
         );
  INV_X1 U10364 ( .A(n9000), .ZN(P1_U3234) );
  NAND2_X1 U10365 ( .A1(n9002), .A2(n9001), .ZN(n9003) );
  XOR2_X1 U10366 ( .A(n9004), .B(n9003), .Z(n9011) );
  NAND2_X1 U10367 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9943) );
  OAI21_X1 U10368 ( .B1(n9005), .B2(n5711), .A(n9943), .ZN(n9006) );
  AOI21_X1 U10369 ( .B1(n9007), .B2(n9284), .A(n9006), .ZN(n9008) );
  OAI21_X1 U10370 ( .B1(n9021), .B2(n9278), .A(n9008), .ZN(n9009) );
  AOI21_X1 U10371 ( .B1(n9447), .B2(n9023), .A(n9009), .ZN(n9010) );
  OAI21_X1 U10372 ( .B1(n9011), .B2(n9025), .A(n9010), .ZN(P1_U3236) );
  NAND2_X1 U10373 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  XOR2_X1 U10374 ( .A(n9015), .B(n9014), .Z(n9026) );
  AND2_X1 U10375 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9050) );
  NOR2_X1 U10376 ( .A1(n9017), .A2(n9016), .ZN(n9018) );
  AOI211_X1 U10377 ( .C1(n9019), .C2(n9327), .A(n9050), .B(n9018), .ZN(n9020)
         );
  OAI21_X1 U10378 ( .B1(n9021), .B2(n9334), .A(n9020), .ZN(n9022) );
  AOI21_X1 U10379 ( .B1(n9340), .B2(n9023), .A(n9022), .ZN(n9024) );
  OAI21_X1 U10380 ( .B1(n9026), .B2(n9025), .A(n9024), .ZN(P1_U3239) );
  MUX2_X1 U10381 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n4859), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10382 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9027), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10383 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9137), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10384 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9028), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10385 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9143), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10386 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9029), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10387 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9204), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10388 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9211), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10389 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9228), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10390 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9212), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10391 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9263), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10392 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9284), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10393 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9298), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10394 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9310), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10395 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9328), .S(P1_U4006), .Z(
        P1_U3571) );
  MUX2_X1 U10396 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9311), .S(P1_U4006), .Z(
        P1_U3570) );
  MUX2_X1 U10397 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9327), .S(P1_U4006), .Z(
        P1_U3569) );
  MUX2_X1 U10398 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9030), .S(P1_U4006), .Z(
        P1_U3568) );
  MUX2_X1 U10399 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9031), .S(P1_U4006), .Z(
        P1_U3567) );
  MUX2_X1 U10400 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9032), .S(P1_U4006), .Z(
        P1_U3566) );
  MUX2_X1 U10401 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9033), .S(P1_U4006), .Z(
        P1_U3565) );
  MUX2_X1 U10402 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9034), .S(P1_U4006), .Z(
        P1_U3564) );
  MUX2_X1 U10403 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9035), .S(P1_U4006), .Z(
        P1_U3563) );
  MUX2_X1 U10404 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9036), .S(P1_U4006), .Z(
        P1_U3562) );
  MUX2_X1 U10405 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9037), .S(P1_U4006), .Z(
        P1_U3561) );
  MUX2_X1 U10406 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9986), .S(P1_U4006), .Z(
        P1_U3560) );
  MUX2_X1 U10407 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9038), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10408 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n10009), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10409 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6542), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10410 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9039), .S(P1_U4006), .Z(
        P1_U3556) );
  INV_X1 U10411 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9054) );
  NOR2_X1 U10412 ( .A1(n9041), .A2(n9040), .ZN(n9043) );
  NOR2_X1 U10413 ( .A1(n9043), .A2(n9042), .ZN(n9055) );
  AOI211_X1 U10414 ( .C1(n9044), .C2(n9335), .A(n9056), .B(n9944), .ZN(n9045)
         );
  INV_X1 U10415 ( .A(n9045), .ZN(n9053) );
  OAI21_X1 U10416 ( .B1(n9047), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9046), .ZN(
        n9062) );
  XNOR2_X1 U10417 ( .A(n9063), .B(n9062), .ZN(n9048) );
  INV_X1 U10418 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9837) );
  NOR2_X1 U10419 ( .A1(n9837), .A2(n9048), .ZN(n9064) );
  AOI211_X1 U10420 ( .C1(n9048), .C2(n9837), .A(n9064), .B(n9907), .ZN(n9049)
         );
  AOI211_X1 U10421 ( .C1(n9950), .C2(n9051), .A(n9050), .B(n9049), .ZN(n9052)
         );
  OAI211_X1 U10422 ( .C1(n9942), .C2(n9054), .A(n9053), .B(n9052), .ZN(
        P1_U3256) );
  NOR2_X1 U10423 ( .A1(n9055), .A2(n9063), .ZN(n9057) );
  OR2_X1 U10424 ( .A1(n9083), .A2(n9058), .ZN(n9060) );
  NAND2_X1 U10425 ( .A1(n9083), .A2(n9058), .ZN(n9059) );
  AND2_X1 U10426 ( .A1(n9060), .A2(n9059), .ZN(n9061) );
  AOI211_X1 U10427 ( .C1(n4439), .C2(n9061), .A(n9078), .B(n9944), .ZN(n9077)
         );
  NOR2_X1 U10428 ( .A1(n9063), .A2(n9062), .ZN(n9065) );
  INV_X1 U10429 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9066) );
  OR2_X1 U10430 ( .A1(n9083), .A2(n9066), .ZN(n9068) );
  NAND2_X1 U10431 ( .A1(n9083), .A2(n9066), .ZN(n9067) );
  AND2_X1 U10432 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  NOR2_X1 U10433 ( .A1(n9070), .A2(n9069), .ZN(n9082) );
  AOI211_X1 U10434 ( .C1(n9070), .C2(n9069), .A(n9082), .B(n9907), .ZN(n9076)
         );
  INV_X1 U10435 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9074) );
  INV_X1 U10436 ( .A(n9071), .ZN(n9073) );
  NAND2_X1 U10437 ( .A1(n9950), .A2(n9083), .ZN(n9072) );
  OAI211_X1 U10438 ( .C1(n9942), .C2(n9074), .A(n9073), .B(n9072), .ZN(n9075)
         );
  OR3_X1 U10439 ( .A1(n9077), .A2(n9076), .A3(n9075), .ZN(P1_U3257) );
  AOI21_X1 U10440 ( .B1(n9083), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9078), .ZN(
        n9081) );
  NAND2_X1 U10441 ( .A1(n9102), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9079) );
  OAI21_X1 U10442 ( .B1(n9102), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9079), .ZN(
        n9080) );
  NOR2_X1 U10443 ( .A1(n9081), .A2(n9080), .ZN(n9095) );
  AOI211_X1 U10444 ( .C1(n9081), .C2(n9080), .A(n9095), .B(n9944), .ZN(n9093)
         );
  INV_X1 U10445 ( .A(n9102), .ZN(n9090) );
  AOI21_X1 U10446 ( .B1(n9083), .B2(P1_REG1_REG_16__SCAN_IN), .A(n9082), .ZN(
        n9086) );
  MUX2_X1 U10447 ( .A(n9084), .B(P1_REG1_REG_17__SCAN_IN), .S(n9102), .Z(n9085) );
  NOR2_X1 U10448 ( .A1(n9086), .A2(n9085), .ZN(n9101) );
  AOI211_X1 U10449 ( .C1(n9086), .C2(n9085), .A(n9101), .B(n9907), .ZN(n9087)
         );
  INV_X1 U10450 ( .A(n9087), .ZN(n9089) );
  NAND2_X1 U10451 ( .A1(P1_REG3_REG_17__SCAN_IN), .A2(P1_U3084), .ZN(n9088) );
  OAI211_X1 U10452 ( .C1(n9091), .C2(n9090), .A(n9089), .B(n9088), .ZN(n9092)
         );
  AOI211_X1 U10453 ( .C1(P1_ADDR_REG_17__SCAN_IN), .C2(n9955), .A(n9093), .B(
        n9092), .ZN(n9094) );
  INV_X1 U10454 ( .A(n9094), .ZN(P1_U3258) );
  AOI21_X1 U10455 ( .B1(n9102), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9095), .ZN(
        n9947) );
  NOR2_X1 U10456 ( .A1(n9951), .A2(n9096), .ZN(n9097) );
  AOI21_X1 U10457 ( .B1(n9951), .B2(n9096), .A(n9097), .ZN(n9946) );
  NOR2_X1 U10458 ( .A1(n9947), .A2(n9946), .ZN(n9945) );
  AOI21_X1 U10459 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9951), .A(n9945), .ZN(
        n9098) );
  XNOR2_X1 U10460 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9098), .ZN(n9109) );
  INV_X1 U10461 ( .A(n9109), .ZN(n9104) );
  AOI22_X1 U10462 ( .A1(n9951), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9100), .B2(
        n9099), .ZN(n9954) );
  NAND2_X1 U10463 ( .A1(n9954), .A2(n9953), .ZN(n9952) );
  OAI21_X1 U10464 ( .B1(n9951), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9952), .ZN(
        n9103) );
  XOR2_X1 U10465 ( .A(n9103), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9106) );
  INV_X1 U10466 ( .A(n9105), .ZN(n9108) );
  AOI21_X1 U10467 ( .B1(n9106), .B2(n9956), .A(n9950), .ZN(n9107) );
  XNOR2_X1 U10468 ( .A(n9390), .B(n9115), .ZN(n9388) );
  NAND2_X1 U10469 ( .A1(n9388), .A2(n10003), .ZN(n9114) );
  NAND2_X1 U10470 ( .A1(n9112), .A2(n9111), .ZN(n9817) );
  NOR2_X1 U10471 ( .A1(n9387), .A2(n9817), .ZN(n9119) );
  AOI21_X1 U10472 ( .B1(n10021), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9119), .ZN(
        n9113) );
  OAI211_X1 U10473 ( .C1(n9390), .C2(n10029), .A(n9114), .B(n9113), .ZN(
        P1_U3261) );
  OAI21_X1 U10474 ( .B1(n9117), .B2(n9116), .A(n9115), .ZN(n9818) );
  NOR2_X1 U10475 ( .A1(n9321), .A2(n9118), .ZN(n9120) );
  AOI211_X1 U10476 ( .C1(n9821), .C2(n9350), .A(n9120), .B(n9119), .ZN(n9121)
         );
  OAI21_X1 U10477 ( .B1(n9818), .B2(n10032), .A(n9121), .ZN(P1_U3262) );
  AOI21_X1 U10478 ( .B1(n9122), .B2(n9128), .A(n9989), .ZN(n9126) );
  OAI22_X1 U10479 ( .A1(n9164), .A2(n10012), .B1(n9123), .B2(n10010), .ZN(
        n9124) );
  AOI21_X1 U10480 ( .B1(n9126), .B2(n9125), .A(n9124), .ZN(n9399) );
  INV_X1 U10481 ( .A(n9400), .ZN(n9134) );
  NAND2_X1 U10482 ( .A1(n9144), .A2(n9396), .ZN(n9129) );
  NAND2_X1 U10483 ( .A1(n9397), .A2(n10003), .ZN(n9132) );
  AOI22_X1 U10484 ( .A1(n10021), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n9130), 
        .B2(n10020), .ZN(n9131) );
  OAI211_X1 U10485 ( .C1(n4719), .C2(n10029), .A(n9132), .B(n9131), .ZN(n9133)
         );
  AOI21_X1 U10486 ( .B1(n9134), .B2(n9363), .A(n9133), .ZN(n9135) );
  OAI21_X1 U10487 ( .B1(n10021), .B2(n9399), .A(n9135), .ZN(P1_U3263) );
  XNOR2_X1 U10488 ( .A(n4420), .B(n9136), .ZN(n9405) );
  AND2_X1 U10489 ( .A1(n9137), .A2(n9985), .ZN(n9142) );
  AOI211_X1 U10490 ( .C1(n9140), .C2(n9139), .A(n9989), .B(n9138), .ZN(n9141)
         );
  INV_X1 U10491 ( .A(n9404), .ZN(n9152) );
  INV_X1 U10492 ( .A(n9155), .ZN(n9146) );
  INV_X1 U10493 ( .A(n9144), .ZN(n9145) );
  AOI21_X1 U10494 ( .B1(n9401), .B2(n9146), .A(n9145), .ZN(n9402) );
  NAND2_X1 U10495 ( .A1(n9402), .A2(n10003), .ZN(n9149) );
  AOI22_X1 U10496 ( .A1(n10021), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9147), 
        .B2(n10020), .ZN(n9148) );
  OAI211_X1 U10497 ( .C1(n9150), .C2(n10029), .A(n9149), .B(n9148), .ZN(n9151)
         );
  AOI21_X1 U10498 ( .B1(n9152), .B2(n9321), .A(n9151), .ZN(n9153) );
  OAI21_X1 U10499 ( .B1(n9323), .B2(n9405), .A(n9153), .ZN(P1_U3264) );
  XOR2_X1 U10500 ( .A(n9162), .B(n9154), .Z(n9410) );
  AOI211_X1 U10501 ( .C1(n9408), .C2(n9168), .A(n10118), .B(n9155), .ZN(n9407)
         );
  INV_X1 U10502 ( .A(n9156), .ZN(n9157) );
  AOI22_X1 U10503 ( .A1(n10021), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9157), 
        .B2(n10020), .ZN(n9158) );
  OAI21_X1 U10504 ( .B1(n9159), .B2(n10029), .A(n9158), .ZN(n9160) );
  AOI21_X1 U10505 ( .B1(n9407), .B2(n9258), .A(n9160), .ZN(n9166) );
  XOR2_X1 U10506 ( .A(n9162), .B(n9161), .Z(n9163) );
  OAI222_X1 U10507 ( .A1(n10010), .A2(n9164), .B1(n10012), .B2(n9186), .C1(
        n9163), .C2(n9989), .ZN(n9406) );
  NAND2_X1 U10508 ( .A1(n9406), .A2(n9321), .ZN(n9165) );
  OAI211_X1 U10509 ( .C1(n9410), .C2(n9323), .A(n9166), .B(n9165), .ZN(
        P1_U3265) );
  XNOR2_X1 U10510 ( .A(n9167), .B(n9173), .ZN(n9416) );
  INV_X1 U10511 ( .A(n9168), .ZN(n9169) );
  AOI21_X1 U10512 ( .B1(n9412), .B2(n9188), .A(n9169), .ZN(n9413) );
  INV_X1 U10513 ( .A(n9412), .ZN(n9171) );
  INV_X1 U10514 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9170) );
  OAI22_X1 U10515 ( .A1(n9171), .A2(n10029), .B1(n9170), .B2(n9321), .ZN(n9180) );
  AOI21_X1 U10516 ( .B1(n4436), .B2(n9173), .A(n9172), .ZN(n9174) );
  OAI222_X1 U10517 ( .A1(n10010), .A2(n9176), .B1(n10012), .B2(n9175), .C1(
        n9989), .C2(n9174), .ZN(n9411) );
  AOI21_X1 U10518 ( .B1(n9177), .B2(n10020), .A(n9411), .ZN(n9178) );
  NOR2_X1 U10519 ( .A1(n9178), .A2(n9387), .ZN(n9179) );
  AOI211_X1 U10520 ( .C1(n9413), .C2(n10003), .A(n9180), .B(n9179), .ZN(n9181)
         );
  OAI21_X1 U10521 ( .B1(n9416), .B2(n9323), .A(n9181), .ZN(P1_U3266) );
  XNOR2_X1 U10522 ( .A(n9182), .B(n9184), .ZN(n9421) );
  AOI21_X1 U10523 ( .B1(n9184), .B2(n9183), .A(n4465), .ZN(n9185) );
  OAI222_X1 U10524 ( .A1(n10012), .A2(n9187), .B1(n10010), .B2(n9186), .C1(
        n9989), .C2(n9185), .ZN(n9417) );
  INV_X1 U10525 ( .A(n9188), .ZN(n9189) );
  AOI211_X1 U10526 ( .C1(n9419), .C2(n4712), .A(n10118), .B(n9189), .ZN(n9418)
         );
  INV_X1 U10527 ( .A(n9418), .ZN(n9193) );
  INV_X1 U10528 ( .A(n9190), .ZN(n9191) );
  OAI22_X1 U10529 ( .A1(n9193), .A2(n9192), .B1(n9994), .B2(n9191), .ZN(n9194)
         );
  OAI21_X1 U10530 ( .B1(n9417), .B2(n9194), .A(n9321), .ZN(n9196) );
  AOI22_X1 U10531 ( .A1(n9419), .A2(n9350), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9387), .ZN(n9195) );
  OAI211_X1 U10532 ( .C1(n9421), .C2(n9323), .A(n9196), .B(n9195), .ZN(
        P1_U3267) );
  XNOR2_X1 U10533 ( .A(n9197), .B(n9203), .ZN(n9426) );
  AOI21_X1 U10534 ( .B1(n9422), .B2(n9220), .A(n9198), .ZN(n9423) );
  INV_X1 U10535 ( .A(n9199), .ZN(n9200) );
  AOI22_X1 U10536 ( .A1(n10021), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9200), 
        .B2(n10020), .ZN(n9201) );
  OAI21_X1 U10537 ( .B1(n4710), .B2(n10029), .A(n9201), .ZN(n9207) );
  XOR2_X1 U10538 ( .A(n9203), .B(n9202), .Z(n9205) );
  AOI222_X1 U10539 ( .A1(n10019), .A2(n9205), .B1(n9228), .B2(n9987), .C1(
        n9204), .C2(n9985), .ZN(n9425) );
  NOR2_X1 U10540 ( .A1(n9425), .A2(n9387), .ZN(n9206) );
  AOI211_X1 U10541 ( .C1(n9423), .C2(n10003), .A(n9207), .B(n9206), .ZN(n9208)
         );
  OAI21_X1 U10542 ( .B1(n9426), .B2(n9323), .A(n9208), .ZN(P1_U3268) );
  NAND2_X1 U10543 ( .A1(n9227), .A2(n9209), .ZN(n9210) );
  XOR2_X1 U10544 ( .A(n9214), .B(n9210), .Z(n9213) );
  AOI222_X1 U10545 ( .A1(n10019), .A2(n9213), .B1(n9212), .B2(n9987), .C1(
        n9211), .C2(n9985), .ZN(n9430) );
  XOR2_X1 U10546 ( .A(n9215), .B(n9214), .Z(n9431) );
  NAND2_X1 U10547 ( .A1(n10021), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9216) );
  OAI21_X1 U10548 ( .B1(n9994), .B2(n9217), .A(n9216), .ZN(n9218) );
  AOI21_X1 U10549 ( .B1(n9427), .B2(n9350), .A(n9218), .ZN(n9222) );
  NAND2_X1 U10550 ( .A1(n9236), .A2(n9427), .ZN(n9219) );
  AND2_X1 U10551 ( .A1(n9220), .A2(n9219), .ZN(n9428) );
  NAND2_X1 U10552 ( .A1(n9428), .A2(n10003), .ZN(n9221) );
  OAI211_X1 U10553 ( .C1(n9431), .C2(n9323), .A(n9222), .B(n9221), .ZN(n9223)
         );
  INV_X1 U10554 ( .A(n9223), .ZN(n9224) );
  OAI21_X1 U10555 ( .B1(n10021), .B2(n9430), .A(n9224), .ZN(P1_U3269) );
  OR2_X1 U10556 ( .A1(n9225), .A2(n4777), .ZN(n9226) );
  NAND2_X1 U10557 ( .A1(n9227), .A2(n9226), .ZN(n9232) );
  NAND2_X1 U10558 ( .A1(n9228), .A2(n9985), .ZN(n9229) );
  OAI21_X1 U10559 ( .B1(n9230), .B2(n10012), .A(n9229), .ZN(n9231) );
  AOI21_X1 U10560 ( .B1(n9232), .B2(n10019), .A(n9231), .ZN(n9435) );
  XNOR2_X1 U10561 ( .A(n9233), .B(n4777), .ZN(n9432) );
  NAND2_X1 U10562 ( .A1(n9432), .A2(n9363), .ZN(n9243) );
  INV_X1 U10563 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9235) );
  OAI22_X1 U10564 ( .A1(n9321), .A2(n9235), .B1(n9234), .B2(n9994), .ZN(n9240)
         );
  OAI211_X1 U10565 ( .C1(n9237), .C2(n9252), .A(n9469), .B(n9236), .ZN(n9433)
         );
  INV_X1 U10566 ( .A(n9258), .ZN(n9238) );
  NOR2_X1 U10567 ( .A1(n9433), .A2(n9238), .ZN(n9239) );
  AOI211_X1 U10568 ( .C1(n9350), .C2(n9241), .A(n9240), .B(n9239), .ZN(n9242)
         );
  OAI211_X1 U10569 ( .C1(n10021), .C2(n9435), .A(n9243), .B(n9242), .ZN(
        P1_U3270) );
  XNOR2_X1 U10570 ( .A(n9244), .B(n9245), .ZN(n9441) );
  XOR2_X1 U10571 ( .A(n9246), .B(n9245), .Z(n9247) );
  OAI222_X1 U10572 ( .A1(n10010), .A2(n9249), .B1(n10012), .B2(n9248), .C1(
        n9247), .C2(n9989), .ZN(n9437) );
  NAND2_X1 U10573 ( .A1(n9437), .A2(n9321), .ZN(n9260) );
  NAND2_X1 U10574 ( .A1(n9266), .A2(n9439), .ZN(n9250) );
  NAND2_X1 U10575 ( .A1(n9250), .A2(n9469), .ZN(n9251) );
  NOR2_X1 U10576 ( .A1(n9252), .A2(n9251), .ZN(n9438) );
  OAI22_X1 U10577 ( .A1(n9321), .A2(n9254), .B1(n9253), .B2(n9994), .ZN(n9257)
         );
  NOR2_X1 U10578 ( .A1(n9255), .A2(n10029), .ZN(n9256) );
  AOI211_X1 U10579 ( .C1(n9438), .C2(n9258), .A(n9257), .B(n9256), .ZN(n9259)
         );
  OAI211_X1 U10580 ( .C1(n9441), .C2(n9323), .A(n9260), .B(n9259), .ZN(
        P1_U3271) );
  XNOR2_X1 U10581 ( .A(n9262), .B(n9261), .ZN(n9264) );
  AOI222_X1 U10582 ( .A1(n10019), .A2(n9264), .B1(n9298), .B2(n9987), .C1(
        n9263), .C2(n9985), .ZN(n9445) );
  OR2_X1 U10583 ( .A1(n9277), .A2(n9270), .ZN(n9265) );
  AND2_X1 U10584 ( .A1(n9266), .A2(n9265), .ZN(n9443) );
  INV_X1 U10585 ( .A(n9267), .ZN(n9268) );
  AOI22_X1 U10586 ( .A1(n10021), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9268), 
        .B2(n10020), .ZN(n9269) );
  OAI21_X1 U10587 ( .B1(n9270), .B2(n10029), .A(n9269), .ZN(n9274) );
  XNOR2_X1 U10588 ( .A(n4774), .B(n9271), .ZN(n9446) );
  NOR2_X1 U10589 ( .A1(n9446), .A2(n9323), .ZN(n9273) );
  AOI211_X1 U10590 ( .C1(n9443), .C2(n10003), .A(n9274), .B(n9273), .ZN(n9275)
         );
  OAI21_X1 U10591 ( .B1(n10021), .B2(n9445), .A(n9275), .ZN(P1_U3272) );
  XNOR2_X1 U10592 ( .A(n9276), .B(n9283), .ZN(n9451) );
  AOI21_X1 U10593 ( .B1(n9447), .B2(n4725), .A(n9277), .ZN(n9448) );
  INV_X1 U10594 ( .A(n9278), .ZN(n9279) );
  AOI22_X1 U10595 ( .A1(n10021), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9279), 
        .B2(n10020), .ZN(n9280) );
  OAI21_X1 U10596 ( .B1(n9281), .B2(n10029), .A(n9280), .ZN(n9287) );
  OAI21_X1 U10597 ( .B1(n4479), .B2(n9283), .A(n9282), .ZN(n9285) );
  AOI222_X1 U10598 ( .A1(n10019), .A2(n9285), .B1(n9310), .B2(n9987), .C1(
        n9284), .C2(n9985), .ZN(n9450) );
  NOR2_X1 U10599 ( .A1(n9450), .A2(n9387), .ZN(n9286) );
  AOI211_X1 U10600 ( .C1(n9448), .C2(n10003), .A(n9287), .B(n9286), .ZN(n9288)
         );
  OAI21_X1 U10601 ( .B1(n9323), .B2(n9451), .A(n9288), .ZN(P1_U3273) );
  XNOR2_X1 U10602 ( .A(n9290), .B(n9289), .ZN(n9456) );
  AOI21_X1 U10603 ( .B1(n9452), .B2(n9314), .A(n9291), .ZN(n9453) );
  INV_X1 U10604 ( .A(n9292), .ZN(n9293) );
  AOI22_X1 U10605 ( .A1(n10021), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9293), 
        .B2(n10020), .ZN(n9294) );
  OAI21_X1 U10606 ( .B1(n4723), .B2(n10029), .A(n9294), .ZN(n9302) );
  OAI211_X1 U10607 ( .C1(n9297), .C2(n9296), .A(n9295), .B(n10019), .ZN(n9300)
         );
  AOI22_X1 U10608 ( .A1(n9987), .A2(n9328), .B1(n9298), .B2(n9985), .ZN(n9299)
         );
  AND2_X1 U10609 ( .A1(n9300), .A2(n9299), .ZN(n9455) );
  NOR2_X1 U10610 ( .A1(n9455), .A2(n9387), .ZN(n9301) );
  AOI211_X1 U10611 ( .C1(n9453), .C2(n10003), .A(n9302), .B(n9301), .ZN(n9303)
         );
  OAI21_X1 U10612 ( .B1(n9323), .B2(n9456), .A(n9303), .ZN(P1_U3274) );
  OAI21_X1 U10613 ( .B1(n9305), .B2(n9306), .A(n9304), .ZN(n9824) );
  NAND3_X1 U10614 ( .A1(n9329), .A2(n9307), .A3(n9306), .ZN(n9308) );
  NAND3_X1 U10615 ( .A1(n9309), .A2(n10019), .A3(n9308), .ZN(n9313) );
  AOI22_X1 U10616 ( .A1(n9987), .A2(n9311), .B1(n9310), .B2(n9985), .ZN(n9312)
         );
  NAND2_X1 U10617 ( .A1(n9313), .A2(n9312), .ZN(n9828) );
  AOI21_X1 U10618 ( .B1(n9337), .B2(n9318), .A(n10118), .ZN(n9315) );
  NAND2_X1 U10619 ( .A1(n9315), .A2(n9314), .ZN(n9825) );
  OAI22_X1 U10620 ( .A1(n9321), .A2(n9058), .B1(n9316), .B2(n9994), .ZN(n9317)
         );
  AOI21_X1 U10621 ( .B1(n9318), .B2(n9350), .A(n9317), .ZN(n9319) );
  OAI21_X1 U10622 ( .B1(n9825), .B2(n9353), .A(n9319), .ZN(n9320) );
  AOI21_X1 U10623 ( .B1(n9828), .B2(n9321), .A(n9320), .ZN(n9322) );
  OAI21_X1 U10624 ( .B1(n9824), .B2(n9323), .A(n9322), .ZN(P1_U3275) );
  NAND2_X1 U10625 ( .A1(n9324), .A2(n9331), .ZN(n9325) );
  NAND2_X1 U10626 ( .A1(n9326), .A2(n9325), .ZN(n9831) );
  AOI22_X1 U10627 ( .A1(n9985), .A2(n9328), .B1(n9327), .B2(n9987), .ZN(n9333)
         );
  OAI211_X1 U10628 ( .C1(n9331), .C2(n9330), .A(n9329), .B(n10019), .ZN(n9332)
         );
  OAI211_X1 U10629 ( .C1(n9831), .C2(n10015), .A(n9333), .B(n9332), .ZN(n9834)
         );
  NAND2_X1 U10630 ( .A1(n9834), .A2(n9321), .ZN(n9342) );
  OAI22_X1 U10631 ( .A1(n9321), .A2(n9335), .B1(n9334), .B2(n9994), .ZN(n9339)
         );
  OR2_X1 U10632 ( .A1(n9346), .A2(n9832), .ZN(n9336) );
  NAND2_X1 U10633 ( .A1(n9337), .A2(n9336), .ZN(n9833) );
  NOR2_X1 U10634 ( .A1(n9833), .A2(n10032), .ZN(n9338) );
  AOI211_X1 U10635 ( .C1(n9350), .C2(n9340), .A(n9339), .B(n9338), .ZN(n9341)
         );
  OAI211_X1 U10636 ( .C1(n9831), .C2(n10027), .A(n9342), .B(n9341), .ZN(
        P1_U3276) );
  XNOR2_X1 U10637 ( .A(n9344), .B(n9343), .ZN(n9842) );
  OAI21_X1 U10638 ( .B1(n9379), .B2(n9840), .A(n9469), .ZN(n9345) );
  OR2_X1 U10639 ( .A1(n9346), .A2(n9345), .ZN(n9838) );
  NAND2_X1 U10640 ( .A1(n10021), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9347) );
  OAI21_X1 U10641 ( .B1(n9994), .B2(n9348), .A(n9347), .ZN(n9349) );
  AOI21_X1 U10642 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9352) );
  OAI21_X1 U10643 ( .B1(n9838), .B2(n9353), .A(n9352), .ZN(n9362) );
  AOI21_X1 U10644 ( .B1(n9355), .B2(n9354), .A(n9989), .ZN(n9360) );
  OAI22_X1 U10645 ( .A1(n9357), .A2(n10010), .B1(n9356), .B2(n10012), .ZN(
        n9358) );
  AOI21_X1 U10646 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9839) );
  NOR2_X1 U10647 ( .A1(n9839), .A2(n9387), .ZN(n9361) );
  AOI211_X1 U10648 ( .C1(n9363), .C2(n9842), .A(n9362), .B(n9361), .ZN(n9364)
         );
  INV_X1 U10649 ( .A(n9364), .ZN(P1_U3277) );
  XNOR2_X1 U10650 ( .A(n9366), .B(n9365), .ZN(n9376) );
  OAI22_X1 U10651 ( .A1(n9368), .A2(n10010), .B1(n9367), .B2(n10012), .ZN(
        n9375) );
  NAND2_X1 U10652 ( .A1(n7430), .A2(n9369), .ZN(n9371) );
  NAND2_X1 U10653 ( .A1(n9371), .A2(n9370), .ZN(n9373) );
  XNOR2_X1 U10654 ( .A(n9373), .B(n9372), .ZN(n9461) );
  NOR2_X1 U10655 ( .A1(n9461), .A2(n10015), .ZN(n9374) );
  AOI211_X1 U10656 ( .C1(n9376), .C2(n10019), .A(n9375), .B(n9374), .ZN(n9460)
         );
  AND2_X1 U10657 ( .A1(n9377), .A2(n9457), .ZN(n9378) );
  NOR2_X1 U10658 ( .A1(n9379), .A2(n9378), .ZN(n9458) );
  INV_X1 U10659 ( .A(n9457), .ZN(n9383) );
  INV_X1 U10660 ( .A(n9380), .ZN(n9381) );
  AOI22_X1 U10661 ( .A1(n9387), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9381), .B2(
        n10020), .ZN(n9382) );
  OAI21_X1 U10662 ( .B1(n9383), .B2(n10029), .A(n9382), .ZN(n9385) );
  NOR2_X1 U10663 ( .A1(n9461), .A2(n10027), .ZN(n9384) );
  AOI211_X1 U10664 ( .C1(n9458), .C2(n10003), .A(n9385), .B(n9384), .ZN(n9386)
         );
  OAI21_X1 U10665 ( .B1(n9460), .B2(n9387), .A(n9386), .ZN(P1_U3278) );
  NAND2_X1 U10666 ( .A1(n9388), .A2(n9469), .ZN(n9389) );
  OAI211_X1 U10667 ( .C1(n9390), .C2(n10116), .A(n9389), .B(n9817), .ZN(n9475)
         );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9475), .S(n4387), .Z(
        P1_U3554) );
  AOI21_X1 U10669 ( .B1(n9822), .B2(n9392), .A(n9391), .ZN(n9393) );
  AOI22_X1 U10670 ( .A1(n9397), .A2(n9469), .B1(n9822), .B2(n9396), .ZN(n9398)
         );
  OAI211_X1 U10671 ( .C1(n9400), .C2(n9823), .A(n9399), .B(n9398), .ZN(n9477)
         );
  MUX2_X1 U10672 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9477), .S(n4387), .Z(
        P1_U3551) );
  AOI22_X1 U10673 ( .A1(n9402), .A2(n9469), .B1(n9822), .B2(n9401), .ZN(n9403)
         );
  OAI211_X1 U10674 ( .C1(n9405), .C2(n9823), .A(n9404), .B(n9403), .ZN(n9478)
         );
  MUX2_X1 U10675 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9478), .S(n4387), .Z(
        P1_U3550) );
  AOI211_X1 U10676 ( .C1(n9822), .C2(n9408), .A(n9407), .B(n9406), .ZN(n9409)
         );
  OAI21_X1 U10677 ( .B1(n9410), .B2(n9823), .A(n9409), .ZN(n9479) );
  MUX2_X1 U10678 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9479), .S(n4387), .Z(
        P1_U3549) );
  INV_X1 U10679 ( .A(n9411), .ZN(n9415) );
  AOI22_X1 U10680 ( .A1(n9413), .A2(n9469), .B1(n9822), .B2(n9412), .ZN(n9414)
         );
  OAI211_X1 U10681 ( .C1(n9416), .C2(n9823), .A(n9415), .B(n9414), .ZN(n9480)
         );
  MUX2_X1 U10682 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9480), .S(n4387), .Z(
        P1_U3548) );
  AOI211_X1 U10683 ( .C1(n9822), .C2(n9419), .A(n9418), .B(n9417), .ZN(n9420)
         );
  OAI21_X1 U10684 ( .B1(n9823), .B2(n9421), .A(n9420), .ZN(n9481) );
  MUX2_X1 U10685 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9481), .S(n4387), .Z(
        P1_U3547) );
  AOI22_X1 U10686 ( .A1(n9423), .A2(n9469), .B1(n9822), .B2(n9422), .ZN(n9424)
         );
  OAI211_X1 U10687 ( .C1(n9426), .C2(n9823), .A(n9425), .B(n9424), .ZN(n9482)
         );
  MUX2_X1 U10688 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9482), .S(n4387), .Z(
        P1_U3546) );
  AOI22_X1 U10689 ( .A1(n9428), .A2(n9469), .B1(n9822), .B2(n9427), .ZN(n9429)
         );
  OAI211_X1 U10690 ( .C1(n9431), .C2(n9823), .A(n9430), .B(n9429), .ZN(n9763)
         );
  MUX2_X1 U10691 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9763), .S(n4387), .Z(
        P1_U3545) );
  INV_X1 U10692 ( .A(n9823), .ZN(n10122) );
  NAND2_X1 U10693 ( .A1(n9432), .A2(n10122), .ZN(n9436) );
  NAND4_X1 U10694 ( .A1(n9436), .A2(n9435), .A3(n9434), .A4(n9433), .ZN(n9764)
         );
  MUX2_X1 U10695 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9764), .S(n4387), .Z(
        P1_U3544) );
  AOI211_X1 U10696 ( .C1(n9822), .C2(n9439), .A(n9438), .B(n9437), .ZN(n9440)
         );
  OAI21_X1 U10697 ( .B1(n9823), .B2(n9441), .A(n9440), .ZN(n9765) );
  MUX2_X1 U10698 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9765), .S(n4387), .Z(
        P1_U3543) );
  AOI22_X1 U10699 ( .A1(n9443), .A2(n9469), .B1(n9822), .B2(n9442), .ZN(n9444)
         );
  OAI211_X1 U10700 ( .C1(n9446), .C2(n9823), .A(n9445), .B(n9444), .ZN(n9766)
         );
  MUX2_X1 U10701 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9766), .S(n4387), .Z(
        P1_U3542) );
  AOI22_X1 U10702 ( .A1(n9448), .A2(n9469), .B1(n9822), .B2(n9447), .ZN(n9449)
         );
  OAI211_X1 U10703 ( .C1(n9823), .C2(n9451), .A(n9450), .B(n9449), .ZN(n9767)
         );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9767), .S(n4387), .Z(
        P1_U3541) );
  AOI22_X1 U10705 ( .A1(n9453), .A2(n9469), .B1(n9822), .B2(n9452), .ZN(n9454)
         );
  OAI211_X1 U10706 ( .C1(n9456), .C2(n9823), .A(n9455), .B(n9454), .ZN(n9768)
         );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9768), .S(n4387), .Z(
        P1_U3540) );
  AOI22_X1 U10708 ( .A1(n9458), .A2(n9469), .B1(n9822), .B2(n9457), .ZN(n9459)
         );
  OAI211_X1 U10709 ( .C1(n9473), .C2(n9461), .A(n9460), .B(n9459), .ZN(n9769)
         );
  MUX2_X1 U10710 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9769), .S(n4387), .Z(
        P1_U3536) );
  AOI211_X1 U10711 ( .C1(n9822), .C2(n9464), .A(n9463), .B(n9462), .ZN(n9465)
         );
  OAI21_X1 U10712 ( .B1(n9823), .B2(n9466), .A(n9465), .ZN(n9770) );
  MUX2_X1 U10713 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9770), .S(n4387), .Z(
        P1_U3535) );
  INV_X1 U10714 ( .A(n9467), .ZN(n9474) );
  AOI22_X1 U10715 ( .A1(n9470), .A2(n9469), .B1(n9822), .B2(n9468), .ZN(n9471)
         );
  OAI211_X1 U10716 ( .C1(n9474), .C2(n9473), .A(n9472), .B(n9471), .ZN(n9771)
         );
  MUX2_X1 U10717 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9771), .S(n4387), .Z(
        P1_U3534) );
  MUX2_X1 U10718 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9475), .S(n10126), .Z(
        P1_U3522) );
  MUX2_X1 U10719 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9476), .S(n10126), .Z(
        P1_U3520) );
  MUX2_X1 U10720 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9477), .S(n10126), .Z(
        P1_U3519) );
  MUX2_X1 U10721 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9478), .S(n10126), .Z(
        P1_U3518) );
  MUX2_X1 U10722 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9479), .S(n10126), .Z(
        P1_U3517) );
  MUX2_X1 U10723 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9480), .S(n10126), .Z(
        P1_U3516) );
  MUX2_X1 U10724 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9481), .S(n10126), .Z(
        P1_U3515) );
  MUX2_X1 U10725 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9482), .S(n10126), .Z(
        n9762) );
  NOR2_X1 U10726 ( .A1(keyinput62), .A2(keyinput92), .ZN(n9483) );
  NAND3_X1 U10727 ( .A1(keyinput59), .A2(keyinput89), .A3(n9483), .ZN(n9541)
         );
  INV_X1 U10728 ( .A(keyinput91), .ZN(n9484) );
  NAND4_X1 U10729 ( .A1(keyinput85), .A2(keyinput49), .A3(keyinput118), .A4(
        n9484), .ZN(n9540) );
  NAND4_X1 U10730 ( .A1(keyinput11), .A2(keyinput77), .A3(keyinput86), .A4(
        keyinput115), .ZN(n9485) );
  NOR3_X1 U10731 ( .A1(keyinput75), .A2(keyinput16), .A3(n9485), .ZN(n9493) );
  NOR2_X1 U10732 ( .A1(keyinput69), .A2(keyinput108), .ZN(n9486) );
  NAND3_X1 U10733 ( .A1(keyinput46), .A2(keyinput51), .A3(n9486), .ZN(n9490)
         );
  NAND4_X1 U10734 ( .A1(keyinput34), .A2(keyinput68), .A3(keyinput37), .A4(
        keyinput106), .ZN(n9489) );
  NAND4_X1 U10735 ( .A1(keyinput41), .A2(keyinput17), .A3(keyinput13), .A4(
        keyinput24), .ZN(n9488) );
  OR4_X1 U10736 ( .A1(keyinput123), .A2(keyinput102), .A3(keyinput73), .A4(
        keyinput90), .ZN(n9487) );
  NOR4_X1 U10737 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n9492)
         );
  INV_X1 U10738 ( .A(keyinput8), .ZN(n9491) );
  NAND4_X1 U10739 ( .A1(keyinput98), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(
        n9539) );
  NOR4_X1 U10740 ( .A1(keyinput28), .A2(keyinput26), .A3(keyinput113), .A4(
        keyinput65), .ZN(n9494) );
  NAND4_X1 U10741 ( .A1(keyinput116), .A2(keyinput5), .A3(keyinput10), .A4(
        n9494), .ZN(n9505) );
  NAND4_X1 U10742 ( .A1(keyinput57), .A2(keyinput9), .A3(keyinput122), .A4(
        keyinput38), .ZN(n9504) );
  NOR2_X1 U10743 ( .A1(keyinput67), .A2(keyinput80), .ZN(n9495) );
  NAND3_X1 U10744 ( .A1(keyinput111), .A2(keyinput25), .A3(n9495), .ZN(n9503)
         );
  AND4_X1 U10745 ( .A1(keyinput101), .A2(keyinput72), .A3(keyinput21), .A4(
        keyinput125), .ZN(n9501) );
  NOR4_X1 U10746 ( .A1(keyinput2), .A2(keyinput103), .A3(keyinput35), .A4(
        keyinput61), .ZN(n9500) );
  NAND2_X1 U10747 ( .A1(keyinput66), .A2(keyinput33), .ZN(n9496) );
  NOR3_X1 U10748 ( .A1(keyinput4), .A2(keyinput45), .A3(n9496), .ZN(n9499) );
  INV_X1 U10749 ( .A(keyinput15), .ZN(n9497) );
  NOR4_X1 U10750 ( .A1(keyinput121), .A2(keyinput96), .A3(keyinput124), .A4(
        n9497), .ZN(n9498) );
  NAND4_X1 U10751 ( .A1(n9501), .A2(n9500), .A3(n9499), .A4(n9498), .ZN(n9502)
         );
  NOR4_X1 U10752 ( .A1(n9505), .A2(n9504), .A3(n9503), .A4(n9502), .ZN(n9537)
         );
  NOR2_X1 U10753 ( .A1(keyinput107), .A2(keyinput42), .ZN(n9506) );
  NAND3_X1 U10754 ( .A1(keyinput71), .A2(keyinput105), .A3(n9506), .ZN(n9518)
         );
  NAND4_X1 U10755 ( .A1(keyinput95), .A2(keyinput7), .A3(keyinput36), .A4(
        keyinput94), .ZN(n9517) );
  NOR2_X1 U10756 ( .A1(keyinput39), .A2(keyinput22), .ZN(n9508) );
  NOR4_X1 U10757 ( .A1(keyinput82), .A2(keyinput14), .A3(keyinput100), .A4(
        keyinput40), .ZN(n9507) );
  NAND4_X1 U10758 ( .A1(n9508), .A2(keyinput84), .A3(keyinput18), .A4(n9507), 
        .ZN(n9516) );
  INV_X1 U10759 ( .A(keyinput55), .ZN(n9509) );
  NOR4_X1 U10760 ( .A1(keyinput97), .A2(keyinput76), .A3(keyinput6), .A4(n9509), .ZN(n9514) );
  NOR4_X1 U10761 ( .A1(keyinput79), .A2(keyinput127), .A3(keyinput117), .A4(
        keyinput43), .ZN(n9513) );
  NAND3_X1 U10762 ( .A1(keyinput114), .A2(keyinput1), .A3(keyinput53), .ZN(
        n9510) );
  NOR2_X1 U10763 ( .A1(keyinput70), .A2(n9510), .ZN(n9512) );
  INV_X1 U10764 ( .A(keyinput47), .ZN(n9594) );
  NOR4_X1 U10765 ( .A1(keyinput78), .A2(keyinput20), .A3(keyinput54), .A4(
        n9594), .ZN(n9511) );
  NAND4_X1 U10766 ( .A1(n9514), .A2(n9513), .A3(n9512), .A4(n9511), .ZN(n9515)
         );
  NOR4_X1 U10767 ( .A1(n9518), .A2(n9517), .A3(n9516), .A4(n9515), .ZN(n9536)
         );
  INV_X1 U10768 ( .A(keyinput87), .ZN(n9519) );
  NAND4_X1 U10769 ( .A1(keyinput81), .A2(keyinput19), .A3(keyinput27), .A4(
        n9519), .ZN(n9526) );
  NOR2_X1 U10770 ( .A1(keyinput109), .A2(keyinput64), .ZN(n9520) );
  NAND3_X1 U10771 ( .A1(keyinput30), .A2(keyinput88), .A3(n9520), .ZN(n9525)
         );
  INV_X1 U10772 ( .A(keyinput104), .ZN(n9521) );
  NAND4_X1 U10773 ( .A1(keyinput120), .A2(keyinput83), .A3(keyinput0), .A4(
        n9521), .ZN(n9524) );
  NOR2_X1 U10774 ( .A1(keyinput74), .A2(keyinput3), .ZN(n9522) );
  NAND3_X1 U10775 ( .A1(keyinput23), .A2(keyinput12), .A3(n9522), .ZN(n9523)
         );
  NOR4_X1 U10776 ( .A1(n9526), .A2(n9525), .A3(n9524), .A4(n9523), .ZN(n9535)
         );
  NOR4_X1 U10777 ( .A1(keyinput48), .A2(keyinput119), .A3(keyinput110), .A4(
        keyinput112), .ZN(n9533) );
  NAND2_X1 U10778 ( .A1(keyinput93), .A2(keyinput60), .ZN(n9527) );
  NOR3_X1 U10779 ( .A1(keyinput56), .A2(keyinput29), .A3(n9527), .ZN(n9532) );
  INV_X1 U10780 ( .A(keyinput126), .ZN(n9528) );
  NOR4_X1 U10781 ( .A1(keyinput31), .A2(keyinput99), .A3(keyinput44), .A4(
        n9528), .ZN(n9531) );
  NAND2_X1 U10782 ( .A1(keyinput50), .A2(keyinput52), .ZN(n9529) );
  NOR3_X1 U10783 ( .A1(keyinput58), .A2(keyinput32), .A3(n9529), .ZN(n9530) );
  AND4_X1 U10784 ( .A1(n9533), .A2(n9532), .A3(n9531), .A4(n9530), .ZN(n9534)
         );
  NAND4_X1 U10785 ( .A1(n9537), .A2(n9536), .A3(n9535), .A4(n9534), .ZN(n9538)
         );
  NOR4_X1 U10786 ( .A1(n9541), .A2(n9540), .A3(n9539), .A4(n9538), .ZN(n9542)
         );
  OAI21_X1 U10787 ( .B1(keyinput63), .B2(n9542), .A(n6367), .ZN(n9760) );
  INV_X1 U10788 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U10789 ( .A1(n10226), .A2(keyinput65), .B1(n9170), .B2(keyinput2), 
        .ZN(n9543) );
  OAI221_X1 U10790 ( .B1(n10226), .B2(keyinput65), .C1(n9170), .C2(keyinput2), 
        .A(n9543), .ZN(n9618) );
  AOI22_X1 U10791 ( .A1(n9545), .A2(keyinput26), .B1(keyinput113), .B2(n5372), 
        .ZN(n9544) );
  OAI221_X1 U10792 ( .B1(n9545), .B2(keyinput26), .C1(n5372), .C2(keyinput113), 
        .A(n9544), .ZN(n9617) );
  INV_X1 U10793 ( .A(keyinput5), .ZN(n9551) );
  INV_X1 U10794 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9548) );
  AOI22_X1 U10795 ( .A1(n9548), .A2(keyinput10), .B1(n9547), .B2(keyinput28), 
        .ZN(n9546) );
  OAI221_X1 U10796 ( .B1(n9548), .B2(keyinput10), .C1(n9547), .C2(keyinput28), 
        .A(n9546), .ZN(n9549) );
  AOI221_X1 U10797 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n9551), .C1(n9550), .C2(
        keyinput5), .A(n9549), .ZN(n9565) );
  INV_X1 U10798 ( .A(keyinput101), .ZN(n9553) );
  AOI22_X1 U10799 ( .A1(n9554), .A2(keyinput103), .B1(P1_ADDR_REG_13__SCAN_IN), 
        .B2(n9553), .ZN(n9552) );
  OAI221_X1 U10800 ( .B1(n9554), .B2(keyinput103), .C1(n9553), .C2(
        P1_ADDR_REG_13__SCAN_IN), .A(n9552), .ZN(n9563) );
  INV_X1 U10801 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U10802 ( .A1(n5102), .A2(keyinput61), .B1(keyinput21), .B2(n10231), 
        .ZN(n9555) );
  OAI221_X1 U10803 ( .B1(n5102), .B2(keyinput61), .C1(n10231), .C2(keyinput21), 
        .A(n9555), .ZN(n9562) );
  INV_X1 U10804 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10108) );
  INV_X1 U10805 ( .A(keyinput72), .ZN(n9557) );
  AOI22_X1 U10806 ( .A1(n10108), .A2(keyinput35), .B1(P1_ADDR_REG_1__SCAN_IN), 
        .B2(n9557), .ZN(n9556) );
  OAI221_X1 U10807 ( .B1(n10108), .B2(keyinput35), .C1(n9557), .C2(
        P1_ADDR_REG_1__SCAN_IN), .A(n9556), .ZN(n9561) );
  XOR2_X1 U10808 ( .A(n5950), .B(keyinput125), .Z(n9559) );
  XNOR2_X1 U10809 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput121), .ZN(n9558) );
  NAND2_X1 U10810 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  NOR4_X1 U10811 ( .A1(n9563), .A2(n9562), .A3(n9561), .A4(n9560), .ZN(n9564)
         );
  OAI211_X1 U10812 ( .C1(keyinput63), .C2(n6367), .A(n9565), .B(n9564), .ZN(
        n9616) );
  AOI22_X1 U10813 ( .A1(n6959), .A2(keyinput14), .B1(n9567), .B2(keyinput100), 
        .ZN(n9566) );
  OAI221_X1 U10814 ( .B1(n6959), .B2(keyinput14), .C1(n9567), .C2(keyinput100), 
        .A(n9566), .ZN(n9577) );
  AOI22_X1 U10815 ( .A1(n9569), .A2(keyinput40), .B1(n6321), .B2(keyinput79), 
        .ZN(n9568) );
  OAI221_X1 U10816 ( .B1(n9569), .B2(keyinput40), .C1(n6321), .C2(keyinput79), 
        .A(n9568), .ZN(n9576) );
  AOI22_X1 U10817 ( .A1(n9066), .A2(keyinput18), .B1(keyinput82), .B2(n9571), 
        .ZN(n9570) );
  OAI221_X1 U10818 ( .B1(n9066), .B2(keyinput18), .C1(n9571), .C2(keyinput82), 
        .A(n9570), .ZN(n9575) );
  XNOR2_X1 U10819 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput22), .ZN(n9573) );
  XNOR2_X1 U10820 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput84), .ZN(n9572) );
  NAND2_X1 U10821 ( .A1(n9573), .A2(n9572), .ZN(n9574) );
  NOR4_X1 U10822 ( .A1(n9577), .A2(n9576), .A3(n9575), .A4(n9574), .ZN(n9614)
         );
  INV_X1 U10823 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10228) );
  INV_X1 U10824 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U10825 ( .A1(n10228), .A2(keyinput7), .B1(n10039), .B2(keyinput71), 
        .ZN(n9578) );
  OAI221_X1 U10826 ( .B1(n10228), .B2(keyinput7), .C1(n10039), .C2(keyinput71), 
        .A(n9578), .ZN(n9590) );
  AOI22_X1 U10827 ( .A1(n9581), .A2(keyinput94), .B1(n9580), .B2(keyinput105), 
        .ZN(n9579) );
  OAI221_X1 U10828 ( .B1(n9581), .B2(keyinput94), .C1(n9580), .C2(keyinput105), 
        .A(n9579), .ZN(n9589) );
  AOI22_X1 U10829 ( .A1(n9584), .A2(keyinput42), .B1(n9583), .B2(keyinput39), 
        .ZN(n9582) );
  OAI221_X1 U10830 ( .B1(n9584), .B2(keyinput42), .C1(n9583), .C2(keyinput39), 
        .A(n9582), .ZN(n9588) );
  XNOR2_X1 U10831 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput107), .ZN(n9586)
         );
  XNOR2_X1 U10832 ( .A(SI_8_), .B(keyinput36), .ZN(n9585) );
  NAND2_X1 U10833 ( .A1(n9586), .A2(n9585), .ZN(n9587) );
  NOR4_X1 U10834 ( .A1(n9590), .A2(n9589), .A3(n9588), .A4(n9587), .ZN(n9613)
         );
  INV_X1 U10835 ( .A(keyinput70), .ZN(n9592) );
  AOI22_X1 U10836 ( .A1(n4666), .A2(keyinput1), .B1(P1_ADDR_REG_7__SCAN_IN), 
        .B2(n9592), .ZN(n9591) );
  OAI221_X1 U10837 ( .B1(n4666), .B2(keyinput1), .C1(n9592), .C2(
        P1_ADDR_REG_7__SCAN_IN), .A(n9591), .ZN(n9602) );
  INV_X1 U10838 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U10839 ( .A1(n10229), .A2(keyinput20), .B1(P1_ADDR_REG_8__SCAN_IN), 
        .B2(n9594), .ZN(n9593) );
  OAI221_X1 U10840 ( .B1(n10229), .B2(keyinput20), .C1(n9594), .C2(
        P1_ADDR_REG_8__SCAN_IN), .A(n9593), .ZN(n9601) );
  INV_X1 U10841 ( .A(keyinput53), .ZN(n9596) );
  AOI22_X1 U10842 ( .A1(n6099), .A2(keyinput54), .B1(P2_WR_REG_SCAN_IN), .B2(
        n9596), .ZN(n9595) );
  OAI221_X1 U10843 ( .B1(n6099), .B2(keyinput54), .C1(n9596), .C2(
        P2_WR_REG_SCAN_IN), .A(n9595), .ZN(n9600) );
  XNOR2_X1 U10844 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput114), .ZN(n9598) );
  XNOR2_X1 U10845 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput49), .ZN(n9597) );
  NAND2_X1 U10846 ( .A1(n9598), .A2(n9597), .ZN(n9599) );
  NOR4_X1 U10847 ( .A1(n9602), .A2(n9601), .A3(n9600), .A4(n9599), .ZN(n9612)
         );
  INV_X1 U10848 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n10038) );
  AOI22_X1 U10849 ( .A1(n6479), .A2(keyinput43), .B1(n10038), .B2(keyinput55), 
        .ZN(n9603) );
  OAI221_X1 U10850 ( .B1(n6479), .B2(keyinput43), .C1(n10038), .C2(keyinput55), 
        .A(n9603), .ZN(n9610) );
  AOI22_X1 U10851 ( .A1(n8756), .A2(keyinput127), .B1(n5071), .B2(keyinput117), 
        .ZN(n9604) );
  OAI221_X1 U10852 ( .B1(n8756), .B2(keyinput127), .C1(n5071), .C2(keyinput117), .A(n9604), .ZN(n9609) );
  AOI22_X1 U10853 ( .A1(n5394), .A2(keyinput6), .B1(n6243), .B2(keyinput78), 
        .ZN(n9605) );
  OAI221_X1 U10854 ( .B1(n5394), .B2(keyinput6), .C1(n6243), .C2(keyinput78), 
        .A(n9605), .ZN(n9608) );
  AOI22_X1 U10855 ( .A1(n5198), .A2(keyinput76), .B1(keyinput97), .B2(n5809), 
        .ZN(n9606) );
  OAI221_X1 U10856 ( .B1(n5198), .B2(keyinput76), .C1(n5809), .C2(keyinput97), 
        .A(n9606), .ZN(n9607) );
  NOR4_X1 U10857 ( .A1(n9610), .A2(n9609), .A3(n9608), .A4(n9607), .ZN(n9611)
         );
  NAND4_X1 U10858 ( .A1(n9614), .A2(n9613), .A3(n9612), .A4(n9611), .ZN(n9615)
         );
  NOR4_X1 U10859 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n9759)
         );
  AOI22_X1 U10860 ( .A1(n5536), .A2(keyinput68), .B1(keyinput37), .B2(n5792), 
        .ZN(n9619) );
  OAI221_X1 U10861 ( .B1(n5536), .B2(keyinput68), .C1(n5792), .C2(keyinput37), 
        .A(n9619), .ZN(n9632) );
  AOI22_X1 U10862 ( .A1(n9622), .A2(keyinput106), .B1(n9621), .B2(keyinput69), 
        .ZN(n9620) );
  OAI221_X1 U10863 ( .B1(n9622), .B2(keyinput106), .C1(n9621), .C2(keyinput69), 
        .A(n9620), .ZN(n9631) );
  INV_X1 U10864 ( .A(keyinput46), .ZN(n9625) );
  INV_X1 U10865 ( .A(keyinput108), .ZN(n9624) );
  AOI22_X1 U10866 ( .A1(n9625), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(
        P1_ADDR_REG_0__SCAN_IN), .B2(n9624), .ZN(n9623) );
  OAI221_X1 U10867 ( .B1(n9625), .B2(P1_ADDR_REG_10__SCAN_IN), .C1(n9624), 
        .C2(P1_ADDR_REG_0__SCAN_IN), .A(n9623), .ZN(n9630) );
  INV_X1 U10868 ( .A(keyinput123), .ZN(n9627) );
  AOI22_X1 U10869 ( .A1(n9628), .A2(keyinput51), .B1(P2_ADDR_REG_17__SCAN_IN), 
        .B2(n9627), .ZN(n9626) );
  OAI221_X1 U10870 ( .B1(n9628), .B2(keyinput51), .C1(n9627), .C2(
        P2_ADDR_REG_17__SCAN_IN), .A(n9626), .ZN(n9629) );
  NOR4_X1 U10871 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n9645)
         );
  AOI22_X1 U10872 ( .A1(n5129), .A2(keyinput124), .B1(keyinput33), .B2(n6403), 
        .ZN(n9633) );
  OAI221_X1 U10873 ( .B1(n5129), .B2(keyinput124), .C1(n6403), .C2(keyinput33), 
        .A(n9633), .ZN(n9643) );
  INV_X1 U10874 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U10875 ( .A1(n9635), .A2(keyinput96), .B1(keyinput15), .B2(n10149), 
        .ZN(n9634) );
  OAI221_X1 U10876 ( .B1(n9635), .B2(keyinput96), .C1(n10149), .C2(keyinput15), 
        .A(n9634), .ZN(n9642) );
  INV_X1 U10877 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n9637) );
  AOI22_X1 U10878 ( .A1(n9637), .A2(keyinput45), .B1(n5869), .B2(keyinput111), 
        .ZN(n9636) );
  OAI221_X1 U10879 ( .B1(n9637), .B2(keyinput45), .C1(n5869), .C2(keyinput111), 
        .A(n9636), .ZN(n9641) );
  INV_X1 U10880 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10063) );
  INV_X1 U10881 ( .A(keyinput66), .ZN(n9639) );
  AOI22_X1 U10882 ( .A1(n10063), .A2(keyinput4), .B1(P2_ADDR_REG_1__SCAN_IN), 
        .B2(n9639), .ZN(n9638) );
  OAI221_X1 U10883 ( .B1(n10063), .B2(keyinput4), .C1(n9639), .C2(
        P2_ADDR_REG_1__SCAN_IN), .A(n9638), .ZN(n9640) );
  NOR4_X1 U10884 ( .A1(n9643), .A2(n9642), .A3(n9641), .A4(n9640), .ZN(n9644)
         );
  NAND2_X1 U10885 ( .A1(n9645), .A2(n9644), .ZN(n9757) );
  INV_X1 U10886 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9648) );
  AOI22_X1 U10887 ( .A1(n9648), .A2(keyinput85), .B1(keyinput91), .B2(n9647), 
        .ZN(n9646) );
  OAI221_X1 U10888 ( .B1(n9648), .B2(keyinput85), .C1(n9647), .C2(keyinput91), 
        .A(n9646), .ZN(n9652) );
  INV_X1 U10889 ( .A(SI_4_), .ZN(n9650) );
  AOI22_X1 U10890 ( .A1(n9650), .A2(keyinput29), .B1(keyinput56), .B2(n5728), 
        .ZN(n9649) );
  OAI221_X1 U10891 ( .B1(n9650), .B2(keyinput29), .C1(n5728), .C2(keyinput56), 
        .A(n9649), .ZN(n9651) );
  NOR2_X1 U10892 ( .A1(n9652), .A2(n9651), .ZN(n9674) );
  INV_X1 U10893 ( .A(SI_11_), .ZN(n9654) );
  INV_X1 U10894 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n10051) );
  AOI22_X1 U10895 ( .A1(n9654), .A2(keyinput115), .B1(n10051), .B2(keyinput60), 
        .ZN(n9653) );
  OAI221_X1 U10896 ( .B1(n9654), .B2(keyinput115), .C1(n10051), .C2(keyinput60), .A(n9653), .ZN(n9657) );
  INV_X1 U10897 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10227) );
  INV_X1 U10898 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10064) );
  AOI22_X1 U10899 ( .A1(n10227), .A2(keyinput62), .B1(n10064), .B2(keyinput89), 
        .ZN(n9655) );
  OAI221_X1 U10900 ( .B1(n10227), .B2(keyinput62), .C1(n10064), .C2(keyinput89), .A(n9655), .ZN(n9656) );
  NOR2_X1 U10901 ( .A1(n9657), .A2(n9656), .ZN(n9673) );
  AOI22_X1 U10902 ( .A1(n5922), .A2(keyinput118), .B1(n9659), .B2(keyinput59), 
        .ZN(n9658) );
  OAI221_X1 U10903 ( .B1(n5922), .B2(keyinput118), .C1(n9659), .C2(keyinput59), 
        .A(n9658), .ZN(n9665) );
  XNOR2_X1 U10904 ( .A(P2_REG1_REG_28__SCAN_IN), .B(keyinput110), .ZN(n9663)
         );
  XNOR2_X1 U10905 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput112), .ZN(n9662) );
  XNOR2_X1 U10906 ( .A(keyinput16), .B(P1_REG3_REG_1__SCAN_IN), .ZN(n9661) );
  XNOR2_X1 U10907 ( .A(keyinput73), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n9660) );
  NAND4_X1 U10908 ( .A1(n9663), .A2(n9662), .A3(n9661), .A4(n9660), .ZN(n9664)
         );
  NOR2_X1 U10909 ( .A1(n9665), .A2(n9664), .ZN(n9672) );
  INV_X1 U10910 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U10911 ( .A1(n10232), .A2(keyinput93), .B1(n5075), .B2(keyinput48), 
        .ZN(n9666) );
  OAI221_X1 U10912 ( .B1(n10232), .B2(keyinput93), .C1(n5075), .C2(keyinput48), 
        .A(n9666), .ZN(n9670) );
  AOI22_X1 U10913 ( .A1(n6389), .A2(keyinput77), .B1(n9668), .B2(keyinput75), 
        .ZN(n9667) );
  OAI221_X1 U10914 ( .B1(n6389), .B2(keyinput77), .C1(n9668), .C2(keyinput75), 
        .A(n9667), .ZN(n9669) );
  NOR2_X1 U10915 ( .A1(n9670), .A2(n9669), .ZN(n9671) );
  NAND4_X1 U10916 ( .A1(n9674), .A2(n9673), .A3(n9672), .A4(n9671), .ZN(n9702)
         );
  AOI22_X1 U10917 ( .A1(n6644), .A2(keyinput8), .B1(keyinput11), .B2(n5200), 
        .ZN(n9675) );
  OAI221_X1 U10918 ( .B1(n6644), .B2(keyinput8), .C1(n5200), .C2(keyinput11), 
        .A(n9675), .ZN(n9676) );
  INV_X1 U10919 ( .A(n9676), .ZN(n9700) );
  AOI22_X1 U10920 ( .A1(n9678), .A2(keyinput24), .B1(keyinput98), .B2(n5196), 
        .ZN(n9677) );
  OAI221_X1 U10921 ( .B1(n9678), .B2(keyinput24), .C1(n5196), .C2(keyinput98), 
        .A(n9677), .ZN(n9679) );
  INV_X1 U10922 ( .A(n9679), .ZN(n9699) );
  INV_X1 U10923 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10052) );
  AOI22_X1 U10924 ( .A1(n10052), .A2(keyinput17), .B1(keyinput13), .B2(n9681), 
        .ZN(n9680) );
  OAI221_X1 U10925 ( .B1(n10052), .B2(keyinput17), .C1(n9681), .C2(keyinput13), 
        .A(n9680), .ZN(n9686) );
  AOI22_X1 U10926 ( .A1(n9684), .A2(keyinput90), .B1(n9683), .B2(keyinput41), 
        .ZN(n9682) );
  OAI221_X1 U10927 ( .B1(n9684), .B2(keyinput90), .C1(n9683), .C2(keyinput41), 
        .A(n9682), .ZN(n9685) );
  NOR2_X1 U10928 ( .A1(n9686), .A2(n9685), .ZN(n9698) );
  XNOR2_X1 U10929 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput92), .ZN(n9690) );
  XNOR2_X1 U10930 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput102), .ZN(n9689) );
  XNOR2_X1 U10931 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput34), .ZN(n9688) );
  XNOR2_X1 U10932 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput104), .ZN(n9687) );
  NAND4_X1 U10933 ( .A1(n9690), .A2(n9689), .A3(n9688), .A4(n9687), .ZN(n9696)
         );
  XNOR2_X1 U10934 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput86), .ZN(n9694) );
  XNOR2_X1 U10935 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput119), .ZN(n9693) );
  XNOR2_X1 U10936 ( .A(P2_IR_REG_27__SCAN_IN), .B(keyinput120), .ZN(n9692) );
  XNOR2_X1 U10937 ( .A(P1_REG1_REG_31__SCAN_IN), .B(keyinput30), .ZN(n9691) );
  NAND4_X1 U10938 ( .A1(n9694), .A2(n9693), .A3(n9692), .A4(n9691), .ZN(n9695)
         );
  NOR2_X1 U10939 ( .A1(n9696), .A2(n9695), .ZN(n9697) );
  NAND4_X1 U10940 ( .A1(n9700), .A2(n9699), .A3(n9698), .A4(n9697), .ZN(n9701)
         );
  NOR2_X1 U10941 ( .A1(n9702), .A2(n9701), .ZN(n9713) );
  INV_X1 U10942 ( .A(keyinput12), .ZN(n9704) );
  OAI22_X1 U10943 ( .A1(n9096), .A2(keyinput83), .B1(n9704), .B2(SI_31_), .ZN(
        n9703) );
  AOI221_X1 U10944 ( .B1(n9096), .B2(keyinput83), .C1(SI_31_), .C2(n9704), .A(
        n9703), .ZN(n9712) );
  INV_X1 U10945 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9707) );
  INV_X1 U10946 ( .A(keyinput74), .ZN(n9706) );
  OAI22_X1 U10947 ( .A1(keyinput3), .A2(n9707), .B1(n9706), .B2(
        P1_ADDR_REG_15__SCAN_IN), .ZN(n9705) );
  AOI221_X1 U10948 ( .B1(n9707), .B2(keyinput3), .C1(n9706), .C2(
        P1_ADDR_REG_15__SCAN_IN), .A(n9705), .ZN(n9711) );
  OAI22_X1 U10949 ( .A1(n9709), .A2(keyinput0), .B1(n5925), .B2(keyinput58), 
        .ZN(n9708) );
  AOI221_X1 U10950 ( .B1(n9709), .B2(keyinput0), .C1(keyinput58), .C2(n5925), 
        .A(n9708), .ZN(n9710) );
  AND4_X1 U10951 ( .A1(n9713), .A2(n9712), .A3(n9711), .A4(n9710), .ZN(n9755)
         );
  AOI22_X1 U10952 ( .A1(n9715), .A2(keyinput109), .B1(keyinput88), .B2(n6406), 
        .ZN(n9714) );
  OAI221_X1 U10953 ( .B1(n9715), .B2(keyinput109), .C1(n6406), .C2(keyinput88), 
        .A(n9714), .ZN(n9726) );
  AOI22_X1 U10954 ( .A1(n5304), .A2(keyinput64), .B1(n9717), .B2(keyinput81), 
        .ZN(n9716) );
  OAI221_X1 U10955 ( .B1(n5304), .B2(keyinput64), .C1(n9717), .C2(keyinput81), 
        .A(n9716), .ZN(n9725) );
  AOI22_X1 U10956 ( .A1(n6600), .A2(keyinput87), .B1(keyinput19), .B2(n9719), 
        .ZN(n9718) );
  OAI221_X1 U10957 ( .B1(n6600), .B2(keyinput87), .C1(n9719), .C2(keyinput19), 
        .A(n9718), .ZN(n9724) );
  AOI22_X1 U10958 ( .A1(n9722), .A2(keyinput27), .B1(n9721), .B2(keyinput23), 
        .ZN(n9720) );
  OAI221_X1 U10959 ( .B1(n9722), .B2(keyinput27), .C1(n9721), .C2(keyinput23), 
        .A(n9720), .ZN(n9723) );
  NOR4_X1 U10960 ( .A1(n9726), .A2(n9725), .A3(n9724), .A4(n9723), .ZN(n9754)
         );
  AOI22_X1 U10961 ( .A1(n9728), .A2(keyinput80), .B1(n4509), .B2(keyinput57), 
        .ZN(n9727) );
  OAI221_X1 U10962 ( .B1(n9728), .B2(keyinput80), .C1(n4509), .C2(keyinput57), 
        .A(n9727), .ZN(n9739) );
  AOI22_X1 U10963 ( .A1(n9731), .A2(keyinput67), .B1(keyinput25), .B2(n9730), 
        .ZN(n9729) );
  OAI221_X1 U10964 ( .B1(n9731), .B2(keyinput67), .C1(n9730), .C2(keyinput25), 
        .A(n9729), .ZN(n9738) );
  AOI22_X1 U10965 ( .A1(n9733), .A2(keyinput38), .B1(keyinput95), .B2(n9335), 
        .ZN(n9732) );
  OAI221_X1 U10966 ( .B1(n9733), .B2(keyinput38), .C1(n9335), .C2(keyinput95), 
        .A(n9732), .ZN(n9737) );
  AOI22_X1 U10967 ( .A1(n9735), .A2(keyinput9), .B1(n10128), .B2(keyinput122), 
        .ZN(n9734) );
  OAI221_X1 U10968 ( .B1(n9735), .B2(keyinput9), .C1(n10128), .C2(keyinput122), 
        .A(n9734), .ZN(n9736) );
  NOR4_X1 U10969 ( .A1(n9739), .A2(n9738), .A3(n9737), .A4(n9736), .ZN(n9753)
         );
  INV_X1 U10970 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U10971 ( .A1(n10280), .A2(keyinput52), .B1(keyinput50), .B2(n6427), 
        .ZN(n9740) );
  OAI221_X1 U10972 ( .B1(n10280), .B2(keyinput52), .C1(n6427), .C2(keyinput50), 
        .A(n9740), .ZN(n9751) );
  INV_X1 U10973 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9843) );
  AOI22_X1 U10974 ( .A1(n9843), .A2(keyinput32), .B1(n9742), .B2(keyinput31), 
        .ZN(n9741) );
  OAI221_X1 U10975 ( .B1(n9843), .B2(keyinput32), .C1(n9742), .C2(keyinput31), 
        .A(n9741), .ZN(n9750) );
  INV_X1 U10976 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U10977 ( .A1(n9744), .A2(keyinput99), .B1(keyinput126), .B2(n10230), 
        .ZN(n9743) );
  OAI221_X1 U10978 ( .B1(n9744), .B2(keyinput99), .C1(n10230), .C2(keyinput126), .A(n9743), .ZN(n9749) );
  AOI22_X1 U10979 ( .A1(n9747), .A2(keyinput116), .B1(keyinput44), .B2(n9746), 
        .ZN(n9745) );
  OAI221_X1 U10980 ( .B1(n9747), .B2(keyinput116), .C1(n9746), .C2(keyinput44), 
        .A(n9745), .ZN(n9748) );
  NOR4_X1 U10981 ( .A1(n9751), .A2(n9750), .A3(n9749), .A4(n9748), .ZN(n9752)
         );
  NAND4_X1 U10982 ( .A1(n9755), .A2(n9754), .A3(n9753), .A4(n9752), .ZN(n9756)
         );
  NOR2_X1 U10983 ( .A1(n9757), .A2(n9756), .ZN(n9758) );
  NAND3_X1 U10984 ( .A1(n9760), .A2(n9759), .A3(n9758), .ZN(n9761) );
  XNOR2_X1 U10985 ( .A(n9762), .B(n9761), .ZN(P1_U3514) );
  MUX2_X1 U10986 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9763), .S(n10126), .Z(
        P1_U3513) );
  MUX2_X1 U10987 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9764), .S(n10126), .Z(
        P1_U3512) );
  MUX2_X1 U10988 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9765), .S(n10126), .Z(
        P1_U3511) );
  MUX2_X1 U10989 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9766), .S(n10126), .Z(
        P1_U3510) );
  MUX2_X1 U10990 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9767), .S(n10126), .Z(
        P1_U3508) );
  MUX2_X1 U10991 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9768), .S(n10126), .Z(
        P1_U3505) );
  MUX2_X1 U10992 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9769), .S(n10126), .Z(
        P1_U3493) );
  MUX2_X1 U10993 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9770), .S(n10126), .Z(
        P1_U3490) );
  MUX2_X1 U10994 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9771), .S(n10126), .Z(
        P1_U3487) );
  NOR4_X1 U10995 ( .A1(n9772), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3084), .A4(
        n5280), .ZN(n9773) );
  AOI21_X1 U10996 ( .B1(n9774), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9773), .ZN(
        n9775) );
  OAI21_X1 U10997 ( .B1(n9776), .B2(n4389), .A(n9775), .ZN(P1_U3322) );
  NAND2_X1 U10998 ( .A1(n9778), .A2(n9777), .ZN(n9780) );
  OAI211_X1 U10999 ( .C1(n9782), .C2(n9781), .A(n9780), .B(n9779), .ZN(
        P1_U3325) );
  MUX2_X1 U11000 ( .A(n9783), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI21_X1 U11001 ( .B1(n9786), .B2(n9785), .A(n9784), .ZN(n9790) );
  OAI22_X1 U11002 ( .A1(n9788), .A2(n9787), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10149), .ZN(n9789) );
  AOI21_X1 U11003 ( .B1(n10168), .B2(n9790), .A(n9789), .ZN(n9793) );
  NAND2_X1 U11004 ( .A1(n10166), .A2(n9791), .ZN(n9792) );
  AND2_X1 U11005 ( .A1(n9793), .A2(n9792), .ZN(n9798) );
  AND2_X1 U11006 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9795) );
  OAI211_X1 U11007 ( .C1(n9796), .C2(n9795), .A(n10151), .B(n9794), .ZN(n9797)
         );
  NAND2_X1 U11008 ( .A1(n9798), .A2(n9797), .ZN(P2_U3246) );
  AOI22_X1 U11009 ( .A1(n10162), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9809) );
  AOI211_X1 U11010 ( .C1(n9801), .C2(n9800), .A(n9799), .B(n10153), .ZN(n9802)
         );
  AOI21_X1 U11011 ( .B1(n10166), .B2(n9803), .A(n9802), .ZN(n9808) );
  OAI211_X1 U11012 ( .C1(n9806), .C2(n9805), .A(n10151), .B(n9804), .ZN(n9807)
         );
  NAND3_X1 U11013 ( .A1(n9809), .A2(n9808), .A3(n9807), .ZN(P2_U3247) );
  OAI22_X1 U11014 ( .A1(n9811), .A2(n10298), .B1(n9810), .B2(n10296), .ZN(
        n9813) );
  AOI211_X1 U11015 ( .C1(n9814), .C2(n10302), .A(n9813), .B(n9812), .ZN(n9816)
         );
  AOI22_X1 U11016 ( .A1(n10319), .A2(n9816), .B1(n7139), .B2(n10317), .ZN(
        P2_U3534) );
  INV_X1 U11017 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9815) );
  AOI22_X1 U11018 ( .A1(n10306), .A2(n9816), .B1(n9815), .B2(n10304), .ZN(
        P2_U3493) );
  INV_X1 U11019 ( .A(n9817), .ZN(n9820) );
  NOR2_X1 U11020 ( .A1(n9818), .A2(n10118), .ZN(n9819) );
  AOI22_X1 U11021 ( .A1(n4387), .A2(n9844), .B1(n5643), .B2(n10134), .ZN(
        P1_U3553) );
  OR2_X1 U11022 ( .A1(n9824), .A2(n9823), .ZN(n9830) );
  OAI21_X1 U11023 ( .B1(n9826), .B2(n10116), .A(n9825), .ZN(n9827) );
  NOR2_X1 U11024 ( .A1(n9828), .A2(n9827), .ZN(n9829) );
  AOI22_X1 U11025 ( .A1(n4387), .A2(n9845), .B1(n9066), .B2(n10134), .ZN(
        P1_U3539) );
  INV_X1 U11026 ( .A(n9831), .ZN(n9836) );
  OAI22_X1 U11027 ( .A1(n9833), .A2(n10118), .B1(n9832), .B2(n10116), .ZN(
        n9835) );
  AOI211_X1 U11028 ( .C1(n10099), .C2(n9836), .A(n9835), .B(n9834), .ZN(n9846)
         );
  AOI22_X1 U11029 ( .A1(n4387), .A2(n9846), .B1(n9837), .B2(n10134), .ZN(
        P1_U3538) );
  OAI211_X1 U11030 ( .C1(n9840), .C2(n10116), .A(n9839), .B(n9838), .ZN(n9841)
         );
  AOI21_X1 U11031 ( .B1(n10122), .B2(n9842), .A(n9841), .ZN(n9848) );
  AOI22_X1 U11032 ( .A1(n4387), .A2(n9848), .B1(n6997), .B2(n10134), .ZN(
        P1_U3537) );
  AOI22_X1 U11033 ( .A1(n10126), .A2(n9844), .B1(n9843), .B2(n10124), .ZN(
        P1_U3521) );
  AOI22_X1 U11034 ( .A1(n10126), .A2(n9845), .B1(n5413), .B2(n10124), .ZN(
        P1_U3502) );
  AOI22_X1 U11035 ( .A1(n10126), .A2(n9846), .B1(n5394), .B2(n10124), .ZN(
        P1_U3499) );
  INV_X1 U11036 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n9847) );
  AOI22_X1 U11037 ( .A1(n10126), .A2(n9848), .B1(n9847), .B2(n10124), .ZN(
        P1_U3496) );
  XNOR2_X1 U11038 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11039 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI211_X1 U11040 ( .C1(n9871), .C2(n9850), .A(n9849), .B(n9944), .ZN(n9855)
         );
  NAND2_X1 U11041 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9853) );
  AOI211_X1 U11042 ( .C1(n9853), .C2(n9852), .A(n9851), .B(n9907), .ZN(n9854)
         );
  AOI211_X1 U11043 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n9855), 
        .B(n9854), .ZN(n9859) );
  INV_X1 U11044 ( .A(n9856), .ZN(n9857) );
  AOI22_X1 U11045 ( .A1(n9955), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(n9857), .B2(
        n9950), .ZN(n9858) );
  NAND2_X1 U11046 ( .A1(n9859), .A2(n9858), .ZN(P1_U3242) );
  AOI22_X1 U11047 ( .A1(n9950), .A2(n9860), .B1(P1_REG3_REG_2__SCAN_IN), .B2(
        P1_U3084), .ZN(n9877) );
  AOI211_X1 U11048 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9907), .ZN(n9868)
         );
  AOI211_X1 U11049 ( .C1(n9866), .C2(n9865), .A(n9864), .B(n9944), .ZN(n9867)
         );
  AOI211_X1 U11050 ( .C1(P1_ADDR_REG_2__SCAN_IN), .C2(n9955), .A(n9868), .B(
        n9867), .ZN(n9876) );
  MUX2_X1 U11051 ( .A(n9871), .B(n9870), .S(n9869), .Z(n9875) );
  OAI211_X1 U11052 ( .C1(n9875), .C2(n9874), .A(n9873), .B(n9872), .ZN(n9888)
         );
  NAND3_X1 U11053 ( .A1(n9877), .A2(n9876), .A3(n9888), .ZN(P1_U3243) );
  XNOR2_X1 U11054 ( .A(n9879), .B(n9878), .ZN(n9880) );
  AOI22_X1 U11055 ( .A1(n9950), .A2(n9881), .B1(n9956), .B2(n9880), .ZN(n9890)
         );
  OAI21_X1 U11056 ( .B1(n9884), .B2(n9883), .A(n9882), .ZN(n9885) );
  AND2_X1 U11057 ( .A1(n9937), .A2(n9885), .ZN(n9886) );
  AOI211_X1 U11058 ( .C1(P1_ADDR_REG_4__SCAN_IN), .C2(n9955), .A(n9887), .B(
        n9886), .ZN(n9889) );
  NAND3_X1 U11059 ( .A1(n9890), .A2(n9889), .A3(n9888), .ZN(P1_U3245) );
  OAI21_X1 U11060 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(n9900) );
  NOR2_X1 U11061 ( .A1(n9895), .A2(n9894), .ZN(n9896) );
  NOR3_X1 U11062 ( .A1(n9907), .A2(n9897), .A3(n9896), .ZN(n9898) );
  AOI211_X1 U11063 ( .C1(n9937), .C2(n9900), .A(n9899), .B(n9898), .ZN(n9903)
         );
  AOI22_X1 U11064 ( .A1(n9955), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n9901), .B2(
        n9950), .ZN(n9902) );
  NAND2_X1 U11065 ( .A1(n9903), .A2(n9902), .ZN(P1_U3246) );
  OAI21_X1 U11066 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9913) );
  AOI211_X1 U11067 ( .C1(n9910), .C2(n9909), .A(n9908), .B(n9907), .ZN(n9911)
         );
  AOI211_X1 U11068 ( .C1(n9937), .C2(n9913), .A(n9912), .B(n9911), .ZN(n9916)
         );
  AOI22_X1 U11069 ( .A1(n9955), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n9914), .B2(
        n9950), .ZN(n9915) );
  NAND2_X1 U11070 ( .A1(n9916), .A2(n9915), .ZN(P1_U3249) );
  AOI211_X1 U11071 ( .C1(n9919), .C2(n9918), .A(n9917), .B(n9944), .ZN(n9920)
         );
  AOI21_X1 U11072 ( .B1(P1_REG3_REG_9__SCAN_IN), .B2(P1_U3084), .A(n9920), 
        .ZN(n9927) );
  OAI21_X1 U11073 ( .B1(n9923), .B2(n9922), .A(n9921), .ZN(n9925) );
  AOI22_X1 U11074 ( .A1(n9925), .A2(n9956), .B1(n9924), .B2(n9950), .ZN(n9926)
         );
  OAI211_X1 U11075 ( .C1(n9942), .C2(n10358), .A(n9927), .B(n9926), .ZN(
        P1_U3250) );
  INV_X1 U11076 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9941) );
  AOI21_X1 U11077 ( .B1(n9950), .B2(n9929), .A(n9928), .ZN(n9940) );
  OAI21_X1 U11078 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n9938) );
  OAI21_X1 U11079 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9936) );
  AOI22_X1 U11080 ( .A1(n9938), .A2(n9956), .B1(n9937), .B2(n9936), .ZN(n9939)
         );
  OAI211_X1 U11081 ( .C1(n9942), .C2(n9941), .A(n9940), .B(n9939), .ZN(
        P1_U3252) );
  INV_X1 U11082 ( .A(n9943), .ZN(n9949) );
  AOI211_X1 U11083 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9944), .ZN(n9948)
         );
  AOI211_X1 U11084 ( .C1(n9951), .C2(n9950), .A(n9949), .B(n9948), .ZN(n9959)
         );
  OAI21_X1 U11085 ( .B1(n9954), .B2(n9953), .A(n9952), .ZN(n9957) );
  AOI22_X1 U11086 ( .A1(n9957), .A2(n9956), .B1(n9955), .B2(
        P1_ADDR_REG_18__SCAN_IN), .ZN(n9958) );
  NAND2_X1 U11087 ( .A1(n9959), .A2(n9958), .ZN(P1_U3259) );
  OAI21_X1 U11088 ( .B1(n9961), .B2(n9963), .A(n9960), .ZN(n9962) );
  INV_X1 U11089 ( .A(n9962), .ZN(n10123) );
  XNOR2_X1 U11090 ( .A(n9964), .B(n9963), .ZN(n9965) );
  OAI222_X1 U11091 ( .A1(n10012), .A2(n9967), .B1(n10010), .B2(n9966), .C1(
        n9965), .C2(n9989), .ZN(n10120) );
  AOI21_X1 U11092 ( .B1(n10123), .B2(n9992), .A(n10120), .ZN(n9979) );
  INV_X1 U11093 ( .A(n9968), .ZN(n10117) );
  NOR2_X1 U11094 ( .A1(n9994), .A2(n9969), .ZN(n9970) );
  AOI21_X1 U11095 ( .B1(n10021), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9970), .ZN(
        n9971) );
  OAI21_X1 U11096 ( .B1(n10029), .B2(n10117), .A(n9971), .ZN(n9972) );
  INV_X1 U11097 ( .A(n9972), .ZN(n9978) );
  INV_X1 U11098 ( .A(n9973), .ZN(n9975) );
  OAI21_X1 U11099 ( .B1(n9975), .B2(n10117), .A(n9974), .ZN(n10119) );
  INV_X1 U11100 ( .A(n10119), .ZN(n9976) );
  AOI22_X1 U11101 ( .A1(n10123), .A2(n10004), .B1(n10003), .B2(n9976), .ZN(
        n9977) );
  OAI211_X1 U11102 ( .C1(n10021), .C2(n9979), .A(n9978), .B(n9977), .ZN(
        P1_U3283) );
  XNOR2_X1 U11103 ( .A(n9984), .B(n9980), .ZN(n10098) );
  NAND2_X1 U11104 ( .A1(n9982), .A2(n9981), .ZN(n9983) );
  XOR2_X1 U11105 ( .A(n9984), .B(n9983), .Z(n9990) );
  AOI22_X1 U11106 ( .A1(n9987), .A2(n10009), .B1(n9986), .B2(n9985), .ZN(n9988) );
  OAI21_X1 U11107 ( .B1(n9990), .B2(n9989), .A(n9988), .ZN(n9991) );
  AOI21_X1 U11108 ( .B1(n9992), .B2(n10098), .A(n9991), .ZN(n10095) );
  NOR2_X1 U11109 ( .A1(n9994), .A2(n9993), .ZN(n9995) );
  AOI21_X1 U11110 ( .B1(n10021), .B2(P1_REG2_REG_4__SCAN_IN), .A(n9995), .ZN(
        n9996) );
  OAI21_X1 U11111 ( .B1(n10029), .B2(n10093), .A(n9996), .ZN(n9997) );
  INV_X1 U11112 ( .A(n9997), .ZN(n10006) );
  NAND2_X1 U11113 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NAND2_X1 U11114 ( .A1(n10001), .A2(n10000), .ZN(n10094) );
  INV_X1 U11115 ( .A(n10094), .ZN(n10002) );
  AOI22_X1 U11116 ( .A1(n10098), .A2(n10004), .B1(n10003), .B2(n10002), .ZN(
        n10005) );
  OAI211_X1 U11117 ( .C1(n10021), .C2(n10095), .A(n10006), .B(n10005), .ZN(
        P1_U3287) );
  OAI21_X1 U11118 ( .B1(n10014), .B2(n10008), .A(n10007), .ZN(n10018) );
  INV_X1 U11119 ( .A(n10009), .ZN(n10011) );
  OAI22_X1 U11120 ( .A1(n5135), .A2(n10012), .B1(n10011), .B2(n10010), .ZN(
        n10017) );
  XNOR2_X1 U11121 ( .A(n10014), .B(n10013), .ZN(n10079) );
  NOR2_X1 U11122 ( .A1(n10079), .A2(n10015), .ZN(n10016) );
  AOI211_X1 U11123 ( .C1(n10019), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10082) );
  AOI22_X1 U11124 ( .A1(n10021), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10020), .ZN(n10035) );
  INV_X1 U11125 ( .A(n10022), .ZN(n10026) );
  NAND2_X1 U11126 ( .A1(n10024), .A2(n10023), .ZN(n10025) );
  NAND2_X1 U11127 ( .A1(n10026), .A2(n10025), .ZN(n10081) );
  OR2_X1 U11128 ( .A1(n10027), .A2(n10079), .ZN(n10031) );
  OR2_X1 U11129 ( .A1(n10029), .A2(n10028), .ZN(n10030) );
  OAI211_X1 U11130 ( .C1(n10081), .C2(n10032), .A(n10031), .B(n10030), .ZN(
        n10033) );
  INV_X1 U11131 ( .A(n10033), .ZN(n10034) );
  OAI211_X1 U11132 ( .C1(n10021), .C2(n10082), .A(n10035), .B(n10034), .ZN(
        P1_U3289) );
  INV_X1 U11133 ( .A(n10036), .ZN(n10037) );
  NOR2_X1 U11134 ( .A1(n10037), .A2(n10072), .ZN(n10062) );
  NOR2_X1 U11135 ( .A1(n10069), .A2(n10038), .ZN(P1_U3292) );
  NOR2_X1 U11136 ( .A1(n10069), .A2(n10039), .ZN(P1_U3293) );
  INV_X1 U11137 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10040) );
  NOR2_X1 U11138 ( .A1(n10069), .A2(n10040), .ZN(P1_U3294) );
  INV_X1 U11139 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10041) );
  NOR2_X1 U11140 ( .A1(n10069), .A2(n10041), .ZN(P1_U3295) );
  INV_X1 U11141 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10042) );
  NOR2_X1 U11142 ( .A1(n10069), .A2(n10042), .ZN(P1_U3296) );
  INV_X1 U11143 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n10043) );
  NOR2_X1 U11144 ( .A1(n10069), .A2(n10043), .ZN(P1_U3297) );
  INV_X1 U11145 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U11146 ( .A1(n10069), .A2(n10044), .ZN(P1_U3298) );
  INV_X1 U11147 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n10045) );
  NOR2_X1 U11148 ( .A1(n10069), .A2(n10045), .ZN(P1_U3299) );
  INV_X1 U11149 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10046) );
  NOR2_X1 U11150 ( .A1(n10069), .A2(n10046), .ZN(P1_U3300) );
  INV_X1 U11151 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n10047) );
  NOR2_X1 U11152 ( .A1(n10062), .A2(n10047), .ZN(P1_U3301) );
  INV_X1 U11153 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n10048) );
  NOR2_X1 U11154 ( .A1(n10062), .A2(n10048), .ZN(P1_U3302) );
  INV_X1 U11155 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n10049) );
  NOR2_X1 U11156 ( .A1(n10062), .A2(n10049), .ZN(P1_U3303) );
  INV_X1 U11157 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10050) );
  NOR2_X1 U11158 ( .A1(n10062), .A2(n10050), .ZN(P1_U3304) );
  NOR2_X1 U11159 ( .A1(n10062), .A2(n10051), .ZN(P1_U3305) );
  NOR2_X1 U11160 ( .A1(n10062), .A2(n10052), .ZN(P1_U3306) );
  INV_X1 U11161 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n10053) );
  NOR2_X1 U11162 ( .A1(n10062), .A2(n10053), .ZN(P1_U3307) );
  INV_X1 U11163 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U11164 ( .A1(n10062), .A2(n10054), .ZN(P1_U3308) );
  INV_X1 U11165 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10055) );
  NOR2_X1 U11166 ( .A1(n10062), .A2(n10055), .ZN(P1_U3309) );
  INV_X1 U11167 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n10056) );
  NOR2_X1 U11168 ( .A1(n10069), .A2(n10056), .ZN(P1_U3310) );
  INV_X1 U11169 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10057) );
  NOR2_X1 U11170 ( .A1(n10069), .A2(n10057), .ZN(P1_U3311) );
  INV_X1 U11171 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10058) );
  NOR2_X1 U11172 ( .A1(n10069), .A2(n10058), .ZN(P1_U3312) );
  INV_X1 U11173 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10059) );
  NOR2_X1 U11174 ( .A1(n10069), .A2(n10059), .ZN(P1_U3313) );
  INV_X1 U11175 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10060) );
  NOR2_X1 U11176 ( .A1(n10069), .A2(n10060), .ZN(P1_U3314) );
  INV_X1 U11177 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10061) );
  NOR2_X1 U11178 ( .A1(n10062), .A2(n10061), .ZN(P1_U3315) );
  NOR2_X1 U11179 ( .A1(n10069), .A2(n10063), .ZN(P1_U3316) );
  NOR2_X1 U11180 ( .A1(n10069), .A2(n10064), .ZN(P1_U3317) );
  INV_X1 U11181 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10065) );
  NOR2_X1 U11182 ( .A1(n10069), .A2(n10065), .ZN(P1_U3318) );
  INV_X1 U11183 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10066) );
  NOR2_X1 U11184 ( .A1(n10069), .A2(n10066), .ZN(P1_U3319) );
  INV_X1 U11185 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10067) );
  NOR2_X1 U11186 ( .A1(n10069), .A2(n10067), .ZN(P1_U3320) );
  INV_X1 U11187 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10068) );
  NOR2_X1 U11188 ( .A1(n10069), .A2(n10068), .ZN(P1_U3321) );
  INV_X1 U11189 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10071) );
  AOI21_X1 U11190 ( .B1(n10072), .B2(n10071), .A(n10070), .ZN(P1_U3440) );
  OAI21_X1 U11191 ( .B1(n10074), .B2(n10116), .A(n10073), .ZN(n10076) );
  AOI211_X1 U11192 ( .C1(n10099), .C2(n10077), .A(n10076), .B(n10075), .ZN(
        n10127) );
  INV_X1 U11193 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10078) );
  AOI22_X1 U11194 ( .A1(n10126), .A2(n10127), .B1(n10078), .B2(n10124), .ZN(
        P1_U3457) );
  INV_X1 U11195 ( .A(n10079), .ZN(n10085) );
  OAI21_X1 U11196 ( .B1(n10081), .B2(n10118), .A(n10080), .ZN(n10084) );
  INV_X1 U11197 ( .A(n10082), .ZN(n10083) );
  AOI211_X1 U11198 ( .C1(n10099), .C2(n10085), .A(n10084), .B(n10083), .ZN(
        n10129) );
  INV_X1 U11199 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U11200 ( .A1(n10126), .A2(n10129), .B1(n10086), .B2(n10124), .ZN(
        P1_U3460) );
  OAI22_X1 U11201 ( .A1(n10088), .A2(n10118), .B1(n10087), .B2(n10116), .ZN(
        n10090) );
  AOI211_X1 U11202 ( .C1(n10099), .C2(n10091), .A(n10090), .B(n10089), .ZN(
        n10130) );
  INV_X1 U11203 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U11204 ( .A1(n10126), .A2(n10130), .B1(n10092), .B2(n10124), .ZN(
        P1_U3463) );
  OAI22_X1 U11205 ( .A1(n10094), .A2(n10118), .B1(n10093), .B2(n10116), .ZN(
        n10097) );
  INV_X1 U11206 ( .A(n10095), .ZN(n10096) );
  AOI211_X1 U11207 ( .C1(n10099), .C2(n10098), .A(n10097), .B(n10096), .ZN(
        n10131) );
  INV_X1 U11208 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U11209 ( .A1(n10126), .A2(n10131), .B1(n10100), .B2(n10124), .ZN(
        P1_U3466) );
  NAND3_X1 U11210 ( .A1(n10102), .A2(n10101), .A3(n10122), .ZN(n10104) );
  OAI211_X1 U11211 ( .C1(n10105), .C2(n10116), .A(n10104), .B(n10103), .ZN(
        n10106) );
  NOR2_X1 U11212 ( .A1(n10107), .A2(n10106), .ZN(n10132) );
  AOI22_X1 U11213 ( .A1(n10126), .A2(n10132), .B1(n10108), .B2(n10124), .ZN(
        P1_U3469) );
  INV_X1 U11214 ( .A(n10109), .ZN(n10111) );
  NAND3_X1 U11215 ( .A1(n10112), .A2(n10111), .A3(n10110), .ZN(n10113) );
  AOI21_X1 U11216 ( .B1(n10122), .B2(n10114), .A(n10113), .ZN(n10133) );
  INV_X1 U11217 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U11218 ( .A1(n10126), .A2(n10133), .B1(n10115), .B2(n10124), .ZN(
        P1_U3475) );
  OAI22_X1 U11219 ( .A1(n10119), .A2(n10118), .B1(n10117), .B2(n10116), .ZN(
        n10121) );
  AOI211_X1 U11220 ( .C1(n10123), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        n10135) );
  INV_X1 U11221 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U11222 ( .A1(n10126), .A2(n10135), .B1(n10125), .B2(n10124), .ZN(
        P1_U3478) );
  AOI22_X1 U11223 ( .A1(n4387), .A2(n10127), .B1(n6235), .B2(n10134), .ZN(
        P1_U3524) );
  AOI22_X1 U11224 ( .A1(n4387), .A2(n10129), .B1(n10128), .B2(n10134), .ZN(
        P1_U3525) );
  AOI22_X1 U11225 ( .A1(n4387), .A2(n10130), .B1(n5162), .B2(n10134), .ZN(
        P1_U3526) );
  AOI22_X1 U11226 ( .A1(n4387), .A2(n10131), .B1(n6330), .B2(n10134), .ZN(
        P1_U3527) );
  AOI22_X1 U11227 ( .A1(n4387), .A2(n10132), .B1(n5196), .B2(n10134), .ZN(
        P1_U3528) );
  AOI22_X1 U11228 ( .A1(n4387), .A2(n10133), .B1(n5231), .B2(n10134), .ZN(
        P1_U3530) );
  AOI22_X1 U11229 ( .A1(n4387), .A2(n10135), .B1(n6358), .B2(n10134), .ZN(
        P1_U3531) );
  NAND2_X1 U11230 ( .A1(n10136), .A2(n5806), .ZN(n10147) );
  NAND2_X1 U11231 ( .A1(n10137), .A2(n10206), .ZN(n10146) );
  OAI21_X1 U11232 ( .B1(n10140), .B2(n10139), .A(n10138), .ZN(n10142) );
  NAND2_X1 U11233 ( .A1(n10142), .A2(n10141), .ZN(n10145) );
  OR2_X1 U11234 ( .A1(n10143), .A2(n10246), .ZN(n10144) );
  AND4_X1 U11235 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10148) );
  OAI21_X1 U11236 ( .B1(n10150), .B2(n10149), .A(n10148), .ZN(P2_U3224) );
  AOI22_X1 U11237 ( .A1(n10151), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n10168), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U11238 ( .A1(n10162), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10157) );
  NOR2_X1 U11239 ( .A1(n10172), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10155) );
  OAI21_X1 U11240 ( .B1(n10153), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10152), .ZN(
        n10154) );
  OAI21_X1 U11241 ( .B1(n10155), .B2(n10154), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10156) );
  OAI211_X1 U11242 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10158), .A(n10157), .B(
        n10156), .ZN(P2_U3245) );
  AOI21_X1 U11243 ( .B1(n10161), .B2(n10160), .A(n10159), .ZN(n10173) );
  AOI22_X1 U11244 ( .A1(n10162), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n10171) );
  OAI21_X1 U11245 ( .B1(n10165), .B2(n10164), .A(n10163), .ZN(n10169) );
  AOI22_X1 U11246 ( .A1(n10169), .A2(n10168), .B1(n10167), .B2(n10166), .ZN(
        n10170) );
  OAI211_X1 U11247 ( .C1(n10173), .C2(n10172), .A(n10171), .B(n10170), .ZN(
        P2_U3258) );
  AOI21_X1 U11248 ( .B1(n10174), .B2(n10179), .A(n6148), .ZN(n10177) );
  AOI21_X1 U11249 ( .B1(n10177), .B2(n10176), .A(n10175), .ZN(n10264) );
  XNOR2_X1 U11250 ( .A(n10178), .B(n10179), .ZN(n10267) );
  XNOR2_X1 U11251 ( .A(n10196), .B(n10182), .ZN(n10263) );
  OAI22_X1 U11252 ( .A1(n10222), .A2(n5822), .B1(n10180), .B2(n10218), .ZN(
        n10181) );
  AOI21_X1 U11253 ( .B1(n10183), .B2(n10182), .A(n10181), .ZN(n10184) );
  OAI21_X1 U11254 ( .B1(n10219), .B2(n10263), .A(n10184), .ZN(n10185) );
  AOI21_X1 U11255 ( .B1(n10267), .B2(n10202), .A(n10185), .ZN(n10186) );
  OAI21_X1 U11256 ( .B1(n10224), .B2(n10264), .A(n10186), .ZN(P2_U3292) );
  XNOR2_X1 U11257 ( .A(n10188), .B(n10187), .ZN(n10192) );
  AOI222_X1 U11258 ( .A1(n10193), .A2(n10192), .B1(n10191), .B2(n10190), .C1(
        n5806), .C2(n10189), .ZN(n10258) );
  XNOR2_X1 U11259 ( .A(n10195), .B(n10194), .ZN(n10261) );
  OAI21_X1 U11260 ( .B1(n10197), .B2(n10256), .A(n10196), .ZN(n10257) );
  OAI22_X1 U11261 ( .A1(n10219), .A2(n10257), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n10218), .ZN(n10198) );
  AOI21_X1 U11262 ( .B1(n10224), .B2(P2_REG2_REG_3__SCAN_IN), .A(n10198), .ZN(
        n10199) );
  OAI21_X1 U11263 ( .B1(n10256), .B2(n10200), .A(n10199), .ZN(n10201) );
  AOI21_X1 U11264 ( .B1(n10202), .B2(n10261), .A(n10201), .ZN(n10203) );
  OAI21_X1 U11265 ( .B1(n10224), .B2(n10258), .A(n10203), .ZN(P2_U3293) );
  XNOR2_X1 U11266 ( .A(n10204), .B(n8401), .ZN(n10250) );
  NOR2_X1 U11267 ( .A1(n10246), .A2(n10205), .ZN(n10212) );
  INV_X1 U11268 ( .A(n10206), .ZN(n10209) );
  XOR2_X1 U11269 ( .A(n8401), .B(n10207), .Z(n10208) );
  OAI222_X1 U11270 ( .A1(n10211), .A2(n5805), .B1(n10210), .B2(n10209), .C1(
        n6148), .C2(n10208), .ZN(n10248) );
  AOI211_X1 U11271 ( .C1(n10213), .C2(n10250), .A(n10212), .B(n10248), .ZN(
        n10223) );
  NAND2_X1 U11272 ( .A1(n10215), .A2(n10214), .ZN(n10216) );
  NAND2_X1 U11273 ( .A1(n10217), .A2(n10216), .ZN(n10247) );
  OAI22_X1 U11274 ( .A1(n10219), .A2(n10247), .B1(n10149), .B2(n10218), .ZN(
        n10220) );
  INV_X1 U11275 ( .A(n10220), .ZN(n10221) );
  OAI221_X1 U11276 ( .B1(n10224), .B2(n10223), .C1(n10222), .C2(n5771), .A(
        n10221), .ZN(P2_U3295) );
  NOR2_X1 U11277 ( .A1(n10234), .A2(n10225), .ZN(n10235) );
  AND2_X1 U11278 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10237), .ZN(P2_U3297) );
  AND2_X1 U11279 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10237), .ZN(P2_U3298) );
  NOR2_X1 U11280 ( .A1(n10235), .A2(n10226), .ZN(P2_U3299) );
  AND2_X1 U11281 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10237), .ZN(P2_U3300) );
  AND2_X1 U11282 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10237), .ZN(P2_U3301) );
  AND2_X1 U11283 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10237), .ZN(P2_U3302) );
  NOR2_X1 U11284 ( .A1(n10235), .A2(n10227), .ZN(P2_U3303) );
  AND2_X1 U11285 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10237), .ZN(P2_U3304) );
  AND2_X1 U11286 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10237), .ZN(P2_U3305) );
  AND2_X1 U11287 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10237), .ZN(P2_U3306) );
  AND2_X1 U11288 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10237), .ZN(P2_U3307) );
  AND2_X1 U11289 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10237), .ZN(P2_U3308) );
  NOR2_X1 U11290 ( .A1(n10235), .A2(n10228), .ZN(P2_U3309) );
  AND2_X1 U11291 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10237), .ZN(P2_U3310) );
  AND2_X1 U11292 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10237), .ZN(P2_U3311) );
  NOR2_X1 U11293 ( .A1(n10235), .A2(n10229), .ZN(P2_U3312) );
  AND2_X1 U11294 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10237), .ZN(P2_U3313) );
  NOR2_X1 U11295 ( .A1(n10235), .A2(n10230), .ZN(P2_U3314) );
  AND2_X1 U11296 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10237), .ZN(P2_U3315) );
  AND2_X1 U11297 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10237), .ZN(P2_U3316) );
  AND2_X1 U11298 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10237), .ZN(P2_U3317) );
  AND2_X1 U11299 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10237), .ZN(P2_U3318) );
  AND2_X1 U11300 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10237), .ZN(P2_U3319) );
  AND2_X1 U11301 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10237), .ZN(P2_U3320) );
  AND2_X1 U11302 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10237), .ZN(P2_U3321) );
  NOR2_X1 U11303 ( .A1(n10235), .A2(n10231), .ZN(P2_U3322) );
  AND2_X1 U11304 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10237), .ZN(P2_U3323) );
  AND2_X1 U11305 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10237), .ZN(P2_U3324) );
  AND2_X1 U11306 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10237), .ZN(P2_U3325) );
  NOR2_X1 U11307 ( .A1(n10235), .A2(n10232), .ZN(P2_U3326) );
  OAI22_X1 U11308 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10235), .B1(n10234), .B2(
        n10233), .ZN(n10236) );
  INV_X1 U11309 ( .A(n10236), .ZN(P2_U3437) );
  AOI22_X1 U11310 ( .A1(n10240), .A2(n10239), .B1(n10238), .B2(n10237), .ZN(
        P2_U3438) );
  OAI21_X1 U11311 ( .B1(n10243), .B2(n10242), .A(n10241), .ZN(n10244) );
  AOI21_X1 U11312 ( .B1(n10245), .B2(n10302), .A(n10244), .ZN(n10307) );
  AOI22_X1 U11313 ( .A1(n10306), .A2(n10307), .B1(n5781), .B2(n10304), .ZN(
        P2_U3451) );
  OAI22_X1 U11314 ( .A1(n10247), .A2(n10298), .B1(n10296), .B2(n10246), .ZN(
        n10249) );
  AOI211_X1 U11315 ( .C1(n10302), .C2(n10250), .A(n10249), .B(n10248), .ZN(
        n10308) );
  AOI22_X1 U11316 ( .A1(n10306), .A2(n10308), .B1(n5772), .B2(n10304), .ZN(
        P2_U3454) );
  OAI22_X1 U11317 ( .A1(n10252), .A2(n10298), .B1(n10251), .B2(n10296), .ZN(
        n10254) );
  AOI211_X1 U11318 ( .C1(n10302), .C2(n10255), .A(n10254), .B(n10253), .ZN(
        n10309) );
  AOI22_X1 U11319 ( .A1(n10306), .A2(n10309), .B1(n5792), .B2(n10304), .ZN(
        P2_U3457) );
  OAI22_X1 U11320 ( .A1(n10257), .A2(n10298), .B1(n10256), .B2(n10296), .ZN(
        n10260) );
  INV_X1 U11321 ( .A(n10258), .ZN(n10259) );
  AOI211_X1 U11322 ( .C1(n10261), .C2(n10302), .A(n10260), .B(n10259), .ZN(
        n10311) );
  AOI22_X1 U11323 ( .A1(n10306), .A2(n10311), .B1(n5810), .B2(n10304), .ZN(
        P2_U3460) );
  OAI22_X1 U11324 ( .A1(n10263), .A2(n10298), .B1(n10262), .B2(n10296), .ZN(
        n10266) );
  INV_X1 U11325 ( .A(n10264), .ZN(n10265) );
  AOI211_X1 U11326 ( .C1(n10302), .C2(n10267), .A(n10266), .B(n10265), .ZN(
        n10312) );
  INV_X1 U11327 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10268) );
  AOI22_X1 U11328 ( .A1(n10306), .A2(n10312), .B1(n10268), .B2(n10304), .ZN(
        P2_U3463) );
  OAI21_X1 U11329 ( .B1(n10270), .B2(n10296), .A(n10269), .ZN(n10272) );
  AOI211_X1 U11330 ( .C1(n10302), .C2(n10273), .A(n10272), .B(n10271), .ZN(
        n10313) );
  INV_X1 U11331 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10274) );
  AOI22_X1 U11332 ( .A1(n10306), .A2(n10313), .B1(n10274), .B2(n10304), .ZN(
        P2_U3466) );
  OAI22_X1 U11333 ( .A1(n10276), .A2(n10298), .B1(n10275), .B2(n10296), .ZN(
        n10278) );
  AOI211_X1 U11334 ( .C1(n10279), .C2(n10302), .A(n10278), .B(n10277), .ZN(
        n10314) );
  AOI22_X1 U11335 ( .A1(n10306), .A2(n10314), .B1(n10280), .B2(n10304), .ZN(
        P2_U3469) );
  OAI22_X1 U11336 ( .A1(n10282), .A2(n10298), .B1(n10281), .B2(n10296), .ZN(
        n10283) );
  AOI211_X1 U11337 ( .C1(n10285), .C2(n10302), .A(n10284), .B(n10283), .ZN(
        n10315) );
  INV_X1 U11338 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10286) );
  AOI22_X1 U11339 ( .A1(n10306), .A2(n10315), .B1(n10286), .B2(n10304), .ZN(
        P2_U3475) );
  INV_X1 U11340 ( .A(n10287), .ZN(n10292) );
  OAI22_X1 U11341 ( .A1(n10289), .A2(n10298), .B1(n10288), .B2(n10296), .ZN(
        n10291) );
  AOI211_X1 U11342 ( .C1(n10293), .C2(n10292), .A(n10291), .B(n10290), .ZN(
        n10316) );
  INV_X1 U11343 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10294) );
  AOI22_X1 U11344 ( .A1(n10306), .A2(n10316), .B1(n10294), .B2(n10304), .ZN(
        P2_U3481) );
  INV_X1 U11345 ( .A(n10295), .ZN(n10297) );
  OAI22_X1 U11346 ( .A1(n10299), .A2(n10298), .B1(n10297), .B2(n10296), .ZN(
        n10301) );
  AOI211_X1 U11347 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10318) );
  INV_X1 U11348 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U11349 ( .A1(n10306), .A2(n10318), .B1(n10305), .B2(n10304), .ZN(
        P2_U3487) );
  AOI22_X1 U11350 ( .A1(n10319), .A2(n10307), .B1(n5780), .B2(n10317), .ZN(
        P2_U3520) );
  AOI22_X1 U11351 ( .A1(n10319), .A2(n10308), .B1(n6403), .B2(n10317), .ZN(
        P2_U3521) );
  AOI22_X1 U11352 ( .A1(n10319), .A2(n10309), .B1(n5790), .B2(n10317), .ZN(
        P2_U3522) );
  INV_X1 U11353 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U11354 ( .A1(n10319), .A2(n10311), .B1(n10310), .B2(n10317), .ZN(
        P2_U3523) );
  AOI22_X1 U11355 ( .A1(n10319), .A2(n10312), .B1(n6406), .B2(n10317), .ZN(
        P2_U3524) );
  AOI22_X1 U11356 ( .A1(n10319), .A2(n10313), .B1(n5838), .B2(n10317), .ZN(
        P2_U3525) );
  AOI22_X1 U11357 ( .A1(n10319), .A2(n10314), .B1(n6427), .B2(n10317), .ZN(
        P2_U3526) );
  AOI22_X1 U11358 ( .A1(n10319), .A2(n10315), .B1(n6511), .B2(n10317), .ZN(
        P2_U3528) );
  AOI22_X1 U11359 ( .A1(n10319), .A2(n10316), .B1(n5909), .B2(n10317), .ZN(
        P2_U3530) );
  AOI22_X1 U11360 ( .A1(n10319), .A2(n10318), .B1(n5936), .B2(n10317), .ZN(
        P2_U3532) );
  INV_X1 U11361 ( .A(n10320), .ZN(n10321) );
  NAND2_X1 U11362 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  XNOR2_X1 U11363 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10323), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11364 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11365 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(ADD_1071_U56) );
  OAI21_X1 U11366 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(ADD_1071_U57) );
  OAI21_X1 U11367 ( .B1(n10332), .B2(n10331), .A(n10330), .ZN(ADD_1071_U58) );
  OAI21_X1 U11368 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(ADD_1071_U59) );
  OAI21_X1 U11369 ( .B1(n10338), .B2(n10337), .A(n10336), .ZN(ADD_1071_U60) );
  OAI21_X1 U11370 ( .B1(n10341), .B2(n10340), .A(n10339), .ZN(ADD_1071_U61) );
  AOI21_X1 U11371 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(ADD_1071_U62) );
  AOI21_X1 U11372 ( .B1(n10347), .B2(n10346), .A(n10345), .ZN(ADD_1071_U63) );
  XOR2_X1 U11373 ( .A(n10348), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11374 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  XOR2_X1 U11375 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10351), .Z(ADD_1071_U51) );
  OAI21_X1 U11376 ( .B1(n10354), .B2(n10353), .A(n10352), .ZN(n10355) );
  XNOR2_X1 U11377 ( .A(n10355), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11378 ( .B1(n10358), .B2(n10357), .A(n10356), .ZN(ADD_1071_U47) );
  XOR2_X1 U11379 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10359), .Z(ADD_1071_U48) );
  XOR2_X1 U11380 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10360), .Z(ADD_1071_U49) );
  XOR2_X1 U11381 ( .A(n10362), .B(n10361), .Z(ADD_1071_U54) );
  XOR2_X1 U11382 ( .A(n10364), .B(n10363), .Z(ADD_1071_U53) );
  XNOR2_X1 U11383 ( .A(n10366), .B(n10365), .ZN(ADD_1071_U52) );
  INV_X2 U8283 ( .A(n6493), .ZN(n6674) );
  CLKBUF_X1 U4895 ( .A(n5336), .Z(n4502) );
  CLKBUF_X1 U4939 ( .A(n5791), .Z(n6110) );
  CLKBUF_X1 U4942 ( .A(n5179), .Z(n6480) );
  CLKBUF_X1 U5001 ( .A(n5719), .Z(n4392) );
endmodule

