

module b22_C_SARLock_k_128_6 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, 
        SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, 
        SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, 
        SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, 
        U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, 
        P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, 
        P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, 
        P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, 
        P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, 
        P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, 
        P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, 
        P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, 
        P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, 
        P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, 
        P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, 
        P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, 
        P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, 
        P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, 
        P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, 
        P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, 
        P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, 
        P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, 
        P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, 
        P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, 
        P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, 
        P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, 
        P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, 
        P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, 
        P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, 
        P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, 
        P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, 
        P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, 
        P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, 
        P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, 
        P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, 
        P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, 
        P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, 
        P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, 
        P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, 
        P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, 
        P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, 
        P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, 
        P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, 
        P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, 
        P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, 
        P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, 
        P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, 
        P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, 
        P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, 
        P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, 
        P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, 
        P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, 
        P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, 
        P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63, keyinput64, keyinput65, keyinput66, keyinput67,
         keyinput68, keyinput69, keyinput70, keyinput71, keyinput72,
         keyinput73, keyinput74, keyinput75, keyinput76, keyinput77,
         keyinput78, keyinput79, keyinput80, keyinput81, keyinput82,
         keyinput83, keyinput84, keyinput85, keyinput86, keyinput87,
         keyinput88, keyinput89, keyinput90, keyinput91, keyinput92,
         keyinput93, keyinput94, keyinput95, keyinput96, keyinput97,
         keyinput98, keyinput99, keyinput100, keyinput101, keyinput102,
         keyinput103, keyinput104, keyinput105, keyinput106, keyinput107,
         keyinput108, keyinput109, keyinput110, keyinput111, keyinput112,
         keyinput113, keyinput114, keyinput115, keyinput116, keyinput117,
         keyinput118, keyinput119, keyinput120, keyinput121, keyinput122,
         keyinput123, keyinput124, keyinput125, keyinput126, keyinput127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438;

  AOI211_X1 U7291 ( .C1(n14899), .C2(n14361), .A(n14195), .B(n14194), .ZN(
        n14365) );
  OR2_X1 U7292 ( .A1(n13302), .A2(n13156), .ZN(n13145) );
  AOI21_X1 U7293 ( .B1(n15228), .B2(n15227), .A(n15226), .ZN(n15245) );
  OAI21_X1 U7294 ( .B1(n15175), .B2(n15174), .A(n15173), .ZN(n15192) );
  INV_X1 U7295 ( .A(n7604), .ZN(n7980) );
  CLKBUF_X2 U7296 ( .A(n7424), .Z(n11036) );
  INV_X4 U7297 ( .A(n13729), .ZN(n9891) );
  INV_X1 U7298 ( .A(n11242), .ZN(n15320) );
  INV_X1 U7300 ( .A(n7558), .ZN(n10733) );
  CLKBUF_X2 U7301 ( .A(n7546), .Z(n12033) );
  AND3_X1 U7302 ( .A1(n7540), .A2(n7539), .A3(n7538), .ZN(n10956) );
  AND2_X1 U7303 ( .A1(n7506), .A2(n12771), .ZN(n7515) );
  NAND2_X1 U7304 ( .A1(n10577), .A2(n9960), .ZN(n12035) );
  NAND2_X2 U7305 ( .A1(n7985), .A2(n7986), .ZN(n10577) );
  INV_X1 U7306 ( .A(n9847), .ZN(n10810) );
  INV_X2 U7307 ( .A(n8789), .ZN(n8414) );
  INV_X2 U7308 ( .A(n8212), .ZN(n8789) );
  AND2_X1 U7309 ( .A1(n7262), .A2(n9313), .ZN(n8981) );
  AOI22_X1 U7310 ( .A1(n13553), .A2(keyinput73), .B1(keyinput68), .B2(n13877), 
        .ZN(n13552) );
  NAND2_X1 U7311 ( .A1(n9866), .A2(n9861), .ZN(n9886) );
  INV_X1 U7312 ( .A(n7515), .ZN(n7826) );
  NAND2_X1 U7313 ( .A1(n7985), .A2(n7986), .ZN(n6550) );
  AND3_X1 U7314 ( .A1(n7554), .A2(n7553), .A3(n7552), .ZN(n11037) );
  INV_X1 U7315 ( .A(n8718), .ZN(n8745) );
  NAND2_X1 U7316 ( .A1(n12110), .A2(n12111), .ZN(n11564) );
  NAND2_X1 U7317 ( .A1(n6868), .A2(n6869), .ZN(n12013) );
  INV_X1 U7318 ( .A(n12484), .ZN(n11922) );
  OR2_X1 U7320 ( .A1(n12350), .A2(n6693), .ZN(n6692) );
  INV_X2 U7321 ( .A(n8563), .ZN(n9770) );
  AND2_X1 U7322 ( .A1(n13379), .A2(n11823), .ZN(n8719) );
  NAND2_X1 U7323 ( .A1(n13798), .A2(n9951), .ZN(n13728) );
  BUF_X1 U7324 ( .A(n9008), .Z(n10033) );
  INV_X1 U7325 ( .A(n10684), .ZN(n9952) );
  NAND2_X1 U7326 ( .A1(n9864), .A2(n10684), .ZN(n9861) );
  CLKBUF_X2 U7327 ( .A(n13679), .Z(n6549) );
  NOR2_X1 U7328 ( .A1(n12696), .A2(n10751), .ZN(n12701) );
  CLKBUF_X3 U7329 ( .A(n7530), .Z(n6547) );
  AND4_X1 U7330 ( .A1(n7609), .A2(n7608), .A3(n7607), .A4(n7606), .ZN(n11746)
         );
  AND3_X1 U7331 ( .A1(n7022), .A2(n7024), .A3(n7532), .ZN(n12698) );
  XNOR2_X1 U7332 ( .A(n7500), .B(P3_IR_REG_30__SCAN_IN), .ZN(n7506) );
  AOI21_X1 U7333 ( .B1(n14129), .B2(n14766), .A(n14128), .ZN(n14340) );
  INV_X1 U7334 ( .A(n11746), .ZN(n12255) );
  NAND4_X1 U7335 ( .A1(n7513), .A2(n7512), .A3(n7511), .A4(n7510), .ZN(n12696)
         );
  CLKBUF_X3 U7336 ( .A(n7986), .Z(n12774) );
  BUF_X1 U7337 ( .A(n10595), .Z(n6546) );
  AND2_X1 U7338 ( .A1(n14070), .A2(n14069), .ZN(n6542) );
  OR2_X1 U7339 ( .A1(n7798), .A2(n6623), .ZN(n6543) );
  NOR2_X2 U7340 ( .A1(n15207), .A2(n15206), .ZN(n15205) );
  XNOR2_X2 U7341 ( .A(n7018), .B(n15214), .ZN(n15206) );
  NAND4_X2 U7342 ( .A1(n9052), .A2(n9051), .A3(n9050), .A4(n9049), .ZN(n13920)
         );
  OAI21_X2 U7343 ( .B1(n13228), .B2(n8866), .A(n9811), .ZN(n13218) );
  INV_X1 U7344 ( .A(n9184), .ZN(n6544) );
  AOI21_X2 U7345 ( .B1(n10707), .B2(n10704), .A(n10999), .ZN(n8360) );
  NAND2_X2 U7346 ( .A1(n7129), .A2(n8329), .ZN(n10707) );
  AND2_X2 U7347 ( .A1(n7693), .A2(n6573), .ZN(n7992) );
  AND4_X2 U7348 ( .A1(n7482), .A2(n7628), .A3(n7026), .A4(n7025), .ZN(n7693)
         );
  OAI21_X2 U7349 ( .B1(n11419), .B2(n7939), .A(n7938), .ZN(n11485) );
  NAND2_X2 U7350 ( .A1(n7937), .A2(n7936), .ZN(n11419) );
  NOR2_X2 U7351 ( .A1(n11432), .A2(n11431), .ZN(n11692) );
  NOR2_X2 U7352 ( .A1(n11521), .A2(n11430), .ZN(n11432) );
  OAI21_X2 U7353 ( .B1(n10865), .B2(n10864), .A(n10863), .ZN(n14799) );
  OR2_X2 U7354 ( .A1(n8690), .A2(n8689), .ZN(n8692) );
  INV_X2 U7355 ( .A(n8719), .ZN(n8563) );
  INV_X4 U7356 ( .A(n9213), .ZN(n9327) );
  AOI21_X2 U7357 ( .B1(n11904), .B2(n6547), .A(n7903), .ZN(n12417) );
  NOR2_X4 U7358 ( .A1(n8206), .A2(n8205), .ZN(n10074) );
  BUF_X2 U7359 ( .A(n9322), .Z(n6545) );
  INV_X1 U7360 ( .A(n9008), .ZN(n9322) );
  XNOR2_X2 U7361 ( .A(n11847), .B(n11845), .ZN(n11919) );
  AOI21_X2 U7362 ( .B1(n11996), .B2(n11843), .A(n11842), .ZN(n11847) );
  OAI21_X2 U7363 ( .B1(n11239), .B2(n7934), .A(n7933), .ZN(n7937) );
  OAI21_X2 U7364 ( .B1(n7929), .B2(n11404), .A(n7928), .ZN(n11239) );
  AOI21_X2 U7365 ( .B1(n15192), .B2(n15191), .A(n15190), .ZN(n15210) );
  OAI21_X2 U7366 ( .B1(n15278), .B2(n6570), .A(n7012), .ZN(n11429) );
  OR2_X2 U7367 ( .A1(n11073), .A2(n11428), .ZN(n6570) );
  NOR2_X2 U7368 ( .A1(n15280), .A2(n15279), .ZN(n15278) );
  OAI21_X2 U7369 ( .B1(n15210), .B2(n15209), .A(n15208), .ZN(n15228) );
  NAND2_X1 U7370 ( .A1(n7160), .A2(n7159), .ZN(n13278) );
  NAND2_X1 U7371 ( .A1(n14164), .A2(n7248), .ZN(n7250) );
  NOR2_X2 U7372 ( .A1(n12414), .A2(n6655), .ZN(n7979) );
  INV_X2 U7373 ( .A(n9807), .ZN(n13090) );
  AND2_X1 U7374 ( .A1(n12364), .A2(n7010), .ZN(n12345) );
  NAND2_X1 U7375 ( .A1(n6942), .A2(n11012), .ZN(n11161) );
  OR2_X1 U7376 ( .A1(n10982), .A2(n11014), .ZN(n11010) );
  NAND2_X1 U7377 ( .A1(n10629), .A2(n10628), .ZN(n7129) );
  INV_X1 U7378 ( .A(n11669), .ZN(n11744) );
  INV_X2 U7379 ( .A(n11036), .ZN(n11898) );
  NAND2_X1 U7380 ( .A1(n13219), .A2(n12982), .ZN(n8306) );
  INV_X1 U7381 ( .A(n12698), .ZN(n10825) );
  INV_X1 U7382 ( .A(n15339), .ZN(n12258) );
  INV_X1 U7383 ( .A(n15341), .ZN(n10506) );
  INV_X1 U7384 ( .A(n12983), .ZN(n10481) );
  AND4_X1 U7385 ( .A1(n7545), .A2(n7544), .A3(n7543), .A4(n7542), .ZN(n15339)
         );
  AND4_X1 U7386 ( .A1(n7595), .A2(n7594), .A3(n7593), .A4(n7592), .ZN(n11667)
         );
  INV_X1 U7387 ( .A(n12985), .ZN(n7134) );
  BUF_X2 U7388 ( .A(n7515), .Z(n10734) );
  CLKBUF_X2 U7389 ( .A(n9071), .Z(n9475) );
  BUF_X2 U7390 ( .A(n8234), .Z(n8662) );
  AND2_X1 U7392 ( .A1(n12769), .A2(n7505), .ZN(n7588) );
  XNOR2_X1 U7393 ( .A(n9010), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9864) );
  OR2_X1 U7394 ( .A1(n8188), .A2(n9960), .ZN(n8693) );
  INV_X1 U7395 ( .A(n7505), .ZN(n12771) );
  NAND2_X1 U7396 ( .A1(n13379), .A2(n8179), .ZN(n8213) );
  XNOR2_X1 U7397 ( .A(n7537), .B(P3_IR_REG_2__SCAN_IN), .ZN(n11119) );
  NOR2_X1 U7398 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8135) );
  OR2_X1 U7399 ( .A1(n9849), .A2(n9848), .ZN(n7304) );
  XNOR2_X1 U7400 ( .A(n8887), .B(n9806), .ZN(n13268) );
  OAI22_X1 U7401 ( .A1(n9450), .A2(n7295), .B1(n9451), .B2(n7296), .ZN(n9464)
         );
  NAND2_X1 U7402 ( .A1(n13278), .A2(n8877), .ZN(n13069) );
  AND2_X1 U7403 ( .A1(n13272), .A2(n13271), .ZN(n6812) );
  NAND2_X1 U7404 ( .A1(n8876), .A2(n7161), .ZN(n7160) );
  NAND2_X1 U7405 ( .A1(n6722), .A2(n14099), .ZN(n14176) );
  AND2_X1 U7406 ( .A1(n6958), .A2(n14335), .ZN(n6836) );
  NAND2_X1 U7407 ( .A1(n7250), .A2(n6607), .ZN(n14120) );
  AOI21_X1 U7408 ( .B1(n12811), .B2(n8647), .A(n8646), .ZN(n8648) );
  NAND2_X1 U7409 ( .A1(n13766), .A2(n13765), .ZN(n13889) );
  AND2_X1 U7410 ( .A1(n7055), .A2(n7063), .ZN(n7054) );
  OR2_X1 U7411 ( .A1(n6576), .A2(n6834), .ZN(n7238) );
  CLKBUF_X1 U7412 ( .A(n14250), .Z(n6721) );
  NAND2_X1 U7413 ( .A1(n11897), .A2(n11896), .ZN(n11913) );
  AOI21_X1 U7414 ( .B1(n6571), .B2(n15323), .A(n8821), .ZN(n6774) );
  NAND2_X1 U7415 ( .A1(n9532), .A2(n14081), .ZN(n14123) );
  OR2_X1 U7416 ( .A1(n7227), .A2(n14100), .ZN(n7222) );
  NAND2_X1 U7417 ( .A1(n6977), .A2(n6975), .ZN(n13117) );
  XNOR2_X1 U7418 ( .A(n7174), .B(n7173), .ZN(n14604) );
  OR2_X1 U7419 ( .A1(n14140), .A2(n6580), .ZN(n7227) );
  NAND2_X1 U7420 ( .A1(n12345), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n12365) );
  CLKBUF_X1 U7421 ( .A(n13165), .Z(n6714) );
  AOI21_X1 U7422 ( .B1(n7978), .B2(n12508), .A(n6614), .ZN(n6797) );
  NAND2_X2 U7423 ( .A1(n8717), .A2(n8716), .ZN(n13280) );
  NAND2_X1 U7424 ( .A1(n6940), .A2(n6938), .ZN(n14302) );
  NAND2_X1 U7425 ( .A1(n9448), .A2(n9447), .ZN(n14343) );
  NAND2_X1 U7426 ( .A1(n12508), .A2(n12516), .ZN(n12507) );
  XNOR2_X1 U7427 ( .A(n11841), .B(n11839), .ZN(n11996) );
  NAND2_X1 U7428 ( .A1(n11934), .A2(n11838), .ZN(n11841) );
  NAND2_X1 U7429 ( .A1(n9413), .A2(n9412), .ZN(n14356) );
  NAND2_X1 U7430 ( .A1(n8692), .A2(n8691), .ZN(n13390) );
  NAND2_X1 U7431 ( .A1(n8655), .A2(n8654), .ZN(n13297) );
  NOR2_X1 U7432 ( .A1(n12307), .A2(n12306), .ZN(n12309) );
  NAND2_X1 U7433 ( .A1(n7356), .A2(n7355), .ZN(n13883) );
  NOR2_X1 U7434 ( .A1(n12287), .A2(n12288), .ZN(n12307) );
  NOR2_X1 U7435 ( .A1(n13023), .A2(n6924), .ZN(n13038) );
  OR2_X1 U7436 ( .A1(n12286), .A2(n7017), .ZN(n7015) );
  OAI21_X1 U7437 ( .B1(n11471), .B2(n8924), .A(n8923), .ZN(n11537) );
  NAND2_X1 U7438 ( .A1(n8621), .A2(n8620), .ZN(n13302) );
  NAND2_X1 U7439 ( .A1(n9381), .A2(n9380), .ZN(n14369) );
  OAI21_X1 U7440 ( .B1(n8619), .B2(n11190), .A(n8123), .ZN(n8125) );
  NAND2_X1 U7441 ( .A1(n11161), .A2(n11160), .ZN(n11220) );
  OR2_X1 U7442 ( .A1(n8120), .A2(n8121), .ZN(n8122) );
  NAND2_X1 U7443 ( .A1(n8120), .A2(n8121), .ZN(n8123) );
  NAND2_X1 U7444 ( .A1(n8616), .A2(n8119), .ZN(n8120) );
  NAND2_X1 U7445 ( .A1(n9324), .A2(n9323), .ZN(n14392) );
  NAND2_X1 U7446 ( .A1(n8537), .A2(n8536), .ZN(n13328) );
  NAND3_X1 U7447 ( .A1(n6814), .A2(n8119), .A3(n8118), .ZN(n8616) );
  NAND2_X1 U7448 ( .A1(n8115), .A2(n13626), .ZN(n6814) );
  OAI21_X2 U7449 ( .B1(n10538), .B2(n9417), .A(n9304), .ZN(n14398) );
  INV_X1 U7450 ( .A(n11477), .ZN(n6548) );
  NAND2_X1 U7451 ( .A1(n8116), .A2(SI_22_), .ZN(n8119) );
  NAND2_X1 U7452 ( .A1(n6723), .A2(n10973), .ZN(n14767) );
  NAND2_X1 U7453 ( .A1(n9237), .A2(n9236), .ZN(n14658) );
  NAND2_X1 U7454 ( .A1(n10360), .A2(n8264), .ZN(n10466) );
  NAND2_X1 U7455 ( .A1(n8494), .A2(n8493), .ZN(n13339) );
  OR2_X1 U7456 ( .A1(n8108), .A2(n10690), .ZN(n8111) );
  NAND2_X1 U7457 ( .A1(n7121), .A2(n7120), .ZN(n10360) );
  NAND2_X1 U7458 ( .A1(n11487), .A2(n12121), .ZN(n15307) );
  NAND2_X1 U7459 ( .A1(n8241), .A2(n8240), .ZN(n7121) );
  NAND2_X1 U7460 ( .A1(n7197), .A2(n7196), .ZN(n10855) );
  NAND2_X1 U7461 ( .A1(n8411), .A2(n8410), .ZN(n13348) );
  OR2_X1 U7462 ( .A1(n11043), .A2(n11040), .ZN(n11269) );
  NOR2_X1 U7463 ( .A1(n10958), .A2(n10957), .ZN(n11043) );
  NAND2_X1 U7464 ( .A1(n7020), .A2(n6594), .ZN(n15258) );
  NAND2_X1 U7465 ( .A1(n8089), .A2(n7315), .ZN(n7314) );
  NAND2_X1 U7466 ( .A1(n7199), .A2(n7198), .ZN(n10853) );
  NAND2_X1 U7467 ( .A1(n6820), .A2(n6818), .ZN(n8089) );
  OR2_X1 U7468 ( .A1(n15242), .A2(n11099), .ZN(n7020) );
  OAI21_X2 U7469 ( .B1(n8796), .B2(n8897), .A(n15050), .ZN(n8784) );
  INV_X2 U7470 ( .A(n15369), .ZN(n15371) );
  NAND2_X1 U7471 ( .A1(n10896), .A2(n9544), .ZN(n14783) );
  NAND2_X1 U7472 ( .A1(n8350), .A2(n8349), .ZN(n15126) );
  NOR2_X1 U7473 ( .A1(n14524), .A2(n14523), .ZN(n14526) );
  OR2_X1 U7474 ( .A1(n7919), .A2(n7927), .ZN(n7929) );
  AND2_X1 U7475 ( .A1(n14782), .A2(n9540), .ZN(n10893) );
  NOR2_X1 U7476 ( .A1(n10826), .A2(n10508), .ZN(n12005) );
  INV_X1 U7477 ( .A(n10869), .ZN(n14800) );
  BUF_X4 U7478 ( .A(n8211), .Z(n8718) );
  NAND2_X1 U7479 ( .A1(n8065), .A2(n8064), .ZN(n8331) );
  INV_X2 U7480 ( .A(n8233), .ZN(n15021) );
  CLKBUF_X1 U7481 ( .A(n10304), .Z(n15018) );
  INV_X1 U7482 ( .A(n11037), .ZN(n15331) );
  NAND2_X1 U7484 ( .A1(n7276), .A2(n7275), .ZN(n9078) );
  NAND2_X2 U7485 ( .A1(n10810), .A2(n7130), .ZN(n8233) );
  XNOR2_X1 U7486 ( .A(n14519), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U7487 ( .A1(n8231), .A2(n8232), .ZN(n10433) );
  AND4_X1 U7488 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n11242)
         );
  INV_X2 U7489 ( .A(n9417), .ZN(n9519) );
  NAND2_X2 U7490 ( .A1(n9860), .A2(n9866), .ZN(n13729) );
  NAND2_X1 U7491 ( .A1(n6946), .A2(n6945), .ZN(n9027) );
  AND4_X1 U7492 ( .A1(n9003), .A2(n9002), .A3(n9001), .A4(n9000), .ZN(n9939)
         );
  NAND4_X1 U7493 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n12985)
         );
  AND2_X2 U7494 ( .A1(n12244), .A2(n12074), .ZN(n12227) );
  AND2_X1 U7495 ( .A1(n8003), .A2(n8026), .ZN(n8008) );
  AND3_X1 U7496 ( .A1(n7569), .A2(n7568), .A3(n7567), .ZN(n11411) );
  OR2_X1 U7497 ( .A1(n8155), .A2(n8154), .ZN(n8159) );
  BUF_X2 U7498 ( .A(n8894), .Z(n9847) );
  INV_X1 U7499 ( .A(n9469), .ZN(n9417) );
  INV_X4 U7500 ( .A(n8658), .ZN(n8956) );
  CLKBUF_X3 U7501 ( .A(n8226), .Z(n9780) );
  AND4_X1 U7502 ( .A1(n8184), .A2(n8183), .A3(n8185), .A4(n8182), .ZN(n8842)
         );
  AND2_X1 U7503 ( .A1(n14970), .A2(n14969), .ZN(n6923) );
  CLKBUF_X2 U7504 ( .A(n9072), .Z(n9477) );
  AND2_X1 U7505 ( .A1(n8162), .A2(n8163), .ZN(n8894) );
  INV_X1 U7506 ( .A(n10692), .ZN(n10816) );
  INV_X1 U7507 ( .A(n8693), .ZN(n8226) );
  NAND2_X1 U7508 ( .A1(n14449), .A2(n14452), .ZN(n9072) );
  AND2_X1 U7509 ( .A1(n6915), .A2(n8059), .ZN(n6912) );
  MUX2_X1 U7510 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8161), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8162) );
  NAND2_X1 U7511 ( .A1(n8048), .A2(n8047), .ZN(n8225) );
  AND2_X1 U7512 ( .A1(n7504), .A2(n12764), .ZN(n7505) );
  NOR2_X1 U7513 ( .A1(n7684), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7700) );
  INV_X1 U7514 ( .A(n8179), .ZN(n11823) );
  XNOR2_X1 U7515 ( .A(n8166), .B(n8165), .ZN(n8783) );
  NAND2_X1 U7516 ( .A1(n8982), .A2(n14442), .ZN(n14452) );
  OR2_X1 U7517 ( .A1(n7503), .A2(n8002), .ZN(n7500) );
  XNOR2_X1 U7518 ( .A(n8177), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8181) );
  OR2_X1 U7519 ( .A1(n8164), .A2(n8333), .ZN(n8166) );
  NAND2_X1 U7520 ( .A1(n7491), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7493) );
  XNOR2_X1 U7521 ( .A(n8978), .B(n8977), .ZN(n8983) );
  MUX2_X1 U7522 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8980), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n8982) );
  OR2_X1 U7523 ( .A1(n7139), .A2(n8333), .ZN(n6813) );
  NAND2_X1 U7524 ( .A1(n13372), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8177) );
  OR2_X1 U7525 ( .A1(n8981), .A2(n14441), .ZN(n8978) );
  OAI21_X1 U7526 ( .B1(n9586), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9583) );
  AND2_X1 U7528 ( .A1(n8976), .A2(n6634), .ZN(n7262) );
  NAND2_X2 U7529 ( .A1(n9960), .A2(P1_U3086), .ZN(n14458) );
  INV_X4 U7530 ( .A(n8043), .ZN(n9960) );
  NAND2_X1 U7531 ( .A1(n7184), .A2(n7182), .ZN(n14511) );
  INV_X1 U7532 ( .A(n8975), .ZN(n8976) );
  NOR2_X1 U7533 ( .A1(n7051), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7050) );
  AND2_X1 U7534 ( .A1(n7185), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14506) );
  AND2_X1 U7535 ( .A1(n8141), .A2(n6809), .ZN(n6807) );
  AND2_X1 U7536 ( .A1(n6811), .A2(n8229), .ZN(n6808) );
  XNOR2_X1 U7537 ( .A(n7526), .B(n7525), .ZN(n10595) );
  AND4_X1 U7538 ( .A1(n7486), .A2(n7485), .A3(n7484), .A4(n7715), .ZN(n7487)
         );
  AND3_X1 U7539 ( .A1(n8973), .A2(n8972), .A3(n8971), .ZN(n9566) );
  AND3_X1 U7540 ( .A1(n7480), .A2(n7481), .A3(n7479), .ZN(n7628) );
  NOR2_X1 U7541 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7486) );
  NOR2_X1 U7542 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_16__SCAN_IN), .ZN(
        n7485) );
  INV_X1 U7543 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7484) );
  INV_X1 U7544 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8333) );
  INV_X1 U7545 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9232) );
  INV_X1 U7546 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9252) );
  INV_X1 U7547 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14610) );
  NOR3_X1 U7548 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .A3(
        P1_IR_REG_15__SCAN_IN), .ZN(n8969) );
  INV_X2 U7549 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7550 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n13570) );
  INV_X4 U7551 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7552 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8136) );
  INV_X1 U7553 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8488) );
  INV_X1 U7554 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9133) );
  NOR2_X1 U7555 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n8146) );
  INV_X1 U7556 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9180) );
  INV_X1 U7557 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n14043) );
  INV_X1 U7558 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7495) );
  INV_X1 U7559 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n8347) );
  AND2_X1 U7560 ( .A1(n8174), .A2(n6811), .ZN(n8205) );
  AND4_X2 U7561 ( .A1(n6808), .A2(n6807), .A3(n8174), .A4(n6810), .ZN(n8332)
         );
  OAI222_X1 U7562 ( .A1(n10100), .A2(P1_U3086), .B1(n14458), .B2(n9990), .C1(
        n9989), .C2(n14455), .ZN(P1_U3354) );
  OAI222_X1 U7563 ( .A1(n13395), .A2(n9982), .B1(n13393), .B2(n9990), .C1(
        P2_U3088), .C2(n14947), .ZN(P2_U3326) );
  NOR2_X2 U7564 ( .A1(n13200), .A2(n13318), .ZN(n13192) );
  INV_X2 U7565 ( .A(n9072), .ZN(n8998) );
  XNOR2_X1 U7566 ( .A(n8211), .B(n10331), .ZN(n8218) );
  NAND4_X1 U7567 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n12984)
         );
  AND2_X1 U7568 ( .A1(n7506), .A2(n7505), .ZN(n7530) );
  OAI21_X2 U7569 ( .B1(n13861), .B2(n6741), .A(n6739), .ZN(n13700) );
  NAND2_X1 U7570 ( .A1(n8888), .A2(n9845), .ZN(n6553) );
  XNOR2_X1 U7571 ( .A(n10417), .B(n10470), .ZN(n10408) );
  NAND2_X2 U7572 ( .A1(n8254), .A2(n8253), .ZN(n10417) );
  AND2_X1 U7573 ( .A1(n7924), .A2(n7923), .ZN(n11404) );
  NOR2_X2 U7574 ( .A1(n14196), .A2(n14356), .ZN(n14181) );
  NOR2_X2 U7575 ( .A1(n8230), .A2(n8249), .ZN(n12992) );
  INV_X1 U7576 ( .A(n8783), .ZN(n6554) );
  INV_X1 U7577 ( .A(n6554), .ZN(n6555) );
  INV_X1 U7578 ( .A(n6554), .ZN(n6556) );
  OR2_X1 U7579 ( .A1(n10299), .A2(n10167), .ZN(n10328) );
  XNOR2_X1 U7580 ( .A(n6553), .B(n10299), .ZN(n8197) );
  OR2_X1 U7581 ( .A1(n7826), .A2(n10593), .ZN(n7518) );
  NAND2_X2 U7582 ( .A1(n12535), .A2(n7963), .ZN(n12519) );
  NOR2_X2 U7583 ( .A1(n14792), .A2(n14788), .ZN(n14793) );
  NAND2_X1 U7584 ( .A1(n10940), .A2(n6957), .ZN(n14792) );
  OR2_X1 U7585 ( .A1(n14381), .A2(n14252), .ZN(n14073) );
  AND2_X1 U7586 ( .A1(n6882), .A2(n6881), .ZN(n6880) );
  NOR2_X1 U7587 ( .A1(n7162), .A2(n6621), .ZN(n7161) );
  INV_X1 U7588 ( .A(n8875), .ZN(n7162) );
  OAI22_X1 U7589 ( .A1(n13116), .A2(n6984), .B1(n6985), .B2(n9807), .ZN(n13081) );
  NAND2_X1 U7590 ( .A1(n13105), .A2(n13090), .ZN(n6984) );
  NAND2_X1 U7591 ( .A1(n9008), .A2(n6610), .ZN(n7231) );
  NAND2_X1 U7592 ( .A1(n11621), .A2(n6602), .ZN(n6940) );
  INV_X1 U7593 ( .A(n14083), .ZN(n6941) );
  OAI211_X1 U7594 ( .C1(n12702), .C2(n12077), .A(n12076), .B(n15345), .ZN(
        n12083) );
  NAND2_X1 U7595 ( .A1(n12145), .A2(n6702), .ZN(n6701) );
  AND2_X1 U7596 ( .A1(n12615), .A2(n6703), .ZN(n6702) );
  NAND2_X1 U7597 ( .A1(n9348), .A2(n6569), .ZN(n7280) );
  INV_X1 U7598 ( .A(n9349), .ZN(n7281) );
  OR2_X1 U7599 ( .A1(n13255), .A2(n6995), .ZN(n6993) );
  OR2_X1 U7600 ( .A1(n7339), .A2(n7338), .ZN(n7337) );
  NAND2_X1 U7601 ( .A1(n11269), .A2(n6878), .ZN(n6877) );
  AND2_X1 U7602 ( .A1(n11392), .A2(n11268), .ZN(n6878) );
  NAND2_X1 U7603 ( .A1(n12407), .A2(n6782), .ZN(n6781) );
  INV_X1 U7604 ( .A(n12417), .ZN(n6782) );
  OR2_X1 U7605 ( .A1(n12438), .A2(n12416), .ZN(n12198) );
  INV_X1 U7606 ( .A(n7048), .ZN(n7043) );
  NAND2_X1 U7607 ( .A1(n6550), .A2(n9981), .ZN(n7546) );
  INV_X1 U7608 ( .A(n7095), .ZN(n7093) );
  AOI21_X1 U7609 ( .B1(n7095), .B2(n6670), .A(n6677), .ZN(n7092) );
  NAND2_X1 U7610 ( .A1(n7081), .A2(n7080), .ZN(n7477) );
  AOI21_X1 U7611 ( .B1(n7083), .B2(n7085), .A(n6676), .ZN(n7080) );
  NAND2_X1 U7612 ( .A1(n7784), .A2(n7083), .ZN(n7081) );
  NAND2_X1 U7613 ( .A1(n6786), .A2(n6785), .ZN(n7460) );
  AOI21_X1 U7614 ( .B1(n6787), .B2(n7072), .A(n6671), .ZN(n6785) );
  AND2_X1 U7615 ( .A1(n7027), .A2(n13570), .ZN(n7026) );
  INV_X1 U7616 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7027) );
  AND2_X1 U7617 ( .A1(n6558), .A2(n8938), .ZN(n6983) );
  NOR2_X1 U7618 ( .A1(n9898), .A2(n9897), .ZN(n6735) );
  INV_X1 U7619 ( .A(n14452), .ZN(n8984) );
  AOI21_X1 U7620 ( .B1(n14192), .B2(n6950), .A(n6947), .ZN(n7230) );
  INV_X1 U7621 ( .A(n14193), .ZN(n6948) );
  NAND2_X1 U7622 ( .A1(n14175), .A2(n6582), .ZN(n6834) );
  NAND2_X1 U7623 ( .A1(n7215), .A2(n7214), .ZN(n14250) );
  NOR2_X1 U7624 ( .A1(n7416), .A2(n14071), .ZN(n7214) );
  NAND2_X1 U7625 ( .A1(n9008), .A2(n9367), .ZN(n9184) );
  NAND2_X1 U7626 ( .A1(n9528), .A2(n10687), .ZN(n9862) );
  NOR2_X1 U7627 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7265) );
  AND2_X1 U7628 ( .A1(n6828), .A2(n7317), .ZN(n6827) );
  AOI21_X1 U7629 ( .B1(n7319), .B2(n7322), .A(n7318), .ZN(n7317) );
  INV_X1 U7630 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8964) );
  XNOR2_X1 U7631 ( .A(P1_ADDR_REG_1__SCAN_IN), .B(P3_ADDR_REG_1__SCAN_IN), 
        .ZN(n14505) );
  XNOR2_X1 U7632 ( .A(n14468), .B(P3_ADDR_REG_5__SCAN_IN), .ZN(n14519) );
  AND2_X1 U7633 ( .A1(n6871), .A2(n11803), .ZN(n6870) );
  NAND2_X1 U7634 ( .A1(n7444), .A2(n6872), .ZN(n6871) );
  INV_X1 U7635 ( .A(n11786), .ZN(n6872) );
  INV_X1 U7636 ( .A(n7444), .ZN(n6873) );
  NAND2_X1 U7637 ( .A1(n10819), .A2(n15341), .ZN(n10953) );
  XNOR2_X1 U7638 ( .A(n12706), .B(n11901), .ZN(n10819) );
  NAND2_X1 U7639 ( .A1(n11968), .A2(n11922), .ZN(n12071) );
  NAND2_X1 U7640 ( .A1(n12483), .A2(n12464), .ZN(n12467) );
  INV_X1 U7641 ( .A(n12033), .ZN(n7800) );
  INV_X1 U7642 ( .A(n12035), .ZN(n12027) );
  INV_X1 U7643 ( .A(n7086), .ZN(n12031) );
  OAI21_X1 U7644 ( .B1(n12021), .B2(n7088), .A(n7087), .ZN(n7086) );
  NAND2_X1 U7645 ( .A1(n14450), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7087) );
  INV_X1 U7646 ( .A(n12022), .ZN(n7088) );
  AND2_X2 U7647 ( .A1(n7992), .A2(n7993), .ZN(n7991) );
  NAND2_X1 U7648 ( .A1(n6771), .A2(n7475), .ZN(n7784) );
  NAND2_X1 U7649 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n13502), .ZN(n7475) );
  NAND2_X1 U7650 ( .A1(n7758), .A2(n7757), .ZN(n6771) );
  INV_X1 U7651 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7479) );
  NAND2_X1 U7652 ( .A1(n8181), .A2(n8179), .ZN(n8212) );
  XNOR2_X1 U7653 ( .A(n13038), .B(n13037), .ZN(n13025) );
  NOR2_X1 U7654 ( .A1(n13081), .A2(n8945), .ZN(n13064) );
  AND2_X1 U7655 ( .A1(n13280), .A2(n8944), .ZN(n8945) );
  AOI21_X1 U7656 ( .B1(n13105), .B2(n6987), .A(n6986), .ZN(n6985) );
  INV_X1 U7657 ( .A(n8941), .ZN(n6987) );
  INV_X1 U7658 ( .A(n8943), .ZN(n6986) );
  NAND2_X1 U7659 ( .A1(n13109), .A2(n8874), .ZN(n8876) );
  AND2_X1 U7660 ( .A1(n8941), .A2(n8940), .ZN(n13118) );
  NAND2_X1 U7661 ( .A1(n8871), .A2(n7166), .ZN(n7165) );
  NOR2_X1 U7662 ( .A1(n6616), .A2(n7167), .ZN(n7166) );
  INV_X1 U7663 ( .A(n8870), .ZN(n7167) );
  NAND2_X1 U7664 ( .A1(n6558), .A2(n6588), .ZN(n6982) );
  AOI21_X1 U7665 ( .B1(n7006), .B2(n7004), .A(n6609), .ZN(n7003) );
  INV_X1 U7666 ( .A(n7006), .ZN(n7005) );
  INV_X1 U7667 ( .A(n8934), .ZN(n7004) );
  AOI21_X1 U7668 ( .B1(n7154), .B2(n7157), .A(n7153), .ZN(n7152) );
  NAND2_X1 U7669 ( .A1(n6805), .A2(n6603), .ZN(n8862) );
  INV_X1 U7670 ( .A(n11368), .ZN(n6805) );
  INV_X1 U7671 ( .A(n9815), .ZN(n10655) );
  INV_X1 U7672 ( .A(n8188), .ZN(n7136) );
  AND2_X1 U7673 ( .A1(n9868), .A2(n9867), .ZN(n10234) );
  OR2_X1 U7674 ( .A1(n9939), .A2(n13729), .ZN(n9868) );
  NAND2_X1 U7675 ( .A1(n13874), .A2(n13875), .ZN(n13873) );
  AOI21_X1 U7676 ( .B1(n11502), .B2(n11501), .A(n11500), .ZN(n11503) );
  AND2_X1 U7677 ( .A1(n11499), .A2(n11498), .ZN(n11500) );
  NAND2_X1 U7678 ( .A1(n8985), .A2(n14452), .ZN(n9071) );
  NOR2_X1 U7679 ( .A1(n9555), .A2(n7252), .ZN(n7248) );
  AOI21_X1 U7680 ( .B1(n7258), .B2(n14262), .A(n7257), .ZN(n7256) );
  INV_X1 U7681 ( .A(n14073), .ZN(n7257) );
  NAND2_X1 U7682 ( .A1(n14307), .A2(n14409), .ZN(n14306) );
  NOR2_X1 U7683 ( .A1(n14305), .A2(n6939), .ZN(n6938) );
  INV_X1 U7684 ( .A(n14087), .ZN(n6939) );
  NAND2_X1 U7685 ( .A1(n14810), .A2(n10874), .ZN(n10871) );
  INV_X1 U7686 ( .A(n14766), .ZN(n14802) );
  INV_X1 U7687 ( .A(n14261), .ZN(n14386) );
  AND3_X2 U7688 ( .A1(n9313), .A2(n8976), .A3(n7264), .ZN(n8995) );
  INV_X1 U7689 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7264) );
  NAND2_X1 U7690 ( .A1(n6568), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U7691 ( .A1(n6761), .A2(n6567), .ZN(n14555) );
  OR2_X1 U7692 ( .A1(n14717), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n7186) );
  OAI21_X1 U7693 ( .B1(n14603), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n6564), .ZN(
        n7174) );
  NAND2_X1 U7694 ( .A1(n7118), .A2(n7117), .ZN(n7116) );
  INV_X1 U7695 ( .A(n8806), .ZN(n7117) );
  NAND2_X1 U7696 ( .A1(n13274), .A2(n8784), .ZN(n7118) );
  NAND2_X1 U7697 ( .A1(n9322), .A2(n13928), .ZN(n6946) );
  OAI22_X1 U7698 ( .A1(n7384), .A2(n7385), .B1(n9611), .B2(n7383), .ZN(n9615)
         );
  INV_X1 U7699 ( .A(n9610), .ZN(n7383) );
  NOR2_X1 U7700 ( .A1(n9612), .A2(n9610), .ZN(n7384) );
  NAND2_X1 U7701 ( .A1(n7412), .A2(n9661), .ZN(n7411) );
  INV_X1 U7702 ( .A(n9671), .ZN(n7403) );
  AOI21_X1 U7703 ( .B1(n6627), .B2(n9693), .A(n9706), .ZN(n7388) );
  AOI21_X1 U7704 ( .B1(n12158), .B2(n12157), .A(n12156), .ZN(n12165) );
  AND2_X1 U7705 ( .A1(n6904), .A2(n9370), .ZN(n6903) );
  OAI21_X1 U7706 ( .B1(n7281), .B2(n7280), .A(n6622), .ZN(n6907) );
  INV_X1 U7707 ( .A(n6905), .ZN(n6902) );
  NAND2_X1 U7708 ( .A1(n9748), .A2(n9750), .ZN(n7394) );
  NAND2_X1 U7709 ( .A1(n9395), .A2(n9394), .ZN(n6900) );
  INV_X1 U7710 ( .A(n9414), .ZN(n7284) );
  NAND2_X1 U7711 ( .A1(n6705), .A2(n6704), .ZN(n12193) );
  AND2_X1 U7712 ( .A1(n12474), .A2(n12192), .ZN(n6704) );
  NAND2_X1 U7713 ( .A1(n12186), .A2(n6706), .ZN(n6705) );
  INV_X1 U7714 ( .A(n8102), .ZN(n6833) );
  NAND2_X1 U7715 ( .A1(n10825), .A2(n15354), .ZN(n12085) );
  NAND2_X1 U7716 ( .A1(n7310), .A2(n6682), .ZN(n9794) );
  NAND2_X1 U7717 ( .A1(n13052), .A2(n9779), .ZN(n7310) );
  INV_X1 U7718 ( .A(n12959), .ZN(n7309) );
  NAND2_X1 U7719 ( .A1(n7307), .A2(n9832), .ZN(n9797) );
  OAI22_X1 U7720 ( .A1(n9795), .A2(n9794), .B1(n9790), .B2(n9791), .ZN(n7307)
         );
  INV_X1 U7721 ( .A(n8908), .ZN(n6995) );
  AND3_X1 U7722 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .A3(
        P2_IR_REG_27__SCAN_IN), .ZN(n8149) );
  INV_X1 U7723 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8141) );
  INV_X1 U7724 ( .A(n8689), .ZN(n7335) );
  AOI21_X1 U7725 ( .B1(n6821), .B2(n6824), .A(n6819), .ZN(n6818) );
  INV_X1 U7726 ( .A(n7437), .ZN(n6819) );
  AND2_X1 U7727 ( .A1(n8963), .A2(n9054), .ZN(n7266) );
  NAND2_X1 U7728 ( .A1(n14465), .A2(n7177), .ZN(n14466) );
  NAND2_X1 U7729 ( .A1(n14516), .A2(n14463), .ZN(n7177) );
  AND3_X1 U7730 ( .A1(n7586), .A2(n7585), .A3(n7584), .ZN(n11386) );
  NAND2_X1 U7731 ( .A1(n11061), .A2(n11060), .ZN(n11062) );
  NAND2_X1 U7732 ( .A1(n15198), .A2(n6599), .ZN(n11126) );
  NAND2_X1 U7733 ( .A1(n15271), .A2(n6800), .ZN(n11136) );
  OR2_X1 U7734 ( .A1(n11134), .A2(n11133), .ZN(n6800) );
  OR2_X1 U7735 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  NOR2_X1 U7736 ( .A1(n12171), .A2(n7046), .ZN(n7045) );
  INV_X1 U7737 ( .A(n12173), .ZN(n7046) );
  NOR2_X1 U7738 ( .A1(n7033), .A2(n11564), .ZN(n7029) );
  INV_X1 U7739 ( .A(n12113), .ZN(n7033) );
  INV_X1 U7740 ( .A(n12116), .ZN(n7031) );
  AND3_X1 U7741 ( .A1(n7618), .A2(n7617), .A3(n7616), .ZN(n7935) );
  NAND2_X1 U7742 ( .A1(n12085), .A2(n12079), .ZN(n15342) );
  INV_X1 U7743 ( .A(n7456), .ZN(n7069) );
  INV_X1 U7744 ( .A(n7458), .ZN(n7073) );
  NOR2_X1 U7745 ( .A1(n7078), .A2(n7075), .ZN(n7074) );
  INV_X1 U7746 ( .A(n7577), .ZN(n7078) );
  INV_X1 U7747 ( .A(n7563), .ZN(n7075) );
  INV_X1 U7748 ( .A(n7453), .ZN(n7077) );
  NAND2_X1 U7749 ( .A1(n8937), .A2(n8936), .ZN(n13165) );
  NAND2_X1 U7750 ( .A1(n6658), .A2(n8927), .ZN(n7000) );
  NOR2_X1 U7751 ( .A1(n8930), .A2(n7002), .ZN(n7001) );
  INV_X1 U7752 ( .A(n8927), .ZN(n7002) );
  INV_X1 U7753 ( .A(n8905), .ZN(n6974) );
  INV_X1 U7754 ( .A(n8904), .ZN(n6972) );
  OAI21_X1 U7755 ( .B1(n10411), .B2(n6974), .A(n10644), .ZN(n6968) );
  OR2_X1 U7756 ( .A1(n12986), .A2(n10331), .ZN(n8903) );
  AND2_X1 U7757 ( .A1(n6555), .A2(n11057), .ZN(n7130) );
  NOR2_X1 U7758 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n8147) );
  NOR2_X1 U7759 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .ZN(
        n8148) );
  INV_X1 U7760 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n8143) );
  NOR2_X1 U7761 ( .A1(n8508), .A2(n8140), .ZN(n7135) );
  INV_X1 U7762 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U7763 ( .A1(n6688), .A2(n6687), .ZN(n8167) );
  BUF_X1 U7764 ( .A(n8533), .Z(n8534) );
  AND2_X1 U7765 ( .A1(n8427), .A2(n8426), .ZN(n8448) );
  NOR2_X1 U7766 ( .A1(n7347), .A2(n7422), .ZN(n7346) );
  INV_X1 U7767 ( .A(n11180), .ZN(n7347) );
  INV_X1 U7768 ( .A(n14328), .ZN(n14044) );
  NOR2_X1 U7769 ( .A1(n14236), .A2(n14096), .ZN(n6934) );
  NAND2_X1 U7770 ( .A1(n6932), .A2(n14095), .ZN(n6931) );
  INV_X1 U7771 ( .A(n14096), .ZN(n6932) );
  INV_X1 U7772 ( .A(n14236), .ZN(n7260) );
  INV_X1 U7773 ( .A(n7236), .ZN(n7235) );
  OAI21_X1 U7774 ( .B1(n11014), .B2(n7237), .A(n11163), .ZN(n7236) );
  INV_X1 U7775 ( .A(n11016), .ZN(n7237) );
  NAND2_X1 U7776 ( .A1(n9028), .A2(n9027), .ZN(n9536) );
  NAND2_X1 U7777 ( .A1(n9939), .A2(n10320), .ZN(n9538) );
  NAND2_X1 U7778 ( .A1(n14149), .A2(n14080), .ZN(n7249) );
  OR2_X1 U7779 ( .A1(n6720), .A2(n9864), .ZN(n9951) );
  AND2_X1 U7780 ( .A1(n9943), .A2(n10320), .ZN(n10864) );
  AND2_X1 U7781 ( .A1(n9566), .A2(n9568), .ZN(n6752) );
  INV_X1 U7782 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9568) );
  INV_X1 U7783 ( .A(n8650), .ZN(n8127) );
  NAND2_X1 U7784 ( .A1(n6916), .A2(n7323), .ZN(n8551) );
  NAND2_X1 U7785 ( .A1(n8507), .A2(n7324), .ZN(n6916) );
  NAND2_X1 U7786 ( .A1(n6830), .A2(n8102), .ZN(n8507) );
  NAND2_X1 U7787 ( .A1(n7314), .A2(n6579), .ZN(n6830) );
  AOI21_X1 U7788 ( .B1(n7329), .B2(n7331), .A(n6620), .ZN(n7327) );
  XNOR2_X1 U7789 ( .A(n8060), .B(SI_6_), .ZN(n8290) );
  NAND2_X1 U7790 ( .A1(n8057), .A2(n8056), .ZN(n8265) );
  XNOR2_X1 U7791 ( .A(n6816), .B(SI_5_), .ZN(n8266) );
  XNOR2_X1 U7792 ( .A(n8051), .B(n6909), .ZN(n8050) );
  INV_X1 U7793 ( .A(SI_3_), .ZN(n6909) );
  AND2_X2 U7794 ( .A1(n7300), .A2(n7299), .ZN(n8043) );
  INV_X1 U7795 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7496) );
  NAND2_X1 U7796 ( .A1(n7183), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7182) );
  NAND2_X1 U7797 ( .A1(n14505), .A2(n14506), .ZN(n7184) );
  XNOR2_X1 U7798 ( .A(n14466), .B(P3_ADDR_REG_4__SCAN_IN), .ZN(n14503) );
  OAI21_X1 U7799 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n14477), .A(n14476), .ZN(
        n14537) );
  NAND2_X1 U7800 ( .A1(n11963), .A2(n11888), .ZN(n11897) );
  AND2_X1 U7801 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  AND2_X1 U7802 ( .A1(n11269), .A2(n11268), .ZN(n11393) );
  INV_X1 U7803 ( .A(n11573), .ZN(n6879) );
  AND2_X1 U7804 ( .A1(n6592), .A2(n11574), .ZN(n6876) );
  AOI21_X1 U7805 ( .B1(n6870), .B2(n6873), .A(n6661), .ZN(n6869) );
  OR2_X1 U7806 ( .A1(n14626), .A2(n12037), .ZN(n12221) );
  AND2_X1 U7807 ( .A1(n12040), .A2(n7064), .ZN(n7063) );
  NAND2_X1 U7808 ( .A1(n7057), .A2(n7060), .ZN(n7055) );
  NAND3_X1 U7809 ( .A1(n8028), .A2(n8027), .A3(n8026), .ZN(n10513) );
  OAI21_X1 U7810 ( .B1(n6546), .B2(n10579), .A(n7433), .ZN(n6799) );
  INV_X1 U7811 ( .A(n10594), .ZN(n10596) );
  OAI21_X1 U7812 ( .B1(n6552), .B2(P3_REG2_REG_2__SCAN_IN), .A(n7009), .ZN(
        n10585) );
  NAND2_X1 U7813 ( .A1(n11119), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7009) );
  NAND2_X1 U7814 ( .A1(n10585), .A2(n10584), .ZN(n11061) );
  XNOR2_X1 U7815 ( .A(n11062), .B(n15180), .ZN(n15166) );
  NAND2_X1 U7816 ( .A1(n15200), .A2(n15199), .ZN(n15198) );
  XNOR2_X1 U7817 ( .A(n11126), .B(n11127), .ZN(n15218) );
  OR2_X1 U7818 ( .A1(n15187), .A2(n6587), .ZN(n7018) );
  NOR2_X1 U7819 ( .A1(n15223), .A2(n7021), .ZN(n11068) );
  NOR2_X1 U7820 ( .A1(n11129), .A2(n11093), .ZN(n7021) );
  INV_X1 U7821 ( .A(n11135), .ZN(n15289) );
  NAND2_X1 U7822 ( .A1(n11072), .A2(n15289), .ZN(n11071) );
  XNOR2_X1 U7823 ( .A(n11136), .B(n11135), .ZN(n15295) );
  NAND2_X1 U7824 ( .A1(n15295), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n15294) );
  OAI21_X1 U7825 ( .B1(n15284), .B2(n15283), .A(n15282), .ZN(n15281) );
  NAND2_X1 U7826 ( .A1(n12313), .A2(n12314), .ZN(n12330) );
  NAND2_X1 U7827 ( .A1(n12330), .A2(n6804), .ZN(n12331) );
  NAND2_X1 U7828 ( .A1(n14590), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6804) );
  NOR2_X1 U7829 ( .A1(n6695), .A2(n6694), .ZN(n6693) );
  INV_X1 U7830 ( .A(n12352), .ZN(n6695) );
  INV_X1 U7831 ( .A(n6692), .ZN(n12379) );
  AND2_X1 U7832 ( .A1(n7899), .A2(n11905), .ZN(n14614) );
  OAI21_X1 U7833 ( .B1(n7979), .B2(n6562), .A(n6774), .ZN(n6773) );
  NAND2_X1 U7834 ( .A1(n12217), .A2(n6781), .ZN(n6780) );
  NOR2_X1 U7835 ( .A1(n12212), .A2(n7062), .ZN(n7061) );
  NAND2_X1 U7836 ( .A1(n7870), .A2(n7869), .ZN(n12438) );
  AND2_X1 U7837 ( .A1(n12067), .A2(n12066), .ZN(n12451) );
  INV_X1 U7838 ( .A(n7039), .ZN(n7038) );
  OAI21_X1 U7839 ( .B1(n12474), .B2(n7040), .A(n12451), .ZN(n7039) );
  INV_X1 U7840 ( .A(n12071), .ZN(n7040) );
  AND2_X1 U7841 ( .A1(n7854), .A2(n12068), .ZN(n7419) );
  NAND2_X1 U7842 ( .A1(n7419), .A2(n12474), .ZN(n12473) );
  NAND2_X1 U7843 ( .A1(n12463), .A2(n12491), .ZN(n12483) );
  NOR2_X1 U7844 ( .A1(n7809), .A2(n7049), .ZN(n7048) );
  INV_X1 U7845 ( .A(n12161), .ZN(n7049) );
  AND2_X1 U7846 ( .A1(n12564), .A2(n12563), .ZN(n12614) );
  AND4_X1 U7847 ( .A1(n7661), .A2(n7660), .A3(n7659), .A4(n7658), .ZN(n11727)
         );
  AND3_X1 U7848 ( .A1(n7650), .A2(n7649), .A3(n7648), .ZN(n12120) );
  NAND2_X1 U7849 ( .A1(n11463), .A2(n12108), .ZN(n7034) );
  AND2_X1 U7850 ( .A1(n12116), .A2(n12115), .ZN(n12113) );
  OR2_X1 U7851 ( .A1(n7558), .A2(n7516), .ZN(n7517) );
  AND2_X1 U7852 ( .A1(n7846), .A2(n7845), .ZN(n11844) );
  OR2_X1 U7853 ( .A1(n8829), .A2(n8024), .ZN(n10517) );
  AND2_X1 U7854 ( .A1(n10513), .A2(n10039), .ZN(n10574) );
  AOI21_X1 U7855 ( .B1(n8808), .B2(n8809), .A(n7089), .ZN(n12021) );
  AND2_X1 U7856 ( .A1(n11814), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n7089) );
  XNOR2_X1 U7857 ( .A(n7490), .B(n7498), .ZN(n7985) );
  OR2_X1 U7858 ( .A1(n7499), .A2(n8002), .ZN(n7490) );
  INV_X1 U7859 ( .A(n7050), .ZN(n6884) );
  NAND2_X1 U7860 ( .A1(n6790), .A2(n6788), .ZN(n7833) );
  OAI21_X1 U7861 ( .B1(n6789), .B2(n7820), .A(n6674), .ZN(n6788) );
  NOR2_X1 U7862 ( .A1(n6792), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n6791) );
  XNOR2_X1 U7863 ( .A(n7477), .B(n10681), .ZN(n7810) );
  XNOR2_X1 U7864 ( .A(n7799), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12375) );
  NAND2_X1 U7865 ( .A1(n7474), .A2(n7473), .ZN(n7758) );
  NAND2_X1 U7866 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n7472), .ZN(n7473) );
  OR2_X1 U7867 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n10386), .ZN(n7467) );
  NAND2_X1 U7868 ( .A1(n6561), .A2(n7102), .ZN(n7101) );
  INV_X1 U7869 ( .A(n7107), .ZN(n7102) );
  AND2_X1 U7870 ( .A1(n6577), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U7871 ( .A1(n7103), .A2(n7104), .ZN(n7465) );
  NAND2_X1 U7872 ( .A1(n7681), .A2(n7107), .ZN(n7103) );
  AND2_X1 U7873 ( .A1(n7536), .A2(n7483), .ZN(n7025) );
  OR2_X1 U7874 ( .A1(n7646), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U7875 ( .A1(n7457), .A2(n7456), .ZN(n7632) );
  XNOR2_X1 U7876 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7631) );
  XNOR2_X1 U7877 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7577) );
  OR2_X1 U7878 ( .A1(n7583), .A2(n7582), .ZN(n15214) );
  XNOR2_X1 U7879 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7563) );
  NAND2_X1 U7880 ( .A1(n7452), .A2(n7451), .ZN(n7564) );
  AND2_X2 U7881 ( .A1(n6854), .A2(n7526), .ZN(n7536) );
  INV_X1 U7882 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6854) );
  INV_X1 U7883 ( .A(n12965), .ZN(n12852) );
  OR2_X1 U7884 ( .A1(n8495), .A2(n12862), .ZN(n8516) );
  INV_X1 U7885 ( .A(n12913), .ZN(n12885) );
  NAND2_X1 U7886 ( .A1(n7129), .A2(n6600), .ZN(n10995) );
  AND2_X1 U7887 ( .A1(n8444), .A2(n8424), .ZN(n7127) );
  OR2_X1 U7888 ( .A1(n8412), .A2(n10550), .ZN(n8433) );
  INV_X1 U7889 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n8432) );
  NOR2_X1 U7890 ( .A1(n9835), .A2(n9774), .ZN(n9836) );
  AND2_X1 U7891 ( .A1(n13024), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6924) );
  NOR2_X1 U7892 ( .A1(n13025), .A2(n13026), .ZN(n13040) );
  XNOR2_X1 U7893 ( .A(n13270), .B(n9778), .ZN(n9806) );
  NAND2_X1 U7894 ( .A1(n8879), .A2(n8878), .ZN(n13063) );
  OR2_X1 U7895 ( .A1(n13274), .A2(n12961), .ZN(n8878) );
  NAND2_X1 U7896 ( .A1(n13116), .A2(n8941), .ZN(n13094) );
  AND2_X1 U7897 ( .A1(n13129), .A2(n6590), .ZN(n7164) );
  NAND2_X1 U7898 ( .A1(n6714), .A2(n6983), .ZN(n6978) );
  NAND2_X1 U7899 ( .A1(n6980), .A2(n6982), .ZN(n6979) );
  INV_X1 U7900 ( .A(n6983), .ZN(n6980) );
  INV_X1 U7901 ( .A(n6982), .ZN(n6981) );
  OR2_X1 U7902 ( .A1(n8580), .A2(n12892), .ZN(n8600) );
  OAI21_X1 U7903 ( .B1(n13205), .B2(n8931), .A(n8932), .ZN(n13188) );
  OR2_X1 U7904 ( .A1(n13188), .A2(n13189), .ZN(n13186) );
  NAND2_X1 U7905 ( .A1(n13216), .A2(n8867), .ZN(n13199) );
  NAND2_X1 U7906 ( .A1(n13218), .A2(n13217), .ZN(n13216) );
  NAND2_X1 U7907 ( .A1(n8926), .A2(n8925), .ZN(n13239) );
  AND2_X1 U7908 ( .A1(n7150), .A2(n8861), .ZN(n7149) );
  OR2_X1 U7909 ( .A1(n11475), .A2(n8863), .ZN(n7148) );
  OR2_X1 U7910 ( .A1(n8433), .A2(n8432), .ZN(n8453) );
  OAI21_X1 U7911 ( .B1(n11347), .B2(n8919), .A(n8920), .ZN(n11373) );
  INV_X1 U7912 ( .A(n11340), .ZN(n6806) );
  AOI21_X1 U7913 ( .B1(n6965), .B2(n6967), .A(n6606), .ZN(n6962) );
  NAND2_X1 U7914 ( .A1(n7133), .A2(n8856), .ZN(n15033) );
  AND2_X1 U7915 ( .A1(n6994), .A2(n8910), .ZN(n6990) );
  INV_X1 U7916 ( .A(n7170), .ZN(n7169) );
  OAI21_X1 U7917 ( .B1(n8851), .B2(n7171), .A(n10655), .ZN(n7170) );
  NAND2_X1 U7918 ( .A1(n13248), .A2(n13255), .ZN(n13247) );
  NAND2_X1 U7919 ( .A1(n8843), .A2(n8902), .ZN(n10303) );
  NAND2_X1 U7920 ( .A1(n10810), .A2(n11057), .ZN(n15043) );
  NAND2_X1 U7921 ( .A1(n8598), .A2(n8597), .ZN(n13312) );
  NAND2_X1 U7922 ( .A1(n8579), .A2(n8578), .ZN(n13318) );
  NAND2_X1 U7923 ( .A1(n7172), .A2(n8851), .ZN(n15104) );
  INV_X1 U7924 ( .A(n15146), .ZN(n15137) );
  NAND2_X1 U7925 ( .A1(n11057), .A2(n9774), .ZN(n15139) );
  AND2_X1 U7926 ( .A1(n9858), .A2(n10054), .ZN(n8802) );
  INV_X1 U7927 ( .A(n8145), .ZN(n7401) );
  OR2_X1 U7928 ( .A1(n8755), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8758) );
  NOR2_X1 U7929 ( .A1(n8778), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8752) );
  NAND2_X1 U7930 ( .A1(n8752), .A2(n8749), .ZN(n8755) );
  INV_X1 U7931 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8749) );
  INV_X1 U7932 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8154) );
  OR2_X1 U7933 ( .A1(n8251), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8268) );
  AND2_X1 U7934 ( .A1(n8205), .A2(n8229), .ZN(n8249) );
  INV_X1 U7935 ( .A(n6735), .ZN(n6731) );
  AND2_X1 U7936 ( .A1(n14657), .A2(n6581), .ZN(n6742) );
  NAND2_X1 U7937 ( .A1(n6750), .A2(n6749), .ZN(n6748) );
  INV_X1 U7938 ( .A(n13883), .ZN(n6750) );
  AOI21_X1 U7939 ( .B1(n7372), .B2(n7374), .A(n6631), .ZN(n7371) );
  AND2_X1 U7940 ( .A1(n13797), .A2(n7373), .ZN(n7372) );
  OR2_X1 U7941 ( .A1(n13890), .A2(n7374), .ZN(n7373) );
  NAND2_X1 U7942 ( .A1(n11178), .A2(n11177), .ZN(n7348) );
  INV_X1 U7943 ( .A(n13752), .ZN(n7354) );
  AND2_X1 U7944 ( .A1(n13846), .A2(n7353), .ZN(n7352) );
  OR2_X1 U7945 ( .A1(n7354), .A2(n13780), .ZN(n7353) );
  NAND2_X1 U7946 ( .A1(n6663), .A2(n7361), .ZN(n13827) );
  NAND2_X1 U7947 ( .A1(n7376), .A2(n6736), .ZN(n6732) );
  NOR2_X1 U7948 ( .A1(n7345), .A2(n6735), .ZN(n6733) );
  INV_X1 U7949 ( .A(n7346), .ZN(n7345) );
  INV_X1 U7950 ( .A(n10929), .ZN(n6738) );
  NAND2_X1 U7951 ( .A1(n7346), .A2(n7344), .ZN(n7343) );
  INV_X1 U7952 ( .A(n11177), .ZN(n7344) );
  AND2_X1 U7953 ( .A1(n11211), .A2(n11208), .ZN(n11209) );
  NAND2_X1 U7954 ( .A1(n7348), .A2(n7346), .ZN(n11210) );
  NOR2_X1 U7955 ( .A1(n10233), .A2(n10234), .ZN(n10232) );
  INV_X1 U7956 ( .A(n7359), .ZN(n7358) );
  OAI21_X1 U7957 ( .B1(n13711), .B2(n7360), .A(n6672), .ZN(n7359) );
  INV_X1 U7958 ( .A(n13837), .ZN(n7360) );
  OR2_X1 U7959 ( .A1(n9890), .A2(n7377), .ZN(n7376) );
  INV_X1 U7960 ( .A(n7378), .ZN(n7377) );
  NAND2_X1 U7961 ( .A1(n7380), .A2(n7378), .ZN(n7375) );
  NOR2_X1 U7962 ( .A1(n7379), .A2(n7381), .ZN(n7380) );
  AOI21_X1 U7963 ( .B1(n6742), .B2(n6740), .A(n13698), .ZN(n6739) );
  INV_X1 U7964 ( .A(n6742), .ZN(n6741) );
  INV_X1 U7965 ( .A(n13862), .ZN(n6740) );
  INV_X1 U7966 ( .A(n9861), .ZN(n9860) );
  INV_X1 U7967 ( .A(n9503), .ZN(n7278) );
  OR2_X1 U7968 ( .A1(n9468), .A2(n9483), .ZN(n6894) );
  INV_X1 U7969 ( .A(n9423), .ZN(n9374) );
  OR2_X1 U7970 ( .A1(n13996), .A2(n6842), .ZN(n6841) );
  AND2_X1 U7971 ( .A1(n14003), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6842) );
  AND2_X1 U7972 ( .A1(n6841), .A2(n6840), .ZN(n14011) );
  INV_X1 U7973 ( .A(n13997), .ZN(n6840) );
  OR2_X1 U7974 ( .A1(n7227), .A2(n14175), .ZN(n7223) );
  INV_X1 U7975 ( .A(n7226), .ZN(n7225) );
  INV_X1 U7976 ( .A(n14140), .ZN(n9555) );
  NOR2_X1 U7977 ( .A1(n7230), .A2(n6580), .ZN(n7224) );
  AOI21_X1 U7978 ( .B1(n7240), .B2(n7243), .A(n6563), .ZN(n7239) );
  INV_X1 U7979 ( .A(n6834), .ZN(n7240) );
  NAND2_X1 U7980 ( .A1(n14206), .A2(n14097), .ZN(n14192) );
  INV_X1 U7981 ( .A(n14077), .ZN(n14226) );
  NAND2_X1 U7982 ( .A1(n6721), .A2(n14095), .ZN(n14237) );
  NAND2_X1 U7983 ( .A1(n6542), .A2(n14071), .ZN(n14263) );
  NOR2_X1 U7984 ( .A1(n14269), .A2(n7217), .ZN(n7216) );
  INV_X1 U7985 ( .A(n14091), .ZN(n7217) );
  NAND2_X1 U7986 ( .A1(n9299), .A2(n9298), .ZN(n14086) );
  OR2_X1 U7987 ( .A1(n13906), .A2(n14661), .ZN(n11620) );
  NAND2_X1 U7988 ( .A1(n11619), .A2(n11618), .ZN(n11621) );
  INV_X1 U7989 ( .A(n11590), .ZN(n11618) );
  NAND2_X1 U7990 ( .A1(n11220), .A2(n11219), .ZN(n11222) );
  NAND2_X1 U7991 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  CLKBUF_X1 U7992 ( .A(n11015), .Z(n10976) );
  INV_X1 U7993 ( .A(n14240), .ZN(n14769) );
  NAND2_X1 U7994 ( .A1(n6544), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6689) );
  AND4_X1 U7995 ( .A1(n9042), .A2(n9041), .A3(n9040), .A4(n9039), .ZN(n10874)
         );
  OR2_X1 U7996 ( .A1(n9072), .A2(n9038), .ZN(n9039) );
  OR2_X1 U7997 ( .A1(n10032), .A2(n10235), .ZN(n14240) );
  INV_X1 U7998 ( .A(n14330), .ZN(n6958) );
  NAND2_X1 U7999 ( .A1(n9938), .A2(n9937), .ZN(n14766) );
  XNOR2_X1 U8000 ( .A(n9491), .B(n9490), .ZN(n13378) );
  AND2_X1 U8001 ( .A1(n8976), .A2(n7265), .ZN(n7261) );
  NOR2_X1 U8002 ( .A1(n8995), .A2(n14441), .ZN(n8990) );
  NOR2_X1 U8003 ( .A1(n8134), .A2(n7340), .ZN(n7339) );
  INV_X1 U8004 ( .A(n8131), .ZN(n7340) );
  NAND3_X1 U8005 ( .A1(n9313), .A2(n9584), .A3(n6752), .ZN(n9586) );
  INV_X1 U8006 ( .A(n8574), .ZN(n8110) );
  NAND2_X1 U8007 ( .A1(n8111), .A2(n8109), .ZN(n8575) );
  NAND2_X1 U8008 ( .A1(n8530), .A2(n8529), .ZN(n8553) );
  OR2_X1 U8009 ( .A1(n9222), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n9223) );
  OR2_X1 U8010 ( .A1(n14519), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U8011 ( .A1(n15430), .A2(n15431), .ZN(n7175) );
  OAI21_X1 U8012 ( .B1(P3_ADDR_REG_10__SCAN_IN), .B2(n14482), .A(n14481), .ZN(
        n14497) );
  AOI21_X1 U8013 ( .B1(P3_ADDR_REG_12__SCAN_IN), .B2(n14757), .A(n14485), .ZN(
        n14492) );
  AND2_X1 U8014 ( .A1(n14495), .A2(n14494), .ZN(n14485) );
  AND4_X1 U8015 ( .A1(n7794), .A2(n7793), .A3(n7792), .A4(n7791), .ZN(n12572)
         );
  NAND2_X1 U8016 ( .A1(n7497), .A2(n7430), .ZN(n11968) );
  INV_X1 U8017 ( .A(n12249), .ZN(n12500) );
  INV_X1 U8018 ( .A(n12005), .ZN(n12000) );
  INV_X1 U8019 ( .A(n11985), .ZN(n12004) );
  INV_X1 U8020 ( .A(n12008), .ZN(n11997) );
  OAI211_X1 U8021 ( .C1(n12236), .C2(n15363), .A(n12235), .B(n12237), .ZN(
        n12238) );
  NAND2_X1 U8022 ( .A1(n12064), .A2(n12063), .ZN(n12237) );
  INV_X1 U8023 ( .A(n10965), .ZN(n12244) );
  NAND2_X1 U8024 ( .A1(n7877), .A2(n7876), .ZN(n12448) );
  NAND2_X1 U8025 ( .A1(n15166), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n15169) );
  AND2_X1 U8026 ( .A1(n11064), .A2(n7019), .ZN(n15187) );
  INV_X1 U8027 ( .A(n15188), .ZN(n7019) );
  AND2_X1 U8028 ( .A1(n7989), .A2(n7988), .ZN(n12411) );
  NAND2_X1 U8029 ( .A1(n7823), .A2(n7822), .ZN(n12514) );
  AND2_X1 U8030 ( .A1(n7711), .A2(n7710), .ZN(n11994) );
  NAND2_X1 U8031 ( .A1(n7859), .A2(n7858), .ZN(n12717) );
  AND2_X1 U8032 ( .A1(n8006), .A2(n8005), .ZN(n10744) );
  AND2_X1 U8033 ( .A1(n8010), .A2(n8009), .ZN(n10814) );
  INV_X1 U8034 ( .A(n13237), .ZN(n13333) );
  NAND2_X1 U8035 ( .A1(n9597), .A2(n15042), .ZN(n7382) );
  NAND2_X1 U8036 ( .A1(n8618), .A2(n8617), .ZN(n13307) );
  INV_X1 U8037 ( .A(n12946), .ZN(n12938) );
  AND2_X1 U8038 ( .A1(n10169), .A2(n15146), .ZN(n12946) );
  NAND2_X1 U8039 ( .A1(n8725), .A2(n8724), .ZN(n12962) );
  NOR2_X1 U8040 ( .A1(n13090), .A2(n7429), .ZN(n7159) );
  OAI21_X1 U8041 ( .B1(n13116), .B2(n6988), .A(n6985), .ZN(n13079) );
  INV_X1 U8042 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10681) );
  NAND2_X1 U8043 ( .A1(n6727), .A2(n13773), .ZN(n6726) );
  NAND2_X1 U8044 ( .A1(n13889), .A2(n13890), .ZN(n6727) );
  INV_X1 U8045 ( .A(n13797), .ZN(n6725) );
  AND2_X1 U8046 ( .A1(n9472), .A2(n9440), .ZN(n14147) );
  NAND2_X1 U8047 ( .A1(n13873), .A2(n13745), .ZN(n13779) );
  NAND2_X1 U8048 ( .A1(n11256), .A2(n11255), .ZN(n11502) );
  NAND2_X1 U8049 ( .A1(n9357), .A2(n9356), .ZN(n14381) );
  AOI21_X1 U8050 ( .B1(n6746), .B2(n13882), .A(n6630), .ZN(n6745) );
  NAND2_X1 U8051 ( .A1(n9257), .A2(n9256), .ZN(n13869) );
  INV_X1 U8052 ( .A(n13915), .ZN(n11509) );
  INV_X1 U8053 ( .A(n14736), .ZN(n13891) );
  OR2_X1 U8054 ( .A1(n13390), .A2(n9417), .ZN(n9419) );
  AND2_X1 U8055 ( .A1(n14725), .A2(n14722), .ZN(n13905) );
  NAND4_X1 U8056 ( .A1(n9923), .A2(n9949), .A3(n9948), .A4(n10315), .ZN(n13908) );
  INV_X1 U8057 ( .A(n9575), .ZN(n6892) );
  AOI21_X1 U8058 ( .B1(n9574), .B2(n9573), .A(n9572), .ZN(n9575) );
  NAND2_X1 U8059 ( .A1(n9571), .A2(n9530), .ZN(n9576) );
  INV_X1 U8060 ( .A(n14239), .ZN(n14094) );
  NOR2_X1 U8061 ( .A1(n10269), .A2(n6605), .ZN(n13969) );
  NAND2_X1 U8062 ( .A1(n13969), .A2(n13970), .ZN(n13968) );
  NAND2_X1 U8063 ( .A1(n13979), .A2(n6665), .ZN(n10371) );
  OAI21_X1 U8064 ( .B1(n14037), .B2(n14036), .A(n6849), .ZN(n6848) );
  AOI21_X1 U8065 ( .B1(n14038), .B2(n14752), .A(n14750), .ZN(n6849) );
  AND2_X1 U8066 ( .A1(n9344), .A2(n9343), .ZN(n14261) );
  INV_X1 U8067 ( .A(n14808), .ZN(n14309) );
  NAND2_X1 U8068 ( .A1(n14113), .A2(n14775), .ZN(n14774) );
  NOR2_X1 U8069 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n7212) );
  XNOR2_X1 U8071 ( .A(n9023), .B(n9022), .ZN(n10687) );
  XNOR2_X1 U8072 ( .A(n14504), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15426) );
  NAND2_X1 U8073 ( .A1(n6769), .A2(n6768), .ZN(n14550) );
  NAND2_X1 U8074 ( .A1(n14710), .A2(n6770), .ZN(n6769) );
  AOI21_X1 U8075 ( .B1(n6767), .B2(n6766), .A(n6765), .ZN(n14713) );
  NAND2_X1 U8076 ( .A1(n6770), .A2(n14549), .ZN(n6765) );
  AND2_X1 U8077 ( .A1(n14704), .A2(n6768), .ZN(n6766) );
  OR2_X1 U8078 ( .A1(n14713), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7188) );
  INV_X1 U8079 ( .A(n7174), .ZN(n14606) );
  INV_X1 U8080 ( .A(n14605), .ZN(n7173) );
  NOR2_X1 U8081 ( .A1(n15042), .A2(n9593), .ZN(n9595) );
  NAND2_X1 U8082 ( .A1(n9629), .A2(n7406), .ZN(n7405) );
  NAND2_X1 U8083 ( .A1(n9639), .A2(n9641), .ZN(n7398) );
  NAND2_X1 U8084 ( .A1(n9650), .A2(n9652), .ZN(n7396) );
  NAND2_X1 U8085 ( .A1(n7294), .A2(n9138), .ZN(n7293) );
  OR2_X1 U8086 ( .A1(n7294), .A2(n9138), .ZN(n7292) );
  OR2_X1 U8087 ( .A1(n12087), .A2(n12219), .ZN(n6711) );
  NAND2_X1 U8088 ( .A1(n9172), .A2(n7290), .ZN(n7289) );
  AND2_X1 U8089 ( .A1(n12097), .A2(n12096), .ZN(n6700) );
  NOR2_X1 U8090 ( .A1(n7389), .A2(n6618), .ZN(n7387) );
  INV_X1 U8091 ( .A(n9693), .ZN(n7389) );
  NAND2_X1 U8092 ( .A1(n9211), .A2(n7287), .ZN(n7286) );
  NAND2_X1 U8093 ( .A1(n9715), .A2(n9717), .ZN(n7392) );
  NAND2_X1 U8094 ( .A1(n7272), .A2(n7271), .ZN(n7270) );
  NAND2_X1 U8095 ( .A1(n9286), .A2(n7273), .ZN(n7272) );
  NAND2_X1 U8096 ( .A1(n9286), .A2(n9300), .ZN(n7271) );
  OR2_X1 U8097 ( .A1(n12146), .A2(n12219), .ZN(n6703) );
  OR2_X1 U8098 ( .A1(n7415), .A2(n9727), .ZN(n7414) );
  INV_X1 U8099 ( .A(n9726), .ZN(n7415) );
  NAND2_X1 U8100 ( .A1(n9371), .A2(n6905), .ZN(n6904) );
  NOR2_X1 U8101 ( .A1(n7282), .A2(n9359), .ZN(n6905) );
  NAND2_X1 U8102 ( .A1(n7409), .A2(n9738), .ZN(n7408) );
  AND2_X1 U8103 ( .A1(n9384), .A2(n7298), .ZN(n7297) );
  INV_X1 U8104 ( .A(n9382), .ZN(n7298) );
  NAND2_X1 U8105 ( .A1(n6707), .A2(n12227), .ZN(n6706) );
  INV_X1 U8106 ( .A(n12188), .ZN(n6707) );
  NAND2_X1 U8107 ( .A1(n9416), .A2(n9414), .ZN(n7283) );
  NAND2_X1 U8108 ( .A1(n7965), .A2(n12464), .ZN(n7975) );
  NOR2_X1 U8109 ( .A1(n7096), .A2(n7843), .ZN(n7095) );
  NOR2_X1 U8110 ( .A1(n7099), .A2(n6670), .ZN(n7096) );
  INV_X1 U8111 ( .A(n7084), .ZN(n7083) );
  OAI21_X1 U8112 ( .B1(n7782), .B2(n7085), .A(n7796), .ZN(n7084) );
  INV_X1 U8113 ( .A(n7476), .ZN(n7085) );
  OAI21_X1 U8114 ( .B1(n13270), .B2(n9779), .A(n7308), .ZN(n9791) );
  NAND2_X1 U8115 ( .A1(n9778), .A2(n9779), .ZN(n7308) );
  NAND2_X1 U8116 ( .A1(n9803), .A2(n9783), .ZN(n9832) );
  AND2_X2 U8117 ( .A1(n8894), .A2(n8783), .ZN(n9593) );
  INV_X1 U8118 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8142) );
  INV_X1 U8119 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8138) );
  AND2_X1 U8120 ( .A1(n9451), .A2(n7296), .ZN(n7295) );
  INV_X1 U8121 ( .A(n9449), .ZN(n7296) );
  NAND2_X1 U8122 ( .A1(n9024), .A2(n7274), .ZN(n7276) );
  NAND2_X1 U8123 ( .A1(n9498), .A2(n10813), .ZN(n7275) );
  AND2_X1 U8124 ( .A1(n9952), .A2(n9862), .ZN(n7274) );
  AND2_X1 U8125 ( .A1(n7320), .A2(n8103), .ZN(n7319) );
  NAND2_X1 U8126 ( .A1(n7321), .A2(n7323), .ZN(n7320) );
  INV_X1 U8127 ( .A(n7324), .ZN(n7321) );
  INV_X1 U8128 ( .A(n8107), .ZN(n7318) );
  INV_X1 U8129 ( .A(n7323), .ZN(n7322) );
  INV_X1 U8130 ( .A(n6832), .ZN(n6831) );
  OAI21_X1 U8131 ( .B1(n6579), .B2(n6833), .A(n7319), .ZN(n6832) );
  NAND2_X1 U8132 ( .A1(n6831), .A2(n6833), .ZN(n6828) );
  NAND2_X1 U8133 ( .A1(n7325), .A2(SI_17_), .ZN(n7324) );
  INV_X1 U8134 ( .A(n8505), .ZN(n7325) );
  NAND2_X1 U8135 ( .A1(n8505), .A2(n10359), .ZN(n7323) );
  INV_X1 U8136 ( .A(SI_16_), .ZN(n8098) );
  AND2_X1 U8137 ( .A1(n6826), .A2(n7436), .ZN(n6825) );
  INV_X1 U8138 ( .A(n7330), .ZN(n7329) );
  OAI21_X1 U8139 ( .B1(n8066), .B2(n7331), .A(n8069), .ZN(n7330) );
  INV_X1 U8140 ( .A(n8068), .ZN(n7331) );
  OAI21_X1 U8141 ( .B1(n9367), .B2(n6713), .A(n6712), .ZN(n8055) );
  NAND2_X1 U8142 ( .A1(n9367), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6712) );
  INV_X1 U8143 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7494) );
  OAI211_X1 U8144 ( .C1(n12217), .C2(n12216), .A(n12215), .B(n12214), .ZN(
        n12225) );
  AND2_X1 U8145 ( .A1(n12232), .A2(n12226), .ZN(n7064) );
  NAND2_X1 U8146 ( .A1(n7536), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U8147 ( .A1(n6697), .A2(n6696), .ZN(n10594) );
  OR2_X1 U8148 ( .A1(n12774), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8149 ( .A1(n12774), .A2(n10617), .ZN(n6696) );
  NAND2_X1 U8150 ( .A1(n15234), .A2(n6801), .ZN(n11130) );
  OR2_X1 U8151 ( .A1(n11129), .A2(n11092), .ZN(n6801) );
  NAND2_X1 U8152 ( .A1(n11694), .A2(n6803), .ZN(n12272) );
  OR2_X1 U8153 ( .A1(n11698), .A2(n14636), .ZN(n6803) );
  NAND2_X1 U8154 ( .A1(n6783), .A2(n6781), .ZN(n6776) );
  NAND2_X1 U8155 ( .A1(n12217), .A2(n6778), .ZN(n6777) );
  NAND2_X1 U8156 ( .A1(n6779), .A2(n6781), .ZN(n6778) );
  OR2_X1 U8157 ( .A1(n7847), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7849) );
  OR2_X1 U8158 ( .A1(n7836), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7847) );
  OR2_X1 U8159 ( .A1(n7669), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7684) );
  INV_X1 U8160 ( .A(n12780), .ZN(n8026) );
  AND2_X1 U8161 ( .A1(n6593), .A2(n7068), .ZN(n7067) );
  NOR2_X1 U8162 ( .A1(P3_IR_REG_25__SCAN_IN), .A2(P3_IR_REG_28__SCAN_IN), .ZN(
        n7068) );
  AND2_X1 U8163 ( .A1(n6593), .A2(n7993), .ZN(n7066) );
  NAND2_X1 U8164 ( .A1(n13394), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7114) );
  INV_X1 U8165 ( .A(n7867), .ZN(n7112) );
  NAND2_X1 U8166 ( .A1(n7489), .A2(n7052), .ZN(n7051) );
  NOR2_X1 U8167 ( .A1(P3_IR_REG_21__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7052) );
  INV_X1 U8168 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n6881) );
  INV_X1 U8169 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n6882) );
  INV_X1 U8170 ( .A(n6674), .ZN(n6792) );
  INV_X1 U8171 ( .A(n7478), .ZN(n6789) );
  OR2_X1 U8172 ( .A1(n7729), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7743) );
  INV_X1 U8173 ( .A(n7105), .ZN(n7104) );
  OAI21_X1 U8174 ( .B1(n7695), .B2(n7106), .A(n7464), .ZN(n7105) );
  NAND2_X1 U8175 ( .A1(n7462), .A2(n7461), .ZN(n7106) );
  NOR2_X1 U8176 ( .A1(n7695), .A2(n7108), .ZN(n7107) );
  INV_X1 U8177 ( .A(n7461), .ZN(n7108) );
  OR2_X1 U8178 ( .A1(n9800), .A2(n13053), .ZN(n9803) );
  NAND2_X1 U8179 ( .A1(n8719), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8185) );
  NOR2_X1 U8180 ( .A1(n13274), .A2(n7204), .ZN(n7203) );
  INV_X1 U8181 ( .A(n7205), .ZN(n7204) );
  NOR2_X1 U8182 ( .A1(n13280), .A2(n13287), .ZN(n7205) );
  AOI21_X1 U8183 ( .B1(n13189), .B2(n8934), .A(n6615), .ZN(n7006) );
  INV_X1 U8184 ( .A(n13178), .ZN(n7153) );
  AOI21_X1 U8185 ( .B1(n7148), .B2(n7146), .A(n9821), .ZN(n7145) );
  INV_X1 U8186 ( .A(n7149), .ZN(n7146) );
  INV_X1 U8187 ( .A(n7148), .ZN(n7147) );
  NOR2_X1 U8188 ( .A1(n15020), .A2(n13348), .ZN(n7210) );
  INV_X1 U8189 ( .A(n6966), .ZN(n6965) );
  OAI21_X1 U8190 ( .B1(n8913), .B2(n6967), .A(n9818), .ZN(n6966) );
  INV_X1 U8191 ( .A(n8914), .ZN(n6967) );
  AND2_X1 U8192 ( .A1(n6993), .A2(n8909), .ZN(n6989) );
  AND2_X1 U8193 ( .A1(n6995), .A2(n8909), .ZN(n6992) );
  NAND2_X1 U8194 ( .A1(n8842), .A2(n10299), .ZN(n8902) );
  NOR2_X1 U8195 ( .A1(n7139), .A2(n7138), .ZN(n7137) );
  NAND2_X1 U8196 ( .A1(n8790), .A2(n8149), .ZN(n7140) );
  NOR2_X1 U8197 ( .A1(n8150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8198 ( .A1(n10653), .A2(n8853), .ZN(n10772) );
  NOR2_X2 U8199 ( .A1(n8534), .A2(n7008), .ZN(n7139) );
  NAND2_X1 U8200 ( .A1(n7401), .A2(n7435), .ZN(n7008) );
  OR2_X1 U8201 ( .A1(n8472), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n8473) );
  AND2_X1 U8202 ( .A1(n8407), .A2(n8406), .ZN(n8427) );
  NOR2_X1 U8203 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6810) );
  INV_X1 U8204 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14463) );
  INV_X1 U8205 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n13500) );
  INV_X1 U8206 ( .A(n10694), .ZN(n7381) );
  NAND2_X1 U8207 ( .A1(n7381), .A2(n7379), .ZN(n7378) );
  NAND2_X1 U8208 ( .A1(n9024), .A2(n9862), .ZN(n9498) );
  OR2_X1 U8209 ( .A1(n9467), .A2(n9483), .ZN(n6895) );
  AND2_X1 U8210 ( .A1(n9265), .A2(n9094), .ZN(n9134) );
  OAI22_X1 U8211 ( .A1(n14140), .A2(n7229), .B1(n14158), .B2(n14149), .ZN(
        n7226) );
  NAND2_X1 U8212 ( .A1(n14181), .A2(n6596), .ZN(n6937) );
  INV_X1 U8213 ( .A(n14338), .ZN(n6935) );
  NOR2_X1 U8214 ( .A1(n14347), .A2(n14343), .ZN(n6936) );
  AND2_X1 U8215 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n9401), .ZN(n9402) );
  INV_X1 U8216 ( .A(n14099), .ZN(n6951) );
  NOR2_X1 U8217 ( .A1(n11171), .A2(n10978), .ZN(n6954) );
  INV_X1 U8218 ( .A(n10889), .ZN(n7247) );
  AND2_X1 U8219 ( .A1(n14793), .A2(n14897), .ZN(n14759) );
  NAND2_X1 U8220 ( .A1(n8884), .A2(n8883), .ZN(n9486) );
  NAND2_X1 U8221 ( .A1(n7335), .A2(n8133), .ZN(n7334) );
  NAND2_X1 U8222 ( .A1(n6629), .A2(n8097), .ZN(n7313) );
  NOR2_X1 U8223 ( .A1(n8096), .A2(n7316), .ZN(n7315) );
  NAND2_X1 U8224 ( .A1(n8097), .A2(n8088), .ZN(n7316) );
  AOI21_X1 U8225 ( .B1(n6825), .B2(n6823), .A(n6822), .ZN(n6821) );
  INV_X1 U8226 ( .A(n8084), .ZN(n6822) );
  INV_X1 U8227 ( .A(n8080), .ZN(n6823) );
  INV_X1 U8228 ( .A(n6825), .ZN(n6824) );
  OR2_X1 U8229 ( .A1(n9148), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9168) );
  NAND2_X1 U8230 ( .A1(n7312), .A2(n8061), .ZN(n6913) );
  CLKBUF_X1 U8231 ( .A(n9065), .Z(n9066) );
  NAND2_X1 U8232 ( .A1(n8043), .A2(n9982), .ZN(n7301) );
  NAND2_X1 U8233 ( .A1(n14461), .A2(n7179), .ZN(n14464) );
  NAND2_X1 U8234 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7180), .ZN(n7179) );
  NAND2_X1 U8235 ( .A1(n7181), .A2(n14467), .ZN(n14468) );
  OR2_X1 U8236 ( .A1(n14503), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n7181) );
  AOI22_X1 U8237 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n14527), .B1(n14528), .B2(
        n14471), .ZN(n14473) );
  OR2_X1 U8238 ( .A1(n14527), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n14471) );
  INV_X1 U8239 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14484) );
  OR2_X1 U8240 ( .A1(n7719), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7733) );
  NAND2_X1 U8241 ( .A1(n12701), .A2(n12078), .ZN(n10821) );
  NAND2_X1 U8242 ( .A1(n11972), .A2(n6604), .ZN(n11934) );
  INV_X1 U8243 ( .A(n11937), .ZN(n6867) );
  INV_X1 U8244 ( .A(n11411), .ZN(n11272) );
  NOR2_X1 U8245 ( .A1(n7803), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7814) );
  AND2_X1 U8246 ( .A1(n7814), .A2(n7813), .ZN(n7824) );
  NAND2_X1 U8247 ( .A1(n11787), .A2(n11786), .ZN(n11989) );
  OR2_X1 U8248 ( .A1(n7789), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7803) );
  NOR4_X1 U8249 ( .A1(n12061), .A2(n12206), .A3(n12060), .A4(n12217), .ZN(
        n12062) );
  AND2_X1 U8250 ( .A1(n7058), .A2(n12218), .ZN(n7057) );
  OR2_X1 U8251 ( .A1(n7061), .A2(n7060), .ZN(n7058) );
  NAND2_X1 U8252 ( .A1(n7515), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7024) );
  NOR2_X1 U8253 ( .A1(n10599), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10782) );
  INV_X1 U8254 ( .A(n6799), .ZN(n6798) );
  INV_X1 U8255 ( .A(n11124), .ZN(n15200) );
  NAND2_X1 U8256 ( .A1(n15217), .A2(n11128), .ZN(n15236) );
  NAND2_X1 U8257 ( .A1(n15236), .A2(n15235), .ZN(n15234) );
  XNOR2_X1 U8258 ( .A(n11130), .B(n11131), .ZN(n15253) );
  OAI21_X1 U8259 ( .B1(n15245), .B2(n15244), .A(n15243), .ZN(n15265) );
  NAND2_X1 U8260 ( .A1(n15258), .A2(n11069), .ZN(n15259) );
  AOI21_X1 U8261 ( .B1(n15265), .B2(n15264), .A(n15263), .ZN(n15284) );
  NAND2_X1 U8262 ( .A1(n15294), .A2(n11137), .ZN(n11138) );
  NOR2_X1 U8263 ( .A1(n11435), .A2(n11434), .ZN(n11528) );
  NAND2_X1 U8264 ( .A1(n11075), .A2(n7013), .ZN(n7012) );
  NAND2_X1 U8265 ( .A1(n11523), .A2(n11448), .ZN(n11449) );
  NAND2_X1 U8266 ( .A1(n11449), .A2(n11450), .ZN(n11694) );
  XNOR2_X1 U8267 ( .A(n12272), .B(n6802), .ZN(n11695) );
  AND2_X1 U8268 ( .A1(n11701), .A2(n11700), .ZN(n12265) );
  NAND2_X1 U8269 ( .A1(n12295), .A2(n12319), .ZN(n7017) );
  AND2_X1 U8270 ( .A1(n12320), .A2(n12319), .ZN(n6690) );
  NAND2_X1 U8271 ( .A1(n7011), .A2(n6694), .ZN(n7010) );
  INV_X1 U8272 ( .A(n12344), .ZN(n7011) );
  INV_X1 U8273 ( .A(n12331), .ZN(n12356) );
  AND2_X1 U8274 ( .A1(n12029), .A2(n12028), .ZN(n12042) );
  OR2_X1 U8275 ( .A1(n14614), .A2(n7900), .ZN(n11904) );
  INV_X1 U8276 ( .A(n12065), .ZN(n12432) );
  NAND2_X1 U8277 ( .A1(n7037), .A2(n7035), .ZN(n12433) );
  AOI21_X1 U8278 ( .B1(n7038), .B2(n7040), .A(n7036), .ZN(n7035) );
  NAND2_X1 U8279 ( .A1(n7419), .A2(n7038), .ZN(n7037) );
  INV_X1 U8280 ( .A(n12066), .ZN(n7036) );
  AND2_X1 U8281 ( .A1(n12068), .A2(n12188), .ZN(n12480) );
  AND2_X1 U8282 ( .A1(n12187), .A2(n12191), .ZN(n12497) );
  AOI21_X1 U8283 ( .B1(n7045), .B2(n7043), .A(n7042), .ZN(n7041) );
  INV_X1 U8284 ( .A(n7045), .ZN(n7044) );
  INV_X1 U8285 ( .A(n12176), .ZN(n7042) );
  NAND2_X1 U8286 ( .A1(n7962), .A2(n7961), .ZN(n12535) );
  INV_X1 U8287 ( .A(n12533), .ZN(n7962) );
  AND2_X1 U8288 ( .A1(n12161), .A2(n12167), .ZN(n12552) );
  NOR2_X1 U8289 ( .A1(n7733), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7751) );
  AND2_X1 U8290 ( .A1(n7751), .A2(n7750), .ZN(n7764) );
  AND4_X1 U8291 ( .A1(n7756), .A2(n7755), .A3(n7754), .A4(n7753), .ZN(n12607)
         );
  OR2_X1 U8292 ( .A1(n7772), .A2(n7771), .ZN(n11776) );
  AND4_X1 U8293 ( .A1(n7690), .A2(n7689), .A3(n7688), .A4(n7687), .ZN(n11799)
         );
  NAND2_X1 U8294 ( .A1(n7668), .A2(n12127), .ZN(n12562) );
  AND2_X1 U8295 ( .A1(n12137), .A2(n12128), .ZN(n12135) );
  OR2_X1 U8296 ( .A1(n7654), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7669) );
  AND3_X1 U8297 ( .A1(n7667), .A2(n7666), .A3(n7665), .ZN(n11634) );
  AOI21_X1 U8298 ( .B1(n12113), .B2(n7032), .A(n7031), .ZN(n7030) );
  INV_X1 U8299 ( .A(n12110), .ZN(n7032) );
  AND2_X1 U8300 ( .A1(n7619), .A2(n11749), .ZN(n7636) );
  OR2_X1 U8301 ( .A1(n7589), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7602) );
  INV_X1 U8302 ( .A(n15352), .ZN(n15328) );
  INV_X1 U8303 ( .A(n15406), .ZN(n14625) );
  NAND2_X1 U8304 ( .A1(n7884), .A2(n7883), .ZN(n12202) );
  AND2_X1 U8305 ( .A1(n7718), .A2(n7717), .ZN(n11800) );
  INV_X1 U8306 ( .A(n11994), .ZN(n14629) );
  OR2_X1 U8307 ( .A1(n15352), .A2(n15400), .ZN(n14640) );
  INV_X1 U8308 ( .A(n10039), .ZN(n10199) );
  OAI21_X1 U8309 ( .B1(n7893), .B2(n7894), .A(n7090), .ZN(n8808) );
  NAND2_X1 U8310 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7091), .ZN(n7090) );
  XNOR2_X1 U8311 ( .A(n8030), .B(n8029), .ZN(n10575) );
  INV_X1 U8312 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U8313 ( .A1(n7466), .A2(n6794), .ZN(n7712) );
  INV_X1 U8314 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7714) );
  AOI21_X1 U8315 ( .B1(n7071), .B2(n6565), .A(n6666), .ZN(n6787) );
  XNOR2_X1 U8316 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7611) );
  NAND2_X1 U8317 ( .A1(n6784), .A2(n7076), .ZN(n7598) );
  AOI21_X1 U8318 ( .B1(n7077), .B2(n7577), .A(n6626), .ZN(n7076) );
  NAND2_X1 U8319 ( .A1(n7564), .A2(n7074), .ZN(n6784) );
  XNOR2_X1 U8320 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7547) );
  AND2_X1 U8321 ( .A1(n8186), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7522) );
  XNOR2_X1 U8322 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7523) );
  OR2_X1 U8323 ( .A1(n8339), .A2(n13652), .ZN(n8354) );
  NAND2_X1 U8324 ( .A1(n11334), .A2(n8420), .ZN(n11362) );
  INV_X1 U8325 ( .A(n12886), .ZN(n12933) );
  OR2_X1 U8326 ( .A1(n10140), .A2(n10139), .ZN(n6922) );
  NAND2_X1 U8327 ( .A1(n6922), .A2(n6921), .ZN(n6920) );
  NAND2_X1 U8328 ( .A1(n10127), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U8329 ( .A1(n14985), .A2(n6928), .ZN(n10499) );
  AND2_X1 U8330 ( .A1(n14990), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6928) );
  NOR2_X1 U8331 ( .A1(n10499), .A2(n10498), .ZN(n10540) );
  NOR2_X1 U8332 ( .A1(n11152), .A2(n6926), .ZN(n11155) );
  AND2_X1 U8333 ( .A1(n11153), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U8334 ( .A1(n11155), .A2(n11154), .ZN(n11657) );
  XNOR2_X1 U8335 ( .A(n11659), .B(n15013), .ZN(n15004) );
  NOR2_X1 U8336 ( .A1(n11657), .A2(n6925), .ZN(n11659) );
  AND2_X1 U8337 ( .A1(n11658), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6925) );
  NAND2_X1 U8338 ( .A1(n9768), .A2(n9767), .ZN(n13052) );
  NAND2_X1 U8339 ( .A1(n13112), .A2(n7203), .ZN(n13071) );
  AND2_X1 U8340 ( .A1(n8738), .A2(n8737), .ZN(n13072) );
  INV_X1 U8341 ( .A(n13105), .ZN(n6988) );
  NAND2_X1 U8342 ( .A1(n13112), .A2(n13103), .ZN(n13098) );
  AOI21_X1 U8343 ( .B1(n6575), .B2(n6981), .A(n6976), .ZN(n6975) );
  NAND2_X1 U8344 ( .A1(n13165), .A2(n6575), .ZN(n6977) );
  INV_X1 U8345 ( .A(n8939), .ZN(n6976) );
  OR2_X1 U8346 ( .A1(n8656), .A2(n13650), .ZN(n8676) );
  NAND2_X1 U8347 ( .A1(n13192), .A2(n13177), .ZN(n13171) );
  AOI21_X1 U8348 ( .B1(n7156), .B2(n7155), .A(n6662), .ZN(n7154) );
  INV_X1 U8349 ( .A(n9808), .ZN(n7155) );
  NAND2_X1 U8350 ( .A1(n8559), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8580) );
  INV_X1 U8351 ( .A(n6999), .ZN(n6998) );
  OAI21_X1 U8352 ( .B1(n8930), .B2(n7000), .A(n8929), .ZN(n6999) );
  NAND2_X1 U8353 ( .A1(n7201), .A2(n7200), .ZN(n13200) );
  INV_X1 U8354 ( .A(n7201), .ZN(n13220) );
  INV_X1 U8355 ( .A(n8516), .ZN(n8514) );
  NOR2_X1 U8356 ( .A1(n11540), .A2(n13339), .ZN(n13229) );
  NAND2_X1 U8357 ( .A1(n7143), .A2(n7141), .ZN(n13228) );
  AOI21_X1 U8358 ( .B1(n7145), .B2(n7147), .A(n7142), .ZN(n7141) );
  NAND2_X1 U8359 ( .A1(n8862), .A2(n7145), .ZN(n7143) );
  INV_X1 U8360 ( .A(n8865), .ZN(n7142) );
  NAND2_X1 U8361 ( .A1(n6548), .A2(n7206), .ZN(n11540) );
  INV_X1 U8362 ( .A(n8453), .ZN(n8452) );
  NAND2_X1 U8363 ( .A1(n7208), .A2(n7207), .ZN(n11477) );
  INV_X1 U8364 ( .A(n11369), .ZN(n7208) );
  NAND2_X1 U8365 ( .A1(n7007), .A2(n8918), .ZN(n11347) );
  NAND2_X1 U8366 ( .A1(n8917), .A2(n6578), .ZN(n7007) );
  NAND2_X1 U8367 ( .A1(n7210), .A2(n7209), .ZN(n11369) );
  NAND2_X1 U8368 ( .A1(n7132), .A2(n8859), .ZN(n11340) );
  INV_X1 U8369 ( .A(n7210), .ZN(n11341) );
  NAND2_X1 U8370 ( .A1(n10850), .A2(n8855), .ZN(n10834) );
  NAND2_X1 U8371 ( .A1(n13257), .A2(n15112), .ZN(n10773) );
  NAND2_X1 U8372 ( .A1(n6970), .A2(n6969), .ZN(n10642) );
  NAND2_X1 U8373 ( .A1(n10395), .A2(n6971), .ZN(n6970) );
  NOR2_X1 U8374 ( .A1(n6974), .A2(n6972), .ZN(n6971) );
  NAND2_X1 U8375 ( .A1(n6973), .A2(n8905), .ZN(n10643) );
  NAND2_X1 U8376 ( .A1(n10412), .A2(n10411), .ZN(n6973) );
  NAND2_X1 U8377 ( .A1(n10395), .A2(n8904), .ZN(n10412) );
  INV_X1 U8378 ( .A(n10392), .ZN(n10396) );
  INV_X1 U8379 ( .A(n10326), .ZN(n10334) );
  NAND2_X1 U8380 ( .A1(n9812), .A2(n8901), .ZN(n10305) );
  NOR2_X1 U8381 ( .A1(n15139), .A2(n9847), .ZN(n8799) );
  OAI21_X1 U8382 ( .B1(n8946), .B2(n12884), .A(n8957), .ZN(n8958) );
  NAND2_X1 U8383 ( .A1(n8371), .A2(n8370), .ZN(n15136) );
  CLKBUF_X1 U8384 ( .A(n8888), .Z(n15119) );
  INV_X1 U8385 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8949) );
  AND2_X1 U8386 ( .A1(n8751), .A2(n8758), .ZN(n8777) );
  XNOR2_X1 U8387 ( .A(n8780), .B(n8779), .ZN(n10054) );
  INV_X1 U8388 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8779) );
  INV_X1 U8389 ( .A(n8614), .ZN(n8118) );
  INV_X1 U8390 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8165) );
  XNOR2_X1 U8391 ( .A(n8168), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9844) );
  CLKBUF_X1 U8392 ( .A(P2_IR_REG_10__SCAN_IN), .Z(n8386) );
  OR2_X1 U8393 ( .A1(n8368), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n8510) );
  INV_X1 U8394 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8269) );
  CLKBUF_X1 U8395 ( .A(n8174), .Z(n8203) );
  NOR2_X1 U8396 ( .A1(n9960), .A2(n9989), .ZN(n6944) );
  INV_X1 U8397 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n13602) );
  OR2_X1 U8398 ( .A1(n9335), .A2(n13856), .ZN(n9350) );
  NAND2_X1 U8399 ( .A1(n9325), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9335) );
  INV_X1 U8400 ( .A(n13727), .ZN(n6751) );
  INV_X1 U8401 ( .A(n13725), .ZN(n6747) );
  NAND2_X1 U8402 ( .A1(n13808), .A2(n13738), .ZN(n13874) );
  NOR2_X1 U8403 ( .A1(n13877), .A2(n9360), .ZN(n9373) );
  XNOR2_X1 U8404 ( .A(n9874), .B(n6549), .ZN(n9875) );
  XNOR2_X1 U8405 ( .A(n9863), .B(n6549), .ZN(n7341) );
  NAND2_X1 U8406 ( .A1(n9483), .A2(n9482), .ZN(n6896) );
  INV_X1 U8407 ( .A(n9070), .ZN(n9213) );
  INV_X1 U8408 ( .A(n9475), .ZN(n9494) );
  NAND2_X1 U8409 ( .A1(n9423), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n8987) );
  OR2_X1 U8410 ( .A1(n9071), .A2(n8999), .ZN(n9002) );
  OR2_X1 U8411 ( .A1(n10254), .A2(n10255), .ZN(n6846) );
  OR2_X1 U8412 ( .A1(n10283), .A2(n10284), .ZN(n6844) );
  XNOR2_X1 U8413 ( .A(n14025), .B(n14024), .ZN(n14013) );
  INV_X1 U8414 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9009) );
  NOR2_X1 U8415 ( .A1(n14011), .A2(n6839), .ZN(n14025) );
  AND2_X1 U8416 ( .A1(n14012), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6839) );
  NAND2_X1 U8417 ( .A1(n9522), .A2(n9521), .ZN(n14049) );
  OR2_X2 U8418 ( .A1(n6937), .A2(n9556), .ZN(n14107) );
  NAND2_X1 U8419 ( .A1(n14181), .A2(n6936), .ZN(n14145) );
  NAND2_X1 U8420 ( .A1(n14181), .A2(n14167), .ZN(n14166) );
  NAND2_X1 U8421 ( .A1(n6960), .A2(n6959), .ZN(n14196) );
  AOI21_X1 U8422 ( .B1(n14221), .B2(n6934), .A(n6659), .ZN(n6933) );
  NAND2_X1 U8423 ( .A1(n14208), .A2(n14207), .ZN(n14206) );
  NAND2_X1 U8424 ( .A1(n6961), .A2(n14231), .ZN(n14227) );
  NOR2_X2 U8425 ( .A1(n14392), .A2(n14293), .ZN(n14271) );
  NOR2_X1 U8426 ( .A1(n9308), .A2(n13602), .ZN(n9309) );
  AND2_X1 U8427 ( .A1(n9309), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9325) );
  NOR2_X1 U8428 ( .A1(n14086), .A2(n11622), .ZN(n14307) );
  NAND2_X1 U8429 ( .A1(n6956), .A2(n6955), .ZN(n11622) );
  OR2_X1 U8430 ( .A1(n9214), .A2(n13533), .ZN(n9245) );
  NAND2_X1 U8431 ( .A1(n9225), .A2(n9224), .ZN(n11605) );
  NAND2_X1 U8432 ( .A1(n9210), .A2(n9209), .ZN(n11494) );
  INV_X1 U8433 ( .A(n13913), .ZN(n13865) );
  AOI21_X1 U8434 ( .B1(n7235), .B2(n7237), .A(n6613), .ZN(n7233) );
  INV_X1 U8435 ( .A(n11011), .ZN(n6942) );
  NAND3_X1 U8436 ( .A1(n6560), .A2(n6953), .A3(n14793), .ZN(n11230) );
  NAND2_X1 U8437 ( .A1(n6560), .A2(n14793), .ZN(n11017) );
  AND2_X1 U8438 ( .A1(n14793), .A2(n6954), .ZN(n14761) );
  OR2_X1 U8439 ( .A1(n9126), .A2(n9125), .ZN(n9141) );
  INV_X1 U8440 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9140) );
  OR2_X1 U8441 ( .A1(n9141), .A2(n9140), .ZN(n9160) );
  NAND2_X1 U8442 ( .A1(n10894), .A2(n10893), .ZN(n10913) );
  AND2_X1 U8443 ( .A1(n9069), .A2(n9068), .ZN(n10943) );
  INV_X1 U8444 ( .A(n10943), .ZN(n10942) );
  NAND2_X1 U8445 ( .A1(n10868), .A2(n9535), .ZN(n14801) );
  NAND2_X1 U8446 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  AND2_X1 U8447 ( .A1(n7250), .A2(n7249), .ZN(n14122) );
  NOR2_X2 U8448 ( .A1(n9951), .A2(n9902), .ZN(n14722) );
  INV_X1 U8449 ( .A(n10988), .ZN(n14899) );
  INV_X1 U8450 ( .A(n14722), .ZN(n14920) );
  INV_X1 U8451 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7263) );
  XNOR2_X1 U8452 ( .A(n9486), .B(n9485), .ZN(n11821) );
  NAND2_X1 U8453 ( .A1(n9313), .A2(n8976), .ZN(n7213) );
  NAND2_X1 U8454 ( .A1(n8692), .A2(n8131), .ZN(n8715) );
  INV_X1 U8455 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9587) );
  NAND2_X1 U8456 ( .A1(n8126), .A2(n8128), .ZN(n8651) );
  XNOR2_X1 U8457 ( .A(n9019), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9528) );
  INV_X1 U8458 ( .A(n9018), .ZN(n9019) );
  INV_X1 U8459 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9022) );
  AND2_X1 U8460 ( .A1(n9255), .A2(n9254), .ZN(n10724) );
  NAND2_X1 U8461 ( .A1(n7328), .A2(n8068), .ZN(n8345) );
  NAND2_X1 U8462 ( .A1(n8331), .A2(n8066), .ZN(n7328) );
  NAND2_X1 U8463 ( .A1(n8265), .A2(n8058), .ZN(n7311) );
  INV_X1 U8464 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7267) );
  INV_X1 U8465 ( .A(n8050), .ZN(n8224) );
  XNOR2_X1 U8466 ( .A(n8041), .B(SI_1_), .ZN(n8170) );
  NAND2_X1 U8467 ( .A1(n6763), .A2(n14509), .ZN(n14512) );
  NAND2_X1 U8468 ( .A1(n15437), .A2(n15438), .ZN(n6763) );
  XNOR2_X1 U8469 ( .A(n14464), .B(n7178), .ZN(n14516) );
  XNOR2_X1 U8470 ( .A(n14503), .B(n14502), .ZN(n14504) );
  INV_X1 U8471 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n14527) );
  NAND2_X1 U8472 ( .A1(n14530), .A2(n14531), .ZN(n14533) );
  INV_X1 U8473 ( .A(n6754), .ZN(n14541) );
  OAI21_X1 U8474 ( .B1(n14591), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6589), .ZN(
        n6754) );
  AOI21_X1 U8475 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(n14479), .A(n14478), .ZN(
        n14499) );
  AOI21_X1 U8476 ( .B1(n14484), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n14483), .ZN(
        n14494) );
  AND2_X1 U8477 ( .A1(n14496), .A2(n14497), .ZN(n14483) );
  OR2_X1 U8478 ( .A1(n14711), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6770) );
  NAND2_X1 U8479 ( .A1(n14711), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n6768) );
  NOR2_X1 U8480 ( .A1(n14557), .A2(n14556), .ZN(n14563) );
  NOR2_X1 U8481 ( .A1(n14720), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n14557) );
  OAI21_X1 U8482 ( .B1(n11787), .B2(n6873), .A(n6870), .ZN(n11825) );
  NAND3_X1 U8483 ( .A1(n11636), .A2(n11637), .A3(n11635), .ZN(n11713) );
  OR2_X1 U8484 ( .A1(n11041), .A2(n11042), .ZN(n11040) );
  NAND2_X1 U8485 ( .A1(n7427), .A2(n10506), .ZN(n10820) );
  NAND2_X1 U8486 ( .A1(n11972), .A2(n11836), .ZN(n11936) );
  AND4_X1 U8487 ( .A1(n7676), .A2(n7675), .A3(n7674), .A4(n7673), .ZN(n11791)
         );
  INV_X1 U8488 ( .A(n12448), .ZN(n12416) );
  NAND2_X1 U8489 ( .A1(n11849), .A2(n11848), .ZN(n11963) );
  AND2_X1 U8490 ( .A1(n6874), .A2(n6879), .ZN(n11575) );
  AND2_X1 U8491 ( .A1(n7812), .A2(n7811), .ZN(n11980) );
  NAND2_X1 U8492 ( .A1(n7835), .A2(n7834), .ZN(n12501) );
  OR2_X1 U8493 ( .A1(n12033), .A2(n13626), .ZN(n7834) );
  INV_X1 U8494 ( .A(n10956), .ZN(n15354) );
  AND2_X1 U8495 ( .A1(n10523), .A2(n10522), .ZN(n11985) );
  AND2_X1 U8496 ( .A1(n6863), .A2(n6862), .ZN(n6861) );
  NAND2_X1 U8497 ( .A1(n11854), .A2(n6864), .ZN(n6863) );
  NAND2_X1 U8498 ( .A1(n6866), .A2(n11885), .ZN(n6862) );
  NAND2_X1 U8499 ( .A1(n11885), .A2(n6657), .ZN(n6864) );
  INV_X1 U8500 ( .A(n6860), .ZN(n6859) );
  OAI21_X1 U8501 ( .B1(n6861), .B2(n6865), .A(n11971), .ZN(n6860) );
  NOR2_X1 U8502 ( .A1(n11885), .A2(n6657), .ZN(n6865) );
  INV_X1 U8503 ( .A(n11858), .ZN(n6856) );
  NAND2_X1 U8504 ( .A1(n10505), .A2(n10574), .ZN(n12014) );
  AND4_X1 U8505 ( .A1(n7725), .A2(n7724), .A3(n7723), .A4(n7722), .ZN(n12606)
         );
  NAND2_X1 U8506 ( .A1(n10828), .A2(n12242), .ZN(n12008) );
  NAND2_X1 U8507 ( .A1(n7892), .A2(n7891), .ZN(n12434) );
  INV_X1 U8508 ( .A(n12606), .ZN(n11982) );
  INV_X1 U8509 ( .A(n11799), .ZN(n12252) );
  INV_X1 U8510 ( .A(n11791), .ZN(n15304) );
  INV_X1 U8511 ( .A(n11727), .ZN(n12253) );
  INV_X1 U8512 ( .A(n11667), .ZN(n12256) );
  OR2_X1 U8513 ( .A1(n7558), .A2(n7509), .ZN(n7510) );
  OR2_X1 U8514 ( .A1(n10513), .A2(n10199), .ZN(n12259) );
  NAND2_X1 U8515 ( .A1(n10788), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10781) );
  OR2_X1 U8516 ( .A1(n10611), .A2(n10781), .ZN(n10613) );
  INV_X1 U8517 ( .A(n11064), .ZN(n15189) );
  INV_X1 U8518 ( .A(n7018), .ZN(n11066) );
  INV_X1 U8519 ( .A(n7020), .ZN(n15241) );
  AOI21_X1 U8520 ( .B1(n15281), .B2(n11115), .A(n11114), .ZN(n11435) );
  NOR2_X1 U8521 ( .A1(n15278), .A2(n11073), .ZN(n11076) );
  XNOR2_X1 U8522 ( .A(n11429), .B(n11447), .ZN(n11522) );
  NOR2_X1 U8523 ( .A1(n7671), .A2(n11522), .ZN(n11521) );
  NAND2_X1 U8524 ( .A1(n10582), .A2(n10581), .ZN(n15300) );
  NOR2_X1 U8525 ( .A1(n12241), .A2(n12259), .ZN(n15285) );
  INV_X1 U8526 ( .A(n12381), .ZN(n6691) );
  OAI21_X1 U8527 ( .B1(n12768), .B2(n12035), .A(n12034), .ZN(n14626) );
  OAI21_X1 U8528 ( .B1(n6775), .B2(n6628), .A(n6772), .ZN(n12397) );
  INV_X1 U8529 ( .A(n7979), .ZN(n6775) );
  INV_X1 U8530 ( .A(n6773), .ZN(n6772) );
  NAND2_X1 U8531 ( .A1(n7056), .A2(n7059), .ZN(n12036) );
  OAI21_X1 U8532 ( .B1(n7419), .B2(n7040), .A(n7038), .ZN(n12454) );
  NAND2_X1 U8533 ( .A1(n12473), .A2(n12071), .ZN(n12452) );
  AND2_X1 U8534 ( .A1(n12450), .A2(n12449), .ZN(n12642) );
  AOI21_X1 U8535 ( .B1(n12470), .B2(n15319), .A(n12469), .ZN(n12471) );
  NAND2_X1 U8536 ( .A1(n7047), .A2(n12173), .ZN(n12530) );
  NAND2_X1 U8537 ( .A1(n7795), .A2(n7048), .ZN(n7047) );
  NAND2_X1 U8538 ( .A1(n7795), .A2(n12161), .ZN(n12541) );
  INV_X1 U8539 ( .A(n15312), .ZN(n14619) );
  NAND2_X1 U8540 ( .A1(n11416), .A2(n12113), .ZN(n11418) );
  NAND2_X1 U8541 ( .A1(n7034), .A2(n12110), .ZN(n11416) );
  NAND2_X2 U8542 ( .A1(n10750), .A2(n15316), .ZN(n15369) );
  INV_X1 U8543 ( .A(n15316), .ZN(n15365) );
  INV_X1 U8544 ( .A(n15356), .ZN(n15363) );
  AND2_X1 U8545 ( .A1(n15369), .A2(n15330), .ZN(n15366) );
  NAND2_X1 U8546 ( .A1(n15333), .A2(n14625), .ZN(n15312) );
  NAND2_X1 U8547 ( .A1(n8836), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n6717) );
  INV_X1 U8548 ( .A(n12202), .ZN(n12711) );
  INV_X1 U8549 ( .A(n11968), .ZN(n12721) );
  NOR2_X1 U8550 ( .A1(n12647), .A2(n12646), .ZN(n12719) );
  AND2_X1 U8551 ( .A1(n12645), .A2(n14640), .ZN(n12646) );
  INV_X1 U8552 ( .A(n11844), .ZN(n12724) );
  INV_X1 U8553 ( .A(n12501), .ZN(n12729) );
  INV_X1 U8554 ( .A(n12514), .ZN(n12733) );
  INV_X1 U8555 ( .A(n11980), .ZN(n12736) );
  INV_X1 U8556 ( .A(n7959), .ZN(n12745) );
  AOI21_X1 U8557 ( .B1(n10357), .B2(n12027), .A(n7762), .ZN(n12749) );
  INV_X1 U8558 ( .A(n11955), .ZN(n12753) );
  INV_X1 U8559 ( .A(n11800), .ZN(n12761) );
  AND2_X1 U8560 ( .A1(n10575), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10039) );
  CLKBUF_X1 U8561 ( .A(n7985), .Z(n11819) );
  NAND2_X1 U8562 ( .A1(n6887), .A2(n6885), .ZN(n12780) );
  AOI21_X1 U8563 ( .B1(n7991), .B2(n6888), .A(n6886), .ZN(n6885) );
  OR3_X1 U8564 ( .A1(n7991), .A2(n6888), .A3(n8002), .ZN(n6887) );
  NOR2_X1 U8565 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_26__SCAN_IN), .ZN(
        n6886) );
  NAND2_X1 U8566 ( .A1(n7997), .A2(n7996), .ZN(n11678) );
  AOI21_X1 U8567 ( .B1(n7995), .B2(P3_IR_REG_25__SCAN_IN), .A(n7994), .ZN(
        n7996) );
  AND2_X1 U8568 ( .A1(n8002), .A2(n7993), .ZN(n7994) );
  NAND2_X1 U8569 ( .A1(n7113), .A2(n7857), .ZN(n7866) );
  NAND2_X1 U8570 ( .A1(n8000), .A2(n7999), .ZN(n11559) );
  INV_X1 U8571 ( .A(n7094), .ZN(n7844) );
  OAI21_X1 U8572 ( .B1(n7833), .B2(n7832), .A(n7097), .ZN(n7094) );
  NAND2_X1 U8573 ( .A1(n7905), .A2(n6557), .ZN(n10965) );
  XNOR2_X1 U8574 ( .A(n7911), .B(n7910), .ZN(n10817) );
  NAND2_X1 U8575 ( .A1(n6793), .A2(n7478), .ZN(n7821) );
  NAND2_X1 U8576 ( .A1(n7810), .A2(n10682), .ZN(n6793) );
  NAND2_X1 U8577 ( .A1(n7082), .A2(n7476), .ZN(n7797) );
  NAND2_X1 U8578 ( .A1(n7784), .A2(n7782), .ZN(n7082) );
  INV_X1 U8579 ( .A(n12375), .ZN(n12391) );
  INV_X1 U8580 ( .A(SI_14_), .ZN(n10120) );
  INV_X1 U8581 ( .A(SI_13_), .ZN(n10029) );
  NAND2_X1 U8582 ( .A1(n7466), .A2(n6795), .ZN(n7706) );
  AND2_X1 U8583 ( .A1(n7466), .A2(n6577), .ZN(n7707) );
  INV_X1 U8584 ( .A(SI_12_), .ZN(n14575) );
  OAI21_X1 U8585 ( .B1(n7681), .B2(n7462), .A(n7461), .ZN(n7696) );
  AND3_X1 U8586 ( .A1(n7629), .A2(n7628), .A3(n7482), .ZN(n7691) );
  NAND2_X1 U8587 ( .A1(n7070), .A2(n7458), .ZN(n7644) );
  NAND2_X1 U8588 ( .A1(n7632), .A2(n7631), .ZN(n7070) );
  AND2_X1 U8589 ( .A1(n7647), .A2(n7677), .ZN(n11135) );
  NAND2_X1 U8590 ( .A1(n7079), .A2(n7453), .ZN(n7578) );
  NAND2_X1 U8591 ( .A1(n7564), .A2(n7563), .ZN(n7079) );
  NAND2_X1 U8592 ( .A1(n7536), .A2(n13570), .ZN(n7549) );
  NAND2_X1 U8593 ( .A1(n7014), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7537) );
  INV_X1 U8594 ( .A(n7536), .ZN(n7014) );
  NAND2_X1 U8595 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7525) );
  NAND2_X1 U8596 ( .A1(n8310), .A2(n8309), .ZN(n10629) );
  AND2_X1 U8597 ( .A1(n8731), .A2(n8712), .ZN(n7128) );
  NAND2_X1 U8598 ( .A1(n12939), .A2(n8712), .ZN(n12783) );
  INV_X1 U8599 ( .A(n10299), .ZN(n8841) );
  NAND2_X1 U8600 ( .A1(n12902), .A2(n8592), .ZN(n12836) );
  NAND2_X1 U8601 ( .A1(n8674), .A2(n8673), .ZN(n13292) );
  NAND2_X1 U8602 ( .A1(n12948), .A2(n8487), .ZN(n12860) );
  NAND2_X1 U8603 ( .A1(n10466), .A2(n10467), .ZN(n10465) );
  INV_X1 U8604 ( .A(n10707), .ZN(n10996) );
  INV_X1 U8605 ( .A(n15043), .ZN(n7131) );
  NAND2_X1 U8606 ( .A1(n11362), .A2(n8424), .ZN(n12907) );
  INV_X1 U8607 ( .A(n12935), .ZN(n12953) );
  NAND2_X1 U8608 ( .A1(n8391), .A2(n8390), .ZN(n15028) );
  INV_X1 U8609 ( .A(n12937), .ZN(n12950) );
  AND2_X1 U8610 ( .A1(n8550), .A2(n8528), .ZN(n7122) );
  NAND2_X1 U8611 ( .A1(n12881), .A2(n8528), .ZN(n12921) );
  OR2_X1 U8612 ( .A1(n8439), .A2(n8438), .ZN(n12975) );
  NAND4_X1 U8613 ( .A1(n8217), .A2(n8216), .A3(n8215), .A4(n8214), .ZN(n12986)
         );
  OR2_X1 U8614 ( .A1(n8212), .A2(n8190), .ZN(n8191) );
  NOR2_X1 U8615 ( .A1(n6923), .A2(n6597), .ZN(n10070) );
  INV_X1 U8616 ( .A(n6922), .ZN(n10138) );
  AND2_X1 U8617 ( .A1(n6920), .A2(n6919), .ZN(n10151) );
  INV_X1 U8618 ( .A(n10124), .ZN(n6919) );
  INV_X1 U8619 ( .A(n6920), .ZN(n10125) );
  NOR2_X1 U8620 ( .A1(n10151), .A2(n6918), .ZN(n10154) );
  AND2_X1 U8621 ( .A1(n10155), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6918) );
  NOR2_X1 U8622 ( .A1(n10540), .A2(n6927), .ZN(n10542) );
  AND2_X1 U8623 ( .A1(n10541), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U8624 ( .A1(n10542), .A2(n10543), .ZN(n10795) );
  NAND2_X1 U8625 ( .A1(n10072), .A2(n13385), .ZN(n15001) );
  NOR2_X1 U8626 ( .A1(n13040), .A2(n13039), .ZN(n13042) );
  AND2_X1 U8627 ( .A1(n10072), .A2(n10071), .ZN(n15009) );
  NAND2_X1 U8628 ( .A1(n7194), .A2(n15021), .ZN(n13264) );
  XNOR2_X1 U8629 ( .A(n13057), .B(n7195), .ZN(n7194) );
  AND2_X1 U8630 ( .A1(n13066), .A2(n13065), .ZN(n13276) );
  NAND2_X1 U8631 ( .A1(n13094), .A2(n13105), .ZN(n13093) );
  AND2_X1 U8632 ( .A1(n7165), .A2(n6590), .ZN(n13130) );
  OAI21_X1 U8633 ( .B1(n6714), .B2(n6981), .A(n6575), .ZN(n13124) );
  NAND2_X1 U8634 ( .A1(n6978), .A2(n6982), .ZN(n13125) );
  NAND2_X1 U8635 ( .A1(n8871), .A2(n8870), .ZN(n13150) );
  NAND2_X1 U8636 ( .A1(n6714), .A2(n8938), .ZN(n13142) );
  NAND2_X1 U8637 ( .A1(n13186), .A2(n8934), .ZN(n13179) );
  NAND2_X1 U8638 ( .A1(n7158), .A2(n9809), .ZN(n13185) );
  NAND2_X1 U8639 ( .A1(n13199), .A2(n9808), .ZN(n7158) );
  OAI21_X1 U8640 ( .B1(n13239), .B2(n6658), .A(n8927), .ZN(n13212) );
  AND2_X1 U8641 ( .A1(n8513), .A2(n8512), .ZN(n13237) );
  NAND2_X1 U8642 ( .A1(n8862), .A2(n7149), .ZN(n7144) );
  NAND2_X1 U8643 ( .A1(n8862), .A2(n8861), .ZN(n11476) );
  NAND2_X1 U8644 ( .A1(n10846), .A2(n8913), .ZN(n6964) );
  NAND2_X1 U8645 ( .A1(n13247), .A2(n8908), .ZN(n10656) );
  NAND2_X1 U8646 ( .A1(n15104), .A2(n8852), .ZN(n10654) );
  INV_X1 U8647 ( .A(n15023), .ZN(n13259) );
  NAND2_X1 U8648 ( .A1(n8210), .A2(n8209), .ZN(n10756) );
  NAND2_X1 U8649 ( .A1(n13264), .A2(n7192), .ZN(n13353) );
  INV_X1 U8650 ( .A(n7193), .ZN(n7192) );
  OAI21_X1 U8651 ( .B1(n7195), .B2(n15146), .A(n13265), .ZN(n7193) );
  AND3_X1 U8652 ( .A1(n13283), .A2(n13282), .A3(n13281), .ZN(n13284) );
  INV_X2 U8653 ( .A(n15153), .ZN(n15155) );
  CLKBUF_X1 U8654 ( .A(n15079), .Z(n15083) );
  AND2_X1 U8655 ( .A1(n8802), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15088) );
  AND2_X1 U8656 ( .A1(n7400), .A2(n7401), .ZN(n7399) );
  AND2_X1 U8657 ( .A1(n7435), .A2(n8178), .ZN(n7400) );
  INV_X1 U8658 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13488) );
  XNOR2_X1 U8659 ( .A(n8759), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13387) );
  NAND2_X1 U8660 ( .A1(n8758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8759) );
  AND2_X1 U8661 ( .A1(n8756), .A2(n8755), .ZN(n11738) );
  INV_X1 U8662 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11056) );
  NOR2_X1 U8663 ( .A1(n8156), .A2(n8157), .ZN(n8158) );
  NOR2_X1 U8664 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n8157) );
  INV_X1 U8665 ( .A(n9844), .ZN(n13047) );
  INV_X1 U8666 ( .A(n11648), .ZN(n15013) );
  INV_X1 U8667 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n13634) );
  INV_X1 U8668 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10174) );
  INV_X1 U8669 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10053) );
  INV_X1 U8670 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10002) );
  NOR2_X1 U8671 ( .A1(n8205), .A2(n8333), .ZN(n8228) );
  NAND2_X1 U8672 ( .A1(n13861), .A2(n13862), .ZN(n6743) );
  NAND2_X1 U8673 ( .A1(n6748), .A2(n13725), .ZN(n13788) );
  NAND2_X1 U8674 ( .A1(n6748), .A2(n6746), .ZN(n13789) );
  NAND2_X1 U8675 ( .A1(n7370), .A2(n7368), .ZN(n7367) );
  AND2_X1 U8676 ( .A1(n7348), .A2(n7349), .ZN(n11179) );
  AND2_X1 U8677 ( .A1(n9870), .A2(n9869), .ZN(n10424) );
  XNOR2_X1 U8678 ( .A(n7341), .B(n9871), .ZN(n10423) );
  NAND2_X1 U8679 ( .A1(n13853), .A2(n13733), .ZN(n13810) );
  NAND2_X1 U8680 ( .A1(n6724), .A2(n7350), .ZN(n13818) );
  AOI21_X1 U8681 ( .B1(n7352), .B2(n7354), .A(n6611), .ZN(n7350) );
  NAND2_X1 U8682 ( .A1(n13779), .A2(n7352), .ZN(n6724) );
  AND2_X1 U8683 ( .A1(n7361), .A2(n7362), .ZN(n13828) );
  NAND2_X1 U8684 ( .A1(n13827), .A2(n13711), .ZN(n13839) );
  NAND2_X1 U8685 ( .A1(n9316), .A2(n9315), .ZN(n14310) );
  NAND2_X1 U8686 ( .A1(n7351), .A2(n13752), .ZN(n13845) );
  NAND2_X1 U8687 ( .A1(n13779), .A2(n13780), .ZN(n7351) );
  AND2_X1 U8688 ( .A1(n11209), .A2(n7343), .ZN(n7342) );
  NAND3_X1 U8689 ( .A1(n6733), .A2(n6732), .A3(n6737), .ZN(n6728) );
  AND2_X1 U8690 ( .A1(n10452), .A2(n10315), .ZN(n14733) );
  NAND2_X1 U8691 ( .A1(n7357), .A2(n7358), .ZN(n7356) );
  INV_X1 U8692 ( .A(n13908), .ZN(n14726) );
  INV_X1 U8693 ( .A(n10874), .ZN(n13921) );
  CLKBUF_X1 U8694 ( .A(n9859), .Z(n13922) );
  INV_X1 U8695 ( .A(n9939), .ZN(n9943) );
  XNOR2_X1 U8696 ( .A(n13928), .B(n6852), .ZN(n13925) );
  XNOR2_X1 U8697 ( .A(n6853), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13928) );
  NAND2_X1 U8698 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6853) );
  NAND2_X1 U8699 ( .A1(n13968), .A2(n6664), .ZN(n10110) );
  NAND2_X1 U8700 ( .A1(n10110), .A2(n10109), .ZN(n10253) );
  INV_X1 U8701 ( .A(n6846), .ZN(n10281) );
  AND2_X1 U8702 ( .A1(n6846), .A2(n6845), .ZN(n10283) );
  NAND2_X1 U8703 ( .A1(n10282), .A2(n14933), .ZN(n6845) );
  INV_X1 U8704 ( .A(n6844), .ZN(n10370) );
  AND2_X1 U8705 ( .A1(n6844), .A2(n6843), .ZN(n13981) );
  NAND2_X1 U8706 ( .A1(n10375), .A2(n14935), .ZN(n6843) );
  OAI21_X1 U8707 ( .B1(n14747), .B2(n14742), .A(n10557), .ZN(n14745) );
  NOR2_X1 U8708 ( .A1(n10371), .A2(n10372), .ZN(n14747) );
  NAND2_X1 U8709 ( .A1(n14745), .A2(n6838), .ZN(n10560) );
  OR2_X1 U8710 ( .A1(n14751), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6838) );
  INV_X1 U8711 ( .A(n6841), .ZN(n13998) );
  NOR2_X1 U8712 ( .A1(n10111), .A2(n10235), .ZN(n14750) );
  OAI21_X1 U8713 ( .B1(n14756), .B2(n14043), .A(n14042), .ZN(n6851) );
  AND2_X1 U8714 ( .A1(n9493), .A2(n9492), .ZN(n14328) );
  NAND2_X1 U8715 ( .A1(n14164), .A2(n7251), .ZN(n14151) );
  NOR2_X1 U8716 ( .A1(n7224), .A2(n7228), .ZN(n14141) );
  AND2_X1 U8717 ( .A1(n14161), .A2(n14160), .ZN(n14353) );
  NAND2_X1 U8718 ( .A1(n7241), .A2(n7240), .ZN(n14173) );
  AND2_X1 U8719 ( .A1(n7241), .A2(n6582), .ZN(n14174) );
  NAND2_X1 U8720 ( .A1(n6576), .A2(n7242), .ZN(n7241) );
  AND2_X1 U8721 ( .A1(n6576), .A2(n14078), .ZN(n14190) );
  AOI21_X1 U8722 ( .B1(n14237), .B2(n14236), .A(n14096), .ZN(n14223) );
  CLKBUF_X1 U8723 ( .A(n14219), .Z(n14220) );
  NAND2_X1 U8724 ( .A1(n14263), .A2(n14072), .ZN(n14235) );
  AND2_X1 U8725 ( .A1(n7215), .A2(n7218), .ZN(n14251) );
  NAND2_X1 U8726 ( .A1(n14092), .A2(n14091), .ZN(n14270) );
  NAND2_X1 U8727 ( .A1(n6940), .A2(n14087), .ZN(n14304) );
  NAND2_X1 U8728 ( .A1(n11621), .A2(n11620), .ZN(n14084) );
  NOR2_X1 U8729 ( .A1(n11583), .A2(n7254), .ZN(n7253) );
  INV_X1 U8730 ( .A(n11295), .ZN(n7254) );
  NAND2_X1 U8731 ( .A1(n7255), .A2(n11295), .ZN(n11296) );
  NAND2_X1 U8732 ( .A1(n10976), .A2(n11014), .ZN(n7234) );
  NAND2_X1 U8733 ( .A1(n10912), .A2(n10916), .ZN(n7246) );
  NAND2_X1 U8734 ( .A1(n14804), .A2(n10871), .ZN(n10873) );
  INV_X1 U8735 ( .A(n14308), .ZN(n14818) );
  OR2_X1 U8736 ( .A1(n10316), .A2(n10036), .ZN(n14775) );
  OR2_X1 U8737 ( .A1(n14833), .A2(n9953), .ZN(n14808) );
  NOR2_X1 U8738 ( .A1(n14833), .A2(n14802), .ZN(n14829) );
  INV_X1 U8739 ( .A(n14940), .ZN(n14937) );
  NAND2_X1 U8740 ( .A1(n14336), .A2(n14766), .ZN(n6837) );
  INV_X1 U8741 ( .A(n14925), .ZN(n14924) );
  INV_X1 U8742 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n14450) );
  NAND2_X1 U8743 ( .A1(n8990), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n8994) );
  NOR2_X1 U8744 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n8991) );
  NAND2_X1 U8745 ( .A1(n7336), .A2(n8133), .ZN(n8881) );
  NAND2_X1 U8746 ( .A1(n8692), .A2(n7339), .ZN(n7336) );
  INV_X1 U8747 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9582) );
  INV_X1 U8748 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11741) );
  XNOR2_X1 U8749 ( .A(n9585), .B(n9584), .ZN(n11743) );
  NOR2_X1 U8750 ( .A1(n10030), .A2(P1_U3086), .ZN(n11379) );
  NAND2_X1 U8751 ( .A1(n7332), .A2(n8111), .ZN(n8577) );
  INV_X1 U8752 ( .A(n7333), .ZN(n7332) );
  NAND2_X1 U8753 ( .A1(n6911), .A2(n8553), .ZN(n10538) );
  NAND2_X1 U8754 ( .A1(n8532), .A2(n8531), .ZN(n6911) );
  INV_X1 U8755 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10443) );
  INV_X1 U8756 ( .A(n11321), .ZN(n11313) );
  INV_X1 U8757 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10386) );
  INV_X1 U8758 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10051) );
  INV_X1 U8759 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10017) );
  INV_X1 U8760 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10004) );
  INV_X1 U8761 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10000) );
  INV_X1 U8762 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14507) );
  XNOR2_X1 U8763 ( .A(n14508), .B(n6764), .ZN(n15437) );
  INV_X1 U8764 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6764) );
  XNOR2_X1 U8765 ( .A(n14512), .B(n6762), .ZN(n14570) );
  INV_X1 U8766 ( .A(n14513), .ZN(n6762) );
  NAND2_X1 U8767 ( .A1(n6757), .A2(n6755), .ZN(n15427) );
  XNOR2_X1 U8768 ( .A(n14533), .B(n7176), .ZN(n15430) );
  INV_X1 U8769 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7176) );
  XNOR2_X1 U8770 ( .A(n14535), .B(n14536), .ZN(n14591) );
  XNOR2_X1 U8771 ( .A(n14541), .B(n14540), .ZN(n14592) );
  INV_X1 U8772 ( .A(n14539), .ZN(n14540) );
  OAI21_X1 U8773 ( .B1(n14545), .B2(n14702), .A(n14699), .ZN(n14705) );
  XNOR2_X1 U8774 ( .A(n14555), .B(n14554), .ZN(n14720) );
  OAI211_X1 U8775 ( .C1(n11947), .C2(n6858), .A(n6857), .B(n6855), .ZN(
        P3_U3180) );
  NAND2_X1 U8776 ( .A1(n6574), .A2(n11971), .ZN(n6858) );
  AOI21_X1 U8777 ( .B1(n6859), .B2(n6861), .A(n6856), .ZN(n6855) );
  NAND2_X1 U8778 ( .A1(n11947), .A2(n6859), .ZN(n6857) );
  NAND2_X1 U8779 ( .A1(n6718), .A2(n6715), .ZN(P3_U3487) );
  INV_X1 U8780 ( .A(n6716), .ZN(n6715) );
  NAND2_X1 U8781 ( .A1(n12627), .A2(n15424), .ZN(n6718) );
  OAI21_X1 U8782 ( .B1(n12628), .B2(n12694), .A(n6717), .ZN(n6716) );
  INV_X1 U8783 ( .A(n8037), .ZN(n8038) );
  OAI21_X1 U8784 ( .B1(n12628), .B2(n12762), .A(n8036), .ZN(n8037) );
  AND2_X1 U8785 ( .A1(n13274), .A2(n12946), .ZN(n7119) );
  NAND2_X1 U8786 ( .A1(n7121), .A2(n8246), .ZN(n10363) );
  NOR2_X1 U8787 ( .A1(n6923), .A2(n14971), .ZN(n14975) );
  INV_X1 U8788 ( .A(n7189), .ZN(P2_U3498) );
  AOI21_X1 U8789 ( .B1(n13353), .B2(n15155), .A(n7190), .ZN(n7189) );
  NOR2_X1 U8790 ( .A1(n15155), .A2(n7191), .ZN(n7190) );
  INV_X1 U8791 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7191) );
  XNOR2_X1 U8792 ( .A(n6726), .B(n6725), .ZN(n13778) );
  NOR2_X1 U8793 ( .A1(n6893), .A2(n9576), .ZN(n6889) );
  OAI211_X1 U8794 ( .C1(n14040), .C2(n14039), .A(n6850), .B(n6847), .ZN(
        P1_U3262) );
  INV_X1 U8795 ( .A(n6851), .ZN(n6850) );
  NAND2_X1 U8796 ( .A1(n6848), .A2(n14039), .ZN(n6847) );
  NOR2_X1 U8797 ( .A1(n14710), .A2(n14711), .ZN(n14709) );
  NOR2_X1 U8798 ( .A1(n14718), .A2(n14717), .ZN(n14716) );
  AND2_X1 U8799 ( .A1(n7188), .A2(n7187), .ZN(n14718) );
  XNOR2_X1 U8800 ( .A(n6753), .B(n6586), .ZN(SUB_1596_U4) );
  OAI21_X1 U8801 ( .B1(n14604), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n6559), .ZN(
        n6753) );
  OR3_X1 U8802 ( .A1(n7908), .A2(P3_IR_REG_22__SCAN_IN), .A3(
        P3_IR_REG_21__SCAN_IN), .ZN(n6557) );
  INV_X1 U8803 ( .A(n7230), .ZN(n14155) );
  INV_X1 U8804 ( .A(n12413), .ZN(n7062) );
  NAND2_X1 U8805 ( .A1(n13897), .A2(n13898), .ZN(n7361) );
  OR2_X1 U8806 ( .A1(n13302), .A2(n12885), .ZN(n6558) );
  INV_X1 U8807 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14441) );
  INV_X1 U8808 ( .A(n9894), .ZN(n7379) );
  OR2_X1 U8809 ( .A1(n14606), .A2(n14605), .ZN(n6559) );
  AND2_X1 U8810 ( .A1(n6954), .A2(n14912), .ZN(n6560) );
  INV_X1 U8811 ( .A(n13906), .ZN(n6955) );
  INV_X1 U8812 ( .A(n7072), .ZN(n7071) );
  OAI21_X1 U8813 ( .B1(n7631), .B2(n7073), .A(n7642), .ZN(n7072) );
  AND2_X1 U8814 ( .A1(n7104), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n6561) );
  OR2_X1 U8815 ( .A1(n6780), .A2(n15347), .ZN(n6562) );
  INV_X1 U8816 ( .A(n13882), .ZN(n6749) );
  AND2_X1 U8817 ( .A1(n14356), .A2(n14159), .ZN(n6563) );
  INV_X2 U8818 ( .A(n9960), .ZN(n9367) );
  OR2_X1 U8819 ( .A1(n14563), .A2(n14562), .ZN(n6564) );
  OR2_X1 U8820 ( .A1(n7073), .A2(n7069), .ZN(n6565) );
  OR2_X1 U8821 ( .A1(n7908), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n6566) );
  NAND2_X1 U8822 ( .A1(n14717), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n6567) );
  OR2_X1 U8823 ( .A1(n14706), .A2(n14705), .ZN(n6568) );
  NAND2_X1 U8824 ( .A1(n9359), .A2(n7282), .ZN(n6569) );
  AND2_X1 U8825 ( .A1(n6777), .A2(n6776), .ZN(n6571) );
  OAI21_X1 U8826 ( .B1(n6949), .B2(n6948), .A(n14100), .ZN(n6947) );
  AND2_X1 U8827 ( .A1(n7203), .A2(n7202), .ZN(n6572) );
  AND2_X1 U8828 ( .A1(n6640), .A2(n7050), .ZN(n6573) );
  NAND2_X1 U8829 ( .A1(n9386), .A2(n9385), .ZN(n14198) );
  INV_X1 U8830 ( .A(n14198), .ZN(n6959) );
  NAND2_X1 U8831 ( .A1(n6743), .A2(n6742), .ZN(n14656) );
  AND2_X1 U8832 ( .A1(n11854), .A2(n11885), .ZN(n6574) );
  INV_X1 U8833 ( .A(n12319), .ZN(n14585) );
  INV_X1 U8834 ( .A(n6670), .ZN(n7097) );
  CLKBUF_X3 U8835 ( .A(n9784), .Z(n9779) );
  AND2_X1 U8836 ( .A1(n13126), .A2(n6979), .ZN(n6575) );
  OR2_X1 U8837 ( .A1(n14203), .A2(n14207), .ZN(n6576) );
  AND2_X1 U8838 ( .A1(n7100), .A2(n7101), .ZN(n6577) );
  INV_X1 U8839 ( .A(n7157), .ZN(n7156) );
  NAND2_X1 U8840 ( .A1(n9809), .A2(n6591), .ZN(n7157) );
  NAND2_X1 U8841 ( .A1(n13348), .A2(n11348), .ZN(n6578) );
  AND2_X1 U8842 ( .A1(n7425), .A2(n7313), .ZN(n6579) );
  NAND2_X1 U8843 ( .A1(n12069), .A2(n12071), .ZN(n7965) );
  INV_X1 U8844 ( .A(n7965), .ZN(n12474) );
  INV_X2 U8845 ( .A(n9960), .ZN(n9981) );
  NAND4_X1 U8846 ( .A1(n8989), .A2(n8988), .A3(n8987), .A4(n8986), .ZN(n9859)
         );
  INV_X1 U8847 ( .A(n12205), .ZN(n6779) );
  AND2_X1 U8848 ( .A1(n14167), .A2(n14101), .ZN(n6580) );
  NAND2_X1 U8849 ( .A1(n13690), .A2(n13689), .ZN(n6581) );
  OR2_X1 U8850 ( .A1(n14198), .A2(n14079), .ZN(n6582) );
  OAI21_X1 U8851 ( .B1(n7598), .B2(n7455), .A(n7454), .ZN(n7610) );
  INV_X1 U8852 ( .A(n7060), .ZN(n7059) );
  OAI21_X1 U8853 ( .B1(n12212), .B2(n7065), .A(n12209), .ZN(n7060) );
  INV_X1 U8854 ( .A(n11129), .ZN(n15231) );
  INV_X1 U8855 ( .A(n13287), .ZN(n13103) );
  OAI21_X1 U8856 ( .B1(n13199), .B2(n7157), .A(n7154), .ZN(n13170) );
  AND2_X1 U8857 ( .A1(n6914), .A2(n6913), .ZN(n8311) );
  AND2_X1 U8858 ( .A1(n7314), .A2(n7313), .ZN(n6583) );
  XNOR2_X1 U8859 ( .A(n13801), .B(n13800), .ZN(n6584) );
  AND2_X1 U8860 ( .A1(n13112), .A2(n7205), .ZN(n6585) );
  XOR2_X1 U8861 ( .A(n14613), .B(n14612), .Z(n6586) );
  INV_X1 U8862 ( .A(n9800), .ZN(n7195) );
  INV_X1 U8863 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n8178) );
  AND4_X2 U8864 ( .A1(n7520), .A2(n7519), .A3(n7518), .A4(n7517), .ZN(n15341)
         );
  NOR2_X1 U8865 ( .A1(n7798), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n6883) );
  AND2_X1 U8866 ( .A1(n15195), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n6587) );
  AND2_X1 U8867 ( .A1(n13302), .A2(n12885), .ZN(n6588) );
  OR2_X1 U8868 ( .A1(n14536), .A2(n14535), .ZN(n6589) );
  OR2_X1 U8869 ( .A1(n13302), .A2(n12913), .ZN(n6590) );
  INV_X1 U8870 ( .A(n9630), .ZN(n7406) );
  OR2_X1 U8871 ( .A1(n13318), .A2(n12968), .ZN(n6591) );
  OR2_X1 U8872 ( .A1(n11391), .A2(n11390), .ZN(n6592) );
  NAND2_X1 U8873 ( .A1(n12218), .A2(n12226), .ZN(n12217) );
  AND2_X1 U8874 ( .A1(n6888), .A2(n7492), .ZN(n6593) );
  XNOR2_X1 U8875 ( .A(n13280), .B(n8944), .ZN(n9807) );
  INV_X1 U8876 ( .A(n14347), .ZN(n14167) );
  NAND2_X1 U8877 ( .A1(n9419), .A2(n9418), .ZN(n14347) );
  NAND2_X1 U8878 ( .A1(n8152), .A2(n8151), .ZN(n13274) );
  NAND2_X1 U8879 ( .A1(n9033), .A2(n8963), .ZN(n9053) );
  OR2_X1 U8880 ( .A1(n11131), .A2(n11068), .ZN(n6594) );
  NOR2_X1 U8881 ( .A1(n12286), .A2(n12285), .ZN(n6595) );
  AND2_X1 U8882 ( .A1(n6936), .A2(n6935), .ZN(n6596) );
  AND2_X1 U8883 ( .A1(n10076), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6597) );
  INV_X1 U8884 ( .A(n6950), .ZN(n6949) );
  NOR2_X1 U8885 ( .A1(n14175), .A2(n6951), .ZN(n6950) );
  AND2_X1 U8886 ( .A1(n8487), .A2(n8502), .ZN(n6598) );
  OR2_X1 U8887 ( .A1(n11125), .A2(n11083), .ZN(n6599) );
  INV_X1 U8888 ( .A(n6961), .ZN(n14238) );
  NOR2_X1 U8889 ( .A1(n14255), .A2(n14381), .ZN(n6961) );
  AND2_X1 U8890 ( .A1(n8329), .A2(n8337), .ZN(n6600) );
  AND2_X1 U8891 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n6601) );
  INV_X1 U8892 ( .A(n11564), .ZN(n12108) );
  NOR2_X1 U8893 ( .A1(n8533), .A2(n8145), .ZN(n8156) );
  AND2_X1 U8894 ( .A1(n9471), .A2(n9470), .ZN(n14333) );
  AND2_X1 U8895 ( .A1(n11620), .A2(n6941), .ZN(n6602) );
  NAND2_X1 U8896 ( .A1(n13344), .A2(n12974), .ZN(n6603) );
  AND2_X1 U8897 ( .A1(n6867), .A2(n11836), .ZN(n6604) );
  INV_X1 U8898 ( .A(n9662), .ZN(n7412) );
  INV_X1 U8899 ( .A(n7126), .ZN(n7125) );
  NAND2_X1 U8900 ( .A1(n11049), .A2(n8364), .ZN(n7126) );
  INV_X1 U8901 ( .A(n7243), .ZN(n7242) );
  NAND2_X1 U8902 ( .A1(n14193), .A2(n14078), .ZN(n7243) );
  AND2_X1 U8903 ( .A1(n10272), .A2(n10106), .ZN(n6605) );
  AND2_X1 U8904 ( .A1(n15136), .A2(n11329), .ZN(n6606) );
  INV_X1 U8905 ( .A(n9739), .ZN(n7409) );
  AND2_X1 U8906 ( .A1(n14121), .A2(n7249), .ZN(n6607) );
  NOR2_X1 U8907 ( .A1(n14650), .A2(n12975), .ZN(n6608) );
  INV_X1 U8908 ( .A(n6737), .ZN(n6736) );
  NAND2_X1 U8909 ( .A1(n7375), .A2(n6738), .ZN(n6737) );
  INV_X1 U8910 ( .A(n7252), .ZN(n7251) );
  AND2_X1 U8911 ( .A1(n13312), .A2(n8935), .ZN(n6609) );
  AND2_X1 U8912 ( .A1(n8997), .A2(n9960), .ZN(n6610) );
  AND2_X1 U8913 ( .A1(n13758), .A2(n13757), .ZN(n6611) );
  INV_X1 U8914 ( .A(n14268), .ZN(n14269) );
  INV_X1 U8915 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7492) );
  AND2_X1 U8916 ( .A1(n14263), .A2(n7258), .ZN(n6612) );
  INV_X1 U8917 ( .A(n6722), .ZN(n6952) );
  OR2_X1 U8918 ( .A1(n14192), .A2(n14193), .ZN(n6722) );
  NOR2_X1 U8919 ( .A1(n14917), .A2(n13915), .ZN(n6613) );
  NOR2_X1 U8920 ( .A1(n12438), .A2(n12448), .ZN(n6614) );
  NOR2_X1 U8921 ( .A1(n13312), .A2(n8935), .ZN(n6615) );
  INV_X1 U8922 ( .A(n7429), .ZN(n7163) );
  INV_X1 U8923 ( .A(n9301), .ZN(n7273) );
  INV_X1 U8924 ( .A(n10973), .ZN(n14763) );
  AND2_X1 U8925 ( .A1(n13302), .A2(n12913), .ZN(n6616) );
  NAND2_X1 U8926 ( .A1(n6783), .A2(n12205), .ZN(n6617) );
  INV_X1 U8927 ( .A(n7229), .ZN(n7228) );
  NAND2_X1 U8928 ( .A1(n14347), .A2(n14102), .ZN(n7229) );
  NAND2_X1 U8929 ( .A1(n7135), .A2(n8332), .ZN(n8533) );
  INV_X1 U8930 ( .A(n8533), .ZN(n6688) );
  NOR2_X1 U8931 ( .A1(n9682), .A2(n7390), .ZN(n6618) );
  OR2_X1 U8932 ( .A1(n7136), .A2(n14947), .ZN(n6619) );
  INV_X1 U8933 ( .A(n9212), .ZN(n7287) );
  AND2_X1 U8934 ( .A1(n7268), .A2(n7267), .ZN(n9033) );
  INV_X1 U8935 ( .A(n9821), .ZN(n11536) );
  AND2_X1 U8936 ( .A1(n8070), .A2(SI_9_), .ZN(n6620) );
  AND2_X1 U8937 ( .A1(n13287), .A2(n12963), .ZN(n6621) );
  INV_X1 U8938 ( .A(n9173), .ZN(n7290) );
  AND2_X1 U8939 ( .A1(n9372), .A2(n6902), .ZN(n6622) );
  INV_X1 U8940 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7488) );
  OR2_X1 U8941 ( .A1(n6884), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n6623) );
  INV_X1 U8942 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n6888) );
  INV_X1 U8943 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7498) );
  AND2_X1 U8944 ( .A1(n7225), .A2(n7222), .ZN(n6624) );
  INV_X1 U8945 ( .A(n7259), .ZN(n7258) );
  NAND2_X1 U8946 ( .A1(n7260), .A2(n14072), .ZN(n7259) );
  NAND2_X1 U8947 ( .A1(n7160), .A2(n7163), .ZN(n6625) );
  AND2_X1 U8948 ( .A1(n9996), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6626) );
  INV_X1 U8949 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9584) );
  NOR2_X1 U8950 ( .A1(n9683), .A2(n9684), .ZN(n6627) );
  OR2_X1 U8951 ( .A1(n6617), .A2(n15347), .ZN(n6628) );
  INV_X1 U8952 ( .A(n12407), .ZN(n12628) );
  NAND2_X1 U8953 ( .A1(n7898), .A2(n7897), .ZN(n12407) );
  OR2_X1 U8954 ( .A1(n8469), .A2(n8095), .ZN(n6629) );
  AND2_X1 U8955 ( .A1(n13726), .A2(n6751), .ZN(n6630) );
  NAND2_X1 U8956 ( .A1(n6883), .A2(n7488), .ZN(n7908) );
  AND2_X1 U8957 ( .A1(n13796), .A2(n13795), .ZN(n6631) );
  AND2_X1 U8958 ( .A1(n13829), .A2(n13837), .ZN(n6632) );
  INV_X1 U8959 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7489) );
  INV_X1 U8960 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U8961 ( .A1(n8876), .A2(n8875), .ZN(n13104) );
  NOR2_X1 U8962 ( .A1(n14788), .A2(n13917), .ZN(n6633) );
  AND2_X1 U8963 ( .A1(n7265), .A2(n7263), .ZN(n6634) );
  NOR2_X1 U8964 ( .A1(n13787), .A2(n6747), .ZN(n6746) );
  INV_X1 U8965 ( .A(n8852), .ZN(n7171) );
  NAND2_X1 U8966 ( .A1(n9014), .A2(n9013), .ZN(n10684) );
  AND2_X1 U8967 ( .A1(n8304), .A2(n8289), .ZN(n6635) );
  AND2_X1 U8968 ( .A1(n8608), .A2(n8592), .ZN(n6636) );
  OR2_X1 U8969 ( .A1(n7412), .A2(n9661), .ZN(n6637) );
  OR2_X1 U8970 ( .A1(n9652), .A2(n9650), .ZN(n6638) );
  OR2_X1 U8971 ( .A1(n9728), .A2(n9726), .ZN(n6639) );
  AND2_X1 U8972 ( .A1(n7487), .A2(n6880), .ZN(n6640) );
  OR2_X1 U8973 ( .A1(n9750), .A2(n9748), .ZN(n6641) );
  OR2_X1 U8974 ( .A1(n7406), .A2(n9629), .ZN(n6642) );
  OR2_X1 U8975 ( .A1(n9738), .A2(n7409), .ZN(n6643) );
  OR2_X1 U8976 ( .A1(n9715), .A2(n9717), .ZN(n6644) );
  OR2_X1 U8977 ( .A1(n9639), .A2(n9641), .ZN(n6645) );
  OR2_X1 U8978 ( .A1(n9671), .A2(n9673), .ZN(n6646) );
  AND2_X1 U8979 ( .A1(n6561), .A2(n7459), .ZN(n6647) );
  OR2_X1 U8980 ( .A1(n7403), .A2(n9672), .ZN(n6648) );
  OR2_X1 U8981 ( .A1(n9211), .A2(n7287), .ZN(n6649) );
  OR2_X1 U8982 ( .A1(n9172), .A2(n7290), .ZN(n6650) );
  INV_X1 U8983 ( .A(n12207), .ZN(n7065) );
  OR2_X1 U8984 ( .A1(n6952), .A2(n6949), .ZN(n6651) );
  INV_X1 U8985 ( .A(n9139), .ZN(n7294) );
  NAND2_X1 U8986 ( .A1(n9415), .A2(n7284), .ZN(n6652) );
  INV_X1 U8987 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U8988 ( .A1(n9300), .A2(n7273), .ZN(n6653) );
  INV_X1 U8989 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6687) );
  OR2_X1 U8990 ( .A1(n14222), .A2(n6931), .ZN(n6654) );
  NOR2_X1 U8991 ( .A1(n12202), .A2(n12434), .ZN(n6655) );
  NAND2_X1 U8992 ( .A1(n13701), .A2(n13702), .ZN(n7362) );
  AND2_X1 U8993 ( .A1(n6877), .A2(n6592), .ZN(n6656) );
  NAND2_X1 U8994 ( .A1(n11946), .A2(n11882), .ZN(n6657) );
  INV_X1 U8995 ( .A(n7588), .ZN(n7604) );
  NOR2_X1 U8996 ( .A1(n13237), .A2(n12971), .ZN(n6658) );
  AND2_X1 U8997 ( .A1(n14375), .A2(n14241), .ZN(n6659) );
  NOR2_X1 U8998 ( .A1(n12608), .A2(n12617), .ZN(n6660) );
  XNOR2_X1 U8999 ( .A(n13700), .B(n13702), .ZN(n13897) );
  OAI21_X1 U9000 ( .B1(n7795), .B2(n7044), .A(n7041), .ZN(n12515) );
  NAND2_X1 U9001 ( .A1(n6963), .A2(n6962), .ZN(n15015) );
  NAND2_X1 U9002 ( .A1(n6964), .A2(n8914), .ZN(n10835) );
  NAND2_X1 U9003 ( .A1(n7144), .A2(n7148), .ZN(n11535) );
  NAND2_X1 U9004 ( .A1(n11989), .A2(n7444), .ZN(n11804) );
  AND2_X1 U9005 ( .A1(n14459), .A2(n10033), .ZN(n14375) );
  INV_X1 U9006 ( .A(n14375), .ZN(n14231) );
  INV_X1 U9007 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7268) );
  INV_X1 U9008 ( .A(n12540), .ZN(n7961) );
  AND2_X1 U9009 ( .A1(n11824), .A2(n12606), .ZN(n6661) );
  AND2_X1 U9010 ( .A1(n13318), .A2(n12968), .ZN(n6662) );
  INV_X1 U9011 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6852) );
  AND2_X1 U9012 ( .A1(n7362), .A2(n13829), .ZN(n6663) );
  OR2_X1 U9013 ( .A1(n13965), .A2(n10108), .ZN(n6664) );
  OR2_X1 U9014 ( .A1(n13983), .A2(n14938), .ZN(n6665) );
  INV_X1 U9015 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n13631) );
  INV_X1 U9016 ( .A(n11428), .ZN(n7013) );
  AND2_X1 U9017 ( .A1(n11443), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n11428) );
  AND2_X1 U9018 ( .A1(n10020), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n6666) );
  INV_X1 U9019 ( .A(n6960), .ZN(n14209) );
  NOR2_X1 U9020 ( .A1(n14227), .A2(n14369), .ZN(n6960) );
  NAND2_X1 U9021 ( .A1(n8886), .A2(n8885), .ZN(n13270) );
  INV_X1 U9022 ( .A(n13270), .ZN(n7202) );
  AND2_X1 U9023 ( .A1(n7358), .A2(n13898), .ZN(n6667) );
  NAND2_X1 U9024 ( .A1(n7026), .A2(n7536), .ZN(n7627) );
  AND2_X1 U9025 ( .A1(n13735), .A2(n13733), .ZN(n6668) );
  AND2_X1 U9026 ( .A1(n6743), .A2(n6581), .ZN(n6669) );
  INV_X1 U9027 ( .A(n7416), .ZN(n7218) );
  AND2_X1 U9028 ( .A1(n6556), .A2(n9844), .ZN(n9774) );
  AND2_X1 U9029 ( .A1(n11056), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6670) );
  INV_X1 U9030 ( .A(n12273), .ZN(n6802) );
  NAND2_X1 U9031 ( .A1(n6875), .A2(n6874), .ZN(n11636) );
  XOR2_X1 U9032 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .Z(n6671) );
  XNOR2_X1 U9033 ( .A(n9588), .B(n9587), .ZN(n9903) );
  NAND2_X1 U9034 ( .A1(n8451), .A2(n8450), .ZN(n13344) );
  INV_X1 U9035 ( .A(n13344), .ZN(n7207) );
  OAI21_X1 U9036 ( .B1(n10669), .B2(n7376), .A(n7375), .ZN(n10928) );
  NAND2_X1 U9037 ( .A1(n10465), .A2(n8289), .ZN(n10478) );
  NOR2_X1 U9038 ( .A1(n10669), .A2(n9890), .ZN(n10693) );
  NAND2_X1 U9039 ( .A1(n6991), .A2(n6990), .ZN(n10766) );
  NAND2_X1 U9040 ( .A1(n7234), .A2(n11016), .ZN(n11164) );
  NAND2_X1 U9041 ( .A1(n7246), .A2(n10889), .ZN(n14781) );
  NAND2_X1 U9042 ( .A1(n8558), .A2(n8557), .ZN(n13323) );
  INV_X1 U9043 ( .A(n13323), .ZN(n7200) );
  NAND2_X1 U9044 ( .A1(n8476), .A2(n8475), .ZN(n12955) );
  INV_X1 U9045 ( .A(n12955), .ZN(n7206) );
  OR2_X1 U9046 ( .A1(n13718), .A2(n13717), .ZN(n6672) );
  INV_X1 U9047 ( .A(n7832), .ZN(n7099) );
  NOR2_X1 U9048 ( .A1(n11076), .A2(n11075), .ZN(n6673) );
  NAND2_X1 U9049 ( .A1(n13489), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n6674) );
  INV_X1 U9050 ( .A(n8133), .ZN(n7338) );
  NAND2_X1 U9051 ( .A1(n9313), .A2(n9566), .ZN(n6675) );
  INV_X1 U9052 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10682) );
  INV_X1 U9053 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10537) );
  AND2_X1 U9054 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n10686), .ZN(n6676) );
  INV_X1 U9055 ( .A(n6956), .ZN(n11592) );
  NOR2_X1 U9056 ( .A1(n11304), .A2(n14658), .ZN(n6956) );
  OR2_X1 U9057 ( .A1(n11526), .A2(n11439), .ZN(n11701) );
  AND2_X1 U9058 ( .A1(n10341), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6677) );
  AND2_X1 U9059 ( .A1(n7337), .A2(n8880), .ZN(n6678) );
  AND2_X1 U9060 ( .A1(n12285), .A2(n14585), .ZN(n6679) );
  AND2_X1 U9061 ( .A1(n11008), .A2(n8364), .ZN(n6680) );
  INV_X1 U9062 ( .A(n7422), .ZN(n7349) );
  INV_X1 U9063 ( .A(n12351), .ZN(n6694) );
  INV_X1 U9064 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7091) );
  INV_X1 U9065 ( .A(n10921), .ZN(n6957) );
  INV_X1 U9066 ( .A(n14917), .ZN(n6953) );
  OR2_X1 U9067 ( .A1(n9866), .A2(n9856), .ZN(n6681) );
  INV_X1 U9068 ( .A(n15347), .ZN(n15323) );
  NAND2_X1 U9069 ( .A1(n8431), .A2(n8430), .ZN(n14650) );
  INV_X1 U9070 ( .A(n14650), .ZN(n7209) );
  NAND2_X1 U9071 ( .A1(n8336), .A2(n8335), .ZN(n15116) );
  INV_X1 U9072 ( .A(n15116), .ZN(n7198) );
  AOI211_X1 U9073 ( .C1(n10821), .C2(n11901), .A(n10824), .B(n10823), .ZN(
        n10955) );
  AND2_X1 U9074 ( .A1(n8021), .A2(n12020), .ZN(n15347) );
  OR2_X1 U9075 ( .A1(n9779), .A2(n7309), .ZN(n6682) );
  AND2_X1 U9076 ( .A1(n7114), .A2(n11741), .ZN(n6683) );
  NAND2_X1 U9077 ( .A1(n6688), .A2(n7399), .ZN(n13372) );
  INV_X1 U9078 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7180) );
  INV_X1 U9079 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7183) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6713) );
  INV_X1 U9081 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n7178) );
  INV_X1 U9082 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7185) );
  INV_X2 U9083 ( .A(n6681), .ZN(P1_U4016) );
  NAND2_X1 U9084 ( .A1(n10030), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9856) );
  OR3_X1 U9085 ( .A1(n9905), .A2(n9903), .A3(n11743), .ZN(n9866) );
  NAND2_X1 U9086 ( .A1(n6685), .A2(n11332), .ZN(n11334) );
  NAND2_X1 U9087 ( .A1(n7123), .A2(n6686), .ZN(n6685) );
  OR2_X1 U9088 ( .A1(n8361), .A2(n7126), .ZN(n6686) );
  NOR2_X2 U9089 ( .A1(n8167), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n8164) );
  NAND3_X1 U9090 ( .A1(n6913), .A2(n6914), .A3(n8062), .ZN(n8065) );
  NAND2_X1 U9091 ( .A1(n8109), .A2(n8110), .ZN(n7333) );
  NAND2_X1 U9092 ( .A1(n6829), .A2(n6827), .ZN(n8108) );
  NAND2_X1 U9093 ( .A1(n8653), .A2(n8128), .ZN(n8672) );
  NAND3_X2 U9094 ( .A1(n9036), .A2(n9037), .A3(n6689), .ZN(n14810) );
  NAND2_X1 U9095 ( .A1(n11302), .A2(n11303), .ZN(n7255) );
  OAI21_X2 U9096 ( .B1(n6542), .B2(n7259), .A(n7256), .ZN(n14219) );
  NAND2_X1 U9097 ( .A1(n10888), .A2(n10887), .ZN(n10912) );
  OR2_X1 U9098 ( .A1(n14329), .A2(n14420), .ZN(n6835) );
  NAND2_X1 U9099 ( .A1(n14120), .A2(n14081), .ZN(n14082) );
  NOR2_X1 U9100 ( .A1(n12318), .A2(n6690), .ZN(n12335) );
  XNOR2_X1 U9101 ( .A(n12380), .B(n6691), .ZN(n12394) );
  XNOR2_X2 U9102 ( .A(n6692), .B(n12382), .ZN(n12353) );
  XNOR2_X1 U9103 ( .A(n11068), .B(n11131), .ZN(n15242) );
  NOR2_X1 U9104 ( .A1(n15205), .A2(n11067), .ZN(n15225) );
  NAND2_X1 U9105 ( .A1(n7016), .A2(n7015), .ZN(n12287) );
  AOI21_X1 U9106 ( .B1(n6698), .B2(n12413), .A(n12203), .ZN(n12204) );
  NAND2_X1 U9107 ( .A1(n12200), .A2(n12199), .ZN(n6698) );
  NAND2_X1 U9108 ( .A1(n6699), .A2(n12104), .ZN(n12109) );
  NAND2_X1 U9109 ( .A1(n12098), .A2(n6700), .ZN(n6699) );
  AOI21_X1 U9110 ( .B1(n6701), .B2(n12148), .A(n12603), .ZN(n12151) );
  NAND2_X1 U9111 ( .A1(n6709), .A2(n6708), .ZN(n12093) );
  NAND2_X1 U9112 ( .A1(n12090), .A2(n12219), .ZN(n6708) );
  INV_X1 U9113 ( .A(n6710), .ZN(n6709) );
  AOI21_X1 U9114 ( .B1(n12089), .B2(n12088), .A(n6711), .ZN(n6710) );
  NAND2_X1 U9115 ( .A1(n7311), .A2(n8059), .ZN(n8291) );
  OAI21_X1 U9116 ( .B1(n13268), .B2(n13351), .A(n6812), .ZN(n13355) );
  NAND2_X2 U9117 ( .A1(n8294), .A2(n8293), .ZN(n15106) );
  OR2_X1 U9118 ( .A1(n11771), .A2(n7945), .ZN(n7947) );
  OAI21_X1 U9119 ( .B1(n12428), .B2(n7977), .A(n6797), .ZN(n6796) );
  NAND2_X1 U9120 ( .A1(n7991), .A2(n6888), .ZN(n7491) );
  NAND2_X1 U9121 ( .A1(n6719), .A2(n9334), .ZN(n9347) );
  NAND2_X1 U9122 ( .A1(n6917), .A2(n7428), .ZN(n6719) );
  NAND4_X1 U9123 ( .A1(n14610), .A2(n7496), .A3(P2_ADDR_REG_19__SCAN_IN), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n7299) );
  AOI21_X1 U9124 ( .B1(n8170), .B2(n8171), .A(n8042), .ZN(n8201) );
  NAND2_X1 U9125 ( .A1(n9396), .A2(n9397), .ZN(n9395) );
  OAI21_X1 U9126 ( .B1(n6890), .B2(n6889), .A(n9591), .ZN(P1_U3242) );
  AOI21_X1 U9127 ( .B1(n6893), .B2(n9578), .A(n6892), .ZN(n6891) );
  NAND2_X1 U9128 ( .A1(n9399), .A2(n9398), .ZN(n6899) );
  OAI22_X1 U9129 ( .A1(n9383), .A2(n7297), .B1(n9384), .B2(n7298), .ZN(n9396)
         );
  AOI21_X1 U9130 ( .B1(n9524), .B2(n9523), .A(n9558), .ZN(n6893) );
  NAND2_X1 U9131 ( .A1(n9020), .A2(n9022), .ZN(n9011) );
  NAND2_X1 U9132 ( .A1(n6898), .A2(n7283), .ZN(n9432) );
  NAND2_X1 U9133 ( .A1(n9432), .A2(n9433), .ZN(n9431) );
  INV_X1 U9134 ( .A(n6891), .ZN(n6890) );
  NAND2_X1 U9135 ( .A1(n9464), .A2(n9463), .ZN(n9466) );
  OAI21_X1 U9136 ( .B1(n6906), .B2(n7281), .A(n6903), .ZN(n6908) );
  INV_X4 U9137 ( .A(n9078), .ZN(n9025) );
  NAND2_X1 U9138 ( .A1(n14767), .A2(n10981), .ZN(n10982) );
  AND3_X4 U9139 ( .A1(n9264), .A2(n8970), .A3(n8969), .ZN(n9313) );
  NAND2_X1 U9140 ( .A1(n6929), .A2(n10895), .ZN(n14785) );
  INV_X1 U9141 ( .A(n14764), .ZN(n6723) );
  NAND2_X1 U9142 ( .A1(n10913), .A2(n14782), .ZN(n6929) );
  NAND2_X1 U9143 ( .A1(n10669), .A2(n6736), .ZN(n6734) );
  NAND3_X1 U9144 ( .A1(n6729), .A2(n7342), .A3(n6728), .ZN(n11256) );
  NAND3_X1 U9145 ( .A1(n6730), .A2(n6732), .A3(n6733), .ZN(n6729) );
  INV_X1 U9146 ( .A(n10669), .ZN(n6730) );
  NAND3_X1 U9147 ( .A1(n6734), .A2(n6732), .A3(n6731), .ZN(n11178) );
  NAND2_X1 U9148 ( .A1(n13883), .A2(n6746), .ZN(n6744) );
  NAND2_X1 U9149 ( .A1(n6744), .A2(n6745), .ZN(n13855) );
  NAND2_X1 U9150 ( .A1(n9313), .A2(n6752), .ZN(n9581) );
  INV_X2 U9151 ( .A(n13728), .ZN(n9892) );
  NAND3_X1 U9152 ( .A1(n13798), .A2(n9951), .A3(n13922), .ZN(n9865) );
  INV_X4 U9153 ( .A(n9886), .ZN(n13798) );
  NAND2_X1 U9154 ( .A1(n7175), .A2(n14534), .ZN(n14535) );
  NAND2_X1 U9155 ( .A1(n6760), .A2(n14518), .ZN(n14522) );
  NOR2_X1 U9156 ( .A1(n15427), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n14524) );
  OAI21_X1 U9157 ( .B1(n6756), .B2(n6759), .A(n14521), .ZN(n6755) );
  INV_X1 U9158 ( .A(n6760), .ZN(n6756) );
  NAND2_X1 U9159 ( .A1(n6758), .A2(n6760), .ZN(n6757) );
  NOR2_X1 U9160 ( .A1(n14521), .A2(n6759), .ZN(n6758) );
  INV_X1 U9161 ( .A(n14518), .ZN(n6759) );
  NAND2_X1 U9162 ( .A1(n15425), .A2(n15426), .ZN(n6760) );
  NAND3_X1 U9163 ( .A1(n7188), .A2(n7186), .A3(n7187), .ZN(n6761) );
  NAND2_X1 U9164 ( .A1(n6767), .A2(n14704), .ZN(n14710) );
  NAND2_X1 U9165 ( .A1(n7979), .A2(n12205), .ZN(n8814) );
  INV_X1 U9166 ( .A(n12217), .ZN(n6783) );
  OAI21_X1 U9167 ( .B1(n7457), .B2(n7072), .A(n6787), .ZN(n7662) );
  NAND2_X1 U9168 ( .A1(n7457), .A2(n6787), .ZN(n6786) );
  NAND2_X1 U9169 ( .A1(n7523), .A2(n7522), .ZN(n7521) );
  NAND2_X1 U9170 ( .A1(n7810), .A2(n6791), .ZN(n6790) );
  NAND2_X1 U9171 ( .A1(n7712), .A2(n7467), .ZN(n7469) );
  INV_X1 U9172 ( .A(n6795), .ZN(n6794) );
  AND2_X2 U9173 ( .A1(n6796), .A2(n7062), .ZN(n12414) );
  NAND2_X1 U9174 ( .A1(n6798), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10619) );
  NAND2_X1 U9175 ( .A1(n6799), .A2(n10617), .ZN(n10618) );
  MUX2_X1 U9176 ( .A(n12781), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  MUX2_X1 U9177 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12781), .S(n10577), .Z(n10511)
         );
  MUX2_X1 U9178 ( .A(n10789), .B(n15181), .S(P3_IR_REG_0__SCAN_IN), .Z(n10790)
         );
  NAND2_X1 U9179 ( .A1(n10407), .A2(n8848), .ZN(n10636) );
  NAND2_X1 U9180 ( .A1(n10409), .A2(n10408), .ZN(n10407) );
  NAND2_X1 U9181 ( .A1(n10391), .A2(n8847), .ZN(n10409) );
  NAND2_X1 U9182 ( .A1(n10393), .A2(n10392), .ZN(n10391) );
  OAI21_X2 U9183 ( .B1(n6806), .B2(n6608), .A(n8860), .ZN(n11368) );
  INV_X1 U9184 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n6809) );
  NOR2_X2 U9185 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n8174) );
  INV_X1 U9186 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6811) );
  XNOR2_X2 U9187 ( .A(n6813), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8179) );
  INV_X1 U9188 ( .A(n8842), .ZN(n12988) );
  NAND2_X2 U9189 ( .A1(n14162), .A2(n14163), .ZN(n14164) );
  NAND2_X1 U9190 ( .A1(n6814), .A2(n8119), .ZN(n9368) );
  INV_X1 U9191 ( .A(n8266), .ZN(n8058) );
  NAND2_X1 U9192 ( .A1(n6817), .A2(n6815), .ZN(n7312) );
  NAND2_X1 U9193 ( .A1(n8266), .A2(n8059), .ZN(n6815) );
  NAND2_X1 U9194 ( .A1(n6816), .A2(SI_5_), .ZN(n8059) );
  MUX2_X1 U9195 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8043), .Z(n6816) );
  INV_X1 U9196 ( .A(n8290), .ZN(n6817) );
  MUX2_X1 U9197 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n9367), .Z(n8060) );
  OAI21_X1 U9198 ( .B1(n8384), .B2(n6824), .A(n6821), .ZN(n8425) );
  NAND2_X1 U9199 ( .A1(n8384), .A2(n6821), .ZN(n6820) );
  OAI21_X1 U9200 ( .B1(n8384), .B2(n8385), .A(n8080), .ZN(n8405) );
  NAND2_X1 U9201 ( .A1(n8385), .A2(n8080), .ZN(n6826) );
  NAND2_X1 U9202 ( .A1(n7314), .A2(n6831), .ZN(n6829) );
  NAND3_X1 U9203 ( .A1(n6837), .A2(n6836), .A3(n6835), .ZN(n14425) );
  INV_X1 U9204 ( .A(n11854), .ZN(n6866) );
  INV_X2 U9205 ( .A(n7424), .ZN(n11901) );
  AOI21_X2 U9206 ( .B1(n10814), .B2(n12063), .A(n10818), .ZN(n7424) );
  NAND2_X1 U9207 ( .A1(n11787), .A2(n6870), .ZN(n6868) );
  NAND2_X1 U9208 ( .A1(n6877), .A2(n6876), .ZN(n6874) );
  AND2_X1 U9209 ( .A1(n6879), .A2(n11576), .ZN(n6875) );
  NAND2_X1 U9210 ( .A1(n7693), .A2(n7487), .ZN(n7798) );
  NAND3_X1 U9211 ( .A1(n6895), .A2(n9482), .A3(n6894), .ZN(n7279) );
  NAND3_X1 U9212 ( .A1(n9484), .A2(n6897), .A3(n6896), .ZN(n9504) );
  NAND3_X1 U9213 ( .A1(n9467), .A2(n9482), .A3(n9468), .ZN(n6897) );
  NAND3_X1 U9214 ( .A1(n9467), .A2(n9468), .A3(n9483), .ZN(n9484) );
  NAND3_X1 U9215 ( .A1(n6900), .A2(n6899), .A3(n6652), .ZN(n6898) );
  INV_X1 U9216 ( .A(n7280), .ZN(n6901) );
  NAND2_X1 U9217 ( .A1(n6901), .A2(n9371), .ZN(n6906) );
  NAND2_X1 U9218 ( .A1(n6908), .A2(n6907), .ZN(n9383) );
  OAI21_X1 U9219 ( .B1(n9960), .B2(n7450), .A(n6910), .ZN(n8051) );
  NAND2_X1 U9220 ( .A1(n9960), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U9221 ( .A1(n8057), .A2(n6912), .ZN(n6914) );
  AND2_X1 U9222 ( .A1(n8056), .A2(n8061), .ZN(n6915) );
  NAND3_X1 U9223 ( .A1(n7269), .A2(n7418), .A3(n6653), .ZN(n6917) );
  NAND2_X1 U9224 ( .A1(n14785), .A2(n10896), .ZN(n10898) );
  INV_X1 U9225 ( .A(n14250), .ZN(n6930) );
  OAI21_X1 U9226 ( .B1(n6930), .B2(n6654), .A(n6933), .ZN(n14208) );
  INV_X1 U9227 ( .A(n6937), .ZN(n14135) );
  AND2_X1 U9228 ( .A1(n7231), .A2(n6943), .ZN(n6945) );
  NAND2_X1 U9229 ( .A1(n9008), .A2(n6944), .ZN(n6943) );
  NOR2_X2 U9230 ( .A1(n10941), .A2(n10942), .ZN(n10940) );
  NAND3_X1 U9231 ( .A1(n9537), .A2(n9535), .A3(n9015), .ZN(n9026) );
  NAND2_X1 U9232 ( .A1(n10846), .A2(n6965), .ZN(n6963) );
  INV_X1 U9233 ( .A(n6968), .ZN(n6969) );
  NAND2_X1 U9234 ( .A1(n13248), .A2(n6989), .ZN(n6991) );
  NAND2_X1 U9235 ( .A1(n6992), .A2(n6993), .ZN(n6994) );
  INV_X2 U9236 ( .A(n8172), .ZN(n8389) );
  OAI211_X2 U9237 ( .C1(n8693), .C2(n9990), .A(n6996), .B(n6619), .ZN(n10299)
         );
  OR2_X1 U9238 ( .A1(n8227), .A2(n9982), .ZN(n6996) );
  NAND2_X1 U9239 ( .A1(n6997), .A2(n6998), .ZN(n13205) );
  NAND2_X1 U9240 ( .A1(n13239), .A2(n7001), .ZN(n6997) );
  OAI21_X1 U9241 ( .B1(n13188), .B2(n7005), .A(n7003), .ZN(n13162) );
  AOI21_X2 U9242 ( .B1(n12365), .B2(n12364), .A(n12363), .ZN(n12373) );
  AOI21_X1 U9243 ( .B1(n12286), .B2(n14585), .A(n6679), .ZN(n7016) );
  NAND2_X1 U9244 ( .A1(n12698), .A2(n10956), .ZN(n12079) );
  OAI21_X1 U9245 ( .B1(n7558), .B2(n7531), .A(n7533), .ZN(n7023) );
  INV_X1 U9246 ( .A(n7023), .ZN(n7022) );
  NAND2_X1 U9247 ( .A1(n11463), .A2(n7029), .ZN(n7028) );
  NAND2_X1 U9248 ( .A1(n7028), .A2(n7030), .ZN(n11484) );
  NAND2_X1 U9249 ( .A1(n7053), .A2(n7054), .ZN(n12041) );
  NAND2_X1 U9250 ( .A1(n12412), .A2(n7057), .ZN(n7053) );
  NAND2_X1 U9251 ( .A1(n12412), .A2(n7061), .ZN(n7056) );
  AOI21_X1 U9252 ( .B1(n12412), .B2(n12413), .A(n12207), .ZN(n8813) );
  AND2_X1 U9253 ( .A1(n7992), .A2(n7066), .ZN(n7499) );
  NAND2_X1 U9254 ( .A1(n7992), .A2(n7067), .ZN(n7501) );
  NOR2_X2 U9256 ( .A1(n11230), .A2(n11494), .ZN(n11232) );
  INV_X2 U9257 ( .A(n10320), .ZN(n10458) );
  OAI21_X1 U9258 ( .B1(n7833), .B2(n7093), .A(n7092), .ZN(n7098) );
  INV_X1 U9259 ( .A(n7098), .ZN(n7855) );
  NAND2_X1 U9260 ( .A1(n7460), .A2(n6647), .ZN(n7100) );
  NAND2_X1 U9261 ( .A1(n7460), .A2(n7459), .ZN(n7681) );
  NAND2_X1 U9262 ( .A1(n7111), .A2(n7109), .ZN(n7879) );
  NAND2_X1 U9263 ( .A1(n7110), .A2(n7114), .ZN(n7109) );
  NAND2_X1 U9264 ( .A1(n7857), .A2(n7112), .ZN(n7110) );
  NAND2_X1 U9265 ( .A1(n7856), .A2(n6683), .ZN(n7111) );
  NAND2_X1 U9266 ( .A1(n7856), .A2(n11741), .ZN(n7113) );
  NAND2_X2 U9267 ( .A1(n12948), .A2(n6598), .ZN(n12878) );
  NAND2_X2 U9268 ( .A1(n12947), .A2(n8483), .ZN(n12948) );
  OAI21_X1 U9269 ( .B1(n8807), .B2(n13274), .A(n7115), .ZN(P2_U3192) );
  AOI21_X1 U9270 ( .B1(n8782), .B2(n7119), .A(n7116), .ZN(n7115) );
  NAND2_X1 U9271 ( .A1(n12902), .A2(n6636), .ZN(n12837) );
  NAND2_X2 U9272 ( .A1(n8588), .A2(n12895), .ZN(n12902) );
  AND2_X1 U9273 ( .A1(n8263), .A2(n8246), .ZN(n7120) );
  NAND2_X1 U9274 ( .A1(n12881), .A2(n7122), .ZN(n12824) );
  NAND2_X2 U9275 ( .A1(n8524), .A2(n12873), .ZN(n12881) );
  INV_X1 U9276 ( .A(n7124), .ZN(n7123) );
  OAI21_X1 U9277 ( .B1(n8360), .B2(n7126), .A(n8383), .ZN(n7124) );
  NAND2_X1 U9278 ( .A1(n11008), .A2(n7125), .ZN(n11048) );
  NAND2_X1 U9279 ( .A1(n8361), .A2(n8360), .ZN(n11008) );
  NAND2_X1 U9280 ( .A1(n11362), .A2(n7127), .ZN(n12794) );
  NAND2_X1 U9281 ( .A1(n12939), .A2(n7128), .ZN(n12785) );
  NAND2_X2 U9282 ( .A1(n12849), .A2(n8708), .ZN(n12939) );
  NAND2_X1 U9283 ( .A1(n10465), .A2(n6635), .ZN(n8310) );
  NAND2_X1 U9284 ( .A1(n7131), .A2(n6554), .ZN(n8897) );
  NAND2_X1 U9285 ( .A1(n7131), .A2(n9850), .ZN(n15146) );
  NOR2_X1 U9286 ( .A1(n7382), .A2(n7131), .ZN(n10168) );
  NAND2_X1 U9287 ( .A1(n11191), .A2(n8858), .ZN(n7132) );
  NAND2_X1 U9288 ( .A1(n15033), .A2(n15032), .ZN(n15031) );
  NAND2_X1 U9289 ( .A1(n10834), .A2(n10836), .ZN(n7133) );
  XNOR2_X1 U9290 ( .A(n7134), .B(n10433), .ZN(n10392) );
  INV_X4 U9291 ( .A(n8227), .ZN(n8694) );
  NAND2_X2 U9292 ( .A1(n7136), .A2(n9960), .ZN(n8227) );
  NAND2_X2 U9293 ( .A1(n7140), .A2(n7137), .ZN(n8188) );
  INV_X1 U9294 ( .A(n8863), .ZN(n7150) );
  NAND2_X1 U9295 ( .A1(n13199), .A2(n7154), .ZN(n7151) );
  NAND2_X1 U9296 ( .A1(n7151), .A2(n7152), .ZN(n8869) );
  NAND2_X1 U9297 ( .A1(n7165), .A2(n7164), .ZN(n13132) );
  NAND2_X1 U9298 ( .A1(n13256), .A2(n8852), .ZN(n7168) );
  NAND2_X1 U9299 ( .A1(n7168), .A2(n7169), .ZN(n10653) );
  INV_X1 U9300 ( .A(n13256), .ZN(n7172) );
  INV_X1 U9301 ( .A(n14714), .ZN(n7187) );
  NOR2_X2 U9302 ( .A1(n10855), .A2(n15136), .ZN(n15022) );
  INV_X1 U9303 ( .A(n15126), .ZN(n7196) );
  INV_X1 U9304 ( .A(n10853), .ZN(n7197) );
  INV_X1 U9305 ( .A(n10773), .ZN(n7199) );
  NOR2_X2 U9306 ( .A1(n13230), .A2(n13328), .ZN(n7201) );
  AND2_X2 U9307 ( .A1(n13112), .A2(n6572), .ZN(n13058) );
  NAND2_X2 U9308 ( .A1(n8996), .A2(n7211), .ZN(n14454) );
  AOI21_X2 U9309 ( .B1(n7213), .B2(n6601), .A(n7212), .ZN(n7211) );
  NAND2_X1 U9310 ( .A1(n14092), .A2(n7216), .ZN(n7215) );
  OAI211_X1 U9311 ( .C1(n14804), .C2(n7219), .A(n10891), .B(n7220), .ZN(n10947) );
  NAND2_X1 U9312 ( .A1(n10947), .A2(n10948), .ZN(n10914) );
  NAND2_X1 U9313 ( .A1(n10872), .A2(n7221), .ZN(n7220) );
  INV_X1 U9314 ( .A(n10872), .ZN(n7219) );
  INV_X1 U9315 ( .A(n10871), .ZN(n7221) );
  NAND2_X1 U9316 ( .A1(n10873), .A2(n10872), .ZN(n10892) );
  OAI21_X2 U9317 ( .B1(n14176), .B2(n7223), .A(n6624), .ZN(n14124) );
  AND2_X2 U9318 ( .A1(n9008), .A2(n9960), .ZN(n9469) );
  INV_X2 U9319 ( .A(n9027), .ZN(n10862) );
  NAND2_X1 U9320 ( .A1(n11015), .A2(n7235), .ZN(n7232) );
  NAND2_X1 U9321 ( .A1(n7232), .A2(n7233), .ZN(n11224) );
  NAND2_X1 U9322 ( .A1(n7238), .A2(n7239), .ZN(n14162) );
  NAND2_X1 U9323 ( .A1(n7245), .A2(n7244), .ZN(n10970) );
  AOI21_X1 U9324 ( .B1(n14783), .B2(n7247), .A(n6633), .ZN(n7244) );
  NAND3_X1 U9325 ( .A1(n10912), .A2(n10916), .A3(n14783), .ZN(n7245) );
  INV_X1 U9326 ( .A(n7250), .ZN(n14150) );
  NOR2_X1 U9327 ( .A1(n14167), .A2(n14102), .ZN(n7252) );
  NAND2_X2 U9328 ( .A1(n7255), .A2(n7253), .ZN(n14676) );
  OAI21_X2 U9329 ( .B1(n14280), .B2(n14068), .A(n14067), .ZN(n14267) );
  OAI21_X2 U9330 ( .B1(n14301), .B2(n14064), .A(n14065), .ZN(n14280) );
  NAND2_X2 U9331 ( .A1(n14062), .A2(n14061), .ZN(n14301) );
  NAND2_X1 U9332 ( .A1(n7261), .A2(n9313), .ZN(n8979) );
  NAND2_X1 U9333 ( .A1(n9033), .A2(n7266), .ZN(n9065) );
  NAND2_X1 U9334 ( .A1(n9287), .A2(n7270), .ZN(n7269) );
  NAND2_X1 U9335 ( .A1(n7277), .A2(n9502), .ZN(n9524) );
  NAND3_X1 U9336 ( .A1(n7279), .A2(n9484), .A3(n7278), .ZN(n7277) );
  INV_X1 U9337 ( .A(n9358), .ZN(n7282) );
  NAND2_X1 U9338 ( .A1(n7285), .A2(n7286), .ZN(n9228) );
  NAND3_X1 U9339 ( .A1(n9194), .A2(n6649), .A3(n9193), .ZN(n7285) );
  NAND2_X1 U9340 ( .A1(n7288), .A2(n7289), .ZN(n9189) );
  NAND3_X1 U9341 ( .A1(n9159), .A2(n6650), .A3(n9158), .ZN(n7288) );
  NAND4_X1 U9342 ( .A1(n8970), .A2(n9264), .A3(n9009), .A4(n8969), .ZN(n9302)
         );
  NOR2_X2 U9343 ( .A1(n9302), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n9020) );
  NAND2_X1 U9344 ( .A1(n7291), .A2(n7293), .ZN(n9154) );
  NAND3_X1 U9345 ( .A1(n9124), .A2(n7292), .A3(n9123), .ZN(n7291) );
  NAND4_X1 U9346 ( .A1(n14043), .A2(n7494), .A3(n7495), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n7300) );
  OAI21_X1 U9347 ( .B1(n8043), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n7301), .ZN(
        n8041) );
  NAND2_X1 U9348 ( .A1(n7302), .A2(n9855), .ZN(P2_U3328) );
  NAND2_X1 U9349 ( .A1(n7303), .A2(n11381), .ZN(n7302) );
  NAND2_X1 U9350 ( .A1(n7305), .A2(n7304), .ZN(n7303) );
  OAI22_X1 U9351 ( .A1(n9849), .A2(n9836), .B1(n9843), .B2(n7306), .ZN(n7305)
         );
  OR2_X1 U9352 ( .A1(n9841), .A2(n9842), .ZN(n7306) );
  NAND2_X1 U9353 ( .A1(n8089), .A2(n8088), .ZN(n8445) );
  NAND2_X1 U9354 ( .A1(n8331), .A2(n7329), .ZN(n7326) );
  NAND2_X1 U9355 ( .A1(n7326), .A2(n7327), .ZN(n8365) );
  NAND3_X1 U9356 ( .A1(n8126), .A2(n8128), .A3(n8127), .ZN(n8653) );
  NAND2_X1 U9357 ( .A1(n8111), .A2(n7333), .ZN(n8594) );
  OAI21_X1 U9358 ( .B1(n8690), .B2(n7334), .A(n6678), .ZN(n8884) );
  OAI22_X1 U9359 ( .A1(n10424), .A2(n10423), .B1(n9871), .B2(n7341), .ZN(
        n10459) );
  NAND2_X1 U9360 ( .A1(n13897), .A2(n6667), .ZN(n7355) );
  NAND2_X1 U9361 ( .A1(n7362), .A2(n6632), .ZN(n7357) );
  INV_X1 U9362 ( .A(n13773), .ZN(n7374) );
  OAI211_X1 U9363 ( .C1(n13889), .C2(n7369), .A(n7365), .B(n7363), .ZN(n13807)
         );
  NAND2_X1 U9364 ( .A1(n13889), .A2(n7364), .ZN(n7363) );
  AND2_X1 U9365 ( .A1(n6584), .A2(n7372), .ZN(n7364) );
  OAI21_X1 U9366 ( .B1(n7371), .B2(n6584), .A(n7366), .ZN(n7365) );
  NAND2_X1 U9367 ( .A1(n7371), .A2(n7367), .ZN(n7366) );
  INV_X1 U9368 ( .A(n7372), .ZN(n7368) );
  NAND2_X1 U9369 ( .A1(n7371), .A2(n7370), .ZN(n7369) );
  INV_X1 U9370 ( .A(n6584), .ZN(n7370) );
  NAND2_X1 U9371 ( .A1(n13853), .A2(n6668), .ZN(n13808) );
  XNOR2_X2 U9372 ( .A(n9583), .B(n9582), .ZN(n9905) );
  INV_X1 U9373 ( .A(n9313), .ZN(n9567) );
  NAND2_X1 U9374 ( .A1(n7382), .A2(n9596), .ZN(n9599) );
  NAND2_X1 U9375 ( .A1(n10302), .A2(n7382), .ZN(n15092) );
  NAND2_X1 U9376 ( .A1(n9609), .A2(n9608), .ZN(n7385) );
  NAND3_X1 U9377 ( .A1(n9681), .A2(n9680), .A3(n7387), .ZN(n7386) );
  NAND2_X1 U9378 ( .A1(n7386), .A2(n7388), .ZN(n9709) );
  INV_X1 U9379 ( .A(n9684), .ZN(n7390) );
  NAND3_X1 U9380 ( .A1(n9714), .A2(n9713), .A3(n6644), .ZN(n7391) );
  NAND2_X1 U9381 ( .A1(n7391), .A2(n7392), .ZN(n9720) );
  NAND3_X1 U9382 ( .A1(n9747), .A2(n9746), .A3(n6641), .ZN(n7393) );
  NAND2_X1 U9383 ( .A1(n7393), .A2(n7394), .ZN(n9753) );
  NAND3_X1 U9384 ( .A1(n9649), .A2(n9648), .A3(n6638), .ZN(n7395) );
  NAND2_X1 U9385 ( .A1(n7395), .A2(n7396), .ZN(n9655) );
  NAND3_X1 U9386 ( .A1(n9638), .A2(n9637), .A3(n6645), .ZN(n7397) );
  NAND2_X1 U9387 ( .A1(n7397), .A2(n7398), .ZN(n9644) );
  NAND3_X1 U9388 ( .A1(n9670), .A2(n9669), .A3(n6646), .ZN(n7402) );
  NAND2_X1 U9389 ( .A1(n7402), .A2(n6648), .ZN(n9676) );
  NAND2_X1 U9390 ( .A1(n7404), .A2(n7405), .ZN(n9633) );
  NAND3_X1 U9391 ( .A1(n9628), .A2(n9627), .A3(n6642), .ZN(n7404) );
  NAND3_X1 U9392 ( .A1(n9736), .A2(n9735), .A3(n6643), .ZN(n7407) );
  NAND2_X1 U9393 ( .A1(n7407), .A2(n7408), .ZN(n9742) );
  NAND3_X1 U9394 ( .A1(n9660), .A2(n9659), .A3(n6637), .ZN(n7410) );
  NAND2_X1 U9395 ( .A1(n7410), .A2(n7411), .ZN(n9665) );
  NAND3_X1 U9396 ( .A1(n9725), .A2(n9724), .A3(n6639), .ZN(n7413) );
  NAND2_X1 U9397 ( .A1(n7413), .A2(n7414), .ZN(n9731) );
  NAND2_X1 U9398 ( .A1(n8123), .A2(n8122), .ZN(n8619) );
  XNOR2_X1 U9399 ( .A(n8748), .B(n8747), .ZN(n8782) );
  OR2_X2 U9400 ( .A1(n13297), .A2(n13145), .ZN(n13133) );
  NAND2_X1 U9401 ( .A1(n13117), .A2(n13118), .ZN(n13116) );
  NAND2_X1 U9402 ( .A1(n11403), .A2(n12092), .ZN(n11402) );
  OR2_X1 U9403 ( .A1(n7922), .A2(n15342), .ZN(n7923) );
  INV_X1 U9404 ( .A(n13272), .ZN(n8960) );
  NAND2_X1 U9405 ( .A1(n10333), .A2(n10334), .ZN(n10332) );
  INV_X1 U9406 ( .A(n7506), .ZN(n12769) );
  NAND2_X1 U9407 ( .A1(n11586), .A2(n11585), .ZN(n11619) );
  NAND2_X1 U9408 ( .A1(n9536), .A2(n9538), .ZN(n10868) );
  AND2_X1 U9409 ( .A1(n14164), .A2(n14165), .ZN(n14351) );
  NAND2_X1 U9410 ( .A1(n10305), .A2(n8902), .ZN(n10333) );
  NAND2_X1 U9411 ( .A1(n9064), .A2(n9063), .ZN(n9081) );
  XNOR2_X1 U9412 ( .A(n14082), .B(n14104), .ZN(n14329) );
  NAND2_X1 U9413 ( .A1(n8998), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n8988) );
  OR2_X1 U9414 ( .A1(n9017), .A2(n14441), .ZN(n9010) );
  MUX2_X1 U9415 ( .A(n14347), .B(n14101), .S(n9025), .Z(n9430) );
  INV_X1 U9416 ( .A(n9720), .ZN(n9723) );
  NAND2_X1 U9417 ( .A1(n8125), .A2(SI_24_), .ZN(n8128) );
  AND2_X1 U9418 ( .A1(n9797), .A2(n9786), .ZN(n9787) );
  INV_X1 U9419 ( .A(n13052), .ZN(n13267) );
  NAND2_X1 U9420 ( .A1(n9486), .A2(n9485), .ZN(n9518) );
  NAND2_X1 U9421 ( .A1(n9866), .A2(n10009), .ZN(n10036) );
  OR2_X1 U9422 ( .A1(n9528), .A2(n10687), .ZN(n9024) );
  OR2_X1 U9423 ( .A1(n6720), .A2(n14824), .ZN(n14401) );
  NAND2_X1 U9424 ( .A1(n9864), .A2(n6720), .ZN(n10032) );
  NAND2_X1 U9425 ( .A1(n8181), .A2(n11823), .ZN(n8234) );
  INV_X1 U9426 ( .A(n8181), .ZN(n13379) );
  XNOR2_X1 U9427 ( .A(n8715), .B(n8714), .ZN(n13384) );
  NAND2_X1 U9428 ( .A1(n10870), .A2(n10869), .ZN(n14804) );
  NAND2_X1 U9429 ( .A1(n8998), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n9003) );
  INV_X1 U9430 ( .A(n15048), .ZN(n13242) );
  AND2_X1 U9431 ( .A1(n8893), .A2(n15050), .ZN(n15038) );
  INV_X1 U9432 ( .A(n15038), .ZN(n15048) );
  AND2_X1 U9433 ( .A1(n14392), .A2(n14093), .ZN(n7416) );
  AND2_X1 U9434 ( .A1(n9330), .A2(n14268), .ZN(n7417) );
  AND2_X1 U9435 ( .A1(n14281), .A2(n9317), .ZN(n7418) );
  INV_X1 U9436 ( .A(n8822), .ZN(n12399) );
  OR2_X1 U9437 ( .A1(n15424), .A2(n13480), .ZN(n7420) );
  INV_X1 U9438 ( .A(n15424), .ZN(n8836) );
  INV_X1 U9439 ( .A(n12694), .ZN(n8838) );
  OR2_X1 U9440 ( .A1(n15412), .A2(n15406), .ZN(n12762) );
  INV_X1 U9441 ( .A(n12762), .ZN(n8823) );
  AND2_X2 U9442 ( .A1(n8034), .A2(n8033), .ZN(n15412) );
  AND2_X1 U9443 ( .A1(n9878), .A2(n9877), .ZN(n7421) );
  AND2_X1 U9444 ( .A1(n11176), .A2(n11175), .ZN(n7422) );
  AND2_X1 U9445 ( .A1(n15304), .A2(n11782), .ZN(n7423) );
  AND2_X1 U9446 ( .A1(n8102), .A2(n8101), .ZN(n7425) );
  INV_X1 U9447 ( .A(n7951), .ZN(n12588) );
  AND2_X1 U9448 ( .A1(n8839), .A2(n7420), .ZN(n7426) );
  AND2_X1 U9449 ( .A1(n11036), .A2(n12706), .ZN(n7427) );
  AND2_X1 U9450 ( .A1(n9331), .A2(n7417), .ZN(n7428) );
  AND2_X1 U9451 ( .A1(n13103), .A2(n12853), .ZN(n7429) );
  OR2_X1 U9452 ( .A1(n12033), .A2(n11558), .ZN(n7430) );
  OR2_X1 U9453 ( .A1(n13683), .A2(n13682), .ZN(n7431) );
  AND2_X1 U9454 ( .A1(n8825), .A2(n8824), .ZN(n7432) );
  OR2_X1 U9455 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10787), .ZN(n7433) );
  AND2_X1 U9456 ( .A1(n8148), .A2(n8147), .ZN(n7434) );
  AND3_X1 U9457 ( .A1(n8148), .A2(n8146), .A3(n8147), .ZN(n7435) );
  AND2_X1 U9458 ( .A1(n8084), .A2(n8083), .ZN(n7436) );
  INV_X1 U9459 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10369) );
  INV_X1 U9460 ( .A(n13393), .ZN(n13380) );
  INV_X1 U9461 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8049) );
  INV_X1 U9462 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7472) );
  INV_X1 U9463 ( .A(n14262), .ZN(n14071) );
  AND2_X1 U9464 ( .A1(n8088), .A2(n8087), .ZN(n7437) );
  INV_X1 U9465 ( .A(n15160), .ZN(n15164) );
  NAND2_X1 U9466 ( .A1(n8744), .A2(n8743), .ZN(n12961) );
  NOR2_X1 U9467 ( .A1(n7775), .A2(n12563), .ZN(n7438) );
  INV_X1 U9468 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n13526) );
  INV_X1 U9469 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n13629) );
  INV_X1 U9470 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10422) );
  INV_X1 U9471 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n13373) );
  AND2_X2 U9472 ( .A1(n7947), .A2(n7946), .ZN(n7439) );
  INV_X1 U9473 ( .A(n12884), .ZN(n12932) );
  NAND2_X1 U9474 ( .A1(n10055), .A2(n10067), .ZN(n12884) );
  INV_X1 U9476 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8002) );
  OR2_X1 U9477 ( .A1(n13268), .A2(n13246), .ZN(n7440) );
  AND4_X1 U9478 ( .A1(n14123), .A2(n9554), .A3(n14177), .A4(n14156), .ZN(n7441) );
  INV_X1 U9479 ( .A(n15319), .ZN(n15338) );
  AND2_X1 U9480 ( .A1(n7987), .A2(n12227), .ZN(n15319) );
  OR2_X1 U9481 ( .A1(n10577), .A2(n6546), .ZN(n7442) );
  INV_X1 U9482 ( .A(n10704), .ZN(n8337) );
  NOR2_X1 U9483 ( .A1(n7943), .A2(n11761), .ZN(n7443) );
  AND2_X1 U9484 ( .A1(n11987), .A2(n11988), .ZN(n7444) );
  AND2_X1 U9485 ( .A1(n12598), .A2(n12147), .ZN(n12615) );
  NAND2_X1 U9486 ( .A1(n12466), .A2(n12465), .ZN(n7445) );
  AND2_X1 U9487 ( .A1(n7849), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7446) );
  INV_X1 U9488 ( .A(n12468), .ZN(n12470) );
  AND2_X1 U9489 ( .A1(n9593), .A2(n9592), .ZN(n9594) );
  MUX2_X1 U9490 ( .A(n12986), .B(n10756), .S(n9784), .Z(n9611) );
  NAND2_X1 U9491 ( .A1(n10868), .A2(n9393), .ZN(n9029) );
  OAI21_X1 U9492 ( .B1(n9081), .B2(n9080), .A(n9079), .ZN(n9083) );
  AND2_X1 U9493 ( .A1(n11583), .A2(n9260), .ZN(n9261) );
  AND2_X1 U9494 ( .A1(n9283), .A2(n9282), .ZN(n9284) );
  INV_X1 U9495 ( .A(n9682), .ZN(n9683) );
  INV_X1 U9496 ( .A(n9721), .ZN(n9722) );
  MUX2_X1 U9497 ( .A(n14198), .B(n14079), .S(n9500), .Z(n9397) );
  MUX2_X1 U9498 ( .A(n14347), .B(n14101), .S(n9500), .Z(n9433) );
  INV_X1 U9499 ( .A(n9743), .ZN(n9744) );
  AND2_X1 U9500 ( .A1(n13118), .A2(n9826), .ZN(n9827) );
  AND2_X1 U9501 ( .A1(n13105), .A2(n9827), .ZN(n9828) );
  AND2_X1 U9502 ( .A1(n13090), .A2(n9828), .ZN(n9829) );
  AND2_X1 U9503 ( .A1(n13063), .A2(n9829), .ZN(n9830) );
  INV_X1 U9504 ( .A(n9558), .ZN(n9559) );
  INV_X1 U9505 ( .A(n11441), .ZN(n11437) );
  INV_X1 U9506 ( .A(n12552), .ZN(n7957) );
  INV_X1 U9507 ( .A(n9881), .ZN(n9882) );
  INV_X1 U9508 ( .A(n14334), .ZN(n14335) );
  NAND2_X1 U9509 ( .A1(n6544), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9056) );
  INV_X1 U9510 ( .A(n8713), .ZN(n8132) );
  INV_X1 U9511 ( .A(SI_15_), .ZN(n8090) );
  INV_X1 U9512 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8963) );
  INV_X1 U9513 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n7699) );
  INV_X1 U9514 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n11939) );
  NAND2_X1 U9515 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  INV_X1 U9516 ( .A(n12414), .ZN(n12415) );
  NOR2_X1 U9517 ( .A1(n7849), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U9518 ( .A1(n7958), .A2(n7957), .ZN(n12549) );
  INV_X1 U9519 ( .A(n12615), .ZN(n7948) );
  NAND2_X1 U9520 ( .A1(n15305), .A2(n7940), .ZN(n11725) );
  INV_X1 U9521 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7483) );
  INV_X1 U9522 ( .A(n9593), .ZN(n9845) );
  INV_X1 U9523 ( .A(n8600), .ZN(n8599) );
  INV_X1 U9524 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10550) );
  INV_X1 U9525 ( .A(n8561), .ZN(n8559) );
  INV_X1 U9526 ( .A(n10303), .ZN(n9812) );
  OAI22_X1 U9527 ( .A1(n9028), .A2(n13729), .B1(n9886), .B2(n10862), .ZN(n9863) );
  NAND2_X1 U9528 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  OAI22_X1 U9529 ( .A1(n9043), .A2(n9886), .B1(n10874), .B2(n13729), .ZN(n9874) );
  INV_X1 U9530 ( .A(n9565), .ZN(n9530) );
  INV_X1 U9531 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9125) );
  INV_X1 U9532 ( .A(n9859), .ZN(n9028) );
  AND2_X1 U9533 ( .A1(n11805), .A2(n11806), .ZN(n11803) );
  INV_X1 U9534 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n7763) );
  OR2_X1 U9535 ( .A1(n7871), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7885) );
  INV_X1 U9536 ( .A(n15261), .ZN(n11069) );
  NOR2_X1 U9537 ( .A1(n11702), .A2(n11703), .ZN(n11700) );
  AND2_X1 U9538 ( .A1(n12293), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12285) );
  NOR2_X1 U9539 ( .A1(n7885), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7899) );
  INV_X1 U9540 ( .A(n12481), .ZN(n12463) );
  AND2_X1 U9541 ( .A1(n12173), .A2(n12172), .ZN(n12540) );
  OR2_X1 U9542 ( .A1(n12614), .A2(n12565), .ZN(n12584) );
  OR2_X1 U9543 ( .A1(n11770), .A2(n7774), .ZN(n12563) );
  INV_X1 U9544 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7635) );
  INV_X1 U9545 ( .A(n10817), .ZN(n12074) );
  INV_X1 U9546 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7993) );
  OR2_X1 U9547 ( .A1(n7743), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7746) );
  INV_X1 U9548 ( .A(n10362), .ZN(n8263) );
  INV_X1 U9549 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8538) );
  NAND2_X2 U9550 ( .A1(n8888), .A2(n9845), .ZN(n8211) );
  NAND2_X1 U9551 ( .A1(n8697), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U9552 ( .A1(n8599), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n8631) );
  NAND2_X1 U9553 ( .A1(n8514), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8539) );
  OR2_X1 U9554 ( .A1(n8373), .A2(n14984), .ZN(n8395) );
  INV_X1 U9555 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n13652) );
  OR2_X1 U9556 ( .A1(n8633), .A2(n12818), .ZN(n8656) );
  NAND2_X1 U9557 ( .A1(n8452), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8479) );
  NAND2_X1 U9558 ( .A1(n13054), .A2(n12959), .ZN(n8957) );
  INV_X1 U9559 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8229) );
  OR2_X1 U9560 ( .A1(n13744), .A2(n13743), .ZN(n13745) );
  OR2_X1 U9561 ( .A1(n13751), .A2(n13750), .ZN(n13752) );
  INV_X1 U9562 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n13533) );
  INV_X1 U9563 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13812) );
  INV_X1 U9564 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14480) );
  OAI22_X1 U9565 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14491), .B1(n14492), 
        .B2(n14486), .ZN(n14548) );
  OR2_X1 U9566 ( .A1(n11827), .A2(n12607), .ZN(n11828) );
  OR2_X1 U9567 ( .A1(n8827), .A2(n8024), .ZN(n10826) );
  AND3_X1 U9568 ( .A1(n7865), .A2(n7864), .A3(n7863), .ZN(n12468) );
  NAND2_X1 U9569 ( .A1(n15169), .A2(n11063), .ZN(n11064) );
  INV_X1 U9570 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n11749) );
  INV_X1 U9571 ( .A(n11701), .ZN(n11704) );
  OR2_X1 U9572 ( .A1(n11819), .A2(n12774), .ZN(n10580) );
  NAND2_X1 U9573 ( .A1(n7842), .A2(n12187), .ZN(n12492) );
  INV_X1 U9574 ( .A(n12580), .ZN(n12554) );
  AND2_X1 U9575 ( .A1(n12149), .A2(n12152), .ZN(n12600) );
  OR2_X1 U9576 ( .A1(n10965), .A2(n7916), .ZN(n8830) );
  INV_X1 U9577 ( .A(n10744), .ZN(n8832) );
  OR2_X1 U9578 ( .A1(n12033), .A2(n12775), .ZN(n7883) );
  NAND3_X1 U9579 ( .A1(n10580), .A2(n12227), .A3(n6550), .ZN(n15340) );
  INV_X1 U9580 ( .A(n11634), .ZN(n15405) );
  AND2_X1 U9581 ( .A1(n10692), .A2(n12375), .ZN(n15356) );
  INV_X1 U9582 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8029) );
  NAND2_X1 U9583 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n13629), .ZN(n7476) );
  NOR2_X1 U9584 ( .A1(n7746), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7759) );
  INV_X1 U9585 ( .A(n12782), .ZN(n8731) );
  INV_X1 U9586 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n12862) );
  INV_X1 U9587 ( .A(n12861), .ZN(n8502) );
  NOR2_X1 U9588 ( .A1(n11057), .A2(n10810), .ZN(n10055) );
  XNOR2_X1 U9589 ( .A(n8643), .B(n8641), .ZN(n12808) );
  OR2_X1 U9590 ( .A1(n8539), .A2(n8538), .ZN(n8561) );
  OR2_X1 U9591 ( .A1(n10166), .A2(n8803), .ZN(n8804) );
  AND2_X1 U9592 ( .A1(n8736), .A2(n8735), .ZN(n8898) );
  INV_X1 U9593 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n14984) );
  AND2_X1 U9594 ( .A1(n10084), .A2(n10068), .ZN(n10072) );
  OR2_X1 U9595 ( .A1(n13333), .A2(n12971), .ZN(n9811) );
  NAND2_X1 U9596 ( .A1(n10055), .A2(n8793), .ZN(n12886) );
  OR2_X1 U9597 ( .A1(n15038), .A2(n8897), .ZN(n13236) );
  NAND2_X1 U9598 ( .A1(n10327), .A2(n10326), .ZN(n10325) );
  OR2_X1 U9599 ( .A1(n13387), .A2(n11738), .ZN(n8765) );
  NAND2_X1 U9600 ( .A1(n8156), .A2(n7434), .ZN(n8790) );
  NAND2_X1 U9601 ( .A1(n11254), .A2(n11253), .ZN(n11255) );
  OR2_X1 U9602 ( .A1(n9289), .A2(n9288), .ZN(n9308) );
  NOR2_X1 U9603 ( .A1(n9160), .A2(n13578), .ZN(n9198) );
  OR2_X1 U9604 ( .A1(n9350), .A2(n13812), .ZN(n9360) );
  INV_X1 U9605 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n13578) );
  INV_X1 U9606 ( .A(n9580), .ZN(n10235) );
  INV_X1 U9607 ( .A(n9947), .ZN(n10425) );
  OR2_X1 U9608 ( .A1(n10032), .A2(n9580), .ZN(n14288) );
  NAND2_X1 U9609 ( .A1(n10867), .A2(n10866), .ZN(n10882) );
  NAND2_X1 U9610 ( .A1(n14812), .A2(n14039), .ZN(n10316) );
  INV_X1 U9611 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n8977) );
  INV_X1 U9612 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14502) );
  INV_X1 U9613 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n14472) );
  OR2_X1 U9614 ( .A1(n10574), .A2(n10573), .ZN(n10588) );
  AOI21_X1 U9615 ( .B1(n11913), .B2(n11912), .A(n11900), .ZN(n11903) );
  NAND2_X1 U9616 ( .A1(n10953), .A2(n10820), .ZN(n10823) );
  INV_X1 U9617 ( .A(n12014), .ZN(n11971) );
  AND2_X1 U9618 ( .A1(n10510), .A2(n10509), .ZN(n12018) );
  AND2_X1 U9619 ( .A1(n10739), .A2(n7984), .ZN(n8812) );
  AND4_X1 U9620 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n12522)
         );
  INV_X1 U9621 ( .A(n15258), .ZN(n15262) );
  INV_X1 U9622 ( .A(n12387), .ZN(n15296) );
  OAI21_X1 U9623 ( .B1(n12472), .B2(n15347), .A(n12471), .ZN(n12647) );
  INV_X1 U9624 ( .A(n15340), .ZN(n15321) );
  NAND2_X1 U9625 ( .A1(n7917), .A2(n8830), .ZN(n15352) );
  NOR2_X1 U9626 ( .A1(n10750), .A2(n15356), .ZN(n15333) );
  INV_X1 U9627 ( .A(n10511), .ZN(n10751) );
  AND3_X1 U9628 ( .A1(n8829), .A2(n8828), .A3(n8827), .ZN(n10747) );
  NAND2_X1 U9629 ( .A1(n10965), .A2(n10817), .ZN(n15406) );
  AND2_X1 U9630 ( .A1(n10965), .A2(n15356), .ZN(n15400) );
  AND2_X1 U9631 ( .A1(n12704), .A2(n12703), .ZN(n15361) );
  NOR2_X1 U9632 ( .A1(n8008), .A2(n10199), .ZN(n10209) );
  INV_X1 U9633 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7910) );
  NOR2_X1 U9634 ( .A1(n7747), .A2(n7759), .ZN(n12341) );
  INV_X1 U9635 ( .A(n15214), .ZN(n11127) );
  NOR2_X1 U9636 ( .A1(n9858), .A2(n9857), .ZN(n10056) );
  OR2_X1 U9637 ( .A1(n10057), .A2(n10056), .ZN(n10084) );
  INV_X1 U9638 ( .A(n15001), .ZN(n14976) );
  AND2_X1 U9639 ( .A1(n8795), .A2(n8794), .ZN(n13065) );
  AND2_X1 U9640 ( .A1(n9809), .A2(n9808), .ZN(n13204) );
  INV_X1 U9641 ( .A(n9818), .ZN(n10836) );
  INV_X1 U9642 ( .A(n13236), .ZN(n15027) );
  INV_X1 U9643 ( .A(n13246), .ZN(n15035) );
  INV_X1 U9644 ( .A(n15084), .ZN(n10313) );
  AND2_X1 U9645 ( .A1(n15119), .A2(n15139), .ZN(n13351) );
  INV_X1 U9646 ( .A(n15119), .ZN(n15143) );
  INV_X1 U9647 ( .A(n13351), .ZN(n15151) );
  AND2_X1 U9648 ( .A1(n8760), .A2(n13387), .ZN(n15051) );
  AND2_X1 U9649 ( .A1(n8766), .A2(n8765), .ZN(n15084) );
  AND2_X1 U9650 ( .A1(n8252), .A2(n8268), .ZN(n10076) );
  NAND2_X1 U9651 ( .A1(n9581), .A2(n9570), .ZN(n10030) );
  NOR2_X1 U9652 ( .A1(n9245), .A2(n9239), .ZN(n9269) );
  AND2_X1 U9653 ( .A1(n14733), .A2(n14771), .ZN(n13901) );
  AND2_X1 U9654 ( .A1(n9922), .A2(n9921), .ZN(n10315) );
  AND2_X1 U9655 ( .A1(n9342), .A2(n9341), .ZN(n14239) );
  AND4_X1 U9656 ( .A1(n9275), .A2(n9274), .A3(n9273), .A4(n9272), .ZN(n14661)
         );
  AND2_X1 U9657 ( .A1(n10042), .A2(n10041), .ZN(n10094) );
  INV_X1 U9658 ( .A(n14750), .ZN(n13984) );
  INV_X1 U9659 ( .A(n14036), .ZN(n14748) );
  INV_X1 U9660 ( .A(n10687), .ZN(n14039) );
  INV_X1 U9661 ( .A(n14177), .ZN(n14175) );
  XNOR2_X1 U9662 ( .A(n14086), .B(n14085), .ZN(n14083) );
  INV_X1 U9663 ( .A(n14288), .ZN(n14771) );
  INV_X1 U9664 ( .A(n14299), .ZN(n14816) );
  INV_X1 U9665 ( .A(n14323), .ZN(n14828) );
  AND3_X1 U9666 ( .A1(n9949), .A2(n10425), .A3(n9948), .ZN(n10452) );
  INV_X1 U9667 ( .A(n14049), .ZN(n14325) );
  AND2_X1 U9668 ( .A1(n10988), .A2(n14401), .ZN(n14420) );
  INV_X1 U9669 ( .A(n14420), .ZN(n14922) );
  AND2_X1 U9670 ( .A1(n9950), .A2(n9949), .ZN(n10318) );
  NAND2_X1 U9671 ( .A1(n9907), .A2(n9906), .ZN(n10007) );
  AND2_X1 U9672 ( .A1(n9095), .A2(n9113), .ZN(n10105) );
  OAI21_X1 U9673 ( .B1(n14544), .B2(n14999), .A(n14593), .ZN(n14701) );
  AND2_X1 U9674 ( .A1(n10589), .A2(n10588), .ZN(n15293) );
  INV_X1 U9675 ( .A(n12018), .ZN(n11979) );
  AND2_X1 U9676 ( .A1(n10739), .A2(n8820), .ZN(n12037) );
  INV_X1 U9677 ( .A(n12607), .ZN(n12251) );
  INV_X1 U9678 ( .A(n15285), .ZN(n15176) );
  AND2_X1 U9679 ( .A1(n12582), .A2(n12581), .ZN(n12683) );
  OR2_X1 U9680 ( .A1(n10748), .A2(n15363), .ZN(n15316) );
  NAND2_X1 U9681 ( .A1(n15424), .A2(n14625), .ZN(n12694) );
  AND2_X2 U9682 ( .A1(n10747), .A2(n8835), .ZN(n15424) );
  INV_X2 U9683 ( .A(n15412), .ZN(n15411) );
  CLKBUF_X1 U9684 ( .A(n10209), .Z(n10225) );
  INV_X1 U9685 ( .A(SI_23_), .ZN(n11190) );
  INV_X1 U9686 ( .A(SI_17_), .ZN(n10359) );
  NAND2_X1 U9687 ( .A1(n9981), .A2(P3_U3151), .ZN(n14574) );
  INV_X1 U9688 ( .A(n10640), .ZN(n15098) );
  OR2_X1 U9689 ( .A1(n9854), .A2(n9853), .ZN(n9855) );
  NAND2_X1 U9690 ( .A1(n8639), .A2(n8638), .ZN(n12966) );
  NAND2_X1 U9691 ( .A1(n8523), .A2(n8522), .ZN(n12971) );
  NAND2_X1 U9692 ( .A1(n10084), .A2(n10058), .ZN(n15014) );
  OR2_X1 U9693 ( .A1(n15038), .A2(n9844), .ZN(n15023) );
  AOI21_X2 U9694 ( .B1(n15143), .B2(n15048), .A(n10651), .ZN(n13246) );
  NAND2_X1 U9695 ( .A1(n15088), .A2(n8799), .ZN(n15050) );
  AND3_X1 U9696 ( .A1(n15109), .A2(n15108), .A3(n15107), .ZN(n15158) );
  OR2_X1 U9697 ( .A1(n10342), .A2(n15084), .ZN(n15153) );
  NOR2_X1 U9698 ( .A1(n15051), .A2(n15086), .ZN(n15079) );
  INV_X1 U9699 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n13489) );
  INV_X1 U9700 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10252) );
  INV_X1 U9701 ( .A(n11605), .ZN(n14598) );
  INV_X1 U9702 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n10341) );
  OAI21_X1 U9703 ( .B1(n14242), .B2(n9374), .A(n9355), .ZN(n14252) );
  NAND2_X1 U9704 ( .A1(n10094), .A2(n14454), .ZN(n14036) );
  NAND2_X1 U9705 ( .A1(n10040), .A2(n10041), .ZN(n14756) );
  OR2_X1 U9706 ( .A1(n14833), .A2(n14039), .ZN(n14308) );
  OR2_X1 U9707 ( .A1(n14833), .A2(n9954), .ZN(n14299) );
  INV_X1 U9708 ( .A(n14774), .ZN(n14315) );
  OR2_X1 U9709 ( .A1(n14833), .A2(n14130), .ZN(n14323) );
  INV_X2 U9710 ( .A(n14774), .ZN(n14833) );
  AND2_X2 U9711 ( .A1(n10453), .A2(n10452), .ZN(n14940) );
  AND4_X1 U9712 ( .A1(n14904), .A2(n14903), .A3(n14902), .A4(n14901), .ZN(
        n14932) );
  AND2_X2 U9713 ( .A1(n10318), .A2(n10453), .ZN(n14925) );
  AND2_X2 U9714 ( .A1(n10008), .A2(n10007), .ZN(n14864) );
  INV_X1 U9715 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11814) );
  INV_X1 U9716 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n13502) );
  INV_X1 U9717 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10175) );
  XNOR2_X1 U9718 ( .A(n14526), .B(n14525), .ZN(n14582) );
  INV_X2 U9719 ( .A(n12259), .ZN(P3_U3897) );
  OAI21_X1 U9720 ( .B1(n8039), .B2(n15412), .A(n8038), .ZN(P3_U3455) );
  INV_X1 U9721 ( .A(n12987), .ZN(P2_U3947) );
  INV_X1 U9722 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U9723 ( .A1(n9982), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7447) );
  NAND2_X1 U9724 ( .A1(n7521), .A2(n7447), .ZN(n7535) );
  XNOR2_X1 U9725 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7534) );
  NAND2_X1 U9726 ( .A1(n7535), .A2(n7534), .ZN(n7449) );
  INV_X1 U9727 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9998) );
  NAND2_X1 U9728 ( .A1(n9998), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7448) );
  NAND2_X1 U9729 ( .A1(n7449), .A2(n7448), .ZN(n7548) );
  NAND2_X1 U9730 ( .A1(n7548), .A2(n7547), .ZN(n7452) );
  INV_X1 U9731 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U9732 ( .A1(n7450), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n7451) );
  INV_X1 U9733 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U9734 ( .A1(n9994), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7453) );
  INV_X1 U9735 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9996) );
  AND2_X1 U9736 ( .A1(n10002), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7455) );
  NAND2_X1 U9737 ( .A1(n10000), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7454) );
  NAND2_X1 U9738 ( .A1(n7610), .A2(n7611), .ZN(n7457) );
  NAND2_X1 U9739 ( .A1(n10004), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7456) );
  NAND2_X1 U9740 ( .A1(n10017), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7458) );
  XNOR2_X1 U9741 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7642) );
  INV_X1 U9742 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10020) );
  INV_X1 U9743 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U9744 ( .A1(n10024), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n7459) );
  AND2_X1 U9745 ( .A1(n10051), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7462) );
  NAND2_X1 U9746 ( .A1(n10053), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n7461) );
  NAND2_X1 U9747 ( .A1(n10175), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n7464) );
  NAND2_X1 U9748 ( .A1(n10174), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n7463) );
  NAND2_X1 U9749 ( .A1(n7464), .A2(n7463), .ZN(n7695) );
  NAND2_X1 U9750 ( .A1(n7465), .A2(n13631), .ZN(n7466) );
  NAND2_X1 U9751 ( .A1(n10386), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9752 ( .A1(n7469), .A2(n7468), .ZN(n7728) );
  XNOR2_X1 U9753 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n7726) );
  NAND2_X1 U9754 ( .A1(n7728), .A2(n7726), .ZN(n7471) );
  NAND2_X1 U9755 ( .A1(n10443), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n7470) );
  NAND2_X1 U9756 ( .A1(n7471), .A2(n7470), .ZN(n7742) );
  XNOR2_X1 U9757 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n7740) );
  NAND2_X1 U9758 ( .A1(n7742), .A2(n7740), .ZN(n7474) );
  AOI22_X1 U9759 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10422), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n13502), .ZN(n7757) );
  AOI22_X1 U9760 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10537), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n13629), .ZN(n7782) );
  INV_X1 U9761 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10686) );
  AOI22_X1 U9762 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n10686), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n13526), .ZN(n7796) );
  NAND2_X1 U9763 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n7477), .ZN(n7478) );
  INV_X1 U9764 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10811) );
  AOI22_X1 U9765 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(n10811), .B2(n13489), .ZN(n7820) );
  INV_X1 U9766 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8117) );
  AOI22_X1 U9767 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n11056), .B2(n8117), .ZN(n7832) );
  INV_X1 U9768 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U9769 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n10341), .B2(n10388), .ZN(n7843) );
  INV_X1 U9770 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11739) );
  XNOR2_X1 U9771 ( .A(n7855), .B(n11739), .ZN(n7856) );
  XOR2_X1 U9772 ( .A(n11741), .B(n7856), .Z(n11561) );
  NOR2_X1 U9773 ( .A1(P3_IR_REG_4__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n7481) );
  NOR2_X1 U9774 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n7480) );
  NOR3_X1 U9775 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .A3(
        P3_IR_REG_11__SCAN_IN), .ZN(n7482) );
  XNOR2_X2 U9776 ( .A(n7493), .B(n7492), .ZN(n7986) );
  NAND2_X1 U9777 ( .A1(n11561), .A2(n12027), .ZN(n7497) );
  INV_X1 U9778 ( .A(SI_24_), .ZN(n11558) );
  NOR2_X2 U9779 ( .A1(n7501), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n7503) );
  NAND2_X1 U9780 ( .A1(n7501), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7502) );
  MUX2_X1 U9781 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7502), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7504) );
  INV_X1 U9782 ( .A(n7503), .ZN(n12764) );
  INV_X1 U9783 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12648) );
  NOR2_X1 U9784 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7571) );
  INV_X1 U9785 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7570) );
  NAND2_X1 U9786 ( .A1(n7571), .A2(n7570), .ZN(n7589) );
  NOR2_X1 U9787 ( .A1(n7602), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7619) );
  NAND2_X1 U9788 ( .A1(n7636), .A2(n7635), .ZN(n7654) );
  NAND2_X1 U9789 ( .A1(n7700), .A2(n7699), .ZN(n7719) );
  INV_X1 U9790 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n7750) );
  NAND2_X1 U9791 ( .A1(n7764), .A2(n7763), .ZN(n7789) );
  INV_X1 U9792 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U9793 ( .A1(n7824), .A2(n11939), .ZN(n7836) );
  OR2_X1 U9794 ( .A1(n7446), .A2(n7861), .ZN(n12475) );
  NAND2_X1 U9795 ( .A1(n12475), .A2(n6551), .ZN(n7508) );
  AOI22_X1 U9796 ( .A1(n10733), .A2(P3_REG0_REG_24__SCAN_IN), .B1(n10734), 
        .B2(P3_REG2_REG_24__SCAN_IN), .ZN(n7507) );
  OAI211_X1 U9797 ( .C1(n7604), .C2(n12648), .A(n7508), .B(n7507), .ZN(n12484)
         );
  NAND2_X1 U9798 ( .A1(n10734), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7513) );
  NAND2_X1 U9799 ( .A1(n6547), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U9800 ( .A1(n7588), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7511) );
  INV_X1 U9801 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n7509) );
  XNOR2_X1 U9802 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .ZN(n7514) );
  NAND2_X1 U9803 ( .A1(n8043), .A2(SI_0_), .ZN(n8187) );
  OAI21_X1 U9804 ( .B1(n9981), .B2(n7514), .A(n8187), .ZN(n12781) );
  NAND2_X1 U9805 ( .A1(n6551), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9806 ( .A1(n7588), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7519) );
  INV_X1 U9807 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10593) );
  INV_X1 U9808 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n7516) );
  OAI21_X1 U9809 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7524) );
  INV_X1 U9810 ( .A(n7524), .ZN(n9964) );
  OR2_X1 U9811 ( .A1(n12035), .A2(n9964), .ZN(n7529) );
  INV_X1 U9812 ( .A(SI_1_), .ZN(n9963) );
  OR2_X1 U9813 ( .A1(n7546), .A2(n9963), .ZN(n7527) );
  INV_X1 U9814 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n7526) );
  AND2_X1 U9815 ( .A1(n7527), .A2(n7442), .ZN(n7528) );
  NAND2_X1 U9816 ( .A1(n7529), .A2(n7528), .ZN(n12706) );
  INV_X1 U9817 ( .A(n12706), .ZN(n10830) );
  NAND2_X1 U9818 ( .A1(n10506), .A2(n10830), .ZN(n12078) );
  NAND2_X1 U9819 ( .A1(n15341), .A2(n12706), .ZN(n12081) );
  NAND2_X1 U9820 ( .A1(n10821), .A2(n12081), .ZN(n15337) );
  NAND2_X1 U9821 ( .A1(n6547), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7533) );
  NAND2_X1 U9822 ( .A1(n7588), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7532) );
  INV_X1 U9823 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10600) );
  INV_X1 U9824 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n7531) );
  OR2_X1 U9825 ( .A1(n7546), .A2(SI_2_), .ZN(n7540) );
  XNOR2_X1 U9826 ( .A(n7535), .B(n7534), .ZN(n9979) );
  OR2_X1 U9827 ( .A1(n12035), .A2(n9979), .ZN(n7539) );
  OR2_X1 U9828 ( .A1(n6550), .A2(n6552), .ZN(n7538) );
  INV_X1 U9829 ( .A(n15342), .ZN(n15345) );
  NAND2_X1 U9830 ( .A1(n15337), .A2(n15345), .ZN(n15336) );
  NAND2_X1 U9831 ( .A1(n15336), .A2(n12079), .ZN(n15318) );
  NAND2_X1 U9832 ( .A1(n7588), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7545) );
  INV_X1 U9833 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15332) );
  NAND2_X1 U9834 ( .A1(n6551), .A2(n15332), .ZN(n7544) );
  INV_X1 U9835 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n11079) );
  OR2_X1 U9836 ( .A1(n7826), .A2(n11079), .ZN(n7543) );
  INV_X1 U9837 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n7541) );
  OR2_X1 U9838 ( .A1(n7558), .A2(n7541), .ZN(n7542) );
  OR2_X1 U9839 ( .A1(n12033), .A2(SI_3_), .ZN(n7554) );
  XNOR2_X1 U9840 ( .A(n7548), .B(n7547), .ZN(n9977) );
  OR2_X1 U9841 ( .A1(n12035), .A2(n9977), .ZN(n7553) );
  NAND2_X1 U9842 ( .A1(n7549), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7550) );
  MUX2_X1 U9843 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7550), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n7551) );
  AND2_X1 U9844 ( .A1(n7551), .A2(n7627), .ZN(n15180) );
  OR2_X1 U9845 ( .A1(n10577), .A2(n15180), .ZN(n7552) );
  NAND2_X1 U9846 ( .A1(n15339), .A2(n11037), .ZN(n12086) );
  NAND2_X1 U9847 ( .A1(n12258), .A2(n15331), .ZN(n12084) );
  AND2_X2 U9848 ( .A1(n12086), .A2(n12084), .ZN(n7919) );
  NAND2_X1 U9849 ( .A1(n15318), .A2(n7919), .ZN(n7555) );
  NAND2_X1 U9850 ( .A1(n7555), .A2(n12086), .ZN(n11403) );
  AND2_X1 U9851 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7556) );
  OR2_X1 U9852 ( .A1(n7556), .A2(n7571), .ZN(n11412) );
  NAND2_X1 U9853 ( .A1(n6547), .A2(n11412), .ZN(n7562) );
  NAND2_X1 U9854 ( .A1(n7588), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7561) );
  OR2_X1 U9855 ( .A1(n7826), .A2(n11065), .ZN(n7560) );
  INV_X1 U9856 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n7557) );
  OR2_X1 U9857 ( .A1(n7558), .A2(n7557), .ZN(n7559) );
  OR2_X1 U9858 ( .A1(n7546), .A2(SI_4_), .ZN(n7569) );
  XNOR2_X1 U9859 ( .A(n7564), .B(n7563), .ZN(n9973) );
  OR2_X1 U9860 ( .A1(n12035), .A2(n9973), .ZN(n7568) );
  NAND2_X1 U9861 ( .A1(n7627), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7566) );
  INV_X1 U9862 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7565) );
  XNOR2_X1 U9863 ( .A(n7566), .B(n7565), .ZN(n15195) );
  INV_X1 U9864 ( .A(n15195), .ZN(n11125) );
  OR2_X1 U9865 ( .A1(n6550), .A2(n11125), .ZN(n7567) );
  NAND2_X1 U9866 ( .A1(n11242), .A2(n11411), .ZN(n12095) );
  NAND2_X1 U9867 ( .A1(n15320), .A2(n11272), .ZN(n12094) );
  NAND2_X1 U9868 ( .A1(n12095), .A2(n12094), .ZN(n11406) );
  INV_X1 U9869 ( .A(n11406), .ZN(n12092) );
  NAND2_X1 U9870 ( .A1(n11402), .A2(n12095), .ZN(n11238) );
  NAND2_X1 U9871 ( .A1(n10734), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U9872 ( .A1(n7588), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7575) );
  OR2_X1 U9873 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  NAND2_X1 U9874 ( .A1(n7589), .A2(n7572), .ZN(n11385) );
  NAND2_X1 U9875 ( .A1(n6547), .A2(n11385), .ZN(n7574) );
  NAND2_X1 U9876 ( .A1(n10733), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7573) );
  NAND4_X1 U9877 ( .A1(n7576), .A2(n7575), .A3(n7574), .A4(n7573), .ZN(n12257)
         );
  INV_X1 U9878 ( .A(n12257), .ZN(n11567) );
  OR2_X1 U9879 ( .A1(n12033), .A2(SI_5_), .ZN(n7586) );
  XNOR2_X1 U9880 ( .A(n7578), .B(n7577), .ZN(n9975) );
  OR2_X1 U9881 ( .A1(n12035), .A2(n9975), .ZN(n7585) );
  NOR2_X1 U9882 ( .A1(n7627), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7581) );
  NOR2_X1 U9883 ( .A1(n7581), .A2(n8002), .ZN(n7579) );
  MUX2_X1 U9884 ( .A(n8002), .B(n7579), .S(P3_IR_REG_5__SCAN_IN), .Z(n7583) );
  INV_X1 U9885 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7580) );
  NAND2_X1 U9886 ( .A1(n7581), .A2(n7580), .ZN(n7613) );
  INV_X1 U9887 ( .A(n7613), .ZN(n7582) );
  OR2_X1 U9888 ( .A1(n6550), .A2(n11127), .ZN(n7584) );
  NAND2_X1 U9889 ( .A1(n11567), .A2(n11386), .ZN(n12100) );
  INV_X1 U9890 ( .A(n11386), .ZN(n11397) );
  NAND2_X1 U9891 ( .A1(n12257), .A2(n11397), .ZN(n12099) );
  NAND2_X1 U9892 ( .A1(n12100), .A2(n12099), .ZN(n11240) );
  INV_X1 U9893 ( .A(n11240), .ZN(n12097) );
  NAND2_X1 U9894 ( .A1(n11238), .A2(n12097), .ZN(n7587) );
  NAND2_X1 U9895 ( .A1(n7587), .A2(n12100), .ZN(n11546) );
  NAND2_X1 U9896 ( .A1(n7588), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7595) );
  NAND2_X1 U9897 ( .A1(n7589), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7590) );
  NAND2_X1 U9898 ( .A1(n7602), .A2(n7590), .ZN(n11681) );
  NAND2_X1 U9899 ( .A1(n6547), .A2(n11681), .ZN(n7594) );
  INV_X1 U9900 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11093) );
  OR2_X1 U9901 ( .A1(n7826), .A2(n11093), .ZN(n7593) );
  INV_X1 U9902 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n7591) );
  OR2_X1 U9903 ( .A1(n7558), .A2(n7591), .ZN(n7592) );
  NAND2_X1 U9904 ( .A1(n7613), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7596) );
  XNOR2_X1 U9905 ( .A(n7596), .B(P3_IR_REG_6__SCAN_IN), .ZN(n11129) );
  XNOR2_X1 U9906 ( .A(n10002), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n7597) );
  XNOR2_X1 U9907 ( .A(n7598), .B(n7597), .ZN(n9966) );
  OR2_X1 U9908 ( .A1(n12035), .A2(n9966), .ZN(n7600) );
  INV_X1 U9909 ( .A(SI_6_), .ZN(n9965) );
  OR2_X1 U9910 ( .A1(n12033), .A2(n9965), .ZN(n7599) );
  OAI211_X1 U9911 ( .C1(n6550), .C2(n15231), .A(n7600), .B(n7599), .ZN(n11568)
         );
  NAND2_X1 U9912 ( .A1(n11667), .A2(n11568), .ZN(n12106) );
  INV_X1 U9913 ( .A(n11568), .ZN(n11687) );
  NAND2_X1 U9914 ( .A1(n12256), .A2(n11687), .ZN(n12105) );
  NAND2_X1 U9915 ( .A1(n12106), .A2(n12105), .ZN(n11547) );
  INV_X1 U9916 ( .A(n11547), .ZN(n12044) );
  NAND2_X1 U9917 ( .A1(n11546), .A2(n12044), .ZN(n7601) );
  NAND2_X1 U9918 ( .A1(n7601), .A2(n12106), .ZN(n11463) );
  AND2_X1 U9919 ( .A1(n7602), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7603) );
  OR2_X1 U9920 ( .A1(n7603), .A2(n7619), .ZN(n11673) );
  NAND2_X1 U9921 ( .A1(n6547), .A2(n11673), .ZN(n7609) );
  NAND2_X1 U9922 ( .A1(n7588), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7608) );
  INV_X1 U9923 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n7605) );
  OR2_X1 U9924 ( .A1(n7558), .A2(n7605), .ZN(n7607) );
  INV_X1 U9925 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n11099) );
  OR2_X1 U9926 ( .A1(n7826), .A2(n11099), .ZN(n7606) );
  OR2_X1 U9927 ( .A1(n12033), .A2(SI_7_), .ZN(n7618) );
  INV_X1 U9928 ( .A(n7611), .ZN(n7612) );
  XNOR2_X1 U9929 ( .A(n7610), .B(n7612), .ZN(n9971) );
  OR2_X1 U9930 ( .A1(n12035), .A2(n9971), .ZN(n7617) );
  OR2_X1 U9931 ( .A1(n7613), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U9932 ( .A1(n7625), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7615) );
  INV_X1 U9933 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7614) );
  XNOR2_X1 U9934 ( .A(n7615), .B(n7614), .ZN(n15249) );
  INV_X1 U9935 ( .A(n15249), .ZN(n11131) );
  OR2_X1 U9936 ( .A1(n10577), .A2(n11131), .ZN(n7616) );
  NAND2_X1 U9937 ( .A1(n11746), .A2(n7935), .ZN(n12110) );
  INV_X1 U9938 ( .A(n7935), .ZN(n11670) );
  NAND2_X1 U9939 ( .A1(n12255), .A2(n11670), .ZN(n12111) );
  NAND2_X1 U9940 ( .A1(n10733), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7624) );
  NAND2_X1 U9941 ( .A1(n10734), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7623) );
  NOR2_X1 U9942 ( .A1(n7619), .A2(n11749), .ZN(n7620) );
  OR2_X1 U9943 ( .A1(n7636), .A2(n7620), .ZN(n11753) );
  NAND2_X1 U9944 ( .A1(n6547), .A2(n11753), .ZN(n7622) );
  NAND2_X1 U9945 ( .A1(n7588), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7621) );
  NAND4_X1 U9946 ( .A1(n7624), .A2(n7623), .A3(n7622), .A4(n7621), .ZN(n12254)
         );
  INV_X1 U9947 ( .A(n12254), .ZN(n11671) );
  OAI21_X1 U9948 ( .B1(n7625), .B2(P3_IR_REG_7__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7626) );
  MUX2_X1 U9949 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7626), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n7630) );
  INV_X1 U9950 ( .A(n7627), .ZN(n7629) );
  NAND2_X1 U9951 ( .A1(n7629), .A2(n7628), .ZN(n7646) );
  NAND2_X1 U9952 ( .A1(n7630), .A2(n7646), .ZN(n15268) );
  XNOR2_X1 U9953 ( .A(n7632), .B(n7631), .ZN(n9967) );
  OR2_X1 U9954 ( .A1(n12035), .A2(n9967), .ZN(n7634) );
  INV_X1 U9955 ( .A(SI_8_), .ZN(n9968) );
  OR2_X1 U9956 ( .A1(n12033), .A2(n9968), .ZN(n7633) );
  OAI211_X1 U9957 ( .C1(n10577), .C2(n15268), .A(n7634), .B(n7633), .ZN(n11565) );
  NAND2_X1 U9958 ( .A1(n11671), .A2(n11565), .ZN(n12116) );
  INV_X1 U9959 ( .A(n11565), .ZN(n11750) );
  NAND2_X1 U9960 ( .A1(n12254), .A2(n11750), .ZN(n12115) );
  NAND2_X1 U9961 ( .A1(n10734), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U9962 ( .A1(n7980), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7640) );
  OR2_X1 U9963 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  NAND2_X1 U9964 ( .A1(n7654), .A2(n7637), .ZN(n11563) );
  NAND2_X1 U9965 ( .A1(n6551), .A2(n11563), .ZN(n7639) );
  NAND2_X1 U9966 ( .A1(n10733), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7638) );
  NAND4_X1 U9967 ( .A1(n7641), .A2(n7640), .A3(n7639), .A4(n7638), .ZN(n15303)
         );
  OR2_X1 U9968 ( .A1(n12033), .A2(SI_9_), .ZN(n7650) );
  INV_X1 U9969 ( .A(n7642), .ZN(n7643) );
  XNOR2_X1 U9970 ( .A(n7644), .B(n7643), .ZN(n9969) );
  OR2_X1 U9971 ( .A1(n12035), .A2(n9969), .ZN(n7649) );
  NAND2_X1 U9972 ( .A1(n7646), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7645) );
  MUX2_X1 U9973 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7645), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7647) );
  OR2_X1 U9974 ( .A1(n6550), .A2(n11135), .ZN(n7648) );
  INV_X1 U9975 ( .A(n12120), .ZN(n11578) );
  NAND2_X1 U9976 ( .A1(n15303), .A2(n11578), .ZN(n7651) );
  NAND2_X1 U9977 ( .A1(n11484), .A2(n7651), .ZN(n7653) );
  INV_X1 U9978 ( .A(n15303), .ZN(n11751) );
  NAND2_X1 U9979 ( .A1(n11751), .A2(n12120), .ZN(n7652) );
  NAND2_X1 U9980 ( .A1(n7653), .A2(n7652), .ZN(n15302) );
  NAND2_X1 U9981 ( .A1(n7654), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7655) );
  AND2_X1 U9982 ( .A1(n7669), .A2(n7655), .ZN(n15317) );
  INV_X1 U9983 ( .A(n15317), .ZN(n7656) );
  NAND2_X1 U9984 ( .A1(n6547), .A2(n7656), .ZN(n7661) );
  NAND2_X1 U9985 ( .A1(n7980), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7660) );
  INV_X1 U9986 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n7657) );
  OR2_X1 U9987 ( .A1(n7558), .A2(n7657), .ZN(n7659) );
  INV_X1 U9988 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n15311) );
  OR2_X1 U9989 ( .A1(n7826), .A2(n15311), .ZN(n7658) );
  XNOR2_X1 U9990 ( .A(n7662), .B(n6671), .ZN(n9983) );
  OR2_X1 U9991 ( .A1(n12035), .A2(n9983), .ZN(n7667) );
  OR2_X1 U9992 ( .A1(n12033), .A2(SI_10_), .ZN(n7666) );
  NAND2_X1 U9993 ( .A1(n7677), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7664) );
  INV_X1 U9994 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7663) );
  XNOR2_X1 U9995 ( .A(n7664), .B(n7663), .ZN(n11443) );
  INV_X1 U9996 ( .A(n11443), .ZN(n11117) );
  OR2_X1 U9997 ( .A1(n10577), .A2(n11117), .ZN(n7665) );
  NAND2_X1 U9998 ( .A1(n12253), .A2(n15405), .ZN(n12134) );
  NAND2_X1 U9999 ( .A1(n15302), .A2(n12134), .ZN(n7668) );
  NAND2_X1 U10000 ( .A1(n11727), .A2(n11634), .ZN(n12127) );
  NAND2_X1 U10001 ( .A1(n7980), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U10002 ( .A1(n7669), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7670) );
  NAND2_X1 U10003 ( .A1(n7684), .A2(n7670), .ZN(n11732) );
  NAND2_X1 U10004 ( .A1(n6551), .A2(n11732), .ZN(n7675) );
  INV_X1 U10005 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n7671) );
  OR2_X1 U10006 ( .A1(n7826), .A2(n7671), .ZN(n7674) );
  INV_X1 U10007 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n7672) );
  OR2_X1 U10008 ( .A1(n7558), .A2(n7672), .ZN(n7673) );
  OAI21_X1 U10009 ( .B1(n7677), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7679) );
  INV_X1 U10010 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7678) );
  XNOR2_X1 U10011 ( .A(n7679), .B(n7678), .ZN(n14573) );
  INV_X1 U10012 ( .A(n14573), .ZN(n11447) );
  XNOR2_X1 U10013 ( .A(n10053), .B(P2_DATAO_REG_11__SCAN_IN), .ZN(n7680) );
  XNOR2_X1 U10014 ( .A(n7681), .B(n7680), .ZN(n14571) );
  OR2_X1 U10015 ( .A1(n12035), .A2(n14571), .ZN(n7683) );
  OR2_X1 U10016 ( .A1(n12033), .A2(SI_11_), .ZN(n7682) );
  OAI211_X1 U10017 ( .C1(n11447), .C2(n6550), .A(n7683), .B(n7682), .ZN(n11731) );
  INV_X1 U10018 ( .A(n11731), .ZN(n11717) );
  NAND2_X1 U10019 ( .A1(n11791), .A2(n11717), .ZN(n12137) );
  NAND2_X1 U10020 ( .A1(n15304), .A2(n11731), .ZN(n12128) );
  NAND2_X1 U10021 ( .A1(n7980), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7690) );
  AND2_X1 U10022 ( .A1(n7684), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n7685) );
  OR2_X1 U10023 ( .A1(n7685), .A2(n7700), .ZN(n11764) );
  NAND2_X1 U10024 ( .A1(n6547), .A2(n11764), .ZN(n7689) );
  INV_X1 U10025 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11765) );
  OR2_X1 U10026 ( .A1(n7826), .A2(n11765), .ZN(n7688) );
  INV_X1 U10027 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n7686) );
  OR2_X1 U10028 ( .A1(n7558), .A2(n7686), .ZN(n7687) );
  NOR2_X1 U10029 ( .A1(n7691), .A2(n8002), .ZN(n7692) );
  MUX2_X1 U10030 ( .A(n8002), .B(n7692), .S(P3_IR_REG_12__SCAN_IN), .Z(n7694)
         );
  OR2_X1 U10031 ( .A1(n7694), .A2(n7693), .ZN(n14580) );
  OR2_X1 U10032 ( .A1(n12033), .A2(n14575), .ZN(n7698) );
  XNOR2_X1 U10033 ( .A(n7696), .B(n7695), .ZN(n14577) );
  OR2_X1 U10034 ( .A1(n12035), .A2(n14577), .ZN(n7697) );
  OAI211_X1 U10035 ( .C1(n10577), .C2(n14580), .A(n7698), .B(n7697), .ZN(
        n11793) );
  INV_X1 U10036 ( .A(n11793), .ZN(n11785) );
  NAND2_X1 U10037 ( .A1(n12252), .A2(n11785), .ZN(n12130) );
  AND2_X1 U10038 ( .A1(n12135), .A2(n12130), .ZN(n11775) );
  NAND2_X1 U10039 ( .A1(n10733), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7705) );
  NAND2_X1 U10040 ( .A1(n10734), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7704) );
  OR2_X1 U10041 ( .A1(n7700), .A2(n7699), .ZN(n7701) );
  NAND2_X1 U10042 ( .A1(n7719), .A2(n7701), .ZN(n11773) );
  NAND2_X1 U10043 ( .A1(n6547), .A2(n11773), .ZN(n7703) );
  NAND2_X1 U10044 ( .A1(n7980), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7702) );
  NAND4_X1 U10045 ( .A1(n7705), .A2(n7704), .A3(n7703), .A4(n7702), .ZN(n12618) );
  OAI21_X1 U10046 ( .B1(n7707), .B2(P1_DATAO_REG_13__SCAN_IN), .A(n7706), .ZN(
        n10028) );
  NAND2_X1 U10047 ( .A1(n10028), .A2(n12027), .ZN(n7711) );
  INV_X1 U10048 ( .A(n10577), .ZN(n7708) );
  OR2_X1 U10049 ( .A1(n7693), .A2(n8002), .ZN(n7709) );
  XNOR2_X1 U10050 ( .A(n7709), .B(n7714), .ZN(n12273) );
  AOI22_X1 U10051 ( .A1(n7800), .A2(n10029), .B1(n7708), .B2(n12273), .ZN(
        n7710) );
  NAND2_X1 U10052 ( .A1(n12618), .A2(n14629), .ZN(n12146) );
  AND2_X1 U10053 ( .A1(n11775), .A2(n12146), .ZN(n12561) );
  XNOR2_X1 U10054 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n7713) );
  XNOR2_X1 U10055 ( .A(n7712), .B(n7713), .ZN(n10119) );
  NAND2_X1 U10056 ( .A1(n10119), .A2(n12027), .ZN(n7718) );
  NAND2_X1 U10057 ( .A1(n7693), .A2(n7714), .ZN(n7729) );
  NAND2_X1 U10058 ( .A1(n7729), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7716) );
  XNOR2_X1 U10059 ( .A(n7716), .B(n7715), .ZN(n12293) );
  AOI22_X1 U10060 ( .A1(n7800), .A2(n10120), .B1(n7708), .B2(n12293), .ZN(
        n7717) );
  NAND2_X1 U10061 ( .A1(n7719), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U10062 ( .A1(n7733), .A2(n7720), .ZN(n12621) );
  NAND2_X1 U10063 ( .A1(n6547), .A2(n12621), .ZN(n7725) );
  NAND2_X1 U10064 ( .A1(n7980), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7724) );
  INV_X1 U10065 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12759) );
  OR2_X1 U10066 ( .A1(n7558), .A2(n12759), .ZN(n7723) );
  INV_X1 U10067 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n7721) );
  OR2_X1 U10068 ( .A1(n7826), .A2(n7721), .ZN(n7722) );
  NAND2_X1 U10069 ( .A1(n12761), .A2(n11982), .ZN(n12147) );
  INV_X1 U10070 ( .A(n12147), .ZN(n12597) );
  INV_X1 U10071 ( .A(n7726), .ZN(n7727) );
  XNOR2_X1 U10072 ( .A(n7728), .B(n7727), .ZN(n14583) );
  NAND2_X1 U10073 ( .A1(n14583), .A2(n12027), .ZN(n7732) );
  NAND2_X1 U10074 ( .A1(n7743), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7730) );
  XNOR2_X1 U10075 ( .A(n7730), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12319) );
  AOI22_X1 U10076 ( .A1(n7800), .A2(SI_15_), .B1(n7708), .B2(n12319), .ZN(
        n7731) );
  NAND2_X1 U10077 ( .A1(n7732), .A2(n7731), .ZN(n12608) );
  NAND2_X1 U10078 ( .A1(n10733), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7739) );
  NAND2_X1 U10079 ( .A1(n10734), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7738) );
  INV_X1 U10080 ( .A(n7751), .ZN(n7735) );
  NAND2_X1 U10081 ( .A1(n7733), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7734) );
  NAND2_X1 U10082 ( .A1(n7735), .A2(n7734), .ZN(n12609) );
  NAND2_X1 U10083 ( .A1(n6547), .A2(n12609), .ZN(n7737) );
  NAND2_X1 U10084 ( .A1(n7980), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7736) );
  NAND4_X1 U10085 ( .A1(n7739), .A2(n7738), .A3(n7737), .A4(n7736), .ZN(n12617) );
  INV_X1 U10086 ( .A(n12617), .ZN(n7777) );
  OR2_X1 U10087 ( .A1(n12608), .A2(n7777), .ZN(n12149) );
  INV_X1 U10088 ( .A(n12149), .ZN(n7779) );
  OR2_X1 U10089 ( .A1(n12597), .A2(n7779), .ZN(n12585) );
  INV_X1 U10090 ( .A(n7740), .ZN(n7741) );
  XNOR2_X1 U10091 ( .A(n7742), .B(n7741), .ZN(n14588) );
  NAND2_X1 U10092 ( .A1(n14588), .A2(n12027), .ZN(n7749) );
  NAND2_X1 U10093 ( .A1(n7746), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7744) );
  MUX2_X1 U10094 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7744), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n7745) );
  INV_X1 U10095 ( .A(n7745), .ZN(n7747) );
  AOI22_X1 U10096 ( .A1(n7800), .A2(SI_16_), .B1(n7708), .B2(n12341), .ZN(
        n7748) );
  NAND2_X1 U10097 ( .A1(n7749), .A2(n7748), .ZN(n11955) );
  NOR2_X1 U10098 ( .A1(n7751), .A2(n7750), .ZN(n7752) );
  OR2_X1 U10099 ( .A1(n7764), .A2(n7752), .ZN(n12592) );
  NAND2_X1 U10100 ( .A1(n6551), .A2(n12592), .ZN(n7756) );
  NAND2_X1 U10101 ( .A1(n7980), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7755) );
  INV_X1 U10102 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12750) );
  OR2_X1 U10103 ( .A1(n7558), .A2(n12750), .ZN(n7754) );
  INV_X1 U10104 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12340) );
  OR2_X1 U10105 ( .A1(n7826), .A2(n12340), .ZN(n7753) );
  OR2_X1 U10106 ( .A1(n11955), .A2(n12607), .ZN(n12155) );
  NAND2_X1 U10107 ( .A1(n11955), .A2(n12607), .ZN(n12153) );
  NAND2_X1 U10108 ( .A1(n12155), .A2(n12153), .ZN(n7951) );
  OR2_X1 U10109 ( .A1(n12585), .A2(n7951), .ZN(n12565) );
  XOR2_X1 U10110 ( .A(n7758), .B(n7757), .Z(n10357) );
  INV_X1 U10111 ( .A(n7759), .ZN(n7785) );
  NAND2_X1 U10112 ( .A1(n7785), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7761) );
  INV_X1 U10113 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7760) );
  XNOR2_X1 U10114 ( .A(n7761), .B(n7760), .ZN(n12351) );
  OAI22_X1 U10115 ( .A1(n12033), .A2(n10359), .B1(n10577), .B2(n12351), .ZN(
        n7762) );
  NAND2_X1 U10116 ( .A1(n10734), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7769) );
  NAND2_X1 U10117 ( .A1(n10733), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7768) );
  OR2_X1 U10118 ( .A1(n7764), .A2(n7763), .ZN(n7765) );
  NAND2_X1 U10119 ( .A1(n7789), .A2(n7765), .ZN(n12573) );
  NAND2_X1 U10120 ( .A1(n6547), .A2(n12573), .ZN(n7767) );
  NAND2_X1 U10121 ( .A1(n7980), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7766) );
  NAND4_X1 U10122 ( .A1(n7769), .A2(n7768), .A3(n7767), .A4(n7766), .ZN(n12580) );
  NAND2_X1 U10123 ( .A1(n12749), .A2(n12580), .ZN(n12159) );
  INV_X1 U10124 ( .A(n12749), .ZN(n7954) );
  NAND2_X1 U10125 ( .A1(n7954), .A2(n12554), .ZN(n12164) );
  NAND2_X1 U10126 ( .A1(n12159), .A2(n12164), .ZN(n12569) );
  INV_X1 U10127 ( .A(n12569), .ZN(n12567) );
  OR2_X1 U10128 ( .A1(n12565), .A2(n12569), .ZN(n7775) );
  INV_X1 U10129 ( .A(n7775), .ZN(n7770) );
  AND2_X1 U10130 ( .A1(n12561), .A2(n7770), .ZN(n7776) );
  INV_X1 U10131 ( .A(n12146), .ZN(n11770) );
  NOR2_X1 U10132 ( .A1(n12618), .A2(n14629), .ZN(n12140) );
  INV_X1 U10133 ( .A(n12140), .ZN(n7773) );
  INV_X1 U10134 ( .A(n12130), .ZN(n7772) );
  NAND2_X1 U10135 ( .A1(n11799), .A2(n11793), .ZN(n12138) );
  AND2_X1 U10136 ( .A1(n12137), .A2(n12138), .ZN(n7771) );
  AND2_X1 U10137 ( .A1(n7773), .A2(n11776), .ZN(n7774) );
  AOI21_X1 U10138 ( .B1(n12562), .B2(n7776), .A(n7438), .ZN(n7781) );
  NAND2_X1 U10139 ( .A1(n11800), .A2(n12606), .ZN(n12598) );
  NAND2_X1 U10140 ( .A1(n12608), .A2(n7777), .ZN(n12152) );
  AND2_X1 U10141 ( .A1(n12598), .A2(n12152), .ZN(n7778) );
  OR2_X1 U10142 ( .A1(n7779), .A2(n7778), .ZN(n12586) );
  OR2_X1 U10143 ( .A1(n7951), .A2(n12586), .ZN(n12583) );
  AND2_X1 U10144 ( .A1(n12153), .A2(n12583), .ZN(n12566) );
  OR2_X1 U10145 ( .A1(n12569), .A2(n12566), .ZN(n7780) );
  NAND3_X1 U10146 ( .A1(n7781), .A2(n12164), .A3(n7780), .ZN(n12548) );
  INV_X1 U10147 ( .A(n7782), .ZN(n7783) );
  XNOR2_X1 U10148 ( .A(n7784), .B(n7783), .ZN(n10405) );
  NAND2_X1 U10149 ( .A1(n10405), .A2(n12027), .ZN(n7788) );
  OAI21_X1 U10150 ( .B1(n7785), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7786) );
  XNOR2_X1 U10151 ( .A(n7786), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U10152 ( .A1(n7800), .A2(SI_18_), .B1(n7708), .B2(n12378), .ZN(
        n7787) );
  NAND2_X1 U10153 ( .A1(n7788), .A2(n7787), .ZN(n7959) );
  NAND2_X1 U10154 ( .A1(n7789), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7790) );
  NAND2_X1 U10155 ( .A1(n7803), .A2(n7790), .ZN(n12556) );
  NAND2_X1 U10156 ( .A1(n6547), .A2(n12556), .ZN(n7794) );
  NAND2_X1 U10157 ( .A1(n7980), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7793) );
  INV_X1 U10158 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12743) );
  OR2_X1 U10159 ( .A1(n7558), .A2(n12743), .ZN(n7792) );
  INV_X1 U10160 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12361) );
  OR2_X1 U10161 ( .A1(n7826), .A2(n12361), .ZN(n7791) );
  OR2_X1 U10162 ( .A1(n7959), .A2(n12572), .ZN(n12161) );
  NAND2_X1 U10163 ( .A1(n7959), .A2(n12572), .ZN(n12167) );
  OR2_X1 U10164 ( .A1(n12548), .A2(n7957), .ZN(n7795) );
  XNOR2_X1 U10165 ( .A(n7797), .B(n7796), .ZN(n10447) );
  NAND2_X1 U10166 ( .A1(n10447), .A2(n12027), .ZN(n7802) );
  INV_X1 U10167 ( .A(SI_19_), .ZN(n10446) );
  NAND2_X1 U10168 ( .A1(n7798), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7799) );
  AOI22_X1 U10169 ( .A1(n7800), .A2(n10446), .B1(n7708), .B2(n12391), .ZN(
        n7801) );
  NAND2_X1 U10170 ( .A1(n7802), .A2(n7801), .ZN(n11933) );
  NAND2_X1 U10171 ( .A1(n10734), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7808) );
  NAND2_X1 U10172 ( .A1(n7980), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7807) );
  AND2_X1 U10173 ( .A1(n7803), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7804) );
  OR2_X1 U10174 ( .A1(n7804), .A2(n7814), .ZN(n12542) );
  NAND2_X1 U10175 ( .A1(n6547), .A2(n12542), .ZN(n7806) );
  NAND2_X1 U10176 ( .A1(n10733), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7805) );
  NAND4_X1 U10177 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n12520) );
  NAND2_X1 U10178 ( .A1(n11933), .A2(n12520), .ZN(n12172) );
  INV_X1 U10179 ( .A(n12172), .ZN(n7809) );
  OR2_X1 U10180 ( .A1(n11933), .A2(n12520), .ZN(n12173) );
  XNOR2_X1 U10181 ( .A(n7810), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U10182 ( .A1(n10689), .A2(n12027), .ZN(n7812) );
  INV_X1 U10183 ( .A(SI_20_), .ZN(n10690) );
  OR2_X1 U10184 ( .A1(n12033), .A2(n10690), .ZN(n7811) );
  NAND2_X1 U10185 ( .A1(n10734), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7819) );
  NAND2_X1 U10186 ( .A1(n7980), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7818) );
  NOR2_X1 U10187 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  OR2_X1 U10188 ( .A1(n7824), .A2(n7815), .ZN(n12525) );
  NAND2_X1 U10189 ( .A1(n6547), .A2(n12525), .ZN(n7817) );
  NAND2_X1 U10190 ( .A1(n10733), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7816) );
  NAND4_X1 U10191 ( .A1(n7819), .A2(n7818), .A3(n7817), .A4(n7816), .ZN(n12536) );
  NAND2_X1 U10192 ( .A1(n11980), .A2(n12536), .ZN(n12176) );
  INV_X1 U10193 ( .A(n12536), .ZN(n11940) );
  NAND2_X1 U10194 ( .A1(n12736), .A2(n11940), .ZN(n12175) );
  NAND2_X1 U10195 ( .A1(n12176), .A2(n12175), .ZN(n12171) );
  XNOR2_X1 U10196 ( .A(n7821), .B(n7820), .ZN(n10763) );
  NAND2_X1 U10197 ( .A1(n10763), .A2(n12027), .ZN(n7823) );
  INV_X1 U10198 ( .A(SI_21_), .ZN(n10764) );
  OR2_X1 U10199 ( .A1(n12033), .A2(n10764), .ZN(n7822) );
  OR2_X1 U10200 ( .A1(n7824), .A2(n11939), .ZN(n7825) );
  NAND2_X1 U10201 ( .A1(n7836), .A2(n7825), .ZN(n11938) );
  NAND2_X1 U10202 ( .A1(n6547), .A2(n11938), .ZN(n7830) );
  NAND2_X1 U10203 ( .A1(n7980), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7829) );
  INV_X1 U10204 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12731) );
  OR2_X1 U10205 ( .A1(n7558), .A2(n12731), .ZN(n7828) );
  INV_X1 U10206 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12512) );
  OR2_X1 U10207 ( .A1(n7826), .A2(n12512), .ZN(n7827) );
  NAND2_X1 U10208 ( .A1(n12514), .A2(n12522), .ZN(n12181) );
  NAND2_X1 U10209 ( .A1(n12515), .A2(n12181), .ZN(n7831) );
  OR2_X1 U10210 ( .A1(n12514), .A2(n12522), .ZN(n12182) );
  NAND2_X1 U10211 ( .A1(n7831), .A2(n12182), .ZN(n12495) );
  XNOR2_X1 U10212 ( .A(n7833), .B(n7832), .ZN(n10967) );
  NAND2_X1 U10213 ( .A1(n10967), .A2(n12027), .ZN(n7835) );
  INV_X1 U10214 ( .A(SI_22_), .ZN(n13626) );
  NAND2_X1 U10215 ( .A1(n10733), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7841) );
  NAND2_X1 U10216 ( .A1(n10734), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10217 ( .A1(n7836), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U10218 ( .A1(n7847), .A2(n7837), .ZN(n12502) );
  NAND2_X1 U10219 ( .A1(n6547), .A2(n12502), .ZN(n7839) );
  NAND2_X1 U10220 ( .A1(n7980), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7838) );
  NAND4_X1 U10221 ( .A1(n7841), .A2(n7840), .A3(n7839), .A4(n7838), .ZN(n12509) );
  INV_X1 U10222 ( .A(n12509), .ZN(n11843) );
  NAND2_X1 U10223 ( .A1(n12501), .A2(n11843), .ZN(n12191) );
  NAND2_X1 U10224 ( .A1(n12495), .A2(n12191), .ZN(n7842) );
  OR2_X1 U10225 ( .A1(n12501), .A2(n11843), .ZN(n12187) );
  XNOR2_X1 U10226 ( .A(n7844), .B(n7843), .ZN(n11188) );
  NAND2_X1 U10227 ( .A1(n11188), .A2(n12027), .ZN(n7846) );
  OR2_X1 U10228 ( .A1(n12033), .A2(n11190), .ZN(n7845) );
  NAND2_X1 U10229 ( .A1(n7847), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U10230 ( .A1(n7849), .A2(n7848), .ZN(n12487) );
  NAND2_X1 U10231 ( .A1(n12487), .A2(n6551), .ZN(n7853) );
  NAND2_X1 U10232 ( .A1(n10733), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7852) );
  NAND2_X1 U10233 ( .A1(n10734), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7851) );
  NAND2_X1 U10234 ( .A1(n7980), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7850) );
  NAND4_X1 U10235 ( .A1(n7853), .A2(n7852), .A3(n7851), .A4(n7850), .ZN(n12249) );
  NAND2_X1 U10236 ( .A1(n11844), .A2(n12249), .ZN(n12068) );
  NAND2_X1 U10237 ( .A1(n12724), .A2(n12500), .ZN(n12188) );
  NAND2_X1 U10238 ( .A1(n12492), .A2(n12480), .ZN(n7854) );
  NAND2_X1 U10239 ( .A1(n12721), .A2(n12484), .ZN(n12069) );
  NAND2_X1 U10240 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7855), .ZN(n7857) );
  INV_X1 U10241 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13394) );
  INV_X1 U10242 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14456) );
  AOI22_X1 U10243 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13394), .B2(n14456), .ZN(n7867) );
  XNOR2_X1 U10244 ( .A(n7866), .B(n7867), .ZN(n11677) );
  NAND2_X1 U10245 ( .A1(n11677), .A2(n12027), .ZN(n7859) );
  INV_X1 U10246 ( .A(SI_25_), .ZN(n11680) );
  OR2_X1 U10247 ( .A1(n12033), .A2(n11680), .ZN(n7858) );
  INV_X1 U10248 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n7860) );
  NAND2_X1 U10249 ( .A1(n7861), .A2(n7860), .ZN(n7871) );
  OR2_X1 U10250 ( .A1(n7861), .A2(n7860), .ZN(n7862) );
  NAND2_X1 U10251 ( .A1(n7871), .A2(n7862), .ZN(n12455) );
  NAND2_X1 U10252 ( .A1(n12455), .A2(n6547), .ZN(n7865) );
  AOI22_X1 U10253 ( .A1(n10733), .A2(P3_REG0_REG_25__SCAN_IN), .B1(n10734), 
        .B2(P3_REG2_REG_25__SCAN_IN), .ZN(n7864) );
  NAND2_X1 U10254 ( .A1(n7980), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n7863) );
  OR2_X1 U10255 ( .A1(n12717), .A2(n12468), .ZN(n12067) );
  NAND2_X1 U10256 ( .A1(n12717), .A2(n12468), .ZN(n12066) );
  INV_X1 U10257 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13388) );
  INV_X1 U10258 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U10259 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n13388), .B2(n11816), .ZN(n7868) );
  XNOR2_X1 U10260 ( .A(n7879), .B(n7868), .ZN(n12777) );
  NAND2_X1 U10261 ( .A1(n12777), .A2(n12027), .ZN(n7870) );
  INV_X1 U10262 ( .A(SI_26_), .ZN(n13476) );
  OR2_X1 U10263 ( .A1(n12033), .A2(n13476), .ZN(n7869) );
  NAND2_X1 U10264 ( .A1(n7871), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n7872) );
  NAND2_X1 U10265 ( .A1(n7885), .A2(n7872), .ZN(n12439) );
  NAND2_X1 U10266 ( .A1(n12439), .A2(n6551), .ZN(n7877) );
  INV_X1 U10267 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12713) );
  NAND2_X1 U10268 ( .A1(n7980), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7874) );
  NAND2_X1 U10269 ( .A1(n10734), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7873) );
  OAI211_X1 U10270 ( .C1(n7558), .C2(n12713), .A(n7874), .B(n7873), .ZN(n7875)
         );
  INV_X1 U10271 ( .A(n7875), .ZN(n7876) );
  NAND2_X1 U10272 ( .A1(n12433), .A2(n12198), .ZN(n7878) );
  NAND2_X1 U10273 ( .A1(n12438), .A2(n12416), .ZN(n12197) );
  NAND2_X1 U10274 ( .A1(n7878), .A2(n12197), .ZN(n12412) );
  NOR2_X1 U10275 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13388), .ZN(n7880) );
  OAI22_X1 U10276 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n11816), .B1(n7880), 
        .B2(n7879), .ZN(n7893) );
  INV_X1 U10277 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13386) );
  AOI22_X1 U10278 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13386), .B2(n7091), .ZN(n7881) );
  INV_X1 U10279 ( .A(n7881), .ZN(n7882) );
  XNOR2_X1 U10280 ( .A(n7893), .B(n7882), .ZN(n12773) );
  NAND2_X1 U10281 ( .A1(n12773), .A2(n12027), .ZN(n7884) );
  INV_X1 U10282 ( .A(SI_27_), .ZN(n12775) );
  INV_X1 U10283 ( .A(n7899), .ZN(n7887) );
  NAND2_X1 U10284 ( .A1(n7885), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n7886) );
  NAND2_X1 U10285 ( .A1(n7887), .A2(n7886), .ZN(n12422) );
  NAND2_X1 U10286 ( .A1(n12422), .A2(n6547), .ZN(n7892) );
  NAND2_X1 U10287 ( .A1(n10733), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10288 ( .A1(n10734), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7889) );
  NAND2_X1 U10289 ( .A1(n7980), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7888) );
  AND3_X1 U10290 ( .A1(n7890), .A2(n7889), .A3(n7888), .ZN(n7891) );
  XNOR2_X1 U10291 ( .A(n12202), .B(n12434), .ZN(n12413) );
  INV_X1 U10292 ( .A(n12434), .ZN(n11906) );
  AND2_X1 U10293 ( .A1(n12202), .A2(n11906), .ZN(n12207) );
  NOR2_X1 U10294 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7091), .ZN(n7894) );
  INV_X1 U10295 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13383) );
  AOI22_X1 U10296 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13383), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11814), .ZN(n7895) );
  INV_X1 U10297 ( .A(n7895), .ZN(n7896) );
  XNOR2_X1 U10298 ( .A(n8808), .B(n7896), .ZN(n11817) );
  NAND2_X1 U10299 ( .A1(n11817), .A2(n12027), .ZN(n7898) );
  INV_X1 U10300 ( .A(SI_28_), .ZN(n11820) );
  OR2_X1 U10301 ( .A1(n12033), .A2(n11820), .ZN(n7897) );
  INV_X1 U10302 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n11905) );
  NOR2_X1 U10303 ( .A1(n7899), .A2(n11905), .ZN(n7900) );
  INV_X1 U10304 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n8035) );
  NAND2_X1 U10305 ( .A1(n7980), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10306 ( .A1(n10734), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7901) );
  OAI211_X1 U10307 ( .C1(n7558), .C2(n8035), .A(n7902), .B(n7901), .ZN(n7903)
         );
  OR2_X1 U10308 ( .A1(n12407), .A2(n12417), .ZN(n12208) );
  NAND2_X1 U10309 ( .A1(n12407), .A2(n12417), .ZN(n12209) );
  NAND2_X1 U10310 ( .A1(n12208), .A2(n12209), .ZN(n12205) );
  XNOR2_X1 U10311 ( .A(n8813), .B(n12205), .ZN(n12408) );
  NAND2_X1 U10312 ( .A1(n6566), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7904) );
  MUX2_X1 U10313 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7904), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n7905) );
  INV_X1 U10314 ( .A(n6883), .ZN(n7906) );
  NAND2_X1 U10315 ( .A1(n7906), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7907) );
  MUX2_X1 U10316 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7907), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n7909) );
  NAND2_X1 U10317 ( .A1(n7909), .A2(n7908), .ZN(n10692) );
  OAI21_X1 U10318 ( .B1(n10965), .B2(n10816), .A(n12375), .ZN(n7912) );
  NAND2_X1 U10319 ( .A1(n7908), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10320 ( .A1(n7912), .A2(n10817), .ZN(n7914) );
  OAI21_X1 U10321 ( .B1(n10816), .B2(n12074), .A(n10965), .ZN(n7913) );
  NAND2_X1 U10322 ( .A1(n7914), .A2(n7913), .ZN(n10516) );
  NAND2_X1 U10323 ( .A1(n10692), .A2(n12391), .ZN(n10815) );
  INV_X1 U10324 ( .A(n10815), .ZN(n12234) );
  AND2_X1 U10325 ( .A1(n15406), .A2(n12234), .ZN(n7915) );
  NAND2_X1 U10326 ( .A1(n10516), .A2(n7915), .ZN(n7917) );
  NAND2_X1 U10327 ( .A1(n10816), .A2(n12391), .ZN(n7916) );
  NAND2_X1 U10328 ( .A1(n12408), .A2(n14640), .ZN(n7990) );
  NAND2_X1 U10329 ( .A1(n15320), .A2(n11411), .ZN(n7925) );
  INV_X1 U10330 ( .A(n7925), .ZN(n7918) );
  NOR2_X1 U10331 ( .A1(n7918), .A2(n11406), .ZN(n7927) );
  NAND2_X1 U10332 ( .A1(n12081), .A2(n12078), .ZN(n12702) );
  NAND2_X1 U10333 ( .A1(n12696), .A2(n10511), .ZN(n12695) );
  NAND2_X1 U10334 ( .A1(n12702), .A2(n12695), .ZN(n15346) );
  NAND2_X1 U10335 ( .A1(n15341), .A2(n10830), .ZN(n15344) );
  NAND2_X1 U10336 ( .A1(n12698), .A2(n15354), .ZN(n7921) );
  AND2_X1 U10337 ( .A1(n15344), .A2(n7921), .ZN(n7920) );
  NAND2_X1 U10338 ( .A1(n15346), .A2(n7920), .ZN(n7924) );
  INV_X1 U10339 ( .A(n7921), .ZN(n7922) );
  NAND2_X1 U10340 ( .A1(n12258), .A2(n11037), .ZN(n11405) );
  AND2_X1 U10341 ( .A1(n11405), .A2(n7925), .ZN(n7926) );
  OR2_X1 U10342 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  NAND2_X1 U10343 ( .A1(n12256), .A2(n11568), .ZN(n7930) );
  NAND2_X1 U10344 ( .A1(n11240), .A2(n7930), .ZN(n7934) );
  INV_X1 U10345 ( .A(n7930), .ZN(n11461) );
  NOR2_X1 U10346 ( .A1(n12257), .A2(n11386), .ZN(n11458) );
  NAND2_X1 U10347 ( .A1(n11458), .A2(n7930), .ZN(n7931) );
  OAI211_X1 U10348 ( .C1(n11547), .C2(n11461), .A(n11564), .B(n7931), .ZN(
        n7932) );
  INV_X1 U10349 ( .A(n7932), .ZN(n7933) );
  NAND2_X1 U10350 ( .A1(n12255), .A2(n7935), .ZN(n7936) );
  AND2_X1 U10351 ( .A1(n12254), .A2(n11565), .ZN(n7939) );
  NAND2_X1 U10352 ( .A1(n11671), .A2(n11750), .ZN(n7938) );
  NAND2_X1 U10353 ( .A1(n15303), .A2(n12120), .ZN(n12121) );
  OAI21_X1 U10354 ( .B1(n15303), .B2(n12120), .A(n12121), .ZN(n12118) );
  OR2_X2 U10355 ( .A1(n11485), .A2(n12118), .ZN(n11487) );
  NAND2_X1 U10356 ( .A1(n12127), .A2(n12134), .ZN(n15306) );
  NAND2_X1 U10357 ( .A1(n15307), .A2(n15306), .ZN(n15305) );
  NAND2_X1 U10358 ( .A1(n12253), .A2(n11634), .ZN(n7940) );
  NAND2_X1 U10359 ( .A1(n11791), .A2(n11731), .ZN(n7941) );
  NAND2_X1 U10360 ( .A1(n11725), .A2(n7941), .ZN(n11760) );
  NAND2_X1 U10361 ( .A1(n15304), .A2(n11717), .ZN(n11759) );
  NAND2_X1 U10362 ( .A1(n12252), .A2(n11793), .ZN(n7942) );
  AND2_X1 U10363 ( .A1(n11759), .A2(n7942), .ZN(n7944) );
  INV_X1 U10364 ( .A(n7942), .ZN(n7943) );
  NAND2_X1 U10365 ( .A1(n12138), .A2(n12130), .ZN(n11761) );
  AOI21_X2 U10366 ( .B1(n11760), .B2(n7944), .A(n7443), .ZN(n11771) );
  AND2_X1 U10367 ( .A1(n12618), .A2(n11994), .ZN(n7945) );
  INV_X1 U10368 ( .A(n12618), .ZN(n11810) );
  NAND2_X1 U10369 ( .A1(n11810), .A2(n14629), .ZN(n7946) );
  NAND2_X2 U10370 ( .A1(n7439), .A2(n7948), .ZN(n12616) );
  NAND2_X1 U10371 ( .A1(n11800), .A2(n11982), .ZN(n12602) );
  NAND2_X1 U10372 ( .A1(n12608), .A2(n12617), .ZN(n7949) );
  AND2_X1 U10373 ( .A1(n12602), .A2(n7949), .ZN(n7950) );
  AOI21_X2 U10374 ( .B1(n12616), .B2(n7950), .A(n6660), .ZN(n12578) );
  NAND2_X1 U10375 ( .A1(n12578), .A2(n7951), .ZN(n7953) );
  NAND2_X1 U10376 ( .A1(n11955), .A2(n12251), .ZN(n7952) );
  NAND2_X1 U10377 ( .A1(n7953), .A2(n7952), .ZN(n12570) );
  NAND2_X1 U10378 ( .A1(n12570), .A2(n12569), .ZN(n7956) );
  NAND2_X1 U10379 ( .A1(n7954), .A2(n12580), .ZN(n7955) );
  NAND2_X1 U10380 ( .A1(n7956), .A2(n7955), .ZN(n12551) );
  INV_X1 U10381 ( .A(n12551), .ZN(n7958) );
  NAND2_X1 U10382 ( .A1(n12745), .A2(n12572), .ZN(n7960) );
  NAND2_X1 U10383 ( .A1(n12549), .A2(n7960), .ZN(n12533) );
  INV_X1 U10384 ( .A(n11933), .ZN(n12740) );
  NAND2_X1 U10385 ( .A1(n12740), .A2(n12520), .ZN(n7963) );
  AND2_X1 U10386 ( .A1(n12736), .A2(n12536), .ZN(n7964) );
  AOI21_X2 U10387 ( .B1(n12519), .B2(n12171), .A(n7964), .ZN(n12508) );
  NAND2_X1 U10388 ( .A1(n12182), .A2(n12181), .ZN(n12516) );
  NAND2_X1 U10389 ( .A1(n12501), .A2(n12509), .ZN(n12461) );
  OR2_X1 U10390 ( .A1(n12480), .A2(n12461), .ZN(n7970) );
  AND2_X1 U10391 ( .A1(n12516), .A2(n7970), .ZN(n7967) );
  NAND2_X1 U10392 ( .A1(n12724), .A2(n12249), .ZN(n12464) );
  INV_X1 U10393 ( .A(n7975), .ZN(n7966) );
  AND2_X1 U10394 ( .A1(n7967), .A2(n7966), .ZN(n12427) );
  NAND2_X1 U10395 ( .A1(n12717), .A2(n12470), .ZN(n12429) );
  NAND2_X1 U10396 ( .A1(n12438), .A2(n12448), .ZN(n7968) );
  AND2_X1 U10397 ( .A1(n12429), .A2(n7968), .ZN(n7969) );
  AND2_X1 U10398 ( .A1(n12427), .A2(n7969), .ZN(n7978) );
  INV_X1 U10399 ( .A(n7969), .ZN(n7977) );
  INV_X1 U10400 ( .A(n7970), .ZN(n7973) );
  NAND2_X1 U10401 ( .A1(n12733), .A2(n12522), .ZN(n12496) );
  OR2_X1 U10402 ( .A1(n12501), .A2(n12509), .ZN(n7971) );
  AND2_X1 U10403 ( .A1(n12496), .A2(n7971), .ZN(n12460) );
  INV_X1 U10404 ( .A(n12480), .ZN(n12491) );
  AND2_X1 U10405 ( .A1(n12460), .A2(n12491), .ZN(n7972) );
  OR2_X1 U10406 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  OR2_X1 U10407 ( .A1(n7975), .A2(n7974), .ZN(n12466) );
  NAND2_X1 U10408 ( .A1(n12721), .A2(n11922), .ZN(n7976) );
  AND2_X1 U10409 ( .A1(n12466), .A2(n7976), .ZN(n12444) );
  INV_X1 U10410 ( .A(n12451), .ZN(n12446) );
  AND2_X1 U10411 ( .A1(n12444), .A2(n12446), .ZN(n12428) );
  OR2_X1 U10412 ( .A1(n10965), .A2(n12391), .ZN(n8021) );
  NAND2_X1 U10413 ( .A1(n12074), .A2(n10816), .ZN(n12020) );
  OAI211_X1 U10414 ( .C1(n7979), .C2(n12205), .A(n8814), .B(n15323), .ZN(n7989) );
  NAND2_X1 U10415 ( .A1(n14614), .A2(n6551), .ZN(n10739) );
  INV_X1 U10416 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n13480) );
  NAND2_X1 U10417 ( .A1(n10733), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10418 ( .A1(n10734), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n7981) );
  OAI211_X1 U10419 ( .C1(n13480), .C2(n7604), .A(n7982), .B(n7981), .ZN(n7983)
         );
  INV_X1 U10420 ( .A(n7983), .ZN(n7984) );
  INV_X1 U10421 ( .A(n8812), .ZN(n12248) );
  NAND2_X1 U10422 ( .A1(n10580), .A2(n10577), .ZN(n7987) );
  AOI22_X1 U10423 ( .A1(n12248), .A2(n15319), .B1(n15321), .B2(n12434), .ZN(
        n7988) );
  NAND2_X1 U10424 ( .A1(n7990), .A2(n12411), .ZN(n12627) );
  INV_X1 U10425 ( .A(n12627), .ZN(n8039) );
  INV_X1 U10426 ( .A(n7991), .ZN(n7997) );
  NOR2_X1 U10427 ( .A1(n7992), .A2(n8002), .ZN(n7995) );
  NAND2_X1 U10428 ( .A1(n6543), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7998) );
  MUX2_X1 U10429 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7998), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n8000) );
  INV_X1 U10430 ( .A(n7992), .ZN(n7999) );
  XNOR2_X1 U10431 ( .A(n11559), .B(P3_B_REG_SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10432 ( .A1(n11678), .A2(n8001), .ZN(n8003) );
  INV_X1 U10433 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U10434 ( .A1(n8008), .A2(n8004), .ZN(n8006) );
  NAND2_X1 U10435 ( .A1(n12780), .A2(n11678), .ZN(n8005) );
  INV_X1 U10436 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n8007) );
  NAND2_X1 U10437 ( .A1(n8008), .A2(n8007), .ZN(n8010) );
  NAND2_X1 U10438 ( .A1(n12780), .A2(n11559), .ZN(n8009) );
  NAND2_X1 U10439 ( .A1(n10744), .A2(n10814), .ZN(n8829) );
  NOR2_X1 U10440 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_12__SCAN_IN), .ZN(
        n8014) );
  NOR4_X1 U10441 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8013) );
  NOR4_X1 U10442 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8012) );
  NOR4_X1 U10443 ( .A1(P3_D_REG_25__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8011) );
  NAND4_X1 U10444 ( .A1(n8014), .A2(n8013), .A3(n8012), .A4(n8011), .ZN(n8020)
         );
  NOR4_X1 U10445 ( .A1(P3_D_REG_21__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8018) );
  NOR4_X1 U10446 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8017) );
  NOR4_X1 U10447 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8016) );
  NOR4_X1 U10448 ( .A1(P3_D_REG_16__SCAN_IN), .A2(P3_D_REG_30__SCAN_IN), .A3(
        P3_D_REG_13__SCAN_IN), .A4(P3_D_REG_23__SCAN_IN), .ZN(n8015) );
  NAND4_X1 U10449 ( .A1(n8018), .A2(n8017), .A3(n8016), .A4(n8015), .ZN(n8019)
         );
  OAI21_X1 U10450 ( .B1(n8020), .B2(n8019), .A(n8008), .ZN(n8826) );
  INV_X1 U10451 ( .A(n8826), .ZN(n8024) );
  INV_X1 U10452 ( .A(n8021), .ZN(n8022) );
  AND2_X1 U10453 ( .A1(n10816), .A2(n10817), .ZN(n12063) );
  NAND2_X1 U10454 ( .A1(n8022), .A2(n12063), .ZN(n10512) );
  INV_X1 U10455 ( .A(n10814), .ZN(n8023) );
  NAND2_X1 U10456 ( .A1(n8832), .A2(n8023), .ZN(n8827) );
  INV_X1 U10457 ( .A(n10516), .ZN(n8025) );
  OAI22_X1 U10458 ( .A1(n10517), .A2(n10512), .B1(n10826), .B2(n8025), .ZN(
        n8031) );
  INV_X1 U10459 ( .A(n11678), .ZN(n8028) );
  INV_X1 U10460 ( .A(n11559), .ZN(n8027) );
  NAND2_X1 U10461 ( .A1(n6557), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8030) );
  NAND2_X1 U10462 ( .A1(n8031), .A2(n10574), .ZN(n8034) );
  INV_X1 U10463 ( .A(n10517), .ZN(n8032) );
  NAND2_X1 U10464 ( .A1(n10574), .A2(n12234), .ZN(n10827) );
  NOR2_X1 U10465 ( .A1(n10827), .A2(n12219), .ZN(n10521) );
  NAND2_X1 U10466 ( .A1(n8032), .A2(n10521), .ZN(n8033) );
  NAND2_X1 U10467 ( .A1(n15412), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8036) );
  INV_X1 U10468 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9989) );
  AND2_X1 U10469 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8040) );
  NAND2_X1 U10470 ( .A1(n9960), .A2(n8040), .ZN(n9007) );
  OAI21_X1 U10471 ( .B1(n8187), .B2(n8186), .A(n9007), .ZN(n8171) );
  NOR2_X1 U10472 ( .A1(n8041), .A2(n9963), .ZN(n8042) );
  INV_X1 U10473 ( .A(n8201), .ZN(n8044) );
  INV_X1 U10474 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9962) );
  MUX2_X1 U10475 ( .A(n9962), .B(n9998), .S(n8043), .Z(n8045) );
  XNOR2_X1 U10476 ( .A(n8045), .B(SI_2_), .ZN(n8202) );
  NAND2_X1 U10477 ( .A1(n8044), .A2(n8202), .ZN(n8048) );
  INV_X1 U10478 ( .A(n8045), .ZN(n8046) );
  NAND2_X1 U10479 ( .A1(n8046), .A2(SI_2_), .ZN(n8047) );
  NAND2_X1 U10480 ( .A1(n8225), .A2(n8050), .ZN(n8053) );
  NAND2_X1 U10481 ( .A1(n8051), .A2(SI_3_), .ZN(n8052) );
  NAND2_X1 U10482 ( .A1(n8053), .A2(n8052), .ZN(n8247) );
  XNOR2_X1 U10483 ( .A(n8055), .B(SI_4_), .ZN(n8248) );
  INV_X1 U10484 ( .A(n8248), .ZN(n8054) );
  NAND2_X1 U10485 ( .A1(n8247), .A2(n8054), .ZN(n8057) );
  NAND2_X1 U10486 ( .A1(n8055), .A2(SI_4_), .ZN(n8056) );
  NAND2_X1 U10487 ( .A1(n8060), .A2(SI_6_), .ZN(n8061) );
  MUX2_X1 U10488 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9367), .Z(n8063) );
  XNOR2_X1 U10489 ( .A(n8063), .B(SI_7_), .ZN(n8312) );
  INV_X1 U10490 ( .A(n8312), .ZN(n8062) );
  NAND2_X1 U10491 ( .A1(n8063), .A2(SI_7_), .ZN(n8064) );
  MUX2_X1 U10492 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9367), .Z(n8067) );
  XNOR2_X1 U10493 ( .A(n8067), .B(SI_8_), .ZN(n8330) );
  INV_X1 U10494 ( .A(n8330), .ZN(n8066) );
  NAND2_X1 U10495 ( .A1(n8067), .A2(SI_8_), .ZN(n8068) );
  MUX2_X1 U10496 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9367), .Z(n8070) );
  XNOR2_X1 U10497 ( .A(n8070), .B(SI_9_), .ZN(n8346) );
  INV_X1 U10498 ( .A(n8346), .ZN(n8069) );
  MUX2_X1 U10499 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9367), .Z(n8366) );
  INV_X1 U10500 ( .A(n8366), .ZN(n8072) );
  INV_X1 U10501 ( .A(SI_10_), .ZN(n8071) );
  NAND2_X1 U10502 ( .A1(n8072), .A2(n8071), .ZN(n8073) );
  NAND2_X1 U10503 ( .A1(n8365), .A2(n8073), .ZN(n8075) );
  NAND2_X1 U10504 ( .A1(n8366), .A2(SI_10_), .ZN(n8074) );
  NAND2_X1 U10505 ( .A1(n8075), .A2(n8074), .ZN(n8384) );
  MUX2_X1 U10506 ( .A(n10051), .B(n10053), .S(n9367), .Z(n8077) );
  INV_X1 U10507 ( .A(SI_11_), .ZN(n8076) );
  NAND2_X1 U10508 ( .A1(n8077), .A2(n8076), .ZN(n8080) );
  INV_X1 U10509 ( .A(n8077), .ZN(n8078) );
  NAND2_X1 U10510 ( .A1(n8078), .A2(SI_11_), .ZN(n8079) );
  NAND2_X1 U10511 ( .A1(n8080), .A2(n8079), .ZN(n8385) );
  MUX2_X1 U10512 ( .A(n10175), .B(n10174), .S(n9367), .Z(n8081) );
  NAND2_X1 U10513 ( .A1(n8081), .A2(n14575), .ZN(n8084) );
  INV_X1 U10514 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U10515 ( .A1(n8082), .A2(SI_12_), .ZN(n8083) );
  MUX2_X1 U10516 ( .A(n13631), .B(n10252), .S(n9367), .Z(n8085) );
  NAND2_X1 U10517 ( .A1(n8085), .A2(n10029), .ZN(n8088) );
  INV_X1 U10518 ( .A(n8085), .ZN(n8086) );
  NAND2_X1 U10519 ( .A1(n8086), .A2(SI_13_), .ZN(n8087) );
  MUX2_X1 U10520 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n8043), .Z(n8467) );
  NOR2_X1 U10521 ( .A1(n8467), .A2(SI_14_), .ZN(n8096) );
  MUX2_X1 U10522 ( .A(n10443), .B(n13634), .S(n8043), .Z(n8091) );
  NAND2_X1 U10523 ( .A1(n8091), .A2(n8090), .ZN(n8097) );
  INV_X1 U10524 ( .A(n8091), .ZN(n8092) );
  NAND2_X1 U10525 ( .A1(n8092), .A2(SI_15_), .ZN(n8093) );
  NAND2_X1 U10526 ( .A1(n8097), .A2(n8093), .ZN(n8469) );
  INV_X1 U10527 ( .A(n8467), .ZN(n8094) );
  NOR2_X1 U10528 ( .A1(n8094), .A2(n10120), .ZN(n8095) );
  MUX2_X1 U10529 ( .A(n7472), .B(n10369), .S(n9981), .Z(n8099) );
  NAND2_X1 U10530 ( .A1(n8099), .A2(n8098), .ZN(n8102) );
  INV_X1 U10531 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10532 ( .A1(n8100), .A2(SI_16_), .ZN(n8101) );
  MUX2_X1 U10533 ( .A(n13502), .B(n10422), .S(n9981), .Z(n8505) );
  MUX2_X1 U10534 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9981), .Z(n8529) );
  MUX2_X1 U10535 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9981), .Z(n8554) );
  AOI22_X1 U10536 ( .A1(SI_18_), .A2(n8529), .B1(n8554), .B2(SI_19_), .ZN(
        n8103) );
  OAI21_X1 U10537 ( .B1(n8529), .B2(SI_18_), .A(SI_19_), .ZN(n8106) );
  INV_X1 U10538 ( .A(n8554), .ZN(n8105) );
  NOR2_X1 U10539 ( .A1(SI_18_), .A2(SI_19_), .ZN(n8104) );
  INV_X1 U10540 ( .A(n8529), .ZN(n8531) );
  AOI22_X1 U10541 ( .A1(n8106), .A2(n8105), .B1(n8104), .B2(n8531), .ZN(n8107)
         );
  NAND2_X1 U10542 ( .A1(n8108), .A2(n10690), .ZN(n8109) );
  MUX2_X1 U10543 ( .A(n10682), .B(n10681), .S(n9981), .Z(n8574) );
  MUX2_X1 U10544 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9981), .Z(n8112) );
  NAND2_X1 U10545 ( .A1(n8112), .A2(SI_21_), .ZN(n8114) );
  OAI21_X1 U10546 ( .B1(SI_21_), .B2(n8112), .A(n8114), .ZN(n8113) );
  INV_X1 U10547 ( .A(n8113), .ZN(n8593) );
  NAND2_X1 U10548 ( .A1(n8594), .A2(n8593), .ZN(n8596) );
  NAND2_X1 U10549 ( .A1(n8596), .A2(n8114), .ZN(n8116) );
  INV_X1 U10550 ( .A(n8116), .ZN(n8115) );
  MUX2_X1 U10551 ( .A(n8117), .B(n11056), .S(n9981), .Z(n8614) );
  MUX2_X1 U10552 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9981), .Z(n8121) );
  INV_X1 U10553 ( .A(n8125), .ZN(n8124) );
  NAND2_X1 U10554 ( .A1(n8124), .A2(n11558), .ZN(n8126) );
  MUX2_X1 U10555 ( .A(n11741), .B(n11739), .S(n9981), .Z(n8650) );
  MUX2_X1 U10556 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9981), .Z(n8129) );
  XNOR2_X1 U10557 ( .A(n8129), .B(SI_25_), .ZN(n8671) );
  OAI22_X2 U10558 ( .A1(n8672), .A2(n8671), .B1(SI_25_), .B2(n8129), .ZN(n8690) );
  MUX2_X1 U10559 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9981), .Z(n8130) );
  NAND2_X1 U10560 ( .A1(n8130), .A2(SI_26_), .ZN(n8131) );
  OAI21_X1 U10561 ( .B1(SI_26_), .B2(n8130), .A(n8131), .ZN(n8689) );
  MUX2_X1 U10562 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9981), .Z(n8713) );
  NOR2_X1 U10563 ( .A1(n8132), .A2(n12775), .ZN(n8134) );
  NAND2_X1 U10564 ( .A1(n8132), .A2(n12775), .ZN(n8133) );
  MUX2_X1 U10565 ( .A(n11814), .B(n13383), .S(n9981), .Z(n8882) );
  XNOR2_X1 U10566 ( .A(n8882), .B(SI_28_), .ZN(n8880) );
  XNOR2_X2 U10567 ( .A(n8881), .B(n8880), .ZN(n9458) );
  INV_X1 U10568 ( .A(n8146), .ZN(n8150) );
  NOR2_X1 U10569 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), 
        .ZN(n8137) );
  NAND4_X1 U10570 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8488), .ZN(n8508)
         );
  NAND3_X1 U10571 ( .A1(n8347), .A2(n8139), .A3(n8138), .ZN(n8140) );
  NOR2_X1 U10572 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8144) );
  NAND4_X1 U10573 ( .A1(n8144), .A2(n8143), .A3(n6687), .A4(n8142), .ZN(n8145)
         );
  NAND2_X1 U10574 ( .A1(n9458), .A2(n9780), .ZN(n8152) );
  NAND2_X1 U10575 ( .A1(n8694), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10576 ( .A1(n8164), .A2(n8165), .ZN(n8160) );
  INV_X1 U10577 ( .A(n8160), .ZN(n8153) );
  NAND2_X1 U10578 ( .A1(n8153), .A2(n8142), .ZN(n8163) );
  NAND2_X1 U10579 ( .A1(n8163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8155) );
  INV_X1 U10580 ( .A(n8156), .ZN(n8778) );
  NAND2_X2 U10581 ( .A1(n8159), .A2(n8158), .ZN(n11057) );
  NAND2_X1 U10582 ( .A1(n8160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8161) );
  XNOR2_X1 U10583 ( .A(n11057), .B(n9593), .ZN(n8169) );
  NAND2_X1 U10584 ( .A1(n8167), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8168) );
  NAND2_X1 U10585 ( .A1(n8169), .A2(n13047), .ZN(n8888) );
  XNOR2_X1 U10586 ( .A(n8170), .B(n8171), .ZN(n9990) );
  INV_X1 U10587 ( .A(n8188), .ZN(n8172) );
  NAND2_X1 U10588 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8173) );
  MUX2_X1 U10589 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8173), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8176) );
  INV_X1 U10590 ( .A(n8203), .ZN(n8175) );
  NAND2_X1 U10591 ( .A1(n8176), .A2(n8175), .ZN(n14947) );
  INV_X1 U10592 ( .A(n14947), .ZN(n10060) );
  INV_X1 U10593 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10349) );
  OR2_X1 U10594 ( .A1(n8212), .A2(n10349), .ZN(n8184) );
  INV_X1 U10595 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8180) );
  OR2_X1 U10596 ( .A1(n8213), .A2(n8180), .ZN(n8183) );
  INV_X1 U10597 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n10354) );
  OR2_X1 U10598 ( .A1(n8234), .A2(n10354), .ZN(n8182) );
  NAND2_X1 U10599 ( .A1(n8233), .A2(n12988), .ZN(n8198) );
  XNOR2_X1 U10600 ( .A(n8197), .B(n8198), .ZN(n11861) );
  XNOR2_X1 U10601 ( .A(n8187), .B(n8186), .ZN(n13397) );
  INV_X1 U10602 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13396) );
  MUX2_X2 U10603 ( .A(n13397), .B(n13396), .S(n8188), .Z(n15042) );
  NAND2_X1 U10604 ( .A1(n8211), .A2(n15042), .ZN(n8196) );
  INV_X1 U10605 ( .A(n15042), .ZN(n10167) );
  NAND2_X1 U10606 ( .A1(n15021), .A2(n10167), .ZN(n8195) );
  NAND2_X1 U10607 ( .A1(n8719), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8194) );
  INV_X1 U10608 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14950) );
  OR2_X1 U10609 ( .A1(n8234), .A2(n14950), .ZN(n8193) );
  INV_X1 U10610 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8189) );
  OR2_X1 U10611 ( .A1(n8213), .A2(n8189), .ZN(n8192) );
  INV_X1 U10612 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n8190) );
  NAND4_X1 U10613 ( .A1(n8194), .A2(n8193), .A3(n8192), .A4(n8191), .ZN(n9597)
         );
  OR2_X1 U10614 ( .A1(n9597), .A2(n15042), .ZN(n10302) );
  AND2_X1 U10615 ( .A1(n8195), .A2(n10302), .ZN(n10172) );
  NAND2_X1 U10616 ( .A1(n8196), .A2(n10172), .ZN(n11860) );
  NAND2_X1 U10617 ( .A1(n11861), .A2(n11860), .ZN(n11859) );
  INV_X1 U10618 ( .A(n8197), .ZN(n8199) );
  NAND2_X1 U10619 ( .A1(n8199), .A2(n8198), .ZN(n8200) );
  NAND2_X1 U10620 ( .A1(n11859), .A2(n8200), .ZN(n10194) );
  XNOR2_X1 U10621 ( .A(n8201), .B(n8202), .ZN(n9961) );
  NAND2_X1 U10622 ( .A1(n9961), .A2(n8226), .ZN(n8210) );
  NOR2_X1 U10623 ( .A1(n8203), .A2(n8333), .ZN(n8204) );
  MUX2_X1 U10624 ( .A(n8333), .B(n8204), .S(P2_IR_REG_2__SCAN_IN), .Z(n8206)
         );
  NAND2_X1 U10625 ( .A1(n8389), .A2(n10074), .ZN(n8207) );
  OAI21_X1 U10626 ( .B1(n8227), .B2(n9998), .A(n8207), .ZN(n8208) );
  INV_X1 U10627 ( .A(n8208), .ZN(n8209) );
  INV_X1 U10628 ( .A(n10756), .ZN(n10331) );
  NAND2_X1 U10629 ( .A1(n8719), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8217) );
  INV_X1 U10630 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10754) );
  OR2_X1 U10631 ( .A1(n8212), .A2(n10754), .ZN(n8216) );
  INV_X1 U10632 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10059) );
  OR2_X1 U10633 ( .A1(n8213), .A2(n10059), .ZN(n8215) );
  INV_X1 U10634 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10073) );
  OR2_X1 U10635 ( .A1(n8234), .A2(n10073), .ZN(n8214) );
  NAND2_X1 U10636 ( .A1(n8233), .A2(n12986), .ZN(n8219) );
  NAND2_X1 U10637 ( .A1(n8218), .A2(n8219), .ZN(n8223) );
  INV_X1 U10638 ( .A(n8218), .ZN(n8221) );
  INV_X1 U10639 ( .A(n8219), .ZN(n8220) );
  NAND2_X1 U10640 ( .A1(n8221), .A2(n8220), .ZN(n8222) );
  AND2_X1 U10641 ( .A1(n8223), .A2(n8222), .ZN(n10195) );
  NAND2_X1 U10642 ( .A1(n10194), .A2(n10195), .ZN(n10193) );
  NAND2_X1 U10643 ( .A1(n10193), .A2(n8223), .ZN(n10227) );
  INV_X1 U10644 ( .A(n10227), .ZN(n8241) );
  XNOR2_X1 U10645 ( .A(n8225), .B(n8224), .ZN(n9985) );
  NAND2_X1 U10646 ( .A1(n9985), .A2(n8226), .ZN(n8232) );
  MUX2_X1 U10647 ( .A(n8333), .B(n8228), .S(P2_IR_REG_3__SCAN_IN), .Z(n8230)
         );
  AOI22_X1 U10648 ( .A1(n8694), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n12992), 
        .B2(n8389), .ZN(n8231) );
  INV_X1 U10649 ( .A(n10433), .ZN(n8896) );
  XNOR2_X1 U10650 ( .A(n8718), .B(n8896), .ZN(n8242) );
  INV_X1 U10651 ( .A(n8233), .ZN(n8274) );
  NAND2_X1 U10652 ( .A1(n8658), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8239) );
  OR2_X1 U10653 ( .A1(n8414), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8238) );
  INV_X1 U10654 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10432) );
  OR2_X1 U10655 ( .A1(n8662), .A2(n10432), .ZN(n8237) );
  INV_X1 U10656 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8235) );
  OR2_X1 U10657 ( .A1(n8563), .A2(n8235), .ZN(n8236) );
  NAND2_X1 U10658 ( .A1(n8233), .A2(n12985), .ZN(n8243) );
  XNOR2_X1 U10659 ( .A(n8242), .B(n8243), .ZN(n10228) );
  INV_X1 U10660 ( .A(n10228), .ZN(n8240) );
  INV_X1 U10661 ( .A(n8242), .ZN(n8245) );
  INV_X1 U10662 ( .A(n8243), .ZN(n8244) );
  NAND2_X1 U10663 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  XNOR2_X1 U10664 ( .A(n8247), .B(n8248), .ZN(n9986) );
  NAND2_X1 U10665 ( .A1(n9986), .A2(n9780), .ZN(n8254) );
  INV_X1 U10666 ( .A(n8249), .ZN(n8251) );
  NAND2_X1 U10667 ( .A1(n8251), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8250) );
  MUX2_X1 U10668 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8250), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8252) );
  AOI22_X1 U10669 ( .A1(n8694), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n10076), 
        .B2(n8389), .ZN(n8253) );
  XNOR2_X1 U10670 ( .A(n8211), .B(n10417), .ZN(n8261) );
  INV_X2 U10671 ( .A(n8662), .ZN(n9769) );
  NAND2_X1 U10672 ( .A1(n9769), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8259) );
  INV_X1 U10673 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10066) );
  OR2_X1 U10674 ( .A1(n8956), .A2(n10066), .ZN(n8258) );
  NAND2_X1 U10675 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8277) );
  OAI21_X1 U10676 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8277), .ZN(n10527) );
  OR2_X1 U10677 ( .A1(n8414), .A2(n10527), .ZN(n8257) );
  INV_X1 U10678 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8255) );
  OR2_X1 U10679 ( .A1(n8563), .A2(n8255), .ZN(n8256) );
  AND2_X1 U10680 ( .A1(n8233), .A2(n12984), .ZN(n8260) );
  OR2_X1 U10681 ( .A1(n8261), .A2(n8260), .ZN(n8264) );
  NAND2_X1 U10682 ( .A1(n8261), .A2(n8260), .ZN(n8262) );
  NAND2_X1 U10683 ( .A1(n8264), .A2(n8262), .ZN(n10362) );
  XNOR2_X1 U10684 ( .A(n8266), .B(n8265), .ZN(n9987) );
  NAND2_X1 U10685 ( .A1(n9987), .A2(n9780), .ZN(n8273) );
  NAND2_X1 U10686 ( .A1(n8268), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8267) );
  MUX2_X1 U10687 ( .A(n8267), .B(P2_IR_REG_31__SCAN_IN), .S(n8269), .Z(n8271)
         );
  INV_X1 U10688 ( .A(n8268), .ZN(n8270) );
  NAND2_X1 U10689 ( .A1(n8270), .A2(n8269), .ZN(n8313) );
  NAND2_X1 U10690 ( .A1(n8271), .A2(n8313), .ZN(n10087) );
  INV_X1 U10691 ( .A(n10087), .ZN(n10126) );
  AOI22_X1 U10692 ( .A1(n8694), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10126), 
        .B2(n8389), .ZN(n8272) );
  NAND2_X1 U10693 ( .A1(n8273), .A2(n8272), .ZN(n10640) );
  XNOR2_X1 U10694 ( .A(n10640), .B(n8745), .ZN(n8284) );
  INV_X2 U10695 ( .A(n8274), .ZN(n13219) );
  NAND2_X1 U10696 ( .A1(n9770), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8283) );
  INV_X1 U10697 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10077) );
  OR2_X1 U10698 ( .A1(n8662), .A2(n10077), .ZN(n8282) );
  INV_X1 U10699 ( .A(n8277), .ZN(n8275) );
  NAND2_X1 U10700 ( .A1(n8275), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8297) );
  INV_X1 U10701 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U10702 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  NAND2_X1 U10703 ( .A1(n8297), .A2(n8278), .ZN(n10638) );
  OR2_X1 U10704 ( .A1(n8414), .A2(n10638), .ZN(n8281) );
  INV_X1 U10705 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n8279) );
  OR2_X1 U10706 ( .A1(n8956), .A2(n8279), .ZN(n8280) );
  NAND4_X1 U10707 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n12983) );
  NAND2_X1 U10708 ( .A1(n13219), .A2(n12983), .ZN(n8285) );
  NAND2_X1 U10709 ( .A1(n8284), .A2(n8285), .ZN(n8289) );
  INV_X1 U10710 ( .A(n8284), .ZN(n8287) );
  INV_X1 U10711 ( .A(n8285), .ZN(n8286) );
  NAND2_X1 U10712 ( .A1(n8287), .A2(n8286), .ZN(n8288) );
  AND2_X1 U10713 ( .A1(n8289), .A2(n8288), .ZN(n10467) );
  XNOR2_X1 U10714 ( .A(n8291), .B(n8290), .ZN(n9999) );
  NAND2_X1 U10715 ( .A1(n9999), .A2(n9780), .ZN(n8294) );
  NAND2_X1 U10716 ( .A1(n8313), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8292) );
  XNOR2_X1 U10717 ( .A(n8292), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U10718 ( .A1(n8694), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10127), 
        .B2(n8389), .ZN(n8293) );
  XNOR2_X1 U10719 ( .A(n15106), .B(n8745), .ZN(n8305) );
  NAND2_X1 U10720 ( .A1(n8658), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8303) );
  INV_X1 U10721 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n13252) );
  OR2_X1 U10722 ( .A1(n8662), .A2(n13252), .ZN(n8302) );
  INV_X1 U10723 ( .A(n8297), .ZN(n8295) );
  NAND2_X1 U10724 ( .A1(n8295), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8319) );
  INV_X1 U10725 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10726 ( .A1(n8297), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U10727 ( .A1(n8319), .A2(n8298), .ZN(n10480) );
  OR2_X1 U10728 ( .A1(n8414), .A2(n10480), .ZN(n8301) );
  INV_X1 U10729 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n8299) );
  OR2_X1 U10730 ( .A1(n8563), .A2(n8299), .ZN(n8300) );
  NAND4_X1 U10731 ( .A1(n8303), .A2(n8302), .A3(n8301), .A4(n8300), .ZN(n12982) );
  XNOR2_X1 U10732 ( .A(n8305), .B(n8306), .ZN(n10479) );
  INV_X1 U10733 ( .A(n10479), .ZN(n8304) );
  INV_X1 U10734 ( .A(n8305), .ZN(n8308) );
  INV_X1 U10735 ( .A(n8306), .ZN(n8307) );
  NAND2_X1 U10736 ( .A1(n8308), .A2(n8307), .ZN(n8309) );
  XNOR2_X1 U10737 ( .A(n8311), .B(n8312), .ZN(n10003) );
  NAND2_X1 U10738 ( .A1(n10003), .A2(n9780), .ZN(n8316) );
  OAI21_X1 U10739 ( .B1(n8313), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8314) );
  XNOR2_X1 U10740 ( .A(n8314), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U10741 ( .A1(n8694), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10155), 
        .B2(n8389), .ZN(n8315) );
  NAND2_X1 U10742 ( .A1(n8316), .A2(n8315), .ZN(n10632) );
  XNOR2_X1 U10743 ( .A(n10632), .B(n8718), .ZN(n8328) );
  NAND2_X1 U10744 ( .A1(n8658), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8325) );
  INV_X1 U10745 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10660) );
  OR2_X1 U10746 ( .A1(n8662), .A2(n10660), .ZN(n8324) );
  INV_X1 U10747 ( .A(n8319), .ZN(n8317) );
  NAND2_X1 U10748 ( .A1(n8317), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8339) );
  INV_X1 U10749 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n8318) );
  NAND2_X1 U10750 ( .A1(n8319), .A2(n8318), .ZN(n8320) );
  NAND2_X1 U10751 ( .A1(n8339), .A2(n8320), .ZN(n10661) );
  OR2_X1 U10752 ( .A1(n8414), .A2(n10661), .ZN(n8323) );
  INV_X1 U10753 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n8321) );
  OR2_X1 U10754 ( .A1(n8563), .A2(n8321), .ZN(n8322) );
  NAND4_X1 U10755 ( .A1(n8325), .A2(n8324), .A3(n8323), .A4(n8322), .ZN(n12981) );
  NAND2_X1 U10756 ( .A1(n13219), .A2(n12981), .ZN(n8326) );
  XNOR2_X1 U10757 ( .A(n8328), .B(n8326), .ZN(n10628) );
  INV_X1 U10758 ( .A(n8326), .ZN(n8327) );
  NAND2_X1 U10759 ( .A1(n8328), .A2(n8327), .ZN(n8329) );
  XNOR2_X1 U10760 ( .A(n8331), .B(n8330), .ZN(n10015) );
  NAND2_X1 U10761 ( .A1(n10015), .A2(n9780), .ZN(n8336) );
  OR2_X1 U10762 ( .A1(n8332), .A2(n8333), .ZN(n8334) );
  XNOR2_X1 U10763 ( .A(n8334), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10184) );
  AOI22_X1 U10764 ( .A1(n8694), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10184), 
        .B2(n8389), .ZN(n8335) );
  XNOR2_X1 U10765 ( .A(n15116), .B(n8718), .ZN(n10704) );
  NAND2_X1 U10766 ( .A1(n9770), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n8344) );
  INV_X1 U10767 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8338) );
  OR2_X1 U10768 ( .A1(n8662), .A2(n8338), .ZN(n8343) );
  NAND2_X1 U10769 ( .A1(n8339), .A2(n13652), .ZN(n8340) );
  NAND2_X1 U10770 ( .A1(n8354), .A2(n8340), .ZN(n10776) );
  OR2_X1 U10771 ( .A1(n8414), .A2(n10776), .ZN(n8342) );
  INV_X1 U10772 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10152) );
  OR2_X1 U10773 ( .A1(n8956), .A2(n10152), .ZN(n8341) );
  NAND4_X1 U10774 ( .A1(n8344), .A2(n8343), .A3(n8342), .A4(n8341), .ZN(n12980) );
  AND2_X1 U10775 ( .A1(n13219), .A2(n12980), .ZN(n10705) );
  NAND2_X1 U10776 ( .A1(n10995), .A2(n10705), .ZN(n8361) );
  XNOR2_X1 U10777 ( .A(n8345), .B(n8346), .ZN(n10019) );
  NAND2_X1 U10778 ( .A1(n10019), .A2(n9780), .ZN(n8350) );
  NAND2_X1 U10779 ( .A1(n8332), .A2(n8347), .ZN(n8368) );
  NAND2_X1 U10780 ( .A1(n8368), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8348) );
  XNOR2_X1 U10781 ( .A(n8348), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10495) );
  AOI22_X1 U10782 ( .A1(n8694), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10495), 
        .B2(n8389), .ZN(n8349) );
  XNOR2_X1 U10783 ( .A(n15126), .B(n8745), .ZN(n8363) );
  NAND2_X1 U10784 ( .A1(n9770), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n8359) );
  INV_X1 U10785 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8351) );
  OR2_X1 U10786 ( .A1(n8662), .A2(n8351), .ZN(n8358) );
  INV_X1 U10787 ( .A(n8354), .ZN(n8352) );
  NAND2_X1 U10788 ( .A1(n8352), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8373) );
  INV_X1 U10789 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10790 ( .A1(n8354), .A2(n8353), .ZN(n8355) );
  NAND2_X1 U10791 ( .A1(n8373), .A2(n8355), .ZN(n11003) );
  OR2_X1 U10792 ( .A1(n8414), .A2(n11003), .ZN(n8357) );
  INV_X1 U10793 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10179) );
  OR2_X1 U10794 ( .A1(n8956), .A2(n10179), .ZN(n8356) );
  NAND4_X1 U10795 ( .A1(n8359), .A2(n8358), .A3(n8357), .A4(n8356), .ZN(n12979) );
  NAND2_X1 U10796 ( .A1(n13219), .A2(n12979), .ZN(n8362) );
  XNOR2_X1 U10797 ( .A(n8363), .B(n8362), .ZN(n10999) );
  NAND2_X1 U10798 ( .A1(n8363), .A2(n8362), .ZN(n8364) );
  XNOR2_X1 U10799 ( .A(n8366), .B(SI_10_), .ZN(n8367) );
  XNOR2_X1 U10800 ( .A(n8365), .B(n8367), .ZN(n10023) );
  NAND2_X1 U10801 ( .A1(n10023), .A2(n9780), .ZN(n8371) );
  NAND2_X1 U10802 ( .A1(n8510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8369) );
  XNOR2_X1 U10803 ( .A(n8369), .B(n8386), .ZN(n14990) );
  AOI22_X1 U10804 ( .A1(n8694), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n14990), 
        .B2(n8389), .ZN(n8370) );
  XNOR2_X1 U10805 ( .A(n15136), .B(n8718), .ZN(n11331) );
  NAND2_X1 U10806 ( .A1(n9770), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8378) );
  INV_X1 U10807 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8372) );
  OR2_X1 U10808 ( .A1(n8662), .A2(n8372), .ZN(n8377) );
  NAND2_X1 U10809 ( .A1(n8373), .A2(n14984), .ZN(n8374) );
  NAND2_X1 U10810 ( .A1(n8395), .A2(n8374), .ZN(n10841) );
  OR2_X1 U10811 ( .A1(n8414), .A2(n10841), .ZN(n8376) );
  INV_X1 U10812 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10496) );
  OR2_X1 U10813 ( .A1(n8956), .A2(n10496), .ZN(n8375) );
  NAND4_X1 U10814 ( .A1(n8378), .A2(n8377), .A3(n8376), .A4(n8375), .ZN(n12978) );
  AND2_X1 U10815 ( .A1(n13219), .A2(n12978), .ZN(n8379) );
  NAND2_X1 U10816 ( .A1(n11331), .A2(n8379), .ZN(n8383) );
  INV_X1 U10817 ( .A(n11331), .ZN(n8381) );
  INV_X1 U10818 ( .A(n8379), .ZN(n8380) );
  NAND2_X1 U10819 ( .A1(n8381), .A2(n8380), .ZN(n8382) );
  AND2_X1 U10820 ( .A1(n8383), .A2(n8382), .ZN(n11049) );
  XNOR2_X1 U10821 ( .A(n8384), .B(n8385), .ZN(n10050) );
  NAND2_X1 U10822 ( .A1(n10050), .A2(n9780), .ZN(n8391) );
  NOR2_X1 U10823 ( .A1(n8510), .A2(n8386), .ZN(n8407) );
  INV_X1 U10824 ( .A(n8407), .ZN(n8387) );
  NAND2_X1 U10825 ( .A1(n8387), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8388) );
  XNOR2_X1 U10826 ( .A(n8388), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U10827 ( .A1(n8694), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10541), 
        .B2(n8389), .ZN(n8390) );
  XNOR2_X1 U10828 ( .A(n15028), .B(n8718), .ZN(n8401) );
  NAND2_X1 U10829 ( .A1(n9770), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8400) );
  INV_X1 U10830 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8392) );
  OR2_X1 U10831 ( .A1(n8662), .A2(n8392), .ZN(n8399) );
  INV_X1 U10832 ( .A(n8395), .ZN(n8393) );
  NAND2_X1 U10833 ( .A1(n8393), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8412) );
  INV_X1 U10834 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10835 ( .A1(n8395), .A2(n8394), .ZN(n8396) );
  NAND2_X1 U10836 ( .A1(n8412), .A2(n8396), .ZN(n15025) );
  OR2_X1 U10837 ( .A1(n8414), .A2(n15025), .ZN(n8398) );
  INV_X1 U10838 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10497) );
  OR2_X1 U10839 ( .A1(n8956), .A2(n10497), .ZN(n8397) );
  NAND4_X1 U10840 ( .A1(n8400), .A2(n8399), .A3(n8398), .A4(n8397), .ZN(n12977) );
  AND2_X1 U10841 ( .A1(n13219), .A2(n12977), .ZN(n8402) );
  NAND2_X1 U10842 ( .A1(n8401), .A2(n8402), .ZN(n8419) );
  INV_X1 U10843 ( .A(n8401), .ZN(n11355) );
  INV_X1 U10844 ( .A(n8402), .ZN(n8403) );
  NAND2_X1 U10845 ( .A1(n11355), .A2(n8403), .ZN(n8404) );
  AND2_X1 U10846 ( .A1(n8419), .A2(n8404), .ZN(n11332) );
  XNOR2_X1 U10847 ( .A(n8405), .B(n7436), .ZN(n10173) );
  NAND2_X1 U10848 ( .A1(n10173), .A2(n9780), .ZN(n8411) );
  INV_X1 U10849 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n8406) );
  INV_X1 U10850 ( .A(n8427), .ZN(n8408) );
  NAND2_X1 U10851 ( .A1(n8408), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8409) );
  XNOR2_X1 U10852 ( .A(n8409), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10796) );
  AOI22_X1 U10853 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n8694), .B1(n10796), 
        .B2(n8389), .ZN(n8410) );
  XNOR2_X1 U10854 ( .A(n13348), .B(n8718), .ZN(n8421) );
  NAND2_X1 U10855 ( .A1(n9769), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n8418) );
  INV_X1 U10856 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n13551) );
  OR2_X1 U10857 ( .A1(n8563), .A2(n13551), .ZN(n8417) );
  NAND2_X1 U10858 ( .A1(n8412), .A2(n10550), .ZN(n8413) );
  NAND2_X1 U10859 ( .A1(n8433), .A2(n8413), .ZN(n11361) );
  OR2_X1 U10860 ( .A1(n8414), .A2(n11361), .ZN(n8416) );
  INV_X1 U10861 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10539) );
  OR2_X1 U10862 ( .A1(n8956), .A2(n10539), .ZN(n8415) );
  NAND4_X1 U10863 ( .A1(n8418), .A2(n8417), .A3(n8416), .A4(n8415), .ZN(n12976) );
  NAND2_X1 U10864 ( .A1(n13219), .A2(n12976), .ZN(n8422) );
  XNOR2_X1 U10865 ( .A(n8421), .B(n8422), .ZN(n11366) );
  AND2_X1 U10866 ( .A1(n11366), .A2(n8419), .ZN(n8420) );
  INV_X1 U10867 ( .A(n8421), .ZN(n8423) );
  NAND2_X1 U10868 ( .A1(n8423), .A2(n8422), .ZN(n8424) );
  XNOR2_X1 U10869 ( .A(n8425), .B(n7437), .ZN(n10226) );
  NAND2_X1 U10870 ( .A1(n10226), .A2(n9780), .ZN(n8431) );
  INV_X1 U10871 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8426) );
  INV_X1 U10872 ( .A(n8448), .ZN(n8428) );
  NAND2_X1 U10873 ( .A1(n8428), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8429) );
  XNOR2_X1 U10874 ( .A(n8429), .B(P2_IR_REG_13__SCAN_IN), .ZN(n11153) );
  AOI22_X1 U10875 ( .A1(n11153), .A2(n8389), .B1(P1_DATAO_REG_13__SCAN_IN), 
        .B2(n8694), .ZN(n8430) );
  XNOR2_X1 U10876 ( .A(n14650), .B(n8718), .ZN(n12795) );
  NAND2_X1 U10877 ( .A1(n8433), .A2(n8432), .ZN(n8434) );
  NAND2_X1 U10878 ( .A1(n8453), .A2(n8434), .ZN(n12905) );
  INV_X1 U10879 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10802) );
  OR2_X1 U10880 ( .A1(n8662), .A2(n10802), .ZN(n8435) );
  OAI21_X1 U10881 ( .B1(n12905), .B2(n8414), .A(n8435), .ZN(n8439) );
  INV_X1 U10882 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10797) );
  INV_X1 U10883 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8436) );
  OR2_X1 U10884 ( .A1(n8563), .A2(n8436), .ZN(n8437) );
  OAI21_X1 U10885 ( .B1(n8956), .B2(n10797), .A(n8437), .ZN(n8438) );
  AND2_X1 U10886 ( .A1(n12975), .A2(n13219), .ZN(n8440) );
  NAND2_X1 U10887 ( .A1(n12795), .A2(n8440), .ZN(n8460) );
  INV_X1 U10888 ( .A(n12795), .ZN(n8442) );
  INV_X1 U10889 ( .A(n8440), .ZN(n8441) );
  NAND2_X1 U10890 ( .A1(n8442), .A2(n8441), .ZN(n8443) );
  NAND2_X1 U10891 ( .A1(n8460), .A2(n8443), .ZN(n12908) );
  INV_X1 U10892 ( .A(n12908), .ZN(n8444) );
  NAND2_X1 U10893 ( .A1(n8445), .A2(n10120), .ZN(n8466) );
  OR2_X1 U10894 ( .A1(n8445), .A2(n10120), .ZN(n8446) );
  NAND2_X1 U10895 ( .A1(n8466), .A2(n8446), .ZN(n8468) );
  XNOR2_X1 U10896 ( .A(n8468), .B(n8467), .ZN(n10385) );
  NAND2_X1 U10897 ( .A1(n10385), .A2(n9780), .ZN(n8451) );
  INV_X1 U10898 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U10899 ( .A1(n8448), .A2(n8447), .ZN(n8472) );
  NAND2_X1 U10900 ( .A1(n8472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8449) );
  XNOR2_X1 U10901 ( .A(n8449), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11658) );
  AOI22_X1 U10902 ( .A1(n11658), .A2(n8389), .B1(P1_DATAO_REG_14__SCAN_IN), 
        .B2(n8694), .ZN(n8450) );
  XNOR2_X1 U10903 ( .A(n13344), .B(n8718), .ZN(n8462) );
  INV_X1 U10904 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8459) );
  INV_X1 U10905 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U10906 ( .A1(n8453), .A2(n12801), .ZN(n8454) );
  NAND2_X1 U10907 ( .A1(n8479), .A2(n8454), .ZN(n12800) );
  OR2_X1 U10908 ( .A1(n12800), .A2(n8414), .ZN(n8458) );
  NAND2_X1 U10909 ( .A1(n9770), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10910 ( .A1(n9769), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8455) );
  AND2_X1 U10911 ( .A1(n8456), .A2(n8455), .ZN(n8457) );
  OAI211_X1 U10912 ( .C1(n8956), .C2(n8459), .A(n8458), .B(n8457), .ZN(n12974)
         );
  NAND2_X1 U10913 ( .A1(n12974), .A2(n13219), .ZN(n8463) );
  XNOR2_X1 U10914 ( .A(n8462), .B(n8463), .ZN(n12797) );
  AND2_X1 U10915 ( .A1(n12797), .A2(n8460), .ZN(n8461) );
  NAND2_X1 U10916 ( .A1(n12794), .A2(n8461), .ZN(n12807) );
  INV_X1 U10917 ( .A(n8462), .ZN(n8464) );
  NAND2_X1 U10918 ( .A1(n8464), .A2(n8463), .ZN(n8465) );
  NAND2_X1 U10919 ( .A1(n12807), .A2(n8465), .ZN(n8484) );
  OAI21_X1 U10920 ( .B1(n8468), .B2(n8467), .A(n8466), .ZN(n8471) );
  INV_X1 U10921 ( .A(n8469), .ZN(n8470) );
  XNOR2_X1 U10922 ( .A(n8471), .B(n8470), .ZN(n10420) );
  NAND2_X1 U10923 ( .A1(n10420), .A2(n9780), .ZN(n8476) );
  NAND2_X1 U10924 ( .A1(n8473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8489) );
  XNOR2_X1 U10925 ( .A(n8489), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11648) );
  NOR2_X1 U10926 ( .A1(n8227), .A2(n13634), .ZN(n8474) );
  AOI21_X1 U10927 ( .B1(n11648), .B2(n8389), .A(n8474), .ZN(n8475) );
  XNOR2_X1 U10928 ( .A(n12955), .B(n8718), .ZN(n8485) );
  XNOR2_X1 U10929 ( .A(n8484), .B(n8485), .ZN(n12947) );
  INV_X1 U10930 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15003) );
  INV_X1 U10931 ( .A(n8479), .ZN(n8477) );
  NAND2_X1 U10932 ( .A1(n8477), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8495) );
  INV_X1 U10933 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8478) );
  NAND2_X1 U10934 ( .A1(n8479), .A2(n8478), .ZN(n8480) );
  NAND2_X1 U10935 ( .A1(n8495), .A2(n8480), .ZN(n12952) );
  OR2_X1 U10936 ( .A1(n12952), .A2(n8414), .ZN(n8482) );
  AOI22_X1 U10937 ( .A1(n9769), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9770), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n8481) );
  OAI211_X1 U10938 ( .C1(n8956), .C2(n15003), .A(n8482), .B(n8481), .ZN(n12973) );
  AND2_X1 U10939 ( .A1(n12973), .A2(n13219), .ZN(n8483) );
  INV_X1 U10940 ( .A(n8484), .ZN(n8486) );
  NAND2_X1 U10941 ( .A1(n8486), .A2(n8485), .ZN(n8487) );
  XNOR2_X1 U10942 ( .A(n6583), .B(n7425), .ZN(n10346) );
  NAND2_X1 U10943 ( .A1(n10346), .A2(n9780), .ZN(n8494) );
  NAND2_X1 U10944 ( .A1(n8489), .A2(n8488), .ZN(n8490) );
  NAND2_X1 U10945 ( .A1(n8490), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8491) );
  XNOR2_X1 U10946 ( .A(n8491), .B(P2_IR_REG_16__SCAN_IN), .ZN(n13005) );
  NOR2_X1 U10947 ( .A1(n8227), .A2(n10369), .ZN(n8492) );
  AOI21_X1 U10948 ( .B1(n13005), .B2(n8389), .A(n8492), .ZN(n8493) );
  XNOR2_X1 U10949 ( .A(n13339), .B(n8745), .ZN(n12875) );
  NAND2_X1 U10950 ( .A1(n8495), .A2(n12862), .ZN(n8496) );
  AND2_X1 U10951 ( .A1(n8516), .A2(n8496), .ZN(n12865) );
  NAND2_X1 U10952 ( .A1(n12865), .A2(n8789), .ZN(n8501) );
  INV_X1 U10953 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11651) );
  NAND2_X1 U10954 ( .A1(n9770), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U10955 ( .A1(n8658), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U10956 ( .C1(n8662), .C2(n11651), .A(n8498), .B(n8497), .ZN(n8499)
         );
  INV_X1 U10957 ( .A(n8499), .ZN(n8500) );
  NAND2_X1 U10958 ( .A1(n8501), .A2(n8500), .ZN(n12972) );
  NAND2_X1 U10959 ( .A1(n12972), .A2(n13219), .ZN(n8503) );
  XNOR2_X1 U10960 ( .A(n12875), .B(n8503), .ZN(n12861) );
  NAND2_X1 U10961 ( .A1(n12875), .A2(n8503), .ZN(n8504) );
  NAND2_X1 U10962 ( .A1(n12878), .A2(n8504), .ZN(n8524) );
  XNOR2_X1 U10963 ( .A(n8505), .B(SI_17_), .ZN(n8506) );
  XNOR2_X1 U10964 ( .A(n8507), .B(n8506), .ZN(n10421) );
  NAND2_X1 U10965 ( .A1(n10421), .A2(n9780), .ZN(n8513) );
  CLKBUF_X1 U10966 ( .A(n8508), .Z(n8509) );
  OAI21_X1 U10967 ( .B1(n8510), .B2(n8509), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8511) );
  XNOR2_X1 U10968 ( .A(n8511), .B(P2_IR_REG_17__SCAN_IN), .ZN(n13024) );
  AOI22_X1 U10969 ( .A1(n8694), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n13024), 
        .B2(n8389), .ZN(n8512) );
  XNOR2_X1 U10970 ( .A(n13237), .B(n8745), .ZN(n8525) );
  INV_X1 U10971 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8515) );
  NAND2_X1 U10972 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  NAND2_X1 U10973 ( .A1(n8539), .A2(n8517), .ZN(n13233) );
  OR2_X1 U10974 ( .A1(n13233), .A2(n8414), .ZN(n8523) );
  INV_X1 U10975 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8520) );
  NAND2_X1 U10976 ( .A1(n9770), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U10977 ( .A1(n9769), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8518) );
  OAI211_X1 U10978 ( .C1(n8520), .C2(n8956), .A(n8519), .B(n8518), .ZN(n8521)
         );
  INV_X1 U10979 ( .A(n8521), .ZN(n8522) );
  NAND2_X1 U10980 ( .A1(n12971), .A2(n13219), .ZN(n8526) );
  XNOR2_X1 U10981 ( .A(n8525), .B(n8526), .ZN(n12873) );
  INV_X1 U10982 ( .A(n8525), .ZN(n8527) );
  NAND2_X1 U10983 ( .A1(n8527), .A2(n8526), .ZN(n8528) );
  XNOR2_X1 U10984 ( .A(n8551), .B(SI_18_), .ZN(n8530) );
  INV_X1 U10985 ( .A(n8530), .ZN(n8532) );
  OR2_X1 U10986 ( .A1(n10538), .A2(n8693), .ZN(n8537) );
  NAND2_X1 U10987 ( .A1(n8534), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8535) );
  XNOR2_X1 U10988 ( .A(n8535), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U10989 ( .A1(n8694), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n13033), 
        .B2(n8389), .ZN(n8536) );
  XNOR2_X1 U10990 ( .A(n13328), .B(n8718), .ZN(n12825) );
  NAND2_X1 U10991 ( .A1(n8539), .A2(n8538), .ZN(n8540) );
  AND2_X1 U10992 ( .A1(n8561), .A2(n8540), .ZN(n13222) );
  NAND2_X1 U10993 ( .A1(n13222), .A2(n8789), .ZN(n8545) );
  INV_X1 U10994 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U10995 ( .A1(n9770), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8542) );
  NAND2_X1 U10996 ( .A1(n9769), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8541) );
  OAI211_X1 U10997 ( .C1(n13026), .C2(n8956), .A(n8542), .B(n8541), .ZN(n8543)
         );
  INV_X1 U10998 ( .A(n8543), .ZN(n8544) );
  NAND2_X1 U10999 ( .A1(n8545), .A2(n8544), .ZN(n12970) );
  AND2_X1 U11000 ( .A1(n12970), .A2(n13219), .ZN(n8546) );
  NAND2_X1 U11001 ( .A1(n12825), .A2(n8546), .ZN(n8569) );
  INV_X1 U11002 ( .A(n12825), .ZN(n8548) );
  INV_X1 U11003 ( .A(n8546), .ZN(n8547) );
  NAND2_X1 U11004 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  NAND2_X1 U11005 ( .A1(n8569), .A2(n8549), .ZN(n12920) );
  INV_X1 U11006 ( .A(n12920), .ZN(n8550) );
  INV_X1 U11007 ( .A(SI_18_), .ZN(n13617) );
  OR2_X1 U11008 ( .A1(n8551), .A2(n13617), .ZN(n8552) );
  NAND2_X1 U11009 ( .A1(n8553), .A2(n8552), .ZN(n8556) );
  XNOR2_X1 U11010 ( .A(n8554), .B(SI_19_), .ZN(n8555) );
  XNOR2_X1 U11011 ( .A(n8556), .B(n8555), .ZN(n10685) );
  NAND2_X1 U11012 ( .A1(n10685), .A2(n9780), .ZN(n8558) );
  AOI22_X1 U11013 ( .A1(n8694), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9844), 
        .B2(n8389), .ZN(n8557) );
  XNOR2_X1 U11014 ( .A(n13323), .B(n8718), .ZN(n8571) );
  INV_X1 U11015 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U11016 ( .A1(n8561), .A2(n8560), .ZN(n8562) );
  NAND2_X1 U11017 ( .A1(n8580), .A2(n8562), .ZN(n13208) );
  OR2_X1 U11018 ( .A1(n13208), .A2(n8414), .ZN(n8568) );
  INV_X1 U11019 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13041) );
  NAND2_X1 U11020 ( .A1(n9769), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n8565) );
  INV_X1 U11021 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n13468) );
  OR2_X1 U11022 ( .A1(n8563), .A2(n13468), .ZN(n8564) );
  OAI211_X1 U11023 ( .C1(n13041), .C2(n8956), .A(n8565), .B(n8564), .ZN(n8566)
         );
  INV_X1 U11024 ( .A(n8566), .ZN(n8567) );
  NAND2_X1 U11025 ( .A1(n8568), .A2(n8567), .ZN(n12969) );
  NAND2_X1 U11026 ( .A1(n12969), .A2(n13219), .ZN(n8572) );
  XNOR2_X1 U11027 ( .A(n8571), .B(n8572), .ZN(n12827) );
  AND2_X1 U11028 ( .A1(n12827), .A2(n8569), .ZN(n8570) );
  NAND2_X1 U11029 ( .A1(n12824), .A2(n8570), .ZN(n12823) );
  INV_X1 U11030 ( .A(n8571), .ZN(n12897) );
  NAND2_X1 U11031 ( .A1(n12897), .A2(n8572), .ZN(n8573) );
  NAND2_X1 U11032 ( .A1(n12823), .A2(n8573), .ZN(n8588) );
  NAND2_X1 U11033 ( .A1(n8575), .A2(n8574), .ZN(n8576) );
  NAND2_X1 U11034 ( .A1(n8577), .A2(n8576), .ZN(n10683) );
  OR2_X1 U11035 ( .A1(n10683), .A2(n8693), .ZN(n8579) );
  NAND2_X1 U11036 ( .A1(n8694), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8578) );
  XNOR2_X1 U11037 ( .A(n13318), .B(n8718), .ZN(n8589) );
  INV_X1 U11038 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U11039 ( .A1(n8580), .A2(n12892), .ZN(n8581) );
  AND2_X1 U11040 ( .A1(n8600), .A2(n8581), .ZN(n13193) );
  NAND2_X1 U11041 ( .A1(n13193), .A2(n8789), .ZN(n8587) );
  INV_X1 U11042 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8584) );
  NAND2_X1 U11043 ( .A1(n9770), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U11044 ( .A1(n8658), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8582) );
  OAI211_X1 U11045 ( .C1(n8662), .C2(n8584), .A(n8583), .B(n8582), .ZN(n8585)
         );
  INV_X1 U11046 ( .A(n8585), .ZN(n8586) );
  NAND2_X1 U11047 ( .A1(n8587), .A2(n8586), .ZN(n12968) );
  NAND2_X1 U11048 ( .A1(n12968), .A2(n13219), .ZN(n8590) );
  XNOR2_X1 U11049 ( .A(n8589), .B(n8590), .ZN(n12895) );
  INV_X1 U11050 ( .A(n8589), .ZN(n8591) );
  NAND2_X1 U11051 ( .A1(n8591), .A2(n8590), .ZN(n8592) );
  OR2_X1 U11052 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U11053 ( .A1(n8596), .A2(n8595), .ZN(n10812) );
  OR2_X1 U11054 ( .A1(n10812), .A2(n8693), .ZN(n8598) );
  NAND2_X1 U11055 ( .A1(n8694), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8597) );
  XNOR2_X1 U11056 ( .A(n13312), .B(n8745), .ZN(n8609) );
  INV_X1 U11057 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12841) );
  NAND2_X1 U11058 ( .A1(n8600), .A2(n12841), .ZN(n8601) );
  NAND2_X1 U11059 ( .A1(n8631), .A2(n8601), .ZN(n13174) );
  OR2_X1 U11060 ( .A1(n13174), .A2(n8414), .ZN(n8607) );
  INV_X1 U11061 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8604) );
  NAND2_X1 U11062 ( .A1(n9770), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n8603) );
  NAND2_X1 U11063 ( .A1(n9769), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8602) );
  OAI211_X1 U11064 ( .C1(n8604), .C2(n8956), .A(n8603), .B(n8602), .ZN(n8605)
         );
  INV_X1 U11065 ( .A(n8605), .ZN(n8606) );
  NAND2_X1 U11066 ( .A1(n8607), .A2(n8606), .ZN(n12967) );
  NAND2_X1 U11067 ( .A1(n12967), .A2(n13219), .ZN(n8610) );
  XNOR2_X1 U11068 ( .A(n8609), .B(n8610), .ZN(n12835) );
  INV_X1 U11069 ( .A(n12835), .ZN(n8608) );
  INV_X1 U11070 ( .A(n8609), .ZN(n8612) );
  INV_X1 U11071 ( .A(n8610), .ZN(n8611) );
  NAND2_X1 U11072 ( .A1(n8612), .A2(n8611), .ZN(n8613) );
  NAND2_X1 U11073 ( .A1(n12837), .A2(n8613), .ZN(n8643) );
  NAND2_X1 U11074 ( .A1(n9368), .A2(n8614), .ZN(n8615) );
  NAND2_X1 U11075 ( .A1(n8616), .A2(n8615), .ZN(n11058) );
  OR2_X1 U11076 ( .A1(n11058), .A2(n8693), .ZN(n8618) );
  NAND2_X1 U11077 ( .A1(n8694), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8617) );
  XNOR2_X1 U11078 ( .A(n13307), .B(n8745), .ZN(n8641) );
  XNOR2_X1 U11079 ( .A(n8619), .B(SI_23_), .ZN(n11378) );
  NAND2_X1 U11080 ( .A1(n11378), .A2(n9780), .ZN(n8621) );
  NAND2_X1 U11081 ( .A1(n8694), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8620) );
  XNOR2_X1 U11082 ( .A(n13302), .B(n8745), .ZN(n12812) );
  INV_X1 U11083 ( .A(n8631), .ZN(n8622) );
  NAND2_X1 U11084 ( .A1(n8622), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8633) );
  INV_X1 U11085 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U11086 ( .A1(n8633), .A2(n12818), .ZN(n8623) );
  NAND2_X1 U11087 ( .A1(n8656), .A2(n8623), .ZN(n13149) );
  OR2_X1 U11088 ( .A1(n13149), .A2(n8414), .ZN(n8629) );
  INV_X1 U11089 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11090 ( .A1(n9770), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8625) );
  NAND2_X1 U11091 ( .A1(n9769), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8624) );
  OAI211_X1 U11092 ( .C1(n8626), .C2(n8956), .A(n8625), .B(n8624), .ZN(n8627)
         );
  INV_X1 U11093 ( .A(n8627), .ZN(n8628) );
  NAND2_X1 U11094 ( .A1(n8629), .A2(n8628), .ZN(n12913) );
  INV_X1 U11095 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U11096 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  NAND2_X1 U11097 ( .A1(n8633), .A2(n8632), .ZN(n12914) );
  OR2_X1 U11098 ( .A1(n12914), .A2(n8414), .ZN(n8639) );
  INV_X1 U11099 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8636) );
  NAND2_X1 U11100 ( .A1(n9770), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8635) );
  NAND2_X1 U11101 ( .A1(n9769), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8634) );
  OAI211_X1 U11102 ( .C1(n8636), .C2(n8956), .A(n8635), .B(n8634), .ZN(n8637)
         );
  INV_X1 U11103 ( .A(n8637), .ZN(n8638) );
  NAND2_X1 U11104 ( .A1(n12966), .A2(n13219), .ZN(n12809) );
  AOI21_X1 U11105 ( .B1(n12812), .B2(n12885), .A(n12809), .ZN(n8640) );
  NAND2_X1 U11106 ( .A1(n12808), .A2(n8640), .ZN(n8649) );
  INV_X1 U11107 ( .A(n8641), .ZN(n8642) );
  AND2_X1 U11108 ( .A1(n8643), .A2(n8642), .ZN(n12811) );
  AND2_X1 U11109 ( .A1(n12913), .A2(n13219), .ZN(n8644) );
  INV_X1 U11110 ( .A(n8644), .ZN(n12815) );
  NAND2_X1 U11111 ( .A1(n12812), .A2(n12815), .ZN(n8647) );
  INV_X1 U11112 ( .A(n12812), .ZN(n8645) );
  AND2_X1 U11113 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U11114 ( .A1(n8649), .A2(n8648), .ZN(n12882) );
  NAND2_X1 U11115 ( .A1(n8651), .A2(n8650), .ZN(n8652) );
  AND2_X1 U11116 ( .A1(n8653), .A2(n8652), .ZN(n11737) );
  NAND2_X1 U11117 ( .A1(n11737), .A2(n9780), .ZN(n8655) );
  NAND2_X1 U11118 ( .A1(n8694), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8654) );
  XNOR2_X1 U11119 ( .A(n13297), .B(n8718), .ZN(n8666) );
  INV_X1 U11120 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13650) );
  NAND2_X1 U11121 ( .A1(n8656), .A2(n13650), .ZN(n8657) );
  AND2_X1 U11122 ( .A1(n8676), .A2(n8657), .ZN(n13135) );
  NAND2_X1 U11123 ( .A1(n13135), .A2(n8789), .ZN(n8665) );
  INV_X1 U11124 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n8661) );
  NAND2_X1 U11125 ( .A1(n9770), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8660) );
  NAND2_X1 U11126 ( .A1(n8658), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8659) );
  OAI211_X1 U11127 ( .C1(n8662), .C2(n8661), .A(n8660), .B(n8659), .ZN(n8663)
         );
  INV_X1 U11128 ( .A(n8663), .ZN(n8664) );
  NAND2_X1 U11129 ( .A1(n8665), .A2(n8664), .ZN(n12965) );
  AND2_X1 U11130 ( .A1(n12965), .A2(n13219), .ZN(n8667) );
  NAND2_X1 U11131 ( .A1(n8666), .A2(n8667), .ZN(n8670) );
  INV_X1 U11132 ( .A(n8666), .ZN(n12848) );
  INV_X1 U11133 ( .A(n8667), .ZN(n8668) );
  NAND2_X1 U11134 ( .A1(n12848), .A2(n8668), .ZN(n8669) );
  AND2_X1 U11135 ( .A1(n8670), .A2(n8669), .ZN(n12883) );
  NAND2_X1 U11136 ( .A1(n12882), .A2(n12883), .ZN(n12845) );
  NAND2_X1 U11137 ( .A1(n12845), .A2(n8670), .ZN(n8688) );
  XNOR2_X1 U11138 ( .A(n8672), .B(n8671), .ZN(n13391) );
  NAND2_X1 U11139 ( .A1(n13391), .A2(n9780), .ZN(n8674) );
  NAND2_X1 U11140 ( .A1(n8694), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8673) );
  XNOR2_X1 U11141 ( .A(n13292), .B(n8718), .ZN(n8684) );
  INV_X1 U11142 ( .A(n8676), .ZN(n8675) );
  NAND2_X1 U11143 ( .A1(n8675), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n8699) );
  INV_X1 U11144 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12854) );
  NAND2_X1 U11145 ( .A1(n8676), .A2(n12854), .ZN(n8677) );
  NAND2_X1 U11146 ( .A1(n8699), .A2(n8677), .ZN(n13115) );
  OR2_X1 U11147 ( .A1(n13115), .A2(n8414), .ZN(n8683) );
  INV_X1 U11148 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11149 ( .A1(n9770), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U11150 ( .A1(n9769), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8678) );
  OAI211_X1 U11151 ( .C1(n8680), .C2(n8956), .A(n8679), .B(n8678), .ZN(n8681)
         );
  INV_X1 U11152 ( .A(n8681), .ZN(n8682) );
  NAND2_X1 U11153 ( .A1(n8683), .A2(n8682), .ZN(n12964) );
  AND2_X1 U11154 ( .A1(n12964), .A2(n13219), .ZN(n8685) );
  NAND2_X1 U11155 ( .A1(n8684), .A2(n8685), .ZN(n8707) );
  INV_X1 U11156 ( .A(n8684), .ZN(n12929) );
  INV_X1 U11157 ( .A(n8685), .ZN(n8686) );
  NAND2_X1 U11158 ( .A1(n12929), .A2(n8686), .ZN(n8687) );
  AND2_X1 U11159 ( .A1(n8707), .A2(n8687), .ZN(n12846) );
  NAND2_X1 U11160 ( .A1(n8688), .A2(n12846), .ZN(n12849) );
  NAND2_X1 U11161 ( .A1(n8690), .A2(n8689), .ZN(n8691) );
  OR2_X1 U11162 ( .A1(n13390), .A2(n8693), .ZN(n8696) );
  NAND2_X1 U11163 ( .A1(n8694), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8695) );
  NAND2_X2 U11164 ( .A1(n8696), .A2(n8695), .ZN(n13287) );
  XNOR2_X1 U11165 ( .A(n13287), .B(n8718), .ZN(n8709) );
  INV_X1 U11166 ( .A(n8699), .ZN(n8697) );
  INV_X1 U11167 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11168 ( .A1(n8699), .A2(n8698), .ZN(n8700) );
  NAND2_X1 U11169 ( .A1(n8734), .A2(n8700), .ZN(n12934) );
  OR2_X1 U11170 ( .A1(n12934), .A2(n8414), .ZN(n8706) );
  INV_X1 U11171 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8703) );
  NAND2_X1 U11172 ( .A1(n9770), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11173 ( .A1(n9769), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8701) );
  OAI211_X1 U11174 ( .C1(n8703), .C2(n8956), .A(n8702), .B(n8701), .ZN(n8704)
         );
  INV_X1 U11175 ( .A(n8704), .ZN(n8705) );
  NAND2_X1 U11176 ( .A1(n8706), .A2(n8705), .ZN(n12963) );
  NAND2_X1 U11177 ( .A1(n12963), .A2(n13219), .ZN(n8710) );
  XNOR2_X1 U11178 ( .A(n8709), .B(n8710), .ZN(n12943) );
  AND2_X1 U11179 ( .A1(n12943), .A2(n8707), .ZN(n8708) );
  INV_X1 U11180 ( .A(n8709), .ZN(n8711) );
  NAND2_X1 U11181 ( .A1(n8711), .A2(n8710), .ZN(n8712) );
  XNOR2_X1 U11182 ( .A(n8713), .B(SI_27_), .ZN(n8714) );
  NAND2_X1 U11183 ( .A1(n13384), .A2(n9780), .ZN(n8717) );
  NAND2_X1 U11184 ( .A1(n8694), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8716) );
  XNOR2_X1 U11185 ( .A(n13280), .B(n8718), .ZN(n8726) );
  XNOR2_X1 U11186 ( .A(n8734), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13086) );
  NAND2_X1 U11187 ( .A1(n13086), .A2(n8789), .ZN(n8725) );
  INV_X1 U11188 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11189 ( .A1(n9770), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U11190 ( .A1(n9769), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8720) );
  OAI211_X1 U11191 ( .C1(n8722), .C2(n8956), .A(n8721), .B(n8720), .ZN(n8723)
         );
  INV_X1 U11192 ( .A(n8723), .ZN(n8724) );
  AND2_X1 U11193 ( .A1(n12962), .A2(n13219), .ZN(n8727) );
  NAND2_X1 U11194 ( .A1(n8726), .A2(n8727), .ZN(n8732) );
  INV_X1 U11195 ( .A(n8726), .ZN(n8729) );
  INV_X1 U11196 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U11197 ( .A1(n8729), .A2(n8728), .ZN(n8730) );
  NAND2_X1 U11198 ( .A1(n8732), .A2(n8730), .ZN(n12782) );
  NAND2_X1 U11199 ( .A1(n12785), .A2(n8732), .ZN(n8748) );
  INV_X1 U11200 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12788) );
  INV_X1 U11201 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8733) );
  OAI21_X1 U11202 ( .B1(n8734), .B2(n12788), .A(n8733), .ZN(n8738) );
  INV_X1 U11203 ( .A(n8734), .ZN(n8736) );
  AND2_X1 U11204 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8735) );
  INV_X1 U11205 ( .A(n8898), .ZN(n8737) );
  NAND2_X1 U11206 ( .A1(n13072), .A2(n8789), .ZN(n8744) );
  INV_X1 U11207 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8741) );
  NAND2_X1 U11208 ( .A1(n9770), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11209 ( .A1(n9769), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8739) );
  OAI211_X1 U11210 ( .C1(n8741), .C2(n8956), .A(n8740), .B(n8739), .ZN(n8742)
         );
  INV_X1 U11211 ( .A(n8742), .ZN(n8743) );
  NAND2_X1 U11212 ( .A1(n12961), .A2(n13219), .ZN(n8746) );
  XNOR2_X1 U11213 ( .A(n8746), .B(n8745), .ZN(n8747) );
  INV_X1 U11214 ( .A(n8782), .ZN(n8781) );
  NAND2_X1 U11215 ( .A1(n8755), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8750) );
  MUX2_X1 U11216 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8750), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8751) );
  INV_X1 U11217 ( .A(n8777), .ZN(n13392) );
  INV_X1 U11218 ( .A(n8752), .ZN(n8753) );
  NAND2_X1 U11219 ( .A1(n8753), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8754) );
  MUX2_X1 U11220 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8754), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8756) );
  INV_X1 U11221 ( .A(P2_B_REG_SCAN_IN), .ZN(n8951) );
  XNOR2_X1 U11222 ( .A(n11738), .B(n8951), .ZN(n8757) );
  NAND2_X1 U11223 ( .A1(n13392), .A2(n8757), .ZN(n8760) );
  INV_X1 U11224 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8761) );
  NAND2_X1 U11225 ( .A1(n15051), .A2(n8761), .ZN(n8763) );
  OR2_X1 U11226 ( .A1(n8777), .A2(n13387), .ZN(n8762) );
  NAND2_X1 U11227 ( .A1(n8763), .A2(n8762), .ZN(n15087) );
  INV_X1 U11228 ( .A(n15087), .ZN(n8891) );
  INV_X1 U11229 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U11230 ( .A1(n15051), .A2(n8764), .ZN(n8766) );
  NOR4_X1 U11231 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n8775) );
  INV_X1 U11232 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n15058) );
  INV_X1 U11233 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n15064) );
  INV_X1 U11234 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n15052) );
  INV_X1 U11235 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n15082) );
  NAND4_X1 U11236 ( .A1(n15058), .A2(n15064), .A3(n15052), .A4(n15082), .ZN(
        n8772) );
  NOR4_X1 U11237 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_18__SCAN_IN), .ZN(n8770) );
  NOR4_X1 U11238 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n8769) );
  NOR4_X1 U11239 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_30__SCAN_IN), .ZN(n8768) );
  NOR4_X1 U11240 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8767) );
  NAND4_X1 U11241 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n8771)
         );
  NOR4_X1 U11242 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        n8772), .A4(n8771), .ZN(n8774) );
  NOR4_X1 U11243 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n8773) );
  NAND3_X1 U11244 ( .A1(n8775), .A2(n8774), .A3(n8773), .ZN(n8776) );
  NAND2_X1 U11245 ( .A1(n15051), .A2(n8776), .ZN(n8890) );
  NAND3_X1 U11246 ( .A1(n8891), .A2(n15084), .A3(n8890), .ZN(n8800) );
  NAND3_X1 U11247 ( .A1(n13387), .A2(n11738), .A3(n8777), .ZN(n9858) );
  NAND2_X1 U11248 ( .A1(n8778), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8780) );
  INV_X1 U11249 ( .A(n15088), .ZN(n15086) );
  OR2_X1 U11250 ( .A1(n8800), .A2(n15086), .ZN(n8796) );
  NOR2_X1 U11251 ( .A1(n8796), .A2(n10055), .ZN(n10169) );
  NAND2_X1 U11252 ( .A1(n6555), .A2(n13047), .ZN(n9850) );
  NAND2_X1 U11253 ( .A1(n8781), .A2(n12946), .ZN(n8807) );
  INV_X1 U11254 ( .A(n9774), .ZN(n15045) );
  INV_X1 U11255 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8787) );
  NAND2_X1 U11256 ( .A1(n9769), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8786) );
  NAND2_X1 U11257 ( .A1(n9770), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8785) );
  OAI211_X1 U11258 ( .C1(n8956), .C2(n8787), .A(n8786), .B(n8785), .ZN(n8788)
         );
  AOI21_X1 U11259 ( .B1(n8898), .B2(n8789), .A(n8788), .ZN(n9778) );
  NAND2_X1 U11260 ( .A1(n8790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8950) );
  NAND2_X1 U11261 ( .A1(n8950), .A2(n8949), .ZN(n8791) );
  NAND2_X1 U11262 ( .A1(n8791), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8792) );
  XNOR2_X1 U11263 ( .A(n8792), .B(P2_IR_REG_28__SCAN_IN), .ZN(n10067) );
  INV_X1 U11264 ( .A(n10067), .ZN(n8793) );
  OR2_X1 U11265 ( .A1(n9778), .A2(n12886), .ZN(n8795) );
  NAND2_X1 U11266 ( .A1(n12962), .A2(n12932), .ZN(n8794) );
  INV_X1 U11267 ( .A(n8796), .ZN(n8798) );
  INV_X1 U11268 ( .A(n9850), .ZN(n8797) );
  NAND2_X1 U11269 ( .A1(n8798), .A2(n8797), .ZN(n12937) );
  INV_X1 U11270 ( .A(n8799), .ZN(n10310) );
  NAND2_X1 U11271 ( .A1(n8800), .A2(n10310), .ZN(n8801) );
  NAND2_X1 U11272 ( .A1(n10055), .A2(n9850), .ZN(n8889) );
  NAND2_X1 U11273 ( .A1(n8801), .A2(n8889), .ZN(n10166) );
  INV_X1 U11274 ( .A(n8802), .ZN(n8803) );
  AND2_X1 U11275 ( .A1(n8804), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12935) );
  AOI22_X1 U11276 ( .A1(n13072), .A2(n12935), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8805) );
  OAI21_X1 U11277 ( .B1(n13065), .B2(n12937), .A(n8805), .ZN(n8806) );
  NAND2_X1 U11278 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13383), .ZN(n8809) );
  INV_X1 U11279 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U11280 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n11822), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n14450), .ZN(n12022) );
  XNOR2_X1 U11281 ( .A(n12021), .B(n12022), .ZN(n12770) );
  NAND2_X1 U11282 ( .A1(n12770), .A2(n12027), .ZN(n8811) );
  INV_X1 U11283 ( .A(SI_29_), .ZN(n13569) );
  OR2_X1 U11284 ( .A1(n12033), .A2(n13569), .ZN(n8810) );
  NAND2_X1 U11285 ( .A1(n8811), .A2(n8810), .ZN(n8822) );
  OR2_X1 U11286 ( .A1(n8822), .A2(n8812), .ZN(n12218) );
  NAND2_X1 U11287 ( .A1(n8822), .A2(n8812), .ZN(n12226) );
  INV_X1 U11288 ( .A(n12208), .ZN(n12212) );
  XOR2_X1 U11289 ( .A(n12217), .B(n12036), .Z(n12401) );
  INV_X1 U11290 ( .A(P3_B_REG_SCAN_IN), .ZN(n8815) );
  OR2_X1 U11291 ( .A1(n11819), .A2(n8815), .ZN(n8816) );
  NAND2_X1 U11292 ( .A1(n15319), .A2(n8816), .ZN(n14615) );
  NAND2_X1 U11293 ( .A1(n7980), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8819) );
  NAND2_X1 U11294 ( .A1(n10733), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8818) );
  NAND2_X1 U11295 ( .A1(n10734), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8817) );
  AND3_X1 U11296 ( .A1(n8819), .A2(n8818), .A3(n8817), .ZN(n8820) );
  OAI22_X1 U11297 ( .A1(n12417), .A2(n15340), .B1(n14615), .B2(n12037), .ZN(
        n8821) );
  AOI21_X1 U11298 ( .B1(n12401), .B2(n14640), .A(n12397), .ZN(n8837) );
  NAND2_X1 U11299 ( .A1(n8822), .A2(n8823), .ZN(n8825) );
  NAND2_X1 U11300 ( .A1(n15412), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8824) );
  OAI21_X1 U11301 ( .B1(n8837), .B2(n15412), .A(n7432), .ZN(P3_U3456) );
  AND2_X1 U11302 ( .A1(n8826), .A2(n10574), .ZN(n8828) );
  NAND2_X1 U11303 ( .A1(n12227), .A2(n10815), .ZN(n10746) );
  NAND2_X1 U11304 ( .A1(n12219), .A2(n8830), .ZN(n10742) );
  AND2_X1 U11305 ( .A1(n10746), .A2(n10742), .ZN(n8834) );
  OAI22_X1 U11306 ( .A1(n15406), .A2(n10816), .B1(n12375), .B2(n10965), .ZN(
        n8831) );
  AOI21_X1 U11307 ( .B1(n8831), .B2(n10815), .A(n12227), .ZN(n8833) );
  MUX2_X1 U11308 ( .A(n8834), .B(n8833), .S(n8832), .Z(n8835) );
  OR2_X1 U11309 ( .A1(n8837), .A2(n8836), .ZN(n8840) );
  NAND2_X1 U11310 ( .A1(n8822), .A2(n8838), .ZN(n8839) );
  NAND2_X1 U11311 ( .A1(n8840), .A2(n7426), .ZN(P3_U3488) );
  NAND2_X1 U11312 ( .A1(n12988), .A2(n8841), .ZN(n8843) );
  NAND2_X1 U11313 ( .A1(n9597), .A2(n10167), .ZN(n10298) );
  NAND2_X1 U11314 ( .A1(n10303), .A2(n10298), .ZN(n10297) );
  OR2_X1 U11315 ( .A1(n12988), .A2(n10299), .ZN(n8844) );
  NAND2_X1 U11316 ( .A1(n10297), .A2(n8844), .ZN(n10327) );
  NAND2_X1 U11317 ( .A1(n12986), .A2(n10331), .ZN(n8845) );
  NAND2_X1 U11318 ( .A1(n8903), .A2(n8845), .ZN(n10326) );
  OR2_X1 U11319 ( .A1(n12986), .A2(n10756), .ZN(n8846) );
  NAND2_X1 U11320 ( .A1(n10325), .A2(n8846), .ZN(n10393) );
  OR2_X1 U11321 ( .A1(n10433), .A2(n12985), .ZN(n8847) );
  INV_X1 U11322 ( .A(n12984), .ZN(n10470) );
  OR2_X1 U11323 ( .A1(n10417), .A2(n12984), .ZN(n8848) );
  OAI21_X1 U11324 ( .B1(n10636), .B2(n10481), .A(n15098), .ZN(n8850) );
  NAND2_X1 U11325 ( .A1(n10636), .A2(n10481), .ZN(n8849) );
  NAND2_X1 U11326 ( .A1(n8850), .A2(n8849), .ZN(n13256) );
  XNOR2_X1 U11327 ( .A(n15106), .B(n12982), .ZN(n13255) );
  INV_X1 U11328 ( .A(n13255), .ZN(n8851) );
  NAND2_X1 U11329 ( .A1(n15106), .A2(n12982), .ZN(n8852) );
  XNOR2_X1 U11330 ( .A(n10632), .B(n12981), .ZN(n9815) );
  NAND2_X1 U11331 ( .A1(n10632), .A2(n12981), .ZN(n8853) );
  XNOR2_X1 U11332 ( .A(n15116), .B(n12980), .ZN(n10767) );
  INV_X1 U11333 ( .A(n10767), .ZN(n10771) );
  NAND2_X1 U11334 ( .A1(n10772), .A2(n10771), .ZN(n10770) );
  NAND2_X1 U11335 ( .A1(n15116), .A2(n12980), .ZN(n8854) );
  NAND2_X1 U11336 ( .A1(n10770), .A2(n8854), .ZN(n10852) );
  INV_X1 U11337 ( .A(n12979), .ZN(n10837) );
  XNOR2_X1 U11338 ( .A(n15126), .B(n10837), .ZN(n10851) );
  NAND2_X1 U11339 ( .A1(n10852), .A2(n10851), .ZN(n10850) );
  NAND2_X1 U11340 ( .A1(n15126), .A2(n12979), .ZN(n8855) );
  XNOR2_X1 U11341 ( .A(n15136), .B(n12978), .ZN(n9818) );
  NAND2_X1 U11342 ( .A1(n15136), .A2(n12978), .ZN(n8856) );
  XNOR2_X1 U11343 ( .A(n15028), .B(n12977), .ZN(n15016) );
  INV_X1 U11344 ( .A(n15016), .ZN(n15032) );
  NAND2_X1 U11345 ( .A1(n15028), .A2(n12977), .ZN(n8857) );
  NAND2_X1 U11346 ( .A1(n15031), .A2(n8857), .ZN(n11191) );
  OR2_X1 U11347 ( .A1(n13348), .A2(n12976), .ZN(n8858) );
  NAND2_X1 U11348 ( .A1(n13348), .A2(n12976), .ZN(n8859) );
  NAND2_X1 U11349 ( .A1(n14650), .A2(n12975), .ZN(n8860) );
  OR2_X1 U11350 ( .A1(n13344), .A2(n12974), .ZN(n8861) );
  INV_X1 U11351 ( .A(n12973), .ZN(n8922) );
  XNOR2_X1 U11352 ( .A(n12955), .B(n8922), .ZN(n11475) );
  NOR2_X1 U11353 ( .A1(n12955), .A2(n12973), .ZN(n8863) );
  NAND2_X1 U11354 ( .A1(n13339), .A2(n12972), .ZN(n8865) );
  OR2_X1 U11355 ( .A1(n13339), .A2(n12972), .ZN(n8864) );
  NAND2_X1 U11356 ( .A1(n8865), .A2(n8864), .ZN(n9821) );
  NAND2_X1 U11357 ( .A1(n13333), .A2(n12971), .ZN(n9810) );
  INV_X1 U11358 ( .A(n9810), .ZN(n8866) );
  INV_X1 U11359 ( .A(n12970), .ZN(n8928) );
  XNOR2_X1 U11360 ( .A(n13328), .B(n8928), .ZN(n13217) );
  OR2_X1 U11361 ( .A1(n13328), .A2(n12970), .ZN(n8867) );
  NAND2_X1 U11362 ( .A1(n13323), .A2(n12969), .ZN(n9808) );
  OR2_X1 U11363 ( .A1(n13323), .A2(n12969), .ZN(n9809) );
  INV_X1 U11364 ( .A(n12967), .ZN(n8935) );
  XNOR2_X1 U11365 ( .A(n13312), .B(n8935), .ZN(n13178) );
  NAND2_X1 U11366 ( .A1(n13312), .A2(n12967), .ZN(n8868) );
  NAND2_X1 U11367 ( .A1(n8869), .A2(n8868), .ZN(n13155) );
  INV_X1 U11368 ( .A(n12966), .ZN(n12817) );
  XNOR2_X1 U11369 ( .A(n13307), .B(n12817), .ZN(n13161) );
  NAND2_X1 U11370 ( .A1(n13155), .A2(n13161), .ZN(n8871) );
  NAND2_X1 U11371 ( .A1(n13307), .A2(n12966), .ZN(n8870) );
  NAND2_X1 U11372 ( .A1(n13297), .A2(n12852), .ZN(n8939) );
  OR2_X1 U11373 ( .A1(n13297), .A2(n12852), .ZN(n8872) );
  NAND2_X1 U11374 ( .A1(n8939), .A2(n8872), .ZN(n13129) );
  NAND2_X1 U11375 ( .A1(n13297), .A2(n12965), .ZN(n8873) );
  NAND2_X1 U11376 ( .A1(n13132), .A2(n8873), .ZN(n13109) );
  OR2_X1 U11377 ( .A1(n13292), .A2(n12964), .ZN(n8874) );
  NAND2_X1 U11378 ( .A1(n13292), .A2(n12964), .ZN(n8875) );
  INV_X1 U11379 ( .A(n12963), .ZN(n12853) );
  INV_X1 U11380 ( .A(n12962), .ZN(n8944) );
  NAND2_X1 U11381 ( .A1(n13280), .A2(n12962), .ZN(n8877) );
  NAND2_X1 U11382 ( .A1(n13274), .A2(n12961), .ZN(n8879) );
  INV_X1 U11383 ( .A(n13063), .ZN(n13068) );
  NAND2_X1 U11384 ( .A1(n13069), .A2(n13068), .ZN(n13067) );
  NAND2_X1 U11385 ( .A1(n13067), .A2(n8879), .ZN(n8887) );
  NAND2_X1 U11386 ( .A1(n8882), .A2(n11820), .ZN(n8883) );
  MUX2_X1 U11387 ( .A(n14450), .B(n11822), .S(n9981), .Z(n9487) );
  XNOR2_X1 U11388 ( .A(n9487), .B(SI_29_), .ZN(n9485) );
  NAND2_X1 U11389 ( .A1(n11821), .A2(n9780), .ZN(n8886) );
  NAND2_X1 U11390 ( .A1(n8694), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8885) );
  NAND3_X1 U11391 ( .A1(n15088), .A2(n8890), .A3(n8889), .ZN(n10312) );
  INV_X1 U11392 ( .A(n10312), .ZN(n8892) );
  NAND3_X1 U11393 ( .A1(n8892), .A2(n8891), .A3(n10313), .ZN(n8893) );
  AND2_X2 U11394 ( .A1(n9847), .A2(n9774), .ZN(n15044) );
  INV_X1 U11395 ( .A(n15044), .ZN(n8895) );
  OR2_X1 U11396 ( .A1(n15038), .A2(n8895), .ZN(n10437) );
  INV_X1 U11397 ( .A(n10437), .ZN(n10651) );
  INV_X1 U11398 ( .A(n13274), .ZN(n13075) );
  INV_X1 U11399 ( .A(n15028), .ZN(n15147) );
  INV_X1 U11400 ( .A(n10632), .ZN(n15112) );
  INV_X1 U11401 ( .A(n10417), .ZN(n10528) );
  NOR2_X1 U11402 ( .A1(n10328), .A2(n10756), .ZN(n10329) );
  AND2_X1 U11403 ( .A1(n10329), .A2(n8896), .ZN(n10415) );
  AND2_X1 U11404 ( .A1(n10528), .A2(n10415), .ZN(n10637) );
  NAND2_X1 U11405 ( .A1(n15098), .A2(n10637), .ZN(n13258) );
  NOR2_X2 U11406 ( .A1(n13258), .A2(n15106), .ZN(n13257) );
  NAND2_X1 U11407 ( .A1(n15147), .A2(n15022), .ZN(n15020) );
  NAND2_X1 U11408 ( .A1(n13229), .A2(n13237), .ZN(n13230) );
  INV_X1 U11409 ( .A(n13312), .ZN(n13177) );
  OR2_X1 U11410 ( .A1(n13307), .A2(n13171), .ZN(n13156) );
  NOR2_X2 U11411 ( .A1(n13292), .A2(n13133), .ZN(n13112) );
  AOI211_X1 U11412 ( .C1(n13270), .C2(n13071), .A(n13219), .B(n13058), .ZN(
        n13269) );
  INV_X1 U11413 ( .A(n15050), .ZN(n13254) );
  AOI22_X1 U11414 ( .A1(n8898), .A2(n13254), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13242), .ZN(n8899) );
  OAI21_X1 U11415 ( .B1(n7202), .B2(n13236), .A(n8899), .ZN(n8900) );
  AOI21_X1 U11416 ( .B1(n13269), .B2(n13259), .A(n8900), .ZN(n8962) );
  INV_X1 U11417 ( .A(n12961), .ZN(n8946) );
  INV_X1 U11418 ( .A(n10302), .ZN(n8901) );
  NAND2_X1 U11419 ( .A1(n10332), .A2(n8903), .ZN(n10397) );
  NAND2_X1 U11420 ( .A1(n10397), .A2(n10396), .ZN(n10395) );
  NAND2_X1 U11421 ( .A1(n7134), .A2(n10433), .ZN(n8904) );
  INV_X1 U11422 ( .A(n10408), .ZN(n10411) );
  NAND2_X1 U11423 ( .A1(n10417), .A2(n10470), .ZN(n8905) );
  NAND2_X1 U11424 ( .A1(n10640), .A2(n10481), .ZN(n8907) );
  OR2_X1 U11425 ( .A1(n10640), .A2(n10481), .ZN(n8906) );
  NAND2_X1 U11426 ( .A1(n8907), .A2(n8906), .ZN(n10635) );
  INV_X1 U11427 ( .A(n10635), .ZN(n10644) );
  NAND2_X1 U11428 ( .A1(n10642), .A2(n8907), .ZN(n13248) );
  INV_X1 U11429 ( .A(n12982), .ZN(n10469) );
  NAND2_X1 U11430 ( .A1(n15106), .A2(n10469), .ZN(n8908) );
  INV_X1 U11431 ( .A(n12981), .ZN(n10708) );
  OR2_X1 U11432 ( .A1(n10632), .A2(n10708), .ZN(n8909) );
  NAND2_X1 U11433 ( .A1(n10632), .A2(n10708), .ZN(n8910) );
  NAND2_X1 U11434 ( .A1(n10766), .A2(n10767), .ZN(n8912) );
  INV_X1 U11435 ( .A(n12980), .ZN(n10997) );
  NAND2_X1 U11436 ( .A1(n15116), .A2(n10997), .ZN(n8911) );
  NAND2_X1 U11437 ( .A1(n8912), .A2(n8911), .ZN(n10846) );
  INV_X1 U11438 ( .A(n10851), .ZN(n8913) );
  NAND2_X1 U11439 ( .A1(n15126), .A2(n10837), .ZN(n8914) );
  INV_X1 U11440 ( .A(n12978), .ZN(n11329) );
  NAND2_X1 U11441 ( .A1(n15015), .A2(n15016), .ZN(n8916) );
  INV_X1 U11442 ( .A(n12977), .ZN(n11354) );
  NAND2_X1 U11443 ( .A1(n15028), .A2(n11354), .ZN(n8915) );
  NAND2_X1 U11444 ( .A1(n8916), .A2(n8915), .ZN(n11197) );
  INV_X1 U11445 ( .A(n11197), .ZN(n8917) );
  INV_X1 U11446 ( .A(n12976), .ZN(n11348) );
  OR2_X1 U11447 ( .A1(n13348), .A2(n11348), .ZN(n8918) );
  INV_X1 U11448 ( .A(n12975), .ZN(n11198) );
  NOR2_X1 U11449 ( .A1(n14650), .A2(n11198), .ZN(n8919) );
  NAND2_X1 U11450 ( .A1(n14650), .A2(n11198), .ZN(n8920) );
  INV_X1 U11451 ( .A(n12974), .ZN(n11349) );
  AND2_X1 U11452 ( .A1(n13344), .A2(n11349), .ZN(n8921) );
  OAI22_X1 U11453 ( .A1(n11373), .A2(n8921), .B1(n11349), .B2(n13344), .ZN(
        n11471) );
  NOR2_X1 U11454 ( .A1(n12955), .A2(n8922), .ZN(n8924) );
  NAND2_X1 U11455 ( .A1(n12955), .A2(n8922), .ZN(n8923) );
  NAND2_X1 U11456 ( .A1(n11537), .A2(n9821), .ZN(n8926) );
  INV_X1 U11457 ( .A(n12972), .ZN(n12874) );
  NAND2_X1 U11458 ( .A1(n13339), .A2(n12874), .ZN(n8925) );
  NAND2_X1 U11459 ( .A1(n13237), .A2(n12971), .ZN(n8927) );
  NOR2_X1 U11460 ( .A1(n13328), .A2(n8928), .ZN(n8930) );
  NAND2_X1 U11461 ( .A1(n13328), .A2(n8928), .ZN(n8929) );
  INV_X1 U11462 ( .A(n12969), .ZN(n12896) );
  AND2_X1 U11463 ( .A1(n13323), .A2(n12896), .ZN(n8931) );
  OR2_X1 U11464 ( .A1(n13323), .A2(n12896), .ZN(n8932) );
  INV_X1 U11465 ( .A(n12968), .ZN(n8933) );
  XNOR2_X1 U11466 ( .A(n13318), .B(n8933), .ZN(n13189) );
  NAND2_X1 U11467 ( .A1(n13318), .A2(n8933), .ZN(n8934) );
  INV_X1 U11468 ( .A(n13162), .ZN(n8937) );
  INV_X1 U11469 ( .A(n13161), .ZN(n8936) );
  OR2_X1 U11470 ( .A1(n13307), .A2(n12817), .ZN(n8938) );
  INV_X1 U11471 ( .A(n13129), .ZN(n13126) );
  INV_X1 U11472 ( .A(n12964), .ZN(n12928) );
  NAND2_X1 U11473 ( .A1(n13292), .A2(n12928), .ZN(n8941) );
  OR2_X1 U11474 ( .A1(n13292), .A2(n12928), .ZN(n8940) );
  NAND2_X1 U11475 ( .A1(n13103), .A2(n12963), .ZN(n8942) );
  NAND2_X1 U11476 ( .A1(n13287), .A2(n12853), .ZN(n8943) );
  AND2_X2 U11477 ( .A1(n8942), .A2(n8943), .ZN(n13105) );
  NAND2_X1 U11478 ( .A1(n13064), .A2(n13063), .ZN(n13062) );
  OAI21_X1 U11479 ( .B1(n8946), .B2(n13274), .A(n13062), .ZN(n8947) );
  XNOR2_X1 U11480 ( .A(n8947), .B(n9806), .ZN(n8959) );
  NAND2_X1 U11481 ( .A1(n9847), .A2(n6554), .ZN(n8948) );
  OAI21_X1 U11482 ( .B1(n11057), .B2(n13047), .A(n8948), .ZN(n10304) );
  XNOR2_X1 U11483 ( .A(n8950), .B(n8949), .ZN(n13385) );
  NOR2_X1 U11484 ( .A1(n13385), .A2(n8951), .ZN(n8952) );
  NOR2_X1 U11485 ( .A1(n12886), .A2(n8952), .ZN(n13054) );
  INV_X1 U11486 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8955) );
  NAND2_X1 U11487 ( .A1(n9769), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8954) );
  NAND2_X1 U11488 ( .A1(n9770), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8953) );
  OAI211_X1 U11489 ( .C1(n8956), .C2(n8955), .A(n8954), .B(n8953), .ZN(n12959)
         );
  AOI21_X2 U11490 ( .B1(n8959), .B2(n15018), .A(n8958), .ZN(n13272) );
  NAND2_X1 U11491 ( .A1(n8960), .A2(n15048), .ZN(n8961) );
  NAND3_X1 U11492 ( .A1(n7440), .A2(n8962), .A3(n8961), .ZN(P2_U3236) );
  INV_X1 U11493 ( .A(n9065), .ZN(n8970) );
  NOR2_X1 U11494 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .ZN(n8966) );
  NOR2_X2 U11495 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8965) );
  NAND4_X1 U11496 ( .A1(n8966), .A2(n8965), .A3(n9252), .A4(n8964), .ZN(n8968)
         );
  INV_X2 U11497 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n13616) );
  NAND4_X1 U11498 ( .A1(n9232), .A2(n13616), .A3(n9180), .A4(n9133), .ZN(n8967) );
  NOR2_X2 U11499 ( .A1(n8968), .A2(n8967), .ZN(n9264) );
  NOR2_X1 U11500 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n8973) );
  NOR2_X1 U11501 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), 
        .ZN(n8972) );
  NOR2_X1 U11502 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n8971) );
  NOR2_X1 U11503 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), 
        .ZN(n8974) );
  NAND4_X1 U11504 ( .A1(n9566), .A2(n8974), .A3(n9587), .A4(n9584), .ZN(n8975)
         );
  BUF_X2 U11505 ( .A(n8983), .Z(n14449) );
  NAND2_X1 U11506 ( .A1(n8979), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8980) );
  INV_X1 U11507 ( .A(n8981), .ZN(n14442) );
  AND2_X2 U11508 ( .A1(n14449), .A2(n8984), .ZN(n9070) );
  NAND2_X1 U11509 ( .A1(n9070), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n8989) );
  INV_X1 U11510 ( .A(n8983), .ZN(n8985) );
  AND2_X4 U11511 ( .A1(n8985), .A2(n8984), .ZN(n9423) );
  INV_X1 U11512 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10089) );
  OR2_X1 U11513 ( .A1(n9071), .A2(n10089), .ZN(n8986) );
  INV_X1 U11514 ( .A(n8979), .ZN(n8992) );
  NOR2_X1 U11515 ( .A1(n8992), .A2(n8991), .ZN(n8993) );
  NAND2_X1 U11516 ( .A1(n8994), .A2(n8993), .ZN(n9580) );
  INV_X1 U11517 ( .A(n8995), .ZN(n8996) );
  NAND2_X2 U11518 ( .A1(n9580), .A2(n14454), .ZN(n9008) );
  INV_X1 U11519 ( .A(n9990), .ZN(n8997) );
  NAND2_X1 U11520 ( .A1(n9859), .A2(n10862), .ZN(n9535) );
  INV_X1 U11521 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8999) );
  NAND2_X1 U11522 ( .A1(n9070), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9001) );
  NAND2_X1 U11523 ( .A1(n9423), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n9000) );
  INV_X1 U11524 ( .A(SI_0_), .ZN(n9005) );
  INV_X1 U11525 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9004) );
  OAI21_X1 U11526 ( .B1(n9981), .B2(n9005), .A(n9004), .ZN(n9006) );
  AND2_X1 U11527 ( .A1(n9007), .A2(n9006), .ZN(n14460) );
  MUX2_X1 U11528 ( .A(P1_IR_REG_0__SCAN_IN), .B(n14460), .S(n10033), .Z(n10320) );
  NOR2_X2 U11529 ( .A1(n9011), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n9017) );
  NAND2_X1 U11530 ( .A1(n9011), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9012) );
  MUX2_X1 U11531 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9012), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n9014) );
  INV_X1 U11532 ( .A(n9017), .ZN(n9013) );
  NAND2_X1 U11533 ( .A1(n9538), .A2(n9861), .ZN(n9015) );
  NAND2_X1 U11534 ( .A1(n9943), .A2(n10458), .ZN(n9537) );
  INV_X1 U11535 ( .A(n9864), .ZN(n10813) );
  INV_X1 U11536 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9016) );
  AOI21_X1 U11537 ( .B1(n9017), .B2(n9016), .A(n14441), .ZN(n9018) );
  INV_X1 U11538 ( .A(n9020), .ZN(n9021) );
  NAND2_X1 U11539 ( .A1(n9021), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11540 ( .A1(n9026), .A2(n9025), .ZN(n9030) );
  CLKBUF_X2 U11541 ( .A(n9078), .Z(n9393) );
  NAND2_X1 U11542 ( .A1(n9030), .A2(n9029), .ZN(n9045) );
  MUX2_X1 U11543 ( .A(n9027), .B(n13922), .S(n9078), .Z(n9032) );
  NAND2_X1 U11544 ( .A1(n13922), .A2(n9027), .ZN(n9031) );
  NAND2_X1 U11545 ( .A1(n9032), .A2(n9031), .ZN(n9044) );
  NAND2_X1 U11546 ( .A1(n9469), .A2(n9961), .ZN(n9037) );
  INV_X1 U11547 ( .A(n9033), .ZN(n9034) );
  NAND2_X1 U11548 ( .A1(n9034), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9035) );
  XNOR2_X1 U11549 ( .A(n9035), .B(P1_IR_REG_2__SCAN_IN), .ZN(n10249) );
  NAND2_X1 U11550 ( .A1(n9322), .A2(n10249), .ZN(n9036) );
  INV_X2 U11551 ( .A(n14810), .ZN(n9043) );
  INV_X1 U11552 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10088) );
  OR2_X1 U11553 ( .A1(n9071), .A2(n10088), .ZN(n9042) );
  NAND2_X1 U11554 ( .A1(n9423), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n9041) );
  NAND2_X1 U11555 ( .A1(n9070), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9040) );
  INV_X1 U11556 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9038) );
  XNOR2_X2 U11557 ( .A(n9043), .B(n10874), .ZN(n10869) );
  NAND3_X1 U11558 ( .A1(n9045), .A2(n9044), .A3(n10869), .ZN(n9059) );
  NAND2_X1 U11559 ( .A1(n13921), .A2(n9043), .ZN(n9046) );
  MUX2_X1 U11560 ( .A(n9046), .B(n10871), .S(n9078), .Z(n9058) );
  INV_X1 U11561 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9047) );
  OR2_X1 U11562 ( .A1(n9072), .A2(n9047), .ZN(n9052) );
  INV_X1 U11563 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11564 ( .A1(n9423), .A2(n9048), .ZN(n9051) );
  NAND2_X1 U11565 ( .A1(n9070), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9050) );
  INV_X1 U11566 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10876) );
  OR2_X1 U11567 ( .A1(n9071), .A2(n10876), .ZN(n9049) );
  NAND2_X1 U11568 ( .A1(n9053), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9055) );
  INV_X1 U11569 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9054) );
  XNOR2_X1 U11570 ( .A(n9055), .B(n9054), .ZN(n13935) );
  NAND2_X1 U11571 ( .A1(n9985), .A2(n9469), .ZN(n9057) );
  INV_X2 U11572 ( .A(n9184), .ZN(n9520) );
  OAI211_X1 U11573 ( .C1(n10033), .C2(n13935), .A(n9057), .B(n9056), .ZN(n9060) );
  XNOR2_X2 U11574 ( .A(n9060), .B(n13920), .ZN(n10872) );
  NAND3_X1 U11575 ( .A1(n9059), .A2(n9058), .A3(n10872), .ZN(n9064) );
  NAND2_X1 U11576 ( .A1(n9078), .A2(n13920), .ZN(n9062) );
  OR2_X1 U11577 ( .A1(n9078), .A2(n13920), .ZN(n9061) );
  MUX2_X1 U11578 ( .A(n9062), .B(n9061), .S(n14721), .Z(n9063) );
  NAND2_X1 U11579 ( .A1(n9986), .A2(n9469), .ZN(n9069) );
  NAND2_X1 U11580 ( .A1(n9066), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9067) );
  XNOR2_X1 U11581 ( .A(n9067), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U11582 ( .A1(n9520), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6545), .B2(
        n13954), .ZN(n9068) );
  NAND2_X1 U11583 ( .A1(n9327), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9077) );
  INV_X1 U11584 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10091) );
  OR2_X1 U11585 ( .A1(n9475), .A2(n10091), .ZN(n9076) );
  NAND2_X1 U11586 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9085) );
  OAI21_X1 U11587 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n9085), .ZN(n10944) );
  OR2_X1 U11588 ( .A1(n9374), .A2(n10944), .ZN(n9075) );
  INV_X1 U11589 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9073) );
  OR2_X1 U11590 ( .A1(n9477), .A2(n9073), .ZN(n9074) );
  AND4_X2 U11591 ( .A1(n9077), .A2(n9076), .A3(n9075), .A4(n9074), .ZN(n10886)
         );
  MUX2_X1 U11592 ( .A(n10943), .B(n10886), .S(n9025), .Z(n9080) );
  INV_X1 U11593 ( .A(n10886), .ZN(n13919) );
  MUX2_X1 U11594 ( .A(n10942), .B(n13919), .S(n9393), .Z(n9079) );
  NAND2_X1 U11595 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U11596 ( .A1(n9083), .A2(n9082), .ZN(n9100) );
  NAND2_X1 U11597 ( .A1(n9327), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9091) );
  INV_X1 U11598 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n9084) );
  NOR2_X1 U11599 ( .A1(n9085), .A2(n9084), .ZN(n9106) );
  AND2_X1 U11600 ( .A1(n9085), .A2(n9084), .ZN(n9086) );
  NOR2_X1 U11601 ( .A1(n9106), .A2(n9086), .ZN(n10697) );
  NAND2_X1 U11602 ( .A1(n9423), .A2(n10697), .ZN(n9090) );
  INV_X1 U11603 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10920) );
  OR2_X1 U11604 ( .A1(n9475), .A2(n10920), .ZN(n9089) );
  INV_X1 U11605 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n9087) );
  OR2_X1 U11606 ( .A1(n9477), .A2(n9087), .ZN(n9088) );
  NAND4_X1 U11607 ( .A1(n9091), .A2(n9090), .A3(n9089), .A4(n9088), .ZN(n13918) );
  NAND2_X1 U11608 ( .A1(n9987), .A2(n9519), .ZN(n9097) );
  NOR2_X1 U11609 ( .A1(n9066), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n9265) );
  INV_X1 U11610 ( .A(n9265), .ZN(n9092) );
  NAND2_X1 U11611 ( .A1(n9092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9093) );
  MUX2_X1 U11612 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9093), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9095) );
  INV_X1 U11613 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n9094) );
  INV_X1 U11614 ( .A(n9134), .ZN(n9113) );
  AOI22_X1 U11615 ( .A1(n9520), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6545), .B2(
        n10105), .ZN(n9096) );
  NAND2_X1 U11616 ( .A1(n9097), .A2(n9096), .ZN(n10921) );
  MUX2_X1 U11617 ( .A(n13918), .B(n10921), .S(n9025), .Z(n9101) );
  NAND2_X1 U11618 ( .A1(n9100), .A2(n9101), .ZN(n9099) );
  MUX2_X1 U11619 ( .A(n10921), .B(n13918), .S(n9025), .Z(n9098) );
  NAND2_X1 U11620 ( .A1(n9099), .A2(n9098), .ZN(n9105) );
  INV_X1 U11621 ( .A(n9100), .ZN(n9103) );
  INV_X1 U11622 ( .A(n9101), .ZN(n9102) );
  NAND2_X1 U11623 ( .A1(n9103), .A2(n9102), .ZN(n9104) );
  NAND2_X1 U11624 ( .A1(n9105), .A2(n9104), .ZN(n9119) );
  NAND2_X1 U11625 ( .A1(n9327), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U11626 ( .A1(n9106), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9126) );
  OR2_X1 U11627 ( .A1(n9106), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9107) );
  AND2_X1 U11628 ( .A1(n9126), .A2(n9107), .ZN(n14789) );
  NAND2_X1 U11629 ( .A1(n9423), .A2(n14789), .ZN(n9111) );
  INV_X1 U11630 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10093) );
  OR2_X1 U11631 ( .A1(n9475), .A2(n10093), .ZN(n9110) );
  INV_X1 U11632 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9108) );
  OR2_X1 U11633 ( .A1(n9477), .A2(n9108), .ZN(n9109) );
  NAND4_X1 U11634 ( .A1(n9112), .A2(n9111), .A3(n9110), .A4(n9109), .ZN(n13917) );
  NAND2_X1 U11635 ( .A1(n9999), .A2(n9519), .ZN(n9116) );
  NAND2_X1 U11636 ( .A1(n9113), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9114) );
  XNOR2_X1 U11637 ( .A(n9114), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U11638 ( .A1(n9520), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6545), .B2(
        n10107), .ZN(n9115) );
  NAND2_X1 U11639 ( .A1(n9116), .A2(n9115), .ZN(n14788) );
  MUX2_X1 U11640 ( .A(n13917), .B(n14788), .S(n9393), .Z(n9120) );
  NAND2_X1 U11641 ( .A1(n9119), .A2(n9120), .ZN(n9118) );
  MUX2_X1 U11642 ( .A(n13917), .B(n14788), .S(n9025), .Z(n9117) );
  NAND2_X1 U11643 ( .A1(n9118), .A2(n9117), .ZN(n9124) );
  INV_X1 U11644 ( .A(n9119), .ZN(n9122) );
  INV_X1 U11645 ( .A(n9120), .ZN(n9121) );
  NAND2_X1 U11646 ( .A1(n9122), .A2(n9121), .ZN(n9123) );
  NAND2_X1 U11647 ( .A1(n9327), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9132) );
  NAND2_X1 U11648 ( .A1(n9126), .A2(n9125), .ZN(n9127) );
  AND2_X1 U11649 ( .A1(n9141), .A2(n9127), .ZN(n9931) );
  NAND2_X1 U11650 ( .A1(n9423), .A2(n9931), .ZN(n9131) );
  INV_X1 U11651 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10904) );
  OR2_X1 U11652 ( .A1(n9475), .A2(n10904), .ZN(n9130) );
  INV_X1 U11653 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9128) );
  OR2_X1 U11654 ( .A1(n9477), .A2(n9128), .ZN(n9129) );
  NAND4_X1 U11655 ( .A1(n9132), .A2(n9131), .A3(n9130), .A4(n9129), .ZN(n14770) );
  NAND2_X1 U11656 ( .A1(n10003), .A2(n9519), .ZN(n9137) );
  NAND2_X1 U11657 ( .A1(n9134), .A2(n9133), .ZN(n9148) );
  NAND2_X1 U11658 ( .A1(n9148), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9135) );
  XNOR2_X1 U11659 ( .A(n9135), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10115) );
  AOI22_X1 U11660 ( .A1(n9520), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6545), .B2(
        n10115), .ZN(n9136) );
  NAND2_X1 U11661 ( .A1(n9137), .A2(n9136), .ZN(n10978) );
  MUX2_X1 U11662 ( .A(n14770), .B(n10978), .S(n9025), .Z(n9139) );
  MUX2_X1 U11663 ( .A(n14770), .B(n10978), .S(n9393), .Z(n9138) );
  NAND2_X1 U11664 ( .A1(n9141), .A2(n9140), .ZN(n9142) );
  NAND2_X1 U11665 ( .A1(n9160), .A2(n9142), .ZN(n14776) );
  OR2_X1 U11666 ( .A1(n9374), .A2(n14776), .ZN(n9147) );
  NAND2_X1 U11667 ( .A1(n9494), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U11668 ( .A1(n9327), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n9145) );
  INV_X1 U11669 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9143) );
  OR2_X1 U11670 ( .A1(n9477), .A2(n9143), .ZN(n9144) );
  NAND4_X1 U11671 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), .ZN(n13916) );
  NAND2_X1 U11672 ( .A1(n10015), .A2(n9519), .ZN(n9151) );
  NAND2_X1 U11673 ( .A1(n9168), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9149) );
  XNOR2_X1 U11674 ( .A(n9149), .B(P1_IR_REG_8__SCAN_IN), .ZN(n10287) );
  AOI22_X1 U11675 ( .A1(n9520), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6545), .B2(
        n10287), .ZN(n9150) );
  NAND2_X1 U11676 ( .A1(n9151), .A2(n9150), .ZN(n11171) );
  MUX2_X1 U11677 ( .A(n13916), .B(n11171), .S(n9393), .Z(n9155) );
  NAND2_X1 U11678 ( .A1(n9154), .A2(n9155), .ZN(n9153) );
  MUX2_X1 U11679 ( .A(n13916), .B(n11171), .S(n9025), .Z(n9152) );
  NAND2_X1 U11680 ( .A1(n9153), .A2(n9152), .ZN(n9159) );
  INV_X1 U11681 ( .A(n9154), .ZN(n9157) );
  INV_X1 U11682 ( .A(n9155), .ZN(n9156) );
  NAND2_X1 U11683 ( .A1(n9157), .A2(n9156), .ZN(n9158) );
  NAND2_X1 U11684 ( .A1(n9327), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n9167) );
  AND2_X1 U11685 ( .A1(n9160), .A2(n13578), .ZN(n9161) );
  NOR2_X1 U11686 ( .A1(n9198), .A2(n9161), .ZN(n11216) );
  NAND2_X1 U11687 ( .A1(n9423), .A2(n11216), .ZN(n9166) );
  INV_X1 U11688 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9162) );
  OR2_X1 U11689 ( .A1(n9475), .A2(n9162), .ZN(n9165) );
  INV_X1 U11690 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9163) );
  OR2_X1 U11691 ( .A1(n9477), .A2(n9163), .ZN(n9164) );
  NAND4_X1 U11692 ( .A1(n9167), .A2(n9166), .A3(n9165), .A4(n9164), .ZN(n14768) );
  NAND2_X1 U11693 ( .A1(n10019), .A2(n9519), .ZN(n9171) );
  NOR2_X1 U11694 ( .A1(n9168), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9207) );
  INV_X1 U11695 ( .A(n9207), .ZN(n9169) );
  NAND2_X1 U11696 ( .A1(n9169), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9181) );
  XNOR2_X1 U11697 ( .A(n9181), .B(P1_IR_REG_9__SCAN_IN), .ZN(n10288) );
  AOI22_X1 U11698 ( .A1(n9520), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6545), .B2(
        n10288), .ZN(n9170) );
  NAND2_X1 U11699 ( .A1(n9171), .A2(n9170), .ZN(n11206) );
  MUX2_X1 U11700 ( .A(n14768), .B(n11206), .S(n9025), .Z(n9173) );
  MUX2_X1 U11701 ( .A(n14768), .B(n11206), .S(n9500), .Z(n9172) );
  NAND2_X1 U11702 ( .A1(n9327), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9179) );
  INV_X1 U11703 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9174) );
  XNOR2_X1 U11704 ( .A(n9198), .B(n9174), .ZN(n11262) );
  NAND2_X1 U11705 ( .A1(n9423), .A2(n11262), .ZN(n9178) );
  INV_X1 U11706 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9175) );
  OR2_X1 U11707 ( .A1(n9477), .A2(n9175), .ZN(n9177) );
  INV_X1 U11708 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10376) );
  OR2_X1 U11709 ( .A1(n9475), .A2(n10376), .ZN(n9176) );
  NAND4_X1 U11710 ( .A1(n9179), .A2(n9178), .A3(n9177), .A4(n9176), .ZN(n13915) );
  NAND2_X1 U11711 ( .A1(n10023), .A2(n9519), .ZN(n9186) );
  NAND2_X1 U11712 ( .A1(n9181), .A2(n9180), .ZN(n9182) );
  NAND2_X1 U11713 ( .A1(n9182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9183) );
  XNOR2_X1 U11714 ( .A(n9183), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U11715 ( .A1(n10377), .A2(n6545), .B1(n9520), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11716 ( .A1(n9186), .A2(n9185), .ZN(n14917) );
  MUX2_X1 U11717 ( .A(n13915), .B(n14917), .S(n9500), .Z(n9190) );
  NAND2_X1 U11718 ( .A1(n9189), .A2(n9190), .ZN(n9188) );
  MUX2_X1 U11719 ( .A(n13915), .B(n14917), .S(n9025), .Z(n9187) );
  NAND2_X1 U11720 ( .A1(n9188), .A2(n9187), .ZN(n9194) );
  INV_X1 U11721 ( .A(n9189), .ZN(n9192) );
  INV_X1 U11722 ( .A(n9190), .ZN(n9191) );
  NAND2_X1 U11723 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  NAND2_X1 U11724 ( .A1(n9327), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9205) );
  NAND2_X1 U11725 ( .A1(n9198), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9196) );
  INV_X1 U11726 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U11727 ( .A1(n9196), .A2(n9195), .ZN(n9199) );
  AND2_X1 U11728 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n9197) );
  NAND2_X1 U11729 ( .A1(n9198), .A2(n9197), .ZN(n9214) );
  AND2_X1 U11730 ( .A1(n9199), .A2(n9214), .ZN(n11511) );
  NAND2_X1 U11731 ( .A1(n9423), .A2(n11511), .ZN(n9204) );
  INV_X1 U11732 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n9200) );
  OR2_X1 U11733 ( .A1(n9477), .A2(n9200), .ZN(n9203) );
  INV_X1 U11734 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9201) );
  OR2_X1 U11735 ( .A1(n9475), .A2(n9201), .ZN(n9202) );
  NAND4_X1 U11736 ( .A1(n9205), .A2(n9204), .A3(n9203), .A4(n9202), .ZN(n13914) );
  NAND2_X1 U11737 ( .A1(n10050), .A2(n9519), .ZN(n9210) );
  NOR2_X1 U11738 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n9206) );
  NAND2_X1 U11739 ( .A1(n9207), .A2(n9206), .ZN(n9222) );
  NAND2_X1 U11740 ( .A1(n9222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9208) );
  XNOR2_X1 U11741 ( .A(n9208), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10562) );
  AOI22_X1 U11742 ( .A1(n10562), .A2(n9322), .B1(n9520), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n9209) );
  MUX2_X1 U11743 ( .A(n13914), .B(n11494), .S(n9025), .Z(n9212) );
  MUX2_X1 U11744 ( .A(n13914), .B(n11494), .S(n9500), .Z(n9211) );
  NAND2_X1 U11745 ( .A1(n9327), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U11746 ( .A1(n9214), .A2(n13533), .ZN(n9215) );
  AND2_X1 U11747 ( .A1(n9245), .A2(n9215), .ZN(n11613) );
  NAND2_X1 U11748 ( .A1(n9423), .A2(n11613), .ZN(n9220) );
  INV_X1 U11749 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n9216) );
  OR2_X1 U11750 ( .A1(n9477), .A2(n9216), .ZN(n9219) );
  INV_X1 U11751 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9217) );
  OR2_X1 U11752 ( .A1(n9475), .A2(n9217), .ZN(n9218) );
  NAND4_X1 U11753 ( .A1(n9221), .A2(n9220), .A3(n9219), .A4(n9218), .ZN(n13913) );
  NAND2_X1 U11754 ( .A1(n10173), .A2(n9469), .ZN(n9225) );
  NAND2_X1 U11755 ( .A1(n9223), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9233) );
  XNOR2_X1 U11756 ( .A(n9233), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14751) );
  AOI22_X1 U11757 ( .A1(n14751), .A2(n6545), .B1(n9520), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9224) );
  MUX2_X1 U11758 ( .A(n13913), .B(n11605), .S(n9500), .Z(n9229) );
  NAND2_X1 U11759 ( .A1(n9228), .A2(n9229), .ZN(n9227) );
  MUX2_X1 U11760 ( .A(n13913), .B(n11605), .S(n9025), .Z(n9226) );
  NAND2_X1 U11761 ( .A1(n9227), .A2(n9226), .ZN(n9263) );
  INV_X1 U11762 ( .A(n9228), .ZN(n9231) );
  INV_X1 U11763 ( .A(n9229), .ZN(n9230) );
  NAND2_X1 U11764 ( .A1(n9231), .A2(n9230), .ZN(n9262) );
  NAND2_X1 U11765 ( .A1(n10385), .A2(n9519), .ZN(n9237) );
  NAND2_X1 U11766 ( .A1(n9233), .A2(n9232), .ZN(n9234) );
  NAND2_X1 U11767 ( .A1(n9234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U11768 ( .A1(n9253), .A2(n9252), .ZN(n9255) );
  NAND2_X1 U11769 ( .A1(n9255), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9235) );
  XNOR2_X1 U11770 ( .A(n9235), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U11771 ( .A1(n11029), .A2(n6545), .B1(n9520), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n9236) );
  INV_X1 U11772 ( .A(n9245), .ZN(n9238) );
  AOI21_X1 U11773 ( .B1(n9238), .B2(P1_REG3_REG_13__SCAN_IN), .A(
        P1_REG3_REG_14__SCAN_IN), .ZN(n9240) );
  NAND2_X1 U11774 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_REG3_REG_14__SCAN_IN), 
        .ZN(n9239) );
  OR2_X1 U11775 ( .A1(n9240), .A2(n9269), .ZN(n14669) );
  OR2_X1 U11776 ( .A1(n9374), .A2(n14669), .ZN(n9244) );
  NAND2_X1 U11777 ( .A1(n9327), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n9243) );
  NAND2_X1 U11778 ( .A1(n8998), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9242) );
  INV_X1 U11779 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11287) );
  OR2_X1 U11780 ( .A1(n9475), .A2(n11287), .ZN(n9241) );
  NAND4_X1 U11781 ( .A1(n9244), .A2(n9243), .A3(n9242), .A4(n9241), .ZN(n13911) );
  XNOR2_X1 U11782 ( .A(n14658), .B(n13911), .ZN(n11583) );
  NAND2_X1 U11783 ( .A1(n9327), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9251) );
  XNOR2_X1 U11784 ( .A(n9245), .B(P1_REG3_REG_13__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U11785 ( .A1(n9423), .A2(n13868), .ZN(n9250) );
  INV_X1 U11786 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9246) );
  OR2_X1 U11787 ( .A1(n9477), .A2(n9246), .ZN(n9249) );
  INV_X1 U11788 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9247) );
  OR2_X1 U11789 ( .A1(n9475), .A2(n9247), .ZN(n9248) );
  NAND4_X1 U11790 ( .A1(n9251), .A2(n9250), .A3(n9249), .A4(n9248), .ZN(n13912) );
  NAND2_X1 U11791 ( .A1(n10226), .A2(n9469), .ZN(n9257) );
  OR2_X1 U11792 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  AOI22_X1 U11793 ( .A1(n10724), .A2(n9322), .B1(n9520), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9256) );
  MUX2_X1 U11794 ( .A(n13912), .B(n13869), .S(n9025), .Z(n9279) );
  NAND2_X1 U11795 ( .A1(n9025), .A2(n13912), .ZN(n9259) );
  NAND2_X1 U11796 ( .A1(n13869), .A2(n9500), .ZN(n9258) );
  NAND3_X1 U11797 ( .A1(n9279), .A2(n9259), .A3(n9258), .ZN(n9260) );
  NAND3_X1 U11798 ( .A1(n9263), .A2(n9262), .A3(n9261), .ZN(n9285) );
  NAND2_X1 U11799 ( .A1(n10420), .A2(n9519), .ZN(n9268) );
  NAND2_X1 U11800 ( .A1(n9265), .A2(n9264), .ZN(n9296) );
  NAND2_X1 U11801 ( .A1(n9296), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9266) );
  XNOR2_X1 U11802 ( .A(n9266), .B(P1_IR_REG_15__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U11803 ( .A1(n9520), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9322), 
        .B2(n11321), .ZN(n9267) );
  NAND2_X1 U11804 ( .A1(n9268), .A2(n9267), .ZN(n13906) );
  NAND2_X1 U11805 ( .A1(n9327), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n9275) );
  INV_X1 U11806 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11593) );
  OR2_X1 U11807 ( .A1(n9475), .A2(n11593), .ZN(n9274) );
  NAND2_X1 U11808 ( .A1(n9269), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9289) );
  OR2_X1 U11809 ( .A1(n9269), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11810 ( .A1(n9289), .A2(n9270), .ZN(n13903) );
  OR2_X1 U11811 ( .A1(n9374), .A2(n13903), .ZN(n9273) );
  INV_X1 U11812 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9271) );
  OR2_X1 U11813 ( .A1(n9477), .A2(n9271), .ZN(n9272) );
  INV_X1 U11814 ( .A(n13911), .ZN(n13864) );
  OR2_X1 U11815 ( .A1(n14658), .A2(n13864), .ZN(n11585) );
  AOI21_X1 U11816 ( .B1(n11620), .B2(n11585), .A(n9500), .ZN(n9278) );
  NAND2_X1 U11817 ( .A1(n13906), .A2(n14661), .ZN(n9534) );
  NAND2_X1 U11818 ( .A1(n14658), .A2(n13864), .ZN(n9276) );
  AOI21_X1 U11819 ( .B1(n9534), .B2(n9276), .A(n9025), .ZN(n9277) );
  NOR2_X1 U11820 ( .A1(n9278), .A2(n9277), .ZN(n9283) );
  INV_X1 U11821 ( .A(n9279), .ZN(n9281) );
  MUX2_X1 U11822 ( .A(n13912), .B(n13869), .S(n9500), .Z(n9280) );
  NAND3_X1 U11823 ( .A1(n11583), .A2(n9281), .A3(n9280), .ZN(n9282) );
  NAND2_X1 U11824 ( .A1(n9285), .A2(n9284), .ZN(n9287) );
  MUX2_X1 U11825 ( .A(n9534), .B(n11620), .S(n9500), .Z(n9286) );
  INV_X1 U11826 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9288) );
  NAND2_X1 U11827 ( .A1(n9289), .A2(n9288), .ZN(n9290) );
  AND2_X1 U11828 ( .A1(n9308), .A2(n9290), .ZN(n13834) );
  NAND2_X1 U11829 ( .A1(n13834), .A2(n9423), .ZN(n9295) );
  NAND2_X1 U11830 ( .A1(n9327), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n9294) );
  INV_X1 U11831 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11324) );
  OR2_X1 U11832 ( .A1(n9475), .A2(n11324), .ZN(n9293) );
  INV_X1 U11833 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9291) );
  OR2_X1 U11834 ( .A1(n9477), .A2(n9291), .ZN(n9292) );
  NAND4_X1 U11835 ( .A1(n9295), .A2(n9294), .A3(n9293), .A4(n9292), .ZN(n14311) );
  NAND2_X1 U11836 ( .A1(n10346), .A2(n9519), .ZN(n9299) );
  OAI21_X1 U11837 ( .B1(n9296), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9297) );
  XNOR2_X1 U11838 ( .A(n9297), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14003) );
  AOI22_X1 U11839 ( .A1(n9520), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n9322), 
        .B2(n14003), .ZN(n9298) );
  MUX2_X1 U11840 ( .A(n14311), .B(n14086), .S(n9025), .Z(n9301) );
  MUX2_X1 U11841 ( .A(n14311), .B(n14086), .S(n9500), .Z(n9300) );
  NAND2_X1 U11842 ( .A1(n9302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9303) );
  XNOR2_X1 U11843 ( .A(n9303), .B(P1_IR_REG_18__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U11844 ( .A1(n9520), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6545), 
        .B2(n14031), .ZN(n9304) );
  NOR2_X1 U11845 ( .A1(n9309), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9305) );
  OR2_X1 U11846 ( .A1(n9325), .A2(n9305), .ZN(n14291) );
  AOI22_X1 U11847 ( .A1(n9327), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n9494), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U11848 ( .A1(n8998), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n9306) );
  OAI211_X1 U11849 ( .C1(n14291), .C2(n9374), .A(n9307), .B(n9306), .ZN(n14313) );
  OR2_X1 U11850 ( .A1(n14398), .A2(n14313), .ZN(n14067) );
  NAND2_X1 U11851 ( .A1(n14398), .A2(n14313), .ZN(n14066) );
  NAND2_X1 U11852 ( .A1(n14067), .A2(n14066), .ZN(n14281) );
  AND2_X1 U11853 ( .A1(n9308), .A2(n13602), .ZN(n9310) );
  OR2_X1 U11854 ( .A1(n9310), .A2(n9309), .ZN(n14314) );
  AOI22_X1 U11855 ( .A1(n9327), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n9494), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n9312) );
  NAND2_X1 U11856 ( .A1(n8998), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n9311) );
  OAI211_X1 U11857 ( .C1(n14314), .C2(n9374), .A(n9312), .B(n9311), .ZN(n14088) );
  NAND2_X1 U11858 ( .A1(n10421), .A2(n9519), .ZN(n9316) );
  NAND2_X1 U11859 ( .A1(n9567), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9314) );
  XNOR2_X1 U11860 ( .A(n9314), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14012) );
  AOI22_X1 U11861 ( .A1(n9520), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n9322), 
        .B2(n14012), .ZN(n9315) );
  MUX2_X1 U11862 ( .A(n14088), .B(n14310), .S(n9500), .Z(n9318) );
  NAND2_X1 U11863 ( .A1(n14310), .A2(n14088), .ZN(n14065) );
  NAND2_X1 U11864 ( .A1(n9318), .A2(n14065), .ZN(n9317) );
  INV_X1 U11865 ( .A(n9318), .ZN(n9319) );
  OR2_X1 U11866 ( .A1(n14310), .A2(n14088), .ZN(n14063) );
  NAND3_X1 U11867 ( .A1(n14281), .A2(n9319), .A3(n14063), .ZN(n9331) );
  NAND2_X1 U11868 ( .A1(n14398), .A2(n9025), .ZN(n9321) );
  OR2_X1 U11869 ( .A1(n14398), .A2(n9025), .ZN(n9320) );
  MUX2_X1 U11870 ( .A(n9321), .B(n9320), .S(n14313), .Z(n9330) );
  NAND2_X1 U11871 ( .A1(n10685), .A2(n9519), .ZN(n9324) );
  AOI22_X1 U11872 ( .A1(n9520), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14039), 
        .B2(n6545), .ZN(n9323) );
  OR2_X1 U11873 ( .A1(n9325), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9326) );
  NAND2_X1 U11874 ( .A1(n9335), .A2(n9326), .ZN(n14272) );
  AOI22_X1 U11875 ( .A1(n9327), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n9494), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n9329) );
  INV_X1 U11876 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n13540) );
  OR2_X1 U11877 ( .A1(n9477), .A2(n13540), .ZN(n9328) );
  OAI211_X1 U11878 ( .C1(n14272), .C2(n9374), .A(n9329), .B(n9328), .ZN(n14290) );
  XNOR2_X1 U11879 ( .A(n14392), .B(n14290), .ZN(n14268) );
  NAND2_X1 U11880 ( .A1(n14290), .A2(n9025), .ZN(n9333) );
  OR2_X1 U11881 ( .A1(n14290), .A2(n9025), .ZN(n9332) );
  MUX2_X1 U11882 ( .A(n9333), .B(n9332), .S(n14392), .Z(n9334) );
  INV_X1 U11883 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n13856) );
  NAND2_X1 U11884 ( .A1(n9335), .A2(n13856), .ZN(n9336) );
  NAND2_X1 U11885 ( .A1(n9350), .A2(n9336), .ZN(n14258) );
  OR2_X1 U11886 ( .A1(n14258), .A2(n9374), .ZN(n9342) );
  INV_X1 U11887 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9339) );
  NAND2_X1 U11888 ( .A1(n9494), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9338) );
  NAND2_X1 U11889 ( .A1(n8998), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9337) );
  OAI211_X1 U11890 ( .C1(n9213), .C2(n9339), .A(n9338), .B(n9337), .ZN(n9340)
         );
  INV_X1 U11891 ( .A(n9340), .ZN(n9341) );
  OR2_X1 U11892 ( .A1(n10683), .A2(n9417), .ZN(n9344) );
  NAND2_X1 U11893 ( .A1(n9520), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9343) );
  MUX2_X1 U11894 ( .A(n14239), .B(n14261), .S(n9025), .Z(n9346) );
  MUX2_X1 U11895 ( .A(n14094), .B(n14386), .S(n9393), .Z(n9345) );
  OAI21_X1 U11896 ( .B1(n9347), .B2(n9346), .A(n9345), .ZN(n9349) );
  NAND2_X1 U11897 ( .A1(n9347), .A2(n9346), .ZN(n9348) );
  NAND2_X1 U11898 ( .A1(n9350), .A2(n13812), .ZN(n9351) );
  NAND2_X1 U11899 ( .A1(n9360), .A2(n9351), .ZN(n14242) );
  INV_X1 U11900 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U11901 ( .A1(n9494), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U11902 ( .A1(n9327), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n9352) );
  OAI211_X1 U11903 ( .C1(n13517), .C2(n9477), .A(n9353), .B(n9352), .ZN(n9354)
         );
  INV_X1 U11904 ( .A(n9354), .ZN(n9355) );
  OR2_X1 U11905 ( .A1(n10812), .A2(n9417), .ZN(n9357) );
  NAND2_X1 U11906 ( .A1(n9520), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n9356) );
  MUX2_X1 U11907 ( .A(n14252), .B(n14381), .S(n9393), .Z(n9359) );
  MUX2_X1 U11908 ( .A(n14252), .B(n14381), .S(n9025), .Z(n9358) );
  INV_X1 U11909 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13877) );
  AOI21_X1 U11910 ( .B1(n9360), .B2(n13877), .A(n9373), .ZN(n14229) );
  NAND2_X1 U11911 ( .A1(n14229), .A2(n9423), .ZN(n9366) );
  INV_X1 U11912 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U11913 ( .A1(n9494), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U11914 ( .A1(n8998), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9361) );
  OAI211_X1 U11915 ( .C1(n9213), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9364)
         );
  INV_X1 U11916 ( .A(n9364), .ZN(n9365) );
  NAND2_X1 U11917 ( .A1(n9366), .A2(n9365), .ZN(n14074) );
  OR2_X1 U11918 ( .A1(n9368), .A2(n9367), .ZN(n9369) );
  XNOR2_X1 U11919 ( .A(n9369), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14459) );
  MUX2_X1 U11920 ( .A(n14074), .B(n14375), .S(n9025), .Z(n9371) );
  MUX2_X1 U11921 ( .A(n14074), .B(n14375), .S(n9500), .Z(n9370) );
  INV_X1 U11922 ( .A(n9371), .ZN(n9372) );
  NAND2_X1 U11923 ( .A1(n9373), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9400) );
  OAI21_X1 U11924 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n9373), .A(n9400), .ZN(
        n14213) );
  OR2_X1 U11925 ( .A1(n9374), .A2(n14213), .ZN(n9379) );
  NAND2_X1 U11926 ( .A1(n9327), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n9378) );
  NAND2_X1 U11927 ( .A1(n9494), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9377) );
  INV_X1 U11928 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9375) );
  OR2_X1 U11929 ( .A1(n9477), .A2(n9375), .ZN(n9376) );
  NAND4_X1 U11930 ( .A1(n9379), .A2(n9378), .A3(n9377), .A4(n9376), .ZN(n14077) );
  NAND2_X1 U11931 ( .A1(n11378), .A2(n9469), .ZN(n9381) );
  NAND2_X1 U11932 ( .A1(n9520), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9380) );
  MUX2_X1 U11933 ( .A(n14077), .B(n14369), .S(n9393), .Z(n9384) );
  MUX2_X1 U11934 ( .A(n14077), .B(n14369), .S(n9025), .Z(n9382) );
  NAND2_X1 U11935 ( .A1(n11737), .A2(n9469), .ZN(n9386) );
  NAND2_X1 U11936 ( .A1(n9520), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n9385) );
  NAND2_X1 U11937 ( .A1(n9327), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n9392) );
  XNOR2_X1 U11938 ( .A(P1_REG3_REG_24__SCAN_IN), .B(n9400), .ZN(n14197) );
  NAND2_X1 U11939 ( .A1(n9423), .A2(n14197), .ZN(n9391) );
  INV_X1 U11940 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9387) );
  OR2_X1 U11941 ( .A1(n9477), .A2(n9387), .ZN(n9390) );
  INV_X1 U11942 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9388) );
  OR2_X1 U11943 ( .A1(n9475), .A2(n9388), .ZN(n9389) );
  NAND4_X1 U11944 ( .A1(n9392), .A2(n9391), .A3(n9390), .A4(n9389), .ZN(n14079) );
  MUX2_X1 U11945 ( .A(n14079), .B(n14198), .S(n9393), .Z(n9394) );
  INV_X1 U11946 ( .A(n9396), .ZN(n9399) );
  INV_X1 U11947 ( .A(n9397), .ZN(n9398) );
  NAND2_X1 U11948 ( .A1(n9327), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n9411) );
  INV_X1 U11949 ( .A(n9400), .ZN(n9401) );
  NAND2_X1 U11950 ( .A1(n9402), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n9421) );
  INV_X1 U11951 ( .A(n9402), .ZN(n9404) );
  INV_X1 U11952 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9403) );
  NAND2_X1 U11953 ( .A1(n9404), .A2(n9403), .ZN(n9405) );
  AND2_X1 U11954 ( .A1(n9421), .A2(n9405), .ZN(n13820) );
  NAND2_X1 U11955 ( .A1(n9423), .A2(n13820), .ZN(n9410) );
  INV_X1 U11956 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9406) );
  OR2_X1 U11957 ( .A1(n9475), .A2(n9406), .ZN(n9409) );
  INV_X1 U11958 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9407) );
  OR2_X1 U11959 ( .A1(n9477), .A2(n9407), .ZN(n9408) );
  NAND4_X1 U11960 ( .A1(n9411), .A2(n9410), .A3(n9409), .A4(n9408), .ZN(n14159) );
  NAND2_X1 U11961 ( .A1(n13391), .A2(n9519), .ZN(n9413) );
  NAND2_X1 U11962 ( .A1(n6544), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n9412) );
  MUX2_X1 U11963 ( .A(n14159), .B(n14356), .S(n9500), .Z(n9415) );
  MUX2_X1 U11964 ( .A(n14159), .B(n14356), .S(n9025), .Z(n9414) );
  INV_X1 U11965 ( .A(n9415), .ZN(n9416) );
  NAND2_X1 U11966 ( .A1(n9520), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U11967 ( .A1(n9070), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n9429) );
  INV_X1 U11968 ( .A(n9421), .ZN(n9420) );
  NAND2_X1 U11969 ( .A1(n9420), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n9439) );
  INV_X1 U11970 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13579) );
  NAND2_X1 U11971 ( .A1(n9421), .A2(n13579), .ZN(n9422) );
  AND2_X1 U11972 ( .A1(n9439), .A2(n9422), .ZN(n14168) );
  NAND2_X1 U11973 ( .A1(n9423), .A2(n14168), .ZN(n9428) );
  INV_X1 U11974 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9424) );
  OR2_X1 U11975 ( .A1(n9475), .A2(n9424), .ZN(n9427) );
  INV_X1 U11976 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9425) );
  OR2_X1 U11977 ( .A1(n9477), .A2(n9425), .ZN(n9426) );
  NAND4_X1 U11978 ( .A1(n9429), .A2(n9428), .A3(n9427), .A4(n9426), .ZN(n14101) );
  NAND2_X1 U11979 ( .A1(n9431), .A2(n9430), .ZN(n9437) );
  INV_X1 U11980 ( .A(n9432), .ZN(n9435) );
  INV_X1 U11981 ( .A(n9433), .ZN(n9434) );
  NAND2_X1 U11982 ( .A1(n9435), .A2(n9434), .ZN(n9436) );
  NAND2_X1 U11983 ( .A1(n9437), .A2(n9436), .ZN(n9450) );
  NAND2_X1 U11984 ( .A1(n9327), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n9446) );
  INV_X1 U11985 ( .A(n9439), .ZN(n9438) );
  NAND2_X1 U11986 ( .A1(n9438), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9472) );
  INV_X1 U11987 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13774) );
  NAND2_X1 U11988 ( .A1(n9439), .A2(n13774), .ZN(n9440) );
  NAND2_X1 U11989 ( .A1(n9423), .A2(n14147), .ZN(n9445) );
  INV_X1 U11990 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9441) );
  OR2_X1 U11991 ( .A1(n9475), .A2(n9441), .ZN(n9444) );
  INV_X1 U11992 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9442) );
  OR2_X1 U11993 ( .A1(n9477), .A2(n9442), .ZN(n9443) );
  NAND4_X1 U11994 ( .A1(n9446), .A2(n9445), .A3(n9444), .A4(n9443), .ZN(n14158) );
  NAND2_X1 U11995 ( .A1(n13384), .A2(n9469), .ZN(n9448) );
  NAND2_X1 U11996 ( .A1(n9520), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n9447) );
  MUX2_X1 U11997 ( .A(n14158), .B(n14343), .S(n9500), .Z(n9451) );
  MUX2_X1 U11998 ( .A(n14158), .B(n14343), .S(n9025), .Z(n9449) );
  INV_X1 U11999 ( .A(n9464), .ZN(n9462) );
  NAND2_X1 U12000 ( .A1(n9070), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n9457) );
  XNOR2_X1 U12001 ( .A(n9472), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n14132) );
  NAND2_X1 U12002 ( .A1(n9423), .A2(n14132), .ZN(n9456) );
  INV_X1 U12003 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9452) );
  OR2_X1 U12004 ( .A1(n9475), .A2(n9452), .ZN(n9455) );
  INV_X1 U12005 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9453) );
  OR2_X1 U12006 ( .A1(n9477), .A2(n9453), .ZN(n9454) );
  NAND4_X1 U12007 ( .A1(n9457), .A2(n9456), .A3(n9455), .A4(n9454), .ZN(n14108) );
  NAND2_X1 U12008 ( .A1(n9458), .A2(n9469), .ZN(n9460) );
  NAND2_X1 U12009 ( .A1(n6544), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n9459) );
  NAND2_X2 U12010 ( .A1(n9460), .A2(n9459), .ZN(n14338) );
  MUX2_X1 U12011 ( .A(n14108), .B(n14338), .S(n9025), .Z(n9463) );
  INV_X1 U12012 ( .A(n9463), .ZN(n9461) );
  NAND2_X1 U12013 ( .A1(n9462), .A2(n9461), .ZN(n9468) );
  MUX2_X1 U12014 ( .A(n14338), .B(n14108), .S(n9025), .Z(n9465) );
  NAND2_X1 U12015 ( .A1(n9466), .A2(n9465), .ZN(n9467) );
  NAND2_X1 U12016 ( .A1(n11821), .A2(n9469), .ZN(n9471) );
  NAND2_X1 U12017 ( .A1(n9520), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n9470) );
  NAND2_X1 U12018 ( .A1(n9070), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n9481) );
  INV_X1 U12019 ( .A(n9472), .ZN(n9473) );
  AND2_X1 U12020 ( .A1(n9473), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U12021 ( .A1(n9423), .A2(n14111), .ZN(n9480) );
  INV_X1 U12022 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9474) );
  OR2_X1 U12023 ( .A1(n9475), .A2(n9474), .ZN(n9479) );
  INV_X1 U12024 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9476) );
  OR2_X1 U12025 ( .A1(n9477), .A2(n9476), .ZN(n9478) );
  NAND4_X1 U12026 ( .A1(n9481), .A2(n9480), .A3(n9479), .A4(n9478), .ZN(n14125) );
  INV_X1 U12027 ( .A(n14125), .ZN(n13804) );
  MUX2_X1 U12028 ( .A(n14333), .B(n13804), .S(n9025), .Z(n9483) );
  INV_X1 U12029 ( .A(n14333), .ZN(n9556) );
  MUX2_X1 U12030 ( .A(n14125), .B(n9556), .S(n9025), .Z(n9482) );
  NAND2_X1 U12031 ( .A1(n9487), .A2(n13569), .ZN(n9506) );
  NAND2_X1 U12032 ( .A1(n9518), .A2(n9506), .ZN(n9491) );
  MUX2_X1 U12033 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9981), .Z(n9488) );
  NAND2_X1 U12034 ( .A1(n9488), .A2(SI_30_), .ZN(n9510) );
  INV_X1 U12035 ( .A(n9488), .ZN(n9489) );
  INV_X1 U12036 ( .A(SI_30_), .ZN(n13654) );
  NAND2_X1 U12037 ( .A1(n9489), .A2(n13654), .ZN(n9507) );
  AND2_X1 U12038 ( .A1(n9510), .A2(n9507), .ZN(n9490) );
  NAND2_X1 U12039 ( .A1(n13378), .A2(n9519), .ZN(n9493) );
  NAND2_X1 U12040 ( .A1(n9520), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9492) );
  AOI222_X1 U12041 ( .A1(n9070), .A2(P1_REG1_REG_30__SCAN_IN), .B1(n9494), 
        .B2(P1_REG2_REG_30__SCAN_IN), .C1(n8998), .C2(P1_REG0_REG_30__SCAN_IN), 
        .ZN(n9531) );
  INV_X1 U12042 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9497) );
  NAND2_X1 U12043 ( .A1(n9494), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9496) );
  NAND2_X1 U12044 ( .A1(n8998), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9495) );
  OAI211_X1 U12045 ( .C1(n9213), .C2(n9497), .A(n9496), .B(n9495), .ZN(n14048)
         );
  AOI22_X1 U12046 ( .A1(n9500), .A2(n14048), .B1(n10813), .B2(n9498), .ZN(
        n9499) );
  OAI22_X1 U12047 ( .A1(n14328), .A2(n9500), .B1(n9531), .B2(n9499), .ZN(n9503) );
  NAND2_X1 U12048 ( .A1(n9864), .A2(n9952), .ZN(n9937) );
  INV_X1 U12049 ( .A(n9531), .ZN(n14110) );
  OAI21_X1 U12050 ( .B1(n14048), .B2(n9937), .A(n14110), .ZN(n9501) );
  MUX2_X1 U12051 ( .A(n14328), .B(n9501), .S(n9025), .Z(n9502) );
  NAND2_X1 U12052 ( .A1(n9504), .A2(n9503), .ZN(n9523) );
  MUX2_X1 U12053 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9981), .Z(n9505) );
  INV_X1 U12054 ( .A(SI_31_), .ZN(n12767) );
  XNOR2_X1 U12055 ( .A(n9505), .B(n12767), .ZN(n9509) );
  NAND2_X1 U12056 ( .A1(n9509), .A2(n9510), .ZN(n9517) );
  NAND2_X1 U12057 ( .A1(n9507), .A2(n9506), .ZN(n9513) );
  NOR2_X1 U12058 ( .A1(n9513), .A2(n9509), .ZN(n9508) );
  NAND2_X1 U12059 ( .A1(n9518), .A2(n9508), .ZN(n9516) );
  INV_X1 U12060 ( .A(n9509), .ZN(n9514) );
  INV_X1 U12061 ( .A(n9510), .ZN(n9511) );
  XNOR2_X1 U12062 ( .A(n9514), .B(n9511), .ZN(n9512) );
  OAI21_X1 U12063 ( .B1(n9514), .B2(n9513), .A(n9512), .ZN(n9515) );
  OAI211_X1 U12064 ( .C1(n9518), .C2(n9517), .A(n9516), .B(n9515), .ZN(n13371)
         );
  NAND2_X1 U12065 ( .A1(n13371), .A2(n9519), .ZN(n9522) );
  NAND2_X1 U12066 ( .A1(n9520), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n9521) );
  XOR2_X1 U12067 ( .A(n14048), .B(n14049), .Z(n9558) );
  INV_X1 U12068 ( .A(n14048), .ZN(n9525) );
  AND2_X1 U12069 ( .A1(n14049), .A2(n9525), .ZN(n9527) );
  NOR2_X1 U12070 ( .A1(n14049), .A2(n9525), .ZN(n9526) );
  MUX2_X1 U12071 ( .A(n9527), .B(n9526), .S(n9025), .Z(n9563) );
  OAI21_X1 U12072 ( .B1(n6720), .B2(n9952), .A(n10032), .ZN(n9529) );
  OR2_X1 U12073 ( .A1(n9861), .A2(n10687), .ZN(n9954) );
  NAND2_X1 U12074 ( .A1(n9529), .A2(n9954), .ZN(n9565) );
  XOR2_X1 U12075 ( .A(n9531), .B(n14044), .Z(n9561) );
  OR2_X1 U12076 ( .A1(n14338), .A2(n14108), .ZN(n9532) );
  NAND2_X1 U12077 ( .A1(n14338), .A2(n14108), .ZN(n14081) );
  INV_X1 U12078 ( .A(n14079), .ZN(n14098) );
  XNOR2_X1 U12079 ( .A(n14198), .B(n14098), .ZN(n14193) );
  XNOR2_X1 U12080 ( .A(n14369), .B(n14226), .ZN(n14204) );
  XNOR2_X1 U12081 ( .A(n14231), .B(n14074), .ZN(n14222) );
  NAND2_X1 U12082 ( .A1(n14381), .A2(n14252), .ZN(n9533) );
  NAND2_X1 U12083 ( .A1(n14073), .A2(n9533), .ZN(n14236) );
  NAND2_X1 U12084 ( .A1(n14063), .A2(n14065), .ZN(n14300) );
  NAND2_X1 U12085 ( .A1(n14300), .A2(n11583), .ZN(n9550) );
  NAND2_X1 U12086 ( .A1(n11620), .A2(n9534), .ZN(n11590) );
  INV_X1 U12087 ( .A(n14311), .ZN(n14085) );
  INV_X1 U12088 ( .A(n13912), .ZN(n14662) );
  XNOR2_X1 U12089 ( .A(n13869), .B(n14662), .ZN(n11303) );
  XNOR2_X1 U12090 ( .A(n11605), .B(n13865), .ZN(n11291) );
  INV_X1 U12091 ( .A(n13914), .ZN(n11260) );
  XNOR2_X1 U12092 ( .A(n11494), .B(n11260), .ZN(n11223) );
  XNOR2_X1 U12093 ( .A(n14917), .B(n11509), .ZN(n11163) );
  XNOR2_X1 U12094 ( .A(n11206), .B(n14768), .ZN(n10983) );
  AND2_X1 U12095 ( .A1(n9536), .A2(n9535), .ZN(n10865) );
  AND2_X1 U12096 ( .A1(n9538), .A2(n9537), .ZN(n10319) );
  AND3_X1 U12097 ( .A1(n10865), .A2(n10319), .A3(n10869), .ZN(n9542) );
  INV_X1 U12098 ( .A(n13918), .ZN(n9539) );
  NAND2_X1 U12099 ( .A1(n10921), .A2(n9539), .ZN(n14782) );
  OR2_X1 U12100 ( .A1(n10921), .A2(n9539), .ZN(n9540) );
  NAND2_X1 U12101 ( .A1(n10886), .A2(n10942), .ZN(n10915) );
  NAND2_X1 U12102 ( .A1(n10943), .A2(n13919), .ZN(n9541) );
  AND2_X1 U12103 ( .A1(n10915), .A2(n9541), .ZN(n10948) );
  NAND4_X1 U12104 ( .A1(n9542), .A2(n10893), .A3(n10948), .A4(n10872), .ZN(
        n9545) );
  INV_X1 U12105 ( .A(n13917), .ZN(n9543) );
  NAND2_X1 U12106 ( .A1(n14788), .A2(n9543), .ZN(n10896) );
  OR2_X1 U12107 ( .A1(n14788), .A2(n9543), .ZN(n9544) );
  NOR2_X1 U12108 ( .A1(n9545), .A2(n14783), .ZN(n9546) );
  XNOR2_X1 U12109 ( .A(n11171), .B(n13916), .ZN(n10973) );
  XNOR2_X1 U12110 ( .A(n10978), .B(n14770), .ZN(n10897) );
  NAND4_X1 U12111 ( .A1(n10983), .A2(n9546), .A3(n10973), .A4(n10897), .ZN(
        n9547) );
  OR4_X1 U12112 ( .A1(n11291), .A2(n11223), .A3(n11163), .A4(n9547), .ZN(n9548) );
  OR4_X1 U12113 ( .A1(n11590), .A2(n14083), .A3(n11303), .A4(n9548), .ZN(n9549) );
  NOR2_X1 U12114 ( .A1(n9550), .A2(n9549), .ZN(n9551) );
  XNOR2_X1 U12115 ( .A(n14386), .B(n14094), .ZN(n14262) );
  NAND4_X1 U12116 ( .A1(n14236), .A2(n9551), .A3(n14281), .A4(n14262), .ZN(
        n9552) );
  OR4_X1 U12117 ( .A1(n14204), .A2(n14269), .A3(n14222), .A4(n9552), .ZN(n9553) );
  NOR2_X1 U12118 ( .A1(n14193), .A2(n9553), .ZN(n9554) );
  XNOR2_X1 U12119 ( .A(n14356), .B(n14159), .ZN(n14177) );
  XNOR2_X1 U12120 ( .A(n14347), .B(n14101), .ZN(n14156) );
  INV_X1 U12121 ( .A(n14158), .ZN(n14080) );
  XNOR2_X1 U12122 ( .A(n14343), .B(n14080), .ZN(n14140) );
  NAND2_X1 U12123 ( .A1(n7441), .A2(n9555), .ZN(n9557) );
  XOR2_X1 U12124 ( .A(n14125), .B(n9556), .Z(n14104) );
  NOR2_X1 U12125 ( .A1(n9557), .A2(n14104), .ZN(n9560) );
  NAND3_X1 U12126 ( .A1(n9561), .A2(n9560), .A3(n9559), .ZN(n9562) );
  XOR2_X1 U12127 ( .A(n14039), .B(n9562), .Z(n9574) );
  NAND2_X1 U12128 ( .A1(n10813), .A2(n9952), .ZN(n9564) );
  INV_X1 U12129 ( .A(n9564), .ZN(n9573) );
  INV_X1 U12130 ( .A(n9563), .ZN(n9571) );
  NAND2_X1 U12131 ( .A1(n9565), .A2(n9564), .ZN(n9577) );
  NAND2_X1 U12132 ( .A1(n6675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9569) );
  MUX2_X1 U12133 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9569), .S(
        P1_IR_REG_23__SCAN_IN), .Z(n9570) );
  INV_X4 U12134 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  OAI21_X1 U12135 ( .B1(n9571), .B2(n9577), .A(n11379), .ZN(n9572) );
  INV_X1 U12136 ( .A(n9577), .ZN(n9578) );
  INV_X1 U12137 ( .A(n10032), .ZN(n9579) );
  NAND2_X1 U12138 ( .A1(n10684), .A2(n10687), .ZN(n9901) );
  AND2_X1 U12139 ( .A1(n9579), .A2(n9901), .ZN(n9947) );
  NAND2_X1 U12140 ( .A1(n9581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9585) );
  NAND2_X1 U12141 ( .A1(n9586), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9588) );
  INV_X1 U12142 ( .A(n9856), .ZN(n10009) );
  NOR4_X1 U12143 ( .A1(n9947), .A2(n14288), .A3(n14454), .A4(n10036), .ZN(
        n9590) );
  INV_X1 U12144 ( .A(n11379), .ZN(n10035) );
  OAI21_X1 U12145 ( .B1(n6720), .B2(n10035), .A(P1_B_REG_SCAN_IN), .ZN(n9589)
         );
  OR2_X1 U12146 ( .A1(n9590), .A2(n9589), .ZN(n9591) );
  NAND2_X1 U12147 ( .A1(n11057), .A2(n9844), .ZN(n9592) );
  NOR2_X1 U12148 ( .A1(n9595), .A2(n9594), .ZN(n9596) );
  NAND2_X2 U12149 ( .A1(n15044), .A2(n11057), .ZN(n9784) );
  OAI211_X1 U12150 ( .C1(n15042), .C2(n9845), .A(n9597), .B(n9784), .ZN(n9598)
         );
  NAND2_X1 U12151 ( .A1(n9599), .A2(n9598), .ZN(n9604) );
  NAND2_X1 U12152 ( .A1(n12988), .A2(n9784), .ZN(n9601) );
  NAND2_X1 U12153 ( .A1(n9777), .A2(n10299), .ZN(n9600) );
  NAND2_X1 U12154 ( .A1(n9601), .A2(n9600), .ZN(n9605) );
  NAND2_X1 U12155 ( .A1(n9604), .A2(n9605), .ZN(n9603) );
  MUX2_X1 U12156 ( .A(n12988), .B(n10299), .S(n9784), .Z(n9602) );
  NAND2_X1 U12157 ( .A1(n9603), .A2(n9602), .ZN(n9609) );
  INV_X1 U12158 ( .A(n9604), .ZN(n9607) );
  INV_X1 U12159 ( .A(n9605), .ZN(n9606) );
  NAND2_X1 U12160 ( .A1(n9607), .A2(n9606), .ZN(n9608) );
  MUX2_X1 U12161 ( .A(n10756), .B(n12986), .S(n9784), .Z(n9610) );
  INV_X1 U12162 ( .A(n9611), .ZN(n9612) );
  MUX2_X1 U12163 ( .A(n10433), .B(n12985), .S(n9784), .Z(n9616) );
  NAND2_X1 U12164 ( .A1(n9615), .A2(n9616), .ZN(n9614) );
  INV_X2 U12165 ( .A(n9784), .ZN(n9777) );
  MUX2_X1 U12166 ( .A(n12985), .B(n10433), .S(n9779), .Z(n9613) );
  NAND2_X1 U12167 ( .A1(n9614), .A2(n9613), .ZN(n9620) );
  INV_X1 U12168 ( .A(n9615), .ZN(n9618) );
  INV_X1 U12169 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U12170 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  NAND2_X1 U12171 ( .A1(n9620), .A2(n9619), .ZN(n9623) );
  MUX2_X1 U12172 ( .A(n12984), .B(n10417), .S(n9779), .Z(n9624) );
  NAND2_X1 U12173 ( .A1(n9623), .A2(n9624), .ZN(n9622) );
  INV_X1 U12174 ( .A(n9784), .ZN(n9737) );
  MUX2_X1 U12175 ( .A(n12984), .B(n10417), .S(n9737), .Z(n9621) );
  NAND2_X1 U12176 ( .A1(n9622), .A2(n9621), .ZN(n9628) );
  INV_X1 U12177 ( .A(n9623), .ZN(n9626) );
  INV_X1 U12178 ( .A(n9624), .ZN(n9625) );
  NAND2_X1 U12179 ( .A1(n9626), .A2(n9625), .ZN(n9627) );
  MUX2_X1 U12180 ( .A(n12983), .B(n10640), .S(n9737), .Z(n9630) );
  MUX2_X1 U12181 ( .A(n12983), .B(n10640), .S(n9779), .Z(n9629) );
  MUX2_X1 U12182 ( .A(n12982), .B(n15106), .S(n9779), .Z(n9634) );
  NAND2_X1 U12183 ( .A1(n9633), .A2(n9634), .ZN(n9632) );
  MUX2_X1 U12184 ( .A(n12982), .B(n15106), .S(n9737), .Z(n9631) );
  NAND2_X1 U12185 ( .A1(n9632), .A2(n9631), .ZN(n9638) );
  INV_X1 U12186 ( .A(n9633), .ZN(n9636) );
  INV_X1 U12187 ( .A(n9634), .ZN(n9635) );
  NAND2_X1 U12188 ( .A1(n9636), .A2(n9635), .ZN(n9637) );
  MUX2_X1 U12189 ( .A(n12981), .B(n10632), .S(n9777), .Z(n9640) );
  MUX2_X1 U12190 ( .A(n12981), .B(n10632), .S(n9779), .Z(n9639) );
  INV_X1 U12191 ( .A(n9640), .ZN(n9641) );
  MUX2_X1 U12192 ( .A(n12980), .B(n15116), .S(n9779), .Z(n9645) );
  NAND2_X1 U12193 ( .A1(n9644), .A2(n9645), .ZN(n9643) );
  MUX2_X1 U12194 ( .A(n12980), .B(n15116), .S(n9777), .Z(n9642) );
  NAND2_X1 U12195 ( .A1(n9643), .A2(n9642), .ZN(n9649) );
  INV_X1 U12196 ( .A(n9644), .ZN(n9647) );
  INV_X1 U12197 ( .A(n9645), .ZN(n9646) );
  NAND2_X1 U12198 ( .A1(n9647), .A2(n9646), .ZN(n9648) );
  MUX2_X1 U12199 ( .A(n12979), .B(n15126), .S(n9777), .Z(n9651) );
  MUX2_X1 U12200 ( .A(n12979), .B(n15126), .S(n9779), .Z(n9650) );
  INV_X1 U12201 ( .A(n9651), .ZN(n9652) );
  MUX2_X1 U12202 ( .A(n12978), .B(n15136), .S(n9779), .Z(n9656) );
  NAND2_X1 U12203 ( .A1(n9655), .A2(n9656), .ZN(n9654) );
  MUX2_X1 U12204 ( .A(n12978), .B(n15136), .S(n9777), .Z(n9653) );
  NAND2_X1 U12205 ( .A1(n9654), .A2(n9653), .ZN(n9660) );
  INV_X1 U12206 ( .A(n9655), .ZN(n9658) );
  INV_X1 U12207 ( .A(n9656), .ZN(n9657) );
  NAND2_X1 U12208 ( .A1(n9658), .A2(n9657), .ZN(n9659) );
  MUX2_X1 U12209 ( .A(n12977), .B(n15028), .S(n9777), .Z(n9662) );
  MUX2_X1 U12210 ( .A(n12977), .B(n15028), .S(n9779), .Z(n9661) );
  MUX2_X1 U12211 ( .A(n12976), .B(n13348), .S(n9779), .Z(n9666) );
  NAND2_X1 U12212 ( .A1(n9665), .A2(n9666), .ZN(n9664) );
  MUX2_X1 U12213 ( .A(n12976), .B(n13348), .S(n9737), .Z(n9663) );
  NAND2_X1 U12214 ( .A1(n9664), .A2(n9663), .ZN(n9670) );
  INV_X1 U12215 ( .A(n9665), .ZN(n9668) );
  INV_X1 U12216 ( .A(n9666), .ZN(n9667) );
  NAND2_X1 U12217 ( .A1(n9668), .A2(n9667), .ZN(n9669) );
  MUX2_X1 U12218 ( .A(n12975), .B(n14650), .S(n9737), .Z(n9672) );
  MUX2_X1 U12219 ( .A(n12975), .B(n14650), .S(n9779), .Z(n9671) );
  INV_X1 U12220 ( .A(n9672), .ZN(n9673) );
  MUX2_X1 U12221 ( .A(n12974), .B(n13344), .S(n9779), .Z(n9677) );
  NAND2_X1 U12222 ( .A1(n9676), .A2(n9677), .ZN(n9675) );
  MUX2_X1 U12223 ( .A(n12974), .B(n13344), .S(n9777), .Z(n9674) );
  NAND2_X1 U12224 ( .A1(n9675), .A2(n9674), .ZN(n9681) );
  INV_X1 U12225 ( .A(n9676), .ZN(n9679) );
  INV_X1 U12226 ( .A(n9677), .ZN(n9678) );
  NAND2_X1 U12227 ( .A1(n9679), .A2(n9678), .ZN(n9680) );
  MUX2_X1 U12228 ( .A(n12973), .B(n12955), .S(n9737), .Z(n9684) );
  MUX2_X1 U12229 ( .A(n12973), .B(n12955), .S(n9779), .Z(n9682) );
  MUX2_X1 U12230 ( .A(n12972), .B(n13339), .S(n9779), .Z(n9702) );
  NAND2_X1 U12231 ( .A1(n9702), .A2(n12971), .ZN(n9685) );
  NAND2_X1 U12232 ( .A1(n12874), .A2(n9779), .ZN(n9687) );
  AOI21_X1 U12233 ( .B1(n9685), .B2(n9687), .A(n13237), .ZN(n9692) );
  INV_X1 U12234 ( .A(n12971), .ZN(n9688) );
  NAND2_X1 U12235 ( .A1(n9702), .A2(n9688), .ZN(n9686) );
  OR2_X1 U12236 ( .A1(n13339), .A2(n9784), .ZN(n9694) );
  AOI21_X1 U12237 ( .B1(n9686), .B2(n9694), .A(n13333), .ZN(n9691) );
  NAND2_X1 U12238 ( .A1(n12971), .A2(n9737), .ZN(n9695) );
  OR2_X1 U12239 ( .A1(n13339), .A2(n9695), .ZN(n9690) );
  INV_X1 U12240 ( .A(n9687), .ZN(n9698) );
  NAND2_X1 U12241 ( .A1(n9698), .A2(n9688), .ZN(n9689) );
  NAND2_X1 U12242 ( .A1(n9690), .A2(n9689), .ZN(n9701) );
  OR3_X1 U12243 ( .A1(n9692), .A2(n9691), .A3(n9701), .ZN(n9693) );
  INV_X1 U12244 ( .A(n9694), .ZN(n9697) );
  INV_X1 U12245 ( .A(n9695), .ZN(n9696) );
  AOI21_X1 U12246 ( .B1(n9702), .B2(n9697), .A(n9696), .ZN(n9705) );
  NAND2_X1 U12247 ( .A1(n9702), .A2(n9698), .ZN(n9699) );
  OAI21_X1 U12248 ( .B1(n9777), .B2(n12971), .A(n9699), .ZN(n9700) );
  NAND2_X1 U12249 ( .A1(n9700), .A2(n13333), .ZN(n9704) );
  NAND2_X1 U12250 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  OAI211_X1 U12251 ( .C1(n9705), .C2(n13333), .A(n9704), .B(n9703), .ZN(n9706)
         );
  MUX2_X1 U12252 ( .A(n12970), .B(n13328), .S(n9779), .Z(n9710) );
  NAND2_X1 U12253 ( .A1(n9709), .A2(n9710), .ZN(n9708) );
  MUX2_X1 U12254 ( .A(n12970), .B(n13328), .S(n9737), .Z(n9707) );
  NAND2_X1 U12255 ( .A1(n9708), .A2(n9707), .ZN(n9714) );
  INV_X1 U12256 ( .A(n9709), .ZN(n9712) );
  INV_X1 U12257 ( .A(n9710), .ZN(n9711) );
  NAND2_X1 U12258 ( .A1(n9712), .A2(n9711), .ZN(n9713) );
  MUX2_X1 U12259 ( .A(n12969), .B(n13323), .S(n9777), .Z(n9716) );
  MUX2_X1 U12260 ( .A(n12969), .B(n13323), .S(n9779), .Z(n9715) );
  INV_X1 U12261 ( .A(n9716), .ZN(n9717) );
  MUX2_X1 U12262 ( .A(n12968), .B(n13318), .S(n9779), .Z(n9721) );
  NAND2_X1 U12263 ( .A1(n9720), .A2(n9721), .ZN(n9719) );
  MUX2_X1 U12264 ( .A(n12968), .B(n13318), .S(n9737), .Z(n9718) );
  NAND2_X1 U12265 ( .A1(n9719), .A2(n9718), .ZN(n9725) );
  NAND2_X1 U12266 ( .A1(n9723), .A2(n9722), .ZN(n9724) );
  MUX2_X1 U12267 ( .A(n12967), .B(n13312), .S(n9777), .Z(n9727) );
  MUX2_X1 U12268 ( .A(n12967), .B(n13312), .S(n9779), .Z(n9726) );
  INV_X1 U12269 ( .A(n9727), .ZN(n9728) );
  MUX2_X1 U12270 ( .A(n12966), .B(n13307), .S(n9779), .Z(n9732) );
  NAND2_X1 U12271 ( .A1(n9731), .A2(n9732), .ZN(n9730) );
  MUX2_X1 U12272 ( .A(n12966), .B(n13307), .S(n9737), .Z(n9729) );
  NAND2_X1 U12273 ( .A1(n9730), .A2(n9729), .ZN(n9736) );
  INV_X1 U12274 ( .A(n9731), .ZN(n9734) );
  INV_X1 U12275 ( .A(n9732), .ZN(n9733) );
  NAND2_X1 U12276 ( .A1(n9734), .A2(n9733), .ZN(n9735) );
  MUX2_X1 U12277 ( .A(n12913), .B(n13302), .S(n9737), .Z(n9739) );
  MUX2_X1 U12278 ( .A(n12913), .B(n13302), .S(n9779), .Z(n9738) );
  MUX2_X1 U12279 ( .A(n12965), .B(n13297), .S(n9779), .Z(n9743) );
  NAND2_X1 U12280 ( .A1(n9742), .A2(n9743), .ZN(n9741) );
  MUX2_X1 U12281 ( .A(n13297), .B(n12965), .S(n9779), .Z(n9740) );
  NAND2_X1 U12282 ( .A1(n9741), .A2(n9740), .ZN(n9747) );
  INV_X1 U12283 ( .A(n9742), .ZN(n9745) );
  NAND2_X1 U12284 ( .A1(n9745), .A2(n9744), .ZN(n9746) );
  MUX2_X1 U12285 ( .A(n12964), .B(n13292), .S(n9737), .Z(n9749) );
  MUX2_X1 U12286 ( .A(n12964), .B(n13292), .S(n9779), .Z(n9748) );
  INV_X1 U12287 ( .A(n9749), .ZN(n9750) );
  MUX2_X1 U12288 ( .A(n12963), .B(n13287), .S(n9779), .Z(n9754) );
  NAND2_X1 U12289 ( .A1(n9753), .A2(n9754), .ZN(n9752) );
  MUX2_X1 U12290 ( .A(n13287), .B(n12963), .S(n9779), .Z(n9751) );
  NAND2_X1 U12291 ( .A1(n9752), .A2(n9751), .ZN(n9758) );
  INV_X1 U12292 ( .A(n9753), .ZN(n9756) );
  INV_X1 U12293 ( .A(n9754), .ZN(n9755) );
  NAND2_X1 U12294 ( .A1(n9756), .A2(n9755), .ZN(n9757) );
  NAND2_X1 U12295 ( .A1(n9758), .A2(n9757), .ZN(n9761) );
  MUX2_X1 U12296 ( .A(n12962), .B(n13280), .S(n9777), .Z(n9762) );
  NAND2_X1 U12297 ( .A1(n9761), .A2(n9762), .ZN(n9760) );
  MUX2_X1 U12298 ( .A(n12962), .B(n13280), .S(n9779), .Z(n9759) );
  NAND2_X1 U12299 ( .A1(n9760), .A2(n9759), .ZN(n9766) );
  INV_X1 U12300 ( .A(n9761), .ZN(n9764) );
  INV_X1 U12301 ( .A(n9762), .ZN(n9763) );
  NAND2_X1 U12302 ( .A1(n9764), .A2(n9763), .ZN(n9765) );
  NAND2_X1 U12303 ( .A1(n9766), .A2(n9765), .ZN(n9788) );
  NAND2_X1 U12304 ( .A1(n13378), .A2(n9780), .ZN(n9768) );
  NAND2_X1 U12305 ( .A1(n8694), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n9767) );
  INV_X1 U12306 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9773) );
  NAND2_X1 U12307 ( .A1(n9769), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9772) );
  NAND2_X1 U12308 ( .A1(n9770), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9771) );
  OAI211_X1 U12309 ( .C1(n8956), .C2(n9773), .A(n9772), .B(n9771), .ZN(n13053)
         );
  NAND2_X1 U12310 ( .A1(n13053), .A2(n9779), .ZN(n9801) );
  INV_X1 U12311 ( .A(n11057), .ZN(n9852) );
  NAND2_X1 U12312 ( .A1(n9852), .A2(n9774), .ZN(n9840) );
  NAND4_X1 U12313 ( .A1(n9801), .A2(n9847), .A3(n9850), .A4(n9840), .ZN(n9775)
         );
  AND2_X1 U12314 ( .A1(n9775), .A2(n12959), .ZN(n9776) );
  AOI21_X1 U12315 ( .B1(n13052), .B2(n9777), .A(n9776), .ZN(n9795) );
  INV_X1 U12316 ( .A(n9778), .ZN(n12960) );
  MUX2_X1 U12317 ( .A(n12960), .B(n13270), .S(n9779), .Z(n9790) );
  NAND2_X1 U12318 ( .A1(n13371), .A2(n9780), .ZN(n9782) );
  NAND2_X1 U12319 ( .A1(n8694), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n9781) );
  NAND2_X1 U12320 ( .A1(n9782), .A2(n9781), .ZN(n9800) );
  NAND2_X1 U12321 ( .A1(n9800), .A2(n13053), .ZN(n9783) );
  MUX2_X1 U12322 ( .A(n13274), .B(n12961), .S(n9779), .Z(n9793) );
  MUX2_X1 U12323 ( .A(n12961), .B(n13274), .S(n9784), .Z(n9789) );
  INV_X1 U12324 ( .A(n9789), .ZN(n9785) );
  NAND2_X1 U12325 ( .A1(n9793), .A2(n9785), .ZN(n9786) );
  NAND2_X1 U12326 ( .A1(n9788), .A2(n9787), .ZN(n9799) );
  NAND2_X1 U12327 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  OAI211_X1 U12328 ( .C1(n9785), .C2(n9793), .A(n9792), .B(n9832), .ZN(n9796)
         );
  AOI22_X1 U12329 ( .A1(n9797), .A2(n9796), .B1(n9795), .B2(n9794), .ZN(n9798)
         );
  NAND2_X1 U12330 ( .A1(n9799), .A2(n9798), .ZN(n9805) );
  NAND2_X1 U12331 ( .A1(n9800), .A2(n9737), .ZN(n9802) );
  NAND3_X1 U12332 ( .A1(n9803), .A2(n9802), .A3(n9801), .ZN(n9804) );
  NAND2_X1 U12333 ( .A1(n9805), .A2(n9804), .ZN(n9849) );
  XOR2_X1 U12334 ( .A(n12959), .B(n13052), .Z(n9834) );
  INV_X1 U12335 ( .A(n9806), .ZN(n9831) );
  XNOR2_X1 U12336 ( .A(n13302), .B(n12885), .ZN(n13151) );
  NAND2_X1 U12337 ( .A1(n9811), .A2(n9810), .ZN(n13238) );
  XNOR2_X1 U12338 ( .A(n14650), .B(n11198), .ZN(n11346) );
  XNOR2_X1 U12339 ( .A(n13348), .B(n12976), .ZN(n11196) );
  NOR2_X1 U12340 ( .A1(n15092), .A2(n6556), .ZN(n9813) );
  NAND4_X1 U12341 ( .A1(n9813), .A2(n10334), .A3(n9812), .A4(n10396), .ZN(
        n9814) );
  NOR3_X1 U12342 ( .A1(n10635), .A2(n10408), .A3(n9814), .ZN(n9816) );
  NAND4_X1 U12343 ( .A1(n10767), .A2(n9816), .A3(n9815), .A4(n13255), .ZN(
        n9817) );
  NOR2_X1 U12344 ( .A1(n10851), .A2(n9817), .ZN(n9819) );
  NAND4_X1 U12345 ( .A1(n11196), .A2(n9819), .A3(n15016), .A4(n9818), .ZN(
        n9820) );
  NOR2_X1 U12346 ( .A1(n11346), .A2(n9820), .ZN(n9822) );
  XNOR2_X1 U12347 ( .A(n13344), .B(n12974), .ZN(n11374) );
  NAND4_X1 U12348 ( .A1(n13238), .A2(n9822), .A3(n11374), .A4(n9821), .ZN(
        n9823) );
  OR4_X1 U12349 ( .A1(n13189), .A2(n13217), .A3(n11475), .A4(n9823), .ZN(n9824) );
  OR4_X1 U12350 ( .A1(n13161), .A2(n13178), .A3(n13204), .A4(n9824), .ZN(n9825) );
  NOR3_X1 U12351 ( .A1(n13129), .A2(n13151), .A3(n9825), .ZN(n9826) );
  NAND3_X1 U12352 ( .A1(n9832), .A2(n9831), .A3(n9830), .ZN(n9833) );
  NOR2_X1 U12353 ( .A1(n9834), .A2(n9833), .ZN(n9837) );
  AOI21_X1 U12354 ( .B1(n9837), .B2(n9844), .A(n9847), .ZN(n9838) );
  INV_X1 U12355 ( .A(n9838), .ZN(n9835) );
  INV_X1 U12356 ( .A(n9837), .ZN(n9839) );
  AOI21_X1 U12357 ( .B1(n13047), .B2(n9839), .A(n9835), .ZN(n9843) );
  INV_X1 U12358 ( .A(n9840), .ZN(n9842) );
  NOR3_X1 U12359 ( .A1(n10810), .A2(n13047), .A3(n6555), .ZN(n9841) );
  OAI21_X1 U12360 ( .B1(n9852), .B2(n9845), .A(n9844), .ZN(n9846) );
  OAI21_X1 U12361 ( .B1(n9847), .B2(n6556), .A(n9846), .ZN(n9848) );
  NOR2_X1 U12362 ( .A1(n10054), .A2(P2_U3088), .ZN(n11381) );
  NOR4_X1 U12363 ( .A1(n15086), .A2(n12884), .A3(n13385), .A4(n9850), .ZN(
        n9854) );
  INV_X1 U12364 ( .A(n11381), .ZN(n9851) );
  OAI21_X1 U12365 ( .B1(n9852), .B2(n9851), .A(P2_B_REG_SCAN_IN), .ZN(n9853)
         );
  INV_X1 U12366 ( .A(n10054), .ZN(n9857) );
  NAND2_X2 U12367 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10056), .ZN(n12987) );
  NAND2_X1 U12368 ( .A1(n9862), .A2(n9861), .ZN(n13679) );
  OAI21_X1 U12369 ( .B1(n10862), .B2(n13729), .A(n9865), .ZN(n9871) );
  OAI222_X1 U12370 ( .A1(n13729), .A2(n10458), .B1(n13728), .B2(n9939), .C1(
        n9866), .C2(n7268), .ZN(n10233) );
  INV_X1 U12371 ( .A(n9866), .ZN(n9927) );
  AOI22_X1 U12372 ( .A1(n13798), .A2(n10320), .B1(n9927), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9867) );
  INV_X1 U12373 ( .A(n10232), .ZN(n9870) );
  NAND2_X1 U12374 ( .A1(n10234), .A2(n6549), .ZN(n9869) );
  NAND2_X1 U12375 ( .A1(n9892), .A2(n13921), .ZN(n9873) );
  NAND2_X1 U12376 ( .A1(n9891), .A2(n14810), .ZN(n9872) );
  NAND2_X1 U12377 ( .A1(n9873), .A2(n9872), .ZN(n9876) );
  XOR2_X1 U12378 ( .A(n9876), .B(n9875), .Z(n10460) );
  INV_X1 U12379 ( .A(n9875), .ZN(n9878) );
  INV_X1 U12380 ( .A(n9876), .ZN(n9877) );
  AOI21_X1 U12381 ( .B1(n10459), .B2(n10460), .A(n7421), .ZN(n14729) );
  AOI22_X1 U12382 ( .A1(n9892), .A2(n13920), .B1(n9891), .B2(n14721), .ZN(
        n9881) );
  AOI22_X1 U12383 ( .A1(n13920), .A2(n9891), .B1(n14721), .B2(n13798), .ZN(
        n9879) );
  XNOR2_X1 U12384 ( .A(n9879), .B(n6549), .ZN(n9880) );
  XOR2_X1 U12385 ( .A(n9881), .B(n9880), .Z(n14728) );
  NAND2_X1 U12386 ( .A1(n14729), .A2(n14728), .ZN(n14727) );
  INV_X1 U12387 ( .A(n9880), .ZN(n9883) );
  NAND2_X1 U12388 ( .A1(n14727), .A2(n9884), .ZN(n9889) );
  OR2_X1 U12389 ( .A1(n10943), .A2(n13729), .ZN(n9885) );
  OAI21_X1 U12390 ( .B1(n10886), .B2(n13728), .A(n9885), .ZN(n9888) );
  XNOR2_X1 U12391 ( .A(n9889), .B(n9888), .ZN(n10670) );
  OAI22_X1 U12392 ( .A1(n10943), .A2(n9886), .B1(n10886), .B2(n13729), .ZN(
        n9887) );
  XOR2_X1 U12393 ( .A(n6549), .B(n9887), .Z(n10671) );
  NOR2_X1 U12394 ( .A1(n10670), .A2(n10671), .ZN(n10669) );
  AND2_X1 U12395 ( .A1(n9889), .A2(n9888), .ZN(n9890) );
  AOI22_X1 U12396 ( .A1(n10921), .A2(n9891), .B1(n9892), .B2(n13918), .ZN(
        n9894) );
  AOI22_X1 U12397 ( .A1(n10921), .A2(n13798), .B1(n9891), .B2(n13918), .ZN(
        n9893) );
  XNOR2_X1 U12398 ( .A(n9893), .B(n6549), .ZN(n10694) );
  AOI22_X1 U12399 ( .A1(n14788), .A2(n13798), .B1(n9891), .B2(n13917), .ZN(
        n9895) );
  XNOR2_X1 U12400 ( .A(n9895), .B(n6549), .ZN(n9897) );
  AND2_X1 U12401 ( .A1(n9892), .A2(n13917), .ZN(n9896) );
  AOI21_X1 U12402 ( .B1(n14788), .B2(n9891), .A(n9896), .ZN(n9898) );
  XNOR2_X1 U12403 ( .A(n9897), .B(n9898), .ZN(n10929) );
  AND2_X1 U12404 ( .A1(n9892), .A2(n14770), .ZN(n9899) );
  AOI21_X1 U12405 ( .B1(n10978), .B2(n9891), .A(n9899), .ZN(n11174) );
  AOI22_X1 U12406 ( .A1(n10978), .A2(n13798), .B1(n9891), .B2(n14770), .ZN(
        n9900) );
  XNOR2_X1 U12407 ( .A(n9900), .B(n6549), .ZN(n11173) );
  XOR2_X1 U12408 ( .A(n11174), .B(n11173), .Z(n11177) );
  XNOR2_X1 U12409 ( .A(n11178), .B(n11177), .ZN(n9924) );
  INV_X1 U12410 ( .A(n9901), .ZN(n9902) );
  AND2_X1 U12411 ( .A1(n14920), .A2(n10032), .ZN(n9923) );
  NAND2_X1 U12412 ( .A1(n9903), .A2(P1_B_REG_SCAN_IN), .ZN(n9904) );
  MUX2_X1 U12413 ( .A(P1_B_REG_SCAN_IN), .B(n9904), .S(n11743), .Z(n9907) );
  INV_X1 U12414 ( .A(n9905), .ZN(n9906) );
  NOR2_X1 U12415 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .ZN(
        n9911) );
  NOR4_X1 U12416 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9910) );
  NOR4_X1 U12417 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9909) );
  NOR4_X1 U12418 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9908) );
  NAND4_X1 U12419 ( .A1(n9911), .A2(n9910), .A3(n9909), .A4(n9908), .ZN(n9917)
         );
  NOR4_X1 U12420 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9915) );
  NOR4_X1 U12421 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9914) );
  NOR4_X1 U12422 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9913) );
  NOR4_X1 U12423 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9912) );
  NAND4_X1 U12424 ( .A1(n9915), .A2(n9914), .A3(n9913), .A4(n9912), .ZN(n9916)
         );
  NOR2_X1 U12425 ( .A1(n9917), .A2(n9916), .ZN(n9918) );
  OR2_X1 U12426 ( .A1(n10007), .A2(n9918), .ZN(n9925) );
  INV_X1 U12427 ( .A(n10036), .ZN(n10008) );
  AND2_X1 U12428 ( .A1(n9925), .A2(n10008), .ZN(n9949) );
  OR2_X1 U12429 ( .A1(n10007), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9920) );
  NAND2_X1 U12430 ( .A1(n9905), .A2(n11743), .ZN(n9919) );
  AND2_X1 U12431 ( .A1(n9920), .A2(n9919), .ZN(n9948) );
  OR2_X1 U12432 ( .A1(n10007), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9922) );
  NAND2_X1 U12433 ( .A1(n9905), .A2(n9903), .ZN(n9921) );
  NOR2_X1 U12434 ( .A1(n9924), .A2(n13908), .ZN(n9936) );
  NAND3_X1 U12435 ( .A1(n10315), .A2(n9948), .A3(n9925), .ZN(n9926) );
  NOR2_X4 U12436 ( .A1(n9951), .A2(n9952), .ZN(n14812) );
  NAND2_X1 U12437 ( .A1(n9926), .A2(n10316), .ZN(n9929) );
  AND2_X1 U12438 ( .A1(n9929), .A2(n10008), .ZN(n14725) );
  AND2_X1 U12439 ( .A1(n13905), .A2(n10978), .ZN(n9935) );
  NOR2_X1 U12440 ( .A1(n9947), .A2(n9927), .ZN(n9928) );
  NAND2_X1 U12441 ( .A1(n9929), .A2(n9928), .ZN(n9930) );
  AOI21_X2 U12442 ( .B1(n9930), .B2(P1_STATE_REG_SCAN_IN), .A(n11379), .ZN(
        n14736) );
  INV_X1 U12443 ( .A(n9931), .ZN(n10906) );
  NOR2_X1 U12444 ( .A1(n14736), .A2(n10906), .ZN(n9934) );
  INV_X1 U12445 ( .A(n13916), .ZN(n11214) );
  NAND2_X1 U12446 ( .A1(n14733), .A2(n14769), .ZN(n14660) );
  NAND2_X1 U12447 ( .A1(n13901), .A2(n13917), .ZN(n9932) );
  NAND2_X1 U12448 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10112) );
  OAI211_X1 U12449 ( .C1(n11214), .C2(n14660), .A(n9932), .B(n10112), .ZN(
        n9933) );
  OR4_X1 U12450 ( .A1(n9936), .A2(n9935), .A3(n9934), .A4(n9933), .ZN(P1_U3213) );
  NAND2_X1 U12451 ( .A1(n6720), .A2(n14039), .ZN(n9938) );
  AOI21_X1 U12452 ( .B1(n10865), .B2(n9943), .A(n14802), .ZN(n9942) );
  NAND2_X1 U12453 ( .A1(n10862), .A2(n10458), .ZN(n14811) );
  OAI21_X1 U12454 ( .B1(n10862), .B2(n10458), .A(n14811), .ZN(n9955) );
  XNOR2_X1 U12455 ( .A(n9028), .B(n9955), .ZN(n9940) );
  OAI21_X1 U12456 ( .B1(n9940), .B2(n14802), .A(n9939), .ZN(n9941) );
  OAI21_X1 U12457 ( .B1(n9942), .B2(n14771), .A(n9941), .ZN(n9946) );
  XNOR2_X1 U12458 ( .A(n10865), .B(n10864), .ZN(n10451) );
  OR2_X1 U12459 ( .A1(n9862), .A2(n9861), .ZN(n9944) );
  NAND2_X1 U12460 ( .A1(n6549), .A2(n9944), .ZN(n14130) );
  OR2_X1 U12461 ( .A1(n14130), .A2(n14039), .ZN(n10988) );
  NAND2_X1 U12462 ( .A1(n10451), .A2(n14899), .ZN(n9945) );
  OAI211_X1 U12463 ( .C1(n10874), .C2(n14240), .A(n9946), .B(n9945), .ZN(
        n10449) );
  NOR2_X1 U12464 ( .A1(n9948), .A2(n9947), .ZN(n9950) );
  NAND2_X1 U12465 ( .A1(n10318), .A2(n10315), .ZN(n14113) );
  MUX2_X1 U12466 ( .A(n10449), .B(P1_REG2_REG_1__SCAN_IN), .S(n14833), .Z(
        n9959) );
  INV_X1 U12467 ( .A(n9951), .ZN(n10321) );
  NAND2_X1 U12468 ( .A1(n10321), .A2(n9952), .ZN(n9953) );
  INV_X1 U12469 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13926) );
  OAI22_X1 U12470 ( .A1(n14808), .A2(n10862), .B1(n14775), .B2(n13926), .ZN(
        n9958) );
  INV_X1 U12471 ( .A(n10451), .ZN(n9956) );
  INV_X1 U12472 ( .A(n14812), .ZN(n14292) );
  OR2_X1 U12473 ( .A1(n9955), .A2(n14292), .ZN(n10448) );
  OAI22_X1 U12474 ( .A1(n9956), .A2(n14299), .B1(n14308), .B2(n10448), .ZN(
        n9957) );
  OR3_X1 U12475 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(P1_U3292) );
  NAND2_X2 U12476 ( .A1(n9981), .A2(P1_U3086), .ZN(n14455) );
  INV_X1 U12477 ( .A(n9961), .ZN(n9997) );
  INV_X1 U12478 ( .A(n10249), .ZN(n10101) );
  OAI222_X1 U12479 ( .A1(n14455), .A2(n9962), .B1(n14458), .B2(n9997), .C1(
        n10101), .C2(P1_U3086), .ZN(P1_U3353) );
  NOR2_X2 U12480 ( .A1(n9981), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14587) );
  INV_X1 U12481 ( .A(n14587), .ZN(n14576) );
  OAI222_X1 U12482 ( .A1(n6546), .A2(P3_U3151), .B1(n14576), .B2(n9964), .C1(
        n9963), .C2(n14574), .ZN(P3_U3294) );
  OAI222_X1 U12483 ( .A1(n15231), .A2(P3_U3151), .B1(n14576), .B2(n9966), .C1(
        n9965), .C2(n14574), .ZN(P3_U3289) );
  OAI222_X1 U12484 ( .A1(P3_U3151), .A2(n15268), .B1(n14574), .B2(n9968), .C1(
        n14576), .C2(n9967), .ZN(P3_U3287) );
  INV_X1 U12485 ( .A(n14574), .ZN(n14586) );
  AOI222_X1 U12486 ( .A1(n9969), .A2(n14587), .B1(SI_9_), .B2(n14586), .C1(
        n11135), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9970) );
  INV_X1 U12487 ( .A(n9970), .ZN(P3_U3286) );
  AOI222_X1 U12488 ( .A1(n9971), .A2(n14587), .B1(SI_7_), .B2(n14586), .C1(
        n11131), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9972) );
  INV_X1 U12489 ( .A(n9972), .ZN(P3_U3288) );
  AOI222_X1 U12490 ( .A1(n9973), .A2(n14587), .B1(n11125), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n14586), .ZN(n9974) );
  INV_X1 U12491 ( .A(n9974), .ZN(P3_U3291) );
  AOI222_X1 U12492 ( .A1(n9975), .A2(n14587), .B1(n11127), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_5_), .C2(n14586), .ZN(n9976) );
  INV_X1 U12493 ( .A(n9976), .ZN(P3_U3290) );
  AOI222_X1 U12494 ( .A1(n9977), .A2(n14587), .B1(n15180), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n14586), .ZN(n9978) );
  INV_X1 U12495 ( .A(n9978), .ZN(P3_U3292) );
  AOI222_X1 U12496 ( .A1(n9979), .A2(n14587), .B1(n6552), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_2_), .C2(n14586), .ZN(n9980) );
  INV_X1 U12497 ( .A(n9980), .ZN(P3_U3293) );
  AND2_X1 U12498 ( .A1(n9960), .A2(P2_U3088), .ZN(n11382) );
  INV_X2 U12499 ( .A(n11382), .ZN(n13395) );
  NAND2_X2 U12500 ( .A1(n9981), .A2(P2_U3088), .ZN(n13393) );
  AOI222_X1 U12501 ( .A1(n9983), .A2(n14587), .B1(SI_10_), .B2(n14586), .C1(
        n11117), .C2(P3_STATE_REG_SCAN_IN), .ZN(n9984) );
  INV_X1 U12502 ( .A(n9984), .ZN(P3_U3285) );
  INV_X1 U12503 ( .A(n9985), .ZN(n9992) );
  OAI222_X1 U12504 ( .A1(n14455), .A2(n8049), .B1(n14458), .B2(n9992), .C1(
        n13935), .C2(P1_U3086), .ZN(P1_U3352) );
  INV_X1 U12505 ( .A(n9986), .ZN(n9993) );
  INV_X1 U12506 ( .A(n13954), .ZN(n13948) );
  OAI222_X1 U12507 ( .A1(n14455), .A2(n6713), .B1(n14458), .B2(n9993), .C1(
        n13948), .C2(P1_U3086), .ZN(P1_U3351) );
  INV_X1 U12508 ( .A(n10105), .ZN(n10272) );
  INV_X1 U12509 ( .A(n9987), .ZN(n9995) );
  INV_X1 U12510 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9988) );
  OAI222_X1 U12511 ( .A1(n10272), .A2(P1_U3086), .B1(n14458), .B2(n9995), .C1(
        n9988), .C2(n14455), .ZN(P1_U3350) );
  INV_X1 U12512 ( .A(n13928), .ZN(n10100) );
  AOI22_X1 U12513 ( .A1(n12992), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n11382), .ZN(n9991) );
  OAI21_X1 U12514 ( .B1(n9992), .B2(n13393), .A(n9991), .ZN(P2_U3324) );
  INV_X1 U12515 ( .A(n10076), .ZN(n14973) );
  OAI222_X1 U12516 ( .A1(n13395), .A2(n9994), .B1(n13393), .B2(n9993), .C1(
        P2_U3088), .C2(n14973), .ZN(P2_U3323) );
  OAI222_X1 U12517 ( .A1(n13395), .A2(n9996), .B1(n13393), .B2(n9995), .C1(
        P2_U3088), .C2(n10087), .ZN(P2_U3322) );
  INV_X1 U12518 ( .A(n10074), .ZN(n14960) );
  OAI222_X1 U12519 ( .A1(n13395), .A2(n9998), .B1(n13393), .B2(n9997), .C1(
        P2_U3088), .C2(n14960), .ZN(P2_U3325) );
  INV_X1 U12520 ( .A(n10107), .ZN(n13965) );
  INV_X1 U12521 ( .A(n9999), .ZN(n10001) );
  OAI222_X1 U12522 ( .A1(n13965), .A2(P1_U3086), .B1(n14458), .B2(n10001), 
        .C1(n10000), .C2(n14455), .ZN(P1_U3349) );
  INV_X1 U12523 ( .A(n10127), .ZN(n10147) );
  OAI222_X1 U12524 ( .A1(n13395), .A2(n10002), .B1(n13393), .B2(n10001), .C1(
        P2_U3088), .C2(n10147), .ZN(P2_U3321) );
  INV_X1 U12525 ( .A(n10115), .ZN(n10258) );
  INV_X1 U12526 ( .A(n10003), .ZN(n10005) );
  OAI222_X1 U12527 ( .A1(n10258), .A2(P1_U3086), .B1(n14458), .B2(n10005), 
        .C1(n10004), .C2(n14455), .ZN(P1_U3348) );
  INV_X1 U12528 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10006) );
  INV_X1 U12529 ( .A(n10155), .ZN(n10134) );
  OAI222_X1 U12530 ( .A1(n13395), .A2(n10006), .B1(n13393), .B2(n10005), .C1(
        P2_U3088), .C2(n10134), .ZN(P2_U3320) );
  INV_X1 U12531 ( .A(n11743), .ZN(n10010) );
  NAND2_X1 U12532 ( .A1(n9905), .A2(n10009), .ZN(n10012) );
  OAI22_X1 U12533 ( .A1(n14864), .A2(P1_D_REG_0__SCAN_IN), .B1(n10010), .B2(
        n10012), .ZN(n10011) );
  INV_X1 U12534 ( .A(n10011), .ZN(P1_U3445) );
  INV_X1 U12535 ( .A(n9903), .ZN(n10013) );
  OAI22_X1 U12536 ( .A1(n14864), .A2(P1_D_REG_1__SCAN_IN), .B1(n10013), .B2(
        n10012), .ZN(n10014) );
  INV_X1 U12537 ( .A(n10014), .ZN(P1_U3446) );
  INV_X1 U12538 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10016) );
  INV_X1 U12539 ( .A(n10015), .ZN(n10018) );
  INV_X1 U12540 ( .A(n10184), .ZN(n10162) );
  OAI222_X1 U12541 ( .A1(n13395), .A2(n10016), .B1(n13393), .B2(n10018), .C1(
        P2_U3088), .C2(n10162), .ZN(P2_U3319) );
  INV_X1 U12542 ( .A(n10287), .ZN(n10282) );
  OAI222_X1 U12543 ( .A1(n10282), .A2(P1_U3086), .B1(n14458), .B2(n10018), 
        .C1(n10017), .C2(n14455), .ZN(P1_U3347) );
  INV_X1 U12544 ( .A(n10288), .ZN(n10375) );
  INV_X1 U12545 ( .A(n10019), .ZN(n10021) );
  OAI222_X1 U12546 ( .A1(n10375), .A2(P1_U3086), .B1(n14458), .B2(n10021), 
        .C1(n10020), .C2(n14455), .ZN(P1_U3346) );
  INV_X1 U12547 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10022) );
  INV_X1 U12548 ( .A(n10495), .ZN(n10188) );
  OAI222_X1 U12549 ( .A1(n13395), .A2(n10022), .B1(n13393), .B2(n10021), .C1(
        P2_U3088), .C2(n10188), .ZN(P2_U3318) );
  INV_X1 U12550 ( .A(n10377), .ZN(n13983) );
  INV_X1 U12551 ( .A(n10023), .ZN(n10026) );
  OAI222_X1 U12552 ( .A1(n13983), .A2(P1_U3086), .B1(n14458), .B2(n10026), 
        .C1(n10024), .C2(n14455), .ZN(P1_U3345) );
  INV_X1 U12553 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10027) );
  INV_X1 U12554 ( .A(n14990), .ZN(n10025) );
  OAI222_X1 U12555 ( .A1(n13395), .A2(n10027), .B1(n13393), .B2(n10026), .C1(
        P2_U3088), .C2(n10025), .ZN(P2_U3317) );
  OAI222_X1 U12556 ( .A1(P3_U3151), .A2(n12273), .B1(n14574), .B2(n10029), 
        .C1(n14576), .C2(n10028), .ZN(P3_U3282) );
  INV_X1 U12557 ( .A(n10030), .ZN(n10031) );
  OR2_X1 U12558 ( .A1(n10032), .A2(n10031), .ZN(n10034) );
  NAND2_X1 U12559 ( .A1(n10034), .A2(n10033), .ZN(n10040) );
  NAND2_X1 U12560 ( .A1(n10036), .A2(n10035), .ZN(n10041) );
  INV_X1 U12561 ( .A(n14756), .ZN(n13987) );
  NOR2_X1 U12562 ( .A1(n13987), .A2(P1_U4016), .ZN(P1_U3085) );
  NAND2_X1 U12563 ( .A1(n10814), .A2(n10039), .ZN(n10037) );
  OAI21_X1 U12564 ( .B1(n10039), .B2(n8007), .A(n10037), .ZN(P3_U3376) );
  NAND2_X1 U12565 ( .A1(n10744), .A2(n10039), .ZN(n10038) );
  OAI21_X1 U12566 ( .B1(n10039), .B2(n8004), .A(n10038), .ZN(P3_U3377) );
  INV_X1 U12567 ( .A(n10040), .ZN(n10042) );
  INV_X1 U12568 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10043) );
  NAND3_X1 U12569 ( .A1(n14748), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10043), .ZN(
        n10049) );
  INV_X1 U12570 ( .A(n14454), .ZN(n10095) );
  NOR2_X1 U12571 ( .A1(n14454), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n10044) );
  NOR2_X1 U12572 ( .A1(n9580), .A2(n10044), .ZN(n10238) );
  OAI21_X1 U12573 ( .B1(n10095), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10238), .ZN(
        n10045) );
  MUX2_X1 U12574 ( .A(n10045), .B(n10238), .S(P1_IR_REG_0__SCAN_IN), .Z(n10046) );
  INV_X1 U12575 ( .A(n10046), .ZN(n10047) );
  AOI22_X1 U12576 ( .A1(n10094), .A2(n10047), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10048) );
  OAI211_X1 U12577 ( .C1(n14756), .C2(n7185), .A(n10049), .B(n10048), .ZN(
        P1_U3243) );
  INV_X1 U12578 ( .A(n10562), .ZN(n10373) );
  INV_X1 U12579 ( .A(n10050), .ZN(n10052) );
  OAI222_X1 U12580 ( .A1(n10373), .A2(P1_U3086), .B1(n14458), .B2(n10052), 
        .C1(n10051), .C2(n14455), .ZN(P1_U3344) );
  INV_X1 U12581 ( .A(n10541), .ZN(n10544) );
  OAI222_X1 U12582 ( .A1(n13395), .A2(n10053), .B1(n13393), .B2(n10052), .C1(
        P2_U3088), .C2(n10544), .ZN(P2_U3316) );
  AOI21_X1 U12583 ( .B1(n10055), .B2(n10054), .A(n8389), .ZN(n10057) );
  NOR2_X1 U12584 ( .A1(n10067), .A2(P2_U3088), .ZN(n10058) );
  XNOR2_X1 U12585 ( .A(n10074), .B(n10059), .ZN(n14959) );
  XNOR2_X1 U12586 ( .A(n14947), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14946) );
  AND2_X1 U12587 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n14945) );
  NAND2_X1 U12588 ( .A1(n14946), .A2(n14945), .ZN(n10062) );
  NAND2_X1 U12589 ( .A1(n10060), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10061) );
  NAND2_X1 U12590 ( .A1(n10062), .A2(n10061), .ZN(n14958) );
  NAND2_X1 U12591 ( .A1(n14959), .A2(n14958), .ZN(n14957) );
  NAND2_X1 U12592 ( .A1(n10074), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U12593 ( .A1(n14957), .A2(n10063), .ZN(n12990) );
  INV_X1 U12594 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10064) );
  XNOR2_X1 U12595 ( .A(n12992), .B(n10064), .ZN(n12991) );
  NAND2_X1 U12596 ( .A1(n12990), .A2(n12991), .ZN(n12989) );
  NAND2_X1 U12597 ( .A1(n12992), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10065) );
  NAND2_X1 U12598 ( .A1(n12989), .A2(n10065), .ZN(n14970) );
  XNOR2_X1 U12599 ( .A(n10076), .B(n10066), .ZN(n14969) );
  XNOR2_X1 U12600 ( .A(n10126), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n10069) );
  NOR2_X1 U12601 ( .A1(n10070), .A2(n10069), .ZN(n10121) );
  NAND2_X1 U12602 ( .A1(n10067), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13381) );
  INV_X1 U12603 ( .A(n13381), .ZN(n10068) );
  AOI211_X1 U12604 ( .C1(n10070), .C2(n10069), .A(n10121), .B(n15001), .ZN(
        n10083) );
  INV_X1 U12605 ( .A(n13385), .ZN(n10071) );
  INV_X1 U12606 ( .A(n15009), .ZN(n14993) );
  MUX2_X1 U12607 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n10073), .S(n10074), .Z(
        n14964) );
  MUX2_X1 U12608 ( .A(n10354), .B(P2_REG2_REG_1__SCAN_IN), .S(n14947), .Z(
        n14952) );
  NAND3_X1 U12609 ( .A1(n14952), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG2_REG_0__SCAN_IN), .ZN(n14951) );
  OAI21_X1 U12610 ( .B1(n14947), .B2(n10354), .A(n14951), .ZN(n14965) );
  NAND2_X1 U12611 ( .A1(n14964), .A2(n14965), .ZN(n14963) );
  NAND2_X1 U12612 ( .A1(n10074), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n12994) );
  MUX2_X1 U12613 ( .A(n10432), .B(P2_REG2_REG_3__SCAN_IN), .S(n12992), .Z(
        n12995) );
  AOI21_X1 U12614 ( .B1(n14963), .B2(n12994), .A(n12995), .ZN(n12993) );
  AOI21_X1 U12615 ( .B1(n12992), .B2(P2_REG2_REG_3__SCAN_IN), .A(n12993), .ZN(
        n14979) );
  INV_X1 U12616 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10075) );
  MUX2_X1 U12617 ( .A(n10075), .B(P2_REG2_REG_4__SCAN_IN), .S(n10076), .Z(
        n14978) );
  NOR2_X1 U12618 ( .A1(n14979), .A2(n14978), .ZN(n14977) );
  AND2_X1 U12619 ( .A1(n10076), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10079) );
  MUX2_X1 U12620 ( .A(n10077), .B(P2_REG2_REG_5__SCAN_IN), .S(n10087), .Z(
        n10078) );
  OAI21_X1 U12621 ( .B1(n14977), .B2(n10079), .A(n10078), .ZN(n10143) );
  INV_X1 U12622 ( .A(n10143), .ZN(n10081) );
  NOR3_X1 U12623 ( .A1(n14977), .A2(n10079), .A3(n10078), .ZN(n10080) );
  NOR3_X1 U12624 ( .A1(n14993), .A2(n10081), .A3(n10080), .ZN(n10082) );
  NOR2_X1 U12625 ( .A1(n10083), .A2(n10082), .ZN(n10086) );
  NOR2_X2 U12626 ( .A1(n10084), .A2(P2_U3088), .ZN(n15007) );
  NOR2_X1 U12627 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8276), .ZN(n10474) );
  AOI21_X1 U12628 ( .B1(n15007), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10474), .ZN(
        n10085) );
  OAI211_X1 U12629 ( .C1(n10087), .C2(n15014), .A(n10086), .B(n10085), .ZN(
        P2_U3219) );
  MUX2_X1 U12630 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10088), .S(n10249), .Z(
        n10241) );
  MUX2_X1 U12631 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n10089), .S(n13928), .Z(
        n13930) );
  AND2_X1 U12632 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13931) );
  NAND2_X1 U12633 ( .A1(n13930), .A2(n13931), .ZN(n13929) );
  NAND2_X1 U12634 ( .A1(n13928), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U12635 ( .A1(n13929), .A2(n10090), .ZN(n10240) );
  AOI22_X1 U12636 ( .A1(n10241), .A2(n10240), .B1(n10249), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n13943) );
  MUX2_X1 U12637 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10876), .S(n13935), .Z(
        n13942) );
  NOR2_X1 U12638 ( .A1(n13943), .A2(n13942), .ZN(n13960) );
  NOR2_X1 U12639 ( .A1(n13935), .A2(n10876), .ZN(n13955) );
  MUX2_X1 U12640 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10091), .S(n13954), .Z(
        n10092) );
  OAI21_X1 U12641 ( .B1(n13960), .B2(n13955), .A(n10092), .ZN(n13958) );
  NAND2_X1 U12642 ( .A1(n13954), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10275) );
  MUX2_X1 U12643 ( .A(n10920), .B(P1_REG2_REG_5__SCAN_IN), .S(n10105), .Z(
        n10274) );
  AOI21_X1 U12644 ( .B1(n13958), .B2(n10275), .A(n10274), .ZN(n13973) );
  NOR2_X1 U12645 ( .A1(n10272), .A2(n10920), .ZN(n13972) );
  MUX2_X1 U12646 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10093), .S(n10107), .Z(
        n13971) );
  OAI21_X1 U12647 ( .B1(n13973), .B2(n13972), .A(n13971), .ZN(n13975) );
  NAND2_X1 U12648 ( .A1(n10107), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10098) );
  MUX2_X1 U12649 ( .A(n10904), .B(P1_REG2_REG_7__SCAN_IN), .S(n10115), .Z(
        n10097) );
  AOI21_X1 U12650 ( .B1(n13975), .B2(n10098), .A(n10097), .ZN(n10265) );
  INV_X1 U12651 ( .A(n10094), .ZN(n10111) );
  NAND2_X1 U12652 ( .A1(n10235), .A2(n10095), .ZN(n10096) );
  NOR2_X2 U12653 ( .A1(n10111), .A2(n10096), .ZN(n14752) );
  NAND3_X1 U12654 ( .A1(n13975), .A2(n10098), .A3(n10097), .ZN(n10099) );
  NAND2_X1 U12655 ( .A1(n14752), .A2(n10099), .ZN(n10118) );
  INV_X1 U12656 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10108) );
  INV_X1 U12657 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n10106) );
  INV_X1 U12658 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n10104) );
  INV_X1 U12659 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10103) );
  INV_X1 U12660 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10102) );
  NAND3_X1 U12661 ( .A1(n13925), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n13923) );
  OAI21_X1 U12662 ( .B1(n6852), .B2(n10100), .A(n13923), .ZN(n10243) );
  MUX2_X1 U12663 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10102), .S(n10249), .Z(
        n10244) );
  NAND2_X1 U12664 ( .A1(n10243), .A2(n10244), .ZN(n10242) );
  OAI21_X1 U12665 ( .B1(n10102), .B2(n10101), .A(n10242), .ZN(n13939) );
  MUX2_X1 U12666 ( .A(n10103), .B(P1_REG1_REG_3__SCAN_IN), .S(n13935), .Z(
        n13940) );
  NAND2_X1 U12667 ( .A1(n13939), .A2(n13940), .ZN(n13938) );
  OAI21_X1 U12668 ( .B1(n10103), .B2(n13935), .A(n13938), .ZN(n13952) );
  MUX2_X1 U12669 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n10104), .S(n13954), .Z(
        n13953) );
  NAND2_X1 U12670 ( .A1(n13952), .A2(n13953), .ZN(n13951) );
  OAI21_X1 U12671 ( .B1(n13948), .B2(n10104), .A(n13951), .ZN(n10270) );
  XNOR2_X1 U12672 ( .A(n10105), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n10271) );
  NOR2_X1 U12673 ( .A1(n10270), .A2(n10271), .ZN(n10269) );
  XOR2_X1 U12674 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n10107), .Z(n13970) );
  INV_X1 U12675 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n14931) );
  MUX2_X1 U12676 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n14931), .S(n10115), .Z(
        n10109) );
  OAI211_X1 U12677 ( .C1(n10110), .C2(n10109), .A(n10253), .B(n14748), .ZN(
        n10117) );
  INV_X1 U12678 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10113) );
  OAI21_X1 U12679 ( .B1(n14756), .B2(n10113), .A(n10112), .ZN(n10114) );
  AOI21_X1 U12680 ( .B1(n14750), .B2(n10115), .A(n10114), .ZN(n10116) );
  OAI211_X1 U12681 ( .C1(n10265), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        P1_U3250) );
  OAI222_X1 U12682 ( .A1(P3_U3151), .A2(n12293), .B1(n14574), .B2(n10120), 
        .C1(n14576), .C2(n10119), .ZN(P3_U3281) );
  AOI21_X1 U12683 ( .B1(n10126), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10121), .ZN(
        n10140) );
  INV_X1 U12684 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10122) );
  MUX2_X1 U12685 ( .A(n10122), .B(P2_REG1_REG_6__SCAN_IN), .S(n10127), .Z(
        n10139) );
  INV_X1 U12686 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10123) );
  MUX2_X1 U12687 ( .A(n10123), .B(P2_REG1_REG_7__SCAN_IN), .S(n10155), .Z(
        n10124) );
  AOI211_X1 U12688 ( .C1(n10125), .C2(n10124), .A(n15001), .B(n10151), .ZN(
        n10137) );
  NAND2_X1 U12689 ( .A1(n10126), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10142) );
  MUX2_X1 U12690 ( .A(n13252), .B(P2_REG2_REG_6__SCAN_IN), .S(n10127), .Z(
        n10141) );
  AOI21_X1 U12691 ( .B1(n10143), .B2(n10142), .A(n10141), .ZN(n10145) );
  NOR2_X1 U12692 ( .A1(n10147), .A2(n13252), .ZN(n10129) );
  MUX2_X1 U12693 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n10660), .S(n10155), .Z(
        n10128) );
  OAI21_X1 U12694 ( .B1(n10145), .B2(n10129), .A(n10128), .ZN(n10158) );
  INV_X1 U12695 ( .A(n10158), .ZN(n10131) );
  NOR3_X1 U12696 ( .A1(n10145), .A2(n10129), .A3(n10128), .ZN(n10130) );
  NOR3_X1 U12697 ( .A1(n10131), .A2(n10130), .A3(n14993), .ZN(n10136) );
  NOR2_X1 U12698 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8318), .ZN(n10132) );
  AOI21_X1 U12699 ( .B1(n15007), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n10132), .ZN(
        n10133) );
  OAI21_X1 U12700 ( .B1(n10134), .B2(n15014), .A(n10133), .ZN(n10135) );
  OR3_X1 U12701 ( .A1(n10137), .A2(n10136), .A3(n10135), .ZN(P2_U3221) );
  AOI211_X1 U12702 ( .C1(n10140), .C2(n10139), .A(n15001), .B(n10138), .ZN(
        n10150) );
  AND3_X1 U12703 ( .A1(n10143), .A2(n10142), .A3(n10141), .ZN(n10144) );
  NOR3_X1 U12704 ( .A1(n10145), .A2(n14993), .A3(n10144), .ZN(n10149) );
  NAND2_X1 U12705 ( .A1(n15007), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10146) );
  NAND2_X1 U12706 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n10484) );
  OAI211_X1 U12707 ( .C1(n15014), .C2(n10147), .A(n10146), .B(n10484), .ZN(
        n10148) );
  OR3_X1 U12708 ( .A1(n10150), .A2(n10149), .A3(n10148), .ZN(P2_U3220) );
  MUX2_X1 U12709 ( .A(n10152), .B(P2_REG1_REG_8__SCAN_IN), .S(n10184), .Z(
        n10153) );
  NOR2_X1 U12710 ( .A1(n10154), .A2(n10153), .ZN(n10178) );
  AOI211_X1 U12711 ( .C1(n10154), .C2(n10153), .A(n15001), .B(n10178), .ZN(
        n10165) );
  NAND2_X1 U12712 ( .A1(n10155), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10157) );
  MUX2_X1 U12713 ( .A(n8338), .B(P2_REG2_REG_8__SCAN_IN), .S(n10184), .Z(
        n10156) );
  AOI21_X1 U12714 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10183) );
  AND3_X1 U12715 ( .A1(n10158), .A2(n10157), .A3(n10156), .ZN(n10159) );
  NOR3_X1 U12716 ( .A1(n10183), .A2(n10159), .A3(n14993), .ZN(n10164) );
  NOR2_X1 U12717 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n13652), .ZN(n10160) );
  AOI21_X1 U12718 ( .B1(n15007), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10160), .ZN(
        n10161) );
  OAI21_X1 U12719 ( .B1(n10162), .B2(n15014), .A(n10161), .ZN(n10163) );
  OR3_X1 U12720 ( .A1(n10165), .A2(n10164), .A3(n10163), .ZN(P2_U3222) );
  OR2_X1 U12721 ( .A1(n10166), .A2(n15086), .ZN(n11863) );
  AOI22_X1 U12722 ( .A1(n8784), .A2(n10167), .B1(n11863), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10171) );
  NOR2_X1 U12723 ( .A1(n8842), .A2(n12886), .ZN(n15040) );
  AOI22_X1 U12724 ( .A1(n12950), .A2(n15040), .B1(n10169), .B2(n10168), .ZN(
        n10170) );
  OAI211_X1 U12725 ( .C1(n12938), .C2(n10172), .A(n10171), .B(n10170), .ZN(
        P2_U3204) );
  INV_X1 U12726 ( .A(n10173), .ZN(n10176) );
  INV_X1 U12727 ( .A(n10796), .ZN(n10801) );
  OAI222_X1 U12728 ( .A1(n13393), .A2(n10176), .B1(n10801), .B2(P2_U3088), 
        .C1(n10174), .C2(n13395), .ZN(P2_U3315) );
  INV_X1 U12729 ( .A(n14751), .ZN(n10177) );
  OAI222_X1 U12730 ( .A1(P1_U3086), .A2(n10177), .B1(n14458), .B2(n10176), 
        .C1(n10175), .C2(n14455), .ZN(P1_U3343) );
  AOI21_X1 U12731 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n10184), .A(n10178), .ZN(
        n10181) );
  MUX2_X1 U12732 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10179), .S(n10495), .Z(
        n10180) );
  NAND2_X1 U12733 ( .A1(n10181), .A2(n10180), .ZN(n10494) );
  OAI21_X1 U12734 ( .B1(n10181), .B2(n10180), .A(n10494), .ZN(n10182) );
  NAND2_X1 U12735 ( .A1(n10182), .A2(n14976), .ZN(n10192) );
  AOI21_X1 U12736 ( .B1(n10184), .B2(P2_REG2_REG_8__SCAN_IN), .A(n10183), .ZN(
        n10186) );
  MUX2_X1 U12737 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8351), .S(n10495), .Z(
        n10185) );
  NAND2_X1 U12738 ( .A1(n10186), .A2(n10185), .ZN(n10489) );
  OAI21_X1 U12739 ( .B1(n10186), .B2(n10185), .A(n10489), .ZN(n10190) );
  NAND2_X1 U12740 ( .A1(n15007), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n10187) );
  NAND2_X1 U12741 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n11001) );
  OAI211_X1 U12742 ( .C1(n15014), .C2(n10188), .A(n10187), .B(n11001), .ZN(
        n10189) );
  AOI21_X1 U12743 ( .B1(n10190), .B2(n15009), .A(n10189), .ZN(n10191) );
  NAND2_X1 U12744 ( .A1(n10192), .A2(n10191), .ZN(P2_U3223) );
  INV_X1 U12745 ( .A(n8784), .ZN(n12926) );
  OAI21_X1 U12746 ( .B1(n10195), .B2(n10194), .A(n10193), .ZN(n10196) );
  NAND2_X1 U12747 ( .A1(n10196), .A2(n12946), .ZN(n10198) );
  OAI22_X1 U12748 ( .A1(n8842), .A2(n12884), .B1(n7134), .B2(n12886), .ZN(
        n10335) );
  AOI22_X1 U12749 ( .A1(n12950), .A2(n10335), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n11863), .ZN(n10197) );
  OAI211_X1 U12750 ( .C1(n10331), .C2(n12926), .A(n10198), .B(n10197), .ZN(
        P2_U3209) );
  INV_X1 U12751 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U12752 ( .A1(n10225), .A2(n10200), .ZN(P3_U3234) );
  INV_X1 U12753 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10201) );
  NOR2_X1 U12754 ( .A1(n10209), .A2(n10201), .ZN(P3_U3235) );
  INV_X1 U12755 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10202) );
  NOR2_X1 U12756 ( .A1(n10209), .A2(n10202), .ZN(P3_U3236) );
  INV_X1 U12757 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n13614) );
  NOR2_X1 U12758 ( .A1(n10209), .A2(n13614), .ZN(P3_U3237) );
  INV_X1 U12759 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U12760 ( .A1(n10209), .A2(n10203), .ZN(P3_U3238) );
  INV_X1 U12761 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10204) );
  NOR2_X1 U12762 ( .A1(n10209), .A2(n10204), .ZN(P3_U3239) );
  INV_X1 U12763 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n13593) );
  NOR2_X1 U12764 ( .A1(n10209), .A2(n13593), .ZN(P3_U3240) );
  INV_X1 U12765 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n10205) );
  NOR2_X1 U12766 ( .A1(n10209), .A2(n10205), .ZN(P3_U3241) );
  INV_X1 U12767 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U12768 ( .A1(n10209), .A2(n10206), .ZN(P3_U3242) );
  INV_X1 U12769 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10207) );
  NOR2_X1 U12770 ( .A1(n10209), .A2(n10207), .ZN(P3_U3243) );
  INV_X1 U12771 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U12772 ( .A1(n10209), .A2(n10208), .ZN(P3_U3244) );
  INV_X1 U12773 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n13633) );
  NOR2_X1 U12774 ( .A1(n10225), .A2(n13633), .ZN(P3_U3253) );
  INV_X1 U12775 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U12776 ( .A1(n10225), .A2(n10210), .ZN(P3_U3254) );
  INV_X1 U12777 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12778 ( .A1(n10225), .A2(n10211), .ZN(P3_U3255) );
  INV_X1 U12779 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U12780 ( .A1(n10225), .A2(n10212), .ZN(P3_U3256) );
  INV_X1 U12781 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U12782 ( .A1(n10225), .A2(n10213), .ZN(P3_U3257) );
  INV_X1 U12783 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12784 ( .A1(n10209), .A2(n10214), .ZN(P3_U3258) );
  INV_X1 U12785 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12786 ( .A1(n10225), .A2(n10215), .ZN(P3_U3259) );
  INV_X1 U12787 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n13463) );
  NOR2_X1 U12788 ( .A1(n10225), .A2(n13463), .ZN(P3_U3260) );
  INV_X1 U12789 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U12790 ( .A1(n10225), .A2(n10216), .ZN(P3_U3261) );
  INV_X1 U12791 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U12792 ( .A1(n10225), .A2(n10217), .ZN(P3_U3262) );
  INV_X1 U12793 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U12794 ( .A1(n10225), .A2(n10218), .ZN(P3_U3263) );
  INV_X1 U12795 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U12796 ( .A1(n10225), .A2(n10219), .ZN(P3_U3245) );
  INV_X1 U12797 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n13628) );
  NOR2_X1 U12798 ( .A1(n10225), .A2(n13628), .ZN(P3_U3246) );
  INV_X1 U12799 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U12800 ( .A1(n10225), .A2(n10220), .ZN(P3_U3247) );
  INV_X1 U12801 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12802 ( .A1(n10225), .A2(n10221), .ZN(P3_U3248) );
  INV_X1 U12803 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12804 ( .A1(n10225), .A2(n10222), .ZN(P3_U3249) );
  INV_X1 U12805 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n13590) );
  NOR2_X1 U12806 ( .A1(n10225), .A2(n13590), .ZN(P3_U3250) );
  INV_X1 U12807 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U12808 ( .A1(n10225), .A2(n10223), .ZN(P3_U3251) );
  INV_X1 U12809 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U12810 ( .A1(n10225), .A2(n10224), .ZN(P3_U3252) );
  INV_X1 U12811 ( .A(n10724), .ZN(n10570) );
  INV_X1 U12812 ( .A(n10226), .ZN(n10251) );
  OAI222_X1 U12813 ( .A1(P1_U3086), .A2(n10570), .B1(n14458), .B2(n10251), 
        .C1(n13631), .C2(n14455), .ZN(P1_U3342) );
  XNOR2_X1 U12814 ( .A(n10227), .B(n10228), .ZN(n10231) );
  INV_X1 U12815 ( .A(n12986), .ZN(n10300) );
  OAI22_X1 U12816 ( .A1(n10300), .A2(n12884), .B1(n10470), .B2(n12886), .ZN(
        n10398) );
  AOI22_X1 U12817 ( .A1(n12950), .A2(n10398), .B1(n8784), .B2(n10433), .ZN(
        n10230) );
  MUX2_X1 U12818 ( .A(n12953), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n10229) );
  OAI211_X1 U12819 ( .C1(n10231), .C2(n12938), .A(n10230), .B(n10229), .ZN(
        P2_U3190) );
  AOI21_X1 U12820 ( .B1(n10234), .B2(n10233), .A(n10232), .ZN(n10455) );
  MUX2_X1 U12821 ( .A(n13931), .B(n10455), .S(n14454), .Z(n10236) );
  NAND2_X1 U12822 ( .A1(n10236), .A2(n10235), .ZN(n10237) );
  OAI211_X1 U12823 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10238), .A(n10237), .B(
        P1_U4016), .ZN(n13964) );
  INV_X1 U12824 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10239) );
  OAI22_X1 U12825 ( .A1(n14756), .A2(n7180), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10239), .ZN(n10248) );
  INV_X1 U12826 ( .A(n14752), .ZN(n13941) );
  XNOR2_X1 U12827 ( .A(n10241), .B(n10240), .ZN(n10246) );
  OAI211_X1 U12828 ( .C1(n10244), .C2(n10243), .A(n14748), .B(n10242), .ZN(
        n10245) );
  OAI21_X1 U12829 ( .B1(n13941), .B2(n10246), .A(n10245), .ZN(n10247) );
  AOI211_X1 U12830 ( .C1(n10249), .C2(n14750), .A(n10248), .B(n10247), .ZN(
        n10250) );
  NAND2_X1 U12831 ( .A1(n13964), .A2(n10250), .ZN(P1_U3245) );
  INV_X1 U12832 ( .A(n11153), .ZN(n11148) );
  OAI222_X1 U12833 ( .A1(n13395), .A2(n10252), .B1(n11148), .B2(P2_U3088), 
        .C1(n13393), .C2(n10251), .ZN(P2_U3314) );
  INV_X1 U12834 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14933) );
  MUX2_X1 U12835 ( .A(n14933), .B(P1_REG1_REG_8__SCAN_IN), .S(n10287), .Z(
        n10255) );
  OAI21_X1 U12836 ( .B1(n14931), .B2(n10258), .A(n10253), .ZN(n10254) );
  AOI21_X1 U12837 ( .B1(n10255), .B2(n10254), .A(n10281), .ZN(n10268) );
  NAND2_X1 U12838 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n11182) );
  INV_X1 U12839 ( .A(n11182), .ZN(n10257) );
  NOR2_X1 U12840 ( .A1(n13984), .A2(n10282), .ZN(n10256) );
  AOI211_X1 U12841 ( .C1(n13987), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10257), .B(
        n10256), .ZN(n10267) );
  NOR2_X1 U12842 ( .A1(n10258), .A2(n10904), .ZN(n10263) );
  INV_X1 U12843 ( .A(n10263), .ZN(n10261) );
  INV_X1 U12844 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10259) );
  MUX2_X1 U12845 ( .A(n10259), .B(P1_REG2_REG_8__SCAN_IN), .S(n10287), .Z(
        n10260) );
  NAND2_X1 U12846 ( .A1(n10261), .A2(n10260), .ZN(n10264) );
  MUX2_X1 U12847 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10259), .S(n10287), .Z(
        n10262) );
  OAI21_X1 U12848 ( .B1(n10265), .B2(n10263), .A(n10262), .ZN(n10291) );
  OAI211_X1 U12849 ( .C1(n10265), .C2(n10264), .A(n10291), .B(n14752), .ZN(
        n10266) );
  OAI211_X1 U12850 ( .C1(n10268), .C2(n14036), .A(n10267), .B(n10266), .ZN(
        P1_U3251) );
  AOI21_X1 U12851 ( .B1(n10271), .B2(n10270), .A(n10269), .ZN(n10280) );
  AND2_X1 U12852 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10699) );
  NOR2_X1 U12853 ( .A1(n13984), .A2(n10272), .ZN(n10273) );
  AOI211_X1 U12854 ( .C1(n13987), .C2(P1_ADDR_REG_5__SCAN_IN), .A(n10699), .B(
        n10273), .ZN(n10279) );
  INV_X1 U12855 ( .A(n13973), .ZN(n10277) );
  NAND3_X1 U12856 ( .A1(n13958), .A2(n10275), .A3(n10274), .ZN(n10276) );
  NAND3_X1 U12857 ( .A1(n14752), .A2(n10277), .A3(n10276), .ZN(n10278) );
  OAI211_X1 U12858 ( .C1(n10280), .C2(n14036), .A(n10279), .B(n10278), .ZN(
        P1_U3248) );
  INV_X1 U12859 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14935) );
  MUX2_X1 U12860 ( .A(n14935), .B(P1_REG1_REG_9__SCAN_IN), .S(n10288), .Z(
        n10284) );
  AOI21_X1 U12861 ( .B1(n10284), .B2(n10283), .A(n10370), .ZN(n10296) );
  NOR2_X1 U12862 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13578), .ZN(n10286) );
  NOR2_X1 U12863 ( .A1(n13984), .A2(n10375), .ZN(n10285) );
  AOI211_X1 U12864 ( .C1(n13987), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10286), .B(
        n10285), .ZN(n10295) );
  NAND2_X1 U12865 ( .A1(n10287), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10290) );
  MUX2_X1 U12866 ( .A(n9162), .B(P1_REG2_REG_9__SCAN_IN), .S(n10288), .Z(
        n10289) );
  AOI21_X1 U12867 ( .B1(n10291), .B2(n10290), .A(n10289), .ZN(n13990) );
  INV_X1 U12868 ( .A(n13990), .ZN(n10293) );
  NAND3_X1 U12869 ( .A1(n10291), .A2(n10290), .A3(n10289), .ZN(n10292) );
  NAND3_X1 U12870 ( .A1(n10293), .A2(n14752), .A3(n10292), .ZN(n10294) );
  OAI211_X1 U12871 ( .C1(n10296), .C2(n14036), .A(n10295), .B(n10294), .ZN(
        P1_U3252) );
  INV_X1 U12872 ( .A(n15139), .ZN(n15124) );
  OAI21_X1 U12873 ( .B1(n10303), .B2(n10298), .A(n10297), .ZN(n10352) );
  OAI211_X1 U12874 ( .C1(n8841), .C2(n15042), .A(n15021), .B(n10328), .ZN(
        n10348) );
  OAI21_X1 U12875 ( .B1(n8841), .B2(n15146), .A(n10348), .ZN(n10309) );
  INV_X1 U12876 ( .A(n9597), .ZN(n10301) );
  OAI22_X1 U12877 ( .A1(n10301), .A2(n12884), .B1(n10300), .B2(n12886), .ZN(
        n11864) );
  NAND2_X1 U12878 ( .A1(n10303), .A2(n10302), .ZN(n10306) );
  INV_X1 U12879 ( .A(n10304), .ZN(n15039) );
  AOI21_X1 U12880 ( .B1(n10306), .B2(n10305), .A(n15039), .ZN(n10307) );
  AOI211_X1 U12881 ( .C1(n15143), .C2(n10352), .A(n11864), .B(n10307), .ZN(
        n10353) );
  INV_X1 U12882 ( .A(n10353), .ZN(n10308) );
  AOI211_X1 U12883 ( .C1(n15124), .C2(n10352), .A(n10309), .B(n10308), .ZN(
        n10343) );
  NAND2_X1 U12884 ( .A1(n15087), .A2(n10310), .ZN(n10311) );
  OR2_X1 U12885 ( .A1(n10312), .A2(n10311), .ZN(n10342) );
  NOR2_X4 U12886 ( .A1(n10342), .A2(n10313), .ZN(n15160) );
  NAND2_X1 U12887 ( .A1(n15164), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10314) );
  OAI21_X1 U12888 ( .B1(n10343), .B2(n15164), .A(n10314), .ZN(P2_U3500) );
  INV_X1 U12889 ( .A(n10315), .ZN(n10317) );
  AND2_X1 U12890 ( .A1(n10317), .A2(n10316), .ZN(n10453) );
  INV_X1 U12891 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n10324) );
  NAND2_X1 U12892 ( .A1(n10684), .A2(n14039), .ZN(n14824) );
  INV_X1 U12893 ( .A(n10319), .ZN(n14827) );
  OAI21_X1 U12894 ( .B1(n14922), .B2(n14766), .A(n14827), .ZN(n10322) );
  NAND2_X1 U12895 ( .A1(n14769), .A2(n13922), .ZN(n14822) );
  NAND2_X1 U12896 ( .A1(n10321), .A2(n10320), .ZN(n14821) );
  NAND3_X1 U12897 ( .A1(n10322), .A2(n14822), .A3(n14821), .ZN(n14422) );
  NAND2_X1 U12898 ( .A1(n14422), .A2(n14925), .ZN(n10323) );
  OAI21_X1 U12899 ( .B1(n14925), .B2(n10324), .A(n10323), .ZN(P1_U3459) );
  OAI21_X1 U12900 ( .B1(n10327), .B2(n10326), .A(n10325), .ZN(n10760) );
  INV_X1 U12901 ( .A(n10328), .ZN(n10330) );
  INV_X1 U12902 ( .A(n10329), .ZN(n10401) );
  OAI211_X1 U12903 ( .C1(n10331), .C2(n10330), .A(n10401), .B(n15021), .ZN(
        n10758) );
  OAI21_X1 U12904 ( .B1(n10331), .B2(n15146), .A(n10758), .ZN(n10338) );
  OAI21_X1 U12905 ( .B1(n10334), .B2(n10333), .A(n10332), .ZN(n10336) );
  AOI21_X1 U12906 ( .B1(n10336), .B2(n15018), .A(n10335), .ZN(n10762) );
  INV_X1 U12907 ( .A(n10762), .ZN(n10337) );
  AOI211_X1 U12908 ( .C1(n15151), .C2(n10760), .A(n10338), .B(n10337), .ZN(
        n15095) );
  NAND2_X1 U12909 ( .A1(n15164), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10339) );
  OAI21_X1 U12910 ( .B1(n15095), .B2(n15164), .A(n10339), .ZN(P2_U3501) );
  NAND2_X1 U12911 ( .A1(n14077), .A2(P1_U4016), .ZN(n10340) );
  OAI21_X1 U12912 ( .B1(P1_U4016), .B2(n10341), .A(n10340), .ZN(P1_U3583) );
  INV_X1 U12913 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10345) );
  OR2_X1 U12914 ( .A1(n10343), .A2(n15153), .ZN(n10344) );
  OAI21_X1 U12915 ( .B1(n15155), .B2(n10345), .A(n10344), .ZN(P2_U3433) );
  INV_X1 U12916 ( .A(n10346), .ZN(n10368) );
  INV_X1 U12917 ( .A(n14455), .ZN(n14444) );
  AOI22_X1 U12918 ( .A1(n14003), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n14444), .ZN(n10347) );
  OAI21_X1 U12919 ( .B1(n10368), .B2(n14458), .A(n10347), .ZN(P1_U3339) );
  NOR2_X1 U12920 ( .A1(n15023), .A2(n10348), .ZN(n10351) );
  OAI22_X1 U12921 ( .A1(n13236), .A2(n8841), .B1(n10349), .B2(n15050), .ZN(
        n10350) );
  AOI211_X1 U12922 ( .C1(n10651), .C2(n10352), .A(n10351), .B(n10350), .ZN(
        n10356) );
  MUX2_X1 U12923 ( .A(n10354), .B(n10353), .S(n15048), .Z(n10355) );
  NAND2_X1 U12924 ( .A1(n10356), .A2(n10355), .ZN(P2_U3264) );
  INV_X1 U12925 ( .A(n10357), .ZN(n10358) );
  OAI222_X1 U12926 ( .A1(P3_U3151), .A2(n12351), .B1(n14574), .B2(n10359), 
        .C1(n14576), .C2(n10358), .ZN(P3_U3278) );
  INV_X1 U12927 ( .A(n10360), .ZN(n10361) );
  AOI21_X1 U12928 ( .B1(n10363), .B2(n10362), .A(n10361), .ZN(n10367) );
  NAND2_X1 U12929 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n14972) );
  OAI22_X1 U12930 ( .A1(n7134), .A2(n12884), .B1(n10481), .B2(n12886), .ZN(
        n10413) );
  NAND2_X1 U12931 ( .A1(n12950), .A2(n10413), .ZN(n10364) );
  OAI211_X1 U12932 ( .C1(n12953), .C2(n10527), .A(n14972), .B(n10364), .ZN(
        n10365) );
  AOI21_X1 U12933 ( .B1(n10417), .B2(n8784), .A(n10365), .ZN(n10366) );
  OAI21_X1 U12934 ( .B1(n10367), .B2(n12938), .A(n10366), .ZN(P2_U3202) );
  INV_X1 U12935 ( .A(n13005), .ZN(n13011) );
  OAI222_X1 U12936 ( .A1(n13395), .A2(n10369), .B1(n13011), .B2(P2_U3088), 
        .C1(n13393), .C2(n10368), .ZN(P2_U3311) );
  INV_X1 U12937 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14693) );
  MUX2_X1 U12938 ( .A(n14693), .B(P1_REG1_REG_11__SCAN_IN), .S(n10562), .Z(
        n10372) );
  INV_X1 U12939 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14938) );
  MUX2_X1 U12940 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n14938), .S(n10377), .Z(
        n13980) );
  NAND2_X1 U12941 ( .A1(n13981), .A2(n13980), .ZN(n13979) );
  AOI21_X1 U12942 ( .B1(n10372), .B2(n10371), .A(n14747), .ZN(n10384) );
  AND2_X1 U12943 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n11506) );
  NOR2_X1 U12944 ( .A1(n13984), .A2(n10373), .ZN(n10374) );
  AOI211_X1 U12945 ( .C1(n13987), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n11506), 
        .B(n10374), .ZN(n10383) );
  NOR2_X1 U12946 ( .A1(n10375), .A2(n9162), .ZN(n13989) );
  MUX2_X1 U12947 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10376), .S(n10377), .Z(
        n13988) );
  OAI21_X1 U12948 ( .B1(n13990), .B2(n13989), .A(n13988), .ZN(n13992) );
  NAND2_X1 U12949 ( .A1(n10377), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10379) );
  MUX2_X1 U12950 ( .A(n9201), .B(P1_REG2_REG_11__SCAN_IN), .S(n10562), .Z(
        n10378) );
  AOI21_X1 U12951 ( .B1(n13992), .B2(n10379), .A(n10378), .ZN(n10561) );
  INV_X1 U12952 ( .A(n10561), .ZN(n10381) );
  NAND3_X1 U12953 ( .A1(n13992), .A2(n10379), .A3(n10378), .ZN(n10380) );
  NAND3_X1 U12954 ( .A1(n10381), .A2(n14752), .A3(n10380), .ZN(n10382) );
  OAI211_X1 U12955 ( .C1(n10384), .C2(n14036), .A(n10383), .B(n10382), .ZN(
        P1_U3254) );
  INV_X1 U12956 ( .A(n11029), .ZN(n11026) );
  INV_X1 U12957 ( .A(n10385), .ZN(n10389) );
  OAI222_X1 U12958 ( .A1(P1_U3086), .A2(n11026), .B1(n14458), .B2(n10389), 
        .C1(n10386), .C2(n14455), .ZN(P1_U3341) );
  NAND2_X1 U12959 ( .A1(n12913), .A2(P2_U3947), .ZN(n10387) );
  OAI21_X1 U12960 ( .B1(n10388), .B2(P2_U3947), .A(n10387), .ZN(P2_U3554) );
  INV_X1 U12961 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10390) );
  INV_X1 U12962 ( .A(n11658), .ZN(n11151) );
  OAI222_X1 U12963 ( .A1(n13395), .A2(n10390), .B1(n11151), .B2(P2_U3088), 
        .C1(n13393), .C2(n10389), .ZN(P2_U3313) );
  OAI21_X1 U12964 ( .B1(n10393), .B2(n10392), .A(n10391), .ZN(n10394) );
  INV_X1 U12965 ( .A(n10394), .ZN(n10438) );
  OAI21_X1 U12966 ( .B1(n10397), .B2(n10396), .A(n10395), .ZN(n10399) );
  AOI21_X1 U12967 ( .B1(n10399), .B2(n15018), .A(n10398), .ZN(n10400) );
  OAI21_X1 U12968 ( .B1(n10438), .B2(n15119), .A(n10400), .ZN(n10429) );
  INV_X1 U12969 ( .A(n10429), .ZN(n10403) );
  AOI211_X1 U12970 ( .C1(n10433), .C2(n10401), .A(n13219), .B(n10415), .ZN(
        n10434) );
  AOI21_X1 U12971 ( .B1(n15137), .B2(n10433), .A(n10434), .ZN(n10402) );
  OAI211_X1 U12972 ( .C1(n10438), .C2(n15139), .A(n10403), .B(n10402), .ZN(
        n10439) );
  NAND2_X1 U12973 ( .A1(n10439), .A2(n15155), .ZN(n10404) );
  OAI21_X1 U12974 ( .B1(n15155), .B2(n8235), .A(n10404), .ZN(P2_U3439) );
  INV_X1 U12975 ( .A(n12378), .ZN(n12382) );
  INV_X1 U12976 ( .A(n10405), .ZN(n10406) );
  OAI222_X1 U12977 ( .A1(P3_U3151), .A2(n12382), .B1(n14574), .B2(n13617), 
        .C1(n14576), .C2(n10406), .ZN(P3_U3277) );
  OAI21_X1 U12978 ( .B1(n10409), .B2(n10408), .A(n10407), .ZN(n10410) );
  INV_X1 U12979 ( .A(n10410), .ZN(n10533) );
  XNOR2_X1 U12980 ( .A(n10412), .B(n10411), .ZN(n10414) );
  AOI21_X1 U12981 ( .B1(n10414), .B2(n15018), .A(n10413), .ZN(n10526) );
  OAI21_X1 U12982 ( .B1(n10528), .B2(n10415), .A(n15021), .ZN(n10416) );
  NOR2_X1 U12983 ( .A1(n10416), .A2(n10637), .ZN(n10530) );
  AOI21_X1 U12984 ( .B1(n15137), .B2(n10417), .A(n10530), .ZN(n10418) );
  OAI211_X1 U12985 ( .C1(n10533), .C2(n13351), .A(n10526), .B(n10418), .ZN(
        n10441) );
  NAND2_X1 U12986 ( .A1(n10441), .A2(n15155), .ZN(n10419) );
  OAI21_X1 U12987 ( .B1(n15155), .B2(n8255), .A(n10419), .ZN(P2_U3442) );
  INV_X1 U12988 ( .A(n10420), .ZN(n10444) );
  OAI222_X1 U12989 ( .A1(n13393), .A2(n10444), .B1(n15013), .B2(P2_U3088), 
        .C1(n13634), .C2(n13395), .ZN(P2_U3312) );
  INV_X1 U12990 ( .A(n10421), .ZN(n10445) );
  INV_X1 U12991 ( .A(n13024), .ZN(n13018) );
  OAI222_X1 U12992 ( .A1(n13393), .A2(n10445), .B1(n13018), .B2(P2_U3088), 
        .C1(n10422), .C2(n13395), .ZN(P2_U3310) );
  XOR2_X1 U12993 ( .A(n10423), .B(n10424), .Z(n10428) );
  INV_X1 U12994 ( .A(n14660), .ZN(n11507) );
  AOI22_X1 U12995 ( .A1(n11507), .A2(n13921), .B1(n13901), .B2(n9943), .ZN(
        n10427) );
  NAND2_X1 U12996 ( .A1(n14725), .A2(n10425), .ZN(n10462) );
  AOI22_X1 U12997 ( .A1(n13905), .A2(n9027), .B1(n10462), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10426) );
  OAI211_X1 U12998 ( .C1(n10428), .C2(n13908), .A(n10427), .B(n10426), .ZN(
        P1_U3222) );
  INV_X1 U12999 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10430) );
  AOI21_X1 U13000 ( .B1(n13254), .B2(n10430), .A(n10429), .ZN(n10431) );
  MUX2_X1 U13001 ( .A(n10432), .B(n10431), .S(n15048), .Z(n10436) );
  AOI22_X1 U13002 ( .A1(n10434), .A2(n13259), .B1(n15027), .B2(n10433), .ZN(
        n10435) );
  OAI211_X1 U13003 ( .C1(n10438), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        P2_U3262) );
  NAND2_X1 U13004 ( .A1(n10439), .A2(n15160), .ZN(n10440) );
  OAI21_X1 U13005 ( .B1(n15160), .B2(n10064), .A(n10440), .ZN(P2_U3502) );
  NAND2_X1 U13006 ( .A1(n10441), .A2(n15160), .ZN(n10442) );
  OAI21_X1 U13007 ( .B1(n15160), .B2(n10066), .A(n10442), .ZN(P2_U3503) );
  OAI222_X1 U13008 ( .A1(P1_U3086), .A2(n11313), .B1(n14458), .B2(n10444), 
        .C1(n10443), .C2(n14455), .ZN(P1_U3340) );
  INV_X1 U13009 ( .A(n14012), .ZN(n14019) );
  OAI222_X1 U13010 ( .A1(P1_U3086), .A2(n14019), .B1(n14458), .B2(n10445), 
        .C1(n13502), .C2(n14455), .ZN(P1_U3338) );
  OAI222_X1 U13011 ( .A1(n14576), .A2(n10447), .B1(n14574), .B2(n10446), .C1(
        P3_U3151), .C2(n12391), .ZN(P3_U3276) );
  INV_X1 U13012 ( .A(n14401), .ZN(n14916) );
  OAI21_X1 U13013 ( .B1(n10862), .B2(n14920), .A(n10448), .ZN(n10450) );
  AOI211_X1 U13014 ( .C1(n14916), .C2(n10451), .A(n10450), .B(n10449), .ZN(
        n14866) );
  NAND2_X1 U13015 ( .A1(n14937), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10454) );
  OAI21_X1 U13016 ( .B1(n14866), .B2(n14937), .A(n10454), .ZN(P1_U3529) );
  INV_X1 U13017 ( .A(n13905), .ZN(n14659) );
  INV_X1 U13018 ( .A(n14733), .ZN(n13832) );
  OAI22_X1 U13019 ( .A1(n10455), .A2(n13908), .B1(n13832), .B2(n14822), .ZN(
        n10456) );
  AOI21_X1 U13020 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n10462), .A(n10456), .ZN(
        n10457) );
  OAI21_X1 U13021 ( .B1(n10458), .B2(n14659), .A(n10457), .ZN(P1_U3232) );
  XNOR2_X1 U13022 ( .A(n10459), .B(n10460), .ZN(n10461) );
  NAND2_X1 U13023 ( .A1(n10461), .A2(n14726), .ZN(n10464) );
  INV_X1 U13024 ( .A(n13920), .ZN(n10890) );
  OAI22_X1 U13025 ( .A1(n10890), .A2(n14240), .B1(n9028), .B2(n14288), .ZN(
        n14806) );
  AOI22_X1 U13026 ( .A1(n10462), .A2(P1_REG3_REG_2__SCAN_IN), .B1(n14733), 
        .B2(n14806), .ZN(n10463) );
  OAI211_X1 U13027 ( .C1(n9043), .C2(n14659), .A(n10464), .B(n10463), .ZN(
        P1_U3237) );
  OAI21_X1 U13028 ( .B1(n10467), .B2(n10466), .A(n10465), .ZN(n10468) );
  NAND2_X1 U13029 ( .A1(n10468), .A2(n12946), .ZN(n10476) );
  OR2_X1 U13030 ( .A1(n10469), .A2(n12886), .ZN(n10472) );
  OR2_X1 U13031 ( .A1(n10470), .A2(n12884), .ZN(n10471) );
  NAND2_X1 U13032 ( .A1(n10472), .A2(n10471), .ZN(n10645) );
  NOR2_X1 U13033 ( .A1(n12953), .A2(n10638), .ZN(n10473) );
  AOI211_X1 U13034 ( .C1(n12950), .C2(n10645), .A(n10474), .B(n10473), .ZN(
        n10475) );
  OAI211_X1 U13035 ( .C1(n15098), .C2(n12926), .A(n10476), .B(n10475), .ZN(
        P2_U3199) );
  INV_X1 U13036 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n13481) );
  NAND2_X1 U13037 ( .A1(n12618), .A2(P3_U3897), .ZN(n10477) );
  OAI21_X1 U13038 ( .B1(P3_U3897), .B2(n13481), .A(n10477), .ZN(P3_U3504) );
  XNOR2_X1 U13039 ( .A(n10478), .B(n10479), .ZN(n10488) );
  INV_X1 U13040 ( .A(n10480), .ZN(n13253) );
  OR2_X1 U13041 ( .A1(n10708), .A2(n12886), .ZN(n10483) );
  OR2_X1 U13042 ( .A1(n10481), .A2(n12884), .ZN(n10482) );
  AND2_X1 U13043 ( .A1(n10483), .A2(n10482), .ZN(n13249) );
  OAI21_X1 U13044 ( .B1(n12937), .B2(n13249), .A(n10484), .ZN(n10485) );
  AOI21_X1 U13045 ( .B1(n13253), .B2(n12935), .A(n10485), .ZN(n10487) );
  NAND2_X1 U13046 ( .A1(n8784), .A2(n15106), .ZN(n10486) );
  OAI211_X1 U13047 ( .C1(n10488), .C2(n12938), .A(n10487), .B(n10486), .ZN(
        P2_U3211) );
  OAI21_X1 U13048 ( .B1(n10495), .B2(P2_REG2_REG_9__SCAN_IN), .A(n10489), .ZN(
        n14994) );
  MUX2_X1 U13049 ( .A(n8372), .B(P2_REG2_REG_10__SCAN_IN), .S(n14990), .Z(
        n14995) );
  NOR2_X1 U13050 ( .A1(n14994), .A2(n14995), .ZN(n14992) );
  AOI21_X1 U13051 ( .B1(n14990), .B2(P2_REG2_REG_10__SCAN_IN), .A(n14992), 
        .ZN(n10491) );
  MUX2_X1 U13052 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n8392), .S(n10541), .Z(
        n10490) );
  NAND2_X1 U13053 ( .A1(n10491), .A2(n10490), .ZN(n10548) );
  OAI21_X1 U13054 ( .B1(n10491), .B2(n10490), .A(n10548), .ZN(n10502) );
  AND2_X1 U13055 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10492) );
  AOI21_X1 U13056 ( .B1(n15007), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10492), 
        .ZN(n10493) );
  OAI21_X1 U13057 ( .B1(n10544), .B2(n15014), .A(n10493), .ZN(n10501) );
  OAI21_X1 U13058 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10495), .A(n10494), .ZN(
        n14986) );
  MUX2_X1 U13059 ( .A(n10496), .B(P2_REG1_REG_10__SCAN_IN), .S(n14990), .Z(
        n14987) );
  NOR2_X1 U13060 ( .A1(n14986), .A2(n14987), .ZN(n14985) );
  MUX2_X1 U13061 ( .A(n10497), .B(P2_REG1_REG_11__SCAN_IN), .S(n10541), .Z(
        n10498) );
  AOI211_X1 U13062 ( .C1(n10499), .C2(n10498), .A(n15001), .B(n10540), .ZN(
        n10500) );
  AOI211_X1 U13063 ( .C1(n15009), .C2(n10502), .A(n10501), .B(n10500), .ZN(
        n10503) );
  INV_X1 U13064 ( .A(n10503), .ZN(P2_U3225) );
  NAND2_X1 U13065 ( .A1(n12696), .A2(n10751), .ZN(n12073) );
  INV_X1 U13066 ( .A(n12073), .ZN(n10504) );
  NOR2_X1 U13067 ( .A1(n12701), .A2(n10504), .ZN(n12045) );
  NAND2_X1 U13068 ( .A1(n10516), .A2(n15406), .ZN(n10675) );
  OAI22_X1 U13069 ( .A1(n10517), .A2(n10675), .B1(n10826), .B2(n10512), .ZN(
        n10505) );
  INV_X1 U13070 ( .A(n10827), .ZN(n10507) );
  NAND2_X1 U13071 ( .A1(n15319), .A2(n10507), .ZN(n10508) );
  NAND2_X1 U13072 ( .A1(n10517), .A2(n15363), .ZN(n10510) );
  NAND2_X1 U13073 ( .A1(n10574), .A2(n14625), .ZN(n10748) );
  INV_X1 U13074 ( .A(n10748), .ZN(n10509) );
  AOI22_X1 U13075 ( .A1(n10506), .A2(n12005), .B1(n12018), .B2(n10511), .ZN(
        n10525) );
  INV_X1 U13076 ( .A(n10512), .ZN(n10515) );
  NAND3_X1 U13077 ( .A1(n10513), .A2(n10575), .A3(n10746), .ZN(n10514) );
  AOI21_X1 U13078 ( .B1(n10826), .B2(n10515), .A(n10514), .ZN(n10519) );
  NAND2_X1 U13079 ( .A1(n10517), .A2(n10516), .ZN(n10518) );
  NAND2_X1 U13080 ( .A1(n10519), .A2(n10518), .ZN(n10520) );
  NAND2_X1 U13081 ( .A1(n10520), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10523) );
  NAND2_X1 U13082 ( .A1(n10521), .A2(n10826), .ZN(n10522) );
  NAND2_X1 U13083 ( .A1(n11985), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10961) );
  NAND2_X1 U13084 ( .A1(n10961), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10524) );
  OAI211_X1 U13085 ( .C1(n12045), .C2(n12014), .A(n10525), .B(n10524), .ZN(
        P3_U3172) );
  MUX2_X1 U13086 ( .A(n10075), .B(n10526), .S(n15048), .Z(n10532) );
  OAI22_X1 U13087 ( .A1(n13236), .A2(n10528), .B1(n15050), .B2(n10527), .ZN(
        n10529) );
  AOI21_X1 U13088 ( .B1(n13259), .B2(n10530), .A(n10529), .ZN(n10531) );
  OAI211_X1 U13089 ( .C1(n13246), .C2(n10533), .A(n10532), .B(n10531), .ZN(
        P2_U3261) );
  INV_X1 U13090 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n13504) );
  INV_X1 U13091 ( .A(n12572), .ZN(n12537) );
  NAND2_X1 U13092 ( .A1(n12537), .A2(P3_U3897), .ZN(n10534) );
  OAI21_X1 U13093 ( .B1(P3_U3897), .B2(n13504), .A(n10534), .ZN(P3_U3509) );
  INV_X1 U13094 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U13095 ( .A1(n12484), .A2(P3_U3897), .ZN(n10535) );
  OAI21_X1 U13096 ( .B1(P3_U3897), .B2(n13565), .A(n10535), .ZN(P3_U3515) );
  INV_X1 U13097 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U13098 ( .A1(n11982), .A2(P3_U3897), .ZN(n10536) );
  OAI21_X1 U13099 ( .B1(P3_U3897), .B2(n13465), .A(n10536), .ZN(P3_U3505) );
  INV_X1 U13100 ( .A(n13033), .ZN(n13037) );
  OAI222_X1 U13101 ( .A1(n13393), .A2(n10538), .B1(n13037), .B2(P2_U3088), 
        .C1(n10537), .C2(n13395), .ZN(P2_U3309) );
  INV_X1 U13102 ( .A(n14031), .ZN(n14024) );
  OAI222_X1 U13103 ( .A1(P1_U3086), .A2(n14024), .B1(n14458), .B2(n10538), 
        .C1(n13629), .C2(n14455), .ZN(P1_U3337) );
  XNOR2_X1 U13104 ( .A(n10796), .B(n10539), .ZN(n10543) );
  OAI21_X1 U13105 ( .B1(n10543), .B2(n10542), .A(n10795), .ZN(n10554) );
  NAND2_X1 U13106 ( .A1(n10544), .A2(n8392), .ZN(n10546) );
  INV_X1 U13107 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10545) );
  MUX2_X1 U13108 ( .A(n10545), .B(P2_REG2_REG_12__SCAN_IN), .S(n10796), .Z(
        n10547) );
  AOI21_X1 U13109 ( .B1(n10548), .B2(n10546), .A(n10547), .ZN(n10800) );
  AND3_X1 U13110 ( .A1(n10548), .A2(n10547), .A3(n10546), .ZN(n10549) );
  OAI21_X1 U13111 ( .B1(n10800), .B2(n10549), .A(n15009), .ZN(n10552) );
  NOR2_X1 U13112 ( .A1(n10550), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11358) );
  AOI21_X1 U13113 ( .B1(n15007), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n11358), 
        .ZN(n10551) );
  OAI211_X1 U13114 ( .C1(n15014), .C2(n10801), .A(n10552), .B(n10551), .ZN(
        n10553) );
  AOI21_X1 U13115 ( .B1(n10554), .B2(n14976), .A(n10553), .ZN(n10555) );
  INV_X1 U13116 ( .A(n10555), .ZN(P2_U3226) );
  INV_X1 U13117 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n13549) );
  NAND2_X1 U13118 ( .A1(n12470), .A2(P3_U3897), .ZN(n10556) );
  OAI21_X1 U13119 ( .B1(P3_U3897), .B2(n13549), .A(n10556), .ZN(P3_U3516) );
  NOR2_X1 U13120 ( .A1(n10562), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n14742) );
  MUX2_X1 U13121 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n14741), .S(n14751), .Z(
        n10557) );
  INV_X1 U13122 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10558) );
  MUX2_X1 U13123 ( .A(n10558), .B(P1_REG1_REG_13__SCAN_IN), .S(n10724), .Z(
        n10559) );
  NOR2_X1 U13124 ( .A1(n10560), .A2(n10559), .ZN(n10723) );
  AOI211_X1 U13125 ( .C1(n10560), .C2(n10559), .A(n10723), .B(n14036), .ZN(
        n10572) );
  AOI21_X1 U13126 ( .B1(n10562), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10561), 
        .ZN(n14739) );
  MUX2_X1 U13127 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9217), .S(n14751), .Z(
        n14740) );
  AND2_X1 U13128 ( .A1(n14739), .A2(n14740), .ZN(n14737) );
  NOR2_X1 U13129 ( .A1(n14751), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10563) );
  NOR2_X1 U13130 ( .A1(n14737), .A2(n10563), .ZN(n10566) );
  MUX2_X1 U13131 ( .A(n9247), .B(P1_REG2_REG_13__SCAN_IN), .S(n10724), .Z(
        n10564) );
  INV_X1 U13132 ( .A(n10564), .ZN(n10565) );
  NAND2_X1 U13133 ( .A1(n10565), .A2(n10566), .ZN(n10718) );
  OAI211_X1 U13134 ( .C1(n10566), .C2(n10565), .A(n14752), .B(n10718), .ZN(
        n10569) );
  INV_X1 U13135 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n13863) );
  NOR2_X1 U13136 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13863), .ZN(n10567) );
  AOI21_X1 U13137 ( .B1(n13987), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10567), 
        .ZN(n10568) );
  OAI211_X1 U13138 ( .C1(n13984), .C2(n10570), .A(n10569), .B(n10568), .ZN(
        n10571) );
  OR2_X1 U13139 ( .A1(n10572), .A2(n10571), .ZN(P1_U3256) );
  OR2_X1 U13140 ( .A1(n10575), .A2(P3_U3151), .ZN(n12246) );
  INV_X1 U13141 ( .A(n12246), .ZN(n10573) );
  NAND2_X1 U13142 ( .A1(n12227), .A2(n10575), .ZN(n10576) );
  AND2_X1 U13143 ( .A1(n10577), .A2(n10576), .ZN(n10587) );
  AND2_X1 U13144 ( .A1(n10588), .A2(n10587), .ZN(n10582) );
  INV_X1 U13145 ( .A(n10582), .ZN(n10578) );
  MUX2_X1 U13146 ( .A(n12259), .B(n10578), .S(n11819), .Z(n15290) );
  INV_X1 U13147 ( .A(n15290), .ZN(n15181) );
  INV_X1 U13148 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n15413) );
  XNOR2_X1 U13149 ( .A(n6552), .B(n15413), .ZN(n11120) );
  NAND2_X1 U13150 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n13500), .ZN(n10787) );
  INV_X1 U13151 ( .A(n10787), .ZN(n10579) );
  INV_X1 U13152 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13153 ( .A1(n10619), .A2(n7433), .ZN(n11118) );
  XNOR2_X1 U13154 ( .A(n11120), .B(n11118), .ZN(n10592) );
  NAND2_X1 U13155 ( .A1(n10582), .A2(n12774), .ZN(n12387) );
  INV_X1 U13156 ( .A(n10580), .ZN(n10581) );
  INV_X1 U13157 ( .A(n15300), .ZN(n12366) );
  INV_X1 U13158 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10599) );
  OAI21_X1 U13159 ( .B1(n6546), .B2(n10782), .A(n10583), .ZN(n10614) );
  OR2_X1 U13160 ( .A1(n10614), .A2(n10593), .ZN(n10616) );
  NAND2_X1 U13161 ( .A1(n10616), .A2(n10583), .ZN(n10584) );
  OAI21_X1 U13162 ( .B1(n10585), .B2(n10584), .A(n11061), .ZN(n10586) );
  NAND2_X1 U13163 ( .A1(n12366), .A2(n10586), .ZN(n10591) );
  INV_X1 U13164 ( .A(n10587), .ZN(n10589) );
  AOI22_X1 U13165 ( .A1(n15293), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10590) );
  OAI211_X1 U13166 ( .C1(n10592), .C2(n12387), .A(n10591), .B(n10590), .ZN(
        n10609) );
  INV_X1 U13167 ( .A(n6546), .ZN(n10626) );
  NAND2_X1 U13168 ( .A1(n10594), .A2(n10626), .ZN(n10605) );
  NAND2_X1 U13169 ( .A1(n10596), .A2(n6546), .ZN(n10597) );
  NAND2_X1 U13170 ( .A1(n10605), .A2(n10597), .ZN(n10611) );
  INV_X1 U13171 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10598) );
  MUX2_X1 U13172 ( .A(n10599), .B(n10598), .S(n12774), .Z(n10788) );
  MUX2_X1 U13173 ( .A(n10600), .B(n15413), .S(n12774), .Z(n10601) );
  NAND2_X1 U13174 ( .A1(n10601), .A2(n6552), .ZN(n11077) );
  INV_X1 U13175 ( .A(n10601), .ZN(n10602) );
  INV_X1 U13176 ( .A(n6552), .ZN(n11059) );
  NAND2_X1 U13177 ( .A1(n10602), .A2(n11059), .ZN(n10603) );
  NAND2_X1 U13178 ( .A1(n11077), .A2(n10603), .ZN(n10604) );
  AOI21_X1 U13179 ( .B1(n10613), .B2(n10605), .A(n10604), .ZN(n15175) );
  INV_X1 U13180 ( .A(n15175), .ZN(n10607) );
  NAND3_X1 U13181 ( .A1(n10613), .A2(n10605), .A3(n10604), .ZN(n10606) );
  INV_X1 U13182 ( .A(n11819), .ZN(n12241) );
  AOI21_X1 U13183 ( .B1(n10607), .B2(n10606), .A(n15176), .ZN(n10608) );
  AOI211_X1 U13184 ( .C1(n15181), .C2(n6552), .A(n10609), .B(n10608), .ZN(
        n10610) );
  INV_X1 U13185 ( .A(n10610), .ZN(P3_U3184) );
  NAND2_X1 U13186 ( .A1(n10611), .A2(n10781), .ZN(n10612) );
  AOI21_X1 U13187 ( .B1(n10613), .B2(n10612), .A(n15176), .ZN(n10625) );
  NAND2_X1 U13188 ( .A1(n10614), .A2(n10593), .ZN(n10615) );
  AND2_X1 U13189 ( .A1(n10616), .A2(n10615), .ZN(n10623) );
  AOI22_X1 U13190 ( .A1(n15293), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10622) );
  NAND2_X1 U13191 ( .A1(n10619), .A2(n10618), .ZN(n10620) );
  NAND2_X1 U13192 ( .A1(n15296), .A2(n10620), .ZN(n10621) );
  OAI211_X1 U13193 ( .C1(n10623), .C2(n15300), .A(n10622), .B(n10621), .ZN(
        n10624) );
  AOI211_X1 U13194 ( .C1(n15181), .C2(n10626), .A(n10625), .B(n10624), .ZN(
        n10627) );
  INV_X1 U13195 ( .A(n10627), .ZN(P3_U3183) );
  XNOR2_X1 U13196 ( .A(n10629), .B(n10628), .ZN(n10634) );
  AOI22_X1 U13197 ( .A1(n12932), .A2(n12982), .B1(n12933), .B2(n12980), .ZN(
        n10657) );
  OAI22_X1 U13198 ( .A1(n12937), .A2(n10657), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8318), .ZN(n10631) );
  NOR2_X1 U13199 ( .A1(n12953), .A2(n10661), .ZN(n10630) );
  AOI211_X1 U13200 ( .C1(n10632), .C2(n8784), .A(n10631), .B(n10630), .ZN(
        n10633) );
  OAI21_X1 U13201 ( .B1(n10634), .B2(n12938), .A(n10633), .ZN(P2_U3185) );
  XNOR2_X1 U13202 ( .A(n10636), .B(n10635), .ZN(n15096) );
  OAI211_X1 U13203 ( .C1(n15098), .C2(n10637), .A(n15021), .B(n13258), .ZN(
        n15097) );
  INV_X1 U13204 ( .A(n10638), .ZN(n10639) );
  AOI22_X1 U13205 ( .A1(n15027), .A2(n10640), .B1(n10639), .B2(n13254), .ZN(
        n10641) );
  OAI21_X1 U13206 ( .B1(n15023), .B2(n15097), .A(n10641), .ZN(n10650) );
  NAND2_X1 U13207 ( .A1(n15096), .A2(n15143), .ZN(n10648) );
  OAI21_X1 U13208 ( .B1(n10644), .B2(n10643), .A(n10642), .ZN(n10646) );
  AOI21_X1 U13209 ( .B1(n10646), .B2(n15018), .A(n10645), .ZN(n10647) );
  NAND2_X1 U13210 ( .A1(n10648), .A2(n10647), .ZN(n15101) );
  MUX2_X1 U13211 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n15101), .S(n15048), .Z(
        n10649) );
  AOI211_X1 U13212 ( .C1(n10651), .C2(n15096), .A(n10650), .B(n10649), .ZN(
        n10652) );
  INV_X1 U13213 ( .A(n10652), .ZN(P2_U3260) );
  OAI21_X1 U13214 ( .B1(n10654), .B2(n10655), .A(n10653), .ZN(n15110) );
  XNOR2_X1 U13215 ( .A(n10656), .B(n10655), .ZN(n10658) );
  OAI21_X1 U13216 ( .B1(n10658), .B2(n15039), .A(n10657), .ZN(n15113) );
  INV_X1 U13217 ( .A(n15113), .ZN(n10659) );
  MUX2_X1 U13218 ( .A(n10660), .B(n10659), .S(n15048), .Z(n10665) );
  OAI211_X1 U13219 ( .C1(n15112), .C2(n13257), .A(n15021), .B(n10773), .ZN(
        n15111) );
  INV_X1 U13220 ( .A(n15111), .ZN(n10663) );
  OAI22_X1 U13221 ( .A1(n15112), .A2(n13236), .B1(n10661), .B2(n15050), .ZN(
        n10662) );
  AOI21_X1 U13222 ( .B1(n10663), .B2(n13259), .A(n10662), .ZN(n10664) );
  OAI211_X1 U13223 ( .C1(n13246), .C2(n15110), .A(n10665), .B(n10664), .ZN(
        P2_U3258) );
  NOR2_X1 U13224 ( .A1(n14920), .A2(n10943), .ZN(n14880) );
  NAND2_X1 U13225 ( .A1(n14769), .A2(n13918), .ZN(n10667) );
  NAND2_X1 U13226 ( .A1(n14771), .A2(n13920), .ZN(n10666) );
  NAND2_X1 U13227 ( .A1(n10667), .A2(n10666), .ZN(n14878) );
  AND2_X1 U13228 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13950) );
  AOI21_X1 U13229 ( .B1(n14733), .B2(n14878), .A(n13950), .ZN(n10668) );
  OAI21_X1 U13230 ( .B1(n14736), .B2(n10944), .A(n10668), .ZN(n10673) );
  AOI211_X1 U13231 ( .C1(n10671), .C2(n10670), .A(n13908), .B(n10669), .ZN(
        n10672) );
  AOI211_X1 U13232 ( .C1(n14725), .C2(n14880), .A(n10673), .B(n10672), .ZN(
        n10674) );
  INV_X1 U13233 ( .A(n10674), .ZN(P1_U3230) );
  AND2_X1 U13234 ( .A1(n10675), .A2(n15347), .ZN(n10676) );
  OR2_X1 U13235 ( .A1(n12045), .A2(n10676), .ZN(n10678) );
  NAND2_X1 U13236 ( .A1(n10506), .A2(n15319), .ZN(n10677) );
  NAND2_X1 U13237 ( .A1(n10678), .A2(n10677), .ZN(n10749) );
  OAI22_X1 U13238 ( .A1(n12694), .A2(n10751), .B1(n15424), .B2(n10598), .ZN(
        n10679) );
  AOI21_X1 U13239 ( .B1(n10749), .B2(n15424), .A(n10679), .ZN(n10680) );
  INV_X1 U13240 ( .A(n10680), .ZN(P3_U3459) );
  OAI222_X1 U13241 ( .A1(n13393), .A2(n10683), .B1(n6555), .B2(P2_U3088), .C1(
        n10681), .C2(n13395), .ZN(P2_U3307) );
  OAI222_X1 U13242 ( .A1(n10684), .A2(P1_U3086), .B1(n14458), .B2(n10683), 
        .C1(n10682), .C2(n14455), .ZN(P1_U3335) );
  INV_X1 U13243 ( .A(n10685), .ZN(n10688) );
  OAI222_X1 U13244 ( .A1(P1_U3086), .A2(n10687), .B1(n14458), .B2(n10688), 
        .C1(n10686), .C2(n14455), .ZN(P1_U3336) );
  OAI222_X1 U13245 ( .A1(n13395), .A2(n13526), .B1(n13393), .B2(n10688), .C1(
        P2_U3088), .C2(n13047), .ZN(P2_U3308) );
  INV_X1 U13246 ( .A(n10689), .ZN(n10691) );
  OAI222_X1 U13247 ( .A1(P3_U3151), .A2(n10692), .B1(n14576), .B2(n10691), 
        .C1(n10690), .C2(n14574), .ZN(P3_U3275) );
  INV_X1 U13248 ( .A(n14725), .ZN(n13848) );
  NAND2_X1 U13249 ( .A1(n10921), .A2(n14722), .ZN(n14886) );
  XNOR2_X1 U13250 ( .A(n10694), .B(n7379), .ZN(n10695) );
  XNOR2_X1 U13251 ( .A(n10693), .B(n10695), .ZN(n10696) );
  NAND2_X1 U13252 ( .A1(n10696), .A2(n14726), .ZN(n10703) );
  INV_X1 U13253 ( .A(n10697), .ZN(n10922) );
  NAND2_X1 U13254 ( .A1(n14769), .A2(n13917), .ZN(n10698) );
  OAI21_X1 U13255 ( .B1(n10886), .B2(n14288), .A(n10698), .ZN(n10918) );
  AOI21_X1 U13256 ( .B1(n14733), .B2(n10918), .A(n10699), .ZN(n10700) );
  OAI21_X1 U13257 ( .B1(n14736), .B2(n10922), .A(n10700), .ZN(n10701) );
  INV_X1 U13258 ( .A(n10701), .ZN(n10702) );
  OAI211_X1 U13259 ( .C1(n13848), .C2(n14886), .A(n10703), .B(n10702), .ZN(
        P1_U3227) );
  XNOR2_X1 U13260 ( .A(n8337), .B(n10705), .ZN(n10706) );
  XNOR2_X1 U13261 ( .A(n10707), .B(n10706), .ZN(n10714) );
  OR2_X1 U13262 ( .A1(n10837), .A2(n12886), .ZN(n10710) );
  OR2_X1 U13263 ( .A1(n10708), .A2(n12884), .ZN(n10709) );
  NAND2_X1 U13264 ( .A1(n10710), .A2(n10709), .ZN(n10768) );
  AOI22_X1 U13265 ( .A1(n12950), .A2(n10768), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10711) );
  OAI21_X1 U13266 ( .B1(n12953), .B2(n10776), .A(n10711), .ZN(n10712) );
  AOI21_X1 U13267 ( .B1(n15116), .B2(n8784), .A(n10712), .ZN(n10713) );
  OAI21_X1 U13268 ( .B1(n10714), .B2(n12938), .A(n10713), .ZN(P2_U3193) );
  NAND2_X1 U13269 ( .A1(n12259), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n10715) );
  OAI21_X1 U13270 ( .B1(n12037), .B2(n12259), .A(n10715), .ZN(P3_U3521) );
  OAI22_X1 U13271 ( .A1(n10751), .A2(n12762), .B1(n15411), .B2(n7509), .ZN(
        n10716) );
  AOI21_X1 U13272 ( .B1(n10749), .B2(n15411), .A(n10716), .ZN(n10717) );
  INV_X1 U13273 ( .A(n10717), .ZN(P3_U3390) );
  NAND2_X1 U13274 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10724), .ZN(n10719) );
  NAND2_X1 U13275 ( .A1(n10719), .A2(n10718), .ZN(n10721) );
  MUX2_X1 U13276 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n11287), .S(n11029), .Z(
        n10720) );
  NAND2_X1 U13277 ( .A1(n10720), .A2(n10721), .ZN(n11025) );
  OAI211_X1 U13278 ( .C1(n10721), .C2(n10720), .A(n14752), .B(n11025), .ZN(
        n10732) );
  INV_X1 U13279 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10722) );
  MUX2_X1 U13280 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10722), .S(n11029), .Z(
        n10726) );
  AOI21_X1 U13281 ( .B1(n10724), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10723), 
        .ZN(n10725) );
  NAND2_X1 U13282 ( .A1(n10726), .A2(n10725), .ZN(n11028) );
  OAI21_X1 U13283 ( .B1(n10726), .B2(n10725), .A(n11028), .ZN(n10730) );
  NAND2_X1 U13284 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14667)
         );
  INV_X1 U13285 ( .A(n14667), .ZN(n10727) );
  AOI21_X1 U13286 ( .B1(n13987), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10727), 
        .ZN(n10728) );
  OAI21_X1 U13287 ( .B1(n13984), .B2(n11026), .A(n10728), .ZN(n10729) );
  AOI21_X1 U13288 ( .B1(n10730), .B2(n14748), .A(n10729), .ZN(n10731) );
  NAND2_X1 U13289 ( .A1(n10732), .A2(n10731), .ZN(P1_U3257) );
  INV_X1 U13290 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n13478) );
  NAND2_X1 U13291 ( .A1(n7980), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13292 ( .A1(n10733), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U13293 ( .A1(n10734), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n10735) );
  AND3_X1 U13294 ( .A1(n10737), .A2(n10736), .A3(n10735), .ZN(n10738) );
  NAND2_X1 U13295 ( .A1(n10739), .A2(n10738), .ZN(n12039) );
  NAND2_X1 U13296 ( .A1(n12039), .A2(P3_U3897), .ZN(n10740) );
  OAI21_X1 U13297 ( .B1(P3_U3897), .B2(n13478), .A(n10740), .ZN(P3_U3522) );
  NAND2_X1 U13298 ( .A1(n12259), .A2(P3_DATAO_REG_28__SCAN_IN), .ZN(n10741) );
  OAI21_X1 U13299 ( .B1(n12417), .B2(n12259), .A(n10741), .ZN(P3_U3519) );
  INV_X1 U13300 ( .A(n10742), .ZN(n10743) );
  XNOR2_X1 U13301 ( .A(n10744), .B(n10743), .ZN(n10745) );
  NAND3_X1 U13302 ( .A1(n10747), .A2(n10746), .A3(n10745), .ZN(n10750) );
  MUX2_X1 U13303 ( .A(n10749), .B(P3_REG2_REG_0__SCAN_IN), .S(n15371), .Z(
        n10753) );
  INV_X1 U13304 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10783) );
  OAI22_X1 U13305 ( .A1(n15312), .A2(n10751), .B1(n15316), .B2(n10783), .ZN(
        n10752) );
  OR2_X1 U13306 ( .A1(n10753), .A2(n10752), .ZN(P3_U3233) );
  OAI22_X1 U13307 ( .A1(n15048), .A2(n10073), .B1(n10754), .B2(n15050), .ZN(
        n10755) );
  AOI21_X1 U13308 ( .B1(n15027), .B2(n10756), .A(n10755), .ZN(n10757) );
  OAI21_X1 U13309 ( .B1(n15023), .B2(n10758), .A(n10757), .ZN(n10759) );
  AOI21_X1 U13310 ( .B1(n15035), .B2(n10760), .A(n10759), .ZN(n10761) );
  OAI21_X1 U13311 ( .B1(n15038), .B2(n10762), .A(n10761), .ZN(P2_U3263) );
  INV_X1 U13312 ( .A(n10763), .ZN(n10765) );
  OAI222_X1 U13313 ( .A1(P3_U3151), .A2(n10817), .B1(n14576), .B2(n10765), 
        .C1(n10764), .C2(n14574), .ZN(P3_U3274) );
  XNOR2_X1 U13314 ( .A(n10766), .B(n10767), .ZN(n10769) );
  AOI21_X1 U13315 ( .B1(n10769), .B2(n15018), .A(n10768), .ZN(n15118) );
  OAI21_X1 U13316 ( .B1(n10772), .B2(n10771), .A(n10770), .ZN(n15120) );
  INV_X1 U13317 ( .A(n15120), .ZN(n15123) );
  AOI21_X1 U13318 ( .B1(n10773), .B2(n15116), .A(n13219), .ZN(n10774) );
  NAND2_X1 U13319 ( .A1(n10774), .A2(n10853), .ZN(n15117) );
  NAND2_X1 U13320 ( .A1(n13242), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10775) );
  OAI21_X1 U13321 ( .B1(n15050), .B2(n10776), .A(n10775), .ZN(n10777) );
  AOI21_X1 U13322 ( .B1(n15116), .B2(n15027), .A(n10777), .ZN(n10778) );
  OAI21_X1 U13323 ( .B1(n15117), .B2(n15023), .A(n10778), .ZN(n10779) );
  AOI21_X1 U13324 ( .B1(n15123), .B2(n15035), .A(n10779), .ZN(n10780) );
  OAI21_X1 U13325 ( .B1(n15038), .B2(n15118), .A(n10780), .ZN(P2_U3257) );
  INV_X1 U13326 ( .A(n10781), .ZN(n10793) );
  NAND3_X1 U13327 ( .A1(n15300), .A2(n12387), .A3(n15176), .ZN(n10792) );
  NAND2_X1 U13328 ( .A1(n12366), .A2(n10782), .ZN(n10786) );
  NOR2_X1 U13329 ( .A1(n10783), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10784) );
  AOI21_X1 U13330 ( .B1(n15293), .B2(P3_ADDR_REG_0__SCAN_IN), .A(n10784), .ZN(
        n10785) );
  OAI211_X1 U13331 ( .C1(n10787), .C2(n12387), .A(n10786), .B(n10785), .ZN(
        n10791) );
  NOR2_X1 U13332 ( .A1(n15176), .A2(n10788), .ZN(n10789) );
  AOI211_X1 U13333 ( .C1(n10793), .C2(n10792), .A(n10791), .B(n10790), .ZN(
        n10794) );
  INV_X1 U13334 ( .A(n10794), .ZN(P3_U3182) );
  OAI21_X1 U13335 ( .B1(n10796), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10795), 
        .ZN(n10799) );
  MUX2_X1 U13336 ( .A(n10797), .B(P2_REG1_REG_13__SCAN_IN), .S(n11153), .Z(
        n10798) );
  NOR2_X1 U13337 ( .A1(n10799), .A2(n10798), .ZN(n11152) );
  AOI211_X1 U13338 ( .C1(n10799), .C2(n10798), .A(n11152), .B(n15001), .ZN(
        n10809) );
  AOI21_X1 U13339 ( .B1(n10545), .B2(n10801), .A(n10800), .ZN(n10804) );
  MUX2_X1 U13340 ( .A(P2_REG2_REG_13__SCAN_IN), .B(n10802), .S(n11153), .Z(
        n10803) );
  NAND2_X1 U13341 ( .A1(n10803), .A2(n10804), .ZN(n11147) );
  OAI211_X1 U13342 ( .C1(n10804), .C2(n10803), .A(n15009), .B(n11147), .ZN(
        n10807) );
  AND2_X1 U13343 ( .A1(P2_U3088), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n10805) );
  AOI21_X1 U13344 ( .B1(n15007), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10805), 
        .ZN(n10806) );
  OAI211_X1 U13345 ( .C1(n15014), .C2(n11148), .A(n10807), .B(n10806), .ZN(
        n10808) );
  OR2_X1 U13346 ( .A1(n10809), .A2(n10808), .ZN(P2_U3227) );
  OAI222_X1 U13347 ( .A1(n13393), .A2(n10812), .B1(n10810), .B2(P2_U3088), 
        .C1(n13489), .C2(n13395), .ZN(P2_U3306) );
  OAI222_X1 U13348 ( .A1(n10813), .A2(P1_U3086), .B1(n14458), .B2(n10812), 
        .C1(n10811), .C2(n14455), .ZN(P1_U3334) );
  INV_X1 U13349 ( .A(n12695), .ZN(n10824) );
  OAI21_X1 U13350 ( .B1(n10817), .B2(n10816), .A(n10815), .ZN(n10818) );
  INV_X1 U13351 ( .A(n12702), .ZN(n12048) );
  NOR3_X1 U13352 ( .A1(n12048), .A2(n12701), .A3(n11036), .ZN(n10822) );
  AOI211_X1 U13353 ( .C1(n10824), .C2(n10823), .A(n10822), .B(n10955), .ZN(
        n10833) );
  INV_X1 U13354 ( .A(n10826), .ZN(n10828) );
  NOR2_X1 U13355 ( .A1(n15340), .A2(n10827), .ZN(n12242) );
  AOI22_X1 U13356 ( .A1(n10825), .A2(n12005), .B1(n11997), .B2(n12696), .ZN(
        n10829) );
  OAI21_X1 U13357 ( .B1(n10830), .B2(n11979), .A(n10829), .ZN(n10831) );
  AOI21_X1 U13358 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(n10961), .A(n10831), .ZN(
        n10832) );
  OAI21_X1 U13359 ( .B1(n10833), .B2(n12014), .A(n10832), .ZN(P3_U3162) );
  XNOR2_X1 U13360 ( .A(n10834), .B(n10836), .ZN(n15140) );
  XNOR2_X1 U13361 ( .A(n10835), .B(n10836), .ZN(n10840) );
  OR2_X1 U13362 ( .A1(n11354), .A2(n12886), .ZN(n10839) );
  OR2_X1 U13363 ( .A1(n10837), .A2(n12884), .ZN(n10838) );
  AND2_X1 U13364 ( .A1(n10839), .A2(n10838), .ZN(n11050) );
  OAI21_X1 U13365 ( .B1(n10840), .B2(n15039), .A(n11050), .ZN(n15134) );
  INV_X1 U13366 ( .A(n15136), .ZN(n11055) );
  AOI211_X1 U13367 ( .C1(n15136), .C2(n10855), .A(n13219), .B(n15022), .ZN(
        n15135) );
  NAND2_X1 U13368 ( .A1(n15135), .A2(n13259), .ZN(n10843) );
  INV_X1 U13369 ( .A(n10841), .ZN(n11052) );
  AOI22_X1 U13370 ( .A1(n13242), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11052), 
        .B2(n13254), .ZN(n10842) );
  OAI211_X1 U13371 ( .C1(n11055), .C2(n13236), .A(n10843), .B(n10842), .ZN(
        n10844) );
  AOI21_X1 U13372 ( .B1(n15134), .B2(n15048), .A(n10844), .ZN(n10845) );
  OAI21_X1 U13373 ( .B1(n15140), .B2(n13246), .A(n10845), .ZN(P2_U3255) );
  XNOR2_X1 U13374 ( .A(n10846), .B(n10851), .ZN(n10849) );
  OR2_X1 U13375 ( .A1(n11329), .A2(n12886), .ZN(n10848) );
  OR2_X1 U13376 ( .A1(n10997), .A2(n12884), .ZN(n10847) );
  AND2_X1 U13377 ( .A1(n10848), .A2(n10847), .ZN(n11002) );
  OAI21_X1 U13378 ( .B1(n10849), .B2(n15039), .A(n11002), .ZN(n15131) );
  INV_X1 U13379 ( .A(n15131), .ZN(n10861) );
  OAI21_X1 U13380 ( .B1(n10852), .B2(n10851), .A(n10850), .ZN(n15129) );
  INV_X1 U13381 ( .A(n15129), .ZN(n15132) );
  NAND2_X1 U13382 ( .A1(n15126), .A2(n10853), .ZN(n10854) );
  NAND3_X1 U13383 ( .A1(n10855), .A2(n15021), .A3(n10854), .ZN(n15128) );
  NAND2_X1 U13384 ( .A1(n13242), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10856) );
  OAI21_X1 U13385 ( .B1(n15050), .B2(n11003), .A(n10856), .ZN(n10857) );
  AOI21_X1 U13386 ( .B1(n15126), .B2(n15027), .A(n10857), .ZN(n10858) );
  OAI21_X1 U13387 ( .B1(n15128), .B2(n15023), .A(n10858), .ZN(n10859) );
  AOI21_X1 U13388 ( .B1(n15132), .B2(n15035), .A(n10859), .ZN(n10860) );
  OAI21_X1 U13389 ( .B1(n15038), .B2(n10861), .A(n10860), .ZN(P2_U3256) );
  NAND2_X1 U13390 ( .A1(n9028), .A2(n10862), .ZN(n10863) );
  NAND2_X1 U13391 ( .A1(n14799), .A2(n14800), .ZN(n10867) );
  NAND2_X1 U13392 ( .A1(n10874), .A2(n9043), .ZN(n10866) );
  XNOR2_X1 U13393 ( .A(n7219), .B(n10882), .ZN(n14877) );
  INV_X1 U13394 ( .A(n14877), .ZN(n10881) );
  INV_X1 U13395 ( .A(n14801), .ZN(n10870) );
  OAI21_X1 U13396 ( .B1(n10873), .B2(n10872), .A(n10892), .ZN(n10875) );
  OAI22_X1 U13397 ( .A1(n10874), .A2(n14288), .B1(n10886), .B2(n14240), .ZN(
        n14732) );
  AOI21_X1 U13398 ( .B1(n10875), .B2(n14766), .A(n14732), .ZN(n14875) );
  MUX2_X1 U13399 ( .A(n14875), .B(n10876), .S(n14833), .Z(n10880) );
  NOR2_X2 U13400 ( .A1(n14811), .A2(n14810), .ZN(n14814) );
  INV_X1 U13401 ( .A(n14721), .ZN(n10883) );
  NAND2_X1 U13402 ( .A1(n14814), .A2(n10883), .ZN(n10941) );
  OAI211_X1 U13403 ( .C1(n14814), .C2(n10883), .A(n10941), .B(n14812), .ZN(
        n14873) );
  INV_X1 U13404 ( .A(n14873), .ZN(n10878) );
  OAI22_X1 U13405 ( .A1(n14808), .A2(n10883), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14775), .ZN(n10877) );
  AOI21_X1 U13406 ( .B1(n14818), .B2(n10878), .A(n10877), .ZN(n10879) );
  OAI211_X1 U13407 ( .C1(n14323), .C2(n10881), .A(n10880), .B(n10879), .ZN(
        P1_U3290) );
  NAND2_X1 U13408 ( .A1(n10882), .A2(n7219), .ZN(n10885) );
  NAND2_X1 U13409 ( .A1(n10890), .A2(n10883), .ZN(n10884) );
  NAND2_X1 U13410 ( .A1(n10885), .A2(n10884), .ZN(n10939) );
  INV_X1 U13411 ( .A(n10948), .ZN(n10938) );
  NAND2_X1 U13412 ( .A1(n10939), .A2(n10938), .ZN(n10888) );
  NAND2_X1 U13413 ( .A1(n10943), .A2(n10886), .ZN(n10887) );
  INV_X1 U13414 ( .A(n10893), .ZN(n10916) );
  OR2_X1 U13415 ( .A1(n10921), .A2(n13918), .ZN(n10889) );
  INV_X1 U13416 ( .A(n10897), .ZN(n10969) );
  XNOR2_X1 U13417 ( .A(n10970), .B(n10969), .ZN(n14900) );
  INV_X1 U13418 ( .A(n14900), .ZN(n10911) );
  NAND2_X1 U13419 ( .A1(n10890), .A2(n14721), .ZN(n10891) );
  NAND2_X1 U13420 ( .A1(n10914), .A2(n10915), .ZN(n10894) );
  INV_X1 U13421 ( .A(n14783), .ZN(n10895) );
  NAND2_X1 U13422 ( .A1(n10898), .A2(n10897), .ZN(n10980) );
  OR2_X1 U13423 ( .A1(n10898), .A2(n10897), .ZN(n10899) );
  NAND2_X1 U13424 ( .A1(n10980), .A2(n10899), .ZN(n10903) );
  NAND2_X1 U13425 ( .A1(n14769), .A2(n13916), .ZN(n10901) );
  NAND2_X1 U13426 ( .A1(n14771), .A2(n13917), .ZN(n10900) );
  NAND2_X1 U13427 ( .A1(n10901), .A2(n10900), .ZN(n10902) );
  AOI21_X1 U13428 ( .B1(n10903), .B2(n14766), .A(n10902), .ZN(n14904) );
  MUX2_X1 U13429 ( .A(n14904), .B(n10904), .S(n14833), .Z(n10910) );
  INV_X1 U13430 ( .A(n10978), .ZN(n14897) );
  OAI21_X1 U13431 ( .B1(n14793), .B2(n14897), .A(n14812), .ZN(n10905) );
  OR2_X1 U13432 ( .A1(n14759), .A2(n10905), .ZN(n14896) );
  INV_X1 U13433 ( .A(n14896), .ZN(n10908) );
  OAI22_X1 U13434 ( .A1(n14808), .A2(n14897), .B1(n14775), .B2(n10906), .ZN(
        n10907) );
  AOI21_X1 U13435 ( .B1(n10908), .B2(n14818), .A(n10907), .ZN(n10909) );
  OAI211_X1 U13436 ( .C1(n14323), .C2(n10911), .A(n10910), .B(n10909), .ZN(
        P1_U3286) );
  XNOR2_X1 U13437 ( .A(n10912), .B(n10916), .ZN(n14889) );
  INV_X1 U13438 ( .A(n14889), .ZN(n10927) );
  NAND3_X1 U13439 ( .A1(n10914), .A2(n10916), .A3(n10915), .ZN(n10917) );
  AOI21_X1 U13440 ( .B1(n10913), .B2(n10917), .A(n14802), .ZN(n10919) );
  NOR2_X1 U13441 ( .A1(n10919), .A2(n10918), .ZN(n14887) );
  MUX2_X1 U13442 ( .A(n10920), .B(n14887), .S(n14774), .Z(n10926) );
  OAI211_X1 U13443 ( .C1(n10940), .C2(n6957), .A(n14812), .B(n14792), .ZN(
        n14885) );
  INV_X1 U13444 ( .A(n14885), .ZN(n10924) );
  OAI22_X1 U13445 ( .A1(n14808), .A2(n6957), .B1(n14775), .B2(n10922), .ZN(
        n10923) );
  AOI21_X1 U13446 ( .B1(n14818), .B2(n10924), .A(n10923), .ZN(n10925) );
  OAI211_X1 U13447 ( .C1(n14323), .C2(n10927), .A(n10926), .B(n10925), .ZN(
        P1_U3288) );
  XOR2_X1 U13448 ( .A(n10928), .B(n10929), .Z(n10936) );
  INV_X1 U13449 ( .A(n14789), .ZN(n10934) );
  NAND2_X1 U13450 ( .A1(n14769), .A2(n14770), .ZN(n10931) );
  NAND2_X1 U13451 ( .A1(n14771), .A2(n13918), .ZN(n10930) );
  NAND2_X1 U13452 ( .A1(n10931), .A2(n10930), .ZN(n14787) );
  AND2_X1 U13453 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n13967) );
  AOI21_X1 U13454 ( .B1(n14733), .B2(n14787), .A(n13967), .ZN(n10933) );
  NAND2_X1 U13455 ( .A1(n13905), .A2(n14788), .ZN(n10932) );
  OAI211_X1 U13456 ( .C1(n14736), .C2(n10934), .A(n10933), .B(n10932), .ZN(
        n10935) );
  AOI21_X1 U13457 ( .B1(n10936), .B2(n14726), .A(n10935), .ZN(n10937) );
  INV_X1 U13458 ( .A(n10937), .ZN(P1_U3239) );
  XNOR2_X1 U13459 ( .A(n10939), .B(n10938), .ZN(n14883) );
  INV_X1 U13460 ( .A(n14883), .ZN(n10952) );
  AOI211_X1 U13461 ( .C1(n10942), .C2(n10941), .A(n14292), .B(n10940), .ZN(
        n14879) );
  NOR2_X1 U13462 ( .A1(n14808), .A2(n10943), .ZN(n10946) );
  OAI22_X1 U13463 ( .A1(n14774), .A2(n10091), .B1(n10944), .B2(n14775), .ZN(
        n10945) );
  AOI211_X1 U13464 ( .C1(n14879), .C2(n14818), .A(n10946), .B(n10945), .ZN(
        n10951) );
  OAI21_X1 U13465 ( .B1(n10948), .B2(n10947), .A(n10914), .ZN(n10949) );
  AND2_X1 U13466 ( .A1(n10949), .A2(n14766), .ZN(n14881) );
  OAI21_X1 U13467 ( .B1(n14881), .B2(n14878), .A(n14774), .ZN(n10950) );
  OAI211_X1 U13468 ( .C1(n10952), .C2(n14323), .A(n10951), .B(n10950), .ZN(
        P1_U3289) );
  INV_X1 U13469 ( .A(n10953), .ZN(n10954) );
  NOR2_X1 U13470 ( .A1(n10955), .A2(n10954), .ZN(n10958) );
  XNOR2_X1 U13471 ( .A(n10956), .B(n11901), .ZN(n11038) );
  XNOR2_X1 U13472 ( .A(n12698), .B(n11038), .ZN(n10957) );
  AOI21_X1 U13473 ( .B1(n10958), .B2(n10957), .A(n11043), .ZN(n10963) );
  NOR2_X1 U13474 ( .A1(n11979), .A2(n15354), .ZN(n10960) );
  OAI22_X1 U13475 ( .A1(n15339), .A2(n12000), .B1(n15341), .B2(n12008), .ZN(
        n10959) );
  AOI211_X1 U13476 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n10961), .A(n10960), .B(
        n10959), .ZN(n10962) );
  OAI21_X1 U13477 ( .B1(n10963), .B2(n12014), .A(n10962), .ZN(P3_U3177) );
  NOR2_X1 U13478 ( .A1(n14574), .A2(SI_22_), .ZN(n10964) );
  AOI21_X1 U13479 ( .B1(n10965), .B2(P3_STATE_REG_SCAN_IN), .A(n10964), .ZN(
        n10966) );
  OAI21_X1 U13480 ( .B1(n10967), .B2(n14576), .A(n10966), .ZN(n10968) );
  INV_X1 U13481 ( .A(n10968), .ZN(P3_U3273) );
  NAND2_X1 U13482 ( .A1(n10970), .A2(n10969), .ZN(n10972) );
  OR2_X1 U13483 ( .A1(n10978), .A2(n14770), .ZN(n10971) );
  NAND2_X1 U13484 ( .A1(n10972), .A2(n10971), .ZN(n14758) );
  NAND2_X1 U13485 ( .A1(n14758), .A2(n14763), .ZN(n10975) );
  OR2_X1 U13486 ( .A1(n11171), .A2(n13916), .ZN(n10974) );
  NAND2_X1 U13487 ( .A1(n10975), .A2(n10974), .ZN(n11015) );
  XNOR2_X1 U13488 ( .A(n10976), .B(n10983), .ZN(n10989) );
  INV_X1 U13489 ( .A(n14770), .ZN(n10977) );
  NAND2_X1 U13490 ( .A1(n10978), .A2(n10977), .ZN(n10979) );
  NAND2_X1 U13491 ( .A1(n10980), .A2(n10979), .ZN(n14764) );
  OR2_X1 U13492 ( .A1(n11171), .A2(n11214), .ZN(n10981) );
  INV_X1 U13493 ( .A(n10982), .ZN(n10984) );
  INV_X1 U13494 ( .A(n10983), .ZN(n11014) );
  OAI21_X1 U13495 ( .B1(n10984), .B2(n10983), .A(n11010), .ZN(n10986) );
  OAI22_X1 U13496 ( .A1(n11214), .A2(n14288), .B1(n11509), .B2(n14240), .ZN(
        n10985) );
  AOI21_X1 U13497 ( .B1(n10986), .B2(n14766), .A(n10985), .ZN(n10987) );
  OAI21_X1 U13498 ( .B1(n10988), .B2(n10989), .A(n10987), .ZN(n14913) );
  INV_X1 U13499 ( .A(n14913), .ZN(n10994) );
  INV_X1 U13500 ( .A(n10989), .ZN(n14915) );
  INV_X1 U13501 ( .A(n11171), .ZN(n14907) );
  INV_X1 U13502 ( .A(n11206), .ZN(n14912) );
  OAI211_X1 U13503 ( .C1(n14761), .C2(n14912), .A(n14812), .B(n11017), .ZN(
        n14911) );
  INV_X1 U13504 ( .A(n14775), .ZN(n14826) );
  AOI22_X1 U13505 ( .A1(n14315), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n11216), 
        .B2(n14826), .ZN(n10991) );
  NAND2_X1 U13506 ( .A1(n11206), .A2(n14309), .ZN(n10990) );
  OAI211_X1 U13507 ( .C1(n14911), .C2(n14308), .A(n10991), .B(n10990), .ZN(
        n10992) );
  AOI21_X1 U13508 ( .B1(n14915), .B2(n14816), .A(n10992), .ZN(n10993) );
  OAI21_X1 U13509 ( .B1(n10994), .B2(n14315), .A(n10993), .ZN(P1_U3284) );
  NAND2_X1 U13510 ( .A1(n12946), .A2(n13219), .ZN(n12927) );
  INV_X1 U13511 ( .A(n10995), .ZN(n10998) );
  OAI33_X1 U13512 ( .A1(n12927), .A2(n10998), .A3(n10997), .B1(n12938), .B2(
        n8337), .B3(n10996), .ZN(n11000) );
  NAND2_X1 U13513 ( .A1(n11000), .A2(n10999), .ZN(n11007) );
  OAI21_X1 U13514 ( .B1(n12937), .B2(n11002), .A(n11001), .ZN(n11005) );
  NOR2_X1 U13515 ( .A1(n12953), .A2(n11003), .ZN(n11004) );
  AOI211_X1 U13516 ( .C1(n15126), .C2(n8784), .A(n11005), .B(n11004), .ZN(
        n11006) );
  OAI211_X1 U13517 ( .C1(n12938), .C2(n11008), .A(n11007), .B(n11006), .ZN(
        P2_U3203) );
  INV_X1 U13518 ( .A(n14768), .ZN(n11183) );
  NAND2_X1 U13519 ( .A1(n11206), .A2(n11183), .ZN(n11009) );
  AOI21_X1 U13520 ( .B1(n11011), .B2(n11163), .A(n14802), .ZN(n11013) );
  INV_X1 U13521 ( .A(n11163), .ZN(n11012) );
  AOI22_X1 U13522 ( .A1(n11013), .A2(n11161), .B1(n14771), .B2(n14768), .ZN(
        n14919) );
  OR2_X1 U13523 ( .A1(n11206), .A2(n14768), .ZN(n11016) );
  XNOR2_X1 U13524 ( .A(n11164), .B(n11163), .ZN(n14923) );
  NAND2_X1 U13525 ( .A1(n11017), .A2(n14917), .ZN(n11018) );
  NAND3_X1 U13526 ( .A1(n11230), .A2(n14812), .A3(n11018), .ZN(n11020) );
  NAND2_X1 U13527 ( .A1(n14769), .A2(n13914), .ZN(n11019) );
  AND2_X1 U13528 ( .A1(n11020), .A2(n11019), .ZN(n14918) );
  AOI22_X1 U13529 ( .A1(n14315), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n11262), 
        .B2(n14826), .ZN(n11022) );
  NAND2_X1 U13530 ( .A1(n14917), .A2(n14309), .ZN(n11021) );
  OAI211_X1 U13531 ( .C1(n14918), .C2(n14308), .A(n11022), .B(n11021), .ZN(
        n11023) );
  AOI21_X1 U13532 ( .B1(n14923), .B2(n14828), .A(n11023), .ZN(n11024) );
  OAI21_X1 U13533 ( .B1(n14919), .B2(n14833), .A(n11024), .ZN(P1_U3283) );
  OAI21_X1 U13534 ( .B1(n11287), .B2(n11026), .A(n11025), .ZN(n11320) );
  XOR2_X1 U13535 ( .A(n11320), .B(n11313), .Z(n11027) );
  NOR2_X1 U13536 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n11027), .ZN(n11322) );
  AOI21_X1 U13537 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n11027), .A(n11322), 
        .ZN(n11035) );
  OAI21_X1 U13538 ( .B1(n11029), .B2(P1_REG1_REG_14__SCAN_IN), .A(n11028), 
        .ZN(n11312) );
  XOR2_X1 U13539 ( .A(n11312), .B(n11313), .Z(n11030) );
  INV_X1 U13540 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14674) );
  NAND2_X1 U13541 ( .A1(n11030), .A2(n14674), .ZN(n11314) );
  OAI21_X1 U13542 ( .B1(n11030), .B2(n14674), .A(n11314), .ZN(n11033) );
  NAND2_X1 U13543 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n13899)
         );
  NAND2_X1 U13544 ( .A1(n13987), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n11031) );
  OAI211_X1 U13545 ( .C1(n13984), .C2(n11313), .A(n13899), .B(n11031), .ZN(
        n11032) );
  AOI21_X1 U13546 ( .B1(n11033), .B2(n14748), .A(n11032), .ZN(n11034) );
  OAI21_X1 U13547 ( .B1(n11035), .B2(n13941), .A(n11034), .ZN(P1_U3258) );
  XNOR2_X1 U13548 ( .A(n11037), .B(n11898), .ZN(n11266) );
  XNOR2_X1 U13549 ( .A(n15339), .B(n11266), .ZN(n11041) );
  INV_X1 U13550 ( .A(n11038), .ZN(n11039) );
  NOR2_X1 U13551 ( .A1(n10825), .A2(n11039), .ZN(n11042) );
  OAI21_X1 U13552 ( .B1(n11043), .B2(n11042), .A(n11041), .ZN(n11044) );
  NAND3_X1 U13553 ( .A1(n11269), .A2(n11971), .A3(n11044), .ZN(n11047) );
  NOR2_X1 U13554 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15332), .ZN(n15170) );
  OAI22_X1 U13555 ( .A1(n11979), .A2(n15331), .B1(n11242), .B2(n12000), .ZN(
        n11045) );
  AOI211_X1 U13556 ( .C1(n11997), .C2(n10825), .A(n15170), .B(n11045), .ZN(
        n11046) );
  OAI211_X1 U13557 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n11985), .A(n11047), .B(
        n11046), .ZN(P3_U3158) );
  OAI211_X1 U13558 ( .C1(n11049), .C2(n6680), .A(n11048), .B(n12946), .ZN(
        n11054) );
  OAI22_X1 U13559 ( .A1(n12937), .A2(n11050), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14984), .ZN(n11051) );
  AOI21_X1 U13560 ( .B1(n11052), .B2(n12935), .A(n11051), .ZN(n11053) );
  OAI211_X1 U13561 ( .C1(n11055), .C2(n12926), .A(n11054), .B(n11053), .ZN(
        P2_U3189) );
  OAI222_X1 U13562 ( .A1(n13393), .A2(n11058), .B1(n11057), .B2(P2_U3088), 
        .C1(n11056), .C2(n13395), .ZN(P2_U3305) );
  NAND2_X1 U13563 ( .A1(n11059), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n11060) );
  INV_X1 U13564 ( .A(n15180), .ZN(n11123) );
  NAND2_X1 U13565 ( .A1(n11062), .A2(n11123), .ZN(n11063) );
  INV_X1 U13566 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11065) );
  AOI22_X1 U13567 ( .A1(n11125), .A2(P3_REG2_REG_4__SCAN_IN), .B1(n11065), 
        .B2(n15195), .ZN(n15188) );
  NOR2_X1 U13568 ( .A1(n11127), .A2(n11066), .ZN(n11067) );
  INV_X1 U13569 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15207) );
  AOI22_X1 U13570 ( .A1(n11129), .A2(P3_REG2_REG_6__SCAN_IN), .B1(n11093), 
        .B2(n15231), .ZN(n15224) );
  NOR2_X1 U13571 ( .A1(n15225), .A2(n15224), .ZN(n15223) );
  INV_X1 U13572 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11425) );
  MUX2_X1 U13573 ( .A(n11425), .B(P3_REG2_REG_8__SCAN_IN), .S(n15268), .Z(
        n15261) );
  NAND2_X1 U13574 ( .A1(n15268), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U13575 ( .A1(n15259), .A2(n11070), .ZN(n11072) );
  INV_X1 U13576 ( .A(n11071), .ZN(n11073) );
  INV_X1 U13577 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n15280) );
  OAI21_X1 U13578 ( .B1(n11072), .B2(n15289), .A(n11071), .ZN(n15279) );
  NAND2_X1 U13579 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n11443), .ZN(n11074) );
  OAI21_X1 U13580 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n11443), .A(n11074), 
        .ZN(n11075) );
  AOI21_X1 U13581 ( .B1(n11076), .B2(n11075), .A(n6673), .ZN(n11146) );
  INV_X1 U13582 ( .A(n11077), .ZN(n15174) );
  INV_X1 U13583 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n11078) );
  MUX2_X1 U13584 ( .A(n11079), .B(n11078), .S(n12774), .Z(n11080) );
  NAND2_X1 U13585 ( .A1(n11080), .A2(n15180), .ZN(n15191) );
  INV_X1 U13586 ( .A(n11080), .ZN(n11081) );
  NAND2_X1 U13587 ( .A1(n11081), .A2(n11123), .ZN(n11082) );
  AND2_X1 U13588 ( .A1(n15191), .A2(n11082), .ZN(n15173) );
  INV_X1 U13589 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n11083) );
  MUX2_X1 U13590 ( .A(n11065), .B(n11083), .S(n12774), .Z(n11084) );
  NAND2_X1 U13591 ( .A1(n11084), .A2(n11125), .ZN(n11087) );
  INV_X1 U13592 ( .A(n11084), .ZN(n11085) );
  NAND2_X1 U13593 ( .A1(n11085), .A2(n15195), .ZN(n11086) );
  NAND2_X1 U13594 ( .A1(n11087), .A2(n11086), .ZN(n15190) );
  INV_X1 U13595 ( .A(n11087), .ZN(n15209) );
  INV_X1 U13596 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n11088) );
  MUX2_X1 U13597 ( .A(n15207), .B(n11088), .S(n12774), .Z(n11089) );
  NAND2_X1 U13598 ( .A1(n11089), .A2(n11127), .ZN(n15227) );
  INV_X1 U13599 ( .A(n11089), .ZN(n11090) );
  NAND2_X1 U13600 ( .A1(n11090), .A2(n15214), .ZN(n11091) );
  AND2_X1 U13601 ( .A1(n15227), .A2(n11091), .ZN(n15208) );
  INV_X1 U13602 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n11092) );
  MUX2_X1 U13603 ( .A(n11093), .B(n11092), .S(n12774), .Z(n11094) );
  NAND2_X1 U13604 ( .A1(n11094), .A2(n11129), .ZN(n11097) );
  INV_X1 U13605 ( .A(n11094), .ZN(n11095) );
  NAND2_X1 U13606 ( .A1(n11095), .A2(n15231), .ZN(n11096) );
  NAND2_X1 U13607 ( .A1(n11097), .A2(n11096), .ZN(n15226) );
  INV_X1 U13608 ( .A(n11097), .ZN(n15244) );
  INV_X1 U13609 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n11098) );
  MUX2_X1 U13610 ( .A(n11099), .B(n11098), .S(n12774), .Z(n11100) );
  NAND2_X1 U13611 ( .A1(n11100), .A2(n11131), .ZN(n15264) );
  INV_X1 U13612 ( .A(n11100), .ZN(n11101) );
  NAND2_X1 U13613 ( .A1(n11101), .A2(n15249), .ZN(n11102) );
  AND2_X1 U13614 ( .A1(n15264), .A2(n11102), .ZN(n15243) );
  INV_X1 U13615 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11133) );
  MUX2_X1 U13616 ( .A(n11425), .B(n11133), .S(n12774), .Z(n11103) );
  INV_X1 U13617 ( .A(n15268), .ZN(n11134) );
  NAND2_X1 U13618 ( .A1(n11103), .A2(n11134), .ZN(n11106) );
  INV_X1 U13619 ( .A(n11103), .ZN(n11104) );
  NAND2_X1 U13620 ( .A1(n11104), .A2(n15268), .ZN(n11105) );
  NAND2_X1 U13621 ( .A1(n11106), .A2(n11105), .ZN(n15263) );
  INV_X1 U13622 ( .A(n11106), .ZN(n15283) );
  INV_X1 U13623 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n11107) );
  MUX2_X1 U13624 ( .A(n15280), .B(n11107), .S(n12774), .Z(n11108) );
  NAND2_X1 U13625 ( .A1(n11108), .A2(n11135), .ZN(n11115) );
  INV_X1 U13626 ( .A(n11108), .ZN(n11109) );
  NAND2_X1 U13627 ( .A1(n11109), .A2(n15289), .ZN(n11110) );
  AND2_X1 U13628 ( .A1(n11115), .A2(n11110), .ZN(n15282) );
  MUX2_X1 U13629 ( .A(n15311), .B(n15422), .S(n12774), .Z(n11111) );
  NAND2_X1 U13630 ( .A1(n11111), .A2(n11117), .ZN(n11433) );
  INV_X1 U13631 ( .A(n11111), .ZN(n11112) );
  NAND2_X1 U13632 ( .A1(n11112), .A2(n11443), .ZN(n11113) );
  NAND2_X1 U13633 ( .A1(n11433), .A2(n11113), .ZN(n11114) );
  AND3_X1 U13634 ( .A1(n15281), .A2(n11115), .A3(n11114), .ZN(n11116) );
  OAI21_X1 U13635 ( .B1(n11435), .B2(n11116), .A(n15285), .ZN(n11145) );
  INV_X1 U13636 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n15422) );
  AOI22_X1 U13637 ( .A1(n11117), .A2(n15422), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n11443), .ZN(n11139) );
  AOI22_X1 U13638 ( .A1(n11129), .A2(n11092), .B1(P3_REG1_REG_6__SCAN_IN), 
        .B2(n15231), .ZN(n15235) );
  AOI22_X1 U13639 ( .A1(n11125), .A2(n11083), .B1(P3_REG1_REG_4__SCAN_IN), 
        .B2(n15195), .ZN(n15199) );
  INV_X1 U13640 ( .A(n11118), .ZN(n11121) );
  OAI22_X1 U13641 ( .A1(n11121), .A2(n11120), .B1(n6552), .B2(n15413), .ZN(
        n11122) );
  XNOR2_X1 U13642 ( .A(n11122), .B(n15180), .ZN(n15182) );
  AOI22_X1 U13643 ( .A1(n15182), .A2(P3_REG1_REG_3__SCAN_IN), .B1(n11123), 
        .B2(n11122), .ZN(n11124) );
  NAND2_X1 U13644 ( .A1(n15214), .A2(n11126), .ZN(n11128) );
  NAND2_X1 U13645 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n15218), .ZN(n15217) );
  NAND2_X1 U13646 ( .A1(n15249), .A2(n11130), .ZN(n11132) );
  NAND2_X1 U13647 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n15253), .ZN(n15252) );
  NAND2_X1 U13648 ( .A1(n11132), .A2(n15252), .ZN(n15273) );
  MUX2_X1 U13649 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n11133), .S(n15268), .Z(
        n15272) );
  NAND2_X1 U13650 ( .A1(n15273), .A2(n15272), .ZN(n15271) );
  NAND2_X1 U13651 ( .A1(n11136), .A2(n15289), .ZN(n11137) );
  NAND2_X1 U13652 ( .A1(n11139), .A2(n11138), .ZN(n11444) );
  OAI21_X1 U13653 ( .B1(n11139), .B2(n11138), .A(n11444), .ZN(n11143) );
  INV_X1 U13654 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n11140) );
  NOR2_X1 U13655 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11140), .ZN(n11640) );
  AOI21_X1 U13656 ( .B1(n15293), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11640), 
        .ZN(n11141) );
  OAI21_X1 U13657 ( .B1(n15290), .B2(n11443), .A(n11141), .ZN(n11142) );
  AOI21_X1 U13658 ( .B1(n11143), .B2(n15296), .A(n11142), .ZN(n11144) );
  OAI211_X1 U13659 ( .C1(n11146), .C2(n15300), .A(n11145), .B(n11144), .ZN(
        P3_U3192) );
  OAI21_X1 U13660 ( .B1(n11148), .B2(n10802), .A(n11147), .ZN(n11643) );
  XNOR2_X1 U13661 ( .A(n11643), .B(n11658), .ZN(n11644) );
  XNOR2_X1 U13662 ( .A(n11644), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n11158) );
  NOR2_X1 U13663 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12801), .ZN(n11149) );
  AOI21_X1 U13664 ( .B1(n15007), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n11149), 
        .ZN(n11150) );
  OAI21_X1 U13665 ( .B1(n11151), .B2(n15014), .A(n11150), .ZN(n11157) );
  XNOR2_X1 U13666 ( .A(n11658), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11154) );
  AOI211_X1 U13667 ( .C1(n11155), .C2(n11154), .A(n11657), .B(n15001), .ZN(
        n11156) );
  AOI211_X1 U13668 ( .C1(n15009), .C2(n11158), .A(n11157), .B(n11156), .ZN(
        n11159) );
  INV_X1 U13669 ( .A(n11159), .ZN(P2_U3228) );
  OR2_X1 U13670 ( .A1(n14917), .A2(n11509), .ZN(n11160) );
  INV_X1 U13671 ( .A(n11223), .ZN(n11219) );
  XNOR2_X1 U13672 ( .A(n11220), .B(n11219), .ZN(n11162) );
  OAI222_X1 U13673 ( .A1(n14240), .A2(n13865), .B1(n11162), .B2(n14802), .C1(
        n14288), .C2(n11509), .ZN(n14690) );
  INV_X1 U13674 ( .A(n14690), .ZN(n11170) );
  XNOR2_X1 U13675 ( .A(n11224), .B(n11223), .ZN(n14692) );
  INV_X1 U13676 ( .A(n11494), .ZN(n14689) );
  XNOR2_X1 U13677 ( .A(n14689), .B(n11230), .ZN(n11165) );
  NAND2_X1 U13678 ( .A1(n11165), .A2(n14812), .ZN(n14688) );
  AOI22_X1 U13679 ( .A1(n14833), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11511), 
        .B2(n14826), .ZN(n11167) );
  NAND2_X1 U13680 ( .A1(n11494), .A2(n14309), .ZN(n11166) );
  OAI211_X1 U13681 ( .C1(n14688), .C2(n14308), .A(n11167), .B(n11166), .ZN(
        n11168) );
  AOI21_X1 U13682 ( .B1(n14692), .B2(n14828), .A(n11168), .ZN(n11169) );
  OAI21_X1 U13683 ( .B1(n11170), .B2(n14833), .A(n11169), .ZN(P1_U3282) );
  AOI22_X1 U13684 ( .A1(n11171), .A2(n9891), .B1(n9892), .B2(n13916), .ZN(
        n11203) );
  AOI22_X1 U13685 ( .A1(n11171), .A2(n13798), .B1(n9891), .B2(n13916), .ZN(
        n11172) );
  XNOR2_X1 U13686 ( .A(n11172), .B(n6549), .ZN(n11204) );
  XOR2_X1 U13687 ( .A(n11203), .B(n11204), .Z(n11180) );
  INV_X1 U13688 ( .A(n11173), .ZN(n11176) );
  INV_X1 U13689 ( .A(n11174), .ZN(n11175) );
  OAI21_X1 U13690 ( .B1(n11180), .B2(n11179), .A(n11210), .ZN(n11181) );
  NAND2_X1 U13691 ( .A1(n11181), .A2(n14726), .ZN(n11187) );
  NOR2_X1 U13692 ( .A1(n14736), .A2(n14776), .ZN(n11185) );
  OAI21_X1 U13693 ( .B1(n14660), .B2(n11183), .A(n11182), .ZN(n11184) );
  AOI211_X1 U13694 ( .C1(n13901), .C2(n14770), .A(n11185), .B(n11184), .ZN(
        n11186) );
  OAI211_X1 U13695 ( .C1(n14907), .C2(n14659), .A(n11187), .B(n11186), .ZN(
        P1_U3221) );
  NAND2_X1 U13696 ( .A1(n11188), .A2(n14587), .ZN(n11189) );
  OAI211_X1 U13697 ( .C1(n11190), .C2(n14574), .A(n11189), .B(n12246), .ZN(
        P3_U3272) );
  XOR2_X1 U13698 ( .A(n11196), .B(n11191), .Z(n13352) );
  INV_X1 U13699 ( .A(n11341), .ZN(n11192) );
  AOI211_X1 U13700 ( .C1(n13348), .C2(n15020), .A(n13219), .B(n11192), .ZN(
        n13347) );
  INV_X1 U13701 ( .A(n13348), .ZN(n11195) );
  INV_X1 U13702 ( .A(n11361), .ZN(n11193) );
  AOI22_X1 U13703 ( .A1(n13242), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n11193), 
        .B2(n13254), .ZN(n11194) );
  OAI21_X1 U13704 ( .B1(n11195), .B2(n13236), .A(n11194), .ZN(n11201) );
  XNOR2_X1 U13705 ( .A(n11197), .B(n11196), .ZN(n11199) );
  OAI22_X1 U13706 ( .A1(n11198), .A2(n12886), .B1(n11354), .B2(n12884), .ZN(
        n11359) );
  AOI21_X1 U13707 ( .B1(n11199), .B2(n15018), .A(n11359), .ZN(n13350) );
  NOR2_X1 U13708 ( .A1(n13350), .A2(n13242), .ZN(n11200) );
  AOI211_X1 U13709 ( .C1(n13347), .C2(n13259), .A(n11201), .B(n11200), .ZN(
        n11202) );
  OAI21_X1 U13710 ( .B1(n13246), .B2(n13352), .A(n11202), .ZN(P2_U3253) );
  NAND2_X1 U13711 ( .A1(n11204), .A2(n11203), .ZN(n11208) );
  AND2_X1 U13712 ( .A1(n11210), .A2(n11208), .ZN(n11212) );
  AND2_X1 U13713 ( .A1(n9892), .A2(n14768), .ZN(n11205) );
  AOI21_X1 U13714 ( .B1(n11206), .B2(n9891), .A(n11205), .ZN(n11252) );
  AOI22_X1 U13715 ( .A1(n11206), .A2(n13798), .B1(n9891), .B2(n14768), .ZN(
        n11207) );
  XNOR2_X1 U13716 ( .A(n11207), .B(n6549), .ZN(n11251) );
  XOR2_X1 U13717 ( .A(n11252), .B(n11251), .Z(n11211) );
  OAI211_X1 U13718 ( .C1(n11212), .C2(n11211), .A(n14726), .B(n11256), .ZN(
        n11218) );
  INV_X1 U13719 ( .A(n13901), .ZN(n14663) );
  AOI22_X1 U13720 ( .A1(n11507), .A2(n13915), .B1(P1_REG3_REG_9__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11213) );
  OAI21_X1 U13721 ( .B1(n11214), .B2(n14663), .A(n11213), .ZN(n11215) );
  AOI21_X1 U13722 ( .B1(n11216), .B2(n13891), .A(n11215), .ZN(n11217) );
  OAI211_X1 U13723 ( .C1(n14912), .C2(n14659), .A(n11218), .B(n11217), .ZN(
        P1_U3231) );
  OR2_X1 U13724 ( .A1(n11494), .A2(n11260), .ZN(n11221) );
  NAND2_X1 U13725 ( .A1(n11222), .A2(n11221), .ZN(n11278) );
  INV_X1 U13726 ( .A(n11291), .ZN(n11277) );
  XNOR2_X1 U13727 ( .A(n11278), .B(n11277), .ZN(n11229) );
  NAND2_X1 U13728 ( .A1(n11224), .A2(n11223), .ZN(n11226) );
  OR2_X1 U13729 ( .A1(n11494), .A2(n13914), .ZN(n11225) );
  NAND2_X1 U13730 ( .A1(n11226), .A2(n11225), .ZN(n11292) );
  XNOR2_X1 U13731 ( .A(n11292), .B(n11291), .ZN(n14601) );
  OAI22_X1 U13732 ( .A1(n11260), .A2(n14288), .B1(n14662), .B2(n14240), .ZN(
        n11227) );
  AOI21_X1 U13733 ( .B1(n14601), .B2(n14899), .A(n11227), .ZN(n11228) );
  OAI21_X1 U13734 ( .B1(n11229), .B2(n14802), .A(n11228), .ZN(n14599) );
  INV_X1 U13735 ( .A(n14599), .ZN(n11237) );
  AND2_X2 U13736 ( .A1(n14598), .A2(n11232), .ZN(n11305) );
  INV_X1 U13737 ( .A(n11305), .ZN(n11231) );
  OAI211_X1 U13738 ( .C1(n14598), .C2(n11232), .A(n11231), .B(n14812), .ZN(
        n14597) );
  AOI22_X1 U13739 ( .A1(n14833), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11613), 
        .B2(n14826), .ZN(n11234) );
  NAND2_X1 U13740 ( .A1(n11605), .A2(n14309), .ZN(n11233) );
  OAI211_X1 U13741 ( .C1(n14597), .C2(n14308), .A(n11234), .B(n11233), .ZN(
        n11235) );
  AOI21_X1 U13742 ( .B1(n14601), .B2(n14816), .A(n11235), .ZN(n11236) );
  OAI21_X1 U13743 ( .B1(n11237), .B2(n14315), .A(n11236), .ZN(P1_U3281) );
  XNOR2_X1 U13744 ( .A(n11238), .B(n11240), .ZN(n11246) );
  INV_X1 U13745 ( .A(n11239), .ZN(n11241) );
  OR2_X1 U13746 ( .A1(n11239), .A2(n12097), .ZN(n11460) );
  OAI21_X1 U13747 ( .B1(n11241), .B2(n11240), .A(n11460), .ZN(n11244) );
  OAI22_X1 U13748 ( .A1(n11242), .A2(n15340), .B1(n11667), .B2(n15338), .ZN(
        n11243) );
  AOI21_X1 U13749 ( .B1(n11244), .B2(n15323), .A(n11243), .ZN(n11245) );
  OAI21_X1 U13750 ( .B1(n15328), .B2(n11246), .A(n11245), .ZN(n15383) );
  INV_X1 U13751 ( .A(n15383), .ZN(n11250) );
  INV_X1 U13752 ( .A(n11246), .ZN(n15385) );
  NAND2_X1 U13753 ( .A1(n12074), .A2(n15356), .ZN(n15357) );
  INV_X1 U13754 ( .A(n15357), .ZN(n15330) );
  NOR2_X1 U13755 ( .A1(n11397), .A2(n15406), .ZN(n15384) );
  AOI22_X1 U13756 ( .A1(n15333), .A2(n15384), .B1(n15365), .B2(n11385), .ZN(
        n11247) );
  OAI21_X1 U13757 ( .B1(n15207), .B2(n15369), .A(n11247), .ZN(n11248) );
  AOI21_X1 U13758 ( .B1(n15385), .B2(n15366), .A(n11248), .ZN(n11249) );
  OAI21_X1 U13759 ( .B1(n11250), .B2(n15371), .A(n11249), .ZN(P3_U3228) );
  INV_X1 U13760 ( .A(n11251), .ZN(n11254) );
  INV_X1 U13761 ( .A(n11252), .ZN(n11253) );
  AND2_X1 U13762 ( .A1(n9892), .A2(n13915), .ZN(n11257) );
  AOI21_X1 U13763 ( .B1(n14917), .B2(n9891), .A(n11257), .ZN(n11497) );
  AOI22_X1 U13764 ( .A1(n14917), .A2(n13798), .B1(n9891), .B2(n13915), .ZN(
        n11258) );
  XNOR2_X1 U13765 ( .A(n11258), .B(n6549), .ZN(n11496) );
  XOR2_X1 U13766 ( .A(n11497), .B(n11496), .Z(n11501) );
  XNOR2_X1 U13767 ( .A(n11502), .B(n11501), .ZN(n11265) );
  NAND2_X1 U13768 ( .A1(n13901), .A2(n14768), .ZN(n11259) );
  NAND2_X1 U13769 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n13982)
         );
  OAI211_X1 U13770 ( .C1(n11260), .C2(n14660), .A(n11259), .B(n13982), .ZN(
        n11261) );
  AOI21_X1 U13771 ( .B1(n11262), .B2(n13891), .A(n11261), .ZN(n11264) );
  NAND2_X1 U13772 ( .A1(n14917), .A2(n13905), .ZN(n11263) );
  OAI211_X1 U13773 ( .C1(n11265), .C2(n13908), .A(n11264), .B(n11263), .ZN(
        P1_U3217) );
  INV_X1 U13774 ( .A(n11412), .ZN(n11276) );
  INV_X1 U13775 ( .A(n11266), .ZN(n11267) );
  NAND2_X1 U13776 ( .A1(n11267), .A2(n12258), .ZN(n11268) );
  XNOR2_X1 U13777 ( .A(n11272), .B(n11901), .ZN(n11270) );
  NOR2_X1 U13778 ( .A1(n15320), .A2(n11270), .ZN(n11387) );
  AOI21_X1 U13779 ( .B1(n15320), .B2(n11270), .A(n11387), .ZN(n11389) );
  NAND2_X1 U13780 ( .A1(n11393), .A2(n11389), .ZN(n11388) );
  OAI21_X1 U13781 ( .B1(n11393), .B2(n11389), .A(n11388), .ZN(n11271) );
  NAND2_X1 U13782 ( .A1(n11271), .A2(n11971), .ZN(n11275) );
  INV_X1 U13783 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n13532) );
  NOR2_X1 U13784 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13532), .ZN(n15197) );
  OAI22_X1 U13785 ( .A1(n11567), .A2(n12000), .B1(n11979), .B2(n11272), .ZN(
        n11273) );
  AOI211_X1 U13786 ( .C1(n11997), .C2(n12258), .A(n15197), .B(n11273), .ZN(
        n11274) );
  OAI211_X1 U13787 ( .C1(n11276), .C2(n11985), .A(n11275), .B(n11274), .ZN(
        P3_U3170) );
  NAND2_X1 U13788 ( .A1(n11278), .A2(n11277), .ZN(n11280) );
  OR2_X1 U13789 ( .A1(n11605), .A2(n13865), .ZN(n11279) );
  NAND2_X1 U13790 ( .A1(n11280), .A2(n11279), .ZN(n11300) );
  INV_X1 U13791 ( .A(n11303), .ZN(n11299) );
  NAND2_X1 U13792 ( .A1(n11300), .A2(n11299), .ZN(n11282) );
  OR2_X1 U13793 ( .A1(n13869), .A2(n14662), .ZN(n11281) );
  NAND2_X1 U13794 ( .A1(n11282), .A2(n11281), .ZN(n11584) );
  INV_X1 U13795 ( .A(n11583), .ZN(n11283) );
  XNOR2_X1 U13796 ( .A(n11584), .B(n11283), .ZN(n11286) );
  NAND2_X1 U13797 ( .A1(n14771), .A2(n13912), .ZN(n11284) );
  OAI21_X1 U13798 ( .B1(n14661), .B2(n14240), .A(n11284), .ZN(n11285) );
  AOI21_X1 U13799 ( .B1(n11286), .B2(n14766), .A(n11285), .ZN(n14682) );
  OAI22_X1 U13800 ( .A1(n14774), .A2(n11287), .B1(n14669), .B2(n14775), .ZN(
        n11290) );
  INV_X1 U13801 ( .A(n13869), .ZN(n14684) );
  NAND2_X1 U13802 ( .A1(n14684), .A2(n11305), .ZN(n11304) );
  AOI21_X1 U13803 ( .B1(n14658), .B2(n11304), .A(n14292), .ZN(n11288) );
  NAND2_X1 U13804 ( .A1(n11288), .A2(n11592), .ZN(n14677) );
  NOR2_X1 U13805 ( .A1(n14677), .A2(n14308), .ZN(n11289) );
  AOI211_X1 U13806 ( .C1(n14309), .C2(n14658), .A(n11290), .B(n11289), .ZN(
        n11298) );
  NAND2_X1 U13807 ( .A1(n11292), .A2(n11291), .ZN(n11294) );
  OR2_X1 U13808 ( .A1(n11605), .A2(n13913), .ZN(n11293) );
  NAND2_X1 U13809 ( .A1(n11294), .A2(n11293), .ZN(n11302) );
  OR2_X1 U13810 ( .A1(n13869), .A2(n13912), .ZN(n11295) );
  NAND2_X1 U13811 ( .A1(n11296), .A2(n11583), .ZN(n14675) );
  NAND3_X1 U13812 ( .A1(n14676), .A2(n14675), .A3(n14828), .ZN(n11297) );
  OAI211_X1 U13813 ( .C1(n14682), .C2(n14315), .A(n11298), .B(n11297), .ZN(
        P1_U3279) );
  XNOR2_X1 U13814 ( .A(n11300), .B(n11299), .ZN(n11301) );
  OAI222_X1 U13815 ( .A1(n14240), .A2(n13864), .B1(n11301), .B2(n14802), .C1(
        n14288), .C2(n13865), .ZN(n14685) );
  INV_X1 U13816 ( .A(n14685), .ZN(n11310) );
  XNOR2_X1 U13817 ( .A(n11302), .B(n11303), .ZN(n14687) );
  OAI211_X1 U13818 ( .C1(n14684), .C2(n11305), .A(n14812), .B(n11304), .ZN(
        n14683) );
  AOI22_X1 U13819 ( .A1(n14833), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n13868), 
        .B2(n14826), .ZN(n11307) );
  NAND2_X1 U13820 ( .A1(n13869), .A2(n14309), .ZN(n11306) );
  OAI211_X1 U13821 ( .C1(n14683), .C2(n14308), .A(n11307), .B(n11306), .ZN(
        n11308) );
  AOI21_X1 U13822 ( .B1(n14687), .B2(n14828), .A(n11308), .ZN(n11309) );
  OAI21_X1 U13823 ( .B1(n11310), .B2(n14833), .A(n11309), .ZN(P1_U3280) );
  INV_X1 U13824 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11311) );
  NAND2_X1 U13825 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13831)
         );
  OAI21_X1 U13826 ( .B1(n14756), .B2(n11311), .A(n13831), .ZN(n11319) );
  NAND2_X1 U13827 ( .A1(n11313), .A2(n11312), .ZN(n11315) );
  NAND2_X1 U13828 ( .A1(n11315), .A2(n11314), .ZN(n11317) );
  XNOR2_X1 U13829 ( .A(n14003), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11316) );
  NOR2_X1 U13830 ( .A1(n11316), .A2(n11317), .ZN(n13996) );
  AOI211_X1 U13831 ( .C1(n11317), .C2(n11316), .A(n13996), .B(n14036), .ZN(
        n11318) );
  AOI211_X1 U13832 ( .C1(n14750), .C2(n14003), .A(n11319), .B(n11318), .ZN(
        n11328) );
  NOR2_X1 U13833 ( .A1(n11321), .A2(n11320), .ZN(n11323) );
  NOR2_X1 U13834 ( .A1(n11323), .A2(n11322), .ZN(n11326) );
  MUX2_X1 U13835 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n11324), .S(n14003), .Z(
        n11325) );
  NAND2_X1 U13836 ( .A1(n11325), .A2(n11326), .ZN(n14004) );
  OAI211_X1 U13837 ( .C1(n11326), .C2(n11325), .A(n14752), .B(n14004), .ZN(
        n11327) );
  NAND2_X1 U13838 ( .A1(n11328), .A2(n11327), .ZN(P1_U3259) );
  OAI22_X1 U13839 ( .A1(n11329), .A2(n12884), .B1(n11348), .B2(n12886), .ZN(
        n15017) );
  AOI22_X1 U13840 ( .A1(n12950), .A2(n15017), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11330) );
  OAI21_X1 U13841 ( .B1(n12953), .B2(n15025), .A(n11330), .ZN(n11338) );
  INV_X1 U13842 ( .A(n12927), .ZN(n12945) );
  NAND3_X1 U13843 ( .A1(n11331), .A2(n12945), .A3(n12978), .ZN(n11336) );
  INV_X1 U13844 ( .A(n11048), .ZN(n11333) );
  OAI21_X1 U13845 ( .B1(n11333), .B2(n11332), .A(n12946), .ZN(n11335) );
  INV_X1 U13846 ( .A(n11334), .ZN(n11357) );
  AOI21_X1 U13847 ( .B1(n11336), .B2(n11335), .A(n11357), .ZN(n11337) );
  AOI211_X1 U13848 ( .C1(n15028), .C2(n8784), .A(n11338), .B(n11337), .ZN(
        n11339) );
  INV_X1 U13849 ( .A(n11339), .ZN(P2_U3208) );
  XOR2_X1 U13850 ( .A(n11340), .B(n11346), .Z(n14654) );
  AOI21_X1 U13851 ( .B1(n14650), .B2(n11341), .A(n13219), .ZN(n11342) );
  NAND2_X1 U13852 ( .A1(n11342), .A2(n11369), .ZN(n14651) );
  NAND2_X1 U13853 ( .A1(n13242), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11343) );
  OAI21_X1 U13854 ( .B1(n15050), .B2(n12905), .A(n11343), .ZN(n11344) );
  AOI21_X1 U13855 ( .B1(n14650), .B2(n15027), .A(n11344), .ZN(n11345) );
  OAI21_X1 U13856 ( .B1(n14651), .B2(n15023), .A(n11345), .ZN(n11352) );
  XNOR2_X1 U13857 ( .A(n11347), .B(n11346), .ZN(n11350) );
  OAI22_X1 U13858 ( .A1(n11349), .A2(n12886), .B1(n11348), .B2(n12884), .ZN(
        n12903) );
  AOI21_X1 U13859 ( .B1(n11350), .B2(n15018), .A(n12903), .ZN(n14652) );
  NOR2_X1 U13860 ( .A1(n14652), .A2(n15038), .ZN(n11351) );
  AOI211_X1 U13861 ( .C1(n14654), .C2(n15035), .A(n11352), .B(n11351), .ZN(
        n11353) );
  INV_X1 U13862 ( .A(n11353), .ZN(P2_U3252) );
  NOR3_X1 U13863 ( .A1(n11355), .A2(n11354), .A3(n12927), .ZN(n11356) );
  AOI21_X1 U13864 ( .B1(n11357), .B2(n12946), .A(n11356), .ZN(n11367) );
  AOI21_X1 U13865 ( .B1(n12950), .B2(n11359), .A(n11358), .ZN(n11360) );
  OAI21_X1 U13866 ( .B1(n12953), .B2(n11361), .A(n11360), .ZN(n11364) );
  NOR2_X1 U13867 ( .A1(n11362), .A2(n12938), .ZN(n11363) );
  AOI211_X1 U13868 ( .C1(n13348), .C2(n8784), .A(n11364), .B(n11363), .ZN(
        n11365) );
  OAI21_X1 U13869 ( .B1(n11367), .B2(n11366), .A(n11365), .ZN(P2_U3196) );
  XOR2_X1 U13870 ( .A(n11368), .B(n11374), .Z(n13346) );
  AOI211_X1 U13871 ( .C1(n13344), .C2(n11369), .A(n13219), .B(n6548), .ZN(
        n13343) );
  NOR2_X1 U13872 ( .A1(n7207), .A2(n13236), .ZN(n11372) );
  INV_X1 U13873 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11370) );
  OAI22_X1 U13874 ( .A1(n15048), .A2(n11370), .B1(n12800), .B2(n15050), .ZN(
        n11371) );
  AOI211_X1 U13875 ( .C1(n13343), .C2(n13259), .A(n11372), .B(n11371), .ZN(
        n11377) );
  XOR2_X1 U13876 ( .A(n11373), .B(n11374), .Z(n11375) );
  AOI22_X1 U13877 ( .A1(n12973), .A2(n12933), .B1(n12932), .B2(n12975), .ZN(
        n12802) );
  OAI21_X1 U13878 ( .B1(n11375), .B2(n15039), .A(n12802), .ZN(n13342) );
  NAND2_X1 U13879 ( .A1(n13342), .A2(n15048), .ZN(n11376) );
  OAI211_X1 U13880 ( .C1(n13346), .C2(n13246), .A(n11377), .B(n11376), .ZN(
        P2_U3251) );
  INV_X1 U13881 ( .A(n11378), .ZN(n11384) );
  AOI21_X1 U13882 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n14444), .A(n11379), 
        .ZN(n11380) );
  OAI21_X1 U13883 ( .B1(n11384), .B2(n14458), .A(n11380), .ZN(P1_U3332) );
  AOI21_X1 U13884 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n11382), .A(n11381), 
        .ZN(n11383) );
  OAI21_X1 U13885 ( .B1(n11384), .B2(n13393), .A(n11383), .ZN(P2_U3304) );
  INV_X1 U13886 ( .A(n11385), .ZN(n11401) );
  XNOR2_X1 U13887 ( .A(n11386), .B(n11901), .ZN(n11566) );
  XNOR2_X1 U13888 ( .A(n11566), .B(n12257), .ZN(n11395) );
  INV_X1 U13889 ( .A(n11387), .ZN(n11390) );
  NAND2_X1 U13890 ( .A1(n11388), .A2(n11390), .ZN(n11394) );
  AND2_X1 U13891 ( .A1(n11389), .A2(n11395), .ZN(n11392) );
  INV_X1 U13892 ( .A(n11395), .ZN(n11391) );
  OAI21_X1 U13893 ( .B1(n11395), .B2(n11394), .A(n6656), .ZN(n11396) );
  NAND2_X1 U13894 ( .A1(n11396), .A2(n11971), .ZN(n11400) );
  AND2_X1 U13895 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n15216) );
  OAI22_X1 U13896 ( .A1(n11979), .A2(n11397), .B1(n11667), .B2(n12000), .ZN(
        n11398) );
  AOI211_X1 U13897 ( .C1(n11997), .C2(n15320), .A(n15216), .B(n11398), .ZN(
        n11399) );
  OAI211_X1 U13898 ( .C1(n11401), .C2(n11985), .A(n11400), .B(n11399), .ZN(
        P3_U3167) );
  OAI21_X1 U13899 ( .B1(n11403), .B2(n12092), .A(n11402), .ZN(n15382) );
  INV_X1 U13900 ( .A(n15382), .ZN(n11415) );
  INV_X1 U13901 ( .A(n15366), .ZN(n11557) );
  OAI22_X1 U13902 ( .A1(n11567), .A2(n15338), .B1(n15339), .B2(n15340), .ZN(
        n11410) );
  INV_X1 U13903 ( .A(n11404), .ZN(n15325) );
  OR2_X1 U13904 ( .A1(n11404), .A2(n7919), .ZN(n15322) );
  NAND2_X1 U13905 ( .A1(n15322), .A2(n11405), .ZN(n11407) );
  XNOR2_X1 U13906 ( .A(n11407), .B(n11406), .ZN(n11408) );
  NOR2_X1 U13907 ( .A1(n11408), .A2(n15347), .ZN(n11409) );
  AOI211_X1 U13908 ( .C1(n15352), .C2(n15382), .A(n11410), .B(n11409), .ZN(
        n15379) );
  MUX2_X1 U13909 ( .A(n11065), .B(n15379), .S(n15369), .Z(n11414) );
  AND2_X1 U13910 ( .A1(n11411), .A2(n14625), .ZN(n15381) );
  AOI22_X1 U13911 ( .A1(n15333), .A2(n15381), .B1(n15365), .B2(n11412), .ZN(
        n11413) );
  OAI211_X1 U13912 ( .C1(n11415), .C2(n11557), .A(n11414), .B(n11413), .ZN(
        P3_U3229) );
  OR2_X1 U13913 ( .A1(n11416), .A2(n12113), .ZN(n11417) );
  NAND2_X1 U13914 ( .A1(n11418), .A2(n11417), .ZN(n15395) );
  XNOR2_X1 U13915 ( .A(n11419), .B(n12113), .ZN(n11420) );
  NAND2_X1 U13916 ( .A1(n11420), .A2(n15323), .ZN(n11422) );
  AOI22_X1 U13917 ( .A1(n12255), .A2(n15321), .B1(n15319), .B2(n15303), .ZN(
        n11421) );
  NAND2_X1 U13918 ( .A1(n11422), .A2(n11421), .ZN(n11423) );
  AOI21_X1 U13919 ( .B1(n15395), .B2(n15352), .A(n11423), .ZN(n15397) );
  AND2_X1 U13920 ( .A1(n11565), .A2(n14625), .ZN(n15394) );
  AOI22_X1 U13921 ( .A1(n15333), .A2(n15394), .B1(n15365), .B2(n11753), .ZN(
        n11424) );
  OAI21_X1 U13922 ( .B1(n11425), .B2(n15369), .A(n11424), .ZN(n11426) );
  AOI21_X1 U13923 ( .B1(n15395), .B2(n15366), .A(n11426), .ZN(n11427) );
  OAI21_X1 U13924 ( .B1(n15397), .B2(n15371), .A(n11427), .ZN(P3_U3225) );
  NOR2_X1 U13925 ( .A1(n11447), .A2(n11429), .ZN(n11430) );
  INV_X1 U13926 ( .A(n14580), .ZN(n11698) );
  AOI22_X1 U13927 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n11698), .B1(n14580), 
        .B2(n11765), .ZN(n11431) );
  AOI21_X1 U13928 ( .B1(n11432), .B2(n11431), .A(n11692), .ZN(n11457) );
  INV_X1 U13929 ( .A(n11433), .ZN(n11434) );
  MUX2_X1 U13930 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12774), .Z(n11436) );
  XNOR2_X1 U13931 ( .A(n11436), .B(n14573), .ZN(n11527) );
  NOR2_X1 U13932 ( .A1(n11528), .A2(n11527), .ZN(n11526) );
  MUX2_X1 U13933 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12774), .Z(n11697) );
  XNOR2_X1 U13934 ( .A(n11697), .B(n14580), .ZN(n11440) );
  INV_X1 U13935 ( .A(n11440), .ZN(n11438) );
  NOR2_X1 U13936 ( .A1(n11436), .A2(n14573), .ZN(n11441) );
  OAI21_X1 U13937 ( .B1(n11526), .B2(n11441), .A(n11440), .ZN(n11442) );
  NAND3_X1 U13938 ( .A1(n11701), .A2(n15285), .A3(n11442), .ZN(n11456) );
  INV_X1 U13939 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14636) );
  AOI22_X1 U13940 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n14580), .B1(n11698), 
        .B2(n14636), .ZN(n11450) );
  NAND2_X1 U13941 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n11443), .ZN(n11445) );
  NAND2_X1 U13942 ( .A1(n11445), .A2(n11444), .ZN(n11446) );
  NAND2_X1 U13943 ( .A1(n14573), .A2(n11446), .ZN(n11448) );
  XNOR2_X1 U13944 ( .A(n11447), .B(n11446), .ZN(n11524) );
  NAND2_X1 U13945 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n11524), .ZN(n11523) );
  OAI21_X1 U13946 ( .B1(n11450), .B2(n11449), .A(n11694), .ZN(n11454) );
  INV_X1 U13947 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11451) );
  NOR2_X1 U13948 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11451), .ZN(n11789) );
  AOI21_X1 U13949 ( .B1(n15293), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n11789), 
        .ZN(n11452) );
  OAI21_X1 U13950 ( .B1(n15290), .B2(n14580), .A(n11452), .ZN(n11453) );
  AOI21_X1 U13951 ( .B1(n11454), .B2(n15296), .A(n11453), .ZN(n11455) );
  OAI211_X1 U13952 ( .C1(n11457), .C2(n15300), .A(n11456), .B(n11455), .ZN(
        P3_U3194) );
  INV_X1 U13953 ( .A(n11458), .ZN(n11459) );
  NAND2_X1 U13954 ( .A1(n11460), .A2(n11459), .ZN(n11548) );
  NOR2_X1 U13955 ( .A1(n11548), .A2(n12044), .ZN(n11551) );
  NOR2_X1 U13956 ( .A1(n11551), .A2(n11461), .ZN(n11462) );
  XNOR2_X1 U13957 ( .A(n11462), .B(n12108), .ZN(n11466) );
  XNOR2_X1 U13958 ( .A(n11463), .B(n12108), .ZN(n15393) );
  OAI22_X1 U13959 ( .A1(n11671), .A2(n15338), .B1(n11667), .B2(n15340), .ZN(
        n11464) );
  AOI21_X1 U13960 ( .B1(n15393), .B2(n15352), .A(n11464), .ZN(n11465) );
  OAI21_X1 U13961 ( .B1(n11466), .B2(n15347), .A(n11465), .ZN(n15391) );
  INV_X1 U13962 ( .A(n15391), .ZN(n11470) );
  NOR2_X1 U13963 ( .A1(n11670), .A2(n15406), .ZN(n15392) );
  AOI22_X1 U13964 ( .A1(n15333), .A2(n15392), .B1(n15365), .B2(n11673), .ZN(
        n11467) );
  OAI21_X1 U13965 ( .B1(n11099), .B2(n15369), .A(n11467), .ZN(n11468) );
  AOI21_X1 U13966 ( .B1(n15393), .B2(n15366), .A(n11468), .ZN(n11469) );
  OAI21_X1 U13967 ( .B1(n11470), .B2(n15371), .A(n11469), .ZN(P3_U3226) );
  XNOR2_X1 U13968 ( .A(n11471), .B(n11475), .ZN(n11474) );
  NAND2_X1 U13969 ( .A1(n12972), .A2(n12933), .ZN(n11473) );
  NAND2_X1 U13970 ( .A1(n12932), .A2(n12974), .ZN(n11472) );
  NAND2_X1 U13971 ( .A1(n11473), .A2(n11472), .ZN(n12949) );
  AOI21_X1 U13972 ( .B1(n11474), .B2(n15018), .A(n12949), .ZN(n11515) );
  XNOR2_X1 U13973 ( .A(n11476), .B(n11475), .ZN(n11517) );
  AOI21_X1 U13974 ( .B1(n12955), .B2(n11477), .A(n13219), .ZN(n11478) );
  NAND2_X1 U13975 ( .A1(n11478), .A2(n11540), .ZN(n11514) );
  NAND2_X1 U13976 ( .A1(n13242), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n11479) );
  OAI21_X1 U13977 ( .B1(n15050), .B2(n12952), .A(n11479), .ZN(n11480) );
  AOI21_X1 U13978 ( .B1(n12955), .B2(n15027), .A(n11480), .ZN(n11481) );
  OAI21_X1 U13979 ( .B1(n11514), .B2(n15023), .A(n11481), .ZN(n11482) );
  AOI21_X1 U13980 ( .B1(n11517), .B2(n15035), .A(n11482), .ZN(n11483) );
  OAI21_X1 U13981 ( .B1(n15038), .B2(n11515), .A(n11483), .ZN(P2_U3250) );
  XNOR2_X1 U13982 ( .A(n11484), .B(n12118), .ZN(n15401) );
  NAND2_X1 U13983 ( .A1(n11485), .A2(n12118), .ZN(n11486) );
  NAND3_X1 U13984 ( .A1(n11487), .A2(n15323), .A3(n11486), .ZN(n11489) );
  AOI22_X1 U13985 ( .A1(n12253), .A2(n15319), .B1(n15321), .B2(n12254), .ZN(
        n11488) );
  NAND2_X1 U13986 ( .A1(n11489), .A2(n11488), .ZN(n11490) );
  AOI21_X1 U13987 ( .B1(n15401), .B2(n15352), .A(n11490), .ZN(n15403) );
  AND2_X1 U13988 ( .A1(n12120), .A2(n14625), .ZN(n15399) );
  AOI22_X1 U13989 ( .A1(n15333), .A2(n15399), .B1(n15365), .B2(n11563), .ZN(
        n11491) );
  OAI21_X1 U13990 ( .B1(n15280), .B2(n15369), .A(n11491), .ZN(n11492) );
  AOI21_X1 U13991 ( .B1(n15401), .B2(n15366), .A(n11492), .ZN(n11493) );
  OAI21_X1 U13992 ( .B1(n15403), .B2(n15371), .A(n11493), .ZN(P3_U3224) );
  AOI22_X1 U13993 ( .A1(n11494), .A2(n9891), .B1(n9892), .B2(n13914), .ZN(
        n11599) );
  AOI22_X1 U13994 ( .A1(n11494), .A2(n13798), .B1(n9891), .B2(n13914), .ZN(
        n11495) );
  XNOR2_X1 U13995 ( .A(n11495), .B(n6549), .ZN(n11600) );
  XOR2_X1 U13996 ( .A(n11599), .B(n11600), .Z(n11504) );
  INV_X1 U13997 ( .A(n11496), .ZN(n11499) );
  INV_X1 U13998 ( .A(n11497), .ZN(n11498) );
  NAND2_X1 U13999 ( .A1(n11503), .A2(n11504), .ZN(n11608) );
  OAI21_X1 U14000 ( .B1(n11504), .B2(n11503), .A(n11608), .ZN(n11505) );
  NAND2_X1 U14001 ( .A1(n11505), .A2(n14726), .ZN(n11513) );
  AOI21_X1 U14002 ( .B1(n11507), .B2(n13913), .A(n11506), .ZN(n11508) );
  OAI21_X1 U14003 ( .B1(n11509), .B2(n14663), .A(n11508), .ZN(n11510) );
  AOI21_X1 U14004 ( .B1(n11511), .B2(n13891), .A(n11510), .ZN(n11512) );
  OAI211_X1 U14005 ( .C1(n14689), .C2(n14659), .A(n11513), .B(n11512), .ZN(
        P1_U3236) );
  OAI211_X1 U14006 ( .C1(n7206), .C2(n15146), .A(n11515), .B(n11514), .ZN(
        n11516) );
  AOI21_X1 U14007 ( .B1(n11517), .B2(n15151), .A(n11516), .ZN(n11520) );
  NAND2_X1 U14008 ( .A1(n15153), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11518) );
  OAI21_X1 U14009 ( .B1(n11520), .B2(n15153), .A(n11518), .ZN(P2_U3475) );
  NAND2_X1 U14010 ( .A1(n15164), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11519) );
  OAI21_X1 U14011 ( .B1(n11520), .B2(n15164), .A(n11519), .ZN(P2_U3514) );
  AOI21_X1 U14012 ( .B1(n7671), .B2(n11522), .A(n11521), .ZN(n11534) );
  OAI21_X1 U14013 ( .B1(P3_REG1_REG_11__SCAN_IN), .B2(n11524), .A(n11523), 
        .ZN(n11532) );
  AND2_X1 U14014 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11716) );
  AOI21_X1 U14015 ( .B1(n15293), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n11716), 
        .ZN(n11525) );
  OAI21_X1 U14016 ( .B1(n15290), .B2(n14573), .A(n11525), .ZN(n11531) );
  AOI21_X1 U14017 ( .B1(n11528), .B2(n11527), .A(n11526), .ZN(n11529) );
  NOR2_X1 U14018 ( .A1(n11529), .A2(n15176), .ZN(n11530) );
  AOI211_X1 U14019 ( .C1(n15296), .C2(n11532), .A(n11531), .B(n11530), .ZN(
        n11533) );
  OAI21_X1 U14020 ( .B1(n11534), .B2(n15300), .A(n11533), .ZN(P3_U3193) );
  XNOR2_X1 U14021 ( .A(n11535), .B(n11536), .ZN(n13341) );
  XNOR2_X1 U14022 ( .A(n11537), .B(n11536), .ZN(n11539) );
  AND2_X1 U14023 ( .A1(n12973), .A2(n12932), .ZN(n11538) );
  AOI21_X1 U14024 ( .B1(n12971), .B2(n12933), .A(n11538), .ZN(n12863) );
  OAI21_X1 U14025 ( .B1(n11539), .B2(n15039), .A(n12863), .ZN(n13337) );
  INV_X1 U14026 ( .A(n13339), .ZN(n11543) );
  AOI211_X1 U14027 ( .C1(n13339), .C2(n11540), .A(n13219), .B(n13229), .ZN(
        n13338) );
  NAND2_X1 U14028 ( .A1(n13338), .A2(n13259), .ZN(n11542) );
  AOI22_X1 U14029 ( .A1(n13242), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n12865), 
        .B2(n13254), .ZN(n11541) );
  OAI211_X1 U14030 ( .C1(n11543), .C2(n13236), .A(n11542), .B(n11541), .ZN(
        n11544) );
  AOI21_X1 U14031 ( .B1(n13337), .B2(n15048), .A(n11544), .ZN(n11545) );
  OAI21_X1 U14032 ( .B1(n13341), .B2(n13246), .A(n11545), .ZN(P2_U3249) );
  XNOR2_X1 U14033 ( .A(n11546), .B(n11547), .ZN(n15387) );
  NAND2_X1 U14034 ( .A1(n11548), .A2(n12044), .ZN(n11549) );
  NAND2_X1 U14035 ( .A1(n11549), .A2(n15323), .ZN(n11550) );
  OR2_X1 U14036 ( .A1(n11551), .A2(n11550), .ZN(n11553) );
  AOI22_X1 U14037 ( .A1(n12255), .A2(n15319), .B1(n15321), .B2(n12257), .ZN(
        n11552) );
  OAI211_X1 U14038 ( .C1(n15328), .C2(n15387), .A(n11553), .B(n11552), .ZN(
        n15388) );
  MUX2_X1 U14039 ( .A(n15388), .B(P3_REG2_REG_6__SCAN_IN), .S(n15371), .Z(
        n11554) );
  INV_X1 U14040 ( .A(n11554), .ZN(n11556) );
  NOR2_X1 U14041 ( .A1(n11687), .A2(n15406), .ZN(n15389) );
  AOI22_X1 U14042 ( .A1(n15333), .A2(n15389), .B1(n15365), .B2(n11681), .ZN(
        n11555) );
  OAI211_X1 U14043 ( .C1(n15387), .C2(n11557), .A(n11556), .B(n11555), .ZN(
        P3_U3227) );
  OAI22_X1 U14044 ( .A1(n11559), .A2(P3_U3151), .B1(n11558), .B2(n14574), .ZN(
        n11560) );
  AOI21_X1 U14045 ( .B1(n11561), .B2(n14587), .A(n11560), .ZN(n11562) );
  INV_X1 U14046 ( .A(n11562), .ZN(P3_U3271) );
  INV_X1 U14047 ( .A(n11563), .ZN(n11582) );
  XNOR2_X1 U14048 ( .A(n12120), .B(n11898), .ZN(n11633) );
  XNOR2_X1 U14049 ( .A(n11633), .B(n15303), .ZN(n11576) );
  XNOR2_X1 U14050 ( .A(n11564), .B(n11901), .ZN(n11669) );
  XNOR2_X1 U14051 ( .A(n11565), .B(n11901), .ZN(n11570) );
  XNOR2_X1 U14052 ( .A(n12254), .B(n11570), .ZN(n11748) );
  NAND2_X1 U14053 ( .A1(n11567), .A2(n11566), .ZN(n11665) );
  XNOR2_X1 U14054 ( .A(n11568), .B(n11901), .ZN(n11666) );
  NAND2_X1 U14055 ( .A1(n11667), .A2(n11666), .ZN(n11569) );
  AND4_X1 U14056 ( .A1(n11744), .A2(n11748), .A3(n11665), .A4(n11569), .ZN(
        n11574) );
  NOR2_X1 U14057 ( .A1(n11667), .A2(n11666), .ZN(n11668) );
  AOI21_X1 U14058 ( .B1(n11668), .B2(n11748), .A(n11669), .ZN(n11572) );
  AOI21_X1 U14059 ( .B1(n12255), .B2(n11748), .A(n11744), .ZN(n11571) );
  OAI22_X1 U14060 ( .A1(n11572), .A2(n11571), .B1(n11671), .B2(n11570), .ZN(
        n11573) );
  OAI21_X1 U14061 ( .B1(n11576), .B2(n11575), .A(n11636), .ZN(n11577) );
  NAND2_X1 U14062 ( .A1(n11577), .A2(n11971), .ZN(n11581) );
  AND2_X1 U14063 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n15292) );
  OAI22_X1 U14064 ( .A1(n11979), .A2(n11578), .B1(n11727), .B2(n12000), .ZN(
        n11579) );
  AOI211_X1 U14065 ( .C1(n11997), .C2(n12254), .A(n15292), .B(n11579), .ZN(
        n11580) );
  OAI211_X1 U14066 ( .C1(n11582), .C2(n11985), .A(n11581), .B(n11580), .ZN(
        P3_U3171) );
  NAND2_X1 U14067 ( .A1(n11584), .A2(n11583), .ZN(n11586) );
  XNOR2_X1 U14068 ( .A(n11619), .B(n11618), .ZN(n11587) );
  OAI222_X1 U14069 ( .A1(n14240), .A2(n14085), .B1(n14288), .B2(n13864), .C1(
        n14802), .C2(n11587), .ZN(n14671) );
  INV_X1 U14070 ( .A(n14671), .ZN(n11598) );
  NAND2_X1 U14071 ( .A1(n14658), .A2(n13911), .ZN(n11588) );
  NAND2_X1 U14072 ( .A1(n14676), .A2(n11588), .ZN(n11589) );
  INV_X1 U14073 ( .A(n11589), .ZN(n11591) );
  OR2_X2 U14074 ( .A1(n11589), .A2(n11618), .ZN(n11617) );
  OAI21_X1 U14075 ( .B1(n11591), .B2(n11590), .A(n11617), .ZN(n14673) );
  OAI211_X1 U14076 ( .C1(n6955), .C2(n6956), .A(n14812), .B(n11622), .ZN(
        n14670) );
  OAI22_X1 U14077 ( .A1(n14774), .A2(n11593), .B1(n13903), .B2(n14775), .ZN(
        n11594) );
  AOI21_X1 U14078 ( .B1(n13906), .B2(n14309), .A(n11594), .ZN(n11595) );
  OAI21_X1 U14079 ( .B1(n14670), .B2(n14308), .A(n11595), .ZN(n11596) );
  AOI21_X1 U14080 ( .B1(n14673), .B2(n14828), .A(n11596), .ZN(n11597) );
  OAI21_X1 U14081 ( .B1(n11598), .B2(n14833), .A(n11597), .ZN(P1_U3278) );
  NAND2_X1 U14082 ( .A1(n11600), .A2(n11599), .ZN(n11606) );
  AND2_X1 U14083 ( .A1(n11608), .A2(n11606), .ZN(n11610) );
  NAND2_X1 U14084 ( .A1(n11605), .A2(n13798), .ZN(n11602) );
  NAND2_X1 U14085 ( .A1(n13913), .A2(n9891), .ZN(n11601) );
  NAND2_X1 U14086 ( .A1(n11602), .A2(n11601), .ZN(n11603) );
  XNOR2_X1 U14087 ( .A(n11603), .B(n6549), .ZN(n13681) );
  AND2_X1 U14088 ( .A1(n9892), .A2(n13913), .ZN(n11604) );
  AOI21_X1 U14089 ( .B1(n11605), .B2(n9891), .A(n11604), .ZN(n13682) );
  XNOR2_X1 U14090 ( .A(n13681), .B(n13682), .ZN(n11609) );
  AND2_X1 U14091 ( .A1(n11609), .A2(n11606), .ZN(n11607) );
  NAND2_X1 U14092 ( .A1(n11608), .A2(n11607), .ZN(n13684) );
  OAI211_X1 U14093 ( .C1(n11610), .C2(n11609), .A(n14726), .B(n13684), .ZN(
        n11615) );
  NAND2_X1 U14094 ( .A1(n13901), .A2(n13914), .ZN(n11611) );
  NAND2_X1 U14095 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14754)
         );
  OAI211_X1 U14096 ( .C1(n14662), .C2(n14660), .A(n11611), .B(n14754), .ZN(
        n11612) );
  AOI21_X1 U14097 ( .B1(n11613), .B2(n13891), .A(n11612), .ZN(n11614) );
  OAI211_X1 U14098 ( .C1(n14598), .C2(n14659), .A(n11615), .B(n11614), .ZN(
        P1_U3224) );
  INV_X1 U14099 ( .A(n14661), .ZN(n13910) );
  OR2_X1 U14100 ( .A1(n13906), .A2(n13910), .ZN(n11616) );
  NAND2_X1 U14101 ( .A1(n11617), .A2(n11616), .ZN(n14060) );
  XOR2_X1 U14102 ( .A(n14060), .B(n14083), .Z(n14421) );
  XNOR2_X1 U14103 ( .A(n14084), .B(n14083), .ZN(n14418) );
  INV_X1 U14104 ( .A(n14086), .ZN(n14415) );
  NAND2_X1 U14105 ( .A1(n11622), .A2(n14086), .ZN(n11623) );
  NAND2_X1 U14106 ( .A1(n11623), .A2(n14812), .ZN(n11624) );
  NOR2_X1 U14107 ( .A1(n14307), .A2(n11624), .ZN(n14417) );
  NAND2_X1 U14108 ( .A1(n14417), .A2(n14818), .ZN(n11630) );
  NAND2_X1 U14109 ( .A1(n14088), .A2(n14769), .ZN(n11626) );
  NAND2_X1 U14110 ( .A1(n13910), .A2(n14771), .ZN(n11625) );
  AND2_X1 U14111 ( .A1(n11626), .A2(n11625), .ZN(n14414) );
  INV_X1 U14112 ( .A(n13834), .ZN(n11627) );
  OAI22_X1 U14113 ( .A1(n14315), .A2(n14414), .B1(n11627), .B2(n14775), .ZN(
        n11628) );
  AOI21_X1 U14114 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n14833), .A(n11628), 
        .ZN(n11629) );
  OAI211_X1 U14115 ( .C1(n14415), .C2(n14808), .A(n11630), .B(n11629), .ZN(
        n11631) );
  AOI21_X1 U14116 ( .B1(n14418), .B2(n14829), .A(n11631), .ZN(n11632) );
  OAI21_X1 U14117 ( .B1(n14421), .B2(n14323), .A(n11632), .ZN(P1_U3277) );
  NAND2_X1 U14118 ( .A1(n11751), .A2(n11633), .ZN(n11635) );
  AND2_X1 U14119 ( .A1(n11636), .A2(n11635), .ZN(n11638) );
  XNOR2_X1 U14120 ( .A(n11634), .B(n11036), .ZN(n11712) );
  XNOR2_X1 U14121 ( .A(n11727), .B(n11712), .ZN(n11637) );
  OAI211_X1 U14122 ( .C1(n11638), .C2(n11637), .A(n11971), .B(n11713), .ZN(
        n11642) );
  OAI22_X1 U14123 ( .A1(n11751), .A2(n12008), .B1(n11979), .B2(n15405), .ZN(
        n11639) );
  AOI211_X1 U14124 ( .C1(n12005), .C2(n15304), .A(n11640), .B(n11639), .ZN(
        n11641) );
  OAI211_X1 U14125 ( .C1(n15317), .C2(n11985), .A(n11642), .B(n11641), .ZN(
        P3_U3157) );
  NAND2_X1 U14126 ( .A1(n11658), .A2(n11643), .ZN(n11647) );
  INV_X1 U14127 ( .A(n11644), .ZN(n11645) );
  NAND2_X1 U14128 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n11645), .ZN(n11646) );
  NAND2_X1 U14129 ( .A1(n11647), .A2(n11646), .ZN(n11649) );
  NAND2_X1 U14130 ( .A1(n11648), .A2(n11649), .ZN(n11650) );
  XNOR2_X1 U14131 ( .A(n15013), .B(n11649), .ZN(n15010) );
  NAND2_X1 U14132 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n15010), .ZN(n15008) );
  NAND2_X1 U14133 ( .A1(n11650), .A2(n15008), .ZN(n11653) );
  MUX2_X1 U14134 ( .A(P2_REG2_REG_16__SCAN_IN), .B(n11651), .S(n13005), .Z(
        n11652) );
  NAND2_X1 U14135 ( .A1(n11652), .A2(n11653), .ZN(n13010) );
  OAI211_X1 U14136 ( .C1(n11653), .C2(n11652), .A(n15009), .B(n13010), .ZN(
        n11656) );
  NOR2_X1 U14137 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12862), .ZN(n11654) );
  AOI21_X1 U14138 ( .B1(n15007), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11654), 
        .ZN(n11655) );
  OAI211_X1 U14139 ( .C1(n15014), .C2(n13011), .A(n11656), .B(n11655), .ZN(
        n11664) );
  NOR2_X1 U14140 ( .A1(n11659), .A2(n15013), .ZN(n11660) );
  NOR2_X1 U14141 ( .A1(n15003), .A2(n15004), .ZN(n15002) );
  NOR2_X1 U14142 ( .A1(n11660), .A2(n15002), .ZN(n11662) );
  XNOR2_X1 U14143 ( .A(n13005), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11661) );
  NOR2_X1 U14144 ( .A1(n11662), .A2(n11661), .ZN(n13004) );
  AOI211_X1 U14145 ( .C1(n11662), .C2(n11661), .A(n13004), .B(n15001), .ZN(
        n11663) );
  OR2_X1 U14146 ( .A1(n11664), .A2(n11663), .ZN(P2_U3230) );
  NAND2_X1 U14147 ( .A1(n6656), .A2(n11665), .ZN(n11683) );
  XNOR2_X1 U14148 ( .A(n11667), .B(n11666), .ZN(n11684) );
  NOR2_X1 U14149 ( .A1(n11683), .A2(n11684), .ZN(n11682) );
  NOR2_X1 U14150 ( .A1(n11682), .A2(n11668), .ZN(n11745) );
  XNOR2_X1 U14151 ( .A(n11745), .B(n11669), .ZN(n11676) );
  AND2_X1 U14152 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n15251) );
  OAI22_X1 U14153 ( .A1(n11671), .A2(n12000), .B1(n11979), .B2(n11670), .ZN(
        n11672) );
  AOI211_X1 U14154 ( .C1(n11997), .C2(n12256), .A(n15251), .B(n11672), .ZN(
        n11675) );
  NAND2_X1 U14155 ( .A1(n12004), .A2(n11673), .ZN(n11674) );
  OAI211_X1 U14156 ( .C1(n11676), .C2(n12014), .A(n11675), .B(n11674), .ZN(
        P3_U3153) );
  INV_X1 U14157 ( .A(n11677), .ZN(n11679) );
  OAI222_X1 U14158 ( .A1(n14574), .A2(n11680), .B1(n14576), .B2(n11679), .C1(
        P3_U3151), .C2(n11678), .ZN(P3_U3270) );
  INV_X1 U14159 ( .A(n11681), .ZN(n11691) );
  AOI211_X1 U14160 ( .C1(n11684), .C2(n11683), .A(n12014), .B(n11682), .ZN(
        n11685) );
  INV_X1 U14161 ( .A(n11685), .ZN(n11690) );
  INV_X1 U14162 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n11686) );
  NOR2_X1 U14163 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11686), .ZN(n15233) );
  OAI22_X1 U14164 ( .A1(n11687), .A2(n11979), .B1(n11746), .B2(n12000), .ZN(
        n11688) );
  AOI211_X1 U14165 ( .C1(n11997), .C2(n12257), .A(n15233), .B(n11688), .ZN(
        n11689) );
  OAI211_X1 U14166 ( .C1(n11691), .C2(n11985), .A(n11690), .B(n11689), .ZN(
        P3_U3179) );
  INV_X1 U14167 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13641) );
  AOI21_X2 U14168 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n14580), .A(n11692), 
        .ZN(n12260) );
  XNOR2_X1 U14169 ( .A(n12260), .B(n6802), .ZN(n11693) );
  NOR2_X1 U14170 ( .A1(n13641), .A2(n11693), .ZN(n12261) );
  AOI21_X1 U14171 ( .B1(n13641), .B2(n11693), .A(n12261), .ZN(n11711) );
  NAND2_X1 U14172 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n11695), .ZN(n12274) );
  OAI21_X1 U14173 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n11695), .A(n12274), 
        .ZN(n11709) );
  AND2_X1 U14174 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n11981) );
  AOI21_X1 U14175 ( .B1(n15293), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n11981), 
        .ZN(n11696) );
  OAI21_X1 U14176 ( .B1(n15290), .B2(n12273), .A(n11696), .ZN(n11708) );
  MUX2_X1 U14177 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12774), .Z(n12264) );
  XNOR2_X1 U14178 ( .A(n12264), .B(n12273), .ZN(n11702) );
  INV_X1 U14179 ( .A(n11697), .ZN(n11699) );
  NOR2_X1 U14180 ( .A1(n11699), .A2(n11698), .ZN(n11703) );
  INV_X1 U14181 ( .A(n12265), .ZN(n11706) );
  OAI21_X1 U14182 ( .B1(n11704), .B2(n11703), .A(n11702), .ZN(n11705) );
  AOI21_X1 U14183 ( .B1(n11706), .B2(n11705), .A(n15176), .ZN(n11707) );
  AOI211_X1 U14184 ( .C1(n15296), .C2(n11709), .A(n11708), .B(n11707), .ZN(
        n11710) );
  OAI21_X1 U14185 ( .B1(n11711), .B2(n15300), .A(n11710), .ZN(P3_U3195) );
  INV_X1 U14186 ( .A(n11712), .ZN(n11714) );
  OAI21_X1 U14187 ( .B1(n11727), .B2(n11714), .A(n11713), .ZN(n11784) );
  XNOR2_X1 U14188 ( .A(n11036), .B(n11731), .ZN(n11781) );
  XNOR2_X1 U14189 ( .A(n11791), .B(n11781), .ZN(n11715) );
  XNOR2_X1 U14190 ( .A(n11784), .B(n11715), .ZN(n11723) );
  NAND2_X1 U14191 ( .A1(n12004), .A2(n11732), .ZN(n11721) );
  AOI21_X1 U14192 ( .B1(n12252), .B2(n12005), .A(n11716), .ZN(n11720) );
  NAND2_X1 U14193 ( .A1(n12018), .A2(n11717), .ZN(n11719) );
  NAND2_X1 U14194 ( .A1(n12253), .A2(n11997), .ZN(n11718) );
  NAND4_X1 U14195 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11722) );
  AOI21_X1 U14196 ( .B1(n11723), .B2(n11971), .A(n11722), .ZN(n11724) );
  INV_X1 U14197 ( .A(n11724), .ZN(P3_U3176) );
  XNOR2_X1 U14198 ( .A(n11725), .B(n12135), .ZN(n11726) );
  NAND2_X1 U14199 ( .A1(n11726), .A2(n15323), .ZN(n11730) );
  OAI22_X1 U14200 ( .A1(n11727), .A2(n15340), .B1(n11799), .B2(n15338), .ZN(
        n11728) );
  INV_X1 U14201 ( .A(n11728), .ZN(n11729) );
  NAND2_X1 U14202 ( .A1(n11730), .A2(n11729), .ZN(n14637) );
  INV_X1 U14203 ( .A(n14637), .ZN(n11736) );
  NAND2_X1 U14204 ( .A1(n12562), .A2(n12135), .ZN(n11757) );
  OAI21_X1 U14205 ( .B1(n12562), .B2(n12135), .A(n11757), .ZN(n14639) );
  AOI21_X2 U14206 ( .B1(n15328), .B2(n15357), .A(n15371), .ZN(n12595) );
  NOR2_X1 U14207 ( .A1(n11731), .A2(n15406), .ZN(n14638) );
  AOI22_X1 U14208 ( .A1(n15333), .A2(n14638), .B1(n15365), .B2(n11732), .ZN(
        n11733) );
  OAI21_X1 U14209 ( .B1(n7671), .B2(n15369), .A(n11733), .ZN(n11734) );
  AOI21_X1 U14210 ( .B1(n14639), .B2(n12595), .A(n11734), .ZN(n11735) );
  OAI21_X1 U14211 ( .B1(n11736), .B2(n15371), .A(n11735), .ZN(P3_U3222) );
  INV_X1 U14212 ( .A(n11737), .ZN(n11742) );
  INV_X1 U14213 ( .A(n11738), .ZN(n11740) );
  OAI222_X1 U14214 ( .A1(n13393), .A2(n11742), .B1(n11740), .B2(P2_U3088), 
        .C1(n11739), .C2(n13395), .ZN(P2_U3303) );
  OAI222_X1 U14215 ( .A1(n11743), .A2(P1_U3086), .B1(n14458), .B2(n11742), 
        .C1(n11741), .C2(n14455), .ZN(P1_U3331) );
  MUX2_X1 U14216 ( .A(n11746), .B(n11745), .S(n11744), .Z(n11747) );
  XOR2_X1 U14217 ( .A(n11748), .B(n11747), .Z(n11756) );
  NOR2_X1 U14218 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11749), .ZN(n15270) );
  OAI22_X1 U14219 ( .A1(n11751), .A2(n12000), .B1(n11979), .B2(n11750), .ZN(
        n11752) );
  AOI211_X1 U14220 ( .C1(n11997), .C2(n12255), .A(n15270), .B(n11752), .ZN(
        n11755) );
  NAND2_X1 U14221 ( .A1(n12004), .A2(n11753), .ZN(n11754) );
  OAI211_X1 U14222 ( .C1(n11756), .C2(n12014), .A(n11755), .B(n11754), .ZN(
        P3_U3161) );
  NAND2_X1 U14223 ( .A1(n11757), .A2(n12137), .ZN(n11758) );
  INV_X1 U14224 ( .A(n11761), .ZN(n12050) );
  XNOR2_X1 U14225 ( .A(n11758), .B(n12050), .ZN(n14635) );
  INV_X1 U14226 ( .A(n14635), .ZN(n11769) );
  INV_X1 U14227 ( .A(n12595), .ZN(n12625) );
  NAND2_X1 U14228 ( .A1(n11760), .A2(n11759), .ZN(n11762) );
  XNOR2_X1 U14229 ( .A(n11762), .B(n11761), .ZN(n11763) );
  OAI222_X1 U14230 ( .A1(n15338), .A2(n11810), .B1(n15340), .B2(n11791), .C1(
        n11763), .C2(n15347), .ZN(n14633) );
  NAND2_X1 U14231 ( .A1(n14633), .A2(n15369), .ZN(n11768) );
  NOR2_X1 U14232 ( .A1(n11785), .A2(n15406), .ZN(n14634) );
  INV_X1 U14233 ( .A(n11764), .ZN(n11796) );
  OAI22_X1 U14234 ( .A1(n15369), .A2(n11765), .B1(n11796), .B2(n15316), .ZN(
        n11766) );
  AOI21_X1 U14235 ( .B1(n15333), .B2(n14634), .A(n11766), .ZN(n11767) );
  OAI211_X1 U14236 ( .C1(n11769), .C2(n12625), .A(n11768), .B(n11767), .ZN(
        P3_U3221) );
  NOR2_X1 U14237 ( .A1(n11770), .A2(n12140), .ZN(n12131) );
  XNOR2_X1 U14238 ( .A(n11771), .B(n12131), .ZN(n11772) );
  AOI222_X1 U14239 ( .A1(n15323), .A2(n11772), .B1(n11982), .B2(n15319), .C1(
        n12252), .C2(n15321), .ZN(n14628) );
  INV_X1 U14240 ( .A(n11773), .ZN(n11986) );
  OAI22_X1 U14241 ( .A1(n15369), .A2(n13641), .B1(n11986), .B2(n15316), .ZN(
        n11774) );
  AOI21_X1 U14242 ( .B1(n14619), .B2(n11994), .A(n11774), .ZN(n11780) );
  NAND2_X1 U14243 ( .A1(n12562), .A2(n11775), .ZN(n11777) );
  NAND2_X1 U14244 ( .A1(n11777), .A2(n11776), .ZN(n11778) );
  XNOR2_X1 U14245 ( .A(n11778), .B(n12131), .ZN(n14631) );
  NAND2_X1 U14246 ( .A1(n14631), .A2(n12595), .ZN(n11779) );
  OAI211_X1 U14247 ( .C1(n14628), .C2(n15371), .A(n11780), .B(n11779), .ZN(
        P3_U3220) );
  NAND2_X1 U14248 ( .A1(n11791), .A2(n11781), .ZN(n11783) );
  INV_X1 U14249 ( .A(n11781), .ZN(n11782) );
  AOI21_X2 U14250 ( .B1(n11784), .B2(n11783), .A(n7423), .ZN(n11787) );
  XNOR2_X1 U14251 ( .A(n11785), .B(n11898), .ZN(n11797) );
  XNOR2_X1 U14252 ( .A(n11797), .B(n11799), .ZN(n11786) );
  OAI21_X1 U14253 ( .B1(n11787), .B2(n11786), .A(n11989), .ZN(n11788) );
  NAND2_X1 U14254 ( .A1(n11788), .A2(n11971), .ZN(n11795) );
  AOI21_X1 U14255 ( .B1(n12618), .B2(n12005), .A(n11789), .ZN(n11790) );
  OAI21_X1 U14256 ( .B1(n11791), .B2(n12008), .A(n11790), .ZN(n11792) );
  AOI21_X1 U14257 ( .B1(n12018), .B2(n11793), .A(n11792), .ZN(n11794) );
  OAI211_X1 U14258 ( .C1(n11796), .C2(n11985), .A(n11795), .B(n11794), .ZN(
        P3_U3164) );
  XNOR2_X1 U14259 ( .A(n11994), .B(n11898), .ZN(n11801) );
  XNOR2_X1 U14260 ( .A(n11801), .B(n12618), .ZN(n11987) );
  INV_X1 U14261 ( .A(n11797), .ZN(n11798) );
  NAND2_X1 U14262 ( .A1(n11799), .A2(n11798), .ZN(n11988) );
  XNOR2_X1 U14263 ( .A(n11800), .B(n11901), .ZN(n11824) );
  XNOR2_X1 U14264 ( .A(n11824), .B(n11982), .ZN(n11805) );
  INV_X1 U14265 ( .A(n11801), .ZN(n11802) );
  NAND2_X1 U14266 ( .A1(n11802), .A2(n12618), .ZN(n11806) );
  INV_X1 U14267 ( .A(n11825), .ZN(n11808) );
  AOI21_X1 U14268 ( .B1(n11804), .B2(n11806), .A(n11805), .ZN(n11807) );
  OAI21_X1 U14269 ( .B1(n11808), .B2(n11807), .A(n11971), .ZN(n11813) );
  INV_X1 U14270 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n13591) );
  NOR2_X1 U14271 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n13591), .ZN(n12278) );
  AOI21_X1 U14272 ( .B1(n12617), .B2(n12005), .A(n12278), .ZN(n11809) );
  OAI21_X1 U14273 ( .B1(n11810), .B2(n12008), .A(n11809), .ZN(n11811) );
  AOI21_X1 U14274 ( .B1(n12621), .B2(n12004), .A(n11811), .ZN(n11812) );
  OAI211_X1 U14275 ( .C1(n11979), .C2(n12761), .A(n11813), .B(n11812), .ZN(
        P3_U3155) );
  INV_X1 U14276 ( .A(n9458), .ZN(n11815) );
  OAI222_X1 U14277 ( .A1(n9580), .A2(P1_U3086), .B1(n14458), .B2(n11815), .C1(
        n11814), .C2(n14455), .ZN(P1_U3327) );
  OAI222_X1 U14278 ( .A1(n9905), .A2(P1_U3086), .B1(n14458), .B2(n13390), .C1(
        n11816), .C2(n14455), .ZN(P1_U3329) );
  INV_X1 U14279 ( .A(n11817), .ZN(n11818) );
  OAI222_X1 U14280 ( .A1(n14574), .A2(n11820), .B1(P3_U3151), .B2(n11819), 
        .C1(n14576), .C2(n11818), .ZN(P3_U3267) );
  INV_X1 U14281 ( .A(n11821), .ZN(n14451) );
  OAI222_X1 U14282 ( .A1(n13393), .A2(n14451), .B1(n11823), .B2(P2_U3088), 
        .C1(n11822), .C2(n13395), .ZN(P2_U3298) );
  XNOR2_X1 U14283 ( .A(n12608), .B(n11036), .ZN(n11826) );
  NOR2_X1 U14284 ( .A1(n11826), .A2(n12617), .ZN(n12009) );
  NAND2_X1 U14285 ( .A1(n11826), .A2(n12617), .ZN(n12010) );
  OAI21_X1 U14286 ( .B1(n12013), .B2(n12009), .A(n12010), .ZN(n11958) );
  XNOR2_X1 U14287 ( .A(n11955), .B(n11901), .ZN(n11827) );
  XNOR2_X1 U14288 ( .A(n11827), .B(n12251), .ZN(n11957) );
  NAND2_X1 U14289 ( .A1(n11958), .A2(n11957), .ZN(n11956) );
  NAND2_X1 U14290 ( .A1(n11956), .A2(n11828), .ZN(n11876) );
  XNOR2_X1 U14291 ( .A(n12749), .B(n11901), .ZN(n11829) );
  XNOR2_X1 U14292 ( .A(n11829), .B(n12554), .ZN(n11875) );
  NAND2_X1 U14293 ( .A1(n11876), .A2(n11875), .ZN(n11874) );
  NAND2_X1 U14294 ( .A1(n11829), .A2(n12580), .ZN(n11830) );
  NAND2_X1 U14295 ( .A1(n11874), .A2(n11830), .ZN(n11869) );
  XNOR2_X1 U14296 ( .A(n12745), .B(n11898), .ZN(n11831) );
  XNOR2_X1 U14297 ( .A(n11831), .B(n12572), .ZN(n11868) );
  NAND2_X1 U14298 ( .A1(n11869), .A2(n11868), .ZN(n11867) );
  NAND2_X1 U14299 ( .A1(n11831), .A2(n12537), .ZN(n11832) );
  NAND2_X1 U14300 ( .A1(n11867), .A2(n11832), .ZN(n11928) );
  XNOR2_X1 U14301 ( .A(n11933), .B(n11898), .ZN(n11833) );
  XOR2_X1 U14302 ( .A(n12520), .B(n11833), .Z(n11927) );
  NAND2_X1 U14303 ( .A1(n11928), .A2(n11927), .ZN(n11926) );
  NAND2_X1 U14304 ( .A1(n11833), .A2(n12520), .ZN(n11834) );
  NAND2_X1 U14305 ( .A1(n11926), .A2(n11834), .ZN(n11974) );
  XNOR2_X1 U14306 ( .A(n11980), .B(n11898), .ZN(n11835) );
  XNOR2_X1 U14307 ( .A(n11835), .B(n11940), .ZN(n11973) );
  NAND2_X1 U14308 ( .A1(n11974), .A2(n11973), .ZN(n11972) );
  NAND2_X1 U14309 ( .A1(n11835), .A2(n12536), .ZN(n11836) );
  XNOR2_X1 U14310 ( .A(n12514), .B(n11898), .ZN(n11837) );
  XNOR2_X1 U14311 ( .A(n11837), .B(n12522), .ZN(n11937) );
  NAND2_X1 U14312 ( .A1(n11837), .A2(n12522), .ZN(n11838) );
  XNOR2_X1 U14313 ( .A(n12501), .B(n11036), .ZN(n11839) );
  INV_X1 U14314 ( .A(n11839), .ZN(n11840) );
  XNOR2_X1 U14315 ( .A(n11844), .B(n11036), .ZN(n11845) );
  NAND2_X1 U14316 ( .A1(n11919), .A2(n12500), .ZN(n11849) );
  INV_X1 U14317 ( .A(n11845), .ZN(n11846) );
  OR2_X1 U14318 ( .A1(n11847), .A2(n11846), .ZN(n11848) );
  XNOR2_X1 U14319 ( .A(n12721), .B(n11898), .ZN(n11850) );
  XNOR2_X1 U14320 ( .A(n11850), .B(n11922), .ZN(n11964) );
  NAND2_X1 U14321 ( .A1(n11963), .A2(n11964), .ZN(n11947) );
  INV_X1 U14322 ( .A(n11850), .ZN(n11851) );
  NAND2_X1 U14323 ( .A1(n11851), .A2(n11922), .ZN(n11946) );
  XNOR2_X1 U14324 ( .A(n12717), .B(n11898), .ZN(n11852) );
  NAND2_X1 U14325 ( .A1(n11852), .A2(n12468), .ZN(n11882) );
  INV_X1 U14326 ( .A(n11882), .ZN(n11853) );
  XNOR2_X1 U14327 ( .A(n11852), .B(n12470), .ZN(n11949) );
  OR2_X1 U14328 ( .A1(n11853), .A2(n11949), .ZN(n11854) );
  XNOR2_X1 U14329 ( .A(n12438), .B(n11898), .ZN(n11881) );
  XNOR2_X1 U14330 ( .A(n11881), .B(n12448), .ZN(n11885) );
  AOI22_X1 U14331 ( .A1(n12470), .A2(n11997), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11856) );
  NAND2_X1 U14332 ( .A1(n12004), .A2(n12439), .ZN(n11855) );
  OAI211_X1 U14333 ( .C1(n11906), .C2(n12000), .A(n11856), .B(n11855), .ZN(
        n11857) );
  AOI21_X1 U14334 ( .B1(n12438), .B2(n12018), .A(n11857), .ZN(n11858) );
  OAI21_X1 U14335 ( .B1(n11861), .B2(n11860), .A(n11859), .ZN(n11862) );
  NAND2_X1 U14336 ( .A1(n11862), .A2(n12946), .ZN(n11866) );
  AOI22_X1 U14337 ( .A1(n12950), .A2(n11864), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n11863), .ZN(n11865) );
  OAI211_X1 U14338 ( .C1(n8841), .C2(n12926), .A(n11866), .B(n11865), .ZN(
        P2_U3194) );
  OAI211_X1 U14339 ( .C1(n11869), .C2(n11868), .A(n11867), .B(n11971), .ZN(
        n11873) );
  INV_X1 U14340 ( .A(n12520), .ZN(n12555) );
  NAND2_X1 U14341 ( .A1(n11997), .A2(n12580), .ZN(n11870) );
  NAND2_X1 U14342 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12358)
         );
  OAI211_X1 U14343 ( .C1(n12555), .C2(n12000), .A(n11870), .B(n12358), .ZN(
        n11871) );
  AOI21_X1 U14344 ( .B1(n12556), .B2(n12004), .A(n11871), .ZN(n11872) );
  OAI211_X1 U14345 ( .C1(n12745), .C2(n11979), .A(n11873), .B(n11872), .ZN(
        P3_U3178) );
  OAI211_X1 U14346 ( .C1(n11876), .C2(n11875), .A(n11874), .B(n11971), .ZN(
        n11880) );
  NAND2_X1 U14347 ( .A1(n12251), .A2(n11997), .ZN(n11877) );
  NAND2_X1 U14348 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12332)
         );
  OAI211_X1 U14349 ( .C1(n12572), .C2(n12000), .A(n11877), .B(n12332), .ZN(
        n11878) );
  AOI21_X1 U14350 ( .B1(n12573), .B2(n12004), .A(n11878), .ZN(n11879) );
  OAI211_X1 U14351 ( .C1(n12749), .C2(n11979), .A(n11880), .B(n11879), .ZN(
        P3_U3168) );
  NAND2_X1 U14352 ( .A1(n11881), .A2(n12416), .ZN(n11884) );
  AND2_X1 U14353 ( .A1(n11882), .A2(n11884), .ZN(n11891) );
  INV_X1 U14354 ( .A(n11891), .ZN(n11883) );
  OR2_X1 U14355 ( .A1(n11883), .A2(n11949), .ZN(n11890) );
  AND2_X1 U14356 ( .A1(n11964), .A2(n11890), .ZN(n11887) );
  INV_X1 U14357 ( .A(n11884), .ZN(n11886) );
  OR2_X1 U14358 ( .A1(n11886), .A2(n11885), .ZN(n11889) );
  AND2_X1 U14359 ( .A1(n11887), .A2(n11889), .ZN(n11888) );
  INV_X1 U14360 ( .A(n11889), .ZN(n11895) );
  INV_X1 U14361 ( .A(n11890), .ZN(n11893) );
  AND2_X1 U14362 ( .A1(n11946), .A2(n11891), .ZN(n11892) );
  OR2_X1 U14363 ( .A1(n11893), .A2(n11892), .ZN(n11894) );
  OR2_X1 U14364 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  XNOR2_X1 U14365 ( .A(n12202), .B(n11898), .ZN(n11899) );
  XNOR2_X1 U14366 ( .A(n11899), .B(n12434), .ZN(n11912) );
  AND2_X1 U14367 ( .A1(n11899), .A2(n11906), .ZN(n11900) );
  XNOR2_X1 U14368 ( .A(n6779), .B(n11901), .ZN(n11902) );
  XNOR2_X1 U14369 ( .A(n11903), .B(n11902), .ZN(n11911) );
  INV_X1 U14370 ( .A(n11904), .ZN(n12405) );
  OAI22_X1 U14371 ( .A1(n11906), .A2(n12008), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11905), .ZN(n11907) );
  AOI21_X1 U14372 ( .B1(n12005), .B2(n12248), .A(n11907), .ZN(n11908) );
  OAI21_X1 U14373 ( .B1(n12405), .B2(n11985), .A(n11908), .ZN(n11909) );
  AOI21_X1 U14374 ( .B1(n12407), .B2(n12018), .A(n11909), .ZN(n11910) );
  OAI21_X1 U14375 ( .B1(n11911), .B2(n12014), .A(n11910), .ZN(P3_U3160) );
  XNOR2_X1 U14376 ( .A(n11913), .B(n11912), .ZN(n11914) );
  NAND2_X1 U14377 ( .A1(n11914), .A2(n11971), .ZN(n11918) );
  INV_X1 U14378 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n13588) );
  OAI22_X1 U14379 ( .A1(n12416), .A2(n12008), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13588), .ZN(n11916) );
  NOR2_X1 U14380 ( .A1(n12417), .A2(n12000), .ZN(n11915) );
  AOI211_X1 U14381 ( .C1(n12422), .C2(n12004), .A(n11916), .B(n11915), .ZN(
        n11917) );
  OAI211_X1 U14382 ( .C1(n12711), .C2(n11979), .A(n11918), .B(n11917), .ZN(
        P3_U3154) );
  XNOR2_X1 U14383 ( .A(n11919), .B(n12249), .ZN(n11925) );
  AOI22_X1 U14384 ( .A1(n11997), .A2(n12509), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11921) );
  NAND2_X1 U14385 ( .A1(n12004), .A2(n12487), .ZN(n11920) );
  OAI211_X1 U14386 ( .C1(n11922), .C2(n12000), .A(n11921), .B(n11920), .ZN(
        n11923) );
  AOI21_X1 U14387 ( .B1(n12724), .B2(n12018), .A(n11923), .ZN(n11924) );
  OAI21_X1 U14388 ( .B1(n11925), .B2(n12014), .A(n11924), .ZN(P3_U3156) );
  OAI211_X1 U14389 ( .C1(n11928), .C2(n11927), .A(n11926), .B(n11971), .ZN(
        n11932) );
  NAND2_X1 U14390 ( .A1(n12536), .A2(n12005), .ZN(n11929) );
  NAND2_X1 U14391 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12390)
         );
  OAI211_X1 U14392 ( .C1(n12572), .C2(n12008), .A(n11929), .B(n12390), .ZN(
        n11930) );
  AOI21_X1 U14393 ( .B1(n12542), .B2(n12004), .A(n11930), .ZN(n11931) );
  OAI211_X1 U14394 ( .C1(n11979), .C2(n11933), .A(n11932), .B(n11931), .ZN(
        P3_U3159) );
  INV_X1 U14395 ( .A(n11934), .ZN(n11935) );
  AOI21_X1 U14396 ( .B1(n11937), .B2(n11936), .A(n11935), .ZN(n11945) );
  INV_X1 U14397 ( .A(n11938), .ZN(n12511) );
  OAI22_X1 U14398 ( .A1(n11940), .A2(n12008), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11939), .ZN(n11941) );
  AOI21_X1 U14399 ( .B1(n12005), .B2(n12509), .A(n11941), .ZN(n11942) );
  OAI21_X1 U14400 ( .B1(n12511), .B2(n11985), .A(n11942), .ZN(n11943) );
  AOI21_X1 U14401 ( .B1(n12514), .B2(n12018), .A(n11943), .ZN(n11944) );
  OAI21_X1 U14402 ( .B1(n11945), .B2(n12014), .A(n11944), .ZN(P3_U3163) );
  NAND2_X1 U14403 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  XOR2_X1 U14404 ( .A(n11949), .B(n11948), .Z(n11954) );
  AOI22_X1 U14405 ( .A1(n12484), .A2(n11997), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11951) );
  NAND2_X1 U14406 ( .A1(n12004), .A2(n12455), .ZN(n11950) );
  OAI211_X1 U14407 ( .C1(n12416), .C2(n12000), .A(n11951), .B(n11950), .ZN(
        n11952) );
  AOI21_X1 U14408 ( .B1(n12717), .B2(n12018), .A(n11952), .ZN(n11953) );
  OAI21_X1 U14409 ( .B1(n11954), .B2(n12014), .A(n11953), .ZN(P3_U3165) );
  OAI211_X1 U14410 ( .C1(n11958), .C2(n11957), .A(n11956), .B(n11971), .ZN(
        n11962) );
  NAND2_X1 U14411 ( .A1(n11997), .A2(n12617), .ZN(n11959) );
  NAND2_X1 U14412 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12315)
         );
  OAI211_X1 U14413 ( .C1(n12554), .C2(n12000), .A(n11959), .B(n12315), .ZN(
        n11960) );
  AOI21_X1 U14414 ( .B1(n12592), .B2(n12004), .A(n11960), .ZN(n11961) );
  OAI211_X1 U14415 ( .C1(n12753), .C2(n11979), .A(n11962), .B(n11961), .ZN(
        P3_U3166) );
  XOR2_X1 U14416 ( .A(n11964), .B(n11963), .Z(n11970) );
  AOI22_X1 U14417 ( .A1(n12249), .A2(n11997), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11966) );
  NAND2_X1 U14418 ( .A1(n12004), .A2(n12475), .ZN(n11965) );
  OAI211_X1 U14419 ( .C1(n12468), .C2(n12000), .A(n11966), .B(n11965), .ZN(
        n11967) );
  AOI21_X1 U14420 ( .B1(n11968), .B2(n12018), .A(n11967), .ZN(n11969) );
  OAI21_X1 U14421 ( .B1(n11970), .B2(n12014), .A(n11969), .ZN(P3_U3169) );
  OAI211_X1 U14422 ( .C1(n11974), .C2(n11973), .A(n11972), .B(n11971), .ZN(
        n11978) );
  AOI22_X1 U14423 ( .A1(n11997), .A2(n12520), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11975) );
  OAI21_X1 U14424 ( .B1(n12522), .B2(n12000), .A(n11975), .ZN(n11976) );
  AOI21_X1 U14425 ( .B1(n12525), .B2(n12004), .A(n11976), .ZN(n11977) );
  OAI211_X1 U14426 ( .C1(n11980), .C2(n11979), .A(n11978), .B(n11977), .ZN(
        P3_U3173) );
  AOI21_X1 U14427 ( .B1(n11982), .B2(n12005), .A(n11981), .ZN(n11984) );
  NAND2_X1 U14428 ( .A1(n12252), .A2(n11997), .ZN(n11983) );
  OAI211_X1 U14429 ( .C1(n11986), .C2(n11985), .A(n11984), .B(n11983), .ZN(
        n11993) );
  INV_X1 U14430 ( .A(n11804), .ZN(n11991) );
  AOI21_X1 U14431 ( .B1(n11989), .B2(n11988), .A(n11987), .ZN(n11990) );
  NOR3_X1 U14432 ( .A1(n11991), .A2(n11990), .A3(n12014), .ZN(n11992) );
  AOI211_X1 U14433 ( .C1(n12018), .C2(n11994), .A(n11993), .B(n11992), .ZN(
        n11995) );
  INV_X1 U14434 ( .A(n11995), .ZN(P3_U3174) );
  XNOR2_X1 U14435 ( .A(n11996), .B(n12509), .ZN(n12003) );
  INV_X1 U14436 ( .A(n12522), .ZN(n12250) );
  AOI22_X1 U14437 ( .A1(n12250), .A2(n11997), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11999) );
  NAND2_X1 U14438 ( .A1(n12004), .A2(n12502), .ZN(n11998) );
  OAI211_X1 U14439 ( .C1(n12500), .C2(n12000), .A(n11999), .B(n11998), .ZN(
        n12001) );
  AOI21_X1 U14440 ( .B1(n12501), .B2(n12018), .A(n12001), .ZN(n12002) );
  OAI21_X1 U14441 ( .B1(n12003), .B2(n12014), .A(n12002), .ZN(P3_U3175) );
  NAND2_X1 U14442 ( .A1(n12004), .A2(n12609), .ZN(n12007) );
  AND2_X1 U14443 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12291) );
  AOI21_X1 U14444 ( .B1(n12251), .B2(n12005), .A(n12291), .ZN(n12006) );
  OAI211_X1 U14445 ( .C1(n12606), .C2(n12008), .A(n12007), .B(n12006), .ZN(
        n12017) );
  INV_X1 U14446 ( .A(n12009), .ZN(n12011) );
  NAND2_X1 U14447 ( .A1(n12011), .A2(n12010), .ZN(n12012) );
  XNOR2_X1 U14448 ( .A(n12013), .B(n12012), .ZN(n12015) );
  NOR2_X1 U14449 ( .A1(n12015), .A2(n12014), .ZN(n12016) );
  AOI211_X1 U14450 ( .C1(n12018), .C2(n12608), .A(n12017), .B(n12016), .ZN(
        n12019) );
  INV_X1 U14451 ( .A(n12019), .ZN(P3_U3181) );
  INV_X1 U14452 ( .A(n12020), .ZN(n12240) );
  OAI21_X1 U14453 ( .B1(P2_DATAO_REG_30__SCAN_IN), .B2(n13488), .A(n12031), 
        .ZN(n12023) );
  NAND2_X1 U14454 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n13488), .ZN(n12030) );
  NAND2_X1 U14455 ( .A1(n12023), .A2(n12030), .ZN(n12026) );
  INV_X1 U14456 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n13374) );
  INV_X1 U14457 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12024) );
  AOI22_X1 U14458 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n13374), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n12024), .ZN(n12025) );
  XNOR2_X1 U14459 ( .A(n12026), .B(n12025), .ZN(n12763) );
  NAND2_X1 U14460 ( .A1(n12763), .A2(n12027), .ZN(n12029) );
  OR2_X1 U14461 ( .A1(n12033), .A2(n12767), .ZN(n12028) );
  OAI21_X1 U14462 ( .B1(n13488), .B2(P2_DATAO_REG_30__SCAN_IN), .A(n12030), 
        .ZN(n12032) );
  XNOR2_X1 U14463 ( .A(n12032), .B(n12031), .ZN(n12768) );
  OR2_X1 U14464 ( .A1(n12033), .A2(n13654), .ZN(n12034) );
  INV_X1 U14465 ( .A(n12039), .ZN(n14616) );
  NAND2_X1 U14466 ( .A1(n14626), .A2(n12037), .ZN(n12220) );
  INV_X1 U14467 ( .A(n12220), .ZN(n12038) );
  AOI21_X1 U14468 ( .B1(n14616), .B2(n14626), .A(n12038), .ZN(n12040) );
  NAND2_X1 U14469 ( .A1(n12042), .A2(n12039), .ZN(n12232) );
  INV_X1 U14470 ( .A(n12042), .ZN(n14622) );
  AND2_X1 U14471 ( .A1(n14622), .A2(n14616), .ZN(n12060) );
  INV_X1 U14472 ( .A(n12060), .ZN(n12229) );
  OAI211_X1 U14473 ( .C1(n12042), .C2(n12221), .A(n12041), .B(n12229), .ZN(
        n12043) );
  XNOR2_X1 U14474 ( .A(n12043), .B(n12375), .ZN(n12239) );
  NAND2_X1 U14475 ( .A1(n12198), .A2(n12197), .ZN(n12065) );
  INV_X1 U14476 ( .A(n12516), .ZN(n12178) );
  NAND4_X1 U14477 ( .A1(n12045), .A2(n12044), .A3(n7919), .A4(n12118), .ZN(
        n12047) );
  INV_X1 U14478 ( .A(n15306), .ZN(n12125) );
  NAND4_X1 U14479 ( .A1(n12097), .A2(n12108), .A3(n12125), .A4(n12113), .ZN(
        n12046) );
  NOR2_X1 U14480 ( .A1(n12047), .A2(n12046), .ZN(n12051) );
  AND4_X1 U14481 ( .A1(n15345), .A2(n12048), .A3(n12092), .A4(n12135), .ZN(
        n12049) );
  AND4_X1 U14482 ( .A1(n12051), .A2(n12050), .A3(n12131), .A4(n12049), .ZN(
        n12052) );
  NAND4_X1 U14483 ( .A1(n12052), .A2(n12600), .A3(n12588), .A4(n12615), .ZN(
        n12053) );
  NOR2_X1 U14484 ( .A1(n12569), .A2(n12053), .ZN(n12054) );
  NAND3_X1 U14485 ( .A1(n12540), .A2(n12552), .A3(n12054), .ZN(n12055) );
  NOR2_X1 U14486 ( .A1(n12171), .A2(n12055), .ZN(n12056) );
  AND4_X1 U14487 ( .A1(n12474), .A2(n12178), .A3(n12497), .A4(n12056), .ZN(
        n12057) );
  NAND4_X1 U14488 ( .A1(n12413), .A2(n12451), .A3(n12480), .A4(n12057), .ZN(
        n12058) );
  NOR2_X1 U14489 ( .A1(n12065), .A2(n12058), .ZN(n12059) );
  NAND3_X1 U14490 ( .A1(n12232), .A2(n6779), .A3(n12059), .ZN(n12061) );
  NAND2_X1 U14491 ( .A1(n12221), .A2(n12220), .ZN(n12206) );
  XNOR2_X1 U14492 ( .A(n12062), .B(n12391), .ZN(n12064) );
  MUX2_X1 U14493 ( .A(n12067), .B(n12066), .S(n12219), .Z(n12196) );
  NAND2_X1 U14494 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  NAND2_X1 U14495 ( .A1(n12070), .A2(n12071), .ZN(n12072) );
  MUX2_X1 U14496 ( .A(n12072), .B(n12071), .S(n12227), .Z(n12194) );
  NAND2_X1 U14497 ( .A1(n12073), .A2(n12227), .ZN(n12077) );
  OAI22_X1 U14498 ( .A1(n12701), .A2(n12074), .B1(n12244), .B2(n12073), .ZN(
        n12075) );
  NAND2_X1 U14499 ( .A1(n12075), .A2(n12081), .ZN(n12076) );
  INV_X1 U14500 ( .A(n12078), .ZN(n12080) );
  OAI211_X1 U14501 ( .C1(n12083), .C2(n12080), .A(n12086), .B(n12079), .ZN(
        n12090) );
  INV_X1 U14502 ( .A(n12081), .ZN(n12082) );
  OR2_X1 U14503 ( .A1(n12083), .A2(n12082), .ZN(n12089) );
  AND2_X1 U14504 ( .A1(n12085), .A2(n12084), .ZN(n12088) );
  INV_X1 U14505 ( .A(n12086), .ZN(n12087) );
  NAND3_X1 U14506 ( .A1(n12258), .A2(n15331), .A3(n12219), .ZN(n12091) );
  NAND3_X1 U14507 ( .A1(n12093), .A2(n12092), .A3(n12091), .ZN(n12098) );
  MUX2_X1 U14508 ( .A(n12095), .B(n12094), .S(n12227), .Z(n12096) );
  NAND2_X1 U14509 ( .A1(n12105), .A2(n12099), .ZN(n12102) );
  NAND2_X1 U14510 ( .A1(n12106), .A2(n12100), .ZN(n12101) );
  MUX2_X1 U14511 ( .A(n12102), .B(n12101), .S(n12227), .Z(n12103) );
  INV_X1 U14512 ( .A(n12103), .ZN(n12104) );
  MUX2_X1 U14513 ( .A(n12106), .B(n12105), .S(n12227), .Z(n12107) );
  NAND3_X1 U14514 ( .A1(n12109), .A2(n12108), .A3(n12107), .ZN(n12114) );
  MUX2_X1 U14515 ( .A(n12111), .B(n12110), .S(n12227), .Z(n12112) );
  NAND3_X1 U14516 ( .A1(n12114), .A2(n12113), .A3(n12112), .ZN(n12119) );
  MUX2_X1 U14517 ( .A(n12116), .B(n12115), .S(n12227), .Z(n12117) );
  NAND3_X1 U14518 ( .A1(n12119), .A2(n12118), .A3(n12117), .ZN(n12124) );
  MUX2_X1 U14519 ( .A(n15303), .B(n12120), .S(n12227), .Z(n12122) );
  NAND2_X1 U14520 ( .A1(n12122), .A2(n12121), .ZN(n12123) );
  NAND2_X1 U14521 ( .A1(n12124), .A2(n12123), .ZN(n12126) );
  NAND2_X1 U14522 ( .A1(n12126), .A2(n12125), .ZN(n12136) );
  NAND3_X1 U14523 ( .A1(n12136), .A2(n12135), .A3(n12127), .ZN(n12129) );
  NAND3_X1 U14524 ( .A1(n12129), .A2(n12128), .A3(n12130), .ZN(n12133) );
  MUX2_X1 U14525 ( .A(n12138), .B(n12130), .S(n12219), .Z(n12132) );
  AND2_X1 U14526 ( .A1(n12132), .A2(n12131), .ZN(n12141) );
  NAND2_X1 U14527 ( .A1(n12133), .A2(n12141), .ZN(n12144) );
  NAND3_X1 U14528 ( .A1(n12136), .A2(n12135), .A3(n12134), .ZN(n12139) );
  NAND3_X1 U14529 ( .A1(n12139), .A2(n12138), .A3(n12137), .ZN(n12142) );
  AOI21_X1 U14530 ( .B1(n12142), .B2(n12141), .A(n12140), .ZN(n12143) );
  MUX2_X1 U14531 ( .A(n12144), .B(n12143), .S(n12219), .Z(n12145) );
  MUX2_X1 U14532 ( .A(n12598), .B(n12147), .S(n12219), .Z(n12148) );
  INV_X1 U14533 ( .A(n12600), .ZN(n12603) );
  AOI21_X1 U14534 ( .B1(n12155), .B2(n12149), .A(n12227), .ZN(n12150) );
  OAI21_X1 U14535 ( .B1(n12151), .B2(n12150), .A(n12153), .ZN(n12158) );
  NAND2_X1 U14536 ( .A1(n12153), .A2(n12152), .ZN(n12154) );
  NAND2_X1 U14537 ( .A1(n12154), .A2(n12227), .ZN(n12157) );
  NOR2_X1 U14538 ( .A1(n12155), .A2(n12219), .ZN(n12156) );
  INV_X1 U14539 ( .A(n12159), .ZN(n12160) );
  NAND2_X1 U14540 ( .A1(n12167), .A2(n12160), .ZN(n12162) );
  AND3_X1 U14541 ( .A1(n12162), .A2(n12227), .A3(n12161), .ZN(n12163) );
  AND2_X1 U14542 ( .A1(n12163), .A2(n12172), .ZN(n12166) );
  OAI22_X1 U14543 ( .A1(n12165), .A2(n12569), .B1(n12166), .B2(n12164), .ZN(
        n12170) );
  INV_X1 U14544 ( .A(n12166), .ZN(n12169) );
  NAND3_X1 U14545 ( .A1(n12173), .A2(n12167), .A3(n12219), .ZN(n12168) );
  AOI22_X1 U14546 ( .A1(n12170), .A2(n12552), .B1(n12169), .B2(n12168), .ZN(
        n12180) );
  INV_X1 U14547 ( .A(n12171), .ZN(n12529) );
  MUX2_X1 U14548 ( .A(n12173), .B(n12172), .S(n12219), .Z(n12174) );
  NAND2_X1 U14549 ( .A1(n12529), .A2(n12174), .ZN(n12179) );
  MUX2_X1 U14550 ( .A(n12176), .B(n12175), .S(n12219), .Z(n12177) );
  OAI211_X1 U14551 ( .C1(n12180), .C2(n12179), .A(n12178), .B(n12177), .ZN(
        n12184) );
  MUX2_X1 U14552 ( .A(n12182), .B(n12181), .S(n12227), .Z(n12183) );
  NAND3_X1 U14553 ( .A1(n12184), .A2(n12497), .A3(n12183), .ZN(n12185) );
  NAND2_X1 U14554 ( .A1(n12185), .A2(n12480), .ZN(n12186) );
  INV_X1 U14555 ( .A(n12187), .ZN(n12189) );
  NAND2_X1 U14556 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  MUX2_X1 U14557 ( .A(n12191), .B(n12190), .S(n12227), .Z(n12192) );
  NAND3_X1 U14558 ( .A1(n12451), .A2(n12194), .A3(n12193), .ZN(n12195) );
  NAND3_X1 U14559 ( .A1(n12432), .A2(n12196), .A3(n12195), .ZN(n12200) );
  MUX2_X1 U14560 ( .A(n12198), .B(n12197), .S(n12227), .Z(n12199) );
  NAND2_X1 U14561 ( .A1(n12434), .A2(n12219), .ZN(n12201) );
  NOR2_X1 U14562 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  OR2_X1 U14563 ( .A1(n12205), .A2(n12204), .ZN(n12216) );
  INV_X1 U14564 ( .A(n12206), .ZN(n12215) );
  NAND2_X1 U14565 ( .A1(n12208), .A2(n12207), .ZN(n12210) );
  NAND2_X1 U14566 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  MUX2_X1 U14567 ( .A(n12212), .B(n12211), .S(n12227), .Z(n12213) );
  NAND2_X1 U14568 ( .A1(n6783), .A2(n12213), .ZN(n12214) );
  INV_X1 U14569 ( .A(n12218), .ZN(n12224) );
  NAND2_X1 U14570 ( .A1(n12220), .A2(n12219), .ZN(n12222) );
  NAND2_X1 U14571 ( .A1(n12222), .A2(n12221), .ZN(n12223) );
  OAI21_X1 U14572 ( .B1(n12225), .B2(n12224), .A(n12223), .ZN(n12231) );
  INV_X1 U14573 ( .A(n12225), .ZN(n12228) );
  NAND3_X1 U14574 ( .A1(n12228), .A2(n12227), .A3(n12226), .ZN(n12230) );
  NAND3_X1 U14575 ( .A1(n12231), .A2(n12230), .A3(n12229), .ZN(n12233) );
  NAND2_X1 U14576 ( .A1(n12233), .A2(n12232), .ZN(n12236) );
  NAND2_X1 U14577 ( .A1(n12236), .A2(n12234), .ZN(n12235) );
  AOI21_X1 U14578 ( .B1(n12240), .B2(n12239), .A(n12238), .ZN(n12247) );
  NAND2_X1 U14579 ( .A1(n12242), .A2(n12241), .ZN(n12243) );
  OAI211_X1 U14580 ( .C1(n12244), .C2(n12246), .A(n12243), .B(P3_B_REG_SCAN_IN), .ZN(n12245) );
  OAI21_X1 U14581 ( .B1(n12247), .B2(n12246), .A(n12245), .ZN(P3_U3296) );
  MUX2_X1 U14582 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12248), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14583 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12434), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14584 ( .A(n12448), .B(P3_DATAO_REG_26__SCAN_IN), .S(n12259), .Z(
        P3_U3517) );
  MUX2_X1 U14585 ( .A(n12249), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12259), .Z(
        P3_U3514) );
  MUX2_X1 U14586 ( .A(n12509), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12259), .Z(
        P3_U3513) );
  MUX2_X1 U14587 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12250), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14588 ( .A(n12536), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12259), .Z(
        P3_U3511) );
  MUX2_X1 U14589 ( .A(n12520), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12259), .Z(
        P3_U3510) );
  MUX2_X1 U14590 ( .A(n12580), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12259), .Z(
        P3_U3508) );
  MUX2_X1 U14591 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12251), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14592 ( .A(n12617), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12259), .Z(
        P3_U3506) );
  MUX2_X1 U14593 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12252), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14594 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n15304), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14595 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12253), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14596 ( .A(n15303), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12259), .Z(
        P3_U3500) );
  MUX2_X1 U14597 ( .A(n12254), .B(P3_DATAO_REG_8__SCAN_IN), .S(n12259), .Z(
        P3_U3499) );
  MUX2_X1 U14598 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12255), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14599 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12256), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14600 ( .A(n12257), .B(P3_DATAO_REG_5__SCAN_IN), .S(n12259), .Z(
        P3_U3496) );
  MUX2_X1 U14601 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n15320), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14602 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12258), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U14603 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n10825), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14604 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n10506), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14605 ( .A(n12696), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12259), .Z(
        P3_U3491) );
  NOR2_X1 U14606 ( .A1(n6802), .A2(n12260), .ZN(n12262) );
  NOR2_X2 U14607 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  XNOR2_X1 U14608 ( .A(n12293), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n12267) );
  NOR2_X2 U14609 ( .A1(n12263), .A2(n12267), .ZN(n12286) );
  AOI21_X1 U14610 ( .B1(n12263), .B2(n12267), .A(n12286), .ZN(n12284) );
  INV_X1 U14611 ( .A(n12264), .ZN(n12266) );
  AOI21_X1 U14612 ( .B1(n6802), .B2(n12266), .A(n12265), .ZN(n12271) );
  INV_X1 U14613 ( .A(n12267), .ZN(n12269) );
  NAND2_X1 U14614 ( .A1(n12293), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12294) );
  OR2_X1 U14615 ( .A1(n12293), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12268) );
  AND2_X1 U14616 ( .A1(n12294), .A2(n12268), .ZN(n12276) );
  MUX2_X1 U14617 ( .A(n12269), .B(n12276), .S(n12774), .Z(n12270) );
  NAND2_X1 U14618 ( .A1(n12271), .A2(n12270), .ZN(n12297) );
  OAI211_X1 U14619 ( .C1(n12271), .C2(n12270), .A(n12297), .B(n15285), .ZN(
        n12283) );
  NAND2_X1 U14620 ( .A1(n12273), .A2(n12272), .ZN(n12275) );
  NAND2_X1 U14621 ( .A1(n12275), .A2(n12274), .ZN(n12277) );
  NAND2_X1 U14622 ( .A1(n12276), .A2(n12277), .ZN(n12289) );
  OAI21_X1 U14623 ( .B1(n12277), .B2(n12276), .A(n12289), .ZN(n12281) );
  AOI21_X1 U14624 ( .B1(n15293), .B2(P3_ADDR_REG_14__SCAN_IN), .A(n12278), 
        .ZN(n12279) );
  OAI21_X1 U14625 ( .B1(n15290), .B2(n12293), .A(n12279), .ZN(n12280) );
  AOI21_X1 U14626 ( .B1(n12281), .B2(n15296), .A(n12280), .ZN(n12282) );
  OAI211_X1 U14627 ( .C1(n12284), .C2(n15300), .A(n12283), .B(n12282), .ZN(
        P3_U3196) );
  INV_X1 U14628 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12288) );
  AOI21_X1 U14629 ( .B1(n12288), .B2(n12287), .A(n12307), .ZN(n12305) );
  NAND2_X1 U14630 ( .A1(n12294), .A2(n12289), .ZN(n12310) );
  XNOR2_X1 U14631 ( .A(n12319), .B(n12310), .ZN(n12290) );
  NAND2_X1 U14632 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12290), .ZN(n12311) );
  OAI21_X1 U14633 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12290), .A(n12311), 
        .ZN(n12303) );
  AOI21_X1 U14634 ( .B1(n15293), .B2(P3_ADDR_REG_15__SCAN_IN), .A(n12291), 
        .ZN(n12292) );
  OAI21_X1 U14635 ( .B1(n15290), .B2(n14585), .A(n12292), .ZN(n12302) );
  NAND2_X1 U14636 ( .A1(n12293), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12295) );
  MUX2_X1 U14637 ( .A(n12295), .B(n12294), .S(n12774), .Z(n12296) );
  NAND2_X1 U14638 ( .A1(n12297), .A2(n12296), .ZN(n12317) );
  XNOR2_X1 U14639 ( .A(n12317), .B(n14585), .ZN(n12299) );
  MUX2_X1 U14640 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12774), .Z(n12298) );
  NOR2_X1 U14641 ( .A1(n12299), .A2(n12298), .ZN(n12318) );
  AOI21_X1 U14642 ( .B1(n12299), .B2(n12298), .A(n12318), .ZN(n12300) );
  NOR2_X1 U14643 ( .A1(n12300), .A2(n15176), .ZN(n12301) );
  AOI211_X1 U14644 ( .C1(n15296), .C2(n12303), .A(n12302), .B(n12301), .ZN(
        n12304) );
  OAI21_X1 U14645 ( .B1(n12305), .B2(n15300), .A(n12304), .ZN(P3_U3197) );
  NOR2_X1 U14646 ( .A1(n12319), .A2(n6595), .ZN(n12306) );
  INV_X1 U14647 ( .A(n12341), .ZN(n14590) );
  AOI22_X1 U14648 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n12341), .B1(n14590), 
        .B2(n12340), .ZN(n12308) );
  NOR2_X1 U14649 ( .A1(n12309), .A2(n12308), .ZN(n12343) );
  AOI21_X1 U14650 ( .B1(n12309), .B2(n12308), .A(n12343), .ZN(n12329) );
  INV_X1 U14651 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U14652 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n14590), .B1(n12341), 
        .B2(n12684), .ZN(n12314) );
  NAND2_X1 U14653 ( .A1(n14585), .A2(n12310), .ZN(n12312) );
  NAND2_X1 U14654 ( .A1(n12312), .A2(n12311), .ZN(n12313) );
  OAI21_X1 U14655 ( .B1(n12314), .B2(n12313), .A(n12330), .ZN(n12327) );
  INV_X1 U14656 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14558) );
  INV_X1 U14657 ( .A(n15293), .ZN(n15172) );
  NAND2_X1 U14658 ( .A1(n15181), .A2(n12341), .ZN(n12316) );
  OAI211_X1 U14659 ( .C1(n14558), .C2(n15172), .A(n12316), .B(n12315), .ZN(
        n12326) );
  INV_X1 U14660 ( .A(n12317), .ZN(n12320) );
  MUX2_X1 U14661 ( .A(n12340), .B(n12684), .S(n12774), .Z(n12321) );
  NOR2_X1 U14662 ( .A1(n12321), .A2(n12341), .ZN(n12334) );
  NAND2_X1 U14663 ( .A1(n12321), .A2(n12341), .ZN(n12333) );
  INV_X1 U14664 ( .A(n12333), .ZN(n12322) );
  NOR2_X1 U14665 ( .A1(n12334), .A2(n12322), .ZN(n12323) );
  XNOR2_X1 U14666 ( .A(n12335), .B(n12323), .ZN(n12324) );
  NOR2_X1 U14667 ( .A1(n12324), .A2(n15176), .ZN(n12325) );
  AOI211_X1 U14668 ( .C1(n15296), .C2(n12327), .A(n12326), .B(n12325), .ZN(
        n12328) );
  OAI21_X1 U14669 ( .B1(n12329), .B2(n15300), .A(n12328), .ZN(P3_U3198) );
  XNOR2_X1 U14670 ( .A(n12331), .B(n12351), .ZN(n12355) );
  XNOR2_X1 U14671 ( .A(n12355), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12349) );
  INV_X1 U14672 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14561) );
  OAI21_X1 U14673 ( .B1(n15172), .B2(n14561), .A(n12332), .ZN(n12339) );
  MUX2_X1 U14674 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12774), .Z(n12352) );
  XNOR2_X1 U14675 ( .A(n12352), .B(n12351), .ZN(n12337) );
  OAI21_X1 U14676 ( .B1(n12335), .B2(n12334), .A(n12333), .ZN(n12336) );
  NOR2_X1 U14677 ( .A1(n12336), .A2(n12337), .ZN(n12350) );
  AOI211_X1 U14678 ( .C1(n12337), .C2(n12336), .A(n15176), .B(n12350), .ZN(
        n12338) );
  AOI211_X1 U14679 ( .C1(n15181), .C2(n6694), .A(n12339), .B(n12338), .ZN(
        n12348) );
  NOR2_X1 U14680 ( .A1(n12341), .A2(n12340), .ZN(n12342) );
  NAND2_X1 U14681 ( .A1(n12344), .A2(n12351), .ZN(n12364) );
  OAI21_X1 U14682 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12345), .A(n12365), 
        .ZN(n12346) );
  NAND2_X1 U14683 ( .A1(n12346), .A2(n12366), .ZN(n12347) );
  OAI211_X1 U14684 ( .C1(n12349), .C2(n12387), .A(n12348), .B(n12347), .ZN(
        P3_U3199) );
  MUX2_X1 U14685 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12774), .Z(n12354) );
  NOR2_X2 U14686 ( .A1(n12353), .A2(n12354), .ZN(n12377) );
  AOI21_X1 U14687 ( .B1(n12354), .B2(n12353), .A(n12377), .ZN(n12370) );
  INV_X1 U14688 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13528) );
  OAI22_X1 U14689 ( .A1(n6694), .A2(n12356), .B1(n12355), .B2(n13528), .ZN(
        n12384) );
  XNOR2_X1 U14690 ( .A(n12378), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12383) );
  XNOR2_X1 U14691 ( .A(n12384), .B(n12383), .ZN(n12360) );
  NAND2_X1 U14692 ( .A1(n15293), .A2(P3_ADDR_REG_18__SCAN_IN), .ZN(n12357) );
  OAI211_X1 U14693 ( .C1(n15290), .C2(n12382), .A(n12358), .B(n12357), .ZN(
        n12359) );
  AOI21_X1 U14694 ( .B1(n12360), .B2(n15296), .A(n12359), .ZN(n12369) );
  OR2_X1 U14695 ( .A1(n12378), .A2(n12361), .ZN(n12371) );
  NAND2_X1 U14696 ( .A1(n12378), .A2(n12361), .ZN(n12362) );
  NAND2_X1 U14697 ( .A1(n12371), .A2(n12362), .ZN(n12363) );
  AND3_X1 U14698 ( .A1(n12365), .A2(n12364), .A3(n12363), .ZN(n12367) );
  OAI21_X1 U14699 ( .B1(n12373), .B2(n12367), .A(n12366), .ZN(n12368) );
  OAI211_X1 U14700 ( .C1(n12370), .C2(n15176), .A(n12369), .B(n12368), .ZN(
        P3_U3200) );
  INV_X1 U14701 ( .A(n12371), .ZN(n12372) );
  NOR2_X1 U14702 ( .A1(n12373), .A2(n12372), .ZN(n12374) );
  XNOR2_X1 U14703 ( .A(n12375), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12376) );
  XNOR2_X1 U14704 ( .A(n12374), .B(n12376), .ZN(n12396) );
  XNOR2_X1 U14705 ( .A(n12375), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12385) );
  MUX2_X1 U14706 ( .A(n12376), .B(n12385), .S(n12774), .Z(n12381) );
  AOI21_X1 U14707 ( .B1(n12379), .B2(n12378), .A(n12377), .ZN(n12380) );
  AOI22_X1 U14708 ( .A1(n12384), .A2(n12383), .B1(P3_REG1_REG_18__SCAN_IN), 
        .B2(n12382), .ZN(n12386) );
  XNOR2_X1 U14709 ( .A(n12386), .B(n12385), .ZN(n12388) );
  NOR2_X1 U14710 ( .A1(n12388), .A2(n12387), .ZN(n12393) );
  NAND2_X1 U14711 ( .A1(n15293), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12389) );
  OAI211_X1 U14712 ( .C1(n15290), .C2(n12391), .A(n12390), .B(n12389), .ZN(
        n12392) );
  AOI211_X1 U14713 ( .C1(n12394), .C2(n15285), .A(n12393), .B(n12392), .ZN(
        n12395) );
  OAI21_X1 U14714 ( .B1(n12396), .B2(n15300), .A(n12395), .ZN(P3_U3201) );
  INV_X1 U14715 ( .A(n12397), .ZN(n12403) );
  AOI22_X1 U14716 ( .A1(n14614), .A2(n15365), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n15371), .ZN(n12398) );
  OAI21_X1 U14717 ( .B1(n12399), .B2(n15312), .A(n12398), .ZN(n12400) );
  AOI21_X1 U14718 ( .B1(n12401), .B2(n12595), .A(n12400), .ZN(n12402) );
  OAI21_X1 U14719 ( .B1(n12403), .B2(n15371), .A(n12402), .ZN(P3_U3204) );
  INV_X1 U14720 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12404) );
  OAI22_X1 U14721 ( .A1(n12405), .A2(n15316), .B1(n15369), .B2(n12404), .ZN(
        n12406) );
  AOI21_X1 U14722 ( .B1(n12407), .B2(n14619), .A(n12406), .ZN(n12410) );
  NAND2_X1 U14723 ( .A1(n12408), .A2(n12595), .ZN(n12409) );
  OAI211_X1 U14724 ( .C1(n12411), .C2(n15371), .A(n12410), .B(n12409), .ZN(
        P3_U3205) );
  XOR2_X1 U14725 ( .A(n12413), .B(n12412), .Z(n12421) );
  OAI21_X1 U14726 ( .B1(n6796), .B2(n7062), .A(n12415), .ZN(n12419) );
  OAI22_X1 U14727 ( .A1(n12417), .A2(n15338), .B1(n12416), .B2(n15340), .ZN(
        n12418) );
  AOI21_X1 U14728 ( .B1(n12419), .B2(n15323), .A(n12418), .ZN(n12420) );
  OAI21_X1 U14729 ( .B1(n12421), .B2(n15328), .A(n12420), .ZN(n12629) );
  INV_X1 U14730 ( .A(n12629), .ZN(n12426) );
  INV_X1 U14731 ( .A(n12421), .ZN(n12630) );
  AOI22_X1 U14732 ( .A1(n12422), .A2(n15365), .B1(n15371), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12423) );
  OAI21_X1 U14733 ( .B1(n12711), .B2(n15312), .A(n12423), .ZN(n12424) );
  AOI21_X1 U14734 ( .B1(n12630), .B2(n15366), .A(n12424), .ZN(n12425) );
  OAI21_X1 U14735 ( .B1(n12426), .B2(n15371), .A(n12425), .ZN(P3_U3206) );
  NAND2_X1 U14736 ( .A1(n12508), .A2(n12427), .ZN(n12465) );
  NAND2_X1 U14737 ( .A1(n12465), .A2(n12428), .ZN(n12445) );
  NAND2_X1 U14738 ( .A1(n12445), .A2(n12429), .ZN(n12430) );
  XNOR2_X1 U14739 ( .A(n12430), .B(n12432), .ZN(n12431) );
  NAND2_X1 U14740 ( .A1(n12431), .A2(n15323), .ZN(n12437) );
  XNOR2_X1 U14741 ( .A(n12433), .B(n12432), .ZN(n12633) );
  NAND2_X1 U14742 ( .A1(n12633), .A2(n15352), .ZN(n12436) );
  AOI22_X1 U14743 ( .A1(n12434), .A2(n15319), .B1(n15321), .B2(n12470), .ZN(
        n12435) );
  NAND3_X1 U14744 ( .A1(n12437), .A2(n12436), .A3(n12435), .ZN(n12637) );
  INV_X1 U14745 ( .A(n12637), .ZN(n12443) );
  INV_X1 U14746 ( .A(n12438), .ZN(n12634) );
  AOI22_X1 U14747 ( .A1(n15371), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n12439), 
        .B2(n15365), .ZN(n12440) );
  OAI21_X1 U14748 ( .B1(n12634), .B2(n15312), .A(n12440), .ZN(n12441) );
  AOI21_X1 U14749 ( .B1(n12633), .B2(n15366), .A(n12441), .ZN(n12442) );
  OAI21_X1 U14750 ( .B1(n12443), .B2(n15371), .A(n12442), .ZN(P3_U3207) );
  AND2_X1 U14751 ( .A1(n12444), .A2(n12465), .ZN(n12447) );
  OAI211_X1 U14752 ( .C1(n12447), .C2(n12446), .A(n12445), .B(n15323), .ZN(
        n12450) );
  AOI22_X1 U14753 ( .A1(n12448), .A2(n15319), .B1(n15321), .B2(n12484), .ZN(
        n12449) );
  OR2_X1 U14754 ( .A1(n12452), .A2(n12451), .ZN(n12453) );
  NAND2_X1 U14755 ( .A1(n12454), .A2(n12453), .ZN(n12640) );
  INV_X1 U14756 ( .A(n12717), .ZN(n12457) );
  AOI22_X1 U14757 ( .A1(n15371), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n15365), 
        .B2(n12455), .ZN(n12456) );
  OAI21_X1 U14758 ( .B1(n12457), .B2(n15312), .A(n12456), .ZN(n12458) );
  AOI21_X1 U14759 ( .B1(n12640), .B2(n12595), .A(n12458), .ZN(n12459) );
  OAI21_X1 U14760 ( .B1(n12642), .B2(n15371), .A(n12459), .ZN(P3_U3208) );
  NAND2_X1 U14761 ( .A1(n12507), .A2(n12460), .ZN(n12462) );
  AND2_X1 U14762 ( .A1(n12462), .A2(n12461), .ZN(n12481) );
  AOI21_X1 U14763 ( .B1(n12474), .B2(n12467), .A(n7445), .ZN(n12472) );
  NOR2_X1 U14764 ( .A1(n12500), .A2(n15340), .ZN(n12469) );
  INV_X1 U14765 ( .A(n12647), .ZN(n12479) );
  OAI21_X1 U14766 ( .B1(n7419), .B2(n12474), .A(n12473), .ZN(n12645) );
  AOI22_X1 U14767 ( .A1(n15371), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15365), 
        .B2(n12475), .ZN(n12476) );
  OAI21_X1 U14768 ( .B1(n12721), .B2(n15312), .A(n12476), .ZN(n12477) );
  AOI21_X1 U14769 ( .B1(n12645), .B2(n12595), .A(n12477), .ZN(n12478) );
  OAI21_X1 U14770 ( .B1(n12479), .B2(n15371), .A(n12478), .ZN(P3_U3209) );
  NAND2_X1 U14771 ( .A1(n12481), .A2(n12480), .ZN(n12482) );
  NAND3_X1 U14772 ( .A1(n12483), .A2(n15323), .A3(n12482), .ZN(n12486) );
  AOI22_X1 U14773 ( .A1(n12484), .A2(n15319), .B1(n15321), .B2(n12509), .ZN(
        n12485) );
  AND2_X1 U14774 ( .A1(n12486), .A2(n12485), .ZN(n12652) );
  INV_X1 U14775 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12489) );
  INV_X1 U14776 ( .A(n12487), .ZN(n12488) );
  OAI22_X1 U14777 ( .A1(n15369), .A2(n12489), .B1(n12488), .B2(n15316), .ZN(
        n12490) );
  AOI21_X1 U14778 ( .B1(n12724), .B2(n14619), .A(n12490), .ZN(n12494) );
  XNOR2_X1 U14779 ( .A(n12492), .B(n12491), .ZN(n12650) );
  NAND2_X1 U14780 ( .A1(n12650), .A2(n12595), .ZN(n12493) );
  OAI211_X1 U14781 ( .C1(n12652), .C2(n15371), .A(n12494), .B(n12493), .ZN(
        P3_U3210) );
  XOR2_X1 U14782 ( .A(n12497), .B(n12495), .Z(n12656) );
  INV_X1 U14783 ( .A(n12656), .ZN(n12506) );
  NAND2_X1 U14784 ( .A1(n12507), .A2(n12496), .ZN(n12498) );
  XNOR2_X1 U14785 ( .A(n12498), .B(n12497), .ZN(n12499) );
  OAI222_X1 U14786 ( .A1(n15338), .A2(n12500), .B1(n15340), .B2(n12522), .C1(
        n15347), .C2(n12499), .ZN(n12655) );
  AOI22_X1 U14787 ( .A1(n15371), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15365), 
        .B2(n12502), .ZN(n12503) );
  OAI21_X1 U14788 ( .B1(n12729), .B2(n15312), .A(n12503), .ZN(n12504) );
  AOI21_X1 U14789 ( .B1(n12655), .B2(n15369), .A(n12504), .ZN(n12505) );
  OAI21_X1 U14790 ( .B1(n12506), .B2(n12625), .A(n12505), .ZN(P3_U3211) );
  OAI21_X1 U14791 ( .B1(n12508), .B2(n12516), .A(n12507), .ZN(n12510) );
  AOI222_X1 U14792 ( .A1(n15323), .A2(n12510), .B1(n12509), .B2(n15319), .C1(
        n12536), .C2(n15321), .ZN(n12659) );
  OAI22_X1 U14793 ( .A1(n15369), .A2(n12512), .B1(n12511), .B2(n15316), .ZN(
        n12513) );
  AOI21_X1 U14794 ( .B1(n12514), .B2(n14619), .A(n12513), .ZN(n12518) );
  XNOR2_X1 U14795 ( .A(n12515), .B(n12516), .ZN(n12661) );
  NAND2_X1 U14796 ( .A1(n12661), .A2(n12595), .ZN(n12517) );
  OAI211_X1 U14797 ( .C1(n12659), .C2(n15371), .A(n12518), .B(n12517), .ZN(
        P3_U3212) );
  XNOR2_X1 U14798 ( .A(n12519), .B(n12529), .ZN(n12524) );
  NAND2_X1 U14799 ( .A1(n12520), .A2(n15321), .ZN(n12521) );
  OAI21_X1 U14800 ( .B1(n12522), .B2(n15338), .A(n12521), .ZN(n12523) );
  AOI21_X1 U14801 ( .B1(n12524), .B2(n15323), .A(n12523), .ZN(n12666) );
  INV_X1 U14802 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12527) );
  INV_X1 U14803 ( .A(n12525), .ZN(n12526) );
  OAI22_X1 U14804 ( .A1(n15369), .A2(n12527), .B1(n12526), .B2(n15316), .ZN(
        n12528) );
  AOI21_X1 U14805 ( .B1(n12736), .B2(n14619), .A(n12528), .ZN(n12532) );
  XNOR2_X1 U14806 ( .A(n12530), .B(n12529), .ZN(n12664) );
  NAND2_X1 U14807 ( .A1(n12664), .A2(n12595), .ZN(n12531) );
  OAI211_X1 U14808 ( .C1(n12666), .C2(n15371), .A(n12532), .B(n12531), .ZN(
        P3_U3213) );
  NAND2_X1 U14809 ( .A1(n12533), .A2(n12540), .ZN(n12534) );
  NAND3_X1 U14810 ( .A1(n12535), .A2(n15323), .A3(n12534), .ZN(n12539) );
  AOI22_X1 U14811 ( .A1(n12537), .A2(n15321), .B1(n15319), .B2(n12536), .ZN(
        n12538) );
  AND2_X1 U14812 ( .A1(n12539), .A2(n12538), .ZN(n12670) );
  XNOR2_X1 U14813 ( .A(n12541), .B(n7961), .ZN(n12669) );
  NAND2_X1 U14814 ( .A1(n12669), .A2(n12595), .ZN(n12547) );
  INV_X1 U14815 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12544) );
  INV_X1 U14816 ( .A(n12542), .ZN(n12543) );
  OAI22_X1 U14817 ( .A1(n15369), .A2(n12544), .B1(n12543), .B2(n15316), .ZN(
        n12545) );
  AOI21_X1 U14818 ( .B1(n12740), .B2(n14619), .A(n12545), .ZN(n12546) );
  OAI211_X1 U14819 ( .C1(n12670), .C2(n15371), .A(n12547), .B(n12546), .ZN(
        P3_U3214) );
  XNOR2_X1 U14820 ( .A(n12548), .B(n12552), .ZN(n12675) );
  INV_X1 U14821 ( .A(n12675), .ZN(n12560) );
  INV_X1 U14822 ( .A(n12549), .ZN(n12550) );
  AOI21_X1 U14823 ( .B1(n12552), .B2(n12551), .A(n12550), .ZN(n12553) );
  OAI222_X1 U14824 ( .A1(n15338), .A2(n12555), .B1(n15340), .B2(n12554), .C1(
        n15347), .C2(n12553), .ZN(n12674) );
  AOI22_X1 U14825 ( .A1(n15371), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n15365), 
        .B2(n12556), .ZN(n12557) );
  OAI21_X1 U14826 ( .B1(n12745), .B2(n15312), .A(n12557), .ZN(n12558) );
  AOI21_X1 U14827 ( .B1(n12674), .B2(n15369), .A(n12558), .ZN(n12559) );
  OAI21_X1 U14828 ( .B1(n12625), .B2(n12560), .A(n12559), .ZN(P3_U3215) );
  NAND2_X1 U14829 ( .A1(n12562), .A2(n12561), .ZN(n12564) );
  NAND2_X1 U14830 ( .A1(n12584), .A2(n12566), .ZN(n12568) );
  XNOR2_X1 U14831 ( .A(n12568), .B(n12567), .ZN(n12679) );
  INV_X1 U14832 ( .A(n12679), .ZN(n12577) );
  XNOR2_X1 U14833 ( .A(n12570), .B(n12569), .ZN(n12571) );
  OAI222_X1 U14834 ( .A1(n15338), .A2(n12572), .B1(n15340), .B2(n12607), .C1(
        n12571), .C2(n15347), .ZN(n12678) );
  AOI22_X1 U14835 ( .A1(n15371), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n15365), 
        .B2(n12573), .ZN(n12574) );
  OAI21_X1 U14836 ( .B1(n12749), .B2(n15312), .A(n12574), .ZN(n12575) );
  AOI21_X1 U14837 ( .B1(n12678), .B2(n15369), .A(n12575), .ZN(n12576) );
  OAI21_X1 U14838 ( .B1(n12625), .B2(n12577), .A(n12576), .ZN(P3_U3216) );
  XNOR2_X1 U14839 ( .A(n12578), .B(n12588), .ZN(n12579) );
  NAND2_X1 U14840 ( .A1(n12579), .A2(n15323), .ZN(n12582) );
  AOI22_X1 U14841 ( .A1(n15321), .A2(n12617), .B1(n12580), .B2(n15319), .ZN(
        n12581) );
  AND2_X1 U14842 ( .A1(n12584), .A2(n12583), .ZN(n12591) );
  OR2_X1 U14843 ( .A1(n12614), .A2(n12585), .ZN(n12587) );
  NAND2_X1 U14844 ( .A1(n12587), .A2(n12586), .ZN(n12589) );
  OR2_X1 U14845 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  NAND2_X1 U14846 ( .A1(n12591), .A2(n12590), .ZN(n12681) );
  AOI22_X1 U14847 ( .A1(n15371), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15365), 
        .B2(n12592), .ZN(n12593) );
  OAI21_X1 U14848 ( .B1(n12753), .B2(n15312), .A(n12593), .ZN(n12594) );
  AOI21_X1 U14849 ( .B1(n12681), .B2(n12595), .A(n12594), .ZN(n12596) );
  OAI21_X1 U14850 ( .B1(n12683), .B2(n15371), .A(n12596), .ZN(P3_U3217) );
  OR2_X1 U14851 ( .A1(n12614), .A2(n12597), .ZN(n12599) );
  NAND2_X1 U14852 ( .A1(n12599), .A2(n12598), .ZN(n12601) );
  XNOR2_X1 U14853 ( .A(n12601), .B(n12600), .ZN(n12687) );
  INV_X1 U14854 ( .A(n12687), .ZN(n12613) );
  NAND2_X1 U14855 ( .A1(n12616), .A2(n12602), .ZN(n12604) );
  XNOR2_X1 U14856 ( .A(n12604), .B(n12603), .ZN(n12605) );
  OAI222_X1 U14857 ( .A1(n15338), .A2(n12607), .B1(n15340), .B2(n12606), .C1(
        n12605), .C2(n15347), .ZN(n12686) );
  INV_X1 U14858 ( .A(n12608), .ZN(n12757) );
  AOI22_X1 U14859 ( .A1(n15371), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n15365), 
        .B2(n12609), .ZN(n12610) );
  OAI21_X1 U14860 ( .B1(n12757), .B2(n15312), .A(n12610), .ZN(n12611) );
  AOI21_X1 U14861 ( .B1(n12686), .B2(n15369), .A(n12611), .ZN(n12612) );
  OAI21_X1 U14862 ( .B1(n12625), .B2(n12613), .A(n12612), .ZN(P3_U3218) );
  XOR2_X1 U14863 ( .A(n12615), .B(n12614), .Z(n12691) );
  INV_X1 U14864 ( .A(n12691), .ZN(n12626) );
  OAI211_X1 U14865 ( .C1(n7439), .C2(n7948), .A(n15323), .B(n12616), .ZN(
        n12620) );
  AOI22_X1 U14866 ( .A1(n15321), .A2(n12618), .B1(n12617), .B2(n15319), .ZN(
        n12619) );
  NAND2_X1 U14867 ( .A1(n12620), .A2(n12619), .ZN(n12690) );
  AOI22_X1 U14868 ( .A1(n15371), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15365), 
        .B2(n12621), .ZN(n12622) );
  OAI21_X1 U14869 ( .B1(n12761), .B2(n15312), .A(n12622), .ZN(n12623) );
  AOI21_X1 U14870 ( .B1(n12690), .B2(n15369), .A(n12623), .ZN(n12624) );
  OAI21_X1 U14871 ( .B1(n12626), .B2(n12625), .A(n12624), .ZN(P3_U3219) );
  INV_X1 U14872 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12631) );
  AOI21_X1 U14873 ( .B1(n15400), .B2(n12630), .A(n12629), .ZN(n12709) );
  MUX2_X1 U14874 ( .A(n12631), .B(n12709), .S(n15424), .Z(n12632) );
  OAI21_X1 U14875 ( .B1(n12711), .B2(n12694), .A(n12632), .ZN(P3_U3486) );
  INV_X1 U14876 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12638) );
  INV_X1 U14877 ( .A(n12633), .ZN(n12635) );
  INV_X1 U14878 ( .A(n15400), .ZN(n15407) );
  OAI22_X1 U14879 ( .A1(n12635), .A2(n15407), .B1(n12634), .B2(n15406), .ZN(
        n12636) );
  NOR2_X1 U14880 ( .A1(n12637), .A2(n12636), .ZN(n12712) );
  MUX2_X1 U14881 ( .A(n12638), .B(n12712), .S(n15424), .Z(n12639) );
  INV_X1 U14882 ( .A(n12639), .ZN(P3_U3485) );
  NAND2_X1 U14883 ( .A1(n12640), .A2(n14640), .ZN(n12641) );
  NAND2_X1 U14884 ( .A1(n12642), .A2(n12641), .ZN(n12715) );
  MUX2_X1 U14885 ( .A(n12715), .B(P3_REG1_REG_25__SCAN_IN), .S(n8836), .Z(
        n12643) );
  AOI21_X1 U14886 ( .B1(n8838), .B2(n12717), .A(n12643), .ZN(n12644) );
  INV_X1 U14887 ( .A(n12644), .ZN(P3_U3484) );
  MUX2_X1 U14888 ( .A(n12648), .B(n12719), .S(n15424), .Z(n12649) );
  OAI21_X1 U14889 ( .B1(n12721), .B2(n12694), .A(n12649), .ZN(P3_U3483) );
  NAND2_X1 U14890 ( .A1(n12650), .A2(n14640), .ZN(n12651) );
  NAND2_X1 U14891 ( .A1(n12652), .A2(n12651), .ZN(n12722) );
  MUX2_X1 U14892 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n12722), .S(n15424), .Z(
        n12653) );
  AOI21_X1 U14893 ( .B1(n8838), .B2(n12724), .A(n12653), .ZN(n12654) );
  INV_X1 U14894 ( .A(n12654), .ZN(P3_U3482) );
  INV_X1 U14895 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12657) );
  AOI21_X1 U14896 ( .B1(n14640), .B2(n12656), .A(n12655), .ZN(n12726) );
  MUX2_X1 U14897 ( .A(n12657), .B(n12726), .S(n15424), .Z(n12658) );
  OAI21_X1 U14898 ( .B1(n12729), .B2(n12694), .A(n12658), .ZN(P3_U3481) );
  INV_X1 U14899 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12662) );
  INV_X1 U14900 ( .A(n12659), .ZN(n12660) );
  AOI21_X1 U14901 ( .B1(n14640), .B2(n12661), .A(n12660), .ZN(n12730) );
  MUX2_X1 U14902 ( .A(n12662), .B(n12730), .S(n15424), .Z(n12663) );
  OAI21_X1 U14903 ( .B1(n12733), .B2(n12694), .A(n12663), .ZN(P3_U3480) );
  NAND2_X1 U14904 ( .A1(n12664), .A2(n14640), .ZN(n12665) );
  NAND2_X1 U14905 ( .A1(n12666), .A2(n12665), .ZN(n12734) );
  MUX2_X1 U14906 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12734), .S(n15424), .Z(
        n12667) );
  AOI21_X1 U14907 ( .B1(n8838), .B2(n12736), .A(n12667), .ZN(n12668) );
  INV_X1 U14908 ( .A(n12668), .ZN(P3_U3479) );
  NAND2_X1 U14909 ( .A1(n12669), .A2(n14640), .ZN(n12671) );
  NAND2_X1 U14910 ( .A1(n12671), .A2(n12670), .ZN(n12738) );
  MUX2_X1 U14911 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12738), .S(n15424), .Z(
        n12672) );
  AOI21_X1 U14912 ( .B1(n8838), .B2(n12740), .A(n12672), .ZN(n12673) );
  INV_X1 U14913 ( .A(n12673), .ZN(P3_U3478) );
  INV_X1 U14914 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12676) );
  AOI21_X1 U14915 ( .B1(n12675), .B2(n14640), .A(n12674), .ZN(n12742) );
  MUX2_X1 U14916 ( .A(n12676), .B(n12742), .S(n15424), .Z(n12677) );
  OAI21_X1 U14917 ( .B1(n12745), .B2(n12694), .A(n12677), .ZN(P3_U3477) );
  AOI21_X1 U14918 ( .B1(n12679), .B2(n14640), .A(n12678), .ZN(n12746) );
  MUX2_X1 U14919 ( .A(n13528), .B(n12746), .S(n15424), .Z(n12680) );
  OAI21_X1 U14920 ( .B1(n12749), .B2(n12694), .A(n12680), .ZN(P3_U3476) );
  NAND2_X1 U14921 ( .A1(n12681), .A2(n14640), .ZN(n12682) );
  AND2_X1 U14922 ( .A1(n12683), .A2(n12682), .ZN(n12751) );
  MUX2_X1 U14923 ( .A(n12684), .B(n12751), .S(n15424), .Z(n12685) );
  OAI21_X1 U14924 ( .B1(n12753), .B2(n12694), .A(n12685), .ZN(P3_U3475) );
  INV_X1 U14925 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12688) );
  AOI21_X1 U14926 ( .B1(n12687), .B2(n14640), .A(n12686), .ZN(n12754) );
  MUX2_X1 U14927 ( .A(n12688), .B(n12754), .S(n15424), .Z(n12689) );
  OAI21_X1 U14928 ( .B1(n12757), .B2(n12694), .A(n12689), .ZN(P3_U3474) );
  INV_X1 U14929 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12692) );
  AOI21_X1 U14930 ( .B1(n12691), .B2(n14640), .A(n12690), .ZN(n12758) );
  MUX2_X1 U14931 ( .A(n12692), .B(n12758), .S(n15424), .Z(n12693) );
  OAI21_X1 U14932 ( .B1(n12694), .B2(n12761), .A(n12693), .ZN(P3_U3473) );
  OAI21_X1 U14933 ( .B1(n12695), .B2(n12702), .A(n15346), .ZN(n12700) );
  NAND2_X1 U14934 ( .A1(n12696), .A2(n15321), .ZN(n12697) );
  OAI21_X1 U14935 ( .B1(n12698), .B2(n15338), .A(n12697), .ZN(n12699) );
  AOI21_X1 U14936 ( .B1(n12700), .B2(n15323), .A(n12699), .ZN(n12704) );
  XNOR2_X1 U14937 ( .A(n12702), .B(n12701), .ZN(n12705) );
  OR2_X1 U14938 ( .A1(n12705), .A2(n15328), .ZN(n12703) );
  INV_X1 U14939 ( .A(n12705), .ZN(n15367) );
  AND2_X1 U14940 ( .A1(n12706), .A2(n14625), .ZN(n15364) );
  AOI21_X1 U14941 ( .B1(n15367), .B2(n15400), .A(n15364), .ZN(n12707) );
  AND2_X1 U14942 ( .A1(n15361), .A2(n12707), .ZN(n15372) );
  INV_X1 U14943 ( .A(n15372), .ZN(n12708) );
  MUX2_X1 U14944 ( .A(n12708), .B(P3_REG1_REG_1__SCAN_IN), .S(n8836), .Z(
        P3_U3460) );
  INV_X1 U14945 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13600) );
  MUX2_X1 U14946 ( .A(n13600), .B(n12709), .S(n15411), .Z(n12710) );
  OAI21_X1 U14947 ( .B1(n12711), .B2(n12762), .A(n12710), .ZN(P3_U3454) );
  MUX2_X1 U14948 ( .A(n12713), .B(n12712), .S(n15411), .Z(n12714) );
  INV_X1 U14949 ( .A(n12714), .ZN(P3_U3453) );
  MUX2_X1 U14950 ( .A(n12715), .B(P3_REG0_REG_25__SCAN_IN), .S(n15412), .Z(
        n12716) );
  AOI21_X1 U14951 ( .B1(n8823), .B2(n12717), .A(n12716), .ZN(n12718) );
  INV_X1 U14952 ( .A(n12718), .ZN(P3_U3452) );
  INV_X1 U14953 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13491) );
  MUX2_X1 U14954 ( .A(n13491), .B(n12719), .S(n15411), .Z(n12720) );
  OAI21_X1 U14955 ( .B1(n12721), .B2(n12762), .A(n12720), .ZN(P3_U3451) );
  MUX2_X1 U14956 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n12722), .S(n15411), .Z(
        n12723) );
  AOI21_X1 U14957 ( .B1(n8823), .B2(n12724), .A(n12723), .ZN(n12725) );
  INV_X1 U14958 ( .A(n12725), .ZN(P3_U3450) );
  INV_X1 U14959 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12727) );
  MUX2_X1 U14960 ( .A(n12727), .B(n12726), .S(n15411), .Z(n12728) );
  OAI21_X1 U14961 ( .B1(n12729), .B2(n12762), .A(n12728), .ZN(P3_U3449) );
  MUX2_X1 U14962 ( .A(n12731), .B(n12730), .S(n15411), .Z(n12732) );
  OAI21_X1 U14963 ( .B1(n12733), .B2(n12762), .A(n12732), .ZN(P3_U3448) );
  MUX2_X1 U14964 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12734), .S(n15411), .Z(
        n12735) );
  AOI21_X1 U14965 ( .B1(n8823), .B2(n12736), .A(n12735), .ZN(n12737) );
  INV_X1 U14966 ( .A(n12737), .ZN(P3_U3447) );
  MUX2_X1 U14967 ( .A(n12738), .B(P3_REG0_REG_19__SCAN_IN), .S(n15412), .Z(
        n12739) );
  AOI21_X1 U14968 ( .B1(n8823), .B2(n12740), .A(n12739), .ZN(n12741) );
  INV_X1 U14969 ( .A(n12741), .ZN(P3_U3446) );
  MUX2_X1 U14970 ( .A(n12743), .B(n12742), .S(n15411), .Z(n12744) );
  OAI21_X1 U14971 ( .B1(n12745), .B2(n12762), .A(n12744), .ZN(P3_U3444) );
  INV_X1 U14972 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12747) );
  MUX2_X1 U14973 ( .A(n12747), .B(n12746), .S(n15411), .Z(n12748) );
  OAI21_X1 U14974 ( .B1(n12749), .B2(n12762), .A(n12748), .ZN(P3_U3441) );
  MUX2_X1 U14975 ( .A(n12751), .B(n12750), .S(n15412), .Z(n12752) );
  OAI21_X1 U14976 ( .B1(n12753), .B2(n12762), .A(n12752), .ZN(P3_U3438) );
  INV_X1 U14977 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12755) );
  MUX2_X1 U14978 ( .A(n12755), .B(n12754), .S(n15411), .Z(n12756) );
  OAI21_X1 U14979 ( .B1(n12757), .B2(n12762), .A(n12756), .ZN(P3_U3435) );
  MUX2_X1 U14980 ( .A(n12759), .B(n12758), .S(n15411), .Z(n12760) );
  OAI21_X1 U14981 ( .B1(n12762), .B2(n12761), .A(n12760), .ZN(P3_U3432) );
  NAND2_X1 U14982 ( .A1(n12763), .A2(n14587), .ZN(n12766) );
  OR4_X1 U14983 ( .A1(n12764), .A2(P3_IR_REG_30__SCAN_IN), .A3(n8002), .A4(
        P3_U3151), .ZN(n12765) );
  OAI211_X1 U14984 ( .C1(n12767), .C2(n14574), .A(n12766), .B(n12765), .ZN(
        P3_U3264) );
  OAI222_X1 U14985 ( .A1(P3_U3151), .A2(n12769), .B1(n14576), .B2(n12768), 
        .C1(n13654), .C2(n14574), .ZN(P3_U3265) );
  INV_X1 U14986 ( .A(n12770), .ZN(n12772) );
  OAI222_X1 U14987 ( .A1(n14574), .A2(n13569), .B1(n14576), .B2(n12772), .C1(
        P3_U3151), .C2(n12771), .ZN(P3_U3266) );
  INV_X1 U14988 ( .A(n12773), .ZN(n12776) );
  OAI222_X1 U14989 ( .A1(n14576), .A2(n12776), .B1(n14574), .B2(n12775), .C1(
        P3_U3151), .C2(n12774), .ZN(P3_U3268) );
  INV_X1 U14990 ( .A(n12777), .ZN(n12778) );
  OAI222_X1 U14991 ( .A1(n12780), .A2(P3_U3151), .B1(n14576), .B2(n12778), 
        .C1(n13476), .C2(n14574), .ZN(P3_U3269) );
  INV_X1 U14992 ( .A(n13280), .ZN(n12793) );
  NAND2_X1 U14993 ( .A1(n12783), .A2(n12782), .ZN(n12784) );
  NAND3_X1 U14994 ( .A1(n12785), .A2(n12946), .A3(n12784), .ZN(n12792) );
  NAND2_X1 U14995 ( .A1(n12961), .A2(n12933), .ZN(n12787) );
  NAND2_X1 U14996 ( .A1(n12963), .A2(n12932), .ZN(n12786) );
  NAND2_X1 U14997 ( .A1(n12787), .A2(n12786), .ZN(n13082) );
  INV_X1 U14998 ( .A(n13086), .ZN(n12789) );
  OAI22_X1 U14999 ( .A1(n12789), .A2(n12953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12788), .ZN(n12790) );
  AOI21_X1 U15000 ( .B1(n13082), .B2(n12950), .A(n12790), .ZN(n12791) );
  OAI211_X1 U15001 ( .C1(n12793), .C2(n12926), .A(n12792), .B(n12791), .ZN(
        P2_U3186) );
  NAND3_X1 U15002 ( .A1(n12795), .A2(n12945), .A3(n12975), .ZN(n12796) );
  OAI21_X1 U15003 ( .B1(n12794), .B2(n12938), .A(n12796), .ZN(n12799) );
  INV_X1 U15004 ( .A(n12797), .ZN(n12798) );
  NAND2_X1 U15005 ( .A1(n12799), .A2(n12798), .ZN(n12806) );
  NOR2_X1 U15006 ( .A1(n12953), .A2(n12800), .ZN(n12804) );
  OAI22_X1 U15007 ( .A1(n12937), .A2(n12802), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12801), .ZN(n12803) );
  AOI211_X1 U15008 ( .C1(n13344), .C2(n8784), .A(n12804), .B(n12803), .ZN(
        n12805) );
  OAI211_X1 U15009 ( .C1(n12807), .C2(n12938), .A(n12806), .B(n12805), .ZN(
        P2_U3187) );
  INV_X1 U15010 ( .A(n13302), .ZN(n12822) );
  INV_X1 U15011 ( .A(n12808), .ZN(n12810) );
  NOR2_X1 U15012 ( .A1(n12810), .A2(n12809), .ZN(n12919) );
  NOR2_X1 U15013 ( .A1(n12919), .A2(n12811), .ZN(n12813) );
  XNOR2_X1 U15014 ( .A(n12813), .B(n12812), .ZN(n12816) );
  OAI22_X1 U15015 ( .A1(n12816), .A2(n12938), .B1(n12885), .B2(n12927), .ZN(
        n12814) );
  OAI21_X1 U15016 ( .B1(n12816), .B2(n12815), .A(n12814), .ZN(n12821) );
  OAI22_X1 U15017 ( .A1(n12852), .A2(n12886), .B1(n12817), .B2(n12884), .ZN(
        n13143) );
  OAI22_X1 U15018 ( .A1(n13149), .A2(n12953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12818), .ZN(n12819) );
  AOI21_X1 U15019 ( .B1(n13143), .B2(n12950), .A(n12819), .ZN(n12820) );
  OAI211_X1 U15020 ( .C1(n12822), .C2(n12926), .A(n12821), .B(n12820), .ZN(
        P2_U3188) );
  NAND3_X1 U15021 ( .A1(n12825), .A2(n12945), .A3(n12970), .ZN(n12826) );
  OAI21_X1 U15022 ( .B1(n12824), .B2(n12938), .A(n12826), .ZN(n12829) );
  INV_X1 U15023 ( .A(n12827), .ZN(n12828) );
  NAND2_X1 U15024 ( .A1(n12829), .A2(n12828), .ZN(n12834) );
  NOR2_X1 U15025 ( .A1(n12953), .A2(n13208), .ZN(n12832) );
  AND2_X1 U15026 ( .A1(n12970), .A2(n12932), .ZN(n12830) );
  AOI21_X1 U15027 ( .B1(n12968), .B2(n12933), .A(n12830), .ZN(n13206) );
  NAND2_X1 U15028 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13050)
         );
  OAI21_X1 U15029 ( .B1(n13206), .B2(n12937), .A(n13050), .ZN(n12831) );
  AOI211_X1 U15030 ( .C1(n13323), .C2(n8784), .A(n12832), .B(n12831), .ZN(
        n12833) );
  OAI211_X1 U15031 ( .C1(n12938), .C2(n12823), .A(n12834), .B(n12833), .ZN(
        P2_U3191) );
  AOI21_X1 U15032 ( .B1(n12836), .B2(n12835), .A(n12938), .ZN(n12838) );
  NAND2_X1 U15033 ( .A1(n12838), .A2(n12837), .ZN(n12844) );
  NAND2_X1 U15034 ( .A1(n12966), .A2(n12933), .ZN(n12840) );
  NAND2_X1 U15035 ( .A1(n12968), .A2(n12932), .ZN(n12839) );
  NAND2_X1 U15036 ( .A1(n12840), .A2(n12839), .ZN(n13180) );
  OAI22_X1 U15037 ( .A1(n12953), .A2(n13174), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12841), .ZN(n12842) );
  AOI21_X1 U15038 ( .B1(n13180), .B2(n12950), .A(n12842), .ZN(n12843) );
  OAI211_X1 U15039 ( .C1(n13177), .C2(n12926), .A(n12844), .B(n12843), .ZN(
        P2_U3195) );
  INV_X1 U15040 ( .A(n13292), .ZN(n12858) );
  INV_X1 U15041 ( .A(n12846), .ZN(n12847) );
  AOI21_X1 U15042 ( .B1(n12845), .B2(n12847), .A(n12938), .ZN(n12851) );
  NOR3_X1 U15043 ( .A1(n12848), .A2(n12852), .A3(n12927), .ZN(n12850) );
  OAI21_X1 U15044 ( .B1(n12851), .B2(n12850), .A(n12849), .ZN(n12857) );
  OAI22_X1 U15045 ( .A1(n12853), .A2(n12886), .B1(n12852), .B2(n12884), .ZN(
        n13119) );
  OAI22_X1 U15046 ( .A1(n13115), .A2(n12953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12854), .ZN(n12855) );
  AOI21_X1 U15047 ( .B1(n13119), .B2(n12950), .A(n12855), .ZN(n12856) );
  OAI211_X1 U15048 ( .C1(n12858), .C2(n12926), .A(n12857), .B(n12856), .ZN(
        P2_U3197) );
  INV_X1 U15049 ( .A(n12878), .ZN(n12859) );
  AOI21_X1 U15050 ( .B1(n12861), .B2(n12860), .A(n12859), .ZN(n12868) );
  OAI22_X1 U15051 ( .A1(n12863), .A2(n12937), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12862), .ZN(n12864) );
  AOI21_X1 U15052 ( .B1(n12865), .B2(n12935), .A(n12864), .ZN(n12867) );
  NAND2_X1 U15053 ( .A1(n13339), .A2(n8784), .ZN(n12866) );
  OAI211_X1 U15054 ( .C1(n12868), .C2(n12938), .A(n12867), .B(n12866), .ZN(
        P2_U3198) );
  NAND2_X1 U15055 ( .A1(n12970), .A2(n12933), .ZN(n12870) );
  NAND2_X1 U15056 ( .A1(n12972), .A2(n12932), .ZN(n12869) );
  NAND2_X1 U15057 ( .A1(n12870), .A2(n12869), .ZN(n13240) );
  AOI22_X1 U15058 ( .A1(n13240), .A2(n12950), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12871) );
  OAI21_X1 U15059 ( .B1(n13233), .B2(n12953), .A(n12871), .ZN(n12872) );
  AOI21_X1 U15060 ( .B1(n13333), .B2(n8784), .A(n12872), .ZN(n12880) );
  INV_X1 U15061 ( .A(n12873), .ZN(n12877) );
  OAI22_X1 U15062 ( .A1(n12875), .A2(n12938), .B1(n12874), .B2(n12927), .ZN(
        n12876) );
  NAND3_X1 U15063 ( .A1(n12878), .A2(n12877), .A3(n12876), .ZN(n12879) );
  OAI211_X1 U15064 ( .C1(n12881), .C2(n12938), .A(n12880), .B(n12879), .ZN(
        P2_U3200) );
  INV_X1 U15065 ( .A(n13297), .ZN(n13138) );
  OAI211_X1 U15066 ( .C1(n12883), .C2(n12882), .A(n12845), .B(n12946), .ZN(
        n12890) );
  OAI22_X1 U15067 ( .A1(n12928), .A2(n12886), .B1(n12885), .B2(n12884), .ZN(
        n13127) );
  INV_X1 U15068 ( .A(n13135), .ZN(n12887) );
  OAI22_X1 U15069 ( .A1(n12887), .A2(n12953), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13650), .ZN(n12888) );
  AOI21_X1 U15070 ( .B1(n13127), .B2(n12950), .A(n12888), .ZN(n12889) );
  OAI211_X1 U15071 ( .C1(n13138), .C2(n12926), .A(n12890), .B(n12889), .ZN(
        P2_U3201) );
  AND2_X1 U15072 ( .A1(n12969), .A2(n12932), .ZN(n12891) );
  AOI21_X1 U15073 ( .B1(n12967), .B2(n12933), .A(n12891), .ZN(n13190) );
  OAI22_X1 U15074 ( .A1(n13190), .A2(n12937), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12892), .ZN(n12894) );
  INV_X1 U15075 ( .A(n13318), .ZN(n13196) );
  NOR2_X1 U15076 ( .A1(n13196), .A2(n12926), .ZN(n12893) );
  AOI211_X1 U15077 ( .C1(n12935), .C2(n13193), .A(n12894), .B(n12893), .ZN(
        n12901) );
  INV_X1 U15078 ( .A(n12895), .ZN(n12899) );
  OAI22_X1 U15079 ( .A1(n12897), .A2(n12938), .B1(n12896), .B2(n12927), .ZN(
        n12898) );
  NAND3_X1 U15080 ( .A1(n12823), .A2(n12899), .A3(n12898), .ZN(n12900) );
  OAI211_X1 U15081 ( .C1(n12902), .C2(n12938), .A(n12901), .B(n12900), .ZN(
        P2_U3205) );
  AOI22_X1 U15082 ( .A1(n12950), .A2(n12903), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12904) );
  OAI21_X1 U15083 ( .B1(n12953), .B2(n12905), .A(n12904), .ZN(n12910) );
  INV_X1 U15084 ( .A(n12794), .ZN(n12906) );
  AOI211_X1 U15085 ( .C1(n12908), .C2(n12907), .A(n12938), .B(n12906), .ZN(
        n12909) );
  AOI211_X1 U15086 ( .C1(n14650), .C2(n8784), .A(n12910), .B(n12909), .ZN(
        n12911) );
  INV_X1 U15087 ( .A(n12911), .ZN(P2_U3206) );
  AOI22_X1 U15088 ( .A1(n12808), .A2(n12946), .B1(n12945), .B2(n12966), .ZN(
        n12918) );
  AND2_X1 U15089 ( .A1(n12967), .A2(n12932), .ZN(n12912) );
  AOI21_X1 U15090 ( .B1(n12913), .B2(n12933), .A(n12912), .ZN(n13163) );
  INV_X1 U15091 ( .A(n12914), .ZN(n13158) );
  AOI22_X1 U15092 ( .A1(n13158), .A2(n12935), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12915) );
  OAI21_X1 U15093 ( .B1(n13163), .B2(n12937), .A(n12915), .ZN(n12916) );
  AOI21_X1 U15094 ( .B1(n13307), .B2(n8784), .A(n12916), .ZN(n12917) );
  OAI21_X1 U15095 ( .B1(n12919), .B2(n12918), .A(n12917), .ZN(P2_U3207) );
  INV_X1 U15096 ( .A(n13328), .ZN(n13225) );
  AOI21_X1 U15097 ( .B1(n12921), .B2(n12920), .A(n12938), .ZN(n12922) );
  NAND2_X1 U15098 ( .A1(n12922), .A2(n12824), .ZN(n12925) );
  AOI22_X1 U15099 ( .A1(n12969), .A2(n12933), .B1(n12932), .B2(n12971), .ZN(
        n13213) );
  NAND2_X1 U15100 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13021)
         );
  OAI21_X1 U15101 ( .B1(n13213), .B2(n12937), .A(n13021), .ZN(n12923) );
  AOI21_X1 U15102 ( .B1(n13222), .B2(n12935), .A(n12923), .ZN(n12924) );
  OAI211_X1 U15103 ( .C1(n13225), .C2(n12926), .A(n12925), .B(n12924), .ZN(
        P2_U3210) );
  INV_X1 U15104 ( .A(n12849), .ZN(n12931) );
  NOR3_X1 U15105 ( .A1(n12929), .A2(n12928), .A3(n12927), .ZN(n12930) );
  AOI21_X1 U15106 ( .B1(n12931), .B2(n12946), .A(n12930), .ZN(n12944) );
  AOI22_X1 U15107 ( .A1(n12962), .A2(n12933), .B1(n12932), .B2(n12964), .ZN(
        n13095) );
  INV_X1 U15108 ( .A(n12934), .ZN(n13101) );
  AOI22_X1 U15109 ( .A1(n13101), .A2(n12935), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12936) );
  OAI21_X1 U15110 ( .B1(n13095), .B2(n12937), .A(n12936), .ZN(n12941) );
  NOR2_X1 U15111 ( .A1(n12939), .A2(n12938), .ZN(n12940) );
  AOI211_X1 U15112 ( .C1(n13287), .C2(n8784), .A(n12941), .B(n12940), .ZN(
        n12942) );
  OAI21_X1 U15113 ( .B1(n12944), .B2(n12943), .A(n12942), .ZN(P2_U3212) );
  AOI22_X1 U15114 ( .A1(n12947), .A2(n12946), .B1(n12945), .B2(n12973), .ZN(
        n12958) );
  INV_X1 U15115 ( .A(n12948), .ZN(n12957) );
  AOI22_X1 U15116 ( .A1(n12950), .A2(n12949), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12951) );
  OAI21_X1 U15117 ( .B1(n12953), .B2(n12952), .A(n12951), .ZN(n12954) );
  AOI21_X1 U15118 ( .B1(n12955), .B2(n8784), .A(n12954), .ZN(n12956) );
  OAI21_X1 U15119 ( .B1(n12958), .B2(n12957), .A(n12956), .ZN(P2_U3213) );
  MUX2_X1 U15120 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13053), .S(P2_U3947), .Z(
        P2_U3562) );
  MUX2_X1 U15121 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n12959), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15122 ( .A(n12960), .B(P2_DATAO_REG_29__SCAN_IN), .S(n12987), .Z(
        P2_U3560) );
  MUX2_X1 U15123 ( .A(n12961), .B(P2_DATAO_REG_28__SCAN_IN), .S(n12987), .Z(
        P2_U3559) );
  MUX2_X1 U15124 ( .A(n12962), .B(P2_DATAO_REG_27__SCAN_IN), .S(n12987), .Z(
        P2_U3558) );
  MUX2_X1 U15125 ( .A(n12963), .B(P2_DATAO_REG_26__SCAN_IN), .S(n12987), .Z(
        P2_U3557) );
  MUX2_X1 U15126 ( .A(n12964), .B(P2_DATAO_REG_25__SCAN_IN), .S(n12987), .Z(
        P2_U3556) );
  MUX2_X1 U15127 ( .A(n12965), .B(P2_DATAO_REG_24__SCAN_IN), .S(n12987), .Z(
        P2_U3555) );
  MUX2_X1 U15128 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n12966), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U15129 ( .A(n12967), .B(P2_DATAO_REG_21__SCAN_IN), .S(n12987), .Z(
        P2_U3552) );
  MUX2_X1 U15130 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n12968), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U15131 ( .A(n12969), .B(P2_DATAO_REG_19__SCAN_IN), .S(n12987), .Z(
        P2_U3550) );
  MUX2_X1 U15132 ( .A(n12970), .B(P2_DATAO_REG_18__SCAN_IN), .S(n12987), .Z(
        P2_U3549) );
  MUX2_X1 U15133 ( .A(n12971), .B(P2_DATAO_REG_17__SCAN_IN), .S(n12987), .Z(
        P2_U3548) );
  MUX2_X1 U15134 ( .A(n12972), .B(P2_DATAO_REG_16__SCAN_IN), .S(n12987), .Z(
        P2_U3547) );
  MUX2_X1 U15135 ( .A(n12973), .B(P2_DATAO_REG_15__SCAN_IN), .S(n12987), .Z(
        P2_U3546) );
  MUX2_X1 U15136 ( .A(n12974), .B(P2_DATAO_REG_14__SCAN_IN), .S(n12987), .Z(
        P2_U3545) );
  MUX2_X1 U15137 ( .A(n12975), .B(P2_DATAO_REG_13__SCAN_IN), .S(n12987), .Z(
        P2_U3544) );
  MUX2_X1 U15138 ( .A(n12976), .B(P2_DATAO_REG_12__SCAN_IN), .S(n12987), .Z(
        P2_U3543) );
  MUX2_X1 U15139 ( .A(n12977), .B(P2_DATAO_REG_11__SCAN_IN), .S(n12987), .Z(
        P2_U3542) );
  MUX2_X1 U15140 ( .A(n12978), .B(P2_DATAO_REG_10__SCAN_IN), .S(n12987), .Z(
        P2_U3541) );
  MUX2_X1 U15141 ( .A(n12979), .B(P2_DATAO_REG_9__SCAN_IN), .S(n12987), .Z(
        P2_U3540) );
  MUX2_X1 U15142 ( .A(n12980), .B(P2_DATAO_REG_8__SCAN_IN), .S(n12987), .Z(
        P2_U3539) );
  MUX2_X1 U15143 ( .A(n12981), .B(P2_DATAO_REG_7__SCAN_IN), .S(n12987), .Z(
        P2_U3538) );
  MUX2_X1 U15144 ( .A(n12982), .B(P2_DATAO_REG_6__SCAN_IN), .S(n12987), .Z(
        P2_U3537) );
  MUX2_X1 U15145 ( .A(n12983), .B(P2_DATAO_REG_5__SCAN_IN), .S(n12987), .Z(
        P2_U3536) );
  MUX2_X1 U15146 ( .A(n12984), .B(P2_DATAO_REG_4__SCAN_IN), .S(n12987), .Z(
        P2_U3535) );
  MUX2_X1 U15147 ( .A(n12985), .B(P2_DATAO_REG_3__SCAN_IN), .S(n12987), .Z(
        P2_U3534) );
  MUX2_X1 U15148 ( .A(n12986), .B(P2_DATAO_REG_2__SCAN_IN), .S(n12987), .Z(
        P2_U3533) );
  MUX2_X1 U15149 ( .A(n12988), .B(P2_DATAO_REG_1__SCAN_IN), .S(n12987), .Z(
        P2_U3532) );
  MUX2_X1 U15150 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n9597), .S(P2_U3947), .Z(
        P2_U3531) );
  OAI211_X1 U15151 ( .C1(n12991), .C2(n12990), .A(n14976), .B(n12989), .ZN(
        n13001) );
  AOI22_X1 U15152 ( .A1(n15007), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3088), .ZN(n13000) );
  INV_X1 U15153 ( .A(n15014), .ZN(n14991) );
  NAND2_X1 U15154 ( .A1(n14991), .A2(n12992), .ZN(n12999) );
  INV_X1 U15155 ( .A(n12993), .ZN(n12997) );
  NAND3_X1 U15156 ( .A1(n14963), .A2(n12995), .A3(n12994), .ZN(n12996) );
  NAND3_X1 U15157 ( .A1(n15009), .A2(n12997), .A3(n12996), .ZN(n12998) );
  NAND4_X1 U15158 ( .A1(n13001), .A2(n13000), .A3(n12999), .A4(n12998), .ZN(
        P2_U3217) );
  AND2_X1 U15159 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13002) );
  AOI21_X1 U15160 ( .B1(n14991), .B2(n13024), .A(n13002), .ZN(n13003) );
  INV_X1 U15161 ( .A(n13003), .ZN(n13009) );
  AOI21_X1 U15162 ( .B1(n13005), .B2(P2_REG1_REG_16__SCAN_IN), .A(n13004), 
        .ZN(n13007) );
  XNOR2_X1 U15163 ( .A(n13024), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n13006) );
  NOR2_X1 U15164 ( .A1(n13007), .A2(n13006), .ZN(n13023) );
  AOI211_X1 U15165 ( .C1(n13007), .C2(n13006), .A(n13023), .B(n15001), .ZN(
        n13008) );
  AOI211_X1 U15166 ( .C1(n15007), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n13009), 
        .B(n13008), .ZN(n13016) );
  OAI21_X1 U15167 ( .B1(n13011), .B2(n11651), .A(n13010), .ZN(n13014) );
  INV_X1 U15168 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13019) );
  NOR2_X1 U15169 ( .A1(n13018), .A2(n13019), .ZN(n13012) );
  AOI21_X1 U15170 ( .B1(n13019), .B2(n13018), .A(n13012), .ZN(n13013) );
  NAND2_X1 U15171 ( .A1(n13013), .A2(n13014), .ZN(n13017) );
  OAI211_X1 U15172 ( .C1(n13014), .C2(n13013), .A(n15009), .B(n13017), .ZN(
        n13015) );
  NAND2_X1 U15173 ( .A1(n13016), .A2(n13015), .ZN(P2_U3231) );
  OAI21_X1 U15174 ( .B1(n13019), .B2(n13018), .A(n13017), .ZN(n13032) );
  XNOR2_X1 U15175 ( .A(n13033), .B(n13032), .ZN(n13020) );
  NOR2_X1 U15176 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13020), .ZN(n13034) );
  AOI21_X1 U15177 ( .B1(n13020), .B2(P2_REG2_REG_18__SCAN_IN), .A(n13034), 
        .ZN(n13031) );
  OAI21_X1 U15178 ( .B1(n15014), .B2(n13037), .A(n13021), .ZN(n13022) );
  AOI21_X1 U15179 ( .B1(n15007), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n13022), 
        .ZN(n13030) );
  INV_X1 U15180 ( .A(n13025), .ZN(n13028) );
  INV_X1 U15181 ( .A(n13040), .ZN(n13027) );
  OAI211_X1 U15182 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n13028), .A(n14976), 
        .B(n13027), .ZN(n13029) );
  OAI211_X1 U15183 ( .C1(n13031), .C2(n14993), .A(n13030), .B(n13029), .ZN(
        P2_U3232) );
  INV_X1 U15184 ( .A(n15007), .ZN(n15000) );
  NOR2_X1 U15185 ( .A1(n13033), .A2(n13032), .ZN(n13035) );
  NOR2_X1 U15186 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  XOR2_X1 U15187 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n13036), .Z(n13046) );
  INV_X1 U15188 ( .A(n13046), .ZN(n13044) );
  NOR2_X1 U15189 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  XOR2_X1 U15190 ( .A(n13042), .B(n13041), .Z(n13045) );
  OAI21_X1 U15191 ( .B1(n13045), .B2(n15001), .A(n15014), .ZN(n13043) );
  AOI21_X1 U15192 ( .B1(n13044), .B2(n15009), .A(n13043), .ZN(n13049) );
  AOI22_X1 U15193 ( .A1(n13046), .A2(n15009), .B1(n14976), .B2(n13045), .ZN(
        n13048) );
  MUX2_X1 U15194 ( .A(n13049), .B(n13048), .S(n13047), .Z(n13051) );
  OAI211_X1 U15195 ( .C1(n7495), .C2(n15000), .A(n13051), .B(n13050), .ZN(
        P2_U3233) );
  NAND2_X1 U15196 ( .A1(n13058), .A2(n13267), .ZN(n13057) );
  NAND2_X1 U15197 ( .A1(n13054), .A2(n13053), .ZN(n13265) );
  NOR2_X1 U15198 ( .A1(n13242), .A2(n13265), .ZN(n13060) );
  NOR2_X1 U15199 ( .A1(n7195), .A2(n13236), .ZN(n13055) );
  AOI211_X1 U15200 ( .C1(n15038), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13060), 
        .B(n13055), .ZN(n13056) );
  OAI21_X1 U15201 ( .B1(n13264), .B2(n15023), .A(n13056), .ZN(P2_U3234) );
  OAI211_X1 U15202 ( .C1(n13058), .C2(n13267), .A(n15021), .B(n13057), .ZN(
        n13266) );
  NOR2_X1 U15203 ( .A1(n13267), .A2(n13236), .ZN(n13059) );
  AOI211_X1 U15204 ( .C1(n15038), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13060), 
        .B(n13059), .ZN(n13061) );
  OAI21_X1 U15205 ( .B1(n15023), .B2(n13266), .A(n13061), .ZN(P2_U3235) );
  OAI211_X1 U15206 ( .C1(n13064), .C2(n13063), .A(n13062), .B(n15018), .ZN(
        n13066) );
  OAI21_X1 U15207 ( .B1(n13069), .B2(n13068), .A(n13067), .ZN(n13277) );
  INV_X1 U15208 ( .A(n13277), .ZN(n13077) );
  OR2_X1 U15209 ( .A1(n13075), .A2(n6585), .ZN(n13070) );
  AND3_X1 U15210 ( .A1(n13071), .A2(n15021), .A3(n13070), .ZN(n13273) );
  NAND2_X1 U15211 ( .A1(n13273), .A2(n13259), .ZN(n13074) );
  AOI22_X1 U15212 ( .A1(n13072), .A2(n13254), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n13242), .ZN(n13073) );
  OAI211_X1 U15213 ( .C1(n13075), .C2(n13236), .A(n13074), .B(n13073), .ZN(
        n13076) );
  AOI21_X1 U15214 ( .B1(n13077), .B2(n15035), .A(n13076), .ZN(n13078) );
  OAI21_X1 U15215 ( .B1(n13276), .B2(n15038), .A(n13078), .ZN(P2_U3237) );
  NOR2_X1 U15216 ( .A1(n13090), .A2(n13079), .ZN(n13080) );
  OR2_X1 U15217 ( .A1(n13081), .A2(n13080), .ZN(n13083) );
  AOI21_X1 U15218 ( .B1(n13083), .B2(n15018), .A(n13082), .ZN(n13285) );
  NAND2_X1 U15219 ( .A1(n13280), .A2(n13098), .ZN(n13084) );
  NAND2_X1 U15220 ( .A1(n13084), .A2(n15021), .ZN(n13085) );
  OR2_X1 U15221 ( .A1(n6585), .A2(n13085), .ZN(n13281) );
  AOI22_X1 U15222 ( .A1(n13086), .A2(n13254), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n13242), .ZN(n13088) );
  NAND2_X1 U15223 ( .A1(n13280), .A2(n15027), .ZN(n13087) );
  OAI211_X1 U15224 ( .C1(n13281), .C2(n15023), .A(n13088), .B(n13087), .ZN(
        n13089) );
  INV_X1 U15225 ( .A(n13089), .ZN(n13092) );
  NAND2_X1 U15226 ( .A1(n6625), .A2(n13090), .ZN(n13279) );
  NAND3_X1 U15227 ( .A1(n13279), .A2(n13278), .A3(n15035), .ZN(n13091) );
  OAI211_X1 U15228 ( .C1(n13285), .C2(n15038), .A(n13092), .B(n13091), .ZN(
        P2_U3238) );
  OAI21_X1 U15229 ( .B1(n13105), .B2(n13094), .A(n13093), .ZN(n13097) );
  INV_X1 U15230 ( .A(n13095), .ZN(n13096) );
  AOI21_X1 U15231 ( .B1(n13097), .B2(n15018), .A(n13096), .ZN(n13288) );
  INV_X1 U15232 ( .A(n13112), .ZN(n13100) );
  INV_X1 U15233 ( .A(n13098), .ZN(n13099) );
  AOI211_X1 U15234 ( .C1(n13287), .C2(n13100), .A(n13219), .B(n13099), .ZN(
        n13286) );
  AOI22_X1 U15235 ( .A1(n13101), .A2(n13254), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13242), .ZN(n13102) );
  OAI21_X1 U15236 ( .B1(n13103), .B2(n13236), .A(n13102), .ZN(n13107) );
  XOR2_X1 U15237 ( .A(n13104), .B(n13105), .Z(n13290) );
  NOR2_X1 U15238 ( .A1(n13290), .A2(n13246), .ZN(n13106) );
  AOI211_X1 U15239 ( .C1(n13286), .C2(n13259), .A(n13107), .B(n13106), .ZN(
        n13108) );
  OAI21_X1 U15240 ( .B1(n15038), .B2(n13288), .A(n13108), .ZN(P2_U3239) );
  XOR2_X1 U15241 ( .A(n13109), .B(n13118), .Z(n13295) );
  NAND2_X1 U15242 ( .A1(n13292), .A2(n13133), .ZN(n13110) );
  NAND2_X1 U15243 ( .A1(n13110), .A2(n15021), .ZN(n13111) );
  NOR2_X1 U15244 ( .A1(n13112), .A2(n13111), .ZN(n13291) );
  NAND2_X1 U15245 ( .A1(n13292), .A2(n15027), .ZN(n13114) );
  NAND2_X1 U15246 ( .A1(n13242), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13113) );
  OAI211_X1 U15247 ( .C1(n15050), .C2(n13115), .A(n13114), .B(n13113), .ZN(
        n13122) );
  OAI21_X1 U15248 ( .B1(n13118), .B2(n13117), .A(n13116), .ZN(n13120) );
  AOI21_X1 U15249 ( .B1(n13120), .B2(n15018), .A(n13119), .ZN(n13294) );
  NOR2_X1 U15250 ( .A1(n13294), .A2(n13242), .ZN(n13121) );
  AOI211_X1 U15251 ( .C1(n13291), .C2(n13259), .A(n13122), .B(n13121), .ZN(
        n13123) );
  OAI21_X1 U15252 ( .B1(n13246), .B2(n13295), .A(n13123), .ZN(P2_U3240) );
  OAI21_X1 U15253 ( .B1(n13126), .B2(n13125), .A(n13124), .ZN(n13128) );
  AOI21_X1 U15254 ( .B1(n13128), .B2(n15018), .A(n13127), .ZN(n13299) );
  OR2_X1 U15255 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  NAND2_X1 U15256 ( .A1(n13132), .A2(n13131), .ZN(n13300) );
  INV_X1 U15257 ( .A(n13300), .ZN(n13140) );
  AOI21_X1 U15258 ( .B1(n13297), .B2(n13145), .A(n13219), .ZN(n13134) );
  AND2_X1 U15259 ( .A1(n13134), .A2(n13133), .ZN(n13296) );
  NAND2_X1 U15260 ( .A1(n13296), .A2(n13259), .ZN(n13137) );
  AOI22_X1 U15261 ( .A1(n13135), .A2(n13254), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n13242), .ZN(n13136) );
  OAI211_X1 U15262 ( .C1(n13138), .C2(n13236), .A(n13137), .B(n13136), .ZN(
        n13139) );
  AOI21_X1 U15263 ( .B1(n13140), .B2(n15035), .A(n13139), .ZN(n13141) );
  OAI21_X1 U15264 ( .B1(n13299), .B2(n15038), .A(n13141), .ZN(P2_U3241) );
  XNOR2_X1 U15265 ( .A(n13142), .B(n13151), .ZN(n13144) );
  AOI21_X1 U15266 ( .B1(n13144), .B2(n15018), .A(n13143), .ZN(n13304) );
  AOI21_X1 U15267 ( .B1(n13302), .B2(n13156), .A(n13219), .ZN(n13146) );
  AND2_X1 U15268 ( .A1(n13146), .A2(n13145), .ZN(n13301) );
  NAND2_X1 U15269 ( .A1(n13302), .A2(n15027), .ZN(n13148) );
  NAND2_X1 U15270 ( .A1(n15038), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n13147) );
  OAI211_X1 U15271 ( .C1(n15050), .C2(n13149), .A(n13148), .B(n13147), .ZN(
        n13153) );
  XNOR2_X1 U15272 ( .A(n13150), .B(n13151), .ZN(n13305) );
  NOR2_X1 U15273 ( .A1(n13305), .A2(n13246), .ZN(n13152) );
  AOI211_X1 U15274 ( .C1(n13301), .C2(n13259), .A(n13153), .B(n13152), .ZN(
        n13154) );
  OAI21_X1 U15275 ( .B1(n15038), .B2(n13304), .A(n13154), .ZN(P2_U3242) );
  XNOR2_X1 U15276 ( .A(n13155), .B(n13161), .ZN(n13310) );
  INV_X1 U15277 ( .A(n13156), .ZN(n13157) );
  AOI211_X1 U15278 ( .C1(n13307), .C2(n13171), .A(n13219), .B(n13157), .ZN(
        n13306) );
  INV_X1 U15279 ( .A(n13307), .ZN(n13160) );
  AOI22_X1 U15280 ( .A1(n13158), .A2(n13254), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13242), .ZN(n13159) );
  OAI21_X1 U15281 ( .B1(n13160), .B2(n13236), .A(n13159), .ZN(n13168) );
  AOI21_X1 U15282 ( .B1(n13162), .B2(n13161), .A(n15039), .ZN(n13166) );
  INV_X1 U15283 ( .A(n13163), .ZN(n13164) );
  AOI21_X1 U15284 ( .B1(n13166), .B2(n6714), .A(n13164), .ZN(n13309) );
  NOR2_X1 U15285 ( .A1(n13309), .A2(n13242), .ZN(n13167) );
  AOI211_X1 U15286 ( .C1(n13306), .C2(n13259), .A(n13168), .B(n13167), .ZN(
        n13169) );
  OAI21_X1 U15287 ( .B1(n13246), .B2(n13310), .A(n13169), .ZN(P2_U3243) );
  XNOR2_X1 U15288 ( .A(n13170), .B(n13178), .ZN(n13315) );
  INV_X1 U15289 ( .A(n13192), .ZN(n13173) );
  INV_X1 U15290 ( .A(n13171), .ZN(n13172) );
  AOI211_X1 U15291 ( .C1(n13312), .C2(n13173), .A(n13219), .B(n13172), .ZN(
        n13311) );
  INV_X1 U15292 ( .A(n13174), .ZN(n13175) );
  AOI22_X1 U15293 ( .A1(n13175), .A2(n13254), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n13242), .ZN(n13176) );
  OAI21_X1 U15294 ( .B1(n13177), .B2(n13236), .A(n13176), .ZN(n13183) );
  XOR2_X1 U15295 ( .A(n13179), .B(n13178), .Z(n13181) );
  AOI21_X1 U15296 ( .B1(n13181), .B2(n15018), .A(n13180), .ZN(n13314) );
  NOR2_X1 U15297 ( .A1(n13314), .A2(n13242), .ZN(n13182) );
  AOI211_X1 U15298 ( .C1(n13311), .C2(n13259), .A(n13183), .B(n13182), .ZN(
        n13184) );
  OAI21_X1 U15299 ( .B1(n13246), .B2(n13315), .A(n13184), .ZN(P2_U3244) );
  XOR2_X1 U15300 ( .A(n13185), .B(n13189), .Z(n13320) );
  INV_X1 U15301 ( .A(n13186), .ZN(n13187) );
  AOI21_X1 U15302 ( .B1(n13189), .B2(n13188), .A(n13187), .ZN(n13191) );
  OAI21_X1 U15303 ( .B1(n13191), .B2(n15039), .A(n13190), .ZN(n13316) );
  AOI211_X1 U15304 ( .C1(n13318), .C2(n13200), .A(n13219), .B(n13192), .ZN(
        n13317) );
  NAND2_X1 U15305 ( .A1(n13317), .A2(n13259), .ZN(n13195) );
  AOI22_X1 U15306 ( .A1(n13193), .A2(n13254), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n13242), .ZN(n13194) );
  OAI211_X1 U15307 ( .C1(n13196), .C2(n13236), .A(n13195), .B(n13194), .ZN(
        n13197) );
  AOI21_X1 U15308 ( .B1(n13316), .B2(n15048), .A(n13197), .ZN(n13198) );
  OAI21_X1 U15309 ( .B1(n13246), .B2(n13320), .A(n13198), .ZN(P2_U3245) );
  XOR2_X1 U15310 ( .A(n13199), .B(n13204), .Z(n13325) );
  INV_X1 U15311 ( .A(n13200), .ZN(n13201) );
  AOI211_X1 U15312 ( .C1(n13323), .C2(n13220), .A(n13219), .B(n13201), .ZN(
        n13322) );
  INV_X1 U15313 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13202) );
  OAI22_X1 U15314 ( .A1(n7200), .A2(n13236), .B1(n13202), .B2(n15048), .ZN(
        n13203) );
  AOI21_X1 U15315 ( .B1(n13322), .B2(n13259), .A(n13203), .ZN(n13211) );
  XNOR2_X1 U15316 ( .A(n13205), .B(n13204), .ZN(n13207) );
  OAI21_X1 U15317 ( .B1(n13207), .B2(n15039), .A(n13206), .ZN(n13321) );
  NOR2_X1 U15318 ( .A1(n13208), .A2(n15050), .ZN(n13209) );
  OAI21_X1 U15319 ( .B1(n13321), .B2(n13209), .A(n15048), .ZN(n13210) );
  OAI211_X1 U15320 ( .C1(n13325), .C2(n13246), .A(n13211), .B(n13210), .ZN(
        P2_U3246) );
  XNOR2_X1 U15321 ( .A(n13212), .B(n13217), .ZN(n13215) );
  INV_X1 U15322 ( .A(n13213), .ZN(n13214) );
  AOI21_X1 U15323 ( .B1(n13215), .B2(n15018), .A(n13214), .ZN(n13330) );
  OAI21_X1 U15324 ( .B1(n13218), .B2(n13217), .A(n13216), .ZN(n13326) );
  AOI21_X1 U15325 ( .B1(n13328), .B2(n13230), .A(n13219), .ZN(n13221) );
  AND2_X1 U15326 ( .A1(n13221), .A2(n13220), .ZN(n13327) );
  NAND2_X1 U15327 ( .A1(n13327), .A2(n13259), .ZN(n13224) );
  AOI22_X1 U15328 ( .A1(n13242), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13222), 
        .B2(n13254), .ZN(n13223) );
  OAI211_X1 U15329 ( .C1(n13225), .C2(n13236), .A(n13224), .B(n13223), .ZN(
        n13226) );
  AOI21_X1 U15330 ( .B1(n13326), .B2(n15035), .A(n13226), .ZN(n13227) );
  OAI21_X1 U15331 ( .B1(n15038), .B2(n13330), .A(n13227), .ZN(P2_U3247) );
  XOR2_X1 U15332 ( .A(n13228), .B(n13238), .Z(n13336) );
  INV_X1 U15333 ( .A(n13229), .ZN(n13232) );
  INV_X1 U15334 ( .A(n13230), .ZN(n13231) );
  AOI211_X1 U15335 ( .C1(n13333), .C2(n13232), .A(n13219), .B(n13231), .ZN(
        n13332) );
  NOR2_X1 U15336 ( .A1(n13233), .A2(n15050), .ZN(n13234) );
  AOI21_X1 U15337 ( .B1(n15038), .B2(P2_REG2_REG_17__SCAN_IN), .A(n13234), 
        .ZN(n13235) );
  OAI21_X1 U15338 ( .B1(n13237), .B2(n13236), .A(n13235), .ZN(n13244) );
  XNOR2_X1 U15339 ( .A(n13239), .B(n13238), .ZN(n13241) );
  AOI21_X1 U15340 ( .B1(n13241), .B2(n15018), .A(n13240), .ZN(n13335) );
  NOR2_X1 U15341 ( .A1(n13335), .A2(n13242), .ZN(n13243) );
  AOI211_X1 U15342 ( .C1(n13332), .C2(n13259), .A(n13244), .B(n13243), .ZN(
        n13245) );
  OAI21_X1 U15343 ( .B1(n13246), .B2(n13336), .A(n13245), .ZN(P2_U3248) );
  OAI21_X1 U15344 ( .B1(n13248), .B2(n13255), .A(n13247), .ZN(n13251) );
  INV_X1 U15345 ( .A(n13249), .ZN(n13250) );
  AOI21_X1 U15346 ( .B1(n13251), .B2(n15018), .A(n13250), .ZN(n15109) );
  MUX2_X1 U15347 ( .A(n13252), .B(n15109), .S(n15048), .Z(n13263) );
  AOI22_X1 U15348 ( .A1(n15027), .A2(n15106), .B1(n13254), .B2(n13253), .ZN(
        n13262) );
  NAND2_X1 U15349 ( .A1(n13256), .A2(n13255), .ZN(n15103) );
  NAND3_X1 U15350 ( .A1(n15104), .A2(n15103), .A3(n15035), .ZN(n13261) );
  AOI211_X1 U15351 ( .C1(n15106), .C2(n13258), .A(n13219), .B(n13257), .ZN(
        n15105) );
  NAND2_X1 U15352 ( .A1(n15105), .A2(n13259), .ZN(n13260) );
  NAND4_X1 U15353 ( .A1(n13263), .A2(n13262), .A3(n13261), .A4(n13260), .ZN(
        P2_U3259) );
  MUX2_X1 U15354 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13353), .S(n15160), .Z(
        P2_U3530) );
  OAI211_X1 U15355 ( .C1(n13267), .C2(n15146), .A(n13266), .B(n13265), .ZN(
        n13354) );
  MUX2_X1 U15356 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13354), .S(n15160), .Z(
        P2_U3529) );
  AOI21_X1 U15357 ( .B1(n15137), .B2(n13270), .A(n13269), .ZN(n13271) );
  MUX2_X1 U15358 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13355), .S(n15160), .Z(
        P2_U3528) );
  AOI21_X1 U15359 ( .B1(n15137), .B2(n13274), .A(n13273), .ZN(n13275) );
  OAI211_X1 U15360 ( .C1(n13351), .C2(n13277), .A(n13276), .B(n13275), .ZN(
        n13356) );
  MUX2_X1 U15361 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13356), .S(n15160), .Z(
        P2_U3527) );
  NAND3_X1 U15362 ( .A1(n13279), .A2(n15151), .A3(n13278), .ZN(n13283) );
  NAND2_X1 U15363 ( .A1(n13280), .A2(n15137), .ZN(n13282) );
  NAND2_X1 U15364 ( .A1(n13285), .A2(n13284), .ZN(n13357) );
  MUX2_X1 U15365 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13357), .S(n15160), .Z(
        P2_U3526) );
  AOI21_X1 U15366 ( .B1(n15137), .B2(n13287), .A(n13286), .ZN(n13289) );
  OAI211_X1 U15367 ( .C1(n13351), .C2(n13290), .A(n13289), .B(n13288), .ZN(
        n13358) );
  MUX2_X1 U15368 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13358), .S(n15160), .Z(
        P2_U3525) );
  AOI21_X1 U15369 ( .B1(n15137), .B2(n13292), .A(n13291), .ZN(n13293) );
  OAI211_X1 U15370 ( .C1(n13295), .C2(n13351), .A(n13294), .B(n13293), .ZN(
        n13359) );
  MUX2_X1 U15371 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13359), .S(n15160), .Z(
        P2_U3524) );
  AOI21_X1 U15372 ( .B1(n15137), .B2(n13297), .A(n13296), .ZN(n13298) );
  OAI211_X1 U15373 ( .C1(n13351), .C2(n13300), .A(n13299), .B(n13298), .ZN(
        n13360) );
  MUX2_X1 U15374 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13360), .S(n15160), .Z(
        P2_U3523) );
  AOI21_X1 U15375 ( .B1(n15137), .B2(n13302), .A(n13301), .ZN(n13303) );
  OAI211_X1 U15376 ( .C1(n13305), .C2(n13351), .A(n13304), .B(n13303), .ZN(
        n13361) );
  MUX2_X1 U15377 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13361), .S(n15160), .Z(
        P2_U3522) );
  AOI21_X1 U15378 ( .B1(n15137), .B2(n13307), .A(n13306), .ZN(n13308) );
  OAI211_X1 U15379 ( .C1(n13310), .C2(n13351), .A(n13309), .B(n13308), .ZN(
        n13362) );
  MUX2_X1 U15380 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13362), .S(n15160), .Z(
        P2_U3521) );
  AOI21_X1 U15381 ( .B1(n15137), .B2(n13312), .A(n13311), .ZN(n13313) );
  OAI211_X1 U15382 ( .C1(n13315), .C2(n13351), .A(n13314), .B(n13313), .ZN(
        n13363) );
  MUX2_X1 U15383 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13363), .S(n15160), .Z(
        P2_U3520) );
  AOI211_X1 U15384 ( .C1(n15137), .C2(n13318), .A(n13317), .B(n13316), .ZN(
        n13319) );
  OAI21_X1 U15385 ( .B1(n13351), .B2(n13320), .A(n13319), .ZN(n13364) );
  MUX2_X1 U15386 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13364), .S(n15160), .Z(
        P2_U3519) );
  AOI211_X1 U15387 ( .C1(n15137), .C2(n13323), .A(n13322), .B(n13321), .ZN(
        n13324) );
  OAI21_X1 U15388 ( .B1(n13325), .B2(n13351), .A(n13324), .ZN(n13365) );
  MUX2_X1 U15389 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13365), .S(n15160), .Z(
        P2_U3518) );
  INV_X1 U15390 ( .A(n13326), .ZN(n13331) );
  AOI21_X1 U15391 ( .B1(n15137), .B2(n13328), .A(n13327), .ZN(n13329) );
  OAI211_X1 U15392 ( .C1(n13331), .C2(n13351), .A(n13330), .B(n13329), .ZN(
        n13366) );
  MUX2_X1 U15393 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13366), .S(n15160), .Z(
        P2_U3517) );
  AOI21_X1 U15394 ( .B1(n15137), .B2(n13333), .A(n13332), .ZN(n13334) );
  OAI211_X1 U15395 ( .C1(n13336), .C2(n13351), .A(n13335), .B(n13334), .ZN(
        n13367) );
  MUX2_X1 U15396 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13367), .S(n15160), .Z(
        P2_U3516) );
  AOI211_X1 U15397 ( .C1(n15137), .C2(n13339), .A(n13338), .B(n13337), .ZN(
        n13340) );
  OAI21_X1 U15398 ( .B1(n13351), .B2(n13341), .A(n13340), .ZN(n13368) );
  MUX2_X1 U15399 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13368), .S(n15160), .Z(
        P2_U3515) );
  AOI211_X1 U15400 ( .C1(n15137), .C2(n13344), .A(n13343), .B(n13342), .ZN(
        n13345) );
  OAI21_X1 U15401 ( .B1(n13351), .B2(n13346), .A(n13345), .ZN(n13369) );
  MUX2_X1 U15402 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n13369), .S(n15160), .Z(
        P2_U3513) );
  AOI21_X1 U15403 ( .B1(n15137), .B2(n13348), .A(n13347), .ZN(n13349) );
  OAI211_X1 U15404 ( .C1(n13352), .C2(n13351), .A(n13350), .B(n13349), .ZN(
        n13370) );
  MUX2_X1 U15405 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13370), .S(n15160), .Z(
        P2_U3511) );
  MUX2_X1 U15406 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13354), .S(n15155), .Z(
        P2_U3497) );
  MUX2_X1 U15407 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13355), .S(n15155), .Z(
        P2_U3496) );
  MUX2_X1 U15408 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13356), .S(n15155), .Z(
        P2_U3495) );
  MUX2_X1 U15409 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13357), .S(n15155), .Z(
        P2_U3494) );
  MUX2_X1 U15410 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13358), .S(n15155), .Z(
        P2_U3493) );
  MUX2_X1 U15411 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13359), .S(n15155), .Z(
        P2_U3492) );
  MUX2_X1 U15412 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13360), .S(n15155), .Z(
        P2_U3491) );
  MUX2_X1 U15413 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13361), .S(n15155), .Z(
        P2_U3490) );
  MUX2_X1 U15414 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13362), .S(n15155), .Z(
        P2_U3489) );
  MUX2_X1 U15415 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13363), .S(n15155), .Z(
        P2_U3488) );
  MUX2_X1 U15416 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13364), .S(n15155), .Z(
        P2_U3487) );
  MUX2_X1 U15417 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13365), .S(n15155), .Z(
        P2_U3486) );
  MUX2_X1 U15418 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13366), .S(n15155), .Z(
        P2_U3484) );
  MUX2_X1 U15419 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13367), .S(n15155), .Z(
        P2_U3481) );
  MUX2_X1 U15420 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13368), .S(n15155), .Z(
        P2_U3478) );
  MUX2_X1 U15421 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n13369), .S(n15155), .Z(
        P2_U3472) );
  MUX2_X1 U15422 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n13370), .S(n15155), .Z(
        P2_U3466) );
  INV_X1 U15423 ( .A(n13371), .ZN(n14446) );
  NAND3_X1 U15424 ( .A1(n13373), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n13375) );
  OAI22_X1 U15425 ( .A1(n13372), .A2(n13375), .B1(n13374), .B2(n13395), .ZN(
        n13376) );
  INV_X1 U15426 ( .A(n13376), .ZN(n13377) );
  OAI21_X1 U15427 ( .B1(n14446), .B2(n13393), .A(n13377), .ZN(P2_U3296) );
  INV_X1 U15428 ( .A(n13378), .ZN(n14448) );
  OAI222_X1 U15429 ( .A1(n13393), .A2(n14448), .B1(n13379), .B2(P2_U3088), 
        .C1(n13488), .C2(n13395), .ZN(P2_U3297) );
  NAND2_X1 U15430 ( .A1(n9458), .A2(n13380), .ZN(n13382) );
  OAI211_X1 U15431 ( .C1(n13395), .C2(n13383), .A(n13382), .B(n13381), .ZN(
        P2_U3299) );
  INV_X1 U15432 ( .A(n13384), .ZN(n14453) );
  OAI222_X1 U15433 ( .A1(n13395), .A2(n13386), .B1(n13393), .B2(n14453), .C1(
        P2_U3088), .C2(n13385), .ZN(P2_U3300) );
  INV_X1 U15434 ( .A(n13387), .ZN(n13389) );
  OAI222_X1 U15435 ( .A1(n13393), .A2(n13390), .B1(n13389), .B2(P2_U3088), 
        .C1(n13388), .C2(n13395), .ZN(P2_U3301) );
  INV_X1 U15436 ( .A(n13391), .ZN(n14457) );
  OAI222_X1 U15437 ( .A1(n13395), .A2(n13394), .B1(n13393), .B2(n14457), .C1(
        P2_U3088), .C2(n13392), .ZN(P2_U3302) );
  MUX2_X1 U15438 ( .A(n13397), .B(n13396), .S(P2_STATE_REG_SCAN_IN), .Z(n13672) );
  NAND4_X1 U15439 ( .A1(keyinput50), .A2(keyinput62), .A3(keyinput113), .A4(
        keyinput14), .ZN(n13413) );
  NOR2_X1 U15440 ( .A1(keyinput40), .A2(keyinput74), .ZN(n13398) );
  NAND3_X1 U15441 ( .A1(keyinput24), .A2(keyinput70), .A3(n13398), .ZN(n13412)
         );
  NOR2_X1 U15442 ( .A1(keyinput90), .A2(keyinput42), .ZN(n13399) );
  NAND3_X1 U15443 ( .A1(keyinput123), .A2(keyinput17), .A3(n13399), .ZN(n13400) );
  NOR3_X1 U15444 ( .A1(keyinput96), .A2(keyinput46), .A3(n13400), .ZN(n13401)
         );
  NAND3_X1 U15445 ( .A1(keyinput64), .A2(keyinput32), .A3(n13401), .ZN(n13411)
         );
  NAND2_X1 U15446 ( .A1(keyinput23), .A2(keyinput71), .ZN(n13402) );
  NOR3_X1 U15447 ( .A1(keyinput66), .A2(keyinput58), .A3(n13402), .ZN(n13409)
         );
  INV_X1 U15448 ( .A(keyinput124), .ZN(n13403) );
  NOR4_X1 U15449 ( .A1(keyinput105), .A2(keyinput111), .A3(keyinput122), .A4(
        n13403), .ZN(n13408) );
  INV_X1 U15450 ( .A(keyinput8), .ZN(n13404) );
  NOR4_X1 U15451 ( .A1(keyinput84), .A2(keyinput99), .A3(keyinput16), .A4(
        n13404), .ZN(n13407) );
  NAND2_X1 U15452 ( .A1(keyinput88), .A2(keyinput26), .ZN(n13405) );
  NOR3_X1 U15453 ( .A1(keyinput125), .A2(keyinput87), .A3(n13405), .ZN(n13406)
         );
  NAND4_X1 U15454 ( .A1(n13409), .A2(n13408), .A3(n13407), .A4(n13406), .ZN(
        n13410) );
  NOR4_X1 U15455 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13461) );
  INV_X1 U15456 ( .A(keyinput54), .ZN(n13416) );
  NOR2_X1 U15457 ( .A1(keyinput95), .A2(keyinput13), .ZN(n13414) );
  NAND3_X1 U15458 ( .A1(keyinput44), .A2(keyinput92), .A3(n13414), .ZN(n13415)
         );
  NOR4_X1 U15459 ( .A1(keyinput104), .A2(keyinput39), .A3(n13416), .A4(n13415), 
        .ZN(n13428) );
  NAND3_X1 U15460 ( .A1(keyinput100), .A2(keyinput76), .A3(keyinput5), .ZN(
        n13417) );
  NOR2_X1 U15461 ( .A1(keyinput7), .A2(n13417), .ZN(n13427) );
  NOR4_X1 U15462 ( .A1(keyinput12), .A2(keyinput52), .A3(keyinput127), .A4(
        keyinput3), .ZN(n13426) );
  INV_X1 U15463 ( .A(keyinput101), .ZN(n13418) );
  NAND4_X1 U15464 ( .A1(keyinput79), .A2(keyinput0), .A3(keyinput30), .A4(
        n13418), .ZN(n13424) );
  OR4_X1 U15465 ( .A1(keyinput86), .A2(keyinput56), .A3(keyinput93), .A4(
        keyinput34), .ZN(n13423) );
  NOR2_X1 U15466 ( .A1(keyinput61), .A2(keyinput35), .ZN(n13419) );
  NAND3_X1 U15467 ( .A1(keyinput18), .A2(keyinput4), .A3(n13419), .ZN(n13422)
         );
  INV_X1 U15468 ( .A(keyinput102), .ZN(n13420) );
  NAND4_X1 U15469 ( .A1(keyinput38), .A2(keyinput41), .A3(keyinput6), .A4(
        n13420), .ZN(n13421) );
  NOR4_X1 U15470 ( .A1(n13424), .A2(n13423), .A3(n13422), .A4(n13421), .ZN(
        n13425) );
  NAND4_X1 U15471 ( .A1(n13428), .A2(n13427), .A3(n13426), .A4(n13425), .ZN(
        n13459) );
  NAND2_X1 U15472 ( .A1(keyinput112), .A2(keyinput57), .ZN(n13429) );
  NOR3_X1 U15473 ( .A1(keyinput85), .A2(keyinput2), .A3(n13429), .ZN(n13435)
         );
  INV_X1 U15474 ( .A(keyinput72), .ZN(n13430) );
  NOR4_X1 U15475 ( .A1(keyinput31), .A2(keyinput59), .A3(keyinput91), .A4(
        n13430), .ZN(n13434) );
  NOR4_X1 U15476 ( .A1(keyinput109), .A2(keyinput51), .A3(keyinput37), .A4(
        keyinput77), .ZN(n13433) );
  NAND3_X1 U15477 ( .A1(keyinput89), .A2(keyinput69), .A3(keyinput80), .ZN(
        n13431) );
  NOR2_X1 U15478 ( .A1(keyinput43), .A2(n13431), .ZN(n13432) );
  NAND4_X1 U15479 ( .A1(n13435), .A2(n13434), .A3(n13433), .A4(n13432), .ZN(
        n13458) );
  NAND3_X1 U15480 ( .A1(keyinput28), .A2(keyinput121), .A3(keyinput116), .ZN(
        n13436) );
  NOR2_X1 U15481 ( .A1(keyinput47), .A2(n13436), .ZN(n13441) );
  NOR4_X1 U15482 ( .A1(keyinput60), .A2(keyinput120), .A3(keyinput11), .A4(
        keyinput63), .ZN(n13440) );
  NOR4_X1 U15483 ( .A1(keyinput27), .A2(keyinput118), .A3(keyinput49), .A4(
        keyinput78), .ZN(n13439) );
  NAND2_X1 U15484 ( .A1(keyinput53), .A2(keyinput110), .ZN(n13437) );
  NOR3_X1 U15485 ( .A1(keyinput20), .A2(keyinput33), .A3(n13437), .ZN(n13438)
         );
  NAND4_X1 U15486 ( .A1(n13441), .A2(n13440), .A3(n13439), .A4(n13438), .ZN(
        n13457) );
  NAND4_X1 U15487 ( .A1(keyinput21), .A2(keyinput15), .A3(keyinput25), .A4(
        keyinput114), .ZN(n13442) );
  NOR3_X1 U15488 ( .A1(keyinput29), .A2(keyinput65), .A3(n13442), .ZN(n13455)
         );
  INV_X1 U15489 ( .A(keyinput36), .ZN(n13443) );
  NAND4_X1 U15490 ( .A1(keyinput83), .A2(keyinput68), .A3(keyinput55), .A4(
        n13443), .ZN(n13453) );
  NOR2_X1 U15491 ( .A1(keyinput19), .A2(keyinput126), .ZN(n13444) );
  NAND3_X1 U15492 ( .A1(keyinput97), .A2(keyinput73), .A3(n13444), .ZN(n13452)
         );
  NOR4_X1 U15493 ( .A1(keyinput48), .A2(keyinput119), .A3(keyinput67), .A4(
        keyinput103), .ZN(n13450) );
  INV_X1 U15494 ( .A(keyinput108), .ZN(n13445) );
  NOR4_X1 U15495 ( .A1(keyinput10), .A2(keyinput45), .A3(keyinput117), .A4(
        n13445), .ZN(n13449) );
  NOR4_X1 U15496 ( .A1(keyinput82), .A2(keyinput22), .A3(keyinput115), .A4(
        keyinput1), .ZN(n13448) );
  INV_X1 U15497 ( .A(keyinput81), .ZN(n13446) );
  NOR4_X1 U15498 ( .A1(keyinput75), .A2(keyinput107), .A3(keyinput106), .A4(
        n13446), .ZN(n13447) );
  NAND4_X1 U15499 ( .A1(n13450), .A2(n13449), .A3(n13448), .A4(n13447), .ZN(
        n13451) );
  NOR3_X1 U15500 ( .A1(n13453), .A2(n13452), .A3(n13451), .ZN(n13454) );
  NAND4_X1 U15501 ( .A1(keyinput94), .A2(keyinput98), .A3(n13455), .A4(n13454), 
        .ZN(n13456) );
  NOR4_X1 U15502 ( .A1(n13459), .A2(n13458), .A3(n13457), .A4(n13456), .ZN(
        n13460) );
  AOI21_X1 U15503 ( .B1(n13461), .B2(n13460), .A(keyinput9), .ZN(n13670) );
  INV_X1 U15504 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U15505 ( .A1(n13463), .A2(keyinput63), .B1(keyinput121), .B2(n15428), .ZN(n13462) );
  OAI221_X1 U15506 ( .B1(n13463), .B2(keyinput63), .C1(n15428), .C2(
        keyinput121), .A(n13462), .ZN(n13474) );
  AOI22_X1 U15507 ( .A1(n8661), .A2(keyinput47), .B1(keyinput20), .B2(n13465), 
        .ZN(n13464) );
  OAI221_X1 U15508 ( .B1(n8661), .B2(keyinput47), .C1(n13465), .C2(keyinput20), 
        .A(n13464), .ZN(n13473) );
  INV_X1 U15509 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U15510 ( .A1(n13468), .A2(keyinput116), .B1(n13467), .B2(keyinput28), .ZN(n13466) );
  OAI221_X1 U15511 ( .B1(n13468), .B2(keyinput116), .C1(n13467), .C2(
        keyinput28), .A(n13466), .ZN(n13472) );
  XOR2_X1 U15512 ( .A(n13863), .B(keyinput120), .Z(n13470) );
  XNOR2_X1 U15513 ( .A(P2_IR_REG_24__SCAN_IN), .B(keyinput11), .ZN(n13469) );
  NAND2_X1 U15514 ( .A1(n13470), .A2(n13469), .ZN(n13471) );
  NOR4_X1 U15515 ( .A1(n13474), .A2(n13473), .A3(n13472), .A4(n13471), .ZN(
        n13513) );
  INV_X1 U15516 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U15517 ( .A1(n14695), .A2(keyinput110), .B1(n13476), .B2(keyinput27), .ZN(n13475) );
  OAI221_X1 U15518 ( .B1(n14695), .B2(keyinput110), .C1(n13476), .C2(
        keyinput27), .A(n13475), .ZN(n13486) );
  INV_X1 U15519 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U15520 ( .A1(n13478), .A2(keyinput118), .B1(n15154), .B2(keyinput53), .ZN(n13477) );
  OAI221_X1 U15521 ( .B1(n13478), .B2(keyinput118), .C1(n15154), .C2(
        keyinput53), .A(n13477), .ZN(n13485) );
  AOI22_X1 U15522 ( .A1(n13481), .A2(keyinput33), .B1(n13480), .B2(keyinput49), 
        .ZN(n13479) );
  OAI221_X1 U15523 ( .B1(n13481), .B2(keyinput33), .C1(n13480), .C2(keyinput49), .A(n13479), .ZN(n13484) );
  AOI22_X1 U15524 ( .A1(n15064), .A2(keyinput78), .B1(keyinput31), .B2(n11311), 
        .ZN(n13482) );
  OAI221_X1 U15525 ( .B1(n15064), .B2(keyinput78), .C1(n11311), .C2(keyinput31), .A(n13482), .ZN(n13483) );
  NOR4_X1 U15526 ( .A1(n13486), .A2(n13485), .A3(n13484), .A4(n13483), .ZN(
        n13512) );
  AOI22_X1 U15527 ( .A1(n13489), .A2(keyinput2), .B1(keyinput69), .B2(n13488), 
        .ZN(n13487) );
  OAI221_X1 U15528 ( .B1(n13489), .B2(keyinput2), .C1(n13488), .C2(keyinput69), 
        .A(n13487), .ZN(n13494) );
  INV_X1 U15529 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14319) );
  AOI22_X1 U15530 ( .A1(n13491), .A2(keyinput59), .B1(keyinput72), .B2(n14319), 
        .ZN(n13490) );
  OAI221_X1 U15531 ( .B1(n13491), .B2(keyinput59), .C1(n14319), .C2(keyinput72), .A(n13490), .ZN(n13493) );
  XOR2_X1 U15532 ( .A(P2_REG2_REG_0__SCAN_IN), .B(keyinput57), .Z(n13492) );
  OR3_X1 U15533 ( .A1(n13494), .A2(n13493), .A3(n13492), .ZN(n13498) );
  INV_X1 U15534 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14850) );
  INV_X1 U15535 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n14546) );
  AOI22_X1 U15536 ( .A1(n14850), .A2(keyinput91), .B1(keyinput85), .B2(n14546), 
        .ZN(n13495) );
  OAI221_X1 U15537 ( .B1(n14850), .B2(keyinput91), .C1(n14546), .C2(keyinput85), .A(n13495), .ZN(n13497) );
  INV_X1 U15538 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14851) );
  XNOR2_X1 U15539 ( .A(n14851), .B(keyinput112), .ZN(n13496) );
  NOR3_X1 U15540 ( .A1(n13498), .A2(n13497), .A3(n13496), .ZN(n13511) );
  AOI22_X1 U15541 ( .A1(P1_U3086), .A2(keyinput80), .B1(n13500), .B2(
        keyinput43), .ZN(n13499) );
  OAI221_X1 U15542 ( .B1(P1_U3086), .B2(keyinput80), .C1(n13500), .C2(
        keyinput43), .A(n13499), .ZN(n13509) );
  AOI22_X1 U15543 ( .A1(n14484), .A2(keyinput89), .B1(n13502), .B2(keyinput109), .ZN(n13501) );
  OAI221_X1 U15544 ( .B1(n14484), .B2(keyinput89), .C1(n13502), .C2(
        keyinput109), .A(n13501), .ZN(n13508) );
  AOI22_X1 U15545 ( .A1(n13504), .A2(keyinput51), .B1(n14450), .B2(keyinput37), 
        .ZN(n13503) );
  OAI221_X1 U15546 ( .B1(n13504), .B2(keyinput51), .C1(n14450), .C2(keyinput37), .A(n13503), .ZN(n13507) );
  AOI22_X1 U15547 ( .A1(n11370), .A2(keyinput77), .B1(n15052), .B2(keyinput10), 
        .ZN(n13505) );
  OAI221_X1 U15548 ( .B1(n11370), .B2(keyinput77), .C1(n15052), .C2(keyinput10), .A(n13505), .ZN(n13506) );
  NOR4_X1 U15549 ( .A1(n13509), .A2(n13508), .A3(n13507), .A4(n13506), .ZN(
        n13510) );
  NAND4_X1 U15550 ( .A1(n13513), .A2(n13512), .A3(n13511), .A4(n13510), .ZN(
        n13668) );
  INV_X1 U15551 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n13515) );
  AOI22_X1 U15552 ( .A1(n13515), .A2(keyinput45), .B1(n10797), .B2(keyinput108), .ZN(n13514) );
  OAI221_X1 U15553 ( .B1(n13515), .B2(keyinput45), .C1(n10797), .C2(
        keyinput108), .A(n13514), .ZN(n13524) );
  INV_X1 U15554 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15093) );
  AOI22_X1 U15555 ( .A1(n13517), .A2(keyinput117), .B1(n15093), .B2(keyinput48), .ZN(n13516) );
  OAI221_X1 U15556 ( .B1(n13517), .B2(keyinput117), .C1(n15093), .C2(
        keyinput48), .A(n13516), .ZN(n13523) );
  XNOR2_X1 U15557 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput119), .ZN(n13521) );
  XNOR2_X1 U15558 ( .A(P3_IR_REG_26__SCAN_IN), .B(keyinput67), .ZN(n13520) );
  XNOR2_X1 U15559 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput94), .ZN(n13519)
         );
  XNOR2_X1 U15560 ( .A(SI_5_), .B(keyinput103), .ZN(n13518) );
  NAND4_X1 U15561 ( .A1(n13521), .A2(n13520), .A3(n13519), .A4(n13518), .ZN(
        n13522) );
  NOR3_X1 U15562 ( .A1(n13524), .A2(n13523), .A3(n13522), .ZN(n13563) );
  AOI22_X1 U15563 ( .A1(n8318), .A2(keyinput98), .B1(n13526), .B2(keyinput21), 
        .ZN(n13525) );
  OAI221_X1 U15564 ( .B1(n8318), .B2(keyinput98), .C1(n13526), .C2(keyinput21), 
        .A(n13525), .ZN(n13537) );
  INV_X1 U15565 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n13529) );
  AOI22_X1 U15566 ( .A1(n13529), .A2(keyinput15), .B1(n13528), .B2(keyinput25), 
        .ZN(n13527) );
  OAI221_X1 U15567 ( .B1(n13529), .B2(keyinput15), .C1(n13528), .C2(keyinput25), .A(n13527), .ZN(n13536) );
  AOI22_X1 U15568 ( .A1(n10876), .A2(keyinput114), .B1(n13396), .B2(keyinput29), .ZN(n13530) );
  OAI221_X1 U15569 ( .B1(n10876), .B2(keyinput114), .C1(n13396), .C2(
        keyinput29), .A(n13530), .ZN(n13535) );
  AOI22_X1 U15570 ( .A1(n13533), .A2(keyinput65), .B1(n13532), .B2(keyinput75), 
        .ZN(n13531) );
  OAI221_X1 U15571 ( .B1(n13533), .B2(keyinput65), .C1(n13532), .C2(keyinput75), .A(n13531), .ZN(n13534) );
  NOR4_X1 U15572 ( .A1(n13537), .A2(n13536), .A3(n13535), .A4(n13534), .ZN(
        n13562) );
  INV_X1 U15573 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14839) );
  AOI22_X1 U15574 ( .A1(n14839), .A2(keyinput1), .B1(n10123), .B2(keyinput19), 
        .ZN(n13538) );
  OAI221_X1 U15575 ( .B1(n14839), .B2(keyinput1), .C1(n10123), .C2(keyinput19), 
        .A(n13538), .ZN(n13547) );
  AOI22_X1 U15576 ( .A1(n11324), .A2(keyinput22), .B1(n13540), .B2(keyinput115), .ZN(n13539) );
  OAI221_X1 U15577 ( .B1(n11324), .B2(keyinput22), .C1(n13540), .C2(
        keyinput115), .A(n13539), .ZN(n13546) );
  XOR2_X1 U15578 ( .A(n8276), .B(keyinput106), .Z(n13544) );
  XNOR2_X1 U15579 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput107), .ZN(n13543)
         );
  XNOR2_X1 U15580 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput81), .ZN(n13542) );
  XNOR2_X1 U15581 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput82), .ZN(n13541)
         );
  NAND4_X1 U15582 ( .A1(n13544), .A2(n13543), .A3(n13542), .A4(n13541), .ZN(
        n13545) );
  NOR3_X1 U15583 ( .A1(n13547), .A2(n13546), .A3(n13545), .ZN(n13561) );
  AOI22_X1 U15584 ( .A1(n14480), .A2(keyinput104), .B1(keyinput55), .B2(n13549), .ZN(n13548) );
  OAI221_X1 U15585 ( .B1(n14480), .B2(keyinput104), .C1(n13549), .C2(
        keyinput55), .A(n13548), .ZN(n13559) );
  AOI22_X1 U15586 ( .A1(n10558), .A2(keyinput83), .B1(n13551), .B2(keyinput36), 
        .ZN(n13550) );
  OAI221_X1 U15587 ( .B1(n10558), .B2(keyinput83), .C1(n13551), .C2(keyinput36), .A(n13550), .ZN(n13558) );
  INV_X1 U15588 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n13553) );
  OAI221_X1 U15589 ( .B1(n13553), .B2(keyinput73), .C1(n13877), .C2(keyinput68), .A(n13552), .ZN(n13557) );
  XOR2_X1 U15590 ( .A(n9474), .B(keyinput97), .Z(n13555) );
  XNOR2_X1 U15591 ( .A(P3_IR_REG_8__SCAN_IN), .B(keyinput126), .ZN(n13554) );
  NAND2_X1 U15592 ( .A1(n13555), .A2(n13554), .ZN(n13556) );
  NOR4_X1 U15593 ( .A1(n13559), .A2(n13558), .A3(n13557), .A4(n13556), .ZN(
        n13560) );
  NAND4_X1 U15594 ( .A1(n13563), .A2(n13562), .A3(n13561), .A4(n13560), .ZN(
        n13667) );
  AOI22_X1 U15595 ( .A1(n13565), .A2(keyinput62), .B1(n14636), .B2(keyinput70), 
        .ZN(n13564) );
  OAI221_X1 U15596 ( .B1(n13565), .B2(keyinput62), .C1(n14636), .C2(keyinput70), .A(n13564), .ZN(n13575) );
  INV_X1 U15597 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n13567) );
  AOI22_X1 U15598 ( .A1(n13567), .A2(keyinput24), .B1(keyinput50), .B2(n9406), 
        .ZN(n13566) );
  OAI221_X1 U15599 ( .B1(n13567), .B2(keyinput24), .C1(n9406), .C2(keyinput50), 
        .A(n13566), .ZN(n13574) );
  AOI22_X1 U15600 ( .A1(n13570), .A2(keyinput14), .B1(keyinput26), .B2(n13569), 
        .ZN(n13568) );
  OAI221_X1 U15601 ( .B1(n13570), .B2(keyinput14), .C1(n13569), .C2(keyinput26), .A(n13568), .ZN(n13573) );
  INV_X1 U15602 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14520) );
  AOI22_X1 U15603 ( .A1(n14520), .A2(keyinput74), .B1(n8004), .B2(keyinput113), 
        .ZN(n13571) );
  OAI221_X1 U15604 ( .B1(n14520), .B2(keyinput74), .C1(n8004), .C2(keyinput113), .A(n13571), .ZN(n13572) );
  NOR4_X1 U15605 ( .A1(n13575), .A2(n13574), .A3(n13573), .A4(n13572), .ZN(
        n13612) );
  INV_X1 U15606 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U15607 ( .A1(n14479), .A2(keyinput66), .B1(n9143), .B2(keyinput23), 
        .ZN(n13576) );
  OAI221_X1 U15608 ( .B1(n14479), .B2(keyinput66), .C1(n9143), .C2(keyinput23), 
        .A(n13576), .ZN(n13586) );
  AOI22_X1 U15609 ( .A1(n13579), .A2(keyinput122), .B1(keyinput71), .B2(n13578), .ZN(n13577) );
  OAI221_X1 U15610 ( .B1(n13579), .B2(keyinput122), .C1(n13578), .C2(
        keyinput71), .A(n13577), .ZN(n13585) );
  XOR2_X1 U15611 ( .A(n8584), .B(keyinput40), .Z(n13583) );
  XNOR2_X1 U15612 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput124), .ZN(n13582) );
  XNOR2_X1 U15613 ( .A(P3_REG0_REG_23__SCAN_IN), .B(keyinput111), .ZN(n13581)
         );
  XNOR2_X1 U15614 ( .A(SI_0_), .B(keyinput58), .ZN(n13580) );
  NAND4_X1 U15615 ( .A1(n13583), .A2(n13582), .A3(n13581), .A4(n13580), .ZN(
        n13584) );
  NOR3_X1 U15616 ( .A1(n13586), .A2(n13585), .A3(n13584), .ZN(n13611) );
  AOI22_X1 U15617 ( .A1(n11651), .A2(keyinput90), .B1(n13588), .B2(keyinput96), 
        .ZN(n13587) );
  OAI221_X1 U15618 ( .B1(n11651), .B2(keyinput90), .C1(n13588), .C2(keyinput96), .A(n13587), .ZN(n13598) );
  AOI22_X1 U15619 ( .A1(n13591), .A2(keyinput32), .B1(n13590), .B2(keyinput123), .ZN(n13589) );
  OAI221_X1 U15620 ( .B1(n13591), .B2(keyinput32), .C1(n13590), .C2(
        keyinput123), .A(n13589), .ZN(n13597) );
  INV_X1 U15621 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14843) );
  AOI22_X1 U15622 ( .A1(n13593), .A2(keyinput42), .B1(keyinput60), .B2(n14843), 
        .ZN(n13592) );
  OAI221_X1 U15623 ( .B1(n13593), .B2(keyinput42), .C1(n14843), .C2(keyinput60), .A(n13592), .ZN(n13596) );
  INV_X1 U15624 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14840) );
  AOI22_X1 U15625 ( .A1(n10064), .A2(keyinput46), .B1(keyinput17), .B2(n14840), 
        .ZN(n13594) );
  OAI221_X1 U15626 ( .B1(n10064), .B2(keyinput46), .C1(n14840), .C2(keyinput17), .A(n13594), .ZN(n13595) );
  NOR4_X1 U15627 ( .A1(n13598), .A2(n13597), .A3(n13596), .A4(n13595), .ZN(
        n13610) );
  AOI22_X1 U15628 ( .A1(n13600), .A2(keyinput87), .B1(keyinput84), .B2(n7557), 
        .ZN(n13599) );
  OAI221_X1 U15629 ( .B1(n13600), .B2(keyinput87), .C1(n7557), .C2(keyinput84), 
        .A(n13599), .ZN(n13608) );
  INV_X1 U15630 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14848) );
  AOI22_X1 U15631 ( .A1(n13602), .A2(keyinput125), .B1(n14848), .B2(keyinput88), .ZN(n13601) );
  OAI221_X1 U15632 ( .B1(n13602), .B2(keyinput125), .C1(n14848), .C2(
        keyinput88), .A(n13601), .ZN(n13607) );
  AOI22_X1 U15633 ( .A1(n7605), .A2(keyinput16), .B1(keyinput64), .B2(n8299), 
        .ZN(n13603) );
  OAI221_X1 U15634 ( .B1(n7605), .B2(keyinput16), .C1(n8299), .C2(keyinput64), 
        .A(n13603), .ZN(n13606) );
  INV_X1 U15635 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14707) );
  INV_X1 U15636 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14838) );
  AOI22_X1 U15637 ( .A1(n14707), .A2(keyinput99), .B1(n14838), .B2(keyinput8), 
        .ZN(n13604) );
  OAI221_X1 U15638 ( .B1(n14707), .B2(keyinput99), .C1(n14838), .C2(keyinput8), 
        .A(n13604), .ZN(n13605) );
  NOR4_X1 U15639 ( .A1(n13608), .A2(n13607), .A3(n13606), .A4(n13605), .ZN(
        n13609) );
  NAND4_X1 U15640 ( .A1(n13612), .A2(n13611), .A3(n13610), .A4(n13609), .ZN(
        n13666) );
  AOI22_X1 U15641 ( .A1(n13614), .A2(keyinput52), .B1(keyinput127), .B2(n14463), .ZN(n13613) );
  OAI221_X1 U15642 ( .B1(n13614), .B2(keyinput52), .C1(n14463), .C2(
        keyinput127), .A(n13613), .ZN(n13624) );
  AOI22_X1 U15643 ( .A1(n13617), .A2(keyinput100), .B1(keyinput86), .B2(n13616), .ZN(n13615) );
  OAI221_X1 U15644 ( .B1(n13617), .B2(keyinput100), .C1(n13616), .C2(
        keyinput86), .A(n13615), .ZN(n13623) );
  XNOR2_X1 U15645 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput5), .ZN(n13621) );
  XNOR2_X1 U15646 ( .A(P3_REG2_REG_0__SCAN_IN), .B(keyinput3), .ZN(n13620) );
  XNOR2_X1 U15647 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput7), .ZN(n13619) );
  XNOR2_X1 U15648 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput76), .ZN(n13618) );
  NAND4_X1 U15649 ( .A1(n13621), .A2(n13620), .A3(n13619), .A4(n13618), .ZN(
        n13622) );
  NOR3_X1 U15650 ( .A1(n13624), .A2(n13623), .A3(n13622), .ZN(n13664) );
  INV_X1 U15651 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14841) );
  NAND2_X1 U15652 ( .A1(n13626), .A2(keyinput44), .ZN(n13625) );
  OAI221_X1 U15653 ( .B1(n14841), .B2(keyinput9), .C1(n13626), .C2(keyinput44), 
        .A(n13625), .ZN(n13638) );
  AOI22_X1 U15654 ( .A1(n13629), .A2(keyinput54), .B1(n13628), .B2(keyinput39), 
        .ZN(n13627) );
  OAI221_X1 U15655 ( .B1(n13629), .B2(keyinput54), .C1(n13628), .C2(keyinput39), .A(n13627), .ZN(n13637) );
  INV_X1 U15656 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14741) );
  AOI22_X1 U15657 ( .A1(n13631), .A2(keyinput13), .B1(keyinput12), .B2(n14741), 
        .ZN(n13630) );
  OAI221_X1 U15658 ( .B1(n13631), .B2(keyinput13), .C1(n14741), .C2(keyinput12), .A(n13630), .ZN(n13636) );
  AOI22_X1 U15659 ( .A1(n13634), .A2(keyinput95), .B1(n13633), .B2(keyinput92), 
        .ZN(n13632) );
  OAI221_X1 U15660 ( .B1(n13634), .B2(keyinput95), .C1(n13633), .C2(keyinput92), .A(n13632), .ZN(n13635) );
  NOR4_X1 U15661 ( .A1(n13638), .A2(n13637), .A3(n13636), .A4(n13635), .ZN(
        n13663) );
  AOI22_X1 U15662 ( .A1(n8235), .A2(keyinput4), .B1(keyinput105), .B2(n10103), 
        .ZN(n13639) );
  OAI221_X1 U15663 ( .B1(n8235), .B2(keyinput4), .C1(n10103), .C2(keyinput105), 
        .A(n13639), .ZN(n13648) );
  AOI22_X1 U15664 ( .A1(n15058), .A2(keyinput38), .B1(n7686), .B2(keyinput41), 
        .ZN(n13640) );
  OAI221_X1 U15665 ( .B1(n15058), .B2(keyinput38), .C1(n7686), .C2(keyinput41), 
        .A(n13640), .ZN(n13647) );
  XOR2_X1 U15666 ( .A(n13641), .B(keyinput6), .Z(n13645) );
  XNOR2_X1 U15667 ( .A(P3_IR_REG_1__SCAN_IN), .B(keyinput61), .ZN(n13644) );
  XNOR2_X1 U15668 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput18), .ZN(n13643) );
  XNOR2_X1 U15669 ( .A(P1_REG3_REG_5__SCAN_IN), .B(keyinput35), .ZN(n13642) );
  NAND4_X1 U15670 ( .A1(n13645), .A2(n13644), .A3(n13643), .A4(n13642), .ZN(
        n13646) );
  NOR3_X1 U15671 ( .A1(n13648), .A2(n13647), .A3(n13646), .ZN(n13662) );
  AOI22_X1 U15672 ( .A1(n13650), .A2(keyinput56), .B1(keyinput93), .B2(n9047), 
        .ZN(n13649) );
  OAI221_X1 U15673 ( .B1(n13650), .B2(keyinput56), .C1(n9047), .C2(keyinput93), 
        .A(n13649), .ZN(n13660) );
  AOI22_X1 U15674 ( .A1(n13652), .A2(keyinput34), .B1(keyinput101), .B2(n9424), 
        .ZN(n13651) );
  OAI221_X1 U15675 ( .B1(n13652), .B2(keyinput34), .C1(n9424), .C2(keyinput101), .A(n13651), .ZN(n13659) );
  AOI22_X1 U15676 ( .A1(n13774), .A2(keyinput79), .B1(n13654), .B2(keyinput0), 
        .ZN(n13653) );
  OAI221_X1 U15677 ( .B1(n13774), .B2(keyinput79), .C1(n13654), .C2(keyinput0), 
        .A(n13653), .ZN(n13658) );
  XNOR2_X1 U15678 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(keyinput102), .ZN(n13656)
         );
  XNOR2_X1 U15679 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput30), .ZN(n13655) );
  NAND2_X1 U15680 ( .A1(n13656), .A2(n13655), .ZN(n13657) );
  NOR4_X1 U15681 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13661) );
  NAND4_X1 U15682 ( .A1(n13664), .A2(n13663), .A3(n13662), .A4(n13661), .ZN(
        n13665) );
  NOR4_X1 U15683 ( .A1(n13668), .A2(n13667), .A3(n13666), .A4(n13665), .ZN(
        n13669) );
  OAI21_X1 U15684 ( .B1(P1_D_REG_24__SCAN_IN), .B2(n13670), .A(n13669), .ZN(
        n13671) );
  XOR2_X1 U15685 ( .A(n13672), .B(n13671), .Z(P2_U3327) );
  NAND2_X1 U15686 ( .A1(n14343), .A2(n13798), .ZN(n13674) );
  NAND2_X1 U15687 ( .A1(n14158), .A2(n9891), .ZN(n13673) );
  NAND2_X1 U15688 ( .A1(n13674), .A2(n13673), .ZN(n13675) );
  XNOR2_X1 U15689 ( .A(n13675), .B(n6549), .ZN(n13794) );
  AOI22_X1 U15690 ( .A1(n14343), .A2(n9891), .B1(n9892), .B2(n14158), .ZN(
        n13795) );
  XNOR2_X1 U15691 ( .A(n13794), .B(n13795), .ZN(n13797) );
  AND2_X1 U15692 ( .A1(n14290), .A2(n9892), .ZN(n13676) );
  AOI21_X1 U15693 ( .B1(n14392), .B2(n9891), .A(n13676), .ZN(n13727) );
  NAND2_X1 U15694 ( .A1(n14392), .A2(n13798), .ZN(n13678) );
  NAND2_X1 U15695 ( .A1(n14290), .A2(n9891), .ZN(n13677) );
  NAND2_X1 U15696 ( .A1(n13678), .A2(n13677), .ZN(n13680) );
  XNOR2_X1 U15697 ( .A(n13680), .B(n6549), .ZN(n13726) );
  INV_X1 U15698 ( .A(n13681), .ZN(n13683) );
  NAND2_X1 U15699 ( .A1(n13684), .A2(n7431), .ZN(n13861) );
  AND2_X1 U15700 ( .A1(n9892), .A2(n13912), .ZN(n13685) );
  AOI21_X1 U15701 ( .B1(n13869), .B2(n9891), .A(n13685), .ZN(n13688) );
  AOI22_X1 U15702 ( .A1(n13869), .A2(n13798), .B1(n9891), .B2(n13912), .ZN(
        n13686) );
  XNOR2_X1 U15703 ( .A(n13686), .B(n6549), .ZN(n13687) );
  XOR2_X1 U15704 ( .A(n13688), .B(n13687), .Z(n13862) );
  INV_X1 U15705 ( .A(n13687), .ZN(n13690) );
  INV_X1 U15706 ( .A(n13688), .ZN(n13689) );
  NAND2_X1 U15707 ( .A1(n14658), .A2(n13798), .ZN(n13692) );
  NAND2_X1 U15708 ( .A1(n13911), .A2(n9891), .ZN(n13691) );
  NAND2_X1 U15709 ( .A1(n13692), .A2(n13691), .ZN(n13693) );
  XNOR2_X1 U15710 ( .A(n13693), .B(n6549), .ZN(n13697) );
  NAND2_X1 U15711 ( .A1(n14658), .A2(n9891), .ZN(n13695) );
  NAND2_X1 U15712 ( .A1(n9892), .A2(n13911), .ZN(n13694) );
  NAND2_X1 U15713 ( .A1(n13695), .A2(n13694), .ZN(n13696) );
  NOR2_X1 U15714 ( .A1(n13697), .A2(n13696), .ZN(n13698) );
  AOI21_X1 U15715 ( .B1(n13697), .B2(n13696), .A(n13698), .ZN(n14657) );
  OAI22_X1 U15716 ( .A1(n6955), .A2(n9886), .B1(n14661), .B2(n13729), .ZN(
        n13699) );
  XNOR2_X1 U15717 ( .A(n13699), .B(n6549), .ZN(n13702) );
  OAI22_X1 U15718 ( .A1(n6955), .A2(n13729), .B1(n14661), .B2(n13728), .ZN(
        n13898) );
  INV_X1 U15719 ( .A(n13700), .ZN(n13701) );
  NAND2_X1 U15720 ( .A1(n14086), .A2(n13798), .ZN(n13704) );
  NAND2_X1 U15721 ( .A1(n14311), .A2(n9891), .ZN(n13703) );
  NAND2_X1 U15722 ( .A1(n13704), .A2(n13703), .ZN(n13705) );
  XNOR2_X1 U15723 ( .A(n13705), .B(n6549), .ZN(n13709) );
  NAND2_X1 U15724 ( .A1(n14086), .A2(n9891), .ZN(n13707) );
  NAND2_X1 U15725 ( .A1(n9892), .A2(n14311), .ZN(n13706) );
  NAND2_X1 U15726 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  NOR2_X1 U15727 ( .A1(n13709), .A2(n13708), .ZN(n13710) );
  AOI21_X1 U15728 ( .B1(n13709), .B2(n13708), .A(n13710), .ZN(n13829) );
  INV_X1 U15729 ( .A(n13710), .ZN(n13711) );
  NAND2_X1 U15730 ( .A1(n14310), .A2(n13798), .ZN(n13713) );
  NAND2_X1 U15731 ( .A1(n14088), .A2(n9891), .ZN(n13712) );
  NAND2_X1 U15732 ( .A1(n13713), .A2(n13712), .ZN(n13714) );
  XNOR2_X1 U15733 ( .A(n13714), .B(n6549), .ZN(n13718) );
  NAND2_X1 U15734 ( .A1(n14310), .A2(n9891), .ZN(n13716) );
  NAND2_X1 U15735 ( .A1(n14088), .A2(n9892), .ZN(n13715) );
  NAND2_X1 U15736 ( .A1(n13716), .A2(n13715), .ZN(n13717) );
  NAND2_X1 U15737 ( .A1(n13718), .A2(n13717), .ZN(n13837) );
  AOI22_X1 U15738 ( .A1(n14398), .A2(n9891), .B1(n9892), .B2(n14313), .ZN(
        n13722) );
  NAND2_X1 U15739 ( .A1(n14398), .A2(n13798), .ZN(n13720) );
  NAND2_X1 U15740 ( .A1(n14313), .A2(n9891), .ZN(n13719) );
  NAND2_X1 U15741 ( .A1(n13720), .A2(n13719), .ZN(n13721) );
  XNOR2_X1 U15742 ( .A(n13721), .B(n6549), .ZN(n13724) );
  XOR2_X1 U15743 ( .A(n13722), .B(n13724), .Z(n13882) );
  INV_X1 U15744 ( .A(n13722), .ZN(n13723) );
  OR2_X1 U15745 ( .A1(n13724), .A2(n13723), .ZN(n13725) );
  XOR2_X1 U15746 ( .A(n13727), .B(n13726), .Z(n13787) );
  OAI22_X1 U15747 ( .A1(n14261), .A2(n13729), .B1(n14239), .B2(n13728), .ZN(
        n13732) );
  OAI22_X1 U15748 ( .A1(n14261), .A2(n9886), .B1(n14239), .B2(n13729), .ZN(
        n13730) );
  XNOR2_X1 U15749 ( .A(n13730), .B(n6549), .ZN(n13731) );
  XOR2_X1 U15750 ( .A(n13732), .B(n13731), .Z(n13854) );
  NAND2_X1 U15751 ( .A1(n13855), .A2(n13854), .ZN(n13853) );
  NAND2_X1 U15752 ( .A1(n13731), .A2(n13732), .ZN(n13733) );
  AOI22_X1 U15753 ( .A1(n14381), .A2(n13798), .B1(n9891), .B2(n14252), .ZN(
        n13734) );
  XNOR2_X1 U15754 ( .A(n13734), .B(n6549), .ZN(n13736) );
  AOI22_X1 U15755 ( .A1(n14381), .A2(n9891), .B1(n9892), .B2(n14252), .ZN(
        n13737) );
  XNOR2_X1 U15756 ( .A(n13736), .B(n13737), .ZN(n13811) );
  INV_X1 U15757 ( .A(n13811), .ZN(n13735) );
  NAND2_X1 U15758 ( .A1(n13736), .A2(n13737), .ZN(n13738) );
  NAND2_X1 U15759 ( .A1(n14375), .A2(n13798), .ZN(n13740) );
  NAND2_X1 U15760 ( .A1(n14074), .A2(n9891), .ZN(n13739) );
  NAND2_X1 U15761 ( .A1(n13740), .A2(n13739), .ZN(n13741) );
  XNOR2_X1 U15762 ( .A(n13741), .B(n6549), .ZN(n13744) );
  AOI22_X1 U15763 ( .A1(n14375), .A2(n9891), .B1(n9892), .B2(n14074), .ZN(
        n13742) );
  XNOR2_X1 U15764 ( .A(n13744), .B(n13742), .ZN(n13875) );
  INV_X1 U15765 ( .A(n13742), .ZN(n13743) );
  NAND2_X1 U15766 ( .A1(n14369), .A2(n13798), .ZN(n13747) );
  NAND2_X1 U15767 ( .A1(n14077), .A2(n9891), .ZN(n13746) );
  NAND2_X1 U15768 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  XNOR2_X1 U15769 ( .A(n13748), .B(n6549), .ZN(n13751) );
  AOI22_X1 U15770 ( .A1(n14369), .A2(n9891), .B1(n9892), .B2(n14077), .ZN(
        n13749) );
  XNOR2_X1 U15771 ( .A(n13751), .B(n13749), .ZN(n13780) );
  INV_X1 U15772 ( .A(n13749), .ZN(n13750) );
  NAND2_X1 U15773 ( .A1(n14198), .A2(n13798), .ZN(n13754) );
  NAND2_X1 U15774 ( .A1(n14079), .A2(n9891), .ZN(n13753) );
  NAND2_X1 U15775 ( .A1(n13754), .A2(n13753), .ZN(n13755) );
  XNOR2_X1 U15776 ( .A(n13755), .B(n6549), .ZN(n13756) );
  AOI22_X1 U15777 ( .A1(n14198), .A2(n9891), .B1(n9892), .B2(n14079), .ZN(
        n13757) );
  XNOR2_X1 U15778 ( .A(n13756), .B(n13757), .ZN(n13846) );
  INV_X1 U15779 ( .A(n13756), .ZN(n13758) );
  NAND2_X1 U15780 ( .A1(n14356), .A2(n13798), .ZN(n13760) );
  NAND2_X1 U15781 ( .A1(n14159), .A2(n9891), .ZN(n13759) );
  NAND2_X1 U15782 ( .A1(n13760), .A2(n13759), .ZN(n13761) );
  XNOR2_X1 U15783 ( .A(n13761), .B(n6549), .ZN(n13762) );
  AOI22_X1 U15784 ( .A1(n14356), .A2(n9891), .B1(n9892), .B2(n14159), .ZN(
        n13763) );
  XNOR2_X1 U15785 ( .A(n13762), .B(n13763), .ZN(n13819) );
  NAND2_X1 U15786 ( .A1(n13818), .A2(n13819), .ZN(n13766) );
  INV_X1 U15787 ( .A(n13762), .ZN(n13764) );
  NAND2_X1 U15788 ( .A1(n13764), .A2(n13763), .ZN(n13765) );
  NAND2_X1 U15789 ( .A1(n14347), .A2(n13798), .ZN(n13768) );
  NAND2_X1 U15790 ( .A1(n14101), .A2(n9891), .ZN(n13767) );
  NAND2_X1 U15791 ( .A1(n13768), .A2(n13767), .ZN(n13769) );
  XNOR2_X1 U15792 ( .A(n13769), .B(n6549), .ZN(n13770) );
  AOI22_X1 U15793 ( .A1(n14347), .A2(n9891), .B1(n9892), .B2(n14101), .ZN(
        n13771) );
  XNOR2_X1 U15794 ( .A(n13770), .B(n13771), .ZN(n13890) );
  INV_X1 U15795 ( .A(n13770), .ZN(n13772) );
  NAND2_X1 U15796 ( .A1(n13772), .A2(n13771), .ZN(n13773) );
  AOI22_X1 U15797 ( .A1(n14771), .A2(n14101), .B1(n14769), .B2(n14108), .ZN(
        n14142) );
  OAI22_X1 U15798 ( .A1(n13832), .A2(n14142), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13774), .ZN(n13775) );
  AOI21_X1 U15799 ( .B1(n14147), .B2(n13891), .A(n13775), .ZN(n13777) );
  NAND2_X1 U15800 ( .A1(n14343), .A2(n13905), .ZN(n13776) );
  OAI211_X1 U15801 ( .C1(n13778), .C2(n13908), .A(n13777), .B(n13776), .ZN(
        P1_U3214) );
  XOR2_X1 U15802 ( .A(n13780), .B(n13779), .Z(n13786) );
  NAND2_X1 U15803 ( .A1(n14074), .A2(n14771), .ZN(n13782) );
  NAND2_X1 U15804 ( .A1(n14769), .A2(n14079), .ZN(n13781) );
  NAND2_X1 U15805 ( .A1(n13782), .A2(n13781), .ZN(n14368) );
  AOI22_X1 U15806 ( .A1(n14368), .A2(n14733), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13783) );
  OAI21_X1 U15807 ( .B1(n14736), .B2(n14213), .A(n13783), .ZN(n13784) );
  AOI21_X1 U15808 ( .B1(n14369), .B2(n13905), .A(n13784), .ZN(n13785) );
  OAI21_X1 U15809 ( .B1(n13786), .B2(n13908), .A(n13785), .ZN(P1_U3216) );
  INV_X1 U15810 ( .A(n14392), .ZN(n14277) );
  AOI21_X1 U15811 ( .B1(n13788), .B2(n13787), .A(n13908), .ZN(n13790) );
  NAND2_X1 U15812 ( .A1(n13790), .A2(n13789), .ZN(n13793) );
  INV_X1 U15813 ( .A(n14313), .ZN(n14090) );
  OAI22_X1 U15814 ( .A1(n14239), .A2(n14240), .B1(n14090), .B2(n14288), .ZN(
        n14391) );
  AND2_X1 U15815 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14041) );
  NOR2_X1 U15816 ( .A1(n14736), .A2(n14272), .ZN(n13791) );
  AOI211_X1 U15817 ( .C1(n14733), .C2(n14391), .A(n14041), .B(n13791), .ZN(
        n13792) );
  OAI211_X1 U15818 ( .C1(n14277), .C2(n14659), .A(n13793), .B(n13792), .ZN(
        P1_U3219) );
  INV_X1 U15819 ( .A(n13794), .ZN(n13796) );
  AOI22_X1 U15820 ( .A1(n14338), .A2(n13798), .B1(n9891), .B2(n14108), .ZN(
        n13801) );
  AOI22_X1 U15821 ( .A1(n14338), .A2(n9891), .B1(n9892), .B2(n14108), .ZN(
        n13799) );
  XNOR2_X1 U15822 ( .A(n13799), .B(n6549), .ZN(n13800) );
  AOI22_X1 U15823 ( .A1(n13901), .A2(n14158), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13803) );
  NAND2_X1 U15824 ( .A1(n13891), .A2(n14132), .ZN(n13802) );
  OAI211_X1 U15825 ( .C1(n13804), .C2(n14660), .A(n13803), .B(n13802), .ZN(
        n13805) );
  AOI21_X1 U15826 ( .B1(n14338), .B2(n13905), .A(n13805), .ZN(n13806) );
  OAI21_X1 U15827 ( .B1(n13807), .B2(n13908), .A(n13806), .ZN(P1_U3220) );
  INV_X1 U15828 ( .A(n13808), .ZN(n13809) );
  AOI21_X1 U15829 ( .B1(n13811), .B2(n13810), .A(n13809), .ZN(n13817) );
  INV_X1 U15830 ( .A(n14074), .ZN(n14241) );
  OAI22_X1 U15831 ( .A1(n14241), .A2(n14660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13812), .ZN(n13813) );
  AOI21_X1 U15832 ( .B1(n13901), .B2(n14094), .A(n13813), .ZN(n13814) );
  OAI21_X1 U15833 ( .B1(n14736), .B2(n14242), .A(n13814), .ZN(n13815) );
  AOI21_X1 U15834 ( .B1(n14381), .B2(n13905), .A(n13815), .ZN(n13816) );
  OAI21_X1 U15835 ( .B1(n13817), .B2(n13908), .A(n13816), .ZN(P1_U3223) );
  XOR2_X1 U15836 ( .A(n13819), .B(n13818), .Z(n13826) );
  INV_X1 U15837 ( .A(n13820), .ZN(n14182) );
  NAND2_X1 U15838 ( .A1(n14771), .A2(n14079), .ZN(n13822) );
  NAND2_X1 U15839 ( .A1(n14769), .A2(n14101), .ZN(n13821) );
  NAND2_X1 U15840 ( .A1(n13822), .A2(n13821), .ZN(n14355) );
  AOI22_X1 U15841 ( .A1(n14733), .A2(n14355), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13823) );
  OAI21_X1 U15842 ( .B1(n14736), .B2(n14182), .A(n13823), .ZN(n13824) );
  AOI21_X1 U15843 ( .B1(n14356), .B2(n13905), .A(n13824), .ZN(n13825) );
  OAI21_X1 U15844 ( .B1(n13826), .B2(n13908), .A(n13825), .ZN(P1_U3225) );
  OAI21_X1 U15845 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n13830) );
  NAND2_X1 U15846 ( .A1(n13830), .A2(n14726), .ZN(n13836) );
  OAI21_X1 U15847 ( .B1(n13832), .B2(n14414), .A(n13831), .ZN(n13833) );
  AOI21_X1 U15848 ( .B1(n13834), .B2(n13891), .A(n13833), .ZN(n13835) );
  OAI211_X1 U15849 ( .C1(n14415), .C2(n14659), .A(n13836), .B(n13835), .ZN(
        P1_U3226) );
  NAND2_X1 U15850 ( .A1(n6672), .A2(n13837), .ZN(n13838) );
  XNOR2_X1 U15851 ( .A(n13839), .B(n13838), .ZN(n13844) );
  NAND2_X1 U15852 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14000)
         );
  OAI21_X1 U15853 ( .B1(n14660), .B2(n14090), .A(n14000), .ZN(n13840) );
  AOI21_X1 U15854 ( .B1(n13901), .B2(n14311), .A(n13840), .ZN(n13841) );
  OAI21_X1 U15855 ( .B1(n14736), .B2(n14314), .A(n13841), .ZN(n13842) );
  AOI21_X1 U15856 ( .B1(n14310), .B2(n13905), .A(n13842), .ZN(n13843) );
  OAI21_X1 U15857 ( .B1(n13844), .B2(n13908), .A(n13843), .ZN(P1_U3228) );
  XOR2_X1 U15858 ( .A(n13846), .B(n13845), .Z(n13852) );
  INV_X1 U15859 ( .A(n14159), .ZN(n14191) );
  AOI22_X1 U15860 ( .A1(n13901), .A2(n14077), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13847) );
  OAI21_X1 U15861 ( .B1(n14191), .B2(n14660), .A(n13847), .ZN(n13850) );
  NAND2_X1 U15862 ( .A1(n14198), .A2(n14722), .ZN(n14364) );
  NOR2_X1 U15863 ( .A1(n14364), .A2(n13848), .ZN(n13849) );
  AOI211_X1 U15864 ( .C1(n14197), .C2(n13891), .A(n13850), .B(n13849), .ZN(
        n13851) );
  OAI21_X1 U15865 ( .B1(n13852), .B2(n13908), .A(n13851), .ZN(P1_U3229) );
  OAI211_X1 U15866 ( .C1(n13855), .C2(n13854), .A(n13853), .B(n14726), .ZN(
        n13860) );
  NOR2_X1 U15867 ( .A1(n14736), .A2(n14258), .ZN(n13858) );
  INV_X1 U15868 ( .A(n14252), .ZN(n14225) );
  OAI22_X1 U15869 ( .A1(n14225), .A2(n14660), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13856), .ZN(n13857) );
  AOI211_X1 U15870 ( .C1(n13901), .C2(n14290), .A(n13858), .B(n13857), .ZN(
        n13859) );
  OAI211_X1 U15871 ( .C1(n14261), .C2(n14659), .A(n13860), .B(n13859), .ZN(
        P1_U3233) );
  XNOR2_X1 U15872 ( .A(n13861), .B(n13862), .ZN(n13872) );
  OAI22_X1 U15873 ( .A1(n14660), .A2(n13864), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13863), .ZN(n13867) );
  NOR2_X1 U15874 ( .A1(n14663), .A2(n13865), .ZN(n13866) );
  AOI211_X1 U15875 ( .C1(n13868), .C2(n13891), .A(n13867), .B(n13866), .ZN(
        n13871) );
  NAND2_X1 U15876 ( .A1(n13869), .A2(n13905), .ZN(n13870) );
  OAI211_X1 U15877 ( .C1(n13872), .C2(n13908), .A(n13871), .B(n13870), .ZN(
        P1_U3234) );
  OAI21_X1 U15878 ( .B1(n13875), .B2(n13874), .A(n13873), .ZN(n13876) );
  NAND2_X1 U15879 ( .A1(n13876), .A2(n14726), .ZN(n13881) );
  OAI22_X1 U15880 ( .A1(n14660), .A2(n14226), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13877), .ZN(n13879) );
  NOR2_X1 U15881 ( .A1(n14225), .A2(n14663), .ZN(n13878) );
  AOI211_X1 U15882 ( .C1(n14229), .C2(n13891), .A(n13879), .B(n13878), .ZN(
        n13880) );
  OAI211_X1 U15883 ( .C1(n14659), .C2(n14231), .A(n13881), .B(n13880), .ZN(
        P1_U3235) );
  XOR2_X1 U15884 ( .A(n13883), .B(n13882), .Z(n13888) );
  INV_X1 U15885 ( .A(n14290), .ZN(n14093) );
  NAND2_X1 U15886 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14015)
         );
  OAI21_X1 U15887 ( .B1(n14660), .B2(n14093), .A(n14015), .ZN(n13884) );
  AOI21_X1 U15888 ( .B1(n13901), .B2(n14088), .A(n13884), .ZN(n13885) );
  OAI21_X1 U15889 ( .B1(n14736), .B2(n14291), .A(n13885), .ZN(n13886) );
  AOI21_X1 U15890 ( .B1(n14398), .B2(n13905), .A(n13886), .ZN(n13887) );
  OAI21_X1 U15891 ( .B1(n13888), .B2(n13908), .A(n13887), .ZN(P1_U3238) );
  XOR2_X1 U15892 ( .A(n13890), .B(n13889), .Z(n13896) );
  AOI22_X1 U15893 ( .A1(n13901), .A2(n14159), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13893) );
  NAND2_X1 U15894 ( .A1(n13891), .A2(n14168), .ZN(n13892) );
  OAI211_X1 U15895 ( .C1(n14080), .C2(n14660), .A(n13893), .B(n13892), .ZN(
        n13894) );
  AOI21_X1 U15896 ( .B1(n14347), .B2(n13905), .A(n13894), .ZN(n13895) );
  OAI21_X1 U15897 ( .B1(n13896), .B2(n13908), .A(n13895), .ZN(P1_U3240) );
  XNOR2_X1 U15898 ( .A(n13897), .B(n13898), .ZN(n13909) );
  OAI21_X1 U15899 ( .B1(n14660), .B2(n14085), .A(n13899), .ZN(n13900) );
  AOI21_X1 U15900 ( .B1(n13901), .B2(n13911), .A(n13900), .ZN(n13902) );
  OAI21_X1 U15901 ( .B1(n14736), .B2(n13903), .A(n13902), .ZN(n13904) );
  AOI21_X1 U15902 ( .B1(n13906), .B2(n13905), .A(n13904), .ZN(n13907) );
  OAI21_X1 U15903 ( .B1(n13909), .B2(n13908), .A(n13907), .ZN(P1_U3241) );
  MUX2_X1 U15904 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14048), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U15905 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14110), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U15906 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14125), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15907 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14108), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U15908 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14158), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U15909 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14101), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15910 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14159), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U15911 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14079), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15912 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14074), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U15913 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14252), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15914 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14094), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15915 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14290), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15916 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14313), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15917 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14088), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15918 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14311), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15919 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n13910), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15920 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13911), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15921 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n13912), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U15922 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13913), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15923 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13914), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15924 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13915), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15925 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14768), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15926 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13916), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U15927 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14770), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U15928 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13917), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U15929 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13918), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15930 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13919), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U15931 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n13920), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U15932 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13921), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U15933 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n13922), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U15934 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9943), .S(P1_U4016), .Z(
        P1_U3560) );
  AND2_X1 U15935 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13924) );
  OAI211_X1 U15936 ( .C1(n13925), .C2(n13924), .A(n14748), .B(n13923), .ZN(
        n13934) );
  OAI22_X1 U15937 ( .A1(n14756), .A2(n7183), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13926), .ZN(n13927) );
  AOI21_X1 U15938 ( .B1(n14750), .B2(n13928), .A(n13927), .ZN(n13933) );
  OAI211_X1 U15939 ( .C1(n13931), .C2(n13930), .A(n14752), .B(n13929), .ZN(
        n13932) );
  NAND3_X1 U15940 ( .A1(n13934), .A2(n13933), .A3(n13932), .ZN(P1_U3244) );
  AND2_X1 U15941 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13937) );
  NOR2_X1 U15942 ( .A1(n13984), .A2(n13935), .ZN(n13936) );
  AOI211_X1 U15943 ( .C1(n13987), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13937), .B(
        n13936), .ZN(n13947) );
  OAI211_X1 U15944 ( .C1(n13940), .C2(n13939), .A(n14748), .B(n13938), .ZN(
        n13946) );
  AOI211_X1 U15945 ( .C1(n13943), .C2(n13942), .A(n13960), .B(n13941), .ZN(
        n13944) );
  INV_X1 U15946 ( .A(n13944), .ZN(n13945) );
  NAND3_X1 U15947 ( .A1(n13947), .A2(n13946), .A3(n13945), .ZN(P1_U3246) );
  NOR2_X1 U15948 ( .A1(n13984), .A2(n13948), .ZN(n13949) );
  AOI211_X1 U15949 ( .C1(n13987), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n13950), .B(
        n13949), .ZN(n13963) );
  OAI211_X1 U15950 ( .C1(n13953), .C2(n13952), .A(n14748), .B(n13951), .ZN(
        n13962) );
  MUX2_X1 U15951 ( .A(n10091), .B(P1_REG2_REG_4__SCAN_IN), .S(n13954), .Z(
        n13957) );
  INV_X1 U15952 ( .A(n13955), .ZN(n13956) );
  NAND2_X1 U15953 ( .A1(n13957), .A2(n13956), .ZN(n13959) );
  OAI211_X1 U15954 ( .C1(n13960), .C2(n13959), .A(n14752), .B(n13958), .ZN(
        n13961) );
  NAND4_X1 U15955 ( .A1(n13964), .A2(n13963), .A3(n13962), .A4(n13961), .ZN(
        P1_U3247) );
  NOR2_X1 U15956 ( .A1(n13984), .A2(n13965), .ZN(n13966) );
  AOI211_X1 U15957 ( .C1(n13987), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n13967), .B(
        n13966), .ZN(n13978) );
  OAI211_X1 U15958 ( .C1(n13970), .C2(n13969), .A(n14748), .B(n13968), .ZN(
        n13977) );
  OR3_X1 U15959 ( .A1(n13973), .A2(n13972), .A3(n13971), .ZN(n13974) );
  NAND3_X1 U15960 ( .A1(n14752), .A2(n13975), .A3(n13974), .ZN(n13976) );
  NAND3_X1 U15961 ( .A1(n13978), .A2(n13977), .A3(n13976), .ZN(P1_U3249) );
  OAI211_X1 U15962 ( .C1(n13981), .C2(n13980), .A(n13979), .B(n14748), .ZN(
        n13995) );
  INV_X1 U15963 ( .A(n13982), .ZN(n13986) );
  NOR2_X1 U15964 ( .A1(n13984), .A2(n13983), .ZN(n13985) );
  AOI211_X1 U15965 ( .C1(n13987), .C2(P1_ADDR_REG_10__SCAN_IN), .A(n13986), 
        .B(n13985), .ZN(n13994) );
  OR3_X1 U15966 ( .A1(n13990), .A2(n13989), .A3(n13988), .ZN(n13991) );
  NAND3_X1 U15967 ( .A1(n13992), .A2(n14752), .A3(n13991), .ZN(n13993) );
  NAND3_X1 U15968 ( .A1(n13995), .A2(n13994), .A3(n13993), .ZN(P1_U3253) );
  XNOR2_X1 U15969 ( .A(n14012), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13997) );
  AOI211_X1 U15970 ( .C1(n13998), .C2(n13997), .A(n14011), .B(n14036), .ZN(
        n13999) );
  INV_X1 U15971 ( .A(n13999), .ZN(n14010) );
  INV_X1 U15972 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14001) );
  OAI21_X1 U15973 ( .B1(n14756), .B2(n14001), .A(n14000), .ZN(n14002) );
  AOI21_X1 U15974 ( .B1(n14750), .B2(n14012), .A(n14002), .ZN(n14009) );
  XNOR2_X1 U15975 ( .A(n14012), .B(n14319), .ZN(n14007) );
  INV_X1 U15976 ( .A(n14003), .ZN(n14005) );
  OAI21_X1 U15977 ( .B1(n14005), .B2(n11324), .A(n14004), .ZN(n14006) );
  NAND2_X1 U15978 ( .A1(n14007), .A2(n14006), .ZN(n14018) );
  OAI211_X1 U15979 ( .C1(n14007), .C2(n14006), .A(n14752), .B(n14018), .ZN(
        n14008) );
  NAND3_X1 U15980 ( .A1(n14010), .A2(n14009), .A3(n14008), .ZN(P1_U3260) );
  INV_X1 U15981 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14405) );
  NOR2_X1 U15982 ( .A1(n14405), .A2(n14013), .ZN(n14027) );
  AOI211_X1 U15983 ( .C1(n14013), .C2(n14405), .A(n14027), .B(n14036), .ZN(
        n14014) );
  INV_X1 U15984 ( .A(n14014), .ZN(n14023) );
  INV_X1 U15985 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14016) );
  OAI21_X1 U15986 ( .B1(n14756), .B2(n14016), .A(n14015), .ZN(n14017) );
  AOI21_X1 U15987 ( .B1(n14750), .B2(n14031), .A(n14017), .ZN(n14022) );
  OAI21_X1 U15988 ( .B1(n14319), .B2(n14019), .A(n14018), .ZN(n14030) );
  XNOR2_X1 U15989 ( .A(n14024), .B(n14030), .ZN(n14020) );
  NAND2_X1 U15990 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n14020), .ZN(n14033) );
  OAI211_X1 U15991 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n14020), .A(n14752), 
        .B(n14033), .ZN(n14021) );
  NAND3_X1 U15992 ( .A1(n14023), .A2(n14022), .A3(n14021), .ZN(P1_U3261) );
  NOR2_X1 U15993 ( .A1(n14025), .A2(n14024), .ZN(n14026) );
  NOR2_X1 U15994 ( .A1(n14027), .A2(n14026), .ZN(n14029) );
  INV_X1 U15995 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14028) );
  XOR2_X1 U15996 ( .A(n14029), .B(n14028), .Z(n14037) );
  NAND2_X1 U15997 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  NAND2_X1 U15998 ( .A1(n14033), .A2(n14032), .ZN(n14034) );
  XOR2_X1 U15999 ( .A(n14034), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14035) );
  AOI22_X1 U16000 ( .A1(n14037), .A2(n14748), .B1(n14752), .B2(n14035), .ZN(
        n14040) );
  INV_X1 U16001 ( .A(n14035), .ZN(n14038) );
  INV_X1 U16002 ( .A(n14041), .ZN(n14042) );
  INV_X1 U16003 ( .A(n14310), .ZN(n14409) );
  OR2_X2 U16004 ( .A1(n14398), .A2(n14306), .ZN(n14293) );
  NAND2_X1 U16005 ( .A1(n14271), .A2(n14261), .ZN(n14255) );
  NOR2_X2 U16006 ( .A1(n14044), .A2(n14107), .ZN(n14052) );
  XNOR2_X1 U16007 ( .A(n14052), .B(n14049), .ZN(n14045) );
  NAND2_X1 U16008 ( .A1(n14045), .A2(n14812), .ZN(n14324) );
  INV_X1 U16009 ( .A(P1_B_REG_SCAN_IN), .ZN(n14046) );
  NOR2_X1 U16010 ( .A1(n14454), .A2(n14046), .ZN(n14047) );
  NOR2_X1 U16011 ( .A1(n14240), .A2(n14047), .ZN(n14109) );
  NAND2_X1 U16012 ( .A1(n14109), .A2(n14048), .ZN(n14326) );
  NOR2_X1 U16013 ( .A1(n14833), .A2(n14326), .ZN(n14055) );
  NOR2_X1 U16014 ( .A1(n14325), .A2(n14808), .ZN(n14050) );
  AOI211_X1 U16015 ( .C1(n14315), .C2(P1_REG2_REG_31__SCAN_IN), .A(n14055), 
        .B(n14050), .ZN(n14051) );
  OAI21_X1 U16016 ( .B1(n14324), .B2(n14308), .A(n14051), .ZN(P1_U3263) );
  INV_X1 U16017 ( .A(n14107), .ZN(n14054) );
  INV_X1 U16018 ( .A(n14052), .ZN(n14053) );
  OAI211_X1 U16019 ( .C1(n14328), .C2(n14054), .A(n14053), .B(n14812), .ZN(
        n14327) );
  NAND2_X1 U16020 ( .A1(n14315), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14057) );
  INV_X1 U16021 ( .A(n14055), .ZN(n14056) );
  OAI211_X1 U16022 ( .C1(n14328), .C2(n14808), .A(n14057), .B(n14056), .ZN(
        n14058) );
  INV_X1 U16023 ( .A(n14058), .ZN(n14059) );
  OAI21_X1 U16024 ( .B1(n14327), .B2(n14308), .A(n14059), .ZN(P1_U3264) );
  INV_X1 U16025 ( .A(n14343), .ZN(n14149) );
  INV_X1 U16026 ( .A(n14101), .ZN(n14102) );
  NAND2_X1 U16027 ( .A1(n14060), .A2(n14083), .ZN(n14062) );
  OR2_X1 U16028 ( .A1(n14086), .A2(n14311), .ZN(n14061) );
  INV_X1 U16029 ( .A(n14063), .ZN(n14064) );
  INV_X1 U16030 ( .A(n14066), .ZN(n14068) );
  NAND2_X1 U16031 ( .A1(n14267), .A2(n14269), .ZN(n14070) );
  OR2_X1 U16032 ( .A1(n14392), .A2(n14290), .ZN(n14069) );
  OR2_X1 U16033 ( .A1(n14261), .A2(n14239), .ZN(n14072) );
  NAND2_X1 U16034 ( .A1(n14219), .A2(n14222), .ZN(n14076) );
  OR2_X1 U16035 ( .A1(n14375), .A2(n14074), .ZN(n14075) );
  NAND2_X1 U16036 ( .A1(n14076), .A2(n14075), .ZN(n14203) );
  INV_X1 U16037 ( .A(n14204), .ZN(n14207) );
  NAND2_X1 U16038 ( .A1(n14369), .A2(n14077), .ZN(n14078) );
  INV_X1 U16039 ( .A(n14156), .ZN(n14163) );
  INV_X1 U16040 ( .A(n14123), .ZN(n14121) );
  NAND2_X1 U16041 ( .A1(n14086), .A2(n14085), .ZN(n14087) );
  INV_X1 U16042 ( .A(n14300), .ZN(n14305) );
  INV_X1 U16043 ( .A(n14088), .ZN(n14289) );
  OR2_X1 U16044 ( .A1(n14310), .A2(n14289), .ZN(n14089) );
  NAND2_X1 U16045 ( .A1(n14302), .A2(n14089), .ZN(n14283) );
  NAND2_X1 U16046 ( .A1(n14283), .A2(n14281), .ZN(n14092) );
  OR2_X1 U16047 ( .A1(n14398), .A2(n14090), .ZN(n14091) );
  NAND2_X1 U16048 ( .A1(n14261), .A2(n14094), .ZN(n14095) );
  NOR2_X1 U16049 ( .A1(n14381), .A2(n14225), .ZN(n14096) );
  INV_X1 U16050 ( .A(n14222), .ZN(n14221) );
  NAND2_X1 U16051 ( .A1(n14369), .A2(n14226), .ZN(n14097) );
  OR2_X1 U16052 ( .A1(n14198), .A2(n14098), .ZN(n14099) );
  NAND2_X1 U16053 ( .A1(n14356), .A2(n14191), .ZN(n14100) );
  INV_X1 U16054 ( .A(n14108), .ZN(n14103) );
  AOI22_X1 U16055 ( .A1(n14124), .A2(n14123), .B1(n14103), .B2(n14338), .ZN(
        n14105) );
  XNOR2_X1 U16056 ( .A(n14105), .B(n14104), .ZN(n14336) );
  OR2_X1 U16057 ( .A1(n14333), .A2(n14135), .ZN(n14106) );
  AND3_X1 U16058 ( .A1(n14107), .A2(n14812), .A3(n14106), .ZN(n14330) );
  NAND2_X1 U16059 ( .A1(n14330), .A2(n14818), .ZN(n14117) );
  NAND2_X1 U16060 ( .A1(n14771), .A2(n14108), .ZN(n14331) );
  NOR2_X1 U16061 ( .A1(n14315), .A2(n14331), .ZN(n14115) );
  NAND2_X1 U16062 ( .A1(n14110), .A2(n14109), .ZN(n14332) );
  INV_X1 U16063 ( .A(n14111), .ZN(n14112) );
  OAI22_X1 U16064 ( .A1(n14332), .A2(n14113), .B1(n14112), .B2(n14775), .ZN(
        n14114) );
  AOI211_X1 U16065 ( .C1(n14315), .C2(P1_REG2_REG_29__SCAN_IN), .A(n14115), 
        .B(n14114), .ZN(n14116) );
  OAI211_X1 U16066 ( .C1(n14333), .C2(n14808), .A(n14117), .B(n14116), .ZN(
        n14118) );
  AOI21_X1 U16067 ( .B1(n14336), .B2(n14829), .A(n14118), .ZN(n14119) );
  OAI21_X1 U16068 ( .B1(n14329), .B2(n14323), .A(n14119), .ZN(P1_U3356) );
  OAI21_X1 U16069 ( .B1(n14122), .B2(n14121), .A(n14120), .ZN(n14341) );
  XNOR2_X1 U16070 ( .A(n14124), .B(n14123), .ZN(n14129) );
  NAND2_X1 U16071 ( .A1(n14125), .A2(n14769), .ZN(n14127) );
  NAND2_X1 U16072 ( .A1(n14158), .A2(n14771), .ZN(n14126) );
  OAI21_X1 U16073 ( .B1(n14130), .B2(n14341), .A(n14340), .ZN(n14131) );
  NAND2_X1 U16074 ( .A1(n14131), .A2(n14774), .ZN(n14139) );
  AOI22_X1 U16075 ( .A1(n14833), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n14132), 
        .B2(n14826), .ZN(n14138) );
  NAND2_X1 U16076 ( .A1(n14338), .A2(n14145), .ZN(n14133) );
  NAND2_X1 U16077 ( .A1(n14133), .A2(n14812), .ZN(n14134) );
  NOR2_X1 U16078 ( .A1(n14135), .A2(n14134), .ZN(n14337) );
  NAND2_X1 U16079 ( .A1(n14337), .A2(n14818), .ZN(n14137) );
  NAND2_X1 U16080 ( .A1(n14338), .A2(n14309), .ZN(n14136) );
  NAND4_X1 U16081 ( .A1(n14139), .A2(n14138), .A3(n14137), .A4(n14136), .ZN(
        P1_U3265) );
  XNOR2_X1 U16082 ( .A(n14141), .B(n14140), .ZN(n14144) );
  INV_X1 U16083 ( .A(n14142), .ZN(n14143) );
  AOI21_X1 U16084 ( .B1(n14144), .B2(n14766), .A(n14143), .ZN(n14345) );
  INV_X1 U16085 ( .A(n14145), .ZN(n14146) );
  AOI211_X1 U16086 ( .C1(n14343), .C2(n14166), .A(n14292), .B(n14146), .ZN(
        n14342) );
  AOI22_X1 U16087 ( .A1(n14315), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n14147), 
        .B2(n14826), .ZN(n14148) );
  OAI21_X1 U16088 ( .B1(n14149), .B2(n14808), .A(n14148), .ZN(n14153) );
  AOI21_X1 U16089 ( .B1(n9555), .B2(n14151), .A(n14150), .ZN(n14346) );
  NOR2_X1 U16090 ( .A1(n14346), .A2(n14323), .ZN(n14152) );
  AOI211_X1 U16091 ( .C1(n14342), .C2(n14818), .A(n14153), .B(n14152), .ZN(
        n14154) );
  OAI21_X1 U16092 ( .B1(n14315), .B2(n14345), .A(n14154), .ZN(P1_U3266) );
  XNOR2_X1 U16093 ( .A(n14155), .B(n14156), .ZN(n14157) );
  NAND2_X1 U16094 ( .A1(n14157), .A2(n14766), .ZN(n14161) );
  AOI22_X1 U16095 ( .A1(n14771), .A2(n14159), .B1(n14769), .B2(n14158), .ZN(
        n14160) );
  OR2_X1 U16096 ( .A1(n14163), .A2(n14162), .ZN(n14165) );
  OAI211_X1 U16097 ( .C1(n14167), .C2(n14181), .A(n14812), .B(n14166), .ZN(
        n14349) );
  AOI22_X1 U16098 ( .A1(n14833), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n14168), 
        .B2(n14826), .ZN(n14170) );
  NAND2_X1 U16099 ( .A1(n14347), .A2(n14309), .ZN(n14169) );
  OAI211_X1 U16100 ( .C1(n14349), .C2(n14308), .A(n14170), .B(n14169), .ZN(
        n14171) );
  AOI21_X1 U16101 ( .B1(n14351), .B2(n14828), .A(n14171), .ZN(n14172) );
  OAI21_X1 U16102 ( .B1(n14353), .B2(n14315), .A(n14172), .ZN(P1_U3267) );
  OAI21_X1 U16103 ( .B1(n14175), .B2(n14174), .A(n14173), .ZN(n14360) );
  INV_X1 U16104 ( .A(n14176), .ZN(n14178) );
  OAI21_X1 U16105 ( .B1(n14178), .B2(n14177), .A(n6651), .ZN(n14357) );
  NAND2_X1 U16106 ( .A1(n14357), .A2(n14829), .ZN(n14189) );
  NAND2_X1 U16107 ( .A1(n14356), .A2(n14196), .ZN(n14179) );
  NAND2_X1 U16108 ( .A1(n14179), .A2(n14812), .ZN(n14180) );
  NOR2_X1 U16109 ( .A1(n14181), .A2(n14180), .ZN(n14354) );
  INV_X1 U16110 ( .A(n14356), .ZN(n14186) );
  INV_X1 U16111 ( .A(n14355), .ZN(n14183) );
  OAI22_X1 U16112 ( .A1(n14315), .A2(n14183), .B1(n14182), .B2(n14775), .ZN(
        n14184) );
  AOI21_X1 U16113 ( .B1(P1_REG2_REG_25__SCAN_IN), .B2(n14315), .A(n14184), 
        .ZN(n14185) );
  OAI21_X1 U16114 ( .B1(n14186), .B2(n14808), .A(n14185), .ZN(n14187) );
  AOI21_X1 U16115 ( .B1(n14354), .B2(n14818), .A(n14187), .ZN(n14188) );
  OAI211_X1 U16116 ( .C1(n14360), .C2(n14323), .A(n14189), .B(n14188), .ZN(
        P1_U3268) );
  XNOR2_X1 U16117 ( .A(n14190), .B(n14193), .ZN(n14361) );
  OAI22_X1 U16118 ( .A1(n14226), .A2(n14288), .B1(n14191), .B2(n14240), .ZN(
        n14195) );
  AOI211_X1 U16119 ( .C1(n14193), .C2(n14192), .A(n14802), .B(n6952), .ZN(
        n14194) );
  OAI211_X1 U16120 ( .C1(n6959), .C2(n6960), .A(n14812), .B(n14196), .ZN(
        n14362) );
  AOI22_X1 U16121 ( .A1(n14833), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14826), 
        .B2(n14197), .ZN(n14200) );
  NAND2_X1 U16122 ( .A1(n14198), .A2(n14309), .ZN(n14199) );
  OAI211_X1 U16123 ( .C1(n14362), .C2(n14308), .A(n14200), .B(n14199), .ZN(
        n14201) );
  AOI21_X1 U16124 ( .B1(n14816), .B2(n14361), .A(n14201), .ZN(n14202) );
  OAI21_X1 U16125 ( .B1(n14365), .B2(n14833), .A(n14202), .ZN(P1_U3269) );
  INV_X1 U16126 ( .A(n14203), .ZN(n14205) );
  OAI21_X1 U16127 ( .B1(n14205), .B2(n14204), .A(n6576), .ZN(n14372) );
  OAI21_X1 U16128 ( .B1(n14208), .B2(n14207), .A(n14206), .ZN(n14366) );
  AOI21_X1 U16129 ( .B1(n14369), .B2(n14227), .A(n14292), .ZN(n14210) );
  AND2_X1 U16130 ( .A1(n14210), .A2(n14209), .ZN(n14367) );
  NAND2_X1 U16131 ( .A1(n14367), .A2(n14818), .ZN(n14216) );
  NAND2_X1 U16132 ( .A1(n14368), .A2(n14774), .ZN(n14212) );
  NAND2_X1 U16133 ( .A1(n14315), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n14211) );
  OAI211_X1 U16134 ( .C1(n14775), .C2(n14213), .A(n14212), .B(n14211), .ZN(
        n14214) );
  AOI21_X1 U16135 ( .B1(n14369), .B2(n14309), .A(n14214), .ZN(n14215) );
  NAND2_X1 U16136 ( .A1(n14216), .A2(n14215), .ZN(n14217) );
  AOI21_X1 U16137 ( .B1(n14366), .B2(n14829), .A(n14217), .ZN(n14218) );
  OAI21_X1 U16138 ( .B1(n14323), .B2(n14372), .A(n14218), .ZN(P1_U3270) );
  XNOR2_X1 U16139 ( .A(n14220), .B(n14221), .ZN(n14377) );
  XNOR2_X1 U16140 ( .A(n14223), .B(n14222), .ZN(n14224) );
  OAI222_X1 U16141 ( .A1(n14240), .A2(n14226), .B1(n14288), .B2(n14225), .C1(
        n14802), .C2(n14224), .ZN(n14373) );
  NAND2_X1 U16142 ( .A1(n14373), .A2(n14774), .ZN(n14234) );
  INV_X1 U16143 ( .A(n14227), .ZN(n14228) );
  AOI211_X1 U16144 ( .C1(n14375), .C2(n14238), .A(n14292), .B(n14228), .ZN(
        n14374) );
  AOI22_X1 U16145 ( .A1(n14833), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14229), 
        .B2(n14826), .ZN(n14230) );
  OAI21_X1 U16146 ( .B1(n14231), .B2(n14808), .A(n14230), .ZN(n14232) );
  AOI21_X1 U16147 ( .B1(n14374), .B2(n14818), .A(n14232), .ZN(n14233) );
  OAI211_X1 U16148 ( .C1(n14377), .C2(n14323), .A(n14234), .B(n14233), .ZN(
        P1_U3271) );
  AOI21_X1 U16149 ( .B1(n14236), .B2(n14235), .A(n6612), .ZN(n14384) );
  XOR2_X1 U16150 ( .A(n14237), .B(n14236), .Z(n14378) );
  NAND2_X1 U16151 ( .A1(n14378), .A2(n14829), .ZN(n14249) );
  AOI211_X1 U16152 ( .C1(n14381), .C2(n14255), .A(n14292), .B(n6961), .ZN(
        n14379) );
  INV_X1 U16153 ( .A(n14381), .ZN(n14246) );
  OAI22_X1 U16154 ( .A1(n14241), .A2(n14240), .B1(n14239), .B2(n14288), .ZN(
        n14380) );
  INV_X1 U16155 ( .A(n14242), .ZN(n14243) );
  AOI22_X1 U16156 ( .A1(n14380), .A2(n14774), .B1(n14243), .B2(n14826), .ZN(
        n14245) );
  NAND2_X1 U16157 ( .A1(n14315), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n14244) );
  OAI211_X1 U16158 ( .C1(n14246), .C2(n14808), .A(n14245), .B(n14244), .ZN(
        n14247) );
  AOI21_X1 U16159 ( .B1(n14379), .B2(n14818), .A(n14247), .ZN(n14248) );
  OAI211_X1 U16160 ( .C1(n14384), .C2(n14323), .A(n14249), .B(n14248), .ZN(
        P1_U3272) );
  OAI211_X1 U16161 ( .C1(n14251), .C2(n14262), .A(n6721), .B(n14766), .ZN(
        n14254) );
  AOI22_X1 U16162 ( .A1(n14252), .A2(n14769), .B1(n14771), .B2(n14290), .ZN(
        n14253) );
  AND2_X1 U16163 ( .A1(n14254), .A2(n14253), .ZN(n14388) );
  INV_X1 U16164 ( .A(n14271), .ZN(n14257) );
  INV_X1 U16165 ( .A(n14255), .ZN(n14256) );
  AOI211_X1 U16166 ( .C1(n14386), .C2(n14257), .A(n14292), .B(n14256), .ZN(
        n14385) );
  INV_X1 U16167 ( .A(n14258), .ZN(n14259) );
  AOI22_X1 U16168 ( .A1(n14315), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n14259), 
        .B2(n14826), .ZN(n14260) );
  OAI21_X1 U16169 ( .B1(n14261), .B2(n14808), .A(n14260), .ZN(n14265) );
  OAI21_X1 U16170 ( .B1(n6542), .B2(n14071), .A(n14263), .ZN(n14389) );
  NOR2_X1 U16171 ( .A1(n14389), .A2(n14323), .ZN(n14264) );
  AOI211_X1 U16172 ( .C1(n14385), .C2(n14818), .A(n14265), .B(n14264), .ZN(
        n14266) );
  OAI21_X1 U16173 ( .B1(n14315), .B2(n14388), .A(n14266), .ZN(P1_U3273) );
  XNOR2_X1 U16174 ( .A(n14267), .B(n14268), .ZN(n14396) );
  XNOR2_X1 U16175 ( .A(n14270), .B(n14269), .ZN(n14393) );
  AOI211_X1 U16176 ( .C1(n14392), .C2(n14293), .A(n14292), .B(n14271), .ZN(
        n14390) );
  NAND2_X1 U16177 ( .A1(n14390), .A2(n14818), .ZN(n14276) );
  INV_X1 U16178 ( .A(n14391), .ZN(n14273) );
  OAI22_X1 U16179 ( .A1(n14273), .A2(n14315), .B1(n14272), .B2(n14775), .ZN(
        n14274) );
  AOI21_X1 U16180 ( .B1(P1_REG2_REG_19__SCAN_IN), .B2(n14315), .A(n14274), 
        .ZN(n14275) );
  OAI211_X1 U16181 ( .C1(n14277), .C2(n14808), .A(n14276), .B(n14275), .ZN(
        n14278) );
  AOI21_X1 U16182 ( .B1(n14393), .B2(n14829), .A(n14278), .ZN(n14279) );
  OAI21_X1 U16183 ( .B1(n14323), .B2(n14396), .A(n14279), .ZN(P1_U3274) );
  XNOR2_X1 U16184 ( .A(n14280), .B(n14281), .ZN(n14285) );
  INV_X1 U16185 ( .A(n14285), .ZN(n14402) );
  INV_X1 U16186 ( .A(n14281), .ZN(n14282) );
  XNOR2_X1 U16187 ( .A(n14283), .B(n14282), .ZN(n14284) );
  NAND2_X1 U16188 ( .A1(n14284), .A2(n14766), .ZN(n14287) );
  NAND2_X1 U16189 ( .A1(n14285), .A2(n14899), .ZN(n14286) );
  OAI211_X1 U16190 ( .C1(n14289), .C2(n14288), .A(n14287), .B(n14286), .ZN(
        n14404) );
  AND2_X1 U16191 ( .A1(n14290), .A2(n14769), .ZN(n14397) );
  OAI21_X1 U16192 ( .B1(n14404), .B2(n14397), .A(n14774), .ZN(n14298) );
  OAI22_X1 U16193 ( .A1(n14774), .A2(n13515), .B1(n14291), .B2(n14775), .ZN(
        n14296) );
  AOI21_X1 U16194 ( .B1(n14398), .B2(n14306), .A(n14292), .ZN(n14294) );
  NAND2_X1 U16195 ( .A1(n14294), .A2(n14293), .ZN(n14399) );
  NOR2_X1 U16196 ( .A1(n14399), .A2(n14308), .ZN(n14295) );
  AOI211_X1 U16197 ( .C1(n14309), .C2(n14398), .A(n14296), .B(n14295), .ZN(
        n14297) );
  OAI211_X1 U16198 ( .C1(n14402), .C2(n14299), .A(n14298), .B(n14297), .ZN(
        P1_U3275) );
  XNOR2_X1 U16199 ( .A(n14301), .B(n14300), .ZN(n14413) );
  INV_X1 U16200 ( .A(n14302), .ZN(n14303) );
  AOI21_X1 U16201 ( .B1(n14305), .B2(n14304), .A(n14303), .ZN(n14411) );
  OAI211_X1 U16202 ( .C1(n14307), .C2(n14409), .A(n14812), .B(n14306), .ZN(
        n14408) );
  NOR2_X1 U16203 ( .A1(n14408), .A2(n14308), .ZN(n14321) );
  NAND2_X1 U16204 ( .A1(n14310), .A2(n14309), .ZN(n14318) );
  AND2_X1 U16205 ( .A1(n14771), .A2(n14311), .ZN(n14312) );
  AOI21_X1 U16206 ( .B1(n14313), .B2(n14769), .A(n14312), .ZN(n14407) );
  OAI22_X1 U16207 ( .A1(n14315), .A2(n14407), .B1(n14314), .B2(n14775), .ZN(
        n14316) );
  INV_X1 U16208 ( .A(n14316), .ZN(n14317) );
  OAI211_X1 U16209 ( .C1(n14774), .C2(n14319), .A(n14318), .B(n14317), .ZN(
        n14320) );
  AOI211_X1 U16210 ( .C1(n14411), .C2(n14829), .A(n14321), .B(n14320), .ZN(
        n14322) );
  OAI21_X1 U16211 ( .B1(n14323), .B2(n14413), .A(n14322), .ZN(P1_U3276) );
  OAI211_X1 U16212 ( .C1(n14325), .C2(n14920), .A(n14324), .B(n14326), .ZN(
        n14423) );
  MUX2_X1 U16213 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14423), .S(n14940), .Z(
        P1_U3559) );
  OAI211_X1 U16214 ( .C1(n14328), .C2(n14920), .A(n14327), .B(n14326), .ZN(
        n14424) );
  MUX2_X1 U16215 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14424), .S(n14940), .Z(
        P1_U3558) );
  OAI211_X1 U16216 ( .C1(n14333), .C2(n14920), .A(n14332), .B(n14331), .ZN(
        n14334) );
  MUX2_X1 U16217 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14425), .S(n14940), .Z(
        P1_U3557) );
  AOI21_X1 U16218 ( .B1(n14722), .B2(n14338), .A(n14337), .ZN(n14339) );
  OAI211_X1 U16219 ( .C1(n14420), .C2(n14341), .A(n14340), .B(n14339), .ZN(
        n14426) );
  MUX2_X1 U16220 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14426), .S(n14940), .Z(
        P1_U3556) );
  AOI21_X1 U16221 ( .B1(n14722), .B2(n14343), .A(n14342), .ZN(n14344) );
  OAI211_X1 U16222 ( .C1(n14346), .C2(n14420), .A(n14345), .B(n14344), .ZN(
        n14427) );
  MUX2_X1 U16223 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14427), .S(n14940), .Z(
        P1_U3555) );
  NAND2_X1 U16224 ( .A1(n14347), .A2(n14722), .ZN(n14348) );
  NAND2_X1 U16225 ( .A1(n14349), .A2(n14348), .ZN(n14350) );
  AOI21_X1 U16226 ( .B1(n14351), .B2(n14922), .A(n14350), .ZN(n14352) );
  NAND2_X1 U16227 ( .A1(n14353), .A2(n14352), .ZN(n14428) );
  MUX2_X1 U16228 ( .A(n14428), .B(P1_REG1_REG_26__SCAN_IN), .S(n14937), .Z(
        P1_U3554) );
  AOI211_X1 U16229 ( .C1(n14722), .C2(n14356), .A(n14355), .B(n14354), .ZN(
        n14359) );
  NAND2_X1 U16230 ( .A1(n14357), .A2(n14766), .ZN(n14358) );
  OAI211_X1 U16231 ( .C1(n14420), .C2(n14360), .A(n14359), .B(n14358), .ZN(
        n14429) );
  MUX2_X1 U16232 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14429), .S(n14940), .Z(
        P1_U3553) );
  NAND2_X1 U16233 ( .A1(n14361), .A2(n14916), .ZN(n14363) );
  NAND4_X1 U16234 ( .A1(n14365), .A2(n14364), .A3(n14363), .A4(n14362), .ZN(
        n14430) );
  MUX2_X1 U16235 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14430), .S(n14940), .Z(
        P1_U3552) );
  NAND2_X1 U16236 ( .A1(n14366), .A2(n14766), .ZN(n14371) );
  AOI211_X1 U16237 ( .C1(n14722), .C2(n14369), .A(n14368), .B(n14367), .ZN(
        n14370) );
  OAI211_X1 U16238 ( .C1(n14372), .C2(n14420), .A(n14371), .B(n14370), .ZN(
        n14431) );
  MUX2_X1 U16239 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14431), .S(n14940), .Z(
        P1_U3551) );
  AOI211_X1 U16240 ( .C1(n14722), .C2(n14375), .A(n14374), .B(n14373), .ZN(
        n14376) );
  OAI21_X1 U16241 ( .B1(n14420), .B2(n14377), .A(n14376), .ZN(n14432) );
  MUX2_X1 U16242 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14432), .S(n14940), .Z(
        P1_U3550) );
  NAND2_X1 U16243 ( .A1(n14378), .A2(n14766), .ZN(n14383) );
  AOI211_X1 U16244 ( .C1(n14722), .C2(n14381), .A(n14380), .B(n14379), .ZN(
        n14382) );
  OAI211_X1 U16245 ( .C1(n14384), .C2(n14420), .A(n14383), .B(n14382), .ZN(
        n14433) );
  MUX2_X1 U16246 ( .A(n14433), .B(P1_REG1_REG_21__SCAN_IN), .S(n14937), .Z(
        P1_U3549) );
  AOI21_X1 U16247 ( .B1(n14722), .B2(n14386), .A(n14385), .ZN(n14387) );
  OAI211_X1 U16248 ( .C1(n14420), .C2(n14389), .A(n14388), .B(n14387), .ZN(
        n14434) );
  MUX2_X1 U16249 ( .A(n14434), .B(P1_REG1_REG_20__SCAN_IN), .S(n14937), .Z(
        P1_U3548) );
  AOI211_X1 U16250 ( .C1(n14722), .C2(n14392), .A(n14391), .B(n14390), .ZN(
        n14395) );
  NAND2_X1 U16251 ( .A1(n14393), .A2(n14766), .ZN(n14394) );
  OAI211_X1 U16252 ( .C1(n14420), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        n14435) );
  MUX2_X1 U16253 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n14435), .S(n14940), .Z(
        P1_U3547) );
  AOI21_X1 U16254 ( .B1(n14398), .B2(n14722), .A(n14397), .ZN(n14400) );
  OAI211_X1 U16255 ( .C1(n14402), .C2(n14401), .A(n14400), .B(n14399), .ZN(
        n14403) );
  NOR2_X1 U16256 ( .A1(n14404), .A2(n14403), .ZN(n14436) );
  MUX2_X1 U16257 ( .A(n14405), .B(n14436), .S(n14940), .Z(n14406) );
  INV_X1 U16258 ( .A(n14406), .ZN(P1_U3546) );
  OAI211_X1 U16259 ( .C1(n14409), .C2(n14920), .A(n14408), .B(n14407), .ZN(
        n14410) );
  AOI21_X1 U16260 ( .B1(n14411), .B2(n14766), .A(n14410), .ZN(n14412) );
  OAI21_X1 U16261 ( .B1(n14420), .B2(n14413), .A(n14412), .ZN(n14439) );
  MUX2_X1 U16262 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14439), .S(n14940), .Z(
        P1_U3545) );
  OAI21_X1 U16263 ( .B1(n14415), .B2(n14920), .A(n14414), .ZN(n14416) );
  AOI211_X1 U16264 ( .C1(n14418), .C2(n14766), .A(n14417), .B(n14416), .ZN(
        n14419) );
  OAI21_X1 U16265 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14440) );
  MUX2_X1 U16266 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14440), .S(n14940), .Z(
        P1_U3544) );
  MUX2_X1 U16267 ( .A(n14422), .B(P1_REG1_REG_0__SCAN_IN), .S(n14937), .Z(
        P1_U3528) );
  MUX2_X1 U16268 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14423), .S(n14925), .Z(
        P1_U3527) );
  MUX2_X1 U16269 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14424), .S(n14925), .Z(
        P1_U3526) );
  MUX2_X1 U16270 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14425), .S(n14925), .Z(
        P1_U3525) );
  MUX2_X1 U16271 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14426), .S(n14925), .Z(
        P1_U3524) );
  MUX2_X1 U16272 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14427), .S(n14925), .Z(
        P1_U3523) );
  MUX2_X1 U16273 ( .A(n14428), .B(P1_REG0_REG_26__SCAN_IN), .S(n14924), .Z(
        P1_U3522) );
  MUX2_X1 U16274 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14429), .S(n14925), .Z(
        P1_U3521) );
  MUX2_X1 U16275 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14430), .S(n14925), .Z(
        P1_U3520) );
  MUX2_X1 U16276 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14431), .S(n14925), .Z(
        P1_U3519) );
  MUX2_X1 U16277 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14432), .S(n14925), .Z(
        P1_U3518) );
  MUX2_X1 U16278 ( .A(n14433), .B(P1_REG0_REG_21__SCAN_IN), .S(n14924), .Z(
        P1_U3517) );
  MUX2_X1 U16279 ( .A(n14434), .B(P1_REG0_REG_20__SCAN_IN), .S(n14924), .Z(
        P1_U3516) );
  MUX2_X1 U16280 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n14435), .S(n14925), .Z(
        P1_U3515) );
  INV_X1 U16281 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14437) );
  MUX2_X1 U16282 ( .A(n14437), .B(n14436), .S(n14925), .Z(n14438) );
  INV_X1 U16283 ( .A(n14438), .ZN(P1_U3513) );
  MUX2_X1 U16284 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14439), .S(n14925), .Z(
        P1_U3510) );
  MUX2_X1 U16285 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14440), .S(n14925), .Z(
        P1_U3507) );
  NOR4_X1 U16286 ( .A1(n14442), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n14441), .ZN(n14443) );
  AOI21_X1 U16287 ( .B1(n14444), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14443), 
        .ZN(n14445) );
  OAI21_X1 U16288 ( .B1(n14446), .B2(n14458), .A(n14445), .ZN(P1_U3324) );
  INV_X1 U16289 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14447) );
  OAI222_X1 U16290 ( .A1(P1_U3086), .A2(n14449), .B1(n14458), .B2(n14448), 
        .C1(n14447), .C2(n14455), .ZN(P1_U3325) );
  OAI222_X1 U16291 ( .A1(P1_U3086), .A2(n14452), .B1(n14458), .B2(n14451), 
        .C1(n14450), .C2(n14455), .ZN(P1_U3326) );
  OAI222_X1 U16292 ( .A1(P1_U3086), .A2(n14454), .B1(n14458), .B2(n14453), 
        .C1(n7091), .C2(n14455), .ZN(P1_U3328) );
  OAI222_X1 U16293 ( .A1(P1_U3086), .A2(n9903), .B1(n14458), .B2(n14457), .C1(
        n14456), .C2(n14455), .ZN(P1_U3330) );
  MUX2_X1 U16294 ( .A(n6720), .B(n14459), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16295 ( .A(n14460), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U16296 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14551) );
  OR2_X1 U16297 ( .A1(n14551), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n14489) );
  NOR2_X1 U16298 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n14546), .ZN(n14488) );
  INV_X1 U16299 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14491) );
  INV_X1 U16300 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14757) );
  XOR2_X1 U16301 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n14757), .Z(n14495) );
  XOR2_X1 U16302 ( .A(n14484), .B(P1_ADDR_REG_11__SCAN_IN), .Z(n14496) );
  INV_X1 U16303 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14482) );
  XOR2_X1 U16304 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(P3_ADDR_REG_9__SCAN_IN), .Z(
        n14538) );
  INV_X1 U16305 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14477) );
  XOR2_X1 U16306 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n14477), .Z(n14500) );
  XOR2_X1 U16307 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14462), .Z(n14510) );
  NAND2_X1 U16308 ( .A1(n14510), .A2(n14511), .ZN(n14461) );
  NAND2_X1 U16309 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14464), .ZN(n14465) );
  NAND2_X1 U16310 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14466), .ZN(n14467) );
  NAND2_X1 U16311 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14468), .ZN(n14470) );
  NAND2_X1 U16312 ( .A1(n14470), .A2(n14469), .ZN(n14528) );
  NAND2_X1 U16313 ( .A1(n14473), .A2(n14472), .ZN(n14475) );
  XOR2_X1 U16314 ( .A(n14473), .B(n14472), .Z(n14532) );
  NAND2_X1 U16315 ( .A1(n14532), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U16316 ( .A1(n14475), .A2(n14474), .ZN(n14501) );
  NAND2_X1 U16317 ( .A1(n14500), .A2(n14501), .ZN(n14476) );
  NOR2_X1 U16318 ( .A1(n14538), .A2(n14537), .ZN(n14478) );
  XNOR2_X1 U16319 ( .A(n14480), .B(n14482), .ZN(n14498) );
  NAND2_X1 U16320 ( .A1(n14499), .A2(n14498), .ZN(n14481) );
  AND2_X1 U16321 ( .A1(n14491), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14486) );
  INV_X1 U16322 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14487) );
  OAI22_X1 U16323 ( .A1(n14488), .A2(n14548), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14487), .ZN(n14552) );
  AOI22_X1 U16324 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14551), .B1(n14489), 
        .B2(n14552), .ZN(n14559) );
  XNOR2_X1 U16325 ( .A(n11311), .B(P3_ADDR_REG_16__SCAN_IN), .ZN(n14490) );
  XOR2_X1 U16326 ( .A(n14559), .B(n14490), .Z(n14554) );
  XOR2_X1 U16327 ( .A(n14491), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n14493) );
  XOR2_X1 U16328 ( .A(n14493), .B(n14492), .Z(n14711) );
  XNOR2_X1 U16329 ( .A(n14495), .B(n14494), .ZN(n14706) );
  XOR2_X1 U16330 ( .A(n14497), .B(n14496), .Z(n14700) );
  XOR2_X1 U16331 ( .A(n14499), .B(n14498), .Z(n14594) );
  XOR2_X1 U16332 ( .A(n14501), .B(n14500), .Z(n14536) );
  INV_X1 U16333 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n14983) );
  OR2_X1 U16334 ( .A1(n14983), .A2(n14504), .ZN(n14518) );
  XNOR2_X1 U16335 ( .A(n14506), .B(n14505), .ZN(n14508) );
  NAND2_X1 U16336 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14508), .ZN(n14509) );
  AOI21_X1 U16337 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14507), .A(n14506), .ZN(
        n15429) );
  NOR2_X1 U16338 ( .A1(n15429), .A2(n15428), .ZN(n15438) );
  XNOR2_X1 U16339 ( .A(n14511), .B(n14510), .ZN(n14513) );
  NAND2_X1 U16340 ( .A1(n14512), .A2(n14513), .ZN(n14515) );
  NAND2_X1 U16341 ( .A1(n14570), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n14514) );
  NAND2_X1 U16342 ( .A1(n14515), .A2(n14514), .ZN(n15434) );
  XOR2_X1 U16343 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14516), .Z(n15433) );
  NOR2_X1 U16344 ( .A1(n15434), .A2(n15433), .ZN(n14517) );
  INV_X1 U16345 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15435) );
  NAND2_X1 U16346 ( .A1(n15434), .A2(n15433), .ZN(n15432) );
  OAI21_X1 U16347 ( .B1(n14517), .B2(n15435), .A(n15432), .ZN(n15425) );
  NOR2_X1 U16348 ( .A1(n14522), .A2(n14521), .ZN(n14523) );
  NAND2_X1 U16349 ( .A1(n14526), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14531) );
  INV_X1 U16350 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n14525) );
  XOR2_X1 U16351 ( .A(n14527), .B(P3_ADDR_REG_6__SCAN_IN), .Z(n14529) );
  XNOR2_X1 U16352 ( .A(n14529), .B(n14528), .ZN(n14581) );
  NAND2_X1 U16353 ( .A1(n14582), .A2(n14581), .ZN(n14530) );
  XOR2_X1 U16354 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14532), .Z(n15431) );
  NAND2_X1 U16355 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14533), .ZN(n14534) );
  XNOR2_X1 U16356 ( .A(n14538), .B(n14537), .ZN(n14539) );
  NAND2_X1 U16357 ( .A1(n14541), .A2(n14539), .ZN(n14543) );
  NAND2_X1 U16358 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n14592), .ZN(n14542) );
  NAND2_X1 U16359 ( .A1(n14543), .A2(n14542), .ZN(n14595) );
  NOR2_X1 U16360 ( .A1(n14594), .A2(n14595), .ZN(n14544) );
  INV_X1 U16361 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14999) );
  NAND2_X1 U16362 ( .A1(n14594), .A2(n14595), .ZN(n14593) );
  NOR2_X1 U16363 ( .A1(n14700), .A2(n14701), .ZN(n14545) );
  INV_X1 U16364 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n14702) );
  NAND2_X1 U16365 ( .A1(n14700), .A2(n14701), .ZN(n14699) );
  NAND2_X1 U16366 ( .A1(n14706), .A2(n14705), .ZN(n14704) );
  XNOR2_X1 U16367 ( .A(n14546), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n14547) );
  XOR2_X1 U16368 ( .A(n14548), .B(n14547), .Z(n14549) );
  NOR2_X1 U16369 ( .A1(n14550), .A2(n14549), .ZN(n14714) );
  XOR2_X1 U16370 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n14551), .Z(n14553) );
  XOR2_X1 U16371 ( .A(n14553), .B(n14552), .Z(n14717) );
  NOR2_X1 U16372 ( .A1(n14555), .A2(n14554), .ZN(n14556) );
  NOR2_X1 U16373 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14558), .ZN(n14560) );
  OAI22_X1 U16374 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n11311), .B1(n14560), 
        .B2(n14559), .ZN(n14564) );
  XOR2_X1 U16375 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14564), .Z(n14565) );
  XOR2_X1 U16376 ( .A(n14561), .B(n14565), .Z(n14562) );
  XNOR2_X1 U16377 ( .A(n14563), .B(n14562), .ZN(n14603) );
  NOR2_X1 U16378 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14564), .ZN(n14567) );
  AND2_X1 U16379 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14565), .ZN(n14566) );
  NOR2_X1 U16380 ( .A1(n14567), .A2(n14566), .ZN(n14607) );
  XOR2_X1 U16381 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n14016), .Z(n14608) );
  XOR2_X1 U16382 ( .A(n14607), .B(n14608), .Z(n14605) );
  XNOR2_X1 U16383 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14604), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16384 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14568) );
  OAI21_X1 U16385 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14568), 
        .ZN(U28) );
  AOI21_X1 U16386 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14569) );
  OAI21_X1 U16387 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14569), 
        .ZN(U29) );
  XOR2_X1 U16388 ( .A(n14570), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  AOI22_X1 U16389 ( .A1(n14571), .A2(n14587), .B1(SI_11_), .B2(n14586), .ZN(
        n14572) );
  OAI21_X1 U16390 ( .B1(P3_U3151), .B2(n14573), .A(n14572), .ZN(P3_U3284) );
  OAI22_X1 U16391 ( .A1(n14577), .A2(n14576), .B1(n14575), .B2(n14574), .ZN(
        n14578) );
  INV_X1 U16392 ( .A(n14578), .ZN(n14579) );
  OAI21_X1 U16393 ( .B1(P3_U3151), .B2(n14580), .A(n14579), .ZN(P3_U3283) );
  XOR2_X1 U16394 ( .A(n14582), .B(n14581), .Z(SUB_1596_U57) );
  AOI22_X1 U16395 ( .A1(n14583), .A2(n14587), .B1(SI_15_), .B2(n14586), .ZN(
        n14584) );
  OAI21_X1 U16396 ( .B1(P3_U3151), .B2(n14585), .A(n14584), .ZN(P3_U3280) );
  AOI22_X1 U16397 ( .A1(n14588), .A2(n14587), .B1(SI_16_), .B2(n14586), .ZN(
        n14589) );
  OAI21_X1 U16398 ( .B1(P3_U3151), .B2(n14590), .A(n14589), .ZN(P3_U3279) );
  XNOR2_X1 U16399 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14591), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16400 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14592), .Z(SUB_1596_U54) );
  OAI21_X1 U16401 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14596) );
  XOR2_X1 U16402 ( .A(n14596), .B(n14999), .Z(SUB_1596_U70) );
  OAI21_X1 U16403 ( .B1(n14598), .B2(n14920), .A(n14597), .ZN(n14600) );
  AOI211_X1 U16404 ( .C1(n14916), .C2(n14601), .A(n14600), .B(n14599), .ZN(
        n14602) );
  AOI22_X1 U16405 ( .A1(n14925), .A2(n14602), .B1(n9216), .B2(n14924), .ZN(
        P1_U3495) );
  AOI22_X1 U16406 ( .A1(n14940), .A2(n14602), .B1(n14741), .B2(n14937), .ZN(
        P1_U3540) );
  XNOR2_X1 U16407 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14603), .ZN(SUB_1596_U63)
         );
  NAND2_X1 U16408 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  OAI21_X1 U16409 ( .B1(n14016), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n14609), 
        .ZN(n14613) );
  XNOR2_X1 U16410 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14611) );
  XNOR2_X1 U16411 ( .A(n14611), .B(n14610), .ZN(n14612) );
  AOI22_X1 U16412 ( .A1(n14622), .A2(n14619), .B1(P3_REG2_REG_31__SCAN_IN), 
        .B2(n15371), .ZN(n14618) );
  AND2_X1 U16413 ( .A1(n14614), .A2(n15365), .ZN(n14617) );
  NOR2_X1 U16414 ( .A1(n14616), .A2(n14615), .ZN(n14624) );
  OAI21_X1 U16415 ( .B1(n14617), .B2(n14624), .A(n15369), .ZN(n14620) );
  NAND2_X1 U16416 ( .A1(n14618), .A2(n14620), .ZN(P3_U3202) );
  AOI22_X1 U16417 ( .A1(n14626), .A2(n14619), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n15371), .ZN(n14621) );
  NAND2_X1 U16418 ( .A1(n14621), .A2(n14620), .ZN(P3_U3203) );
  AOI21_X1 U16419 ( .B1(n14622), .B2(n14625), .A(n14624), .ZN(n14642) );
  INV_X1 U16420 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14623) );
  AOI22_X1 U16421 ( .A1(n15424), .A2(n14642), .B1(n14623), .B2(n8836), .ZN(
        P3_U3490) );
  AOI21_X1 U16422 ( .B1(n14626), .B2(n14625), .A(n14624), .ZN(n14644) );
  INV_X1 U16423 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14627) );
  AOI22_X1 U16424 ( .A1(n15424), .A2(n14644), .B1(n14627), .B2(n8836), .ZN(
        P3_U3489) );
  OAI21_X1 U16425 ( .B1(n15406), .B2(n14629), .A(n14628), .ZN(n14630) );
  AOI21_X1 U16426 ( .B1(n14631), .B2(n14640), .A(n14630), .ZN(n14646) );
  INV_X1 U16427 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14632) );
  AOI22_X1 U16428 ( .A1(n15424), .A2(n14646), .B1(n14632), .B2(n8836), .ZN(
        P3_U3472) );
  AOI211_X1 U16429 ( .C1(n14635), .C2(n14640), .A(n14634), .B(n14633), .ZN(
        n14648) );
  AOI22_X1 U16430 ( .A1(n15424), .A2(n14648), .B1(n14636), .B2(n8836), .ZN(
        P3_U3471) );
  AOI211_X1 U16431 ( .C1(n14640), .C2(n14639), .A(n14638), .B(n14637), .ZN(
        n14649) );
  INV_X1 U16432 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14641) );
  AOI22_X1 U16433 ( .A1(n15424), .A2(n14649), .B1(n14641), .B2(n8836), .ZN(
        P3_U3470) );
  INV_X1 U16434 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14643) );
  AOI22_X1 U16435 ( .A1(n15412), .A2(n14643), .B1(n14642), .B2(n15411), .ZN(
        P3_U3458) );
  INV_X1 U16436 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14645) );
  AOI22_X1 U16437 ( .A1(n15412), .A2(n14645), .B1(n14644), .B2(n15411), .ZN(
        P3_U3457) );
  INV_X1 U16438 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14647) );
  AOI22_X1 U16439 ( .A1(n15412), .A2(n14647), .B1(n14646), .B2(n15411), .ZN(
        P3_U3429) );
  AOI22_X1 U16440 ( .A1(n15412), .A2(n7686), .B1(n14648), .B2(n15411), .ZN(
        P3_U3426) );
  AOI22_X1 U16441 ( .A1(n15412), .A2(n7672), .B1(n14649), .B2(n15411), .ZN(
        P3_U3423) );
  OAI211_X1 U16442 ( .C1(n7209), .C2(n15146), .A(n14652), .B(n14651), .ZN(
        n14653) );
  AOI21_X1 U16443 ( .B1(n14654), .B2(n15151), .A(n14653), .ZN(n14655) );
  AOI22_X1 U16444 ( .A1(n15160), .A2(n14655), .B1(n10797), .B2(n15164), .ZN(
        P2_U3512) );
  AOI22_X1 U16445 ( .A1(n15155), .A2(n14655), .B1(n8436), .B2(n15153), .ZN(
        P2_U3469) );
  OAI21_X1 U16446 ( .B1(n14657), .B2(n6669), .A(n14656), .ZN(n14666) );
  INV_X1 U16447 ( .A(n14658), .ZN(n14679) );
  NOR2_X1 U16448 ( .A1(n14679), .A2(n14659), .ZN(n14665) );
  OAI22_X1 U16449 ( .A1(n14663), .A2(n14662), .B1(n14661), .B2(n14660), .ZN(
        n14664) );
  AOI211_X1 U16450 ( .C1(n14666), .C2(n14726), .A(n14665), .B(n14664), .ZN(
        n14668) );
  OAI211_X1 U16451 ( .C1(n14736), .C2(n14669), .A(n14668), .B(n14667), .ZN(
        P1_U3215) );
  OAI21_X1 U16452 ( .B1(n6955), .B2(n14920), .A(n14670), .ZN(n14672) );
  AOI211_X1 U16453 ( .C1(n14922), .C2(n14673), .A(n14672), .B(n14671), .ZN(
        n14694) );
  AOI22_X1 U16454 ( .A1(n14940), .A2(n14694), .B1(n14674), .B2(n14937), .ZN(
        P1_U3543) );
  NAND3_X1 U16455 ( .A1(n14676), .A2(n14675), .A3(n14922), .ZN(n14678) );
  OAI211_X1 U16456 ( .C1(n14679), .C2(n14920), .A(n14678), .B(n14677), .ZN(
        n14680) );
  INV_X1 U16457 ( .A(n14680), .ZN(n14681) );
  AND2_X1 U16458 ( .A1(n14682), .A2(n14681), .ZN(n14696) );
  AOI22_X1 U16459 ( .A1(n14940), .A2(n14696), .B1(n10722), .B2(n14937), .ZN(
        P1_U3542) );
  OAI21_X1 U16460 ( .B1(n14684), .B2(n14920), .A(n14683), .ZN(n14686) );
  AOI211_X1 U16461 ( .C1(n14687), .C2(n14922), .A(n14686), .B(n14685), .ZN(
        n14697) );
  AOI22_X1 U16462 ( .A1(n14940), .A2(n14697), .B1(n10558), .B2(n14937), .ZN(
        P1_U3541) );
  OAI21_X1 U16463 ( .B1(n14689), .B2(n14920), .A(n14688), .ZN(n14691) );
  AOI211_X1 U16464 ( .C1(n14692), .C2(n14922), .A(n14691), .B(n14690), .ZN(
        n14698) );
  AOI22_X1 U16465 ( .A1(n14940), .A2(n14698), .B1(n14693), .B2(n14937), .ZN(
        P1_U3539) );
  AOI22_X1 U16466 ( .A1(n14925), .A2(n14694), .B1(n9271), .B2(n14924), .ZN(
        P1_U3504) );
  AOI22_X1 U16467 ( .A1(n14925), .A2(n14696), .B1(n14695), .B2(n14924), .ZN(
        P1_U3501) );
  AOI22_X1 U16468 ( .A1(n14925), .A2(n14697), .B1(n9246), .B2(n14924), .ZN(
        P1_U3498) );
  AOI22_X1 U16469 ( .A1(n14925), .A2(n14698), .B1(n9200), .B2(n14924), .ZN(
        P1_U3492) );
  OAI21_X1 U16470 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14703) );
  XOR2_X1 U16471 ( .A(n14703), .B(n14702), .Z(SUB_1596_U69) );
  OAI21_X1 U16472 ( .B1(n14706), .B2(n14705), .A(n14704), .ZN(n14708) );
  XOR2_X1 U16473 ( .A(n14708), .B(n14707), .Z(SUB_1596_U68) );
  AOI21_X1 U16474 ( .B1(n14711), .B2(n14710), .A(n14709), .ZN(n14712) );
  XOR2_X1 U16475 ( .A(n14712), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  NOR2_X1 U16476 ( .A1(n14714), .A2(n14713), .ZN(n14715) );
  XOR2_X1 U16477 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n14715), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16478 ( .B1(n14718), .B2(n14717), .A(n14716), .ZN(n14719) );
  XOR2_X1 U16479 ( .A(n14719), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  XNOR2_X1 U16480 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14720), .ZN(SUB_1596_U64)
         );
  NAND2_X1 U16481 ( .A1(n14722), .A2(n14721), .ZN(n14872) );
  INV_X1 U16482 ( .A(n14872), .ZN(n14724) );
  AOI22_X1 U16483 ( .A1(n14725), .A2(n14724), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14735) );
  OAI211_X1 U16484 ( .C1(n14729), .C2(n14728), .A(n14727), .B(n14726), .ZN(
        n14730) );
  INV_X1 U16485 ( .A(n14730), .ZN(n14731) );
  AOI21_X1 U16486 ( .B1(n14733), .B2(n14732), .A(n14731), .ZN(n14734) );
  OAI211_X1 U16487 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n14736), .A(n14735), .B(
        n14734), .ZN(P1_U3218) );
  INV_X1 U16488 ( .A(n14737), .ZN(n14738) );
  OAI21_X1 U16489 ( .B1(n14740), .B2(n14739), .A(n14738), .ZN(n14753) );
  MUX2_X1 U16490 ( .A(n14741), .B(P1_REG1_REG_12__SCAN_IN), .S(n14751), .Z(
        n14744) );
  INV_X1 U16491 ( .A(n14742), .ZN(n14743) );
  NAND2_X1 U16492 ( .A1(n14744), .A2(n14743), .ZN(n14746) );
  OAI21_X1 U16493 ( .B1(n14747), .B2(n14746), .A(n14745), .ZN(n14749) );
  AOI222_X1 U16494 ( .A1(n14753), .A2(n14752), .B1(n14751), .B2(n14750), .C1(
        n14749), .C2(n14748), .ZN(n14755) );
  OAI211_X1 U16495 ( .C1(n14757), .C2(n14756), .A(n14755), .B(n14754), .ZN(
        P1_U3255) );
  XNOR2_X1 U16496 ( .A(n14758), .B(n14763), .ZN(n14905) );
  OAI21_X1 U16497 ( .B1(n14759), .B2(n14907), .A(n14812), .ZN(n14760) );
  OR2_X1 U16498 ( .A1(n14761), .A2(n14760), .ZN(n14906) );
  INV_X1 U16499 ( .A(n14906), .ZN(n14762) );
  AOI22_X1 U16500 ( .A1(n14905), .A2(n14828), .B1(n14818), .B2(n14762), .ZN(
        n14780) );
  NAND2_X1 U16501 ( .A1(n14764), .A2(n14763), .ZN(n14765) );
  NAND3_X1 U16502 ( .A1(n14767), .A2(n14766), .A3(n14765), .ZN(n14773) );
  AOI22_X1 U16503 ( .A1(n14771), .A2(n14770), .B1(n14769), .B2(n14768), .ZN(
        n14772) );
  NAND2_X1 U16504 ( .A1(n14773), .A2(n14772), .ZN(n14910) );
  MUX2_X1 U16505 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14910), .S(n14774), .Z(
        n14778) );
  OAI22_X1 U16506 ( .A1(n14907), .A2(n14808), .B1(n14776), .B2(n14775), .ZN(
        n14777) );
  NOR2_X1 U16507 ( .A1(n14778), .A2(n14777), .ZN(n14779) );
  NAND2_X1 U16508 ( .A1(n14780), .A2(n14779), .ZN(P1_U3285) );
  XNOR2_X1 U16509 ( .A(n14781), .B(n14783), .ZN(n14895) );
  NAND3_X1 U16510 ( .A1(n10913), .A2(n14783), .A3(n14782), .ZN(n14784) );
  AOI21_X1 U16511 ( .B1(n14785), .B2(n14784), .A(n14802), .ZN(n14786) );
  AOI211_X1 U16512 ( .C1(n14899), .C2(n14895), .A(n14787), .B(n14786), .ZN(
        n14892) );
  INV_X1 U16513 ( .A(n14788), .ZN(n14891) );
  AOI22_X1 U16514 ( .A1(n14833), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n14789), 
        .B2(n14826), .ZN(n14790) );
  OAI21_X1 U16515 ( .B1(n14808), .B2(n14891), .A(n14790), .ZN(n14791) );
  INV_X1 U16516 ( .A(n14791), .ZN(n14798) );
  INV_X1 U16517 ( .A(n14792), .ZN(n14795) );
  INV_X1 U16518 ( .A(n14793), .ZN(n14794) );
  OAI211_X1 U16519 ( .C1(n14891), .C2(n14795), .A(n14794), .B(n14812), .ZN(
        n14890) );
  INV_X1 U16520 ( .A(n14890), .ZN(n14796) );
  AOI22_X1 U16521 ( .A1(n14895), .A2(n14816), .B1(n14818), .B2(n14796), .ZN(
        n14797) );
  OAI211_X1 U16522 ( .C1(n14833), .C2(n14892), .A(n14798), .B(n14797), .ZN(
        P1_U3287) );
  XNOR2_X1 U16523 ( .A(n14800), .B(n14799), .ZN(n14871) );
  NAND2_X1 U16524 ( .A1(n14801), .A2(n14800), .ZN(n14803) );
  AOI21_X1 U16525 ( .B1(n14804), .B2(n14803), .A(n14802), .ZN(n14805) );
  AOI211_X1 U16526 ( .C1(n14899), .C2(n14871), .A(n14806), .B(n14805), .ZN(
        n14868) );
  AOI22_X1 U16527 ( .A1(n14833), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n14826), .ZN(n14807) );
  OAI21_X1 U16528 ( .B1(n14808), .B2(n9043), .A(n14807), .ZN(n14809) );
  INV_X1 U16529 ( .A(n14809), .ZN(n14820) );
  NAND2_X1 U16530 ( .A1(n14811), .A2(n14810), .ZN(n14813) );
  NAND2_X1 U16531 ( .A1(n14813), .A2(n14812), .ZN(n14815) );
  OR2_X1 U16532 ( .A1(n14815), .A2(n14814), .ZN(n14867) );
  INV_X1 U16533 ( .A(n14867), .ZN(n14817) );
  AOI22_X1 U16534 ( .A1(n14818), .A2(n14817), .B1(n14816), .B2(n14871), .ZN(
        n14819) );
  OAI211_X1 U16535 ( .C1(n14833), .C2(n14868), .A(n14820), .B(n14819), .ZN(
        P1_U3291) );
  INV_X1 U16536 ( .A(n14821), .ZN(n14825) );
  INV_X1 U16537 ( .A(n14822), .ZN(n14823) );
  AOI21_X1 U16538 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n14832) );
  AOI22_X1 U16539 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(n14833), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(n14826), .ZN(n14831) );
  OAI21_X1 U16540 ( .B1(n14829), .B2(n14828), .A(n14827), .ZN(n14830) );
  OAI211_X1 U16541 ( .C1(n14833), .C2(n14832), .A(n14831), .B(n14830), .ZN(
        P1_U3293) );
  INV_X1 U16542 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14834) );
  NOR2_X1 U16543 ( .A1(n14864), .A2(n14834), .ZN(P1_U3294) );
  INV_X1 U16544 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14835) );
  NOR2_X1 U16545 ( .A1(n14864), .A2(n14835), .ZN(P1_U3295) );
  INV_X1 U16546 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14836) );
  NOR2_X1 U16547 ( .A1(n14864), .A2(n14836), .ZN(P1_U3296) );
  INV_X1 U16548 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14837) );
  NOR2_X1 U16549 ( .A1(n14864), .A2(n14837), .ZN(P1_U3297) );
  NOR2_X1 U16550 ( .A1(n14864), .A2(n14838), .ZN(P1_U3298) );
  NOR2_X1 U16551 ( .A1(n14864), .A2(n14839), .ZN(P1_U3299) );
  NOR2_X1 U16552 ( .A1(n14864), .A2(n14840), .ZN(P1_U3300) );
  NOR2_X1 U16553 ( .A1(n14864), .A2(n14841), .ZN(P1_U3301) );
  INV_X1 U16554 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14842) );
  NOR2_X1 U16555 ( .A1(n14864), .A2(n14842), .ZN(P1_U3302) );
  NOR2_X1 U16556 ( .A1(n14864), .A2(n14843), .ZN(P1_U3303) );
  INV_X1 U16557 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14844) );
  NOR2_X1 U16558 ( .A1(n14864), .A2(n14844), .ZN(P1_U3304) );
  INV_X1 U16559 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14845) );
  NOR2_X1 U16560 ( .A1(n14864), .A2(n14845), .ZN(P1_U3305) );
  INV_X1 U16561 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14846) );
  NOR2_X1 U16562 ( .A1(n14864), .A2(n14846), .ZN(P1_U3306) );
  INV_X1 U16563 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14847) );
  NOR2_X1 U16564 ( .A1(n14864), .A2(n14847), .ZN(P1_U3307) );
  NOR2_X1 U16565 ( .A1(n14864), .A2(n14848), .ZN(P1_U3308) );
  INV_X1 U16566 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14849) );
  NOR2_X1 U16567 ( .A1(n14864), .A2(n14849), .ZN(P1_U3309) );
  NOR2_X1 U16568 ( .A1(n14864), .A2(n14850), .ZN(P1_U3310) );
  NOR2_X1 U16569 ( .A1(n14864), .A2(n14851), .ZN(P1_U3311) );
  INV_X1 U16570 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14852) );
  NOR2_X1 U16571 ( .A1(n14864), .A2(n14852), .ZN(P1_U3312) );
  INV_X1 U16572 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14853) );
  NOR2_X1 U16573 ( .A1(n14864), .A2(n14853), .ZN(P1_U3313) );
  INV_X1 U16574 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14854) );
  NOR2_X1 U16575 ( .A1(n14864), .A2(n14854), .ZN(P1_U3314) );
  INV_X1 U16576 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14855) );
  NOR2_X1 U16577 ( .A1(n14864), .A2(n14855), .ZN(P1_U3315) );
  INV_X1 U16578 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14856) );
  NOR2_X1 U16579 ( .A1(n14864), .A2(n14856), .ZN(P1_U3316) );
  INV_X1 U16580 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14857) );
  NOR2_X1 U16581 ( .A1(n14864), .A2(n14857), .ZN(P1_U3317) );
  INV_X1 U16582 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14858) );
  NOR2_X1 U16583 ( .A1(n14864), .A2(n14858), .ZN(P1_U3318) );
  INV_X1 U16584 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14859) );
  NOR2_X1 U16585 ( .A1(n14864), .A2(n14859), .ZN(P1_U3319) );
  INV_X1 U16586 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14860) );
  NOR2_X1 U16587 ( .A1(n14864), .A2(n14860), .ZN(P1_U3320) );
  INV_X1 U16588 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14861) );
  NOR2_X1 U16589 ( .A1(n14864), .A2(n14861), .ZN(P1_U3321) );
  INV_X1 U16590 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14862) );
  NOR2_X1 U16591 ( .A1(n14864), .A2(n14862), .ZN(P1_U3322) );
  INV_X1 U16592 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14863) );
  NOR2_X1 U16593 ( .A1(n14864), .A2(n14863), .ZN(P1_U3323) );
  INV_X1 U16594 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14865) );
  AOI22_X1 U16595 ( .A1(n14925), .A2(n14866), .B1(n14865), .B2(n14924), .ZN(
        P1_U3462) );
  OAI21_X1 U16596 ( .B1(n9043), .B2(n14920), .A(n14867), .ZN(n14870) );
  INV_X1 U16597 ( .A(n14868), .ZN(n14869) );
  AOI211_X1 U16598 ( .C1(n14916), .C2(n14871), .A(n14870), .B(n14869), .ZN(
        n14926) );
  AOI22_X1 U16599 ( .A1(n14925), .A2(n14926), .B1(n9038), .B2(n14924), .ZN(
        P1_U3465) );
  NAND2_X1 U16600 ( .A1(n14877), .A2(n14899), .ZN(n14874) );
  NAND4_X1 U16601 ( .A1(n14875), .A2(n14874), .A3(n14873), .A4(n14872), .ZN(
        n14876) );
  AOI21_X1 U16602 ( .B1(n14916), .B2(n14877), .A(n14876), .ZN(n14927) );
  AOI22_X1 U16603 ( .A1(n14925), .A2(n14927), .B1(n9047), .B2(n14924), .ZN(
        P1_U3468) );
  OR4_X1 U16604 ( .A1(n14881), .A2(n14880), .A3(n14879), .A4(n14878), .ZN(
        n14882) );
  AOI21_X1 U16605 ( .B1(n14922), .B2(n14883), .A(n14882), .ZN(n14928) );
  AOI22_X1 U16606 ( .A1(n14925), .A2(n14928), .B1(n9073), .B2(n14924), .ZN(
        P1_U3471) );
  NAND2_X1 U16607 ( .A1(n14889), .A2(n14899), .ZN(n14884) );
  NAND4_X1 U16608 ( .A1(n14887), .A2(n14886), .A3(n14885), .A4(n14884), .ZN(
        n14888) );
  AOI21_X1 U16609 ( .B1(n14916), .B2(n14889), .A(n14888), .ZN(n14929) );
  AOI22_X1 U16610 ( .A1(n14925), .A2(n14929), .B1(n9087), .B2(n14924), .ZN(
        P1_U3474) );
  OAI21_X1 U16611 ( .B1(n14891), .B2(n14920), .A(n14890), .ZN(n14894) );
  INV_X1 U16612 ( .A(n14892), .ZN(n14893) );
  AOI211_X1 U16613 ( .C1(n14916), .C2(n14895), .A(n14894), .B(n14893), .ZN(
        n14930) );
  AOI22_X1 U16614 ( .A1(n14925), .A2(n14930), .B1(n9108), .B2(n14924), .ZN(
        P1_U3477) );
  OAI21_X1 U16615 ( .B1(n14897), .B2(n14920), .A(n14896), .ZN(n14898) );
  INV_X1 U16616 ( .A(n14898), .ZN(n14903) );
  NAND2_X1 U16617 ( .A1(n14900), .A2(n14916), .ZN(n14902) );
  NAND2_X1 U16618 ( .A1(n14900), .A2(n14899), .ZN(n14901) );
  AOI22_X1 U16619 ( .A1(n14925), .A2(n14932), .B1(n9128), .B2(n14924), .ZN(
        P1_U3480) );
  AND2_X1 U16620 ( .A1(n14905), .A2(n14922), .ZN(n14909) );
  OAI21_X1 U16621 ( .B1(n14907), .B2(n14920), .A(n14906), .ZN(n14908) );
  NOR3_X1 U16622 ( .A1(n14910), .A2(n14909), .A3(n14908), .ZN(n14934) );
  AOI22_X1 U16623 ( .A1(n14925), .A2(n14934), .B1(n9143), .B2(n14924), .ZN(
        P1_U3483) );
  OAI21_X1 U16624 ( .B1(n14912), .B2(n14920), .A(n14911), .ZN(n14914) );
  AOI211_X1 U16625 ( .C1(n14916), .C2(n14915), .A(n14914), .B(n14913), .ZN(
        n14936) );
  AOI22_X1 U16626 ( .A1(n14925), .A2(n14936), .B1(n9163), .B2(n14924), .ZN(
        P1_U3486) );
  OAI211_X1 U16627 ( .C1(n6953), .C2(n14920), .A(n14919), .B(n14918), .ZN(
        n14921) );
  AOI21_X1 U16628 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14939) );
  AOI22_X1 U16629 ( .A1(n14925), .A2(n14939), .B1(n9175), .B2(n14924), .ZN(
        P1_U3489) );
  AOI22_X1 U16630 ( .A1(n14940), .A2(n14926), .B1(n10102), .B2(n14937), .ZN(
        P1_U3530) );
  AOI22_X1 U16631 ( .A1(n14940), .A2(n14927), .B1(n10103), .B2(n14937), .ZN(
        P1_U3531) );
  AOI22_X1 U16632 ( .A1(n14940), .A2(n14928), .B1(n10104), .B2(n14937), .ZN(
        P1_U3532) );
  AOI22_X1 U16633 ( .A1(n14940), .A2(n14929), .B1(n10106), .B2(n14937), .ZN(
        P1_U3533) );
  AOI22_X1 U16634 ( .A1(n14940), .A2(n14930), .B1(n10108), .B2(n14937), .ZN(
        P1_U3534) );
  AOI22_X1 U16635 ( .A1(n14940), .A2(n14932), .B1(n14931), .B2(n14937), .ZN(
        P1_U3535) );
  AOI22_X1 U16636 ( .A1(n14940), .A2(n14934), .B1(n14933), .B2(n14937), .ZN(
        P1_U3536) );
  AOI22_X1 U16637 ( .A1(n14940), .A2(n14936), .B1(n14935), .B2(n14937), .ZN(
        P1_U3537) );
  AOI22_X1 U16638 ( .A1(n14940), .A2(n14939), .B1(n14938), .B2(n14937), .ZN(
        P1_U3538) );
  NOR2_X1 U16639 ( .A1(n15007), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16640 ( .A1(n14976), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15009), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U16641 ( .A1(n15007), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14943) );
  OAI22_X1 U16642 ( .A1(n14993), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n15001), .ZN(n14941) );
  OAI21_X1 U16643 ( .B1(n14991), .B2(n14941), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n14942) );
  OAI211_X1 U16644 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n14944), .A(n14943), .B(
        n14942), .ZN(P2_U3214) );
  AOI22_X1 U16645 ( .A1(n15007), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14956) );
  XNOR2_X1 U16646 ( .A(n14946), .B(n14945), .ZN(n14948) );
  OAI22_X1 U16647 ( .A1(n15001), .A2(n14948), .B1(n14947), .B2(n15014), .ZN(
        n14949) );
  INV_X1 U16648 ( .A(n14949), .ZN(n14955) );
  NOR2_X1 U16649 ( .A1(n14950), .A2(n13396), .ZN(n14953) );
  OAI211_X1 U16650 ( .C1(n14953), .C2(n14952), .A(n15009), .B(n14951), .ZN(
        n14954) );
  NAND3_X1 U16651 ( .A1(n14956), .A2(n14955), .A3(n14954), .ZN(P2_U3215) );
  AOI22_X1 U16652 ( .A1(n15007), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14968) );
  OAI21_X1 U16653 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n14961) );
  OAI22_X1 U16654 ( .A1(n15001), .A2(n14961), .B1(n14960), .B2(n15014), .ZN(
        n14962) );
  INV_X1 U16655 ( .A(n14962), .ZN(n14967) );
  OAI211_X1 U16656 ( .C1(n14965), .C2(n14964), .A(n15009), .B(n14963), .ZN(
        n14966) );
  NAND3_X1 U16657 ( .A1(n14968), .A2(n14967), .A3(n14966), .ZN(P2_U3216) );
  NOR2_X1 U16658 ( .A1(n14970), .A2(n14969), .ZN(n14971) );
  OAI21_X1 U16659 ( .B1(n15014), .B2(n14973), .A(n14972), .ZN(n14974) );
  AOI21_X1 U16660 ( .B1(n14976), .B2(n14975), .A(n14974), .ZN(n14982) );
  AOI211_X1 U16661 ( .C1(n14979), .C2(n14978), .A(n14977), .B(n14993), .ZN(
        n14980) );
  INV_X1 U16662 ( .A(n14980), .ZN(n14981) );
  OAI211_X1 U16663 ( .C1(n15000), .C2(n14983), .A(n14982), .B(n14981), .ZN(
        P2_U3218) );
  NOR2_X1 U16664 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14984), .ZN(n14989) );
  AOI211_X1 U16665 ( .C1(n14987), .C2(n14986), .A(n15001), .B(n14985), .ZN(
        n14988) );
  AOI211_X1 U16666 ( .C1(n14991), .C2(n14990), .A(n14989), .B(n14988), .ZN(
        n14998) );
  AOI211_X1 U16667 ( .C1(n14995), .C2(n14994), .A(n14993), .B(n14992), .ZN(
        n14996) );
  INV_X1 U16668 ( .A(n14996), .ZN(n14997) );
  OAI211_X1 U16669 ( .C1(n15000), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        P2_U3224) );
  AND2_X1 U16670 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n15006) );
  AOI211_X1 U16671 ( .C1(n15004), .C2(n15003), .A(n15002), .B(n15001), .ZN(
        n15005) );
  AOI211_X1 U16672 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n15007), .A(n15006), 
        .B(n15005), .ZN(n15012) );
  OAI211_X1 U16673 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n15010), .A(n15009), 
        .B(n15008), .ZN(n15011) );
  OAI211_X1 U16674 ( .C1(n15014), .C2(n15013), .A(n15012), .B(n15011), .ZN(
        P2_U3229) );
  XNOR2_X1 U16675 ( .A(n15015), .B(n15016), .ZN(n15019) );
  AOI21_X1 U16676 ( .B1(n15019), .B2(n15018), .A(n15017), .ZN(n15148) );
  OAI211_X1 U16677 ( .C1(n15147), .C2(n15022), .A(n15021), .B(n15020), .ZN(
        n15145) );
  OR2_X1 U16678 ( .A1(n15145), .A2(n15023), .ZN(n15030) );
  NAND2_X1 U16679 ( .A1(n15038), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n15024) );
  OAI21_X1 U16680 ( .B1(n15050), .B2(n15025), .A(n15024), .ZN(n15026) );
  AOI21_X1 U16681 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15029) );
  AND2_X1 U16682 ( .A1(n15030), .A2(n15029), .ZN(n15037) );
  OAI21_X1 U16683 ( .B1(n15033), .B2(n15032), .A(n15031), .ZN(n15034) );
  INV_X1 U16684 ( .A(n15034), .ZN(n15152) );
  NAND2_X1 U16685 ( .A1(n15152), .A2(n15035), .ZN(n15036) );
  OAI211_X1 U16686 ( .C1(n15038), .C2(n15148), .A(n15037), .B(n15036), .ZN(
        P2_U3254) );
  NAND2_X1 U16687 ( .A1(n15119), .A2(n15039), .ZN(n15041) );
  AOI21_X1 U16688 ( .B1(n15092), .B2(n15041), .A(n15040), .ZN(n15089) );
  NOR2_X1 U16689 ( .A1(n15043), .A2(n15042), .ZN(n15091) );
  AOI22_X1 U16690 ( .A1(n15091), .A2(n15045), .B1(n15092), .B2(n15044), .ZN(
        n15046) );
  NAND3_X1 U16691 ( .A1(n15048), .A2(n15089), .A3(n15046), .ZN(n15047) );
  OAI21_X1 U16692 ( .B1(n15048), .B2(P2_REG2_REG_0__SCAN_IN), .A(n15047), .ZN(
        n15049) );
  OAI21_X1 U16693 ( .B1(n15050), .B2(n8190), .A(n15049), .ZN(P2_U3265) );
  NOR2_X1 U16694 ( .A1(n15083), .A2(n15052), .ZN(P2_U3266) );
  INV_X1 U16695 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15053) );
  NOR2_X1 U16696 ( .A1(n15083), .A2(n15053), .ZN(P2_U3267) );
  INV_X1 U16697 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n15054) );
  NOR2_X1 U16698 ( .A1(n15083), .A2(n15054), .ZN(P2_U3268) );
  INV_X1 U16699 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n15055) );
  NOR2_X1 U16700 ( .A1(n15079), .A2(n15055), .ZN(P2_U3269) );
  INV_X1 U16701 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n15056) );
  NOR2_X1 U16702 ( .A1(n15079), .A2(n15056), .ZN(P2_U3270) );
  INV_X1 U16703 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n15057) );
  NOR2_X1 U16704 ( .A1(n15079), .A2(n15057), .ZN(P2_U3271) );
  NOR2_X1 U16705 ( .A1(n15079), .A2(n15058), .ZN(P2_U3272) );
  INV_X1 U16706 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n15059) );
  NOR2_X1 U16707 ( .A1(n15079), .A2(n15059), .ZN(P2_U3273) );
  INV_X1 U16708 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n15060) );
  NOR2_X1 U16709 ( .A1(n15079), .A2(n15060), .ZN(P2_U3274) );
  INV_X1 U16710 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n15061) );
  NOR2_X1 U16711 ( .A1(n15079), .A2(n15061), .ZN(P2_U3275) );
  INV_X1 U16712 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n15062) );
  NOR2_X1 U16713 ( .A1(n15079), .A2(n15062), .ZN(P2_U3276) );
  INV_X1 U16714 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n15063) );
  NOR2_X1 U16715 ( .A1(n15079), .A2(n15063), .ZN(P2_U3277) );
  NOR2_X1 U16716 ( .A1(n15083), .A2(n15064), .ZN(P2_U3278) );
  INV_X1 U16717 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n15065) );
  NOR2_X1 U16718 ( .A1(n15083), .A2(n15065), .ZN(P2_U3279) );
  INV_X1 U16719 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n15066) );
  NOR2_X1 U16720 ( .A1(n15083), .A2(n15066), .ZN(P2_U3280) );
  INV_X1 U16721 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n15067) );
  NOR2_X1 U16722 ( .A1(n15083), .A2(n15067), .ZN(P2_U3281) );
  INV_X1 U16723 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n15068) );
  NOR2_X1 U16724 ( .A1(n15083), .A2(n15068), .ZN(P2_U3282) );
  INV_X1 U16725 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n15069) );
  NOR2_X1 U16726 ( .A1(n15083), .A2(n15069), .ZN(P2_U3283) );
  INV_X1 U16727 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n15070) );
  NOR2_X1 U16728 ( .A1(n15083), .A2(n15070), .ZN(P2_U3284) );
  INV_X1 U16729 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n15071) );
  NOR2_X1 U16730 ( .A1(n15083), .A2(n15071), .ZN(P2_U3285) );
  INV_X1 U16731 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U16732 ( .A1(n15083), .A2(n15072), .ZN(P2_U3286) );
  INV_X1 U16733 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n15073) );
  NOR2_X1 U16734 ( .A1(n15083), .A2(n15073), .ZN(P2_U3287) );
  INV_X1 U16735 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n15074) );
  NOR2_X1 U16736 ( .A1(n15083), .A2(n15074), .ZN(P2_U3288) );
  INV_X1 U16737 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n15075) );
  NOR2_X1 U16738 ( .A1(n15083), .A2(n15075), .ZN(P2_U3289) );
  INV_X1 U16739 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n15076) );
  NOR2_X1 U16740 ( .A1(n15079), .A2(n15076), .ZN(P2_U3290) );
  INV_X1 U16741 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n15077) );
  NOR2_X1 U16742 ( .A1(n15083), .A2(n15077), .ZN(P2_U3291) );
  INV_X1 U16743 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n15078) );
  NOR2_X1 U16744 ( .A1(n15079), .A2(n15078), .ZN(P2_U3292) );
  INV_X1 U16745 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n15080) );
  NOR2_X1 U16746 ( .A1(n15083), .A2(n15080), .ZN(P2_U3293) );
  INV_X1 U16747 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n15081) );
  NOR2_X1 U16748 ( .A1(n15083), .A2(n15081), .ZN(P2_U3294) );
  NOR2_X1 U16749 ( .A1(n15083), .A2(n15082), .ZN(P2_U3295) );
  OAI22_X1 U16750 ( .A1(n15086), .A2(n15084), .B1(P2_D_REG_0__SCAN_IN), .B2(
        n15088), .ZN(n15085) );
  INV_X1 U16751 ( .A(n15085), .ZN(P2_U3416) );
  AOI22_X1 U16752 ( .A1(n15088), .A2(n15087), .B1(n8761), .B2(n15086), .ZN(
        P2_U3417) );
  INV_X1 U16753 ( .A(n15089), .ZN(n15090) );
  AOI211_X1 U16754 ( .C1(n15124), .C2(n15092), .A(n15091), .B(n15090), .ZN(
        n15156) );
  AOI22_X1 U16755 ( .A1(n15155), .A2(n15156), .B1(n15093), .B2(n15153), .ZN(
        P2_U3430) );
  INV_X1 U16756 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15094) );
  AOI22_X1 U16757 ( .A1(n15155), .A2(n15095), .B1(n15094), .B2(n15153), .ZN(
        P2_U3436) );
  AND2_X1 U16758 ( .A1(n15096), .A2(n15124), .ZN(n15100) );
  OAI21_X1 U16759 ( .B1(n15098), .B2(n15146), .A(n15097), .ZN(n15099) );
  NOR3_X1 U16760 ( .A1(n15101), .A2(n15100), .A3(n15099), .ZN(n15157) );
  INV_X1 U16761 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U16762 ( .A1(n15155), .A2(n15157), .B1(n15102), .B2(n15153), .ZN(
        P2_U3445) );
  NAND3_X1 U16763 ( .A1(n15104), .A2(n15103), .A3(n15151), .ZN(n15108) );
  AOI21_X1 U16764 ( .B1(n15137), .B2(n15106), .A(n15105), .ZN(n15107) );
  AOI22_X1 U16765 ( .A1(n15155), .A2(n15158), .B1(n8299), .B2(n15153), .ZN(
        P2_U3448) );
  INV_X1 U16766 ( .A(n15110), .ZN(n15115) );
  OAI21_X1 U16767 ( .B1(n15112), .B2(n15146), .A(n15111), .ZN(n15114) );
  AOI211_X1 U16768 ( .C1(n15115), .C2(n15151), .A(n15114), .B(n15113), .ZN(
        n15159) );
  AOI22_X1 U16769 ( .A1(n15155), .A2(n15159), .B1(n8321), .B2(n15153), .ZN(
        P2_U3451) );
  OAI21_X1 U16770 ( .B1(n7198), .B2(n15146), .A(n15117), .ZN(n15122) );
  OAI21_X1 U16771 ( .B1(n15120), .B2(n15119), .A(n15118), .ZN(n15121) );
  AOI211_X1 U16772 ( .C1(n15124), .C2(n15123), .A(n15122), .B(n15121), .ZN(
        n15161) );
  INV_X1 U16773 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n15125) );
  AOI22_X1 U16774 ( .A1(n15155), .A2(n15161), .B1(n15125), .B2(n15153), .ZN(
        P2_U3454) );
  NAND2_X1 U16775 ( .A1(n15126), .A2(n15137), .ZN(n15127) );
  OAI211_X1 U16776 ( .C1(n15129), .C2(n15139), .A(n15128), .B(n15127), .ZN(
        n15130) );
  AOI211_X1 U16777 ( .C1(n15143), .C2(n15132), .A(n15131), .B(n15130), .ZN(
        n15162) );
  INV_X1 U16778 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15133) );
  AOI22_X1 U16779 ( .A1(n15155), .A2(n15162), .B1(n15133), .B2(n15153), .ZN(
        P2_U3457) );
  INV_X1 U16780 ( .A(n15140), .ZN(n15142) );
  AOI211_X1 U16781 ( .C1(n15137), .C2(n15136), .A(n15135), .B(n15134), .ZN(
        n15138) );
  OAI21_X1 U16782 ( .B1(n15140), .B2(n15139), .A(n15138), .ZN(n15141) );
  AOI21_X1 U16783 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n15163) );
  INV_X1 U16784 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n15144) );
  AOI22_X1 U16785 ( .A1(n15155), .A2(n15163), .B1(n15144), .B2(n15153), .ZN(
        P2_U3460) );
  OAI21_X1 U16786 ( .B1(n15147), .B2(n15146), .A(n15145), .ZN(n15150) );
  INV_X1 U16787 ( .A(n15148), .ZN(n15149) );
  AOI211_X1 U16788 ( .C1(n15152), .C2(n15151), .A(n15150), .B(n15149), .ZN(
        n15165) );
  AOI22_X1 U16789 ( .A1(n15155), .A2(n15165), .B1(n15154), .B2(n15153), .ZN(
        P2_U3463) );
  AOI22_X1 U16790 ( .A1(n15160), .A2(n15156), .B1(n8189), .B2(n15164), .ZN(
        P2_U3499) );
  AOI22_X1 U16791 ( .A1(n15160), .A2(n15157), .B1(n8279), .B2(n15164), .ZN(
        P2_U3504) );
  AOI22_X1 U16792 ( .A1(n15160), .A2(n15158), .B1(n10122), .B2(n15164), .ZN(
        P2_U3505) );
  AOI22_X1 U16793 ( .A1(n15160), .A2(n15159), .B1(n10123), .B2(n15164), .ZN(
        P2_U3506) );
  AOI22_X1 U16794 ( .A1(n15160), .A2(n15161), .B1(n10152), .B2(n15164), .ZN(
        P2_U3507) );
  AOI22_X1 U16795 ( .A1(n15160), .A2(n15162), .B1(n10179), .B2(n15164), .ZN(
        P2_U3508) );
  AOI22_X1 U16796 ( .A1(n15160), .A2(n15163), .B1(n10496), .B2(n15164), .ZN(
        P2_U3509) );
  AOI22_X1 U16797 ( .A1(n15160), .A2(n15165), .B1(n10497), .B2(n15164), .ZN(
        P2_U3510) );
  NOR2_X1 U16798 ( .A1(P3_U3897), .A2(n15293), .ZN(P3_U3150) );
  INV_X1 U16799 ( .A(n15166), .ZN(n15167) );
  NAND2_X1 U16800 ( .A1(n15167), .A2(n11079), .ZN(n15168) );
  AND2_X1 U16801 ( .A1(n15169), .A2(n15168), .ZN(n15186) );
  INV_X1 U16802 ( .A(n15170), .ZN(n15171) );
  OAI21_X1 U16803 ( .B1(n15172), .B2(n7178), .A(n15171), .ZN(n15179) );
  OR3_X1 U16804 ( .A1(n15175), .A2(n15174), .A3(n15173), .ZN(n15177) );
  AOI21_X1 U16805 ( .B1(n15192), .B2(n15177), .A(n15176), .ZN(n15178) );
  AOI211_X1 U16806 ( .C1(n15181), .C2(n15180), .A(n15179), .B(n15178), .ZN(
        n15185) );
  XNOR2_X1 U16807 ( .A(n15182), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n15183) );
  NAND2_X1 U16808 ( .A1(n15296), .A2(n15183), .ZN(n15184) );
  OAI211_X1 U16809 ( .C1(n15186), .C2(n15300), .A(n15185), .B(n15184), .ZN(
        P3_U3185) );
  AOI21_X1 U16810 ( .B1(n15189), .B2(n15188), .A(n15187), .ZN(n15204) );
  AND3_X1 U16811 ( .A1(n15192), .A2(n15191), .A3(n15190), .ZN(n15193) );
  OAI21_X1 U16812 ( .B1(n15210), .B2(n15193), .A(n15285), .ZN(n15194) );
  OAI21_X1 U16813 ( .B1(n15290), .B2(n15195), .A(n15194), .ZN(n15196) );
  AOI211_X1 U16814 ( .C1(P3_ADDR_REG_4__SCAN_IN), .C2(n15293), .A(n15197), .B(
        n15196), .ZN(n15203) );
  OAI21_X1 U16815 ( .B1(n15200), .B2(n15199), .A(n15198), .ZN(n15201) );
  NAND2_X1 U16816 ( .A1(n15296), .A2(n15201), .ZN(n15202) );
  OAI211_X1 U16817 ( .C1(n15204), .C2(n15300), .A(n15203), .B(n15202), .ZN(
        P3_U3186) );
  AOI21_X1 U16818 ( .B1(n15207), .B2(n15206), .A(n15205), .ZN(n15222) );
  INV_X1 U16819 ( .A(n15228), .ZN(n15212) );
  NOR3_X1 U16820 ( .A1(n15210), .A2(n15209), .A3(n15208), .ZN(n15211) );
  OAI21_X1 U16821 ( .B1(n15212), .B2(n15211), .A(n15285), .ZN(n15213) );
  OAI21_X1 U16822 ( .B1(n15290), .B2(n15214), .A(n15213), .ZN(n15215) );
  AOI211_X1 U16823 ( .C1(P3_ADDR_REG_5__SCAN_IN), .C2(n15293), .A(n15216), .B(
        n15215), .ZN(n15221) );
  OAI21_X1 U16824 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n15218), .A(n15217), .ZN(
        n15219) );
  NAND2_X1 U16825 ( .A1(n15296), .A2(n15219), .ZN(n15220) );
  OAI211_X1 U16826 ( .C1(n15222), .C2(n15300), .A(n15221), .B(n15220), .ZN(
        P3_U3187) );
  AOI21_X1 U16827 ( .B1(n15225), .B2(n15224), .A(n15223), .ZN(n15240) );
  AND3_X1 U16828 ( .A1(n15228), .A2(n15227), .A3(n15226), .ZN(n15229) );
  OAI21_X1 U16829 ( .B1(n15245), .B2(n15229), .A(n15285), .ZN(n15230) );
  OAI21_X1 U16830 ( .B1(n15290), .B2(n15231), .A(n15230), .ZN(n15232) );
  AOI211_X1 U16831 ( .C1(P3_ADDR_REG_6__SCAN_IN), .C2(n15293), .A(n15233), .B(
        n15232), .ZN(n15239) );
  OAI21_X1 U16832 ( .B1(n15236), .B2(n15235), .A(n15234), .ZN(n15237) );
  NAND2_X1 U16833 ( .A1(n15296), .A2(n15237), .ZN(n15238) );
  OAI211_X1 U16834 ( .C1(n15240), .C2(n15300), .A(n15239), .B(n15238), .ZN(
        P3_U3188) );
  AOI21_X1 U16835 ( .B1(n11099), .B2(n15242), .A(n15241), .ZN(n15257) );
  INV_X1 U16836 ( .A(n15265), .ZN(n15247) );
  NOR3_X1 U16837 ( .A1(n15245), .A2(n15244), .A3(n15243), .ZN(n15246) );
  OAI21_X1 U16838 ( .B1(n15247), .B2(n15246), .A(n15285), .ZN(n15248) );
  OAI21_X1 U16839 ( .B1(n15290), .B2(n15249), .A(n15248), .ZN(n15250) );
  AOI211_X1 U16840 ( .C1(P3_ADDR_REG_7__SCAN_IN), .C2(n15293), .A(n15251), .B(
        n15250), .ZN(n15256) );
  OAI21_X1 U16841 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n15253), .A(n15252), .ZN(
        n15254) );
  NAND2_X1 U16842 ( .A1(n15296), .A2(n15254), .ZN(n15255) );
  OAI211_X1 U16843 ( .C1(n15257), .C2(n15300), .A(n15256), .B(n15255), .ZN(
        P3_U3189) );
  INV_X1 U16844 ( .A(n15259), .ZN(n15260) );
  AOI21_X1 U16845 ( .B1(n15262), .B2(n15261), .A(n15260), .ZN(n15277) );
  AND3_X1 U16846 ( .A1(n15265), .A2(n15264), .A3(n15263), .ZN(n15266) );
  OAI21_X1 U16847 ( .B1(n15284), .B2(n15266), .A(n15285), .ZN(n15267) );
  OAI21_X1 U16848 ( .B1(n15290), .B2(n15268), .A(n15267), .ZN(n15269) );
  AOI211_X1 U16849 ( .C1(P3_ADDR_REG_8__SCAN_IN), .C2(n15293), .A(n15270), .B(
        n15269), .ZN(n15276) );
  OAI21_X1 U16850 ( .B1(n15273), .B2(n15272), .A(n15271), .ZN(n15274) );
  NAND2_X1 U16851 ( .A1(n15274), .A2(n15296), .ZN(n15275) );
  OAI211_X1 U16852 ( .C1(n15277), .C2(n15300), .A(n15276), .B(n15275), .ZN(
        P3_U3190) );
  AOI21_X1 U16853 ( .B1(n15280), .B2(n15279), .A(n15278), .ZN(n15301) );
  INV_X1 U16854 ( .A(n15281), .ZN(n15287) );
  NOR3_X1 U16855 ( .A1(n15284), .A2(n15283), .A3(n15282), .ZN(n15286) );
  OAI21_X1 U16856 ( .B1(n15287), .B2(n15286), .A(n15285), .ZN(n15288) );
  OAI21_X1 U16857 ( .B1(n15290), .B2(n15289), .A(n15288), .ZN(n15291) );
  AOI211_X1 U16858 ( .C1(P3_ADDR_REG_9__SCAN_IN), .C2(n15293), .A(n15292), .B(
        n15291), .ZN(n15299) );
  OAI21_X1 U16859 ( .B1(n15295), .B2(P3_REG1_REG_9__SCAN_IN), .A(n15294), .ZN(
        n15297) );
  NAND2_X1 U16860 ( .A1(n15297), .A2(n15296), .ZN(n15298) );
  OAI211_X1 U16861 ( .C1(n15301), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        P3_U3191) );
  XNOR2_X1 U16862 ( .A(n15302), .B(n15306), .ZN(n15408) );
  AOI22_X1 U16863 ( .A1(n15304), .A2(n15319), .B1(n15321), .B2(n15303), .ZN(
        n15309) );
  OAI211_X1 U16864 ( .C1(n15307), .C2(n15306), .A(n15305), .B(n15323), .ZN(
        n15308) );
  OAI211_X1 U16865 ( .C1(n15408), .C2(n15328), .A(n15309), .B(n15308), .ZN(
        n15410) );
  INV_X1 U16866 ( .A(n15410), .ZN(n15310) );
  OAI21_X1 U16867 ( .B1(n15357), .B2(n15408), .A(n15310), .ZN(n15314) );
  OAI22_X1 U16868 ( .A1(n15312), .A2(n15405), .B1(n15311), .B2(n15369), .ZN(
        n15313) );
  AOI21_X1 U16869 ( .B1(n15314), .B2(n15369), .A(n15313), .ZN(n15315) );
  OAI21_X1 U16870 ( .B1(n15317), .B2(n15316), .A(n15315), .ZN(P3_U3223) );
  XOR2_X1 U16871 ( .A(n15318), .B(n7919), .Z(n15329) );
  INV_X1 U16872 ( .A(n15329), .ZN(n15378) );
  AOI22_X1 U16873 ( .A1(n15321), .A2(n10825), .B1(n15320), .B2(n15319), .ZN(
        n15327) );
  INV_X1 U16874 ( .A(n7919), .ZN(n15324) );
  OAI211_X1 U16875 ( .C1(n15325), .C2(n15324), .A(n15323), .B(n15322), .ZN(
        n15326) );
  OAI211_X1 U16876 ( .C1(n15329), .C2(n15328), .A(n15327), .B(n15326), .ZN(
        n15376) );
  AOI21_X1 U16877 ( .B1(n15330), .B2(n15378), .A(n15376), .ZN(n15335) );
  NOR2_X1 U16878 ( .A1(n15331), .A2(n15406), .ZN(n15377) );
  AOI22_X1 U16879 ( .A1(n15333), .A2(n15377), .B1(n15365), .B2(n15332), .ZN(
        n15334) );
  OAI221_X1 U16880 ( .B1(n15371), .B2(n15335), .C1(n15369), .C2(n11079), .A(
        n15334), .ZN(P3_U3230) );
  OAI21_X1 U16881 ( .B1(n15337), .B2(n15345), .A(n15336), .ZN(n15375) );
  OAI22_X1 U16882 ( .A1(n15341), .A2(n15340), .B1(n15339), .B2(n15338), .ZN(
        n15351) );
  NAND2_X1 U16883 ( .A1(n15346), .A2(n15344), .ZN(n15343) );
  NAND2_X1 U16884 ( .A1(n15343), .A2(n15342), .ZN(n15349) );
  NAND3_X1 U16885 ( .A1(n15346), .A2(n15345), .A3(n15344), .ZN(n15348) );
  AOI21_X1 U16886 ( .B1(n15349), .B2(n15348), .A(n15347), .ZN(n15350) );
  AOI211_X1 U16887 ( .C1(n15352), .C2(n15375), .A(n15351), .B(n15350), .ZN(
        n15353) );
  INV_X1 U16888 ( .A(n15353), .ZN(n15373) );
  INV_X1 U16889 ( .A(n15375), .ZN(n15358) );
  NOR2_X1 U16890 ( .A1(n15354), .A2(n15406), .ZN(n15374) );
  INV_X1 U16891 ( .A(n15374), .ZN(n15355) );
  OAI22_X1 U16892 ( .A1(n15358), .A2(n15357), .B1(n15356), .B2(n15355), .ZN(
        n15359) );
  AOI211_X1 U16893 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15365), .A(n15373), .B(
        n15359), .ZN(n15360) );
  AOI22_X1 U16894 ( .A1(n15371), .A2(n10600), .B1(n15360), .B2(n15369), .ZN(
        P3_U3231) );
  INV_X1 U16895 ( .A(n15361), .ZN(n15362) );
  AOI21_X1 U16896 ( .B1(n15364), .B2(n15363), .A(n15362), .ZN(n15370) );
  AOI22_X1 U16897 ( .A1(n15367), .A2(n15366), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n15365), .ZN(n15368) );
  OAI221_X1 U16898 ( .B1(n15371), .B2(n15370), .C1(n15369), .C2(n10593), .A(
        n15368), .ZN(P3_U3232) );
  AOI22_X1 U16899 ( .A1(n15412), .A2(n7516), .B1(n15372), .B2(n15411), .ZN(
        P3_U3393) );
  AOI211_X1 U16900 ( .C1(n15400), .C2(n15375), .A(n15374), .B(n15373), .ZN(
        n15414) );
  AOI22_X1 U16901 ( .A1(n15412), .A2(n7531), .B1(n15414), .B2(n15411), .ZN(
        P3_U3396) );
  AOI211_X1 U16902 ( .C1(n15378), .C2(n15400), .A(n15377), .B(n15376), .ZN(
        n15415) );
  AOI22_X1 U16903 ( .A1(n15412), .A2(n7541), .B1(n15415), .B2(n15411), .ZN(
        P3_U3399) );
  INV_X1 U16904 ( .A(n15379), .ZN(n15380) );
  AOI211_X1 U16905 ( .C1(n15400), .C2(n15382), .A(n15381), .B(n15380), .ZN(
        n15416) );
  AOI22_X1 U16906 ( .A1(n15412), .A2(n7557), .B1(n15416), .B2(n15411), .ZN(
        P3_U3402) );
  INV_X1 U16907 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15386) );
  AOI211_X1 U16908 ( .C1(n15385), .C2(n15400), .A(n15384), .B(n15383), .ZN(
        n15417) );
  AOI22_X1 U16909 ( .A1(n15412), .A2(n15386), .B1(n15417), .B2(n15411), .ZN(
        P3_U3405) );
  INV_X1 U16910 ( .A(n15387), .ZN(n15390) );
  AOI211_X1 U16911 ( .C1(n15390), .C2(n15400), .A(n15389), .B(n15388), .ZN(
        n15418) );
  AOI22_X1 U16912 ( .A1(n15412), .A2(n7591), .B1(n15418), .B2(n15411), .ZN(
        P3_U3408) );
  AOI211_X1 U16913 ( .C1(n15393), .C2(n15400), .A(n15392), .B(n15391), .ZN(
        n15419) );
  AOI22_X1 U16914 ( .A1(n15412), .A2(n7605), .B1(n15419), .B2(n15411), .ZN(
        P3_U3411) );
  INV_X1 U16915 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15398) );
  AOI21_X1 U16916 ( .B1(n15395), .B2(n15400), .A(n15394), .ZN(n15396) );
  AND2_X1 U16917 ( .A1(n15397), .A2(n15396), .ZN(n15420) );
  AOI22_X1 U16918 ( .A1(n15412), .A2(n15398), .B1(n15420), .B2(n15411), .ZN(
        P3_U3414) );
  INV_X1 U16919 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15404) );
  AOI21_X1 U16920 ( .B1(n15401), .B2(n15400), .A(n15399), .ZN(n15402) );
  AND2_X1 U16921 ( .A1(n15403), .A2(n15402), .ZN(n15421) );
  AOI22_X1 U16922 ( .A1(n15412), .A2(n15404), .B1(n15421), .B2(n15411), .ZN(
        P3_U3417) );
  OAI22_X1 U16923 ( .A1(n15408), .A2(n15407), .B1(n15406), .B2(n15405), .ZN(
        n15409) );
  NOR2_X1 U16924 ( .A1(n15410), .A2(n15409), .ZN(n15423) );
  AOI22_X1 U16925 ( .A1(n15412), .A2(n7657), .B1(n15423), .B2(n15411), .ZN(
        P3_U3420) );
  AOI22_X1 U16926 ( .A1(n15424), .A2(n15414), .B1(n15413), .B2(n8836), .ZN(
        P3_U3461) );
  AOI22_X1 U16927 ( .A1(n15424), .A2(n15415), .B1(n11078), .B2(n8836), .ZN(
        P3_U3462) );
  AOI22_X1 U16928 ( .A1(n15424), .A2(n15416), .B1(n11083), .B2(n8836), .ZN(
        P3_U3463) );
  AOI22_X1 U16929 ( .A1(n15424), .A2(n15417), .B1(n11088), .B2(n8836), .ZN(
        P3_U3464) );
  AOI22_X1 U16930 ( .A1(n15424), .A2(n15418), .B1(n11092), .B2(n8836), .ZN(
        P3_U3465) );
  AOI22_X1 U16931 ( .A1(n15424), .A2(n15419), .B1(n11098), .B2(n8836), .ZN(
        P3_U3466) );
  AOI22_X1 U16932 ( .A1(n15424), .A2(n15420), .B1(n11133), .B2(n8836), .ZN(
        P3_U3467) );
  AOI22_X1 U16933 ( .A1(n15424), .A2(n15421), .B1(n11107), .B2(n8836), .ZN(
        P3_U3468) );
  AOI22_X1 U16934 ( .A1(n15424), .A2(n15423), .B1(n15422), .B2(n8836), .ZN(
        P3_U3469) );
  XOR2_X1 U16935 ( .A(n15426), .B(n15425), .Z(SUB_1596_U59) );
  XNOR2_X1 U16936 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n15427), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16937 ( .B1(n15429), .B2(n15428), .A(n15438), .ZN(SUB_1596_U53) );
  XOR2_X1 U16938 ( .A(n15431), .B(n15430), .Z(SUB_1596_U56) );
  OAI21_X1 U16939 ( .B1(n15434), .B2(n15433), .A(n15432), .ZN(n15436) );
  XOR2_X1 U16940 ( .A(n15436), .B(n15435), .Z(SUB_1596_U60) );
  XOR2_X1 U16941 ( .A(n15438), .B(n15437), .Z(SUB_1596_U5) );
  INV_X2 U7391 ( .A(n8213), .ZN(n8658) );
  INV_X1 U7299 ( .A(n12227), .ZN(n12219) );
  CLKBUF_X1 U7319 ( .A(n9393), .Z(n9500) );
  CLKBUF_X1 U7483 ( .A(n9060), .Z(n14721) );
  CLKBUF_X1 U7527 ( .A(n7530), .Z(n6551) );
  NAND2_X2 U8070 ( .A1(n12769), .A2(n12771), .ZN(n7558) );
  CLKBUF_X2 U9255 ( .A(n11119), .Z(n6552) );
  CLKBUF_X1 U9475 ( .A(n9528), .Z(n6720) );
endmodule

