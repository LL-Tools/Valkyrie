

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025;

  XNOR2_X1 U11164 ( .A(n14601), .B(n14602), .ZN(n15498) );
  OR2_X1 U11165 ( .A1(n13621), .A2(n13620), .ZN(n13809) );
  AND2_X1 U11166 ( .A1(n9794), .A2(n13361), .ZN(n11525) );
  AND2_X1 U11167 ( .A1(n12831), .A2(n10013), .ZN(n10387) );
  AND2_X1 U11169 ( .A1(n14686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10439) );
  AND2_X1 U11170 ( .A1(n14685), .A2(n16039), .ZN(n10455) );
  AND2_X1 U11171 ( .A1(n9745), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10528) );
  AND2_X1 U11172 ( .A1(n9736), .A2(n16039), .ZN(n14503) );
  BUF_X2 U11173 ( .A(n17461), .Z(n17479) );
  CLKBUF_X2 U11174 ( .A(n12265), .Z(n9722) );
  CLKBUF_X1 U11175 ( .A(n11286), .Z(n12081) );
  CLKBUF_X1 U11176 ( .A(n11701), .Z(n12056) );
  CLKBUF_X1 U11177 ( .A(n11306), .Z(n11739) );
  CLKBUF_X1 U11178 ( .A(n11261), .Z(n12076) );
  CLKBUF_X2 U11179 ( .A(n11718), .Z(n9747) );
  CLKBUF_X2 U11181 ( .A(n11508), .Z(n12475) );
  BUF_X1 U11182 ( .A(n12315), .Z(n17439) );
  INV_X1 U11183 ( .A(n10151), .ZN(n9734) );
  NOR2_X1 U11184 ( .A1(n11428), .A2(n11356), .ZN(n13135) );
  NAND2_X1 U11185 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18921) );
  INV_X2 U11186 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n19096) );
  AND4_X1 U11187 ( .A1(n11339), .A2(n11338), .A3(n11337), .A4(n11336), .ZN(
        n11345) );
  OR2_X1 U11188 ( .A1(n11260), .A2(n11259), .ZN(n11291) );
  INV_X1 U11189 ( .A(n10980), .ZN(n16683) );
  AND2_X1 U11190 ( .A1(n11230), .A2(n11232), .ZN(n11455) );
  AND2_X1 U11191 ( .A1(n11233), .A2(n11232), .ZN(n11508) );
  AND2_X2 U11192 ( .A1(n12903), .A2(n11230), .ZN(n11261) );
  NAND2_X1 U11193 ( .A1(n10237), .A2(n10236), .ZN(n13890) );
  CLKBUF_X1 U11194 ( .A(n20673), .Z(n9720) );
  NOR2_X1 U11195 ( .A1(n20632), .A2(n20691), .ZN(n20673) );
  CLKBUF_X1 U11196 ( .A(n18603), .Z(n9721) );
  NOR2_X1 U11197 ( .A1(n18700), .A2(n18561), .ZN(n18603) );
  AOI21_X1 U11198 ( .B1(n19880), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n9740), .ZN(n10407) );
  INV_X1 U11199 ( .A(n10854), .ZN(n11205) );
  BUF_X1 U11200 ( .A(n13846), .Z(n14508) );
  AND2_X1 U11201 ( .A1(n9746), .A2(n16039), .ZN(n10477) );
  AOI21_X1 U11202 ( .B1(n10344), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10345), .ZN(n10863) );
  INV_X1 U11203 ( .A(n11821), .ZN(n12513) );
  AND4_X1 U11204 ( .A1(n11277), .A2(n11276), .A3(n11275), .A4(n11274), .ZN(
        n11278) );
  AND3_X1 U11205 ( .A1(n10305), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10980), 
        .ZN(n14570) );
  NAND2_X1 U11206 ( .A1(n10054), .A2(n10052), .ZN(n10980) );
  NAND2_X1 U11207 ( .A1(n13993), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13992) );
  INV_X1 U11209 ( .A(n10166), .ZN(n17409) );
  NAND2_X1 U11210 ( .A1(n19109), .A2(n19103), .ZN(n17188) );
  NAND2_X1 U11211 ( .A1(n11428), .A2(n13479), .ZN(n13172) );
  INV_X1 U11212 ( .A(n11601), .ZN(n15097) );
  INV_X1 U11213 ( .A(n13479), .ZN(n13292) );
  NOR2_X1 U11214 ( .A1(n13982), .A2(n13981), .ZN(n14092) );
  NAND2_X1 U11215 ( .A1(n10300), .A2(n10979), .ZN(n14444) );
  INV_X1 U11217 ( .A(n18947), .ZN(n18930) );
  INV_X1 U11218 ( .A(n14308), .ZN(n14341) );
  NAND2_X1 U11219 ( .A1(n15089), .A2(n15090), .ZN(n15061) );
  AND2_X1 U11220 ( .A1(n15307), .A2(n15306), .ZN(n15309) );
  NAND2_X1 U11221 ( .A1(n11781), .A2(n11780), .ZN(n12607) );
  INV_X1 U11222 ( .A(n10973), .ZN(n13430) );
  INV_X1 U11223 ( .A(n16211), .ZN(n18485) );
  INV_X1 U11224 ( .A(n18016), .ZN(n17943) );
  INV_X1 U11225 ( .A(n19132), .ZN(n17729) );
  INV_X1 U11226 ( .A(n20221), .ZN(n20277) );
  INV_X1 U11227 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20616) );
  AOI211_X1 U11228 ( .C1(n15922), .C2(n16635), .A(n15921), .B(n15920), .ZN(
        n15928) );
  AOI211_X1 U11229 ( .C1(n19220), .C2(n16635), .A(n15932), .B(n15931), .ZN(
        n15935) );
  INV_X4 U11231 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16647) );
  NOR2_X2 U11232 ( .A1(n15046), .A2(n15186), .ZN(n15010) );
  AND2_X4 U11233 ( .A1(n10211), .A2(n10210), .ZN(n10267) );
  INV_X2 U11234 ( .A(n17670), .ZN(n12367) );
  NAND2_X2 U11235 ( .A1(n11427), .A2(n11426), .ZN(n13659) );
  NOR2_X2 U11236 ( .A1(n13553), .A2(n13555), .ZN(n13554) );
  NAND2_X2 U11237 ( .A1(n15503), .A2(n14577), .ZN(n14601) );
  AND3_X2 U11238 ( .A1(n18959), .A2(n19133), .A3(n16135), .ZN(n16214) );
  NOR2_X2 U11239 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11234) );
  AND2_X1 U11240 ( .A1(n11233), .A2(n12903), .ZN(n11718) );
  NOR2_X4 U11241 ( .A1(n10356), .A2(n16008), .ZN(n19910) );
  AOI21_X2 U11242 ( .B1(n15918), .B2(n16624), .A(n15937), .ZN(n15930) );
  XNOR2_X2 U11243 ( .A(n10585), .B(n10961), .ZN(n16536) );
  NAND2_X2 U11244 ( .A1(n10584), .A2(n13520), .ZN(n10585) );
  NAND2_X2 U11245 ( .A1(n10622), .A2(n10846), .ZN(n10838) );
  NOR2_X1 U11246 ( .A1(n12146), .A2(n12145), .ZN(n12265) );
  NOR2_X2 U11247 ( .A1(n10386), .A2(n10385), .ZN(n10548) );
  XNOR2_X2 U11248 ( .A(n9859), .B(n11435), .ZN(n13284) );
  NOR2_X2 U11249 ( .A1(n15493), .A2(n15492), .ZN(n15491) );
  AND2_X2 U11250 ( .A1(n11224), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11230) );
  INV_X1 U11251 ( .A(n12253), .ZN(n9724) );
  XNOR2_X1 U11252 ( .A(n9780), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14458) );
  OR2_X1 U11253 ( .A1(n15633), .A2(n9775), .ZN(n15621) );
  CLKBUF_X1 U11255 ( .A(n14773), .Z(n14774) );
  NAND2_X1 U11256 ( .A1(n11587), .A2(n16315), .ZN(n14005) );
  AND2_X1 U11257 ( .A1(n10171), .A2(n9832), .ZN(n15558) );
  NAND2_X1 U11258 ( .A1(n13907), .A2(n9815), .ZN(n15525) );
  AND2_X1 U11259 ( .A1(n10575), .A2(n10574), .ZN(n10588) );
  OR2_X1 U11260 ( .A1(n13271), .A2(n13187), .ZN(n13399) );
  INV_X2 U11261 ( .A(n18162), .ZN(n18119) );
  AND2_X2 U11262 ( .A1(n10388), .A2(n10384), .ZN(n10547) );
  AND2_X2 U11263 ( .A1(n10388), .A2(n10387), .ZN(n10549) );
  BUF_X1 U11264 ( .A(n11765), .Z(n9748) );
  NAND2_X1 U11265 ( .A1(n13279), .A2(n11434), .ZN(n11475) );
  NAND2_X1 U11266 ( .A1(n13428), .A2(n13427), .ZN(n19387) );
  OR2_X1 U11267 ( .A1(n13412), .A2(n13411), .ZN(n13414) );
  NOR2_X1 U11268 ( .A1(n15360), .A2(n15630), .ZN(n15363) );
  NAND2_X1 U11269 ( .A1(n11349), .A2(n11291), .ZN(n12515) );
  NOR2_X1 U11270 ( .A1(n18496), .A2(n18516), .ZN(n12364) );
  INV_X4 U11271 ( .A(n10855), .ZN(n9725) );
  NAND2_X1 U11273 ( .A1(n18485), .A2(n17647), .ZN(n12345) );
  INV_X4 U11274 ( .A(n9739), .ZN(n19514) );
  NAND2_X1 U11275 ( .A1(n11360), .A2(n11291), .ZN(n12791) );
  CLKBUF_X2 U11276 ( .A(n10996), .Z(n14442) );
  INV_X2 U11277 ( .A(n11356), .ZN(n13034) );
  INV_X1 U11278 ( .A(n13472), .ZN(n13282) );
  AND4_X1 U11279 ( .A1(n11265), .A2(n11264), .A3(n11263), .A4(n11262), .ZN(
        n11281) );
  CLKBUF_X2 U11280 ( .A(n12188), .Z(n17355) );
  BUF_X2 U11281 ( .A(n11552), .Z(n9730) );
  BUF_X2 U11282 ( .A(n12318), .Z(n17311) );
  AND2_X2 U11283 ( .A1(n16033), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10563) );
  CLKBUF_X2 U11284 ( .A(n11298), .Z(n12051) );
  CLKBUF_X2 U11285 ( .A(n11299), .Z(n12057) );
  CLKBUF_X2 U11286 ( .A(n11455), .Z(n12494) );
  BUF_X2 U11287 ( .A(n10187), .Z(n9738) );
  INV_X4 U11288 ( .A(n9777), .ZN(n17454) );
  BUF_X2 U11289 ( .A(n10188), .Z(n16033) );
  CLKBUF_X2 U11290 ( .A(n11297), .Z(n12050) );
  OR2_X1 U11291 ( .A1(n19085), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12140) );
  OR2_X1 U11292 ( .A1(n12142), .A2(n18921), .ZN(n9777) );
  INV_X1 U11293 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9935) );
  AOI211_X1 U11294 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n15833), .A(
        n15822), .B(n15821), .ZN(n15823) );
  AOI211_X1 U11295 ( .C1(n15800), .C2(n16624), .A(n15799), .B(n15798), .ZN(
        n15801) );
  NAND2_X1 U11296 ( .A1(n9923), .A2(n15621), .ZN(n15820) );
  INV_X1 U11297 ( .A(n10060), .ZN(n15808) );
  AOI211_X1 U11298 ( .C1(n14458), .C2(n19475), .A(n14439), .B(n14438), .ZN(
        n14440) );
  OR2_X1 U11299 ( .A1(n15812), .A2(n19500), .ZN(n10051) );
  NAND2_X1 U11300 ( .A1(n10058), .A2(n9855), .ZN(n10060) );
  AOI22_X1 U11301 ( .A1(n15607), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n10740), .B2(n10739), .ZN(n10742) );
  INV_X1 U11302 ( .A(n15620), .ZN(n9924) );
  CLKBUF_X1 U11303 ( .A(n15633), .Z(n15845) );
  AND2_X1 U11304 ( .A1(n9905), .A2(n9904), .ZN(n11190) );
  OAI21_X1 U11305 ( .B1(n9874), .B2(n9873), .A(n10160), .ZN(n15011) );
  OAI21_X1 U11306 ( .B1(n12488), .B2(n14720), .A(n14708), .ZN(n14947) );
  OR3_X1 U11307 ( .A1(n14989), .A2(n15169), .A3(n15001), .ZN(n10159) );
  AND2_X1 U11308 ( .A1(n14841), .A2(n14825), .ZN(n14915) );
  AND2_X1 U11309 ( .A1(n14923), .A2(n14922), .ZN(n16233) );
  OR2_X1 U11310 ( .A1(n14923), .A2(n14839), .ZN(n14916) );
  NAND2_X1 U11311 ( .A1(n14375), .A2(n15054), .ZN(n10133) );
  NAND2_X1 U11312 ( .A1(n10650), .A2(n9830), .ZN(n15645) );
  NOR2_X1 U11313 ( .A1(n15804), .A2(n10047), .ZN(n10046) );
  OR2_X1 U11314 ( .A1(n15346), .A2(n15345), .ZN(n15797) );
  NAND2_X1 U11315 ( .A1(n10135), .A2(n10137), .ZN(n15089) );
  NOR3_X1 U11316 ( .A1(n15379), .A2(n10095), .A3(n10094), .ZN(n15346) );
  NAND2_X1 U11317 ( .A1(n10835), .A2(n10834), .ZN(n16533) );
  NAND2_X1 U11318 ( .A1(n14005), .A2(n11593), .ZN(n9871) );
  OR2_X1 U11319 ( .A1(n10850), .A2(n16609), .ZN(n10851) );
  OR2_X1 U11320 ( .A1(n16532), .A2(n10840), .ZN(n10841) );
  OR2_X1 U11321 ( .A1(n10846), .A2(n11020), .ZN(n10850) );
  AND2_X1 U11322 ( .A1(n10725), .A2(n10735), .ZN(n14424) );
  NOR2_X1 U11323 ( .A1(n9870), .A2(n9799), .ZN(n9869) );
  NOR2_X1 U11324 ( .A1(n15109), .A2(n15111), .ZN(n11606) );
  OR2_X1 U11325 ( .A1(n18040), .A2(n18265), .ZN(n17967) );
  OR2_X2 U11326 ( .A1(n13399), .A2(n13398), .ZN(n13461) );
  NOR2_X2 U11327 ( .A1(n19851), .A2(n19758), .ZN(n20046) );
  OR2_X1 U11328 ( .A1(n11601), .A2(n15231), .ZN(n16298) );
  AND2_X1 U11329 ( .A1(n10620), .A2(n10619), .ZN(n10840) );
  NAND2_X1 U11330 ( .A1(n9788), .A2(n11805), .ZN(n13144) );
  AOI21_X1 U11331 ( .B1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n19702), .A(
        n10409), .ZN(n10425) );
  OAI21_X1 U11332 ( .B1(n13062), .B2(n13063), .A(n13007), .ZN(n19549) );
  XNOR2_X1 U11333 ( .A(n11576), .B(n11575), .ZN(n11835) );
  OR2_X1 U11334 ( .A1(n10608), .A2(n10607), .ZN(n10620) );
  NAND2_X1 U11335 ( .A1(n11562), .A2(n11561), .ZN(n11576) );
  NAND2_X1 U11336 ( .A1(n13105), .A2(n13104), .ZN(n13110) );
  OR2_X1 U11337 ( .A1(n13006), .A2(n10085), .ZN(n10083) );
  XNOR2_X1 U11338 ( .A(n9877), .B(n11547), .ZN(n11814) );
  NAND2_X1 U11339 ( .A1(n13004), .A2(n13003), .ZN(n13063) );
  NAND2_X1 U11340 ( .A1(n18964), .A2(n19128), .ZN(n16819) );
  INV_X1 U11341 ( .A(n11525), .ZN(n11523) );
  AND2_X1 U11342 ( .A1(n13099), .A2(n13098), .ZN(n13105) );
  INV_X1 U11343 ( .A(n10548), .ZN(n19570) );
  OR2_X1 U11344 ( .A1(n12948), .A2(n12947), .ZN(n13004) );
  OR2_X1 U11345 ( .A1(n13005), .A2(n13001), .ZN(n13002) );
  AND2_X1 U11346 ( .A1(n13091), .A2(n13067), .ZN(n13099) );
  NAND2_X1 U11347 ( .A1(n13000), .A2(n12999), .ZN(n13005) );
  AND2_X1 U11348 ( .A1(n15992), .A2(n9817), .ZN(n16595) );
  CLKBUF_X1 U11349 ( .A(n14941), .Z(n16282) );
  CLKBUF_X1 U11350 ( .A(n12543), .Z(n16284) );
  XNOR2_X1 U11351 ( .A(n11475), .B(n20962), .ZN(n13456) );
  INV_X1 U11352 ( .A(n10382), .ZN(n10388) );
  NOR2_X1 U11353 ( .A1(n10690), .A2(n10662), .ZN(n9937) );
  NOR2_X1 U11354 ( .A1(n13578), .A2(n13034), .ZN(n20574) );
  NAND2_X1 U11355 ( .A1(n11773), .A2(n11774), .ZN(n11477) );
  NAND2_X1 U11356 ( .A1(n11776), .A2(n11393), .ZN(n11773) );
  NAND2_X1 U11357 ( .A1(n18081), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18080) );
  OAI21_X1 U11358 ( .B1(n11449), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11462), 
        .ZN(n11479) );
  AND2_X1 U11359 ( .A1(n10363), .A2(n19481), .ZN(n10364) );
  CLKBUF_X1 U11360 ( .A(n12610), .Z(n13629) );
  NAND2_X1 U11361 ( .A1(n13139), .A2(n13138), .ZN(n20282) );
  XNOR2_X1 U11362 ( .A(n10355), .B(n10362), .ZN(n12831) );
  INV_X2 U11363 ( .A(n17703), .ZN(n17721) );
  OR2_X1 U11364 ( .A1(n11447), .A2(n11446), .ZN(n11448) );
  NAND2_X1 U11365 ( .A1(n11447), .A2(n11446), .ZN(n12952) );
  OR2_X1 U11366 ( .A1(n11777), .A2(n11468), .ZN(n11774) );
  AND2_X1 U11367 ( .A1(n10352), .A2(n10349), .ZN(n19481) );
  OR2_X1 U11368 ( .A1(n13075), .A2(n11790), .ZN(n11791) );
  INV_X2 U11369 ( .A(n15537), .ZN(n9726) );
  NAND2_X1 U11370 ( .A1(n11440), .A2(n11439), .ZN(n11447) );
  AND2_X1 U11371 ( .A1(n10099), .A2(n10865), .ZN(n10098) );
  NAND2_X1 U11372 ( .A1(n11467), .A2(n11466), .ZN(n11777) );
  CLKBUF_X1 U11373 ( .A(n10346), .Z(n10352) );
  NAND2_X1 U11374 ( .A1(n11787), .A2(n10118), .ZN(n11467) );
  XNOR2_X1 U11375 ( .A(n10862), .B(n10863), .ZN(n10861) );
  OR2_X1 U11376 ( .A1(n13345), .A2(n9952), .ZN(n13621) );
  NAND2_X1 U11377 ( .A1(n10343), .A2(n10342), .ZN(n10862) );
  NOR2_X1 U11378 ( .A1(n18117), .A2(n18116), .ZN(n18115) );
  OAI21_X1 U11379 ( .B1(n11441), .B2(n12894), .A(n11445), .ZN(n11446) );
  NAND2_X1 U11380 ( .A1(n10111), .A2(n10112), .ZN(n11410) );
  NAND2_X1 U11381 ( .A1(n13414), .A2(n10992), .ZN(n11000) );
  INV_X2 U11382 ( .A(n9741), .ZN(n10936) );
  XNOR2_X1 U11383 ( .A(n10065), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18117) );
  AND2_X1 U11384 ( .A1(n15363), .A2(n9994), .ZN(n15587) );
  NAND4_X2 U11385 ( .A1(n9779), .A2(n10633), .A3(n11199), .A4(n10579), .ZN(
        n10725) );
  CLKBUF_X1 U11386 ( .A(n12671), .Z(n12750) );
  NAND2_X1 U11387 ( .A1(n12958), .A2(n12957), .ZN(n12956) );
  AND2_X1 U11388 ( .A1(n10578), .A2(n10580), .ZN(n9940) );
  AND2_X1 U11389 ( .A1(n10341), .A2(n10340), .ZN(n10343) );
  AOI21_X1 U11390 ( .B1(n11365), .B2(n10114), .A(n10113), .ZN(n10112) );
  OR2_X1 U11391 ( .A1(n10978), .A2(n10977), .ZN(n12958) );
  OAI211_X1 U11392 ( .C1(n11379), .C2(n11378), .A(n11377), .B(n11376), .ZN(
        n11408) );
  AND2_X1 U11393 ( .A1(n10317), .A2(n10316), .ZN(n10318) );
  AND2_X1 U11394 ( .A1(n10331), .A2(n10330), .ZN(n10332) );
  NAND2_X1 U11395 ( .A1(n11170), .A2(n12725), .ZN(n10306) );
  INV_X1 U11396 ( .A(n11205), .ZN(n14432) );
  AND2_X1 U11397 ( .A1(n12355), .A2(n12340), .ZN(n12417) );
  AND2_X1 U11398 ( .A1(n10282), .A2(n10281), .ZN(n11170) );
  INV_X2 U11399 ( .A(n10855), .ZN(n10339) );
  INV_X2 U11400 ( .A(n11038), .ZN(n11215) );
  NAND3_X1 U11401 ( .A1(n10946), .A2(n10043), .A3(n10042), .ZN(n10855) );
  NOR2_X1 U11402 ( .A1(n17665), .A2(n12367), .ZN(n12372) );
  AND2_X1 U11403 ( .A1(n14342), .A2(n11674), .ZN(n12779) );
  INV_X1 U11404 ( .A(n11038), .ZN(n9727) );
  NAND2_X1 U11405 ( .A1(n12787), .A2(n11353), .ZN(n13044) );
  NAND2_X1 U11406 ( .A1(n13172), .A2(n13438), .ZN(n14342) );
  AND3_X1 U11407 ( .A1(n13495), .A2(n13135), .A3(n13297), .ZN(n12787) );
  OR2_X1 U11408 ( .A1(n9862), .A2(n13172), .ZN(n13052) );
  AND2_X1 U11409 ( .A1(n13481), .A2(n12777), .ZN(n11357) );
  INV_X1 U11410 ( .A(n10285), .ZN(n10946) );
  NAND2_X1 U11411 ( .A1(n14308), .A2(n14313), .ZN(n14332) );
  AND2_X1 U11412 ( .A1(n10298), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U11413 ( .A1(n10976), .A2(n9740), .ZN(n11140) );
  INV_X1 U11414 ( .A(n12343), .ZN(n18510) );
  NAND2_X1 U11415 ( .A1(n9792), .A2(n9758), .ZN(n17670) );
  INV_X1 U11416 ( .A(n17661), .ZN(n12373) );
  NAND2_X1 U11417 ( .A1(n13292), .A2(n13472), .ZN(n20700) );
  BUF_X2 U11418 ( .A(n16683), .Z(n9739) );
  NOR2_X1 U11419 ( .A1(n12187), .A2(n12186), .ZN(n18161) );
  AND2_X2 U11420 ( .A1(n10278), .A2(n10973), .ZN(n10300) );
  NAND2_X1 U11421 ( .A1(n10980), .A2(n19503), .ZN(n10502) );
  INV_X1 U11422 ( .A(n19503), .ZN(n20179) );
  NAND2_X2 U11423 ( .A1(n11250), .A2(n11249), .ZN(n11352) );
  NAND2_X2 U11424 ( .A1(n10039), .A2(n10037), .ZN(n19503) );
  NAND2_X1 U11425 ( .A1(n10198), .A2(n10199), .ZN(n10278) );
  AND4_X1 U11426 ( .A1(n11248), .A2(n11247), .A3(n11246), .A4(n11245), .ZN(
        n11249) );
  AND2_X1 U11427 ( .A1(n11240), .A2(n11239), .ZN(n11371) );
  AND4_X1 U11428 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11326) );
  AND4_X1 U11429 ( .A1(n11314), .A2(n11313), .A3(n11312), .A4(n11311), .ZN(
        n11325) );
  AND4_X1 U11430 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .ZN(
        n11250) );
  AND4_X1 U11431 ( .A1(n11322), .A2(n11321), .A3(n11320), .A4(n11319), .ZN(
        n11323) );
  AND4_X1 U11432 ( .A1(n11228), .A2(n11227), .A3(n11226), .A4(n11225), .ZN(
        n11240) );
  AND4_X1 U11433 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11347) );
  AND4_X1 U11434 ( .A1(n11269), .A2(n11268), .A3(n11267), .A4(n11266), .ZN(
        n11280) );
  AND4_X1 U11435 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n11346) );
  NOR2_X1 U11436 ( .A1(n13531), .A2(n16520), .ZN(n13534) );
  NAND2_X1 U11437 ( .A1(n10040), .A2(n16039), .ZN(n10039) );
  NAND2_X1 U11438 ( .A1(n10038), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10037) );
  AND2_X1 U11439 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  AND4_X1 U11440 ( .A1(n11343), .A2(n11342), .A3(n11341), .A4(n11340), .ZN(
        n11344) );
  INV_X2 U11441 ( .A(n17714), .ZN(n17722) );
  AND4_X1 U11442 ( .A1(n11273), .A2(n11272), .A3(n11271), .A4(n11270), .ZN(
        n11279) );
  NAND2_X2 U11443 ( .A1(n19069), .A2(n19014), .ZN(n19072) );
  INV_X2 U11444 ( .A(n16804), .ZN(U215) );
  INV_X2 U11445 ( .A(n19428), .ZN(n19454) );
  BUF_X2 U11446 ( .A(n12188), .Z(n17462) );
  INV_X1 U11447 ( .A(n12168), .ZN(n12253) );
  INV_X2 U11448 ( .A(n10151), .ZN(n17471) );
  BUF_X2 U11449 ( .A(n12318), .Z(n17481) );
  INV_X1 U11450 ( .A(n12901), .ZN(n12470) );
  INV_X1 U11451 ( .A(n12901), .ZN(n9743) );
  AND3_X1 U11452 ( .A1(n10174), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10173), .ZN(n10178) );
  BUF_X2 U11453 ( .A(n12191), .Z(n9729) );
  NOR2_X2 U11454 ( .A1(n12146), .A2(n12142), .ZN(n12316) );
  NOR2_X4 U11455 ( .A1(n12145), .A2(n12144), .ZN(n17461) );
  INV_X1 U11456 ( .A(n9934), .ZN(n9745) );
  NOR2_X1 U11457 ( .A1(n12143), .A2(n18921), .ZN(n12168) );
  INV_X2 U11458 ( .A(n16808), .ZN(n16810) );
  NAND2_X2 U11459 ( .A1(n10783), .A2(n9935), .ZN(n9934) );
  NAND2_X1 U11460 ( .A1(n19085), .A2(n19096), .ZN(n12145) );
  AND2_X2 U11461 ( .A1(n16020), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14524) );
  NAND2_X1 U11462 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19103), .ZN(
        n12146) );
  AND2_X2 U11463 ( .A1(n16020), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9736) );
  NAND2_X1 U11464 ( .A1(n19085), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12143) );
  AND2_X1 U11465 ( .A1(n11223), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11233) );
  INV_X2 U11466 ( .A(n18455), .ZN(n9731) );
  AND2_X1 U11467 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11232) );
  NOR2_X2 U11468 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13231) );
  NOR2_X2 U11469 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16020) );
  AND2_X1 U11470 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16017) );
  NAND2_X1 U11471 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18948) );
  CLKBUF_X1 U11472 ( .A(n10629), .Z(n9732) );
  NAND2_X1 U11473 ( .A1(n10939), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9733) );
  INV_X2 U11474 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11229) );
  NAND2_X1 U11475 ( .A1(n20352), .A2(n20351), .ZN(n20354) );
  AND3_X1 U11476 ( .A1(n10280), .A2(n10300), .A3(n10279), .ZN(n10794) );
  NOR2_X4 U11477 ( .A1(n14755), .A2(n14756), .ZN(n14740) );
  NAND2_X2 U11478 ( .A1(n14773), .A2(n14775), .ZN(n14755) );
  OR2_X1 U11479 ( .A1(n12144), .A2(n12143), .ZN(n10151) );
  OR2_X1 U11480 ( .A1(n9741), .A2(n10522), .ZN(n10342) );
  OR2_X2 U11481 ( .A1(n9733), .A2(n10329), .ZN(n9804) );
  NOR2_X2 U11482 ( .A1(n15525), .A2(n15526), .ZN(n14516) );
  NAND2_X2 U11483 ( .A1(n14705), .A2(n14308), .ZN(n13168) );
  NAND2_X1 U11484 ( .A1(n10353), .A2(n10354), .ZN(n10362) );
  NAND2_X1 U11485 ( .A1(n9918), .A2(n9796), .ZN(n10036) );
  AOI221_X1 U11486 ( .B1(n17512), .B2(n17523), .C1(n17647), .C2(n17523), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17514) );
  NOR4_X4 U11487 ( .A1(n19132), .A2(n18485), .A3(n16212), .A4(n18983), .ZN(
        n17523) );
  NAND2_X2 U11488 ( .A1(n9879), .A2(n9918), .ZN(n10815) );
  AND2_X2 U11489 ( .A1(n10463), .A2(n10825), .ZN(n9879) );
  NAND2_X2 U11490 ( .A1(n13008), .A2(n10212), .ZN(n10276) );
  AND2_X1 U11491 ( .A1(n16020), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9735) );
  OAI21_X2 U11492 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n14437), .A(n14429), 
        .ZN(n15347) );
  INV_X2 U11493 ( .A(n13890), .ZN(n10268) );
  NAND2_X2 U11494 ( .A1(n9804), .A2(n10332), .ZN(n10335) );
  NOR2_X2 U11495 ( .A1(n15679), .A2(n15678), .ZN(n15873) );
  AND2_X2 U11496 ( .A1(n14858), .A2(n14859), .ZN(n14824) );
  NOR2_X2 U11497 ( .A1(n14271), .A2(n14931), .ZN(n14858) );
  OAI21_X1 U11498 ( .B1(n11441), .B2(n11229), .A(n11482), .ZN(n13283) );
  NAND2_X2 U11499 ( .A1(n10304), .A2(n10303), .ZN(n10939) );
  INV_X2 U11500 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10077) );
  AND2_X4 U11501 ( .A1(n10783), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10188) );
  AND2_X2 U11502 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10783) );
  INV_X2 U11503 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10487) );
  OR2_X2 U11504 ( .A1(n13284), .A2(n11380), .ZN(n20420) );
  INV_X2 U11505 ( .A(n9934), .ZN(n9746) );
  NAND2_X1 U11506 ( .A1(n10939), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U11507 ( .A1(n10939), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9742) );
  INV_X2 U11508 ( .A(n9749), .ZN(n10013) );
  INV_X2 U11510 ( .A(n9934), .ZN(n14534) );
  AND3_X4 U11511 ( .A1(n10487), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10240) );
  XNOR2_X1 U11512 ( .A(n11479), .B(n11477), .ZN(n11765) );
  XNOR2_X2 U11513 ( .A(n11410), .B(n11409), .ZN(n11787) );
  BUF_X2 U11514 ( .A(n10374), .Z(n13064) );
  BUF_X1 U11515 ( .A(n10369), .Z(n9749) );
  XNOR2_X1 U11516 ( .A(n10351), .B(n10350), .ZN(n10369) );
  OR2_X1 U11517 ( .A1(n10374), .A2(n10360), .ZN(n10555) );
  OR2_X1 U11518 ( .A1(n10370), .A2(n10374), .ZN(n10543) );
  OR2_X1 U11519 ( .A1(n10374), .A2(n10366), .ZN(n19764) );
  NOR2_X2 U11520 ( .A1(n11355), .A2(n11327), .ZN(n12720) );
  NAND4_X2 U11521 ( .A1(n9865), .A2(n9864), .A3(n9866), .A4(n9863), .ZN(n11355) );
  INV_X1 U11522 ( .A(n9742), .ZN(n9751) );
  NAND2_X1 U11523 ( .A1(n12791), .A2(n11292), .ZN(n9866) );
  OR2_X1 U11524 ( .A1(n14308), .A2(n13438), .ZN(n14238) );
  NOR2_X1 U11525 ( .A1(n10980), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10979) );
  INV_X1 U11526 ( .A(n11358), .ZN(n11674) );
  NOR2_X1 U11527 ( .A1(n9961), .A2(n9962), .ZN(n9960) );
  INV_X1 U11528 ( .A(n11547), .ZN(n9962) );
  NAND2_X1 U11529 ( .A1(n14989), .A2(n15171), .ZN(n14381) );
  OAI21_X1 U11530 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n15009) );
  NAND2_X1 U11531 ( .A1(n9808), .A2(n11601), .ZN(n10130) );
  INV_X1 U11532 ( .A(n15054), .ZN(n10132) );
  NAND2_X1 U11533 ( .A1(n14375), .A2(n9808), .ZN(n10131) );
  NAND2_X1 U11534 ( .A1(n11292), .A2(n11428), .ZN(n9865) );
  NAND2_X1 U11535 ( .A1(n11359), .A2(n11428), .ZN(n9863) );
  OAI21_X1 U11536 ( .B1(n13034), .B2(n9862), .A(n9860), .ZN(n9864) );
  NAND2_X1 U11537 ( .A1(n14601), .A2(n10076), .ZN(n10073) );
  AND2_X1 U11538 ( .A1(n10031), .A2(n13864), .ZN(n10030) );
  AND2_X1 U11539 ( .A1(n9806), .A2(n9752), .ZN(n9903) );
  INV_X1 U11540 ( .A(n10845), .ZN(n10057) );
  AOI21_X1 U11541 ( .B1(n10845), .B2(n15989), .A(n15984), .ZN(n10056) );
  INV_X1 U11542 ( .A(n14444), .ZN(n11211) );
  AND4_X1 U11543 ( .A1(n11318), .A2(n11317), .A3(n11316), .A4(n11315), .ZN(
        n11324) );
  OR2_X1 U11544 ( .A1(n12484), .A2(n20939), .ZN(n13487) );
  OR3_X1 U11545 ( .A1(n9955), .A2(n13808), .A3(n13966), .ZN(n9954) );
  NAND2_X1 U11546 ( .A1(n10710), .A2(n9822), .ZN(n10717) );
  AND2_X1 U11547 ( .A1(n10813), .A2(n16682), .ZN(n11173) );
  NAND2_X1 U11548 ( .A1(n12828), .A2(n12827), .ZN(n12943) );
  OR2_X1 U11549 ( .A1(n19549), .A2(n20161), .ZN(n19877) );
  AND2_X1 U11550 ( .A1(n9980), .A2(n17171), .ZN(n16848) );
  OR2_X1 U11551 ( .A1(n16858), .A2(n16859), .ZN(n9980) );
  NOR2_X1 U11552 ( .A1(n9990), .A2(n9993), .ZN(n9989) );
  INV_X1 U11553 ( .A(n9991), .ZN(n9990) );
  OAI21_X1 U11554 ( .B1(n12445), .B2(n9897), .A(n9896), .ZN(n17793) );
  NAND2_X1 U11555 ( .A1(n9898), .A2(n18075), .ZN(n9897) );
  NAND2_X1 U11556 ( .A1(n12549), .A2(n9898), .ZN(n9896) );
  INV_X1 U11557 ( .A(n17794), .ZN(n9898) );
  NAND2_X1 U11558 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17907), .ZN(
        n17882) );
  XNOR2_X1 U11559 ( .A(n15369), .B(n11217), .ZN(n16423) );
  AND4_X1 U11560 ( .A1(n10481), .A2(n10480), .A3(n10479), .A4(n10478), .ZN(
        n10482) );
  NOR2_X1 U11561 ( .A1(n15096), .A2(n10136), .ZN(n10134) );
  OR2_X1 U11562 ( .A1(n10139), .A2(n10140), .ZN(n10136) );
  INV_X1 U11563 ( .A(n11595), .ZN(n10140) );
  INV_X1 U11564 ( .A(n11605), .ZN(n10139) );
  AND2_X1 U11565 ( .A1(n11560), .A2(n11559), .ZN(n11563) );
  AND2_X1 U11566 ( .A1(n11410), .A2(n11408), .ZN(n11380) );
  INV_X1 U11567 ( .A(n11369), .ZN(n10113) );
  NOR2_X1 U11568 ( .A1(n11223), .A2(n10118), .ZN(n10117) );
  OAI21_X1 U11569 ( .B1(n11355), .B2(n13135), .A(n13282), .ZN(n11364) );
  OAI21_X1 U11570 ( .B1(n12515), .B2(n12769), .A(n13044), .ZN(n11354) );
  NAND2_X1 U11571 ( .A1(n11367), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11435) );
  NAND2_X1 U11572 ( .A1(n10492), .A2(n10491), .ZN(n10494) );
  NAND2_X1 U11573 ( .A1(n10505), .A2(n10503), .ZN(n10492) );
  XNOR2_X1 U11574 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10493) );
  AND2_X1 U11575 ( .A1(n10494), .A2(n10493), .ZN(n10524) );
  CLKBUF_X1 U11576 ( .A(n14524), .Z(n14681) );
  NAND4_X1 U11577 ( .A1(n10278), .A2(n13430), .A3(n13008), .A4(n10267), .ZN(
        n10285) );
  NAND2_X1 U11578 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10015) );
  NAND2_X1 U11579 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10016) );
  INV_X1 U11580 ( .A(n10431), .ZN(n10434) );
  NAND2_X1 U11581 ( .A1(n10796), .A2(n10267), .ZN(n10804) );
  NAND2_X1 U11582 ( .A1(n10013), .A2(n10364), .ZN(n10371) );
  NAND2_X1 U11583 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12142) );
  AND2_X1 U11584 ( .A1(n12373), .A2(n12372), .ZN(n12377) );
  INV_X1 U11585 ( .A(n14783), .ZN(n9969) );
  AND2_X1 U11586 ( .A1(n9811), .A2(n14798), .ZN(n9970) );
  AND2_X1 U11587 ( .A1(n12072), .A2(n14921), .ZN(n12073) );
  NAND2_X1 U11588 ( .A1(n14359), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12509) );
  NOR2_X1 U11589 ( .A1(n11291), .A2(n20616), .ZN(n11766) );
  NAND2_X1 U11590 ( .A1(n13872), .A2(n9768), .ZN(n14253) );
  INV_X1 U11591 ( .A(n11955), .ZN(n11943) );
  NOR2_X1 U11592 ( .A1(n11360), .A2(n20616), .ZN(n11955) );
  NAND2_X1 U11593 ( .A1(n9871), .A2(n9869), .ZN(n15139) );
  INV_X1 U11594 ( .A(n11594), .ZN(n9870) );
  INV_X1 U11595 ( .A(n14059), .ZN(n9955) );
  AOI21_X1 U11596 ( .B1(n11431), .B2(n11622), .A(n13732), .ZN(n10127) );
  NAND2_X1 U11597 ( .A1(n13284), .A2(n11380), .ZN(n11440) );
  INV_X1 U11598 ( .A(n11477), .ZN(n11478) );
  NAND2_X1 U11599 ( .A1(n12610), .A2(n10118), .ZN(n11494) );
  INV_X1 U11600 ( .A(n19503), .ZN(n10071) );
  AOI21_X1 U11601 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20142), .A(
        n10524), .ZN(n10744) );
  INV_X1 U11602 ( .A(n9937), .ZN(n10681) );
  NOR2_X1 U11603 ( .A1(n10693), .A2(n10684), .ZN(n10687) );
  NOR4_X2 U11604 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13846) );
  OR2_X1 U11605 ( .A1(n14575), .A2(n14576), .ZN(n14577) );
  AND2_X1 U11606 ( .A1(n10028), .A2(n10027), .ZN(n10026) );
  INV_X1 U11607 ( .A(n15401), .ZN(n10027) );
  AND2_X1 U11608 ( .A1(n15416), .A2(n15569), .ZN(n10028) );
  INV_X1 U11609 ( .A(n14071), .ZN(n10090) );
  AND2_X1 U11610 ( .A1(n10707), .A2(n9913), .ZN(n9912) );
  NAND2_X1 U11611 ( .A1(n15427), .A2(n10102), .ZN(n10101) );
  NOR2_X1 U11612 ( .A1(n15440), .A2(n15413), .ZN(n10102) );
  NAND2_X1 U11613 ( .A1(n15709), .A2(n9854), .ZN(n15667) );
  AND2_X1 U11614 ( .A1(n11144), .A2(n15956), .ZN(n10031) );
  NOR2_X1 U11615 ( .A1(n10092), .A2(n13878), .ZN(n10091) );
  INV_X1 U11616 ( .A(n13819), .ZN(n10092) );
  NOR2_X1 U11617 ( .A1(n15967), .A2(n10146), .ZN(n10145) );
  INV_X1 U11618 ( .A(n10638), .ZN(n10146) );
  NAND2_X1 U11620 ( .A1(n10338), .A2(n10337), .ZN(n9925) );
  OR2_X1 U11621 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  INV_X1 U11622 ( .A(n13014), .ZN(n10099) );
  INV_X1 U11623 ( .A(n10816), .ZN(n9930) );
  OR2_X1 U11624 ( .A1(n9750), .A2(n12831), .ZN(n10383) );
  OR2_X1 U11625 ( .A1(n10374), .A2(n19481), .ZN(n10386) );
  NAND2_X1 U11626 ( .A1(n10055), .A2(n16039), .ZN(n10054) );
  NAND2_X1 U11627 ( .A1(n10053), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10052) );
  NAND2_X1 U11628 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19109), .ZN(
        n12144) );
  NOR2_X1 U11629 ( .A1(n17188), .A2(n12140), .ZN(n12315) );
  NAND2_X1 U11630 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17862), .ZN(
        n17837) );
  OR2_X1 U11631 ( .A1(n18064), .A2(n12431), .ZN(n17973) );
  INV_X1 U11632 ( .A(n10062), .ZN(n12242) );
  NAND2_X1 U11633 ( .A1(n18090), .A2(n12385), .ZN(n12389) );
  NOR2_X1 U11634 ( .A1(n12238), .A2(n18115), .ZN(n12240) );
  INV_X1 U11635 ( .A(n10065), .ZN(n12236) );
  NOR2_X1 U11636 ( .A1(n9891), .A2(n12237), .ZN(n12239) );
  OR2_X1 U11637 ( .A1(n16216), .A2(n12344), .ZN(n12414) );
  OR2_X1 U11638 ( .A1(n12406), .A2(n12413), .ZN(n12418) );
  OR2_X1 U11639 ( .A1(n12337), .A2(n18919), .ZN(n16053) );
  NAND2_X1 U11640 ( .A1(n17678), .A2(n17728), .ZN(n12357) );
  AND2_X1 U11641 ( .A1(n20696), .A2(n13478), .ZN(n14892) );
  AND2_X1 U11642 ( .A1(n12924), .A2(n13032), .ZN(n13133) );
  AND2_X1 U11643 ( .A1(n20616), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12512) );
  INV_X1 U11644 ( .A(n14710), .ZN(n9965) );
  AND2_X1 U11645 ( .A1(n13487), .A2(n12485), .ZN(n15003) );
  OR2_X1 U11646 ( .A1(n12115), .A2(n14763), .ZN(n12127) );
  NAND2_X1 U11647 ( .A1(n11680), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12074) );
  OR2_X1 U11648 ( .A1(n11848), .A2(n20970), .ZN(n11853) );
  NAND2_X1 U11649 ( .A1(n13403), .A2(n11503), .ZN(n20352) );
  NAND2_X1 U11650 ( .A1(n10133), .A2(n15186), .ZN(n14376) );
  NOR2_X1 U11651 ( .A1(n14374), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9873) );
  INV_X1 U11652 ( .A(n11613), .ZN(n9874) );
  NAND2_X1 U11653 ( .A1(n16384), .A2(n9953), .ZN(n9952) );
  NOR2_X1 U11654 ( .A1(n13617), .A2(n13344), .ZN(n9953) );
  OR2_X1 U11655 ( .A1(n13345), .A2(n9950), .ZN(n16386) );
  NAND2_X1 U11656 ( .A1(n16384), .A2(n9951), .ZN(n9950) );
  INV_X1 U11657 ( .A(n13344), .ZN(n9951) );
  NAND2_X1 U11658 ( .A1(n13039), .A2(n13038), .ZN(n13054) );
  OR2_X1 U11659 ( .A1(n13037), .A2(n13036), .ZN(n13038) );
  NAND2_X1 U11660 ( .A1(n20420), .A2(n11440), .ZN(n12612) );
  OR2_X1 U11661 ( .A1(n9862), .A2(n13472), .ZN(n11327) );
  AND2_X1 U11662 ( .A1(n12611), .A2(n13370), .ZN(n20493) );
  INV_X1 U11663 ( .A(n13740), .ZN(n20448) );
  NOR2_X1 U11664 ( .A1(n13746), .A2(n14154), .ZN(n20454) );
  NOR2_X1 U11665 ( .A1(n11195), .A2(n11194), .ZN(n11198) );
  AND2_X1 U11666 ( .A1(n10709), .A2(n10708), .ZN(n10710) );
  NAND2_X1 U11667 ( .A1(n10711), .A2(n10725), .ZN(n10709) );
  INV_X1 U11668 ( .A(n13122), .ZN(n10085) );
  AND2_X1 U11669 ( .A1(n14675), .A2(n10082), .ZN(n10080) );
  AND2_X1 U11670 ( .A1(n11023), .A2(n11022), .ZN(n15993) );
  OR2_X1 U11671 ( .A1(n11008), .A2(n11007), .ZN(n13417) );
  NOR2_X1 U11672 ( .A1(n9999), .A2(n9996), .ZN(n9994) );
  INV_X1 U11673 ( .A(n10839), .ZN(n16532) );
  XNOR2_X1 U11674 ( .A(n9936), .B(n10929), .ZN(n15618) );
  NAND2_X1 U11675 ( .A1(n10729), .A2(n10626), .ZN(n9936) );
  OR2_X1 U11676 ( .A1(n15423), .A2(n11020), .ZN(n10714) );
  NAND2_X1 U11677 ( .A1(n9772), .A2(n10143), .ZN(n10142) );
  NAND2_X1 U11678 ( .A1(n10650), .A2(n9771), .ZN(n10141) );
  NOR2_X1 U11679 ( .A1(n15645), .A2(n15753), .ZN(n15648) );
  INV_X1 U11680 ( .A(n15993), .ZN(n11024) );
  NAND2_X1 U11681 ( .A1(n9761), .A2(n13992), .ZN(n9926) );
  NAND2_X1 U11682 ( .A1(n9876), .A2(n13447), .ZN(n9901) );
  AND2_X1 U11683 ( .A1(n10098), .A2(n10100), .ZN(n13019) );
  NAND2_X1 U11684 ( .A1(n10523), .A2(n10522), .ZN(n13446) );
  AOI21_X1 U11685 ( .B1(n12831), .B2(n12994), .A(n12830), .ZN(n12832) );
  NAND2_X1 U11686 ( .A1(n20145), .A2(n20153), .ZN(n19820) );
  NAND2_X1 U11687 ( .A1(n15465), .A2(n20153), .ZN(n19672) );
  OR2_X1 U11688 ( .A1(n19549), .A2(n19548), .ZN(n19851) );
  NAND2_X1 U11689 ( .A1(n15465), .A2(n19573), .ZN(n19758) );
  INV_X1 U11690 ( .A(n19758), .ZN(n19994) );
  NAND2_X1 U11691 ( .A1(n16044), .A2(n12862), .ZN(n12863) );
  INV_X1 U11692 ( .A(n19999), .ZN(n19913) );
  INV_X1 U11693 ( .A(n16816), .ZN(n18959) );
  INV_X1 U11694 ( .A(n17853), .ZN(n9977) );
  NOR2_X1 U11695 ( .A1(n16910), .A2(n9816), .ZN(n9974) );
  INV_X1 U11696 ( .A(n9989), .ZN(n9987) );
  INV_X1 U11697 ( .A(n16215), .ZN(n17524) );
  NAND2_X1 U11698 ( .A1(n12341), .A2(n12422), .ZN(n17728) );
  AND2_X1 U11699 ( .A1(n17987), .A2(n9766), .ZN(n17907) );
  NOR2_X1 U11700 ( .A1(n18074), .A2(n20850), .ZN(n18073) );
  NAND2_X1 U11701 ( .A1(n12444), .A2(n16151), .ZN(n12445) );
  AND2_X1 U11702 ( .A1(n17913), .A2(n9894), .ZN(n17849) );
  AND2_X1 U11703 ( .A1(n12440), .A2(n9895), .ZN(n9894) );
  AND2_X1 U11704 ( .A1(n12435), .A2(n10156), .ZN(n12436) );
  OR2_X1 U11705 ( .A1(n17956), .A2(n18280), .ZN(n12435) );
  XNOR2_X1 U11706 ( .A(n12240), .B(n10064), .ZN(n18104) );
  OR2_X1 U11707 ( .A1(n18104), .A2(n18105), .ZN(n10063) );
  OR2_X1 U11708 ( .A1(n18134), .A2(n18133), .ZN(n10066) );
  NOR2_X1 U11709 ( .A1(n13479), .A2(n13472), .ZN(n13495) );
  AND2_X1 U11710 ( .A1(n13149), .A2(n12802), .ZN(n20696) );
  CLKBUF_X1 U11711 ( .A(n12612), .Z(n12613) );
  NAND3_X1 U11712 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20152), .A3(n19999), 
        .ZN(n13256) );
  XNOR2_X1 U11713 ( .A(n15346), .B(n14428), .ZN(n16422) );
  AOI21_X1 U11714 ( .B1(n16423), .B2(n16621), .A(n10154), .ZN(n11219) );
  NOR2_X1 U11715 ( .A1(n15611), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15809) );
  OAI21_X1 U11716 ( .B1(n15807), .B2(n19491), .A(n10048), .ZN(n10047) );
  AOI21_X1 U11717 ( .B1(n15811), .B2(n15810), .A(n10049), .ZN(n10048) );
  NAND2_X1 U11718 ( .A1(n9924), .A2(n10929), .ZN(n9923) );
  INV_X1 U11719 ( .A(n16639), .ZN(n19500) );
  OR2_X1 U11720 ( .A1(n12943), .A2(n12839), .ZN(n20161) );
  INV_X1 U11721 ( .A(n20050), .ZN(n19538) );
  OAI21_X1 U11722 ( .B1(n16848), .B2(n9842), .A(n9762), .ZN(n9978) );
  AND2_X1 U11723 ( .A1(n16853), .A2(n17208), .ZN(n9979) );
  INV_X1 U11724 ( .A(n17182), .ZN(n17181) );
  NOR2_X2 U11725 ( .A1(n19079), .A2(n17185), .ZN(n17182) );
  NOR2_X1 U11726 ( .A1(n12218), .A2(n12217), .ZN(n17655) );
  AOI21_X1 U11727 ( .B1(n12574), .B2(n18034), .A(n12568), .ZN(n12569) );
  INV_X1 U11728 ( .A(n12567), .ZN(n12568) );
  NAND2_X1 U11729 ( .A1(n17830), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17814) );
  INV_X1 U11730 ( .A(n18079), .ZN(n18034) );
  NAND2_X1 U11731 ( .A1(n12557), .A2(n18131), .ZN(n18042) );
  INV_X1 U11732 ( .A(n18042), .ZN(n18076) );
  OR2_X1 U11733 ( .A1(n16819), .A2(n17729), .ZN(n18167) );
  AOI21_X1 U11734 ( .B1(n18439), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10162), .ZN(n12446) );
  AOI21_X1 U11735 ( .B1(n17803), .B2(n18961), .A(n10067), .ZN(n18168) );
  INV_X1 U11736 ( .A(n10068), .ZN(n10067) );
  AOI21_X1 U11737 ( .B1(n17804), .B2(n18339), .A(n10069), .ZN(n10068) );
  NAND2_X1 U11738 ( .A1(n18176), .A2(n10070), .ZN(n10069) );
  INV_X1 U11739 ( .A(n18454), .ZN(n18439) );
  NOR2_X1 U11740 ( .A1(n18193), .A2(n18461), .ZN(n18460) );
  NOR2_X1 U11741 ( .A1(n18956), .A2(n18461), .ZN(n18458) );
  NAND2_X1 U11742 ( .A1(n11372), .A2(n11291), .ZN(n11675) );
  AND2_X1 U11743 ( .A1(n13886), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10412) );
  NAND2_X1 U11744 ( .A1(n10411), .A2(n10410), .ZN(n10413) );
  NAND2_X1 U11745 ( .A1(n10323), .A2(n10322), .ZN(n10325) );
  AOI22_X1 U11746 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U11747 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10245) );
  AOI21_X1 U11748 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18934), .A(
        n12399), .ZN(n12401) );
  AND2_X1 U11749 ( .A1(n11617), .A2(n11616), .ZN(n11648) );
  NOR2_X1 U11750 ( .A1(n11624), .A2(n11625), .ZN(n11623) );
  OR2_X1 U11751 ( .A1(n11420), .A2(n11419), .ZN(n11581) );
  OR2_X1 U11752 ( .A1(n11535), .A2(n11534), .ZN(n11566) );
  NAND2_X1 U11753 ( .A1(n9861), .A2(n13034), .ZN(n9860) );
  NAND2_X1 U11754 ( .A1(n11360), .A2(n11352), .ZN(n9861) );
  AOI22_X1 U11755 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11303) );
  OR2_X1 U11756 ( .A1(n11492), .A2(n11491), .ZN(n11539) );
  OR2_X1 U11757 ( .A1(n11348), .A2(n10118), .ZN(n11450) );
  AOI21_X1 U11758 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16172), .A(
        n11623), .ZN(n11660) );
  NAND3_X1 U11759 ( .A1(n13472), .A2(n11348), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11662) );
  NAND2_X1 U11760 ( .A1(n20159), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10489) );
  AOI21_X1 U11761 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(n9850), .ZN(n14655) );
  AOI21_X1 U11762 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n9851), .ZN(n14668) );
  AOI21_X1 U11763 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A(n9840), .ZN(n14610) );
  AOI21_X1 U11764 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A(n9838), .ZN(n14585) );
  AOI21_X1 U11765 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n9839), .ZN(n14594) );
  AOI21_X1 U11766 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n9836), .ZN(n14566) );
  AOI21_X1 U11767 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A(n9837), .ZN(n14557) );
  AOI21_X1 U11768 ( .B1(n14524), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A(
        n9825), .ZN(n14499) );
  AOI21_X1 U11769 ( .B1(n9736), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A(n9826), 
        .ZN(n14491) );
  OR2_X1 U11770 ( .A1(n10402), .A2(n10401), .ZN(n10498) );
  NOR2_X1 U11771 ( .A1(n10036), .A2(n10589), .ZN(n10621) );
  AND4_X1 U11772 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10484) );
  AND4_X1 U11773 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n10485) );
  AND4_X1 U11774 ( .A1(n10476), .A2(n10475), .A3(n10474), .A4(n10473), .ZN(
        n10483) );
  OR2_X1 U11775 ( .A1(n10450), .A2(n10449), .ZN(n10818) );
  AND2_X1 U11776 ( .A1(n10800), .A2(n10973), .ZN(n10225) );
  AOI22_X1 U11777 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U11778 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U11779 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U11780 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U11781 ( .A1(n10374), .A2(n10365), .ZN(n10557) );
  NAND2_X1 U11782 ( .A1(n10748), .A2(n10489), .ZN(n10505) );
  AND2_X1 U11783 ( .A1(n10491), .A2(n10490), .ZN(n10503) );
  OR2_X1 U11784 ( .A1(n10754), .A2(n10747), .ZN(n10748) );
  NOR2_X1 U11785 ( .A1(n17655), .A2(n12383), .ZN(n12387) );
  AND2_X1 U11786 ( .A1(n9967), .A2(n14720), .ZN(n9966) );
  AND2_X1 U11787 ( .A1(n9968), .A2(n14742), .ZN(n9967) );
  INV_X1 U11788 ( .A(n12131), .ZN(n9968) );
  INV_X1 U11789 ( .A(n14809), .ZN(n9971) );
  AND2_X1 U11790 ( .A1(n9964), .A2(n9831), .ZN(n9963) );
  OR2_X1 U11791 ( .A1(n9768), .A2(n9812), .ZN(n9964) );
  AND3_X1 U11792 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(n11816), .ZN(n11815) );
  NAND2_X1 U11793 ( .A1(n11525), .A2(n11524), .ZN(n9877) );
  NOR2_X1 U11794 ( .A1(n9959), .A2(n14760), .ZN(n9958) );
  INV_X1 U11795 ( .A(n14771), .ZN(n9959) );
  NAND2_X1 U11796 ( .A1(n9946), .A2(n9944), .ZN(n14827) );
  NOR2_X1 U11797 ( .A1(n9767), .A2(n9945), .ZN(n9944) );
  INV_X1 U11798 ( .A(n14912), .ZN(n9945) );
  AND2_X1 U11799 ( .A1(n15278), .A2(n10138), .ZN(n10137) );
  NAND2_X1 U11800 ( .A1(n9764), .A2(n11605), .ZN(n10138) );
  OR2_X1 U11801 ( .A1(n11601), .A2(n11607), .ZN(n15118) );
  NAND2_X1 U11802 ( .A1(n20354), .A2(n10108), .ZN(n10107) );
  OR2_X1 U11803 ( .A1(n11558), .A2(n11557), .ZN(n11579) );
  INV_X1 U11804 ( .A(n11563), .ZN(n11561) );
  INV_X1 U11805 ( .A(n11564), .ZN(n11562) );
  AND2_X1 U11806 ( .A1(n11407), .A2(n10125), .ZN(n10124) );
  NAND2_X1 U11807 ( .A1(n10128), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10125) );
  OR2_X1 U11808 ( .A1(n11392), .A2(n11391), .ZN(n11464) );
  OR2_X1 U11809 ( .A1(n13472), .A2(n10118), .ZN(n11463) );
  NAND2_X1 U11810 ( .A1(n11381), .A2(n10118), .ZN(n11776) );
  XNOR2_X1 U11811 ( .A(n12952), .B(n13283), .ZN(n12610) );
  NAND2_X1 U11812 ( .A1(n11367), .A2(n10114), .ZN(n10111) );
  NOR2_X1 U11813 ( .A1(n11224), .A2(n10118), .ZN(n10114) );
  AND4_X1 U11814 ( .A1(n12785), .A2(n12784), .A3(n12783), .A4(n12883), .ZN(
        n13051) );
  AND2_X1 U11815 ( .A1(n11480), .A2(n13594), .ZN(n13826) );
  NAND2_X1 U11816 ( .A1(n10115), .A2(n10116), .ZN(n9859) );
  AOI21_X1 U11817 ( .B1(n11365), .B2(n10117), .A(n11366), .ZN(n10116) );
  NAND2_X1 U11818 ( .A1(n11367), .A2(n10117), .ZN(n10115) );
  NOR2_X1 U11819 ( .A1(n11662), .A2(n11622), .ZN(n11659) );
  NAND2_X1 U11820 ( .A1(n11450), .A2(n11463), .ZN(n11651) );
  INV_X1 U11821 ( .A(n13236), .ZN(n16163) );
  OR2_X1 U11822 ( .A1(n10524), .A2(n10495), .ZN(n10745) );
  AND3_X1 U11823 ( .A1(n12700), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10744), .ZN(n10746) );
  INV_X1 U11824 ( .A(n10623), .ZN(n9938) );
  NAND2_X1 U11825 ( .A1(n9937), .A2(n9829), .ZN(n10675) );
  NAND2_X1 U11826 ( .A1(n10687), .A2(n10659), .ZN(n10690) );
  AND2_X1 U11827 ( .A1(n11197), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10684) );
  NAND2_X1 U11828 ( .A1(n10642), .A2(n13107), .ZN(n10645) );
  NAND2_X1 U11829 ( .A1(n10725), .A2(n10640), .ZN(n10642) );
  NAND2_X1 U11830 ( .A1(n10639), .A2(n13103), .ZN(n10640) );
  AND3_X1 U11831 ( .A1(n9779), .A2(n10633), .A3(n10579), .ZN(n10639) );
  NAND2_X1 U11832 ( .A1(n10579), .A2(n9940), .ZN(n10624) );
  NAND2_X1 U11833 ( .A1(n11214), .A2(n10020), .ZN(n10019) );
  NOR2_X1 U11834 ( .A1(n10022), .A2(n11167), .ZN(n10020) );
  NAND2_X1 U11835 ( .A1(n14445), .A2(n14441), .ZN(n10022) );
  NAND2_X1 U11836 ( .A1(n9843), .A2(n10018), .ZN(n10017) );
  INV_X1 U11837 ( .A(n11167), .ZN(n10018) );
  AOI21_X1 U11838 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(n9853), .ZN(n14677) );
  AOI21_X1 U11839 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n9852), .ZN(n14683) );
  AOI21_X1 U11840 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A(n9848), .ZN(n14636) );
  AOI21_X1 U11841 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n9849), .ZN(n14645) );
  AOI21_X1 U11842 ( .B1(n14681), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n9841), .ZN(n14619) );
  NOR2_X1 U11843 ( .A1(n15508), .A2(n14547), .ZN(n14575) );
  AND2_X1 U11844 ( .A1(n9770), .A2(n10087), .ZN(n10086) );
  INV_X1 U11845 ( .A(n14088), .ZN(n10087) );
  NAND2_X1 U11846 ( .A1(n10299), .A2(n10298), .ZN(n10945) );
  NOR2_X1 U11847 ( .A1(n15386), .A2(n9998), .ZN(n9997) );
  INV_X1 U11848 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9998) );
  NOR2_X1 U11849 ( .A1(n15705), .A2(n10007), .ZN(n10006) );
  NOR2_X1 U11850 ( .A1(n16511), .A2(n10003), .ZN(n10002) );
  NOR2_X1 U11851 ( .A1(n16542), .A2(n10012), .ZN(n10011) );
  INV_X1 U11852 ( .A(n13504), .ZN(n10010) );
  NOR2_X1 U11853 ( .A1(n9906), .A2(n9908), .ZN(n9904) );
  OR2_X1 U11854 ( .A1(n15618), .A2(n15623), .ZN(n9906) );
  AND2_X1 U11855 ( .A1(n15901), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9919) );
  OR2_X1 U11856 ( .A1(n19214), .A2(n10677), .ZN(n15651) );
  OR2_X1 U11857 ( .A1(n13544), .A2(n11020), .ZN(n10651) );
  NOR2_X1 U11858 ( .A1(n10618), .A2(n10617), .ZN(n11017) );
  OR2_X1 U11859 ( .A1(n10462), .A2(n10461), .ZN(n10823) );
  NOR2_X1 U11860 ( .A1(n10434), .A2(n10014), .ZN(n10435) );
  NAND2_X1 U11861 ( .A1(n9789), .A2(n10268), .ZN(n10290) );
  INV_X1 U11862 ( .A(n10303), .ZN(n16019) );
  INV_X1 U11863 ( .A(n10383), .ZN(n10384) );
  AOI22_X1 U11864 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U11865 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U11866 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U11867 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U11868 ( .A1(n17188), .A2(n12145), .ZN(n12318) );
  OR2_X2 U11869 ( .A1(n12142), .A2(n17188), .ZN(n17267) );
  OR2_X1 U11870 ( .A1(n17188), .A2(n12143), .ZN(n10166) );
  OR2_X1 U11871 ( .A1(n12145), .A2(n18921), .ZN(n9776) );
  NOR2_X1 U11872 ( .A1(n19135), .A2(n16818), .ZN(n12632) );
  NOR2_X1 U11873 ( .A1(n18155), .A2(n9992), .ZN(n9991) );
  INV_X1 U11874 ( .A(n18107), .ZN(n17126) );
  INV_X1 U11875 ( .A(n12433), .ZN(n12429) );
  NAND2_X1 U11876 ( .A1(n18080), .A2(n12391), .ZN(n12433) );
  NAND2_X1 U11877 ( .A1(n12387), .A2(n12386), .ZN(n12451) );
  NAND2_X1 U11878 ( .A1(n10063), .A2(n9798), .ZN(n10062) );
  NAND2_X1 U11879 ( .A1(n18112), .A2(n12375), .ZN(n12380) );
  XNOR2_X1 U11880 ( .A(n12377), .B(n9891), .ZN(n12374) );
  NAND2_X1 U11881 ( .A1(n10066), .A2(n9795), .ZN(n10065) );
  AOI21_X1 U11882 ( .B1(n12360), .B2(n12359), .A(n12358), .ZN(n18918) );
  NOR2_X1 U11883 ( .A1(n17729), .A2(n18485), .ZN(n17726) );
  NOR2_X1 U11884 ( .A1(n17533), .A2(n12338), .ZN(n17725) );
  INV_X1 U11885 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20834) );
  AND2_X1 U11886 ( .A1(n14247), .A2(n14246), .ZN(n14249) );
  INV_X1 U11887 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20970) );
  NOR2_X1 U11888 ( .A1(n11348), .A2(n11352), .ZN(n13136) );
  NAND2_X1 U11889 ( .A1(n13182), .A2(n11796), .ZN(n13145) );
  AND2_X1 U11890 ( .A1(n11359), .A2(n11291), .ZN(n13077) );
  INV_X1 U11891 ( .A(n14279), .ZN(n13197) );
  INV_X1 U11892 ( .A(n12127), .ZN(n11684) );
  INV_X1 U11893 ( .A(n12112), .ZN(n11682) );
  OAI21_X1 U11894 ( .B1(n13475), .B2(n15022), .A(n12122), .ZN(n14756) );
  NAND2_X1 U11895 ( .A1(n11681), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12099) );
  INV_X1 U11896 ( .A(n12096), .ZN(n11681) );
  OR2_X1 U11897 ( .A1(n12099), .A2(n14787), .ZN(n12112) );
  AND2_X1 U11898 ( .A1(n12011), .A2(n12010), .ZN(n14826) );
  AND2_X1 U11899 ( .A1(n11679), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12026) );
  INV_X1 U11900 ( .A(n12068), .ZN(n11679) );
  NOR2_X1 U11901 ( .A1(n11991), .A2(n15102), .ZN(n12069) );
  NAND2_X1 U11902 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n12069), .ZN(
        n12068) );
  AND2_X1 U11903 ( .A1(n12071), .A2(n12070), .ZN(n14921) );
  NOR2_X1 U11904 ( .A1(n11946), .A2(n16250), .ZN(n11977) );
  NAND2_X1 U11905 ( .A1(n11977), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11991) );
  NAND2_X1 U11906 ( .A1(n11930), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11946) );
  AND2_X1 U11907 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n11910), .ZN(
        n11926) );
  AND2_X1 U11908 ( .A1(n11878), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11883) );
  NOR2_X1 U11909 ( .A1(n11853), .A2(n20969), .ZN(n11878) );
  AND3_X1 U11910 ( .A1(n11852), .A2(n11851), .A3(n11850), .ZN(n13788) );
  CLKBUF_X1 U11911 ( .A(n13786), .Z(n13787) );
  AND2_X1 U11912 ( .A1(n11815), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11831) );
  AOI21_X1 U11913 ( .B1(n11828), .B2(n11955), .A(n11827), .ZN(n13437) );
  CLKBUF_X1 U11914 ( .A(n13351), .Z(n13352) );
  NAND2_X1 U11915 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11798) );
  NOR2_X1 U11916 ( .A1(n20834), .A2(n11798), .ZN(n11816) );
  OR2_X1 U11917 ( .A1(n16187), .A2(n20197), .ZN(n13037) );
  NAND2_X1 U11918 ( .A1(n9858), .A2(n13456), .ZN(n13457) );
  NOR2_X1 U11919 ( .A1(n14743), .A2(n14730), .ZN(n14729) );
  AND2_X1 U11920 ( .A1(n15220), .A2(n14407), .ZN(n15157) );
  NAND2_X1 U11921 ( .A1(n14770), .A2(n9956), .ZN(n14743) );
  NOR2_X1 U11922 ( .A1(n9957), .A2(n14745), .ZN(n9956) );
  INV_X1 U11923 ( .A(n9958), .ZN(n9957) );
  NAND2_X1 U11924 ( .A1(n14770), .A2(n9958), .ZN(n14758) );
  NOR2_X1 U11925 ( .A1(n14810), .A2(n14794), .ZN(n14795) );
  INV_X1 U11926 ( .A(n10133), .ZN(n15046) );
  OR2_X1 U11927 ( .A1(n14828), .A2(n14812), .ZN(n14810) );
  OAI21_X1 U11928 ( .B1(n15063), .B2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15097), .ZN(n15054) );
  NAND2_X1 U11929 ( .A1(n9948), .A2(n9947), .ZN(n14828) );
  INV_X1 U11930 ( .A(n14830), .ZN(n9947) );
  INV_X1 U11931 ( .A(n14827), .ZN(n9948) );
  NAND2_X1 U11932 ( .A1(n11611), .A2(n10121), .ZN(n15063) );
  AND2_X1 U11933 ( .A1(n11610), .A2(n20987), .ZN(n10121) );
  INV_X1 U11934 ( .A(n11610), .ZN(n10119) );
  NOR2_X1 U11935 ( .A1(n14862), .A2(n9767), .ZN(n14913) );
  NAND2_X1 U11936 ( .A1(n9946), .A2(n9949), .ZN(n14926) );
  XNOR2_X1 U11937 ( .A(n11601), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15090) );
  NAND2_X1 U11938 ( .A1(n15121), .A2(n15118), .ZN(n16296) );
  NOR2_X2 U11939 ( .A1(n14275), .A2(n14274), .ZN(n14934) );
  AND2_X1 U11940 ( .A1(n14243), .A2(n14242), .ZN(n14258) );
  AND2_X1 U11941 ( .A1(n14237), .A2(n14236), .ZN(n15307) );
  CLKBUF_X1 U11942 ( .A(n15139), .Z(n15140) );
  AND2_X1 U11943 ( .A1(n13961), .A2(n13960), .ZN(n13966) );
  AND2_X1 U11944 ( .A1(n13964), .A2(n13963), .ZN(n14059) );
  AND3_X1 U11945 ( .A1(n13807), .A2(n14238), .A3(n13806), .ZN(n13808) );
  NAND2_X1 U11946 ( .A1(n16314), .A2(n16316), .ZN(n11587) );
  INV_X1 U11947 ( .A(n11522), .ZN(n10110) );
  AND2_X1 U11948 ( .A1(n13441), .A2(n13440), .ZN(n16384) );
  AND3_X1 U11949 ( .A1(n13343), .A2(n14238), .A3(n13342), .ZN(n13344) );
  XNOR2_X1 U11950 ( .A(n11433), .B(n11432), .ZN(n13278) );
  AND2_X1 U11951 ( .A1(n13054), .A2(n16159), .ZN(n15293) );
  OR2_X1 U11952 ( .A1(n13361), .A2(n9794), .ZN(n11495) );
  OAI22_X1 U11953 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15335), .B1(n13243), 
        .B2(n20702), .ZN(n13239) );
  NAND2_X1 U11954 ( .A1(n9868), .A2(n9867), .ZN(n15329) );
  AND2_X2 U11955 ( .A1(n12894), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12903) );
  INV_X1 U11956 ( .A(n11352), .ZN(n13297) );
  OR2_X1 U11957 ( .A1(n12607), .A2(n13246), .ZN(n14149) );
  NAND2_X1 U11958 ( .A1(n12607), .A2(n13246), .ZN(n13639) );
  INV_X1 U11959 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n16172) );
  AOI221_X1 U11960 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10744), 
        .C1(n12700), .C2(n10744), .A(n10743), .ZN(n10781) );
  NOR2_X1 U11961 ( .A1(n10746), .A2(n10745), .ZN(n10777) );
  NAND2_X1 U11962 ( .A1(n10733), .A2(n10734), .ZN(n11195) );
  AND2_X1 U11963 ( .A1(n10723), .A2(n14424), .ZN(n10729) );
  OR2_X1 U11964 ( .A1(n10717), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10724) );
  NOR2_X1 U11965 ( .A1(n10724), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10728) );
  NAND2_X1 U11966 ( .A1(n10666), .A2(n10665), .ZN(n10711) );
  NOR2_X1 U11967 ( .A1(n10675), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10666) );
  AND2_X1 U11968 ( .A1(n10670), .A2(n10672), .ZN(n19201) );
  AND2_X1 U11969 ( .A1(n11197), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U11970 ( .A1(n10654), .A2(n9941), .ZN(n10693) );
  NOR2_X1 U11971 ( .A1(n10691), .A2(n9942), .ZN(n9941) );
  NAND2_X1 U11972 ( .A1(n10654), .A2(n10655), .ZN(n9943) );
  NAND2_X1 U11973 ( .A1(n10725), .A2(n10656), .ZN(n10654) );
  NOR2_X1 U11974 ( .A1(n10645), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10647) );
  INV_X1 U11975 ( .A(n15556), .ZN(n10025) );
  INV_X1 U11976 ( .A(n14625), .ZN(n10072) );
  NAND2_X1 U11977 ( .A1(n10171), .A2(n10026), .ZN(n15557) );
  NOR2_X1 U11978 ( .A1(n15519), .A2(n14517), .ZN(n15510) );
  AND2_X1 U11979 ( .A1(n14516), .A2(n14546), .ZN(n14517) );
  NOR2_X1 U11980 ( .A1(n15510), .A2(n15509), .ZN(n15508) );
  NAND2_X1 U11981 ( .A1(n13554), .A2(n9814), .ZN(n13982) );
  INV_X1 U11982 ( .A(n13910), .ZN(n10029) );
  NAND2_X1 U11983 ( .A1(n13907), .A2(n9770), .ZN(n14087) );
  AND2_X1 U11984 ( .A1(n19387), .A2(n13431), .ZN(n13717) );
  NAND2_X1 U11985 ( .A1(n15343), .A2(n14428), .ZN(n10093) );
  NAND2_X1 U11986 ( .A1(n10097), .A2(n10096), .ZN(n10095) );
  INV_X1 U11987 ( .A(n10937), .ZN(n10096) );
  INV_X1 U11988 ( .A(n15380), .ZN(n10097) );
  OR2_X1 U11989 ( .A1(n15379), .A2(n15380), .ZN(n15382) );
  NAND2_X1 U11990 ( .A1(n15363), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15365) );
  NAND2_X1 U11991 ( .A1(n15363), .A2(n9997), .ZN(n15349) );
  NAND2_X1 U11992 ( .A1(n15350), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15360) );
  NOR2_X1 U11993 ( .A1(n15358), .A2(n16487), .ZN(n15350) );
  NAND2_X1 U11994 ( .A1(n15359), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15358) );
  NOR2_X1 U11995 ( .A1(n15356), .A2(n15443), .ZN(n15359) );
  NAND2_X1 U11996 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n15357), .ZN(
        n15356) );
  AND2_X1 U11997 ( .A1(n14215), .A2(n10005), .ZN(n15357) );
  AND2_X1 U11998 ( .A1(n9769), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10005) );
  NAND2_X1 U11999 ( .A1(n14215), .A2(n9769), .ZN(n15353) );
  AND2_X1 U12000 ( .A1(n9763), .A2(n14199), .ZN(n10089) );
  NAND2_X1 U12001 ( .A1(n14215), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14214) );
  NOR2_X1 U12002 ( .A1(n14212), .A2(n19228), .ZN(n14215) );
  AND2_X1 U12003 ( .A1(n13534), .A2(n10001), .ZN(n14213) );
  AND2_X1 U12004 ( .A1(n9755), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10001) );
  NAND2_X1 U12005 ( .A1(n14213), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14212) );
  NAND2_X1 U12006 ( .A1(n13534), .A2(n9755), .ZN(n13549) );
  NAND2_X1 U12007 ( .A1(n13534), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13533) );
  AND2_X1 U12008 ( .A1(n10010), .A2(n9759), .ZN(n13532) );
  NAND2_X1 U12009 ( .A1(n10010), .A2(n10011), .ZN(n13529) );
  NOR2_X1 U12010 ( .A1(n13504), .A2(n16542), .ZN(n13530) );
  OR2_X1 U12011 ( .A1(n19320), .A2(n13797), .ZN(n9902) );
  INV_X1 U12012 ( .A(n13793), .ZN(n9900) );
  NOR2_X1 U12013 ( .A1(n13603), .A2(n13449), .ZN(n13505) );
  NAND2_X1 U12014 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13449) );
  NOR2_X1 U12015 ( .A1(n15379), .A2(n10095), .ZN(n15344) );
  INV_X1 U12016 ( .A(n15633), .ZN(n10058) );
  NOR2_X1 U12017 ( .A1(n15810), .A2(n10929), .ZN(n10059) );
  NOR2_X1 U12018 ( .A1(n11190), .A2(n11186), .ZN(n10738) );
  INV_X1 U12019 ( .A(n10050), .ZN(n10049) );
  AOI21_X1 U12020 ( .B1(n15806), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15805), .ZN(n10050) );
  AND2_X1 U12021 ( .A1(n10730), .A2(n15634), .ZN(n15623) );
  NAND2_X1 U12022 ( .A1(n15412), .A2(n10922), .ZN(n15513) );
  AOI21_X1 U12023 ( .B1(n9756), .B2(n9913), .A(n9910), .ZN(n9909) );
  INV_X1 U12024 ( .A(n15852), .ZN(n9910) );
  INV_X1 U12025 ( .A(n15412), .ZN(n15515) );
  CLKBUF_X1 U12026 ( .A(n14221), .Z(n15533) );
  AND2_X1 U12027 ( .A1(n13554), .A2(n10031), .ZN(n13865) );
  NAND2_X1 U12028 ( .A1(n13820), .A2(n10091), .ZN(n14072) );
  AND2_X1 U12029 ( .A1(n13554), .A2(n15956), .ZN(n15954) );
  AND2_X1 U12030 ( .A1(n15764), .A2(n10145), .ZN(n10144) );
  INV_X1 U12031 ( .A(n15777), .ZN(n10848) );
  INV_X1 U12032 ( .A(n15778), .ZN(n10849) );
  NAND2_X1 U12033 ( .A1(n9914), .A2(n10841), .ZN(n13993) );
  NAND2_X1 U12034 ( .A1(n9930), .A2(n9929), .ZN(n10831) );
  INV_X1 U12035 ( .A(n13451), .ZN(n9929) );
  INV_X1 U12036 ( .A(n13417), .ZN(n11009) );
  XNOR2_X1 U12037 ( .A(n12956), .B(n10991), .ZN(n13412) );
  AND2_X1 U12038 ( .A1(n10998), .A2(n10997), .ZN(n12810) );
  INV_X1 U12039 ( .A(n15347), .ZN(n19331) );
  CLKBUF_X1 U12040 ( .A(n10783), .Z(n10784) );
  NAND2_X1 U12041 ( .A1(n19549), .A2(n19548), .ZN(n19757) );
  NOR2_X2 U12042 ( .A1(n13715), .A2(n13256), .ZN(n19532) );
  NOR2_X2 U12043 ( .A1(n13716), .A2(n13256), .ZN(n19531) );
  INV_X1 U12044 ( .A(n17726), .ZN(n12344) );
  INV_X1 U12045 ( .A(n19145), .ZN(n19135) );
  OAI22_X1 U12046 ( .A1(n18193), .A2(n18962), .B1(n18956), .B2(n12556), .ZN(
        n18964) );
  NAND2_X1 U12047 ( .A1(n9975), .A2(n9973), .ZN(n9972) );
  INV_X1 U12048 ( .A(n17842), .ZN(n9973) );
  AND2_X1 U12049 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17363), .ZN(n17346) );
  NOR2_X1 U12050 ( .A1(n17498), .A2(n17380), .ZN(n17421) );
  INV_X1 U12051 ( .A(n12324), .ZN(n9883) );
  AOI21_X1 U12052 ( .B1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17472), .A(
        n9882), .ZN(n9881) );
  INV_X1 U12053 ( .A(n12326), .ZN(n9882) );
  INV_X1 U12054 ( .A(n9778), .ZN(n17473) );
  INV_X1 U12055 ( .A(n12196), .ZN(n9893) );
  NAND2_X1 U12056 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n9892) );
  OAI21_X1 U12057 ( .B1(n16214), .B2(n16213), .A(n19128), .ZN(n16215) );
  NAND2_X1 U12058 ( .A1(n16719), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12562) );
  NOR2_X1 U12059 ( .A1(n17837), .A2(n17838), .ZN(n17823) );
  NAND2_X1 U12060 ( .A1(n17987), .A2(n9754), .ZN(n17918) );
  NOR2_X1 U12061 ( .A1(n17960), .A2(n9983), .ZN(n9982) );
  INV_X1 U12062 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9983) );
  NAND2_X1 U12063 ( .A1(n17987), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17959) );
  NOR2_X1 U12064 ( .A1(n18004), .A2(n18006), .ZN(n17987) );
  AOI21_X1 U12065 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17944), .A(
        n18862), .ZN(n18005) );
  NOR2_X1 U12066 ( .A1(n17046), .A2(n17055), .ZN(n18030) );
  NOR2_X1 U12067 ( .A1(n18095), .A2(n18028), .ZN(n18066) );
  INV_X1 U12068 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18028) );
  NAND2_X1 U12069 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n17126), .ZN(
        n18095) );
  AND2_X1 U12070 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17137) );
  NOR2_X1 U12071 ( .A1(n18119), .A2(n18121), .ZN(n18051) );
  NOR2_X1 U12072 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16149), .ZN(
        n16198) );
  NOR3_X1 U12073 ( .A1(n16150), .A2(n16151), .A3(n16713), .ZN(n16199) );
  NOR2_X1 U12074 ( .A1(n17803), .A2(n16201), .ZN(n16709) );
  NOR2_X1 U12075 ( .A1(n17793), .A2(n18956), .ZN(n12462) );
  AOI21_X1 U12076 ( .B1(n18426), .B2(n12441), .A(n12452), .ZN(n10070) );
  NAND2_X1 U12077 ( .A1(n17843), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17803) );
  NOR2_X1 U12078 ( .A1(n17821), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17820) );
  OR2_X1 U12079 ( .A1(n18340), .A2(n9833), .ZN(n17844) );
  NOR2_X1 U12080 ( .A1(n17851), .A2(n18286), .ZN(n18192) );
  AND2_X1 U12081 ( .A1(n17913), .A2(n17900), .ZN(n17938) );
  AOI21_X1 U12082 ( .B1(n17997), .B2(n12432), .A(n10158), .ZN(n17955) );
  AND2_X1 U12083 ( .A1(n17973), .A2(n17997), .ZN(n10158) );
  INV_X1 U12084 ( .A(n18329), .ZN(n18319) );
  NOR2_X1 U12085 ( .A1(n18319), .A2(n18338), .ZN(n18321) );
  NAND2_X1 U12086 ( .A1(n18943), .A2(n18930), .ZN(n18351) );
  NAND2_X1 U12087 ( .A1(n18080), .A2(n9797), .ZN(n18064) );
  XNOR2_X1 U12088 ( .A(n10062), .B(n10061), .ZN(n18094) );
  INV_X1 U12089 ( .A(n12243), .ZN(n10061) );
  XNOR2_X1 U12090 ( .A(n12380), .B(n12379), .ZN(n18102) );
  INV_X1 U12091 ( .A(n12381), .ZN(n12379) );
  NAND2_X1 U12092 ( .A1(n18102), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18101) );
  NAND2_X1 U12093 ( .A1(n9888), .A2(n9889), .ZN(n18113) );
  NAND2_X1 U12094 ( .A1(n9890), .A2(n18128), .ZN(n9888) );
  OR2_X1 U12095 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9890) );
  XNOR2_X1 U12096 ( .A(n12374), .B(n18417), .ZN(n18114) );
  NAND2_X1 U12097 ( .A1(n18113), .A2(n18114), .ZN(n18112) );
  OR2_X1 U12098 ( .A1(n18920), .A2(n12338), .ZN(n16054) );
  OAI21_X2 U12099 ( .B1(n18919), .B2(n18922), .A(n18918), .ZN(n18928) );
  INV_X1 U12100 ( .A(n18193), .ZN(n18961) );
  OAI21_X1 U12101 ( .B1(n12418), .B2(n12412), .A(n12419), .ZN(n16816) );
  OAI211_X1 U12102 ( .C1(n12421), .C2(n12420), .A(n12419), .B(n12418), .ZN(
        n18962) );
  NAND2_X1 U12103 ( .A1(n18160), .A2(n18152), .ZN(n18151) );
  XNOR2_X1 U12104 ( .A(n17670), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18152) );
  NOR2_X1 U12105 ( .A1(n12357), .A2(n9885), .ZN(n12356) );
  AND2_X1 U12106 ( .A1(n12342), .A2(n19132), .ZN(n9885) );
  INV_X1 U12107 ( .A(n12356), .ZN(n18922) );
  INV_X1 U12108 ( .A(n12339), .ZN(n18496) );
  NOR2_X1 U12109 ( .A1(n12284), .A2(n12283), .ZN(n18501) );
  NAND2_X1 U12110 ( .A1(n18986), .A2(n18483), .ZN(n18562) );
  OAI21_X1 U12111 ( .B1(n12798), .B2(n12797), .A(n11291), .ZN(n16176) );
  AOI21_X1 U12112 ( .B1(n14289), .B2(n14288), .A(n14287), .ZN(n20709) );
  INV_X1 U12113 ( .A(n20269), .ZN(n20257) );
  NOR2_X2 U12114 ( .A1(n14892), .A2(n13489), .ZN(n20221) );
  NAND2_X1 U12115 ( .A1(n13486), .A2(n13474), .ZN(n20271) );
  INV_X1 U12116 ( .A(n16272), .ZN(n20263) );
  INV_X1 U12117 ( .A(n20271), .ZN(n16239) );
  OR2_X1 U12118 ( .A1(n13498), .A2(n20233), .ZN(n20272) );
  INV_X1 U12119 ( .A(n14936), .ZN(n20706) );
  NAND2_X1 U12120 ( .A1(n20282), .A2(n14940), .ZN(n14936) );
  INV_X1 U12121 ( .A(n14290), .ZN(n16280) );
  INV_X1 U12122 ( .A(n20321), .ZN(n20297) );
  INV_X2 U12123 ( .A(n20310), .ZN(n20318) );
  CLKBUF_X1 U12124 ( .A(n20296), .Z(n20319) );
  INV_X1 U12125 ( .A(n20346), .ZN(n13200) );
  INV_X1 U12126 ( .A(n14066), .ZN(n20279) );
  INV_X1 U12127 ( .A(n20361), .ZN(n16303) );
  OR2_X1 U12128 ( .A1(n13037), .A2(n16175), .ZN(n20203) );
  INV_X1 U12129 ( .A(n20203), .ZN(n20356) );
  XNOR2_X1 U12130 ( .A(n14992), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15156) );
  NAND2_X1 U12131 ( .A1(n10159), .A2(n14991), .ZN(n14992) );
  NOR2_X1 U12132 ( .A1(n11614), .A2(n15011), .ZN(n11615) );
  XNOR2_X1 U12133 ( .A(n9872), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15185) );
  NOR2_X1 U12134 ( .A1(n15011), .A2(n15019), .ZN(n9872) );
  NAND2_X1 U12135 ( .A1(n15075), .A2(n10122), .ZN(n15076) );
  NOR2_X1 U12136 ( .A1(n10120), .A2(n10119), .ZN(n10123) );
  NAND2_X1 U12137 ( .A1(n20354), .A2(n11522), .ZN(n16322) );
  NAND2_X1 U12138 ( .A1(n13054), .A2(n13045), .ZN(n20392) );
  AND2_X1 U12139 ( .A1(n13054), .A2(n13043), .ZN(n16379) );
  INV_X1 U12140 ( .A(n20392), .ZN(n20374) );
  NAND2_X1 U12141 ( .A1(n13659), .A2(n11577), .ZN(n10126) );
  INV_X1 U12142 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20549) );
  INV_X1 U12143 ( .A(n13659), .ZN(n13246) );
  INV_X1 U12144 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20788) );
  INV_X1 U12145 ( .A(n20400), .ZN(n13349) );
  INV_X1 U12146 ( .A(n12930), .ZN(n15335) );
  INV_X1 U12147 ( .A(n12517), .ZN(n13233) );
  INV_X1 U12148 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20961) );
  NOR2_X1 U12149 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15334) );
  INV_X1 U12150 ( .A(n20401), .ZN(n20417) );
  NOR2_X2 U12151 ( .A1(n20424), .A2(n14149), .ZN(n20443) );
  OAI21_X1 U12152 ( .B1(n20455), .B2(n20486), .A(n20454), .ZN(n20489) );
  NOR2_X2 U12153 ( .A1(n20525), .A2(n14149), .ZN(n20544) );
  NOR2_X1 U12154 ( .A1(n13746), .A2(n13445), .ZN(n20597) );
  INV_X1 U12155 ( .A(n20562), .ZN(n20608) );
  NOR2_X1 U12156 ( .A1(n13286), .A2(n13746), .ZN(n20553) );
  NOR2_X1 U12157 ( .A1(n13293), .A2(n13746), .ZN(n20567) );
  NOR2_X1 U12158 ( .A1(n13307), .A2(n13746), .ZN(n20573) );
  NOR2_X1 U12159 ( .A1(n13579), .A2(n13746), .ZN(n20585) );
  NOR2_X1 U12160 ( .A1(n13357), .A2(n13746), .ZN(n20591) );
  INV_X1 U12161 ( .A(n13780), .ZN(n20598) );
  INV_X1 U12162 ( .A(n14106), .ZN(n14146) );
  INV_X1 U12163 ( .A(n20553), .ZN(n14169) );
  INV_X1 U12164 ( .A(n20573), .ZN(n14185) );
  INV_X1 U12165 ( .A(n20579), .ZN(n14177) );
  INV_X1 U12166 ( .A(n20585), .ZN(n14196) );
  INV_X1 U12167 ( .A(n20591), .ZN(n14189) );
  INV_X1 U12168 ( .A(n20604), .ZN(n14181) );
  INV_X1 U12169 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n20182) );
  NOR2_X1 U12170 ( .A1(n12690), .A2(n12667), .ZN(n20188) );
  NAND2_X1 U12171 ( .A1(n16426), .A2(n16427), .ZN(n16425) );
  NAND2_X1 U12172 ( .A1(n15368), .A2(n15603), .ZN(n16407) );
  NAND2_X1 U12173 ( .A1(n16450), .A2(n16451), .ZN(n16449) );
  NAND2_X1 U12174 ( .A1(n15397), .A2(n15629), .ZN(n15396) );
  OR2_X1 U12175 ( .A1(n10710), .A2(n9822), .ZN(n10713) );
  NAND2_X1 U12176 ( .A1(n15426), .A2(n16494), .ZN(n15425) );
  INV_X1 U12177 ( .A(n19323), .ZN(n19339) );
  INV_X1 U12178 ( .A(n19346), .ZN(n19315) );
  AND2_X1 U12179 ( .A1(n13004), .A2(n12949), .ZN(n15465) );
  INV_X1 U12180 ( .A(n19342), .ZN(n19324) );
  OR2_X1 U12181 ( .A1(n11080), .A2(n11079), .ZN(n13267) );
  NAND2_X1 U12182 ( .A1(n13007), .A2(n13006), .ZN(n13123) );
  AOI21_X1 U12183 ( .B1(n9835), .B2(n15480), .A(n10080), .ZN(n10079) );
  OR2_X1 U12184 ( .A1(n15480), .A2(n14694), .ZN(n10081) );
  AND2_X1 U12185 ( .A1(n13717), .A2(n13716), .ZN(n19356) );
  INV_X1 U12186 ( .A(n15577), .ZN(n16472) );
  OR2_X1 U12187 ( .A1(n16472), .A2(n13717), .ZN(n19376) );
  INV_X1 U12188 ( .A(n20161), .ZN(n19548) );
  AND2_X1 U12189 ( .A1(n12724), .A2(n20178), .ZN(n19458) );
  NOR2_X1 U12190 ( .A1(n12670), .A2(n19514), .ZN(n12717) );
  XNOR2_X1 U12192 ( .A(n13503), .B(n13502), .ZN(n14437) );
  NAND2_X1 U12193 ( .A1(n10024), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10023) );
  INV_X1 U12194 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16542) );
  NAND2_X1 U12195 ( .A1(n12871), .A2(n12865), .ZN(n16541) );
  INV_X1 U12196 ( .A(n16541), .ZN(n19473) );
  AOI21_X1 U12197 ( .B1(n14450), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14449), .ZN(n14451) );
  XNOR2_X1 U12198 ( .A(n10060), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14371) );
  OAI21_X1 U12199 ( .B1(n15923), .B2(n9933), .A(n9931), .ZN(n15933) );
  NOR2_X1 U12200 ( .A1(n16624), .A2(n15924), .ZN(n9933) );
  AND2_X1 U12201 ( .A1(n15945), .A2(n9932), .ZN(n9931) );
  NAND2_X1 U12202 ( .A1(n10962), .A2(n15944), .ZN(n9932) );
  NOR2_X1 U12203 ( .A1(n15988), .A2(n11179), .ZN(n16581) );
  NAND2_X1 U12204 ( .A1(n10147), .A2(n10638), .ZN(n15966) );
  AND2_X1 U12205 ( .A1(n15992), .A2(n11024), .ZN(n16607) );
  CLKBUF_X1 U12206 ( .A(n19461), .Z(n19326) );
  NAND2_X1 U12207 ( .A1(n13446), .A2(n9901), .ZN(n13794) );
  NAND2_X1 U12208 ( .A1(n10100), .A2(n10865), .ZN(n13015) );
  INV_X1 U12209 ( .A(n12831), .ZN(n19492) );
  NAND2_X1 U12210 ( .A1(n10957), .A2(n15925), .ZN(n15952) );
  INV_X1 U12211 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20166) );
  INV_X1 U12212 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20159) );
  AND2_X1 U12213 ( .A1(n12946), .A2(n12834), .ZN(n20153) );
  INV_X1 U12214 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20149) );
  INV_X1 U12215 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20142) );
  INV_X1 U12216 ( .A(n20153), .ZN(n19573) );
  INV_X1 U12217 ( .A(n15465), .ZN(n20145) );
  INV_X1 U12218 ( .A(n16688), .ZN(n16044) );
  INV_X1 U12219 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12700) );
  INV_X1 U12220 ( .A(n19668), .ZN(n19635) );
  NOR2_X1 U12221 ( .A1(n19700), .A2(n19758), .ZN(n19783) );
  NOR2_X1 U12222 ( .A1(n19877), .A2(n19820), .ZN(n19853) );
  OAI21_X1 U12223 ( .B1(n19939), .B2(n19670), .A(n19917), .ZN(n19942) );
  INV_X1 U12224 ( .A(n20016), .ZN(n19973) );
  INV_X1 U12225 ( .A(n20022), .ZN(n19955) );
  INV_X1 U12226 ( .A(n20034), .ZN(n19979) );
  INV_X1 U12227 ( .A(n20040), .ZN(n19983) );
  INV_X1 U12228 ( .A(n20051), .ZN(n19941) );
  INV_X1 U12229 ( .A(n19932), .ZN(n20025) );
  INV_X1 U12230 ( .A(n19935), .ZN(n20031) );
  NAND2_X1 U12231 ( .A1(n19502), .A2(n19994), .ZN(n20050) );
  INV_X1 U12232 ( .A(n19946), .ZN(n20045) );
  INV_X1 U12233 ( .A(n12667), .ZN(n16682) );
  AND2_X1 U12234 ( .A1(n12859), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16688) );
  CLKBUF_X1 U12235 ( .A(n20119), .Z(n20115) );
  NOR2_X1 U12236 ( .A1(n18958), .A2(n17727), .ZN(n19146) );
  INV_X1 U12237 ( .A(n9980), .ZN(n16857) );
  NOR2_X1 U12238 ( .A1(n16902), .A2(n17853), .ZN(n16901) );
  NOR2_X1 U12239 ( .A1(n16910), .A2(n9816), .ZN(n16902) );
  NAND2_X1 U12240 ( .A1(n16719), .A2(n9986), .ZN(n9985) );
  OR2_X1 U12241 ( .A1(n16719), .A2(n16846), .ZN(n9988) );
  NOR2_X1 U12242 ( .A1(n9987), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9986) );
  INV_X1 U12243 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17055) );
  INV_X1 U12244 ( .A(n17199), .ZN(n17185) );
  NAND4_X1 U12245 ( .A1(n18455), .A2(n19126), .A3(n18992), .A4(n18981), .ZN(
        n17199) );
  NOR2_X1 U12246 ( .A1(n16921), .A2(n17259), .ZN(n17264) );
  AND3_X1 U12247 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(n17404), .ZN(n17376) );
  NAND2_X1 U12248 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17376), .ZN(n17375) );
  INV_X1 U12249 ( .A(n17406), .ZN(n17404) );
  NOR2_X1 U12250 ( .A1(n17751), .A2(n17553), .ZN(n17547) );
  NAND2_X1 U12251 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17557), .ZN(n17553) );
  NOR2_X1 U12252 ( .A1(n17733), .A2(n17600), .ZN(n17601) );
  INV_X1 U12253 ( .A(n12368), .ZN(n17665) );
  INV_X1 U12254 ( .A(n17675), .ZN(n17674) );
  INV_X1 U12255 ( .A(n17671), .ZN(n17666) );
  NOR3_X1 U12256 ( .A1(n17678), .A2(n19130), .A3(n17727), .ZN(n17712) );
  NOR2_X1 U12257 ( .A1(n17796), .A2(n17797), .ZN(n16719) );
  NOR2_X1 U12258 ( .A1(n12450), .A2(n12549), .ZN(n17795) );
  NOR2_X1 U12259 ( .A1(n17967), .A2(n9847), .ZN(n17830) );
  NOR2_X1 U12260 ( .A1(n17882), .A2(n12560), .ZN(n17862) );
  INV_X1 U12261 ( .A(n17967), .ZN(n17950) );
  OR2_X1 U12262 ( .A1(n18340), .A2(n9823), .ZN(n18285) );
  OAI21_X1 U12263 ( .B1(n18079), .B2(n18338), .A(n9884), .ZN(n18060) );
  OR2_X1 U12264 ( .A1(n18340), .A2(n18167), .ZN(n9884) );
  NAND2_X1 U12265 ( .A1(n17648), .A2(n18131), .ZN(n18079) );
  NOR2_X1 U12266 ( .A1(n18083), .A2(n18069), .ZN(n18067) );
  INV_X1 U12267 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18069) );
  INV_X1 U12268 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18083) );
  NAND2_X1 U12269 ( .A1(n17137), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18107) );
  INV_X1 U12270 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17152) );
  NOR2_X1 U12271 ( .A1(n16819), .A2(n19132), .ZN(n18131) );
  INV_X1 U12272 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18150) );
  NOR2_X1 U12273 ( .A1(n17944), .A2(n17943), .ZN(n18146) );
  OR2_X1 U12274 ( .A1(n18722), .A2(n18562), .ZN(n18826) );
  INV_X1 U12275 ( .A(n18167), .ZN(n18154) );
  INV_X1 U12276 ( .A(n18146), .ZN(n18156) );
  INV_X1 U12277 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19088) );
  NOR2_X1 U12278 ( .A1(n17804), .A2(n16201), .ZN(n16712) );
  NAND2_X1 U12279 ( .A1(n17913), .A2(n12440), .ZN(n17850) );
  NOR2_X1 U12280 ( .A1(n18304), .A2(n17994), .ZN(n18287) );
  NAND2_X1 U12281 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18287), .ZN(
        n18286) );
  INV_X1 U12282 ( .A(n18351), .ZN(n18323) );
  INV_X1 U12283 ( .A(n18339), .ZN(n18376) );
  INV_X1 U12284 ( .A(n10063), .ZN(n18103) );
  INV_X1 U12285 ( .A(n10066), .ZN(n18132) );
  NAND2_X1 U12286 ( .A1(n12356), .A2(n18923), .ZN(n18947) );
  INV_X1 U12287 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18938) );
  AOI211_X1 U12288 ( .C1(n19128), .C2(n18945), .A(n18484), .B(n16139), .ZN(
        n19110) );
  INV_X1 U12289 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16143) );
  CLKBUF_X1 U12290 ( .A(n16806), .Z(n16804) );
  OAI21_X1 U12291 ( .B1(n15824), .B2(n16514), .A(n9920), .ZN(P2_U2988) );
  AOI21_X1 U12292 ( .B1(n16442), .B2(n19480), .A(n15622), .ZN(n9922) );
  AOI21_X1 U12293 ( .B1(n15592), .B2(n16624), .A(n11204), .ZN(n11222) );
  INV_X1 U12294 ( .A(n10045), .ZN(n10044) );
  INV_X1 U12295 ( .A(n9978), .ZN(n16844) );
  OAI21_X1 U12296 ( .B1(n12589), .B2(n18167), .A(n12569), .ZN(n12570) );
  OAI21_X1 U12297 ( .B1(n12589), .B2(n16147), .A(n12588), .ZN(n12590) );
  AOI21_X1 U12298 ( .B1(n12448), .B2(n18438), .A(n12447), .ZN(n12449) );
  OAI21_X1 U12299 ( .B1(n17819), .B2(n18358), .A(n12446), .ZN(n12447) );
  AND2_X1 U12300 ( .A1(n13002), .A2(n13011), .ZN(n13062) );
  INV_X1 U12301 ( .A(n10278), .ZN(n11199) );
  NAND2_X1 U12302 ( .A1(n13872), .A2(n13956), .ZN(n13955) );
  OR3_X1 U12303 ( .A1(n15423), .A2(n11020), .A3(n10715), .ZN(n9752) );
  AND2_X1 U12304 ( .A1(n14824), .A2(n9811), .ZN(n14797) );
  NAND2_X1 U12305 ( .A1(n10171), .A2(n10028), .ZN(n15400) );
  NAND2_X1 U12306 ( .A1(n15709), .A2(n15901), .ZN(n9753) );
  NOR2_X1 U12307 ( .A1(n15633), .A2(n15634), .ZN(n15620) );
  AND2_X1 U12308 ( .A1(n9982), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9754) );
  AND2_X1 U12309 ( .A1(n10002), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9755) );
  NAND4_X1 U12310 ( .A1(n15658), .A2(n10706), .A3(n15674), .A4(n15695), .ZN(
        n9756) );
  OAI21_X1 U12311 ( .B1(n11367), .B2(n11365), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11441) );
  AND2_X1 U12312 ( .A1(n11024), .A2(n16608), .ZN(n9757) );
  AND4_X1 U12313 ( .A1(n9893), .A2(n12198), .A3(n12197), .A4(n9892), .ZN(n9758) );
  AND2_X1 U12314 ( .A1(n10011), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9759) );
  AND2_X1 U12315 ( .A1(n10390), .A2(n10389), .ZN(n9760) );
  AND2_X1 U12316 ( .A1(n10845), .A2(n15984), .ZN(n9761) );
  NOR2_X1 U12317 ( .A1(n16843), .A2(n9979), .ZN(n9762) );
  AND2_X1 U12318 ( .A1(n10091), .A2(n10090), .ZN(n9763) );
  AND2_X1 U12319 ( .A1(n15097), .A2(n9844), .ZN(n9764) );
  AND2_X1 U12320 ( .A1(n10628), .A2(n9813), .ZN(n9765) );
  AND2_X1 U12321 ( .A1(n9754), .A2(n9981), .ZN(n9766) );
  NAND2_X1 U12322 ( .A1(n15992), .A2(n9757), .ZN(n15973) );
  NAND2_X1 U12323 ( .A1(n18916), .A2(n18323), .ZN(n18370) );
  INV_X1 U12324 ( .A(n18370), .ZN(n9886) );
  OR2_X1 U12325 ( .A1(n14924), .A2(n14842), .ZN(n9767) );
  AND2_X1 U12326 ( .A1(n13956), .A2(n11887), .ZN(n9768) );
  AND2_X1 U12327 ( .A1(n10006), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n9769) );
  AND2_X1 U12328 ( .A1(n13906), .A2(n9846), .ZN(n9770) );
  AND2_X1 U12329 ( .A1(n10143), .A2(n9830), .ZN(n9771) );
  NAND2_X1 U12330 ( .A1(n15646), .A2(n15754), .ZN(n9772) );
  OR2_X1 U12331 ( .A1(n9974), .A2(n9976), .ZN(n9773) );
  OR3_X1 U12332 ( .A1(n13809), .A2(n9955), .A3(n13808), .ZN(n13965) );
  OR2_X1 U12333 ( .A1(n9823), .A2(n17851), .ZN(n9774) );
  AND2_X2 U12334 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12893) );
  OR2_X1 U12335 ( .A1(n15634), .A2(n10929), .ZN(n9775) );
  AND2_X2 U12336 ( .A1(n10240), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10456) );
  NAND2_X1 U12337 ( .A1(n12655), .A2(n14570), .ZN(n10854) );
  OR3_X1 U12338 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19085), .A3(
        n18948), .ZN(n9778) );
  INV_X1 U12339 ( .A(n11291), .ZN(n14940) );
  AND2_X1 U12340 ( .A1(n9940), .A2(n9938), .ZN(n9779) );
  NAND2_X1 U12341 ( .A1(n10629), .A2(n9765), .ZN(n10147) );
  OR3_X1 U12342 ( .A1(n15633), .A2(n9775), .A3(n10023), .ZN(n9780) );
  OR3_X1 U12343 ( .A1(n15379), .A2(n10095), .A3(n10093), .ZN(n9781) );
  INV_X1 U12344 ( .A(n10278), .ZN(n10212) );
  XNOR2_X1 U12345 ( .A(n9781), .B(n14435), .ZN(n14462) );
  INV_X1 U12346 ( .A(n9862), .ZN(n11678) );
  NAND2_X1 U12347 ( .A1(n13577), .A2(n11352), .ZN(n9862) );
  AND2_X1 U12348 ( .A1(n10133), .A2(n15097), .ZN(n9782) );
  NAND2_X1 U12349 ( .A1(n14824), .A2(n9970), .ZN(n14782) );
  NAND2_X1 U12350 ( .A1(n14824), .A2(n12073), .ZN(n14808) );
  NOR2_X1 U12351 ( .A1(n18340), .A2(n18303), .ZN(n9783) );
  OR2_X1 U12352 ( .A1(n11166), .A2(n11167), .ZN(n9784) );
  OR2_X1 U12353 ( .A1(n15481), .A2(n15480), .ZN(n9785) );
  INV_X2 U12354 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16039) );
  OR2_X1 U12355 ( .A1(n12140), .A2(n18921), .ZN(n9786) );
  AND3_X1 U12356 ( .A1(n13443), .A2(n14238), .A3(n13442), .ZN(n13617) );
  AND2_X1 U12357 ( .A1(n10147), .A2(n10145), .ZN(n15761) );
  OR2_X1 U12358 ( .A1(n11166), .A2(n10019), .ZN(n9787) );
  OR2_X1 U12359 ( .A1(n11797), .A2(n11943), .ZN(n9788) );
  OR2_X1 U12360 ( .A1(n10288), .A2(n19503), .ZN(n9789) );
  NOR2_X1 U12361 ( .A1(n18340), .A2(n9774), .ZN(n9790) );
  NAND2_X1 U12362 ( .A1(n13062), .A2(n13063), .ZN(n13007) );
  AOI21_X1 U12363 ( .B1(n15738), .B2(n10707), .A(n9756), .ZN(n15850) );
  NAND2_X1 U12364 ( .A1(n10141), .A2(n10142), .ZN(n15738) );
  AND2_X1 U12365 ( .A1(n15645), .A2(n15646), .ZN(n15752) );
  AND2_X1 U12366 ( .A1(n10716), .A2(n9752), .ZN(n9791) );
  AND4_X1 U12367 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n9792) );
  AND2_X1 U12368 ( .A1(n15709), .A2(n9919), .ZN(n15666) );
  AND4_X1 U12369 ( .A1(n10553), .A2(n10552), .A3(n10551), .A4(n10550), .ZN(
        n9793) );
  AND2_X1 U12370 ( .A1(n10950), .A2(n10273), .ZN(n10312) );
  NAND2_X1 U12371 ( .A1(n9905), .A2(n9907), .ZN(n15616) );
  NAND2_X1 U12372 ( .A1(n9787), .A2(n10021), .ZN(n16416) );
  AND2_X1 U12373 ( .A1(n11479), .A2(n11478), .ZN(n9794) );
  INV_X1 U12374 ( .A(n10650), .ZN(n16501) );
  OR2_X1 U12375 ( .A1(n12235), .A2(n12392), .ZN(n9795) );
  NAND2_X1 U12376 ( .A1(n13457), .A2(n11476), .ZN(n11502) );
  AND2_X1 U12377 ( .A1(n10463), .A2(n9917), .ZN(n9796) );
  AND2_X1 U12378 ( .A1(n12391), .A2(n20850), .ZN(n9797) );
  OR2_X1 U12379 ( .A1(n12240), .A2(n10064), .ZN(n9798) );
  NOR2_X1 U12380 ( .A1(n11601), .A2(n14053), .ZN(n9799) );
  AND2_X1 U12381 ( .A1(n14230), .A2(n14229), .ZN(n9800) );
  NOR2_X1 U12382 ( .A1(n15513), .A2(n15399), .ZN(n15398) );
  OR2_X1 U12383 ( .A1(n11613), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9801) );
  AND2_X1 U12384 ( .A1(n10171), .A2(n15416), .ZN(n15415) );
  NAND2_X1 U12385 ( .A1(n10327), .A2(n10326), .ZN(n10353) );
  AND2_X1 U12386 ( .A1(n10379), .A2(n10378), .ZN(n9802) );
  NAND2_X1 U12387 ( .A1(n15139), .A2(n11595), .ZN(n15095) );
  OR2_X1 U12388 ( .A1(n10838), .A2(n10839), .ZN(n9803) );
  INV_X1 U12389 ( .A(n9908), .ZN(n9907) );
  NOR2_X1 U12390 ( .A1(n15637), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9908) );
  NOR2_X1 U12391 ( .A1(n15535), .A2(n10101), .ZN(n15412) );
  INV_X1 U12392 ( .A(n11359), .ZN(n9867) );
  NAND2_X1 U12393 ( .A1(n11371), .A2(n11352), .ZN(n11359) );
  NAND2_X1 U12394 ( .A1(n9911), .A2(n9909), .ZN(n16480) );
  OR2_X1 U12395 ( .A1(n15808), .A2(n19490), .ZN(n9805) );
  OR2_X1 U12396 ( .A1(n10720), .A2(n15840), .ZN(n9806) );
  INV_X1 U12397 ( .A(n11546), .ZN(n10109) );
  AND2_X2 U12398 ( .A1(n11234), .A2(n12893), .ZN(n11386) );
  NAND2_X1 U12399 ( .A1(n19514), .A2(n19670), .ZN(n11038) );
  INV_X1 U12400 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10118) );
  INV_X1 U12401 ( .A(n12376), .ZN(n9891) );
  NAND2_X1 U12402 ( .A1(n14770), .A2(n14771), .ZN(n14757) );
  NAND2_X1 U12403 ( .A1(n13554), .A2(n10030), .ZN(n13863) );
  NOR2_X1 U12404 ( .A1(n13537), .A2(n13538), .ZN(n13536) );
  NAND2_X1 U12405 ( .A1(n13820), .A2(n13819), .ZN(n13818) );
  AND2_X1 U12406 ( .A1(n13534), .A2(n10002), .ZN(n9807) );
  NOR2_X2 U12407 ( .A1(n17648), .A2(n12451), .ZN(n18075) );
  NAND2_X1 U12408 ( .A1(n15097), .A2(n14374), .ZN(n9808) );
  AND2_X1 U12409 ( .A1(n13786), .A2(n13873), .ZN(n13872) );
  AND2_X1 U12410 ( .A1(n13820), .A2(n10089), .ZN(n14198) );
  AND2_X1 U12411 ( .A1(n13820), .A2(n9763), .ZN(n9809) );
  INV_X1 U12412 ( .A(n15851), .ZN(n9913) );
  NAND2_X1 U12413 ( .A1(n9878), .A2(n11572), .ZN(n16314) );
  NAND2_X1 U12414 ( .A1(n9871), .A2(n11594), .ZN(n14052) );
  AND2_X1 U12415 ( .A1(n14934), .A2(n14933), .ZN(n14863) );
  AND3_X1 U12416 ( .A1(n11358), .A2(n11371), .A3(n13136), .ZN(n12786) );
  INV_X1 U12417 ( .A(n14862), .ZN(n9946) );
  OR3_X1 U12418 ( .A1(n15535), .A2(n10103), .A3(n15440), .ZN(n9810) );
  INV_X1 U12419 ( .A(n11611), .ZN(n10120) );
  NAND2_X1 U12420 ( .A1(n16322), .A2(n16321), .ZN(n16320) );
  AND2_X1 U12421 ( .A1(n10276), .A2(n10288), .ZN(n10796) );
  AND2_X1 U12422 ( .A1(n12073), .A2(n9971), .ZN(n9811) );
  OR2_X1 U12423 ( .A1(n17946), .A2(n18075), .ZN(n17913) );
  NAND2_X1 U12424 ( .A1(n13405), .A2(n13404), .ZN(n13403) );
  AND2_X1 U12425 ( .A1(n13956), .A2(n11899), .ZN(n9812) );
  AND2_X1 U12426 ( .A1(n15773), .A2(n15982), .ZN(n9813) );
  INV_X1 U12427 ( .A(n14924), .ZN(n9949) );
  AND2_X1 U12428 ( .A1(n10030), .A2(n10029), .ZN(n9814) );
  AND2_X1 U12429 ( .A1(n10086), .A2(n15530), .ZN(n9815) );
  INV_X1 U12430 ( .A(n13436), .ZN(n11837) );
  INV_X1 U12432 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16528) );
  NAND2_X1 U12433 ( .A1(n9779), .A2(n10579), .ZN(n9939) );
  INV_X1 U12434 ( .A(n10129), .ZN(n10128) );
  NAND2_X1 U12435 ( .A1(n11393), .A2(n13479), .ZN(n10129) );
  AND2_X1 U12436 ( .A1(n14795), .A2(n14784), .ZN(n14770) );
  NAND2_X1 U12437 ( .A1(n14215), .A2(n10006), .ZN(n10009) );
  AND2_X1 U12438 ( .A1(n9757), .A2(n15975), .ZN(n9817) );
  AND2_X1 U12439 ( .A1(n9969), .A2(n9970), .ZN(n9818) );
  AND2_X1 U12440 ( .A1(n9966), .A2(n9965), .ZN(n9819) );
  OR2_X1 U12441 ( .A1(n10538), .A2(n10537), .ZN(n10542) );
  INV_X1 U12442 ( .A(n10486), .ZN(n11020) );
  NOR2_X1 U12444 ( .A1(n15309), .A2(n15308), .ZN(n9820) );
  AND2_X1 U12445 ( .A1(n13192), .A2(n13191), .ZN(n13467) );
  NAND2_X1 U12446 ( .A1(n13907), .A2(n13906), .ZN(n13979) );
  AND2_X1 U12447 ( .A1(n13418), .A2(n13421), .ZN(n13419) );
  NOR2_X1 U12448 ( .A1(n13068), .A2(n13069), .ZN(n13067) );
  INV_X1 U12449 ( .A(n17919), .ZN(n9981) );
  INV_X2 U12450 ( .A(n17171), .ZN(n9816) );
  INV_X1 U12451 ( .A(n18075), .ZN(n17997) );
  NOR2_X1 U12452 ( .A1(n13809), .A2(n13808), .ZN(n9821) );
  NAND2_X1 U12453 ( .A1(n11197), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n9822) );
  OR2_X1 U12454 ( .A1(n18303), .A2(n18298), .ZN(n9823) );
  INV_X1 U12455 ( .A(n10655), .ZN(n9942) );
  NAND2_X1 U12456 ( .A1(n13999), .A2(n11021), .ZN(n15992) );
  NOR2_X1 U12457 ( .A1(n13345), .A2(n13344), .ZN(n9824) );
  NOR2_X2 U12458 ( .A1(n12263), .A2(n12262), .ZN(n19132) );
  NOR2_X1 U12459 ( .A1(n13415), .A2(n11009), .ZN(n13418) );
  NAND2_X1 U12460 ( .A1(n13508), .A2(n11018), .ZN(n13998) );
  AND2_X1 U12461 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n9825) );
  AND2_X1 U12462 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n9826)
         );
  AND2_X1 U12463 ( .A1(n13907), .A2(n10086), .ZN(n9827) );
  AND2_X1 U12464 ( .A1(n10126), .A2(n11431), .ZN(n9828) );
  NAND2_X1 U12465 ( .A1(n11197), .A2(n10664), .ZN(n9829) );
  INV_X1 U12466 ( .A(n10041), .ZN(n16018) );
  INV_X1 U12467 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10064) );
  NAND2_X1 U12468 ( .A1(n15363), .A2(n9995), .ZN(n10000) );
  NOR2_X1 U12469 ( .A1(n13809), .A2(n9954), .ZN(n14237) );
  INV_X1 U12470 ( .A(n15343), .ZN(n10094) );
  AND2_X1 U12471 ( .A1(n10658), .A2(n16571), .ZN(n15753) );
  INV_X1 U12472 ( .A(n15753), .ZN(n10143) );
  INV_X1 U12473 ( .A(n9976), .ZN(n9975) );
  NOR2_X1 U12474 ( .A1(n9816), .A2(n9977), .ZN(n9976) );
  NAND2_X1 U12475 ( .A1(n10651), .A2(n16594), .ZN(n9830) );
  INV_X1 U12476 ( .A(n9996), .ZN(n9995) );
  NAND2_X1 U12477 ( .A1(n9997), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9996) );
  AND2_X1 U12478 ( .A1(n14286), .A2(n14257), .ZN(n9831) );
  AND2_X1 U12479 ( .A1(n10026), .A2(n10025), .ZN(n9832) );
  OR2_X1 U12480 ( .A1(n9774), .A2(n9895), .ZN(n9833) );
  INV_X1 U12481 ( .A(n20691), .ZN(n20693) );
  NAND2_X2 U12482 ( .A1(n12770), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20691) );
  NAND2_X1 U12483 ( .A1(n11231), .A2(n12893), .ZN(n12901) );
  AND2_X1 U12484 ( .A1(n16719), .A2(n9991), .ZN(n9834) );
  NOR2_X1 U12485 ( .A1(n14675), .A2(n10082), .ZN(n9835) );
  AND2_X1 U12486 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n9836) );
  AND2_X1 U12487 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n9837)
         );
  AND2_X1 U12488 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n9838)
         );
  AND2_X1 U12489 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n9839) );
  AND2_X1 U12490 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n9840)
         );
  AND2_X1 U12491 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n9841) );
  OR2_X1 U12492 ( .A1(n17101), .A2(n16849), .ZN(n9842) );
  AND2_X1 U12493 ( .A1(n11214), .A2(n14441), .ZN(n9843) );
  OR2_X1 U12494 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9844) );
  INV_X1 U12495 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9992) );
  INV_X1 U12496 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10012) );
  INV_X1 U12497 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10008) );
  AND2_X1 U12498 ( .A1(n17987), .A2(n9982), .ZN(n9845) );
  OR2_X1 U12499 ( .A1(n13978), .A2(n13977), .ZN(n9846) );
  OR3_X1 U12500 ( .A1(n17851), .A2(n18191), .A3(n9895), .ZN(n9847) );
  AND2_X1 U12501 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9848)
         );
  AND2_X1 U12502 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n9849) );
  AND2_X1 U12503 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n9850)
         );
  AND2_X1 U12504 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n9851) );
  AND2_X1 U12505 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n9852) );
  AND2_X1 U12506 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n9853)
         );
  AND2_X1 U12507 ( .A1(n9919), .A2(n11181), .ZN(n9854) );
  AND2_X1 U12508 ( .A1(n10059), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9855) );
  AND2_X1 U12509 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n9856) );
  INV_X1 U12510 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9895) );
  INV_X1 U12511 ( .A(n14694), .ZN(n10082) );
  INV_X1 U12512 ( .A(n14456), .ZN(n10024) );
  INV_X1 U12513 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n9993) );
  INV_X1 U12514 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9984) );
  INV_X1 U12515 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9999) );
  INV_X1 U12516 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10007) );
  INV_X1 U12517 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10004) );
  INV_X1 U12518 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10003) );
  NAND3_X2 U12519 ( .A1(n18986), .A2(n19143), .A3(n19144), .ZN(n18455) );
  NOR2_X1 U12520 ( .A1(n13578), .A2(n13292), .ZN(n9857) );
  NAND2_X1 U12521 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13239), .ZN(n13578) );
  AOI222_X1 U12522 ( .A1(n9720), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20669), .ZN(n20640) );
  AOI222_X1 U12523 ( .A1(n9720), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20669), .ZN(n20638) );
  AOI222_X1 U12524 ( .A1(n9720), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20669), .ZN(n20636) );
  INV_X1 U12525 ( .A(n17184), .ZN(n18992) );
  NOR4_X2 U12526 ( .A1(n20214), .A2(n20213), .A3(n20212), .A4(n20211), .ZN(
        n20687) );
  NOR4_X2 U12527 ( .A1(n16138), .A2(n16214), .A3(n16137), .A4(n16136), .ZN(
        n18966) );
  AND2_X4 U12528 ( .A1(n12893), .A2(n11232), .ZN(n12489) );
  NOR2_X1 U12529 ( .A1(n13456), .A2(n9858), .ZN(n20387) );
  NAND2_X1 U12530 ( .A1(n11474), .A2(n11473), .ZN(n9858) );
  INV_X2 U12531 ( .A(n11371), .ZN(n11360) );
  INV_X2 U12532 ( .A(n11348), .ZN(n13577) );
  INV_X1 U12533 ( .A(n11292), .ZN(n9868) );
  INV_X1 U12534 ( .A(n11449), .ZN(n12611) );
  AND2_X1 U12535 ( .A1(n12903), .A2(n12893), .ZN(n11552) );
  NAND2_X2 U12536 ( .A1(n20282), .A2(n11291), .ZN(n14939) );
  OAI21_X2 U12537 ( .B1(n15703), .B2(n15704), .A(n15654), .ZN(n15698) );
  NAND2_X2 U12538 ( .A1(n9875), .A2(n15651), .ZN(n15703) );
  OR2_X2 U12539 ( .A1(n15714), .A2(n15713), .ZN(n9875) );
  OAI21_X2 U12540 ( .B1(n15723), .B2(n15650), .A(n15722), .ZN(n15714) );
  OAI21_X2 U12541 ( .B1(n15732), .B2(n15649), .A(n15729), .ZN(n15723) );
  NAND2_X1 U12542 ( .A1(n13446), .A2(n9876), .ZN(n13448) );
  NAND2_X1 U12543 ( .A1(n10521), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9876) );
  NAND2_X1 U12544 ( .A1(n10134), .A2(n15139), .ZN(n10135) );
  NAND3_X1 U12545 ( .A1(n10107), .A2(n10105), .A3(n11571), .ZN(n9878) );
  AND2_X2 U12546 ( .A1(n10147), .A2(n10144), .ZN(n10650) );
  OAI21_X2 U12547 ( .B1(n9879), .B2(n9918), .A(n10815), .ZN(n10816) );
  AND2_X2 U12548 ( .A1(n10404), .A2(n10403), .ZN(n9918) );
  INV_X2 U12549 ( .A(n17647), .ZN(n18516) );
  OR2_X2 U12550 ( .A1(n9880), .A2(n12323), .ZN(n17647) );
  NAND3_X1 U12551 ( .A1(n9883), .A2(n9881), .A3(n12325), .ZN(n9880) );
  INV_X2 U12552 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n19085) );
  INV_X2 U12553 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n19103) );
  INV_X2 U12554 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n19109) );
  NAND2_X2 U12555 ( .A1(n9886), .A2(n19132), .ZN(n18193) );
  OAI21_X1 U12556 ( .B1(n18144), .B2(n9887), .A(n18143), .ZN(n18442) );
  NAND2_X1 U12557 ( .A1(n18144), .A2(n9887), .ZN(n18143) );
  XNOR2_X1 U12558 ( .A(n12370), .B(n18436), .ZN(n9887) );
  NOR2_X1 U12559 ( .A1(n18128), .A2(n18129), .ZN(n18127) );
  NAND2_X1 U12560 ( .A1(n18129), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9889) );
  NOR3_X2 U12561 ( .A1(n17938), .A2(n17849), .A3(n18200), .ZN(n17833) );
  NOR2_X1 U12562 ( .A1(n12445), .A2(n17997), .ZN(n12450) );
  NAND2_X1 U12563 ( .A1(n9899), .A2(n9902), .ZN(n16537) );
  NAND3_X1 U12564 ( .A1(n9901), .A2(n13446), .A3(n9900), .ZN(n9899) );
  NAND2_X1 U12565 ( .A1(n16537), .A2(n16536), .ZN(n10587) );
  NAND2_X1 U12566 ( .A1(n10716), .A2(n9903), .ZN(n9905) );
  NAND2_X1 U12567 ( .A1(n15738), .A2(n9912), .ZN(n9911) );
  OAI21_X2 U12568 ( .B1(n10816), .B2(n10626), .A(n13607), .ZN(n10521) );
  NAND2_X1 U12569 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  OR2_X1 U12570 ( .A1(n10842), .A2(n10838), .ZN(n9915) );
  NAND2_X1 U12571 ( .A1(n9803), .A2(n10842), .ZN(n9916) );
  AND2_X1 U12572 ( .A1(n10825), .A2(n10542), .ZN(n9917) );
  NAND2_X2 U12573 ( .A1(n15780), .A2(n10851), .ZN(n15709) );
  INV_X1 U12574 ( .A(n9921), .ZN(n9920) );
  OAI21_X1 U12575 ( .B1(n15820), .B2(n19464), .A(n9922), .ZN(n9921) );
  NAND2_X1 U12576 ( .A1(n9925), .A2(n10861), .ZN(n10100) );
  XNOR2_X2 U12577 ( .A(n9925), .B(n10861), .ZN(n10374) );
  NAND2_X1 U12578 ( .A1(n9927), .A2(n9926), .ZN(n15778) );
  NAND2_X1 U12579 ( .A1(n9928), .A2(n15985), .ZN(n9927) );
  OAI21_X1 U12580 ( .B1(n10057), .B2(n13993), .A(n10056), .ZN(n9928) );
  NAND2_X1 U12581 ( .A1(n13992), .A2(n10845), .ZN(n15987) );
  NOR2_X2 U12582 ( .A1(n15717), .A2(n15710), .ZN(n15923) );
  AND3_X4 U12583 ( .A1(n16647), .A2(n10088), .A3(n9935), .ZN(n10187) );
  MUX2_X1 U12584 ( .A(n16006), .B(n16036), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n16001) );
  AND2_X2 U12585 ( .A1(n9738), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10438) );
  INV_X1 U12586 ( .A(n9939), .ZN(n10635) );
  NAND2_X1 U12587 ( .A1(n9943), .A2(n10691), .ZN(n10692) );
  NAND2_X1 U12588 ( .A1(n9943), .A2(n10657), .ZN(n19248) );
  NAND2_X1 U12589 ( .A1(n11351), .A2(n12517), .ZN(n13041) );
  OR2_X2 U12590 ( .A1(n11354), .A2(n13041), .ZN(n11367) );
  NAND2_X1 U12591 ( .A1(n11525), .A2(n9960), .ZN(n11564) );
  INV_X1 U12592 ( .A(n11524), .ZN(n9961) );
  NAND2_X1 U12594 ( .A1(n14740), .A2(n9966), .ZN(n14708) );
  AND2_X1 U12595 ( .A1(n14740), .A2(n9967), .ZN(n12488) );
  NAND2_X1 U12596 ( .A1(n14740), .A2(n14742), .ZN(n12130) );
  AND2_X2 U12597 ( .A1(n14740), .A2(n9819), .ZN(n14709) );
  AND2_X2 U12598 ( .A1(n14824), .A2(n9818), .ZN(n14773) );
  NOR2_X1 U12599 ( .A1(n9974), .A2(n9972), .ZN(n16894) );
  OAI211_X2 U12600 ( .C1(n9989), .C2(n16846), .A(n9988), .B(n9985), .ZN(n17171) );
  INV_X1 U12601 ( .A(n10000), .ZN(n15366) );
  INV_X1 U12602 ( .A(n10009), .ZN(n15354) );
  NAND3_X1 U12603 ( .A1(n10010), .A2(n9759), .A3(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13531) );
  NAND3_X1 U12604 ( .A1(n10433), .A2(n10016), .A3(n10015), .ZN(n10014) );
  NOR2_X2 U12605 ( .A1(n15667), .A2(n16543), .ZN(n15641) );
  OAI21_X1 U12606 ( .B1(n11166), .B2(n10017), .A(n14446), .ZN(n10021) );
  NOR3_X2 U12607 ( .A1(n11166), .A2(n11167), .A3(n15370), .ZN(n15369) );
  NOR3_X1 U12608 ( .A1(n15633), .A2(n14456), .A3(n9775), .ZN(n15600) );
  INV_X2 U12609 ( .A(n10766), .ZN(n10941) );
  NAND2_X1 U12611 ( .A1(n10033), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10032) );
  NAND4_X1 U12612 ( .A1(n10264), .A2(n10261), .A3(n10262), .A4(n10263), .ZN(
        n10033) );
  NAND2_X1 U12613 ( .A1(n10035), .A2(n16039), .ZN(n10034) );
  NAND4_X1 U12614 ( .A1(n10260), .A2(n10257), .A3(n10258), .A4(n10259), .ZN(
        n10035) );
  XNOR2_X1 U12615 ( .A(n10036), .B(n10588), .ZN(n10836) );
  NAND4_X1 U12616 ( .A1(n10252), .A2(n10251), .A3(n10249), .A4(n10250), .ZN(
        n10038) );
  NAND4_X1 U12617 ( .A1(n10256), .A2(n10255), .A3(n10253), .A4(n10254), .ZN(
        n10040) );
  NAND3_X1 U12618 ( .A1(n10946), .A2(n10043), .A3(n10298), .ZN(n10041) );
  INV_X2 U12619 ( .A(n10502), .ZN(n10043) );
  NAND2_X1 U12620 ( .A1(n10051), .A2(n10044), .ZN(P2_U3019) );
  OAI21_X1 U12621 ( .B1(n15809), .B2(n9805), .A(n10046), .ZN(n10045) );
  NAND2_X2 U12622 ( .A1(n10849), .A2(n10848), .ZN(n15780) );
  NAND2_X2 U12623 ( .A1(n15641), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15633) );
  NAND4_X1 U12624 ( .A1(n10248), .A2(n10245), .A3(n10246), .A4(n10247), .ZN(
        n10053) );
  NAND4_X1 U12625 ( .A1(n10244), .A2(n10241), .A3(n10242), .A4(n10243), .ZN(
        n10055) );
  NAND2_X1 U12626 ( .A1(n10071), .A2(n16683), .ZN(n10297) );
  NAND2_X1 U12627 ( .A1(n15498), .A2(n15497), .ZN(n15496) );
  NAND2_X1 U12628 ( .A1(n15496), .A2(n10073), .ZN(n10075) );
  NAND3_X1 U12629 ( .A1(n15496), .A2(n10073), .A3(n10072), .ZN(n10074) );
  NAND2_X1 U12630 ( .A1(n14628), .A2(n10074), .ZN(n15493) );
  NAND2_X1 U12631 ( .A1(n10075), .A2(n14625), .ZN(n14628) );
  INV_X1 U12632 ( .A(n14602), .ZN(n10076) );
  AND2_X1 U12633 ( .A1(n10276), .A2(n10941), .ZN(n10265) );
  NAND2_X2 U12634 ( .A1(n10185), .A2(n10184), .ZN(n10305) );
  AND3_X4 U12635 ( .A1(n10487), .A2(n10077), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14684) );
  NAND2_X1 U12636 ( .A1(n15481), .A2(n9835), .ZN(n10078) );
  OAI211_X1 U12637 ( .C1(n15481), .C2(n10081), .A(n10079), .B(n10078), .ZN(
        n14703) );
  OAI21_X1 U12638 ( .B1(n14703), .B2(n15539), .A(n14702), .ZN(P2_U2857) );
  NAND2_X1 U12639 ( .A1(n10084), .A2(n10083), .ZN(n13192) );
  NAND4_X1 U12640 ( .A1(n13002), .A2(n13011), .A3(n13063), .A4(n13122), .ZN(
        n10084) );
  INV_X2 U12641 ( .A(n10267), .ZN(n10287) );
  AND2_X2 U12642 ( .A1(n10941), .A2(n10267), .ZN(n10279) );
  INV_X1 U12643 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10088) );
  NAND3_X1 U12644 ( .A1(n10098), .A2(n13020), .A3(n10100), .ZN(n13068) );
  NOR2_X1 U12645 ( .A1(n15535), .A2(n15440), .ZN(n15442) );
  INV_X1 U12646 ( .A(n15427), .ZN(n10103) );
  OAI21_X1 U12647 ( .B1(n20354), .B2(n10106), .A(n10104), .ZN(n13723) );
  AOI21_X1 U12648 ( .B1(n16321), .B2(n10110), .A(n10109), .ZN(n10104) );
  NAND2_X1 U12649 ( .A1(n10106), .A2(n11546), .ZN(n10105) );
  INV_X1 U12650 ( .A(n16321), .ZN(n10106) );
  NOR2_X1 U12651 ( .A1(n10109), .A2(n10110), .ZN(n10108) );
  NAND2_X1 U12652 ( .A1(n10123), .A2(n15097), .ZN(n10122) );
  OAI21_X1 U12653 ( .B1(n11381), .B2(n10129), .A(n10124), .ZN(n11433) );
  OAI21_X2 U12654 ( .B1(n13659), .B2(n11430), .A(n10127), .ZN(n11432) );
  NAND2_X1 U12655 ( .A1(n14377), .A2(n15009), .ZN(n14989) );
  NAND4_X1 U12656 ( .A1(n10280), .A2(n10300), .A3(n19503), .A4(n10279), .ZN(
        n16686) );
  NAND2_X1 U12657 ( .A1(n9732), .A2(n10628), .ZN(n15771) );
  INV_X1 U12658 ( .A(n13351), .ZN(n11830) );
  OR2_X1 U12659 ( .A1(n12368), .A2(n12230), .ZN(n12229) );
  AOI21_X1 U12660 ( .B1(n15007), .B2(n14067), .A(n15006), .ZN(n15008) );
  NOR2_X1 U12661 ( .A1(n18161), .A2(n12367), .ZN(n12230) );
  OR2_X2 U12662 ( .A1(n11305), .A2(n11304), .ZN(n11356) );
  INV_X1 U12663 ( .A(n15430), .ZN(n15446) );
  AND2_X2 U12664 ( .A1(n15430), .A2(n11155), .ZN(n10171) );
  AND2_X2 U12665 ( .A1(n11229), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11231) );
  NAND2_X1 U12666 ( .A1(n11291), .A2(n11348), .ZN(n11292) );
  NAND2_X1 U12667 ( .A1(n19481), .A2(n12994), .ZN(n12828) );
  INV_X1 U12668 ( .A(n19481), .ZN(n19347) );
  NAND2_X1 U12669 ( .A1(n10272), .A2(n10287), .ZN(n10800) );
  OAI211_X1 U12670 ( .C1(n9742), .C2(n12964), .A(n10315), .B(n10314), .ZN(
        n10347) );
  AND2_X1 U12671 ( .A1(n9750), .A2(n10359), .ZN(n10373) );
  AND2_X1 U12672 ( .A1(n19387), .A2(n13430), .ZN(n19416) );
  OR2_X1 U12673 ( .A1(n9726), .A2(n13430), .ZN(n15539) );
  INV_X1 U12674 ( .A(n10945), .ZN(n10947) );
  AOI22_X1 U12675 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10255) );
  NAND2_X1 U12676 ( .A1(n9748), .A2(n13362), .ZN(n20496) );
  INV_X1 U12677 ( .A(n13613), .ZN(n11836) );
  AND2_X1 U12678 ( .A1(n10836), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10839) );
  AOI21_X1 U12679 ( .B1(n11835), .B2(n11955), .A(n11834), .ZN(n13613) );
  OAI22_X1 U12680 ( .A1(n10557), .A2(n14588), .B1(n14579), .B2(n19764), .ZN(
        n10367) );
  NAND2_X1 U12681 ( .A1(n10212), .A2(n10305), .ZN(n10272) );
  NAND2_X1 U12682 ( .A1(n13278), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13279) );
  AND4_X1 U12683 ( .A1(n10421), .A2(n10420), .A3(n10419), .A4(n10418), .ZN(
        n10422) );
  OR2_X1 U12684 ( .A1(n10374), .A2(n10371), .ZN(n10416) );
  NAND2_X1 U12685 ( .A1(n10374), .A2(n19347), .ZN(n10382) );
  AND3_X1 U12686 ( .A1(n12549), .A2(n18378), .A3(n17794), .ZN(n10148) );
  NOR2_X1 U12687 ( .A1(n17820), .A2(n12443), .ZN(n10149) );
  OR3_X1 U12688 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17887), .ZN(n10150) );
  INV_X1 U12689 ( .A(n12434), .ZN(n17998) );
  OR2_X2 U12690 ( .A1(n12140), .A2(n12144), .ZN(n10152) );
  INV_X1 U12691 ( .A(n10152), .ZN(n12189) );
  NAND2_X1 U12692 ( .A1(n11173), .A2(n11172), .ZN(n19487) );
  INV_X1 U12693 ( .A(n19487), .ZN(n16621) );
  AND2_X1 U12694 ( .A1(n11173), .A2(n20171), .ZN(n16624) );
  OR4_X1 U12695 ( .A1(n15789), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14457), .A4(n14456), .ZN(n10153) );
  OR2_X1 U12696 ( .A1(n11218), .A2(n15589), .ZN(n10154) );
  AND2_X1 U12697 ( .A1(n11185), .A2(n11184), .ZN(n10155) );
  AND2_X2 U12698 ( .A1(n20203), .A2(n12133), .ZN(n20350) );
  NAND2_X1 U12699 ( .A1(n9800), .A2(n11962), .ZN(n14271) );
  OR2_X1 U12700 ( .A1(n17997), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10156) );
  OR2_X1 U12701 ( .A1(n17833), .A2(n17997), .ZN(n10157) );
  INV_X1 U12702 ( .A(n13715), .ZN(n13716) );
  INV_X1 U12703 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12430) );
  OR2_X1 U12704 ( .A1(n15097), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10160) );
  AND3_X1 U12705 ( .A1(n14460), .A2(n10153), .A3(n14459), .ZN(n10161) );
  AND2_X1 U12706 ( .A1(n18444), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n10162) );
  INV_X1 U12707 ( .A(n14270), .ZN(n11962) );
  INV_X1 U12708 ( .A(n12791), .ZN(n11353) );
  AND2_X1 U12709 ( .A1(n12864), .A2(n9739), .ZN(n19475) );
  AND4_X1 U12710 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n10163) );
  OR2_X1 U12711 ( .A1(n15231), .A2(n15230), .ZN(n10164) );
  INV_X1 U12712 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18365) );
  INV_X1 U12713 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20969) );
  OR2_X1 U12714 ( .A1(n16151), .A2(n12451), .ZN(n10165) );
  INV_X1 U12715 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19151) );
  NAND2_X1 U12716 ( .A1(n13115), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10167) );
  NOR2_X1 U12717 ( .A1(n13120), .A2(n13119), .ZN(n10168) );
  INV_X1 U12718 ( .A(n20254), .ZN(n20349) );
  INV_X1 U12719 ( .A(n12316), .ZN(n12156) );
  AND4_X1 U12720 ( .A1(n11290), .A2(n11289), .A3(n11288), .A4(n11287), .ZN(
        n10169) );
  OR2_X1 U12721 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13475) );
  OR2_X1 U12722 ( .A1(n14444), .A2(n10986), .ZN(n10170) );
  INV_X1 U12723 ( .A(n16416), .ZN(n14453) );
  NAND2_X1 U12724 ( .A1(n12811), .A2(n12810), .ZN(n12812) );
  AND4_X1 U12725 ( .A1(n11285), .A2(n11284), .A3(n11283), .A4(n11282), .ZN(
        n10172) );
  BUF_X1 U12726 ( .A(n13172), .Z(n14313) );
  NAND2_X1 U12727 ( .A1(n10278), .A2(n10305), .ZN(n10288) );
  INV_X1 U12728 ( .A(n11648), .ZN(n11620) );
  AND2_X1 U12729 ( .A1(n11649), .A2(n11621), .ZN(n11624) );
  AOI22_X1 U12730 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10190) );
  AND2_X1 U12731 ( .A1(n20549), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11636) );
  OR2_X1 U12732 ( .A1(n11514), .A2(n11513), .ZN(n11538) );
  NAND2_X1 U12733 ( .A1(n20149), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10491) );
  AND2_X1 U12734 ( .A1(n14524), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10437) );
  INV_X1 U12735 ( .A(n15431), .ZN(n11155) );
  NOR2_X1 U12736 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11661), .ZN(
        n12521) );
  INV_X1 U12737 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12894) );
  AND4_X1 U12738 ( .A1(n11238), .A2(n11237), .A3(n11236), .A4(n11235), .ZN(
        n11239) );
  AND2_X1 U12739 ( .A1(n10305), .A2(n13890), .ZN(n10280) );
  OR2_X1 U12740 ( .A1(n10573), .A2(n10572), .ZN(n10577) );
  INV_X1 U12741 ( .A(n10437), .ZN(n11099) );
  INV_X1 U12742 ( .A(n14451), .ZN(n14452) );
  AOI22_X1 U12743 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10181) );
  NOR2_X1 U12744 ( .A1(n12421), .A2(n12407), .ZN(n12399) );
  AND2_X1 U12745 ( .A1(n14826), .A2(n14825), .ZN(n12072) );
  NAND2_X1 U12746 ( .A1(n11682), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12115) );
  INV_X1 U12747 ( .A(n12029), .ZN(n11680) );
  INV_X1 U12748 ( .A(n14254), .ZN(n11899) );
  INV_X1 U12749 ( .A(n14226), .ZN(n11887) );
  NOR2_X1 U12750 ( .A1(n11608), .A2(n16296), .ZN(n15278) );
  AND2_X1 U12751 ( .A1(n12884), .A2(n12883), .ZN(n13028) );
  INV_X1 U12752 ( .A(n11662), .ZN(n11665) );
  NAND2_X1 U12753 ( .A1(n10647), .A2(n13272), .ZN(n10656) );
  AND2_X1 U12754 ( .A1(n10170), .A2(n10987), .ZN(n10991) );
  INV_X1 U12755 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20937) );
  NOR2_X1 U12756 ( .A1(n12146), .A2(n12140), .ZN(n12191) );
  INV_X1 U12757 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12455) );
  NAND2_X1 U12758 ( .A1(n12377), .A2(n12376), .ZN(n12383) );
  INV_X1 U12759 ( .A(n12792), .ZN(n11349) );
  INV_X1 U12760 ( .A(n20696), .ZN(n13496) );
  INV_X1 U12761 ( .A(n13178), .ZN(n13175) );
  INV_X1 U12762 ( .A(n12509), .ZN(n12482) );
  INV_X1 U12763 ( .A(n13185), .ZN(n11795) );
  NOR2_X1 U12764 ( .A1(n13487), .A2(n14711), .ZN(n13488) );
  NAND2_X1 U12765 ( .A1(n11684), .A2(n11683), .ZN(n12484) );
  OR2_X1 U12766 ( .A1(n12074), .A2(n14815), .ZN(n12096) );
  INV_X1 U12767 ( .A(n11882), .ZN(n11910) );
  NAND2_X1 U12768 ( .A1(n15097), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11612) );
  NAND2_X1 U12769 ( .A1(n9856), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11609) );
  NOR2_X1 U12770 ( .A1(n11601), .A2(n11602), .ZN(n15111) );
  OR2_X1 U12771 ( .A1(n11601), .A2(n15313), .ZN(n15121) );
  AND2_X1 U12772 ( .A1(n13054), .A2(n13053), .ZN(n15232) );
  OAI21_X1 U12773 ( .B1(n14191), .B2(n16406), .A(n14161), .ZN(n14190) );
  INV_X1 U12774 ( .A(n14152), .ZN(n20421) );
  INV_X1 U12775 ( .A(n14133), .ZN(n14141) );
  NAND2_X1 U12776 ( .A1(n10541), .A2(n10540), .ZN(n10578) );
  AND2_X1 U12777 ( .A1(n13121), .A2(n10168), .ZN(n13122) );
  NAND2_X1 U12778 ( .A1(n12826), .A2(n19670), .ZN(n12998) );
  AND2_X1 U12779 ( .A1(n14546), .A2(n14545), .ZN(n14547) );
  NAND2_X1 U12780 ( .A1(n15587), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13503) );
  INV_X1 U12781 ( .A(n15516), .ZN(n10922) );
  AND2_X1 U12782 ( .A1(n10652), .A2(n16580), .ZN(n15967) );
  OAI21_X1 U12783 ( .B1(n10990), .B2(n11140), .A(n10989), .ZN(n13411) );
  INV_X1 U12784 ( .A(n19492), .ZN(n16008) );
  INV_X1 U12785 ( .A(n18501), .ZN(n16052) );
  INV_X1 U12786 ( .A(n17609), .ZN(n17575) );
  INV_X2 U12787 ( .A(n10152), .ZN(n17455) );
  NAND2_X1 U12788 ( .A1(n12433), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12434) );
  NOR2_X1 U12789 ( .A1(n18163), .A2(n18119), .ZN(n17944) );
  NAND2_X1 U12790 ( .A1(n18351), .A2(n12455), .ZN(n12456) );
  INV_X1 U12791 ( .A(n17913), .ZN(n17886) );
  NAND2_X1 U12792 ( .A1(n12353), .A2(n12364), .ZN(n12338) );
  OR2_X1 U12793 ( .A1(n14414), .A2(n20614), .ZN(n13497) );
  NAND2_X1 U12794 ( .A1(n13486), .A2(n13485), .ZN(n16272) );
  INV_X1 U12795 ( .A(n14294), .ZN(n14236) );
  OAI21_X1 U12796 ( .B1(n13475), .B2(n14731), .A(n11764), .ZN(n12131) );
  NAND2_X1 U12797 ( .A1(n12026), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12029) );
  NAND2_X1 U12798 ( .A1(n14824), .A2(n14921), .ZN(n14923) );
  AND2_X1 U12799 ( .A1(n11926), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11930) );
  AOI21_X1 U12800 ( .B1(n11813), .B2(n11955), .A(n11812), .ZN(n13347) );
  NOR2_X1 U12801 ( .A1(n15001), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14382) );
  OR2_X1 U12802 ( .A1(n15293), .A2(n15232), .ZN(n14387) );
  INV_X1 U12803 ( .A(n14387), .ZN(n15304) );
  AND2_X1 U12804 ( .A1(n11673), .A2(n11672), .ZN(n16187) );
  INV_X1 U12805 ( .A(n14148), .ZN(n14193) );
  OR2_X1 U12806 ( .A1(n20496), .A2(n14149), .ZN(n13920) );
  OR2_X1 U12807 ( .A1(n20496), .A2(n13639), .ZN(n13951) );
  OAI21_X1 U12808 ( .B1(n14046), .B2(n16406), .A(n12624), .ZN(n14045) );
  OR2_X1 U12809 ( .A1(n11797), .A2(n9748), .ZN(n20525) );
  INV_X1 U12810 ( .A(n13239), .ZN(n13746) );
  AOI21_X1 U12811 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20549), .A(n13746), 
        .ZN(n20557) );
  NAND2_X1 U12812 ( .A1(n11494), .A2(n11493), .ZN(n13361) );
  AND2_X1 U12813 ( .A1(n15938), .A2(n13712), .ZN(n11144) );
  OR2_X1 U12814 ( .A1(n20188), .A2(n13514), .ZN(n19305) );
  INV_X1 U12815 ( .A(n19357), .ZN(n15581) );
  INV_X1 U12816 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13603) );
  OR3_X1 U12817 ( .A1(n19248), .A2(n11020), .A3(n16571), .ZN(n15754) );
  INV_X1 U12818 ( .A(n10542), .ZN(n11010) );
  NAND2_X1 U12819 ( .A1(n10767), .A2(n10765), .ZN(n12859) );
  CLKBUF_X1 U12820 ( .A(n10799), .Z(n16656) );
  INV_X1 U12821 ( .A(n19533), .ZN(n19525) );
  AOI22_X1 U12822 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n18934), .B2(n19103), .ZN(
        n12421) );
  NOR2_X1 U12823 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17062), .ZN(n17061) );
  NOR2_X1 U12824 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17110), .ZN(n17079) );
  INV_X1 U12825 ( .A(n17178), .ZN(n17173) );
  NOR3_X1 U12826 ( .A1(n16057), .A2(n17319), .A3(n17318), .ZN(n17290) );
  NOR2_X1 U12827 ( .A1(n17674), .A2(n17525), .ZN(n17526) );
  NOR2_X1 U12828 ( .A1(n18191), .A2(n17846), .ZN(n17845) );
  NAND2_X1 U12829 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18051), .ZN(n18016) );
  NOR2_X1 U12830 ( .A1(n12246), .A2(n12250), .ZN(n12252) );
  AOI21_X1 U12831 ( .B1(n12587), .B2(n18438), .A(n12586), .ZN(n12588) );
  AND2_X1 U12832 ( .A1(n12580), .A2(n12456), .ZN(n12457) );
  NAND2_X1 U12833 ( .A1(n12439), .A2(n10150), .ZN(n12440) );
  INV_X2 U12834 ( .A(n18928), .ZN(n18916) );
  INV_X1 U12835 ( .A(n12390), .ZN(n12388) );
  AOI211_X1 U12836 ( .C1(n12427), .C2(n18957), .A(n16136), .B(n12426), .ZN(
        n12428) );
  INV_X1 U12837 ( .A(n18963), .ZN(n18943) );
  INV_X1 U12838 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18934) );
  INV_X1 U12839 ( .A(n12340), .ZN(n18491) );
  AND2_X1 U12840 ( .A1(n16239), .A2(n14813), .ZN(n16219) );
  NOR2_X2 U12841 ( .A1(n14892), .A2(n13497), .ZN(n20233) );
  AND2_X1 U12842 ( .A1(n13486), .A2(n13480), .ZN(n20253) );
  INV_X1 U12843 ( .A(n16289), .ZN(n14985) );
  INV_X1 U12844 ( .A(n13200), .ZN(n20323) );
  INV_X2 U12845 ( .A(n13181), .ZN(n20345) );
  AND2_X1 U12846 ( .A1(n13181), .A2(n13292), .ZN(n20346) );
  AOI21_X1 U12847 ( .B1(n14917), .B2(n14916), .A(n14915), .ZN(n16286) );
  INV_X1 U12848 ( .A(n14923), .ZN(n14841) );
  AND2_X1 U12849 ( .A1(n14285), .A2(n14286), .ZN(n14287) );
  NAND2_X1 U12850 ( .A1(n11883), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11882) );
  NAND2_X1 U12851 ( .A1(n11831), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11848) );
  AND2_X1 U12852 ( .A1(n13074), .A2(n11793), .ZN(n13080) );
  AND2_X1 U12853 ( .A1(n15269), .A2(n14406), .ZN(n15220) );
  AND2_X1 U12854 ( .A1(n14055), .A2(n13735), .ZN(n16370) );
  NOR2_X1 U12855 ( .A1(n15304), .A2(n15324), .ZN(n20382) );
  NOR2_X1 U12856 ( .A1(n16406), .A2(n16187), .ZN(n12930) );
  OAI22_X1 U12857 ( .A1(n13831), .A2(n13834), .B1(n13828), .B2(n20450), .ZN(
        n20416) );
  NAND2_X1 U12858 ( .A1(n13626), .A2(n11797), .ZN(n20424) );
  NOR2_X1 U12859 ( .A1(n20424), .A2(n13639), .ZN(n14148) );
  INV_X1 U12860 ( .A(n20456), .ZN(n20488) );
  INV_X1 U12861 ( .A(n13920), .ZN(n20515) );
  AND2_X1 U12862 ( .A1(n20493), .A2(n15333), .ZN(n13922) );
  INV_X1 U12863 ( .A(n13951), .ZN(n13583) );
  INV_X1 U12864 ( .A(n13668), .ZN(n13783) );
  NOR2_X1 U12865 ( .A1(n12607), .A2(n13659), .ZN(n13740) );
  INV_X1 U12866 ( .A(n20525), .ZN(n13660) );
  OAI211_X1 U12867 ( .C1(n13750), .C2(n13749), .A(n20454), .B(n13748), .ZN(
        n13774) );
  INV_X1 U12868 ( .A(n13741), .ZN(n13773) );
  NOR2_X1 U12869 ( .A1(n13312), .A2(n13746), .ZN(n20579) );
  NOR2_X1 U12870 ( .A1(n13615), .A2(n13746), .ZN(n20604) );
  INV_X1 U12871 ( .A(n13830), .ZN(n20414) );
  INV_X1 U12872 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20614) );
  OR2_X1 U12873 ( .A1(n20059), .A2(n20182), .ZN(n12667) );
  NAND2_X1 U12874 ( .A1(n13518), .A2(n13517), .ZN(n19342) );
  INV_X1 U12875 ( .A(n19308), .ZN(n19341) );
  INV_X1 U12876 ( .A(n19306), .ZN(n19351) );
  OR2_X1 U12877 ( .A1(n11112), .A2(n11111), .ZN(n13465) );
  OR2_X1 U12878 ( .A1(n11034), .A2(n11033), .ZN(n13115) );
  INV_X1 U12879 ( .A(n15539), .ZN(n15527) );
  AND2_X1 U12880 ( .A1(n13717), .A2(n13715), .ZN(n19357) );
  INV_X1 U12881 ( .A(n19390), .ZN(n19417) );
  INV_X1 U12882 ( .A(n10755), .ZN(n12725) );
  INV_X1 U12883 ( .A(n12727), .ZN(n16411) );
  NAND2_X1 U12884 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n13505), .ZN(
        n13504) );
  AND2_X1 U12885 ( .A1(n16541), .A2(n19472), .ZN(n16530) );
  XNOR2_X1 U12886 ( .A(n10738), .B(n10740), .ZN(n15607) );
  AND2_X1 U12887 ( .A1(n16581), .A2(n11180), .ZN(n15892) );
  INV_X1 U12888 ( .A(n19491), .ZN(n16635) );
  AND2_X1 U12889 ( .A1(n11173), .A2(n16658), .ZN(n15924) );
  AND2_X1 U12890 ( .A1(n11173), .A2(n20170), .ZN(n16639) );
  AND2_X1 U12891 ( .A1(n12863), .A2(n19151), .ZN(n19999) );
  OAI21_X1 U12892 ( .B1(n19507), .B2(n19537), .A(n19999), .ZN(n19540) );
  NAND2_X1 U12893 ( .A1(n19549), .A2(n20161), .ZN(n19700) );
  NOR2_X1 U12894 ( .A1(n19820), .A2(n19757), .ZN(n19574) );
  OAI21_X1 U12895 ( .B1(n19641), .B2(n19670), .A(n19640), .ZN(n19665) );
  NAND2_X1 U12896 ( .A1(n20145), .A2(n19573), .ZN(n20132) );
  AOI22_X1 U12897 ( .A1(n19798), .A2(n19797), .B1(n19796), .B2(n20182), .ZN(
        n19814) );
  INV_X1 U12898 ( .A(n19847), .ZN(n19838) );
  OAI21_X1 U12899 ( .B1(n19856), .B2(n19871), .A(n19999), .ZN(n19873) );
  NOR2_X2 U12900 ( .A1(n19851), .A2(n20132), .ZN(n19904) );
  NOR2_X1 U12901 ( .A1(n19877), .A2(n20132), .ZN(n19912) );
  INV_X1 U12902 ( .A(n20004), .ZN(n19967) );
  AND2_X1 U12903 ( .A1(n19514), .A2(n19525), .ZN(n20005) );
  INV_X1 U12904 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16011) );
  INV_X1 U12905 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20061) );
  NOR2_X1 U12906 ( .A1(n19060), .A2(n16833), .ZN(n16877) );
  INV_X1 U12907 ( .A(n17196), .ZN(n17165) );
  NOR2_X1 U12908 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17006), .ZN(n16987) );
  NOR2_X1 U12909 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17030), .ZN(n17016) );
  NOR2_X1 U12910 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17052), .ZN(n17034) );
  NOR2_X1 U12911 ( .A1(n18977), .A2(n12648), .ZN(n17178) );
  NOR2_X1 U12912 ( .A1(n17292), .A2(n17291), .ZN(n17265) );
  INV_X1 U12913 ( .A(n17375), .ZN(n17363) );
  NAND2_X1 U12914 ( .A1(n17523), .A2(n17379), .ZN(n17498) );
  NOR2_X1 U12915 ( .A1(n16055), .A2(n16138), .ZN(n16212) );
  INV_X1 U12916 ( .A(n17544), .ZN(n17539) );
  NOR2_X1 U12917 ( .A1(n17736), .A2(n17596), .ZN(n17591) );
  NAND2_X1 U12918 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17610), .ZN(n17609) );
  NOR2_X1 U12919 ( .A1(n17774), .A2(n17639), .ZN(n17634) );
  AND2_X1 U12920 ( .A1(n18929), .A2(n17524), .ZN(n17671) );
  NAND2_X1 U12921 ( .A1(n19128), .A2(n18959), .ZN(n17727) );
  INV_X1 U12922 ( .A(n17781), .ZN(n17786) );
  NAND2_X1 U12923 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18035), .ZN(
        n18338) );
  INV_X1 U12924 ( .A(n17799), .ZN(n12466) );
  NOR2_X1 U12925 ( .A1(n17947), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17946) );
  INV_X1 U12926 ( .A(n18358), .ZN(n18378) );
  NAND2_X1 U12927 ( .A1(n18101), .A2(n12382), .ZN(n18091) );
  NOR2_X2 U12928 ( .A1(n12428), .A2(n18983), .ZN(n18438) );
  INV_X1 U12929 ( .A(n18438), .ZN(n18461) );
  INV_X1 U12930 ( .A(U212), .ZN(n16770) );
  OR2_X1 U12931 ( .A1(n13037), .A2(n12515), .ZN(n13149) );
  INV_X1 U12932 ( .A(n20253), .ZN(n20267) );
  INV_X1 U12933 ( .A(n20233), .ZN(n20242) );
  INV_X1 U12934 ( .A(n16233), .ZN(n14981) );
  OAI21_X2 U12935 ( .B1(n13149), .B2(n12529), .A(n12528), .ZN(n14290) );
  NAND2_X1 U12936 ( .A1(n20321), .A2(n20698), .ZN(n20310) );
  OR2_X1 U12937 ( .A1(n13037), .A2(n12967), .ZN(n20321) );
  NOR2_X1 U12938 ( .A1(n13149), .A2(n13148), .ZN(n13181) );
  OAI21_X1 U12939 ( .B1(n14841), .B2(n14840), .A(n14916), .ZN(n15088) );
  OAI21_X1 U12940 ( .B1(n14287), .B2(n14257), .A(n14256), .ZN(n15129) );
  INV_X1 U12941 ( .A(n14067), .ZN(n15147) );
  AND2_X1 U12942 ( .A1(n14392), .A2(n14390), .ZN(n16348) );
  INV_X1 U12943 ( .A(n16379), .ZN(n20385) );
  INV_X1 U12944 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16166) );
  OR2_X1 U12945 ( .A1(n20424), .A2(n20448), .ZN(n20447) );
  AOI22_X1 U12946 ( .A1(n14160), .A2(n14156), .B1(n14154), .B2(n14153), .ZN(
        n14197) );
  NAND2_X1 U12947 ( .A1(n13628), .A2(n13627), .ZN(n20456) );
  OR2_X1 U12948 ( .A1(n20496), .A2(n20448), .ZN(n20519) );
  AOI22_X1 U12949 ( .A1(n13925), .A2(n13922), .B1(n14103), .B2(n14153), .ZN(
        n13954) );
  OR2_X1 U12950 ( .A1(n20496), .A2(n13369), .ZN(n13668) );
  NAND2_X1 U12951 ( .A1(n13660), .A2(n13740), .ZN(n20548) );
  AOI22_X1 U12952 ( .A1(n12623), .A2(n12618), .B1(n14154), .B2(n14104), .ZN(
        n14051) );
  NAND2_X1 U12953 ( .A1(n13660), .A2(n12608), .ZN(n14048) );
  INV_X1 U12954 ( .A(n20567), .ZN(n14173) );
  INV_X1 U12955 ( .A(n20597), .ZN(n14165) );
  OR2_X1 U12956 ( .A1(n14099), .A2(n20448), .ZN(n20612) );
  OR2_X1 U12957 ( .A1(n14099), .A2(n14149), .ZN(n20562) );
  OR2_X1 U12958 ( .A1(n14099), .A2(n13639), .ZN(n14106) );
  OR2_X1 U12959 ( .A1(n16657), .A2(n12656), .ZN(n12670) );
  NAND2_X1 U12960 ( .A1(n16411), .A2(n16684), .ZN(n19323) );
  AND2_X1 U12961 ( .A1(n12836), .A2(n16682), .ZN(n15537) );
  AND2_X1 U12962 ( .A1(n19360), .A2(n19390), .ZN(n19385) );
  NAND2_X1 U12963 ( .A1(n19387), .A2(n13429), .ZN(n19390) );
  INV_X1 U12964 ( .A(n19376), .ZN(n19422) );
  OR2_X1 U12965 ( .A1(n19458), .A2(n19454), .ZN(n19424) );
  INV_X1 U12966 ( .A(n19458), .ZN(n19456) );
  INV_X1 U12967 ( .A(n12717), .ZN(n12727) );
  INV_X1 U12968 ( .A(n19475), .ZN(n19464) );
  INV_X1 U12969 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16520) );
  INV_X1 U12970 ( .A(n16530), .ZN(n19471) );
  INV_X1 U12971 ( .A(n11220), .ZN(n11221) );
  INV_X1 U12972 ( .A(n16624), .ZN(n19490) );
  OR2_X1 U12973 ( .A1(n19820), .A2(n19700), .ZN(n19569) );
  INV_X1 U12974 ( .A(n19574), .ZN(n19598) );
  OR2_X1 U12975 ( .A1(n19757), .A2(n20132), .ZN(n19668) );
  INV_X1 U12976 ( .A(n19783), .ZN(n19756) );
  OR2_X1 U12977 ( .A1(n19758), .A2(n19757), .ZN(n19818) );
  NAND2_X1 U12978 ( .A1(n19788), .A2(n19787), .ZN(n19847) );
  INV_X1 U12979 ( .A(n19853), .ZN(n19876) );
  INV_X1 U12980 ( .A(n19912), .ZN(n19945) );
  AND2_X1 U12981 ( .A1(n13255), .A2(n13254), .ZN(n19966) );
  INV_X1 U12982 ( .A(n19976), .ZN(n20028) );
  NAND2_X1 U12983 ( .A1(n12344), .A2(n12346), .ZN(n19145) );
  INV_X1 U12984 ( .A(n17197), .ZN(n17163) );
  NOR2_X1 U12985 ( .A1(n16885), .A2(n17239), .ZN(n17243) );
  NOR2_X1 U12986 ( .A1(n16892), .A2(n17249), .ZN(n17253) );
  AND2_X1 U12987 ( .A1(n17523), .A2(n17647), .ZN(n17520) );
  INV_X1 U12988 ( .A(n17607), .ZN(n17582) );
  NOR2_X1 U12989 ( .A1(n12228), .A2(n12227), .ZN(n17648) );
  NOR2_X1 U12990 ( .A1(n12208), .A2(n12207), .ZN(n17661) );
  INV_X1 U12991 ( .A(n17692), .ZN(n17696) );
  INV_X1 U12992 ( .A(n17712), .ZN(n17724) );
  AOI221_X1 U12993 ( .B1(n19004), .B2(n18976), .C1(n17728), .C2(n18976), .A(
        n17727), .ZN(n17755) );
  INV_X1 U12994 ( .A(n17779), .ZN(n17788) );
  INV_X1 U12995 ( .A(n12570), .ZN(n12571) );
  OR2_X1 U12996 ( .A1(n17967), .A2(n18233), .ZN(n17929) );
  INV_X1 U12997 ( .A(n18060), .ZN(n18040) );
  OAI21_X2 U12998 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19127), .A(n16819), 
        .ZN(n18162) );
  NOR2_X1 U12999 ( .A1(n10148), .A2(n12466), .ZN(n12467) );
  NAND2_X1 U13000 ( .A1(n12557), .A2(n18458), .ZN(n18358) );
  OAI21_X1 U13001 ( .B1(n18300), .B2(n18264), .A(n18438), .ZN(n18366) );
  INV_X1 U13002 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18932) );
  OR3_X1 U13003 ( .A1(n18989), .A2(n18988), .A3(n18987), .ZN(n18990) );
  INV_X1 U13004 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19079) );
  INV_X1 U13005 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19012) );
  AND2_X1 U13006 ( .A1(n12541), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14279)
         );
  INV_X1 U13007 ( .A(n16775), .ZN(n16772) );
  OAI211_X1 U13008 ( .C1(n15594), .C2(n19500), .A(n11222), .B(n11221), .ZN(
        P2_U3016) );
  AOI22_X1 U13009 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9735), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10174) );
  AND3_X4 U13010 ( .A1(n16647), .A2(n10077), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14685) );
  AOI22_X1 U13011 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10173) );
  AND2_X4 U13012 ( .A1(n16017), .A2(n16647), .ZN(n14686) );
  AOI22_X1 U13013 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10175) );
  NAND2_X1 U13014 ( .A1(n10178), .A2(n10177), .ZN(n10185) );
  AOI22_X1 U13015 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10240), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10179) );
  AND2_X1 U13016 ( .A1(n10179), .A2(n16039), .ZN(n10183) );
  AOI22_X1 U13017 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13018 ( .A1(n14684), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10180) );
  NAND4_X1 U13019 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n10184) );
  AOI22_X1 U13020 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10240), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10186) );
  AND2_X1 U13021 ( .A1(n10186), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10192) );
  AOI22_X1 U13022 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13023 ( .A1(n14684), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10189) );
  NAND4_X1 U13024 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10199) );
  AOI22_X1 U13025 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10240), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10194) );
  AOI22_X1 U13026 ( .A1(n14684), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10193) );
  AND3_X1 U13027 ( .A1(n10194), .A2(n16039), .A3(n10193), .ZN(n10197) );
  AOI22_X1 U13028 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13029 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10195) );
  NAND3_X1 U13030 ( .A1(n10197), .A2(n10196), .A3(n10195), .ZN(n10198) );
  AOI22_X1 U13031 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10203) );
  AOI22_X1 U13032 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13033 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10201) );
  NAND4_X1 U13034 ( .A1(n10203), .A2(n10202), .A3(n10201), .A4(n10200), .ZN(
        n10204) );
  NAND2_X1 U13035 ( .A1(n10204), .A2(n16039), .ZN(n10211) );
  AOI22_X1 U13036 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13037 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13038 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10205) );
  NAND4_X1 U13039 ( .A1(n10208), .A2(n10207), .A3(n10206), .A4(n10205), .ZN(
        n10209) );
  NAND2_X1 U13040 ( .A1(n10209), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10210) );
  AOI22_X1 U13041 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U13042 ( .A1(n14684), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13043 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10240), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10214) );
  NAND4_X1 U13044 ( .A1(n10216), .A2(n10215), .A3(n10214), .A4(n10213), .ZN(
        n10217) );
  NAND2_X1 U13045 ( .A1(n10217), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10224) );
  AOI22_X1 U13046 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10221) );
  AOI22_X1 U13047 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10240), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10220) );
  AOI22_X1 U13048 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14686), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10218) );
  NAND4_X1 U13049 ( .A1(n10221), .A2(n10220), .A3(n10219), .A4(n10218), .ZN(
        n10222) );
  NAND2_X1 U13050 ( .A1(n10222), .A2(n16039), .ZN(n10223) );
  NAND2_X2 U13051 ( .A1(n10224), .A2(n10223), .ZN(n10973) );
  NAND2_X1 U13052 ( .A1(n10804), .A2(n10225), .ZN(n10943) );
  AOI22_X1 U13053 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13054 ( .A1(n14684), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U13055 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10240), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10227) );
  NAND4_X1 U13056 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10230) );
  NAND2_X1 U13057 ( .A1(n10230), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10237) );
  AOI22_X1 U13058 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U13059 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10240), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10232) );
  AOI22_X1 U13060 ( .A1(n14684), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10231) );
  NAND4_X1 U13061 ( .A1(n10234), .A2(n10233), .A3(n10232), .A4(n10231), .ZN(
        n10235) );
  NAND2_X1 U13062 ( .A1(n10235), .A2(n16039), .ZN(n10236) );
  NAND2_X1 U13063 ( .A1(n10943), .A2(n13890), .ZN(n10239) );
  INV_X2 U13064 ( .A(n10305), .ZN(n13008) );
  NAND2_X1 U13065 ( .A1(n10285), .A2(n10268), .ZN(n10238) );
  NAND2_X1 U13066 ( .A1(n10239), .A2(n10238), .ZN(n10310) );
  AOI22_X1 U13067 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13068 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10243) );
  AOI22_X1 U13069 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10242) );
  AOI22_X1 U13070 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14534), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13071 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13072 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13073 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13074 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13075 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13076 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U13077 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10256) );
  AOI22_X1 U13078 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13079 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U13080 ( .A1(n10310), .A2(n10043), .ZN(n10274) );
  MUX2_X1 U13081 ( .A(n13008), .B(n10973), .S(n10287), .Z(n10266) );
  AOI22_X1 U13082 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13083 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13084 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U13085 ( .A1(n10188), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10257) );
  AOI22_X1 U13086 ( .A1(n10187), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9736), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10264) );
  AOI22_X1 U13087 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10263) );
  AOI22_X1 U13088 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U13089 ( .A1(n10272), .A2(n13890), .ZN(n10289) );
  NAND3_X1 U13090 ( .A1(n10266), .A2(n10265), .A3(n10289), .ZN(n10271) );
  NAND4_X1 U13091 ( .A1(n10268), .A2(n10267), .A3(n10766), .A4(n10973), .ZN(
        n10269) );
  NOR2_X2 U13092 ( .A1(n10269), .A2(n10276), .ZN(n10296) );
  INV_X1 U13093 ( .A(n10296), .ZN(n10270) );
  NAND3_X1 U13094 ( .A1(n10271), .A2(n20179), .A3(n10270), .ZN(n10950) );
  NAND3_X1 U13095 ( .A1(n10285), .A2(n9739), .A3(n10272), .ZN(n10311) );
  NAND2_X1 U13096 ( .A1(n10311), .A2(n20179), .ZN(n10273) );
  NAND2_X1 U13097 ( .A1(n10274), .A2(n10312), .ZN(n10275) );
  NAND2_X1 U13098 ( .A1(n10275), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10283) );
  INV_X1 U13099 ( .A(n10276), .ZN(n10277) );
  NAND4_X1 U13100 ( .A1(n13890), .A2(n10277), .A3(n10279), .A4(n10973), .ZN(
        n10814) );
  NAND3_X1 U13101 ( .A1(n10814), .A2(n10941), .A3(n19514), .ZN(n10282) );
  INV_X1 U13102 ( .A(n10794), .ZN(n10281) );
  NAND2_X1 U13103 ( .A1(n19503), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10755) );
  NAND2_X2 U13104 ( .A1(n10283), .A2(n10306), .ZN(n10344) );
  NAND2_X1 U13105 ( .A1(n10043), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10284) );
  AND2_X2 U13106 ( .A1(n10268), .A2(n10941), .ZN(n10298) );
  INV_X1 U13107 ( .A(n10298), .ZN(n10954) );
  NOR2_X1 U13108 ( .A1(n10284), .A2(n10954), .ZN(n10286) );
  OAI22_X1 U13109 ( .A1(n10344), .A2(n10286), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n10339), .ZN(n10295) );
  NAND2_X1 U13110 ( .A1(n10297), .A2(n10502), .ZN(n12660) );
  NAND3_X1 U13111 ( .A1(n12660), .A2(n10973), .A3(n10287), .ZN(n10292) );
  NAND2_X1 U13112 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  NOR2_X2 U13113 ( .A1(n10292), .A2(n10291), .ZN(n10940) );
  NAND2_X1 U13114 ( .A1(n10940), .A2(n10298), .ZN(n10303) );
  NAND2_X1 U13115 ( .A1(n19151), .A2(n16011), .ZN(n20187) );
  NOR2_X1 U13116 ( .A1(n20187), .A2(n20166), .ZN(n10293) );
  AOI21_X1 U13117 ( .B1(n16019), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10293), 
        .ZN(n10294) );
  NAND2_X1 U13118 ( .A1(n10295), .A2(n10294), .ZN(n10348) );
  NAND2_X1 U13119 ( .A1(n10296), .A2(n20179), .ZN(n10799) );
  NAND2_X1 U13120 ( .A1(n10799), .A2(n16686), .ZN(n11169) );
  INV_X1 U13121 ( .A(n10297), .ZN(n10299) );
  NAND2_X1 U13122 ( .A1(n10300), .A2(n13008), .ZN(n10301) );
  NOR2_X1 U13123 ( .A1(n10945), .A2(n10301), .ZN(n10302) );
  OR2_X2 U13124 ( .A1(n11169), .A2(n10302), .ZN(n10320) );
  NAND2_X1 U13125 ( .A1(n10320), .A2(n9739), .ZN(n10304) );
  INV_X1 U13126 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12964) );
  INV_X1 U13127 ( .A(n16686), .ZN(n12655) );
  INV_X1 U13128 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n10985) );
  OAI21_X1 U13129 ( .B1(n10854), .B2(n10985), .A(n10306), .ZN(n10309) );
  INV_X1 U13130 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U13131 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10307) );
  OAI211_X1 U13132 ( .C1(n10855), .C2(n12840), .A(n20187), .B(n10307), .ZN(
        n10308) );
  NOR2_X1 U13133 ( .A1(n10309), .A2(n10308), .ZN(n10315) );
  NAND2_X1 U13134 ( .A1(n10310), .A2(n10311), .ZN(n10955) );
  NAND2_X1 U13135 ( .A1(n10955), .A2(n10312), .ZN(n10313) );
  NAND2_X1 U13136 ( .A1(n10313), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U13137 ( .A1(n10348), .A2(n10347), .ZN(n10346) );
  NAND2_X1 U13138 ( .A1(n9751), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10319) );
  AOI22_X1 U13139 ( .A1(n9725), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10317) );
  NAND2_X1 U13140 ( .A1(n11205), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10316) );
  NAND2_X1 U13141 ( .A1(n10319), .A2(n10318), .ZN(n10324) );
  NAND2_X1 U13142 ( .A1(n10344), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10323) );
  NOR2_X1 U13143 ( .A1(n20187), .A2(n20159), .ZN(n10321) );
  AOI21_X1 U13144 ( .B1(n10320), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10321), 
        .ZN(n10322) );
  NAND2_X1 U13145 ( .A1(n10324), .A2(n10325), .ZN(n10354) );
  NAND2_X1 U13146 ( .A1(n10346), .A2(n10354), .ZN(n10328) );
  INV_X1 U13147 ( .A(n10324), .ZN(n10327) );
  INV_X1 U13148 ( .A(n10325), .ZN(n10326) );
  NAND2_X1 U13149 ( .A1(n10328), .A2(n10353), .ZN(n10351) );
  INV_X1 U13150 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13151 ( .A1(n9725), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10331) );
  NAND2_X1 U13152 ( .A1(n11205), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10330) );
  OAI21_X1 U13153 ( .B1(n20149), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16011), 
        .ZN(n10333) );
  AOI21_X1 U13154 ( .B1(n10344), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10333), .ZN(n10334) );
  XNOR2_X2 U13155 ( .A(n10335), .B(n10334), .ZN(n10350) );
  NAND2_X1 U13156 ( .A1(n10351), .A2(n10350), .ZN(n10338) );
  INV_X1 U13157 ( .A(n10334), .ZN(n10336) );
  AOI22_X1 U13158 ( .A1(n10339), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10341) );
  NAND2_X1 U13159 ( .A1(n11205), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10340) );
  NOR2_X1 U13160 ( .A1(n20187), .A2(n20142), .ZN(n10345) );
  OR2_X1 U13161 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  OR2_X2 U13162 ( .A1(n10386), .A2(n10013), .ZN(n10380) );
  INV_X1 U13163 ( .A(n10352), .ZN(n10355) );
  NOR2_X2 U13164 ( .A1(n10380), .A2(n19492), .ZN(n19702) );
  NAND2_X1 U13165 ( .A1(n10388), .A2(n9750), .ZN(n10356) );
  AOI22_X1 U13166 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19702), .B1(
        n19910), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10392) );
  INV_X1 U13167 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14589) );
  NAND2_X1 U13168 ( .A1(n19481), .A2(n10362), .ZN(n10358) );
  OR2_X1 U13169 ( .A1(n9750), .A2(n10358), .ZN(n10370) );
  INV_X1 U13170 ( .A(n10370), .ZN(n10357) );
  NAND2_X1 U13171 ( .A1(n10357), .A2(n10374), .ZN(n10554) );
  INV_X1 U13172 ( .A(n10358), .ZN(n10359) );
  INV_X1 U13173 ( .A(n10373), .ZN(n10360) );
  INV_X1 U13174 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10361) );
  OAI22_X1 U13175 ( .A1(n14589), .A2(n10554), .B1(n10555), .B2(n10361), .ZN(
        n10368) );
  INV_X1 U13176 ( .A(n10362), .ZN(n10363) );
  NAND2_X1 U13177 ( .A1(n9750), .A2(n10364), .ZN(n10366) );
  INV_X1 U13178 ( .A(n10366), .ZN(n10365) );
  INV_X1 U13179 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14588) );
  INV_X1 U13180 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14579) );
  NOR2_X1 U13181 ( .A1(n10368), .A2(n10367), .ZN(n10379) );
  INV_X1 U13182 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11069) );
  INV_X1 U13183 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14580) );
  OAI22_X1 U13184 ( .A1(n11069), .A2(n10416), .B1(n10543), .B2(n14580), .ZN(
        n10377) );
  INV_X1 U13185 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11068) );
  INV_X1 U13186 ( .A(n10371), .ZN(n10372) );
  NAND2_X1 U13187 ( .A1(n10372), .A2(n10374), .ZN(n10405) );
  NAND2_X1 U13188 ( .A1(n10374), .A2(n10373), .ZN(n13252) );
  INV_X1 U13189 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10375) );
  OAI22_X1 U13190 ( .A1(n11068), .A2(n10405), .B1(n13252), .B2(n10375), .ZN(
        n10376) );
  NOR2_X1 U13191 ( .A1(n10377), .A2(n10376), .ZN(n10378) );
  NOR2_X2 U13192 ( .A1(n10380), .A2(n16008), .ZN(n10560) );
  NAND2_X1 U13193 ( .A1(n12831), .A2(n9750), .ZN(n10381) );
  NOR2_X2 U13194 ( .A1(n10382), .A2(n10381), .ZN(n13886) );
  AOI22_X1 U13195 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10560), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10391) );
  NOR2_X2 U13196 ( .A1(n10386), .A2(n10383), .ZN(n10546) );
  AOI22_X1 U13197 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10546), .B1(
        n10547), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10390) );
  INV_X1 U13198 ( .A(n10387), .ZN(n10385) );
  AOI22_X1 U13199 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10548), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10389) );
  NAND4_X1 U13200 ( .A1(n10392), .A2(n9802), .A3(n10391), .A4(n9760), .ZN(
        n10404) );
  AOI22_X1 U13201 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10437), .B1(
        n10438), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10396) );
  AOI22_X1 U13202 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10395) );
  AND2_X2 U13203 ( .A1(n16033), .A2(n16039), .ZN(n10432) );
  AOI22_X1 U13204 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10563), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13205 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10477), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10393) );
  NAND4_X1 U13206 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10402) );
  AND2_X1 U13207 ( .A1(n14684), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10426) );
  AOI22_X1 U13208 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10455), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10400) );
  AND2_X2 U13209 ( .A1(n10240), .A2(n16039), .ZN(n13847) );
  AND2_X1 U13210 ( .A1(n14684), .A2(n16039), .ZN(n10444) );
  AOI22_X1 U13211 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n13847), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10399) );
  AND2_X1 U13212 ( .A1(n14686), .A2(n16039), .ZN(n10472) );
  AND2_X1 U13213 ( .A1(n14685), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13848) );
  AOI22_X1 U13214 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10472), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10398) );
  AOI22_X1 U13215 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n14508), .ZN(n10397) );
  NAND4_X1 U13216 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10401) );
  INV_X1 U13217 ( .A(n10498), .ZN(n11006) );
  NAND2_X1 U13218 ( .A1(n11006), .A2(n9739), .ZN(n10403) );
  INV_X1 U13219 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10408) );
  INV_X1 U13220 ( .A(n10405), .ZN(n19880) );
  INV_X1 U13221 ( .A(n10554), .ZN(n19824) );
  NAND2_X1 U13222 ( .A1(n19824), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10406) );
  OAI211_X1 U13223 ( .C1(n19570), .C2(n10408), .A(n10407), .B(n10406), .ZN(
        n10409) );
  AOI22_X1 U13224 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10560), .B1(
        n19910), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10424) );
  NAND2_X1 U13225 ( .A1(n10549), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10411) );
  NAND2_X1 U13226 ( .A1(n10546), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10410) );
  NOR2_X1 U13227 ( .A1(n10413), .A2(n10412), .ZN(n10423) );
  INV_X1 U13228 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10414) );
  INV_X1 U13229 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14519) );
  OAI22_X1 U13230 ( .A1(n10414), .A2(n10555), .B1(n19764), .B2(n14519), .ZN(
        n10415) );
  INV_X1 U13231 ( .A(n10415), .ZN(n10421) );
  INV_X1 U13232 ( .A(n10416), .ZN(n19605) );
  INV_X1 U13233 ( .A(n10557), .ZN(n19990) );
  AOI22_X1 U13234 ( .A1(n19605), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n19990), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10420) );
  INV_X1 U13235 ( .A(n10543), .ZN(n19543) );
  INV_X1 U13236 ( .A(n13252), .ZN(n10417) );
  AOI22_X1 U13237 ( .A1(n19543), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10417), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10419) );
  NAND2_X1 U13238 ( .A1(n10547), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10418) );
  NAND4_X1 U13239 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        n10463) );
  AOI22_X1 U13240 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10430) );
  AOI22_X1 U13241 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10429) );
  AOI22_X1 U13242 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10428) );
  AOI22_X1 U13243 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13846), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U13244 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13245 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13246 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10433) );
  NAND3_X1 U13247 ( .A1(n10163), .A2(n10436), .A3(n10435), .ZN(n10817) );
  AOI22_X1 U13248 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13249 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13250 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10441) );
  AOI22_X1 U13251 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10440) );
  NAND4_X1 U13252 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10450) );
  AOI22_X1 U13253 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13255 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13256 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n14508), .ZN(n10445) );
  NAND4_X1 U13257 ( .A1(n10448), .A2(n10447), .A3(n10446), .A4(n10445), .ZN(
        n10449) );
  NAND2_X1 U13258 ( .A1(n10817), .A2(n10818), .ZN(n10821) );
  AOI22_X1 U13259 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14503), .B1(
        n10438), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10454) );
  AOI22_X1 U13260 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10453) );
  AOI22_X1 U13261 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13262 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10451) );
  NAND4_X1 U13263 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10462) );
  AOI22_X1 U13264 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10455), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10460) );
  AOI22_X1 U13265 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10472), .B1(
        n10456), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10459) );
  AOI22_X1 U13266 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10444), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10458) );
  AOI22_X1 U13267 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n14508), .ZN(n10457) );
  NAND4_X1 U13268 ( .A1(n10460), .A2(n10459), .A3(n10458), .A4(n10457), .ZN(
        n10461) );
  INV_X1 U13269 ( .A(n10823), .ZN(n10993) );
  OAI21_X1 U13270 ( .B1(n10821), .B2(n19514), .A(n10993), .ZN(n10825) );
  NAND2_X1 U13271 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10467) );
  NAND2_X1 U13272 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13273 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10465) );
  NAND2_X1 U13274 ( .A1(n10439), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10464) );
  NAND2_X1 U13275 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10471) );
  NAND2_X1 U13276 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13277 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13278 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14508), .ZN(
        n10468) );
  NAND2_X1 U13279 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10476) );
  NAND2_X1 U13280 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10475) );
  NAND2_X1 U13281 ( .A1(n13848), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10474) );
  NAND2_X1 U13282 ( .A1(n10455), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10473) );
  NAND2_X1 U13283 ( .A1(n10432), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10481) );
  NAND2_X1 U13284 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10480) );
  NAND2_X1 U13285 ( .A1(n10563), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10479) );
  NAND2_X1 U13286 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10478) );
  NAND4_X1 U13287 ( .A1(n10485), .A2(n10484), .A3(n10483), .A4(n10482), .ZN(
        n10486) );
  NAND2_X1 U13288 ( .A1(n10487), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10488) );
  NAND2_X1 U13289 ( .A1(n10489), .A2(n10488), .ZN(n10754) );
  NAND2_X1 U13290 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20166), .ZN(
        n10747) );
  NAND2_X1 U13291 ( .A1(n16647), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10490) );
  NOR2_X1 U13292 ( .A1(n10494), .A2(n10493), .ZN(n10495) );
  INV_X1 U13293 ( .A(n10745), .ZN(n10496) );
  NOR2_X1 U13294 ( .A1(n10043), .A2(n10496), .ZN(n10497) );
  MUX2_X1 U13295 ( .A(n10497), .B(P2_EBX_REG_3__SCAN_IN), .S(n11197), .Z(
        n10501) );
  AND2_X1 U13296 ( .A1(n11199), .A2(n10043), .ZN(n10539) );
  INV_X1 U13297 ( .A(n10539), .ZN(n10499) );
  NOR2_X1 U13298 ( .A1(n10499), .A2(n10498), .ZN(n10500) );
  NOR2_X1 U13299 ( .A1(n10501), .A2(n10500), .ZN(n10509) );
  INV_X1 U13300 ( .A(n10503), .ZN(n10504) );
  XNOR2_X1 U13301 ( .A(n10505), .B(n10504), .ZN(n10769) );
  NAND2_X1 U13302 ( .A1(n10502), .A2(n10769), .ZN(n10775) );
  MUX2_X1 U13303 ( .A(n10775), .B(P2_EBX_REG_2__SCAN_IN), .S(n11197), .Z(
        n10507) );
  NAND2_X1 U13304 ( .A1(n10539), .A2(n10823), .ZN(n10506) );
  NAND2_X1 U13305 ( .A1(n10507), .A2(n10506), .ZN(n10518) );
  NOR2_X1 U13306 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n10508) );
  MUX2_X1 U13307 ( .A(n10818), .B(n10508), .S(n11197), .Z(n10517) );
  AND3_X2 U13308 ( .A1(n10509), .A2(n10518), .A3(n10517), .ZN(n10579) );
  INV_X1 U13309 ( .A(n10579), .ZN(n10513) );
  INV_X1 U13310 ( .A(n10509), .ZN(n10511) );
  NAND2_X1 U13311 ( .A1(n10518), .A2(n10517), .ZN(n10510) );
  NAND2_X1 U13312 ( .A1(n10511), .A2(n10510), .ZN(n10512) );
  NAND2_X1 U13313 ( .A1(n10513), .A2(n10512), .ZN(n13607) );
  OAI21_X1 U13314 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20166), .A(
        n10747), .ZN(n10789) );
  INV_X1 U13315 ( .A(n10789), .ZN(n10750) );
  MUX2_X1 U13316 ( .A(n10750), .B(n10817), .S(n10043), .Z(n10773) );
  INV_X4 U13317 ( .A(n11199), .ZN(n11197) );
  MUX2_X1 U13318 ( .A(n10773), .B(P2_EBX_REG_0__SCAN_IN), .S(n11197), .Z(
        n19340) );
  NAND2_X1 U13319 ( .A1(n19340), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12955) );
  INV_X1 U13320 ( .A(n10517), .ZN(n10515) );
  NAND3_X1 U13321 ( .A1(n11197), .A2(P2_EBX_REG_0__SCAN_IN), .A3(
        P2_EBX_REG_1__SCAN_IN), .ZN(n10514) );
  NAND2_X1 U13322 ( .A1(n10515), .A2(n10514), .ZN(n15469) );
  NOR2_X1 U13323 ( .A1(n12955), .A2(n15469), .ZN(n10516) );
  NAND2_X1 U13324 ( .A1(n12955), .A2(n15469), .ZN(n12915) );
  OAI21_X1 U13325 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10516), .A(
        n12915), .ZN(n12809) );
  XNOR2_X1 U13326 ( .A(n10518), .B(n10517), .ZN(n15456) );
  XNOR2_X1 U13327 ( .A(n15456), .B(n10329), .ZN(n12808) );
  OR2_X1 U13328 ( .A1(n12809), .A2(n12808), .ZN(n12873) );
  INV_X1 U13329 ( .A(n15456), .ZN(n10519) );
  NAND2_X1 U13330 ( .A1(n10519), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10520) );
  AND2_X1 U13331 ( .A1(n12873), .A2(n10520), .ZN(n13447) );
  INV_X1 U13332 ( .A(n10521), .ZN(n10523) );
  INV_X1 U13333 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10522) );
  NOR2_X1 U13334 ( .A1(n10746), .A2(n10043), .ZN(n10526) );
  INV_X1 U13335 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10525) );
  MUX2_X1 U13336 ( .A(n10526), .B(n10525), .S(n11197), .Z(n10527) );
  INV_X1 U13337 ( .A(n10527), .ZN(n10541) );
  AOI22_X1 U13338 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10532) );
  AOI22_X1 U13339 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13340 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10530) );
  AOI22_X1 U13341 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10529) );
  NAND4_X1 U13342 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10538) );
  AOI22_X1 U13343 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10536) );
  INV_X1 U13344 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20774) );
  AOI22_X1 U13345 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13346 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U13347 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14508), .ZN(n10533) );
  NAND4_X1 U13348 ( .A1(n10536), .A2(n10535), .A3(n10534), .A4(n10533), .ZN(
        n10537) );
  NAND2_X1 U13349 ( .A1(n10539), .A2(n10542), .ZN(n10540) );
  XNOR2_X1 U13350 ( .A(n10579), .B(n10578), .ZN(n19320) );
  INV_X1 U13351 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13797) );
  XNOR2_X1 U13352 ( .A(n19320), .B(n13797), .ZN(n13793) );
  AOI22_X1 U13353 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19702), .B1(
        n19910), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10553) );
  INV_X1 U13354 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11100) );
  INV_X1 U13355 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14631) );
  OAI22_X1 U13356 ( .A1(n11100), .A2(n10416), .B1(n10543), .B2(n14631), .ZN(
        n10545) );
  INV_X1 U13357 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11098) );
  INV_X1 U13358 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13264) );
  OAI22_X1 U13359 ( .A1(n11098), .A2(n10405), .B1(n13252), .B2(n13264), .ZN(
        n10544) );
  NOR2_X1 U13360 ( .A1(n10545), .A2(n10544), .ZN(n10552) );
  AOI22_X1 U13361 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n10546), .B1(
        n10547), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13362 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n10548), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10550) );
  INV_X1 U13363 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14640) );
  INV_X1 U13364 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10556) );
  OAI22_X1 U13365 ( .A1(n14640), .A2(n10554), .B1(n10555), .B2(n10556), .ZN(
        n10559) );
  INV_X1 U13366 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14630) );
  INV_X1 U13367 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14639) );
  OAI22_X1 U13368 ( .A1(n14630), .A2(n19764), .B1(n10557), .B2(n14639), .ZN(
        n10558) );
  NOR2_X1 U13369 ( .A1(n10559), .A2(n10558), .ZN(n10562) );
  AOI22_X1 U13370 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n10560), .B1(
        n13886), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10561) );
  NAND3_X1 U13371 ( .A1(n9793), .A2(n10562), .A3(n10561), .ZN(n10575) );
  AOI22_X1 U13372 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10567) );
  AOI22_X1 U13373 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10566) );
  AOI22_X1 U13374 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10565) );
  AOI22_X1 U13375 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10564) );
  NAND4_X1 U13376 ( .A1(n10567), .A2(n10566), .A3(n10565), .A4(n10564), .ZN(
        n10573) );
  AOI22_X1 U13377 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13378 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13847), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13379 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13380 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14508), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10568) );
  NAND4_X1 U13381 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10572) );
  INV_X1 U13382 ( .A(n10577), .ZN(n11014) );
  NAND2_X1 U13383 ( .A1(n11014), .A2(n9740), .ZN(n10574) );
  NAND2_X1 U13384 ( .A1(n10836), .A2(n11020), .ZN(n10584) );
  INV_X1 U13385 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10576) );
  MUX2_X1 U13386 ( .A(n10577), .B(n10576), .S(n11197), .Z(n10580) );
  NAND2_X1 U13387 ( .A1(n10579), .A2(n10578), .ZN(n10582) );
  INV_X1 U13388 ( .A(n10580), .ZN(n10581) );
  NAND2_X1 U13389 ( .A1(n10582), .A2(n10581), .ZN(n10583) );
  NAND2_X1 U13390 ( .A1(n10624), .A2(n10583), .ZN(n13520) );
  INV_X1 U13391 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10961) );
  NAND2_X1 U13392 ( .A1(n10585), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10586) );
  NAND2_X1 U13393 ( .A1(n10587), .A2(n10586), .ZN(n13990) );
  INV_X1 U13394 ( .A(n10588), .ZN(n10589) );
  NAND2_X1 U13395 ( .A1(n13886), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10593) );
  NAND2_X1 U13396 ( .A1(n19702), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n10592) );
  NAND2_X1 U13397 ( .A1(n10560), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10591) );
  NAND2_X1 U13398 ( .A1(n19910), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10590) );
  NAND4_X1 U13399 ( .A1(n10593), .A2(n10592), .A3(n10591), .A4(n10590), .ZN(
        n10608) );
  AOI22_X1 U13400 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10546), .B1(
        n10549), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10606) );
  AOI22_X1 U13401 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10548), .B1(
        n10547), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10605) );
  INV_X1 U13402 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10594) );
  INV_X1 U13403 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14661) );
  OAI22_X1 U13404 ( .A1(n10594), .A2(n10405), .B1(n10554), .B2(n14661), .ZN(
        n10597) );
  INV_X1 U13405 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14650) );
  INV_X1 U13406 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10595) );
  OAI22_X1 U13407 ( .A1(n14650), .A2(n10543), .B1(n19764), .B2(n10595), .ZN(
        n10596) );
  NOR2_X1 U13408 ( .A1(n10597), .A2(n10596), .ZN(n10604) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10598) );
  INV_X1 U13410 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14659) );
  OAI22_X1 U13411 ( .A1(n10598), .A2(n10555), .B1(n10557), .B2(n14659), .ZN(
        n10602) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10600) );
  INV_X1 U13413 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10599) );
  OAI22_X1 U13414 ( .A1(n10600), .A2(n10416), .B1(n13252), .B2(n10599), .ZN(
        n10601) );
  NOR2_X1 U13415 ( .A1(n10602), .A2(n10601), .ZN(n10603) );
  NAND4_X1 U13416 ( .A1(n10606), .A2(n10605), .A3(n10604), .A4(n10603), .ZN(
        n10607) );
  AOI22_X1 U13417 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10612) );
  AOI22_X1 U13418 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U13419 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10610) );
  AOI22_X1 U13420 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10609) );
  NAND4_X1 U13421 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n10618) );
  AOI22_X1 U13422 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13423 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10615) );
  AOI22_X1 U13424 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10614) );
  AOI22_X1 U13425 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n14508), .ZN(n10613) );
  NAND4_X1 U13426 ( .A1(n10616), .A2(n10615), .A3(n10614), .A4(n10613), .ZN(
        n10617) );
  NAND2_X1 U13427 ( .A1(n11017), .A2(n9739), .ZN(n10619) );
  OR2_X1 U13428 ( .A1(n10621), .A2(n10840), .ZN(n10622) );
  NAND2_X1 U13429 ( .A1(n10621), .A2(n10840), .ZN(n10846) );
  INV_X1 U13430 ( .A(n11020), .ZN(n10626) );
  MUX2_X1 U13431 ( .A(n11017), .B(P2_EBX_REG_6__SCAN_IN), .S(n11197), .Z(
        n10623) );
  NAND2_X1 U13432 ( .A1(n10624), .A2(n10623), .ZN(n10625) );
  NAND2_X1 U13433 ( .A1(n9939), .A2(n10625), .ZN(n19307) );
  OAI21_X1 U13434 ( .B1(n10838), .B2(n10626), .A(n19307), .ZN(n10627) );
  INV_X1 U13435 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15989) );
  XNOR2_X1 U13436 ( .A(n10627), .B(n15989), .ZN(n13991) );
  NAND2_X1 U13437 ( .A1(n13990), .A2(n13991), .ZN(n10629) );
  NAND2_X1 U13438 ( .A1(n10627), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10628) );
  INV_X1 U13439 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10630) );
  MUX2_X1 U13440 ( .A(n10486), .B(n10630), .S(n11197), .Z(n10633) );
  AND2_X1 U13441 ( .A1(n11197), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10631) );
  XNOR2_X1 U13442 ( .A(n10639), .B(n10631), .ZN(n19284) );
  AND2_X1 U13443 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10632) );
  NAND2_X1 U13444 ( .A1(n19284), .A2(n10632), .ZN(n15773) );
  INV_X1 U13445 ( .A(n10633), .ZN(n10634) );
  XNOR2_X1 U13446 ( .A(n10635), .B(n10634), .ZN(n19297) );
  NAND2_X1 U13447 ( .A1(n19297), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15982) );
  NAND2_X1 U13448 ( .A1(n19284), .A2(n10626), .ZN(n10636) );
  INV_X1 U13449 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16609) );
  NAND2_X1 U13450 ( .A1(n10636), .A2(n16609), .ZN(n15774) );
  INV_X1 U13451 ( .A(n19297), .ZN(n10637) );
  INV_X1 U13452 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15984) );
  NAND2_X1 U13453 ( .A1(n10637), .A2(n15984), .ZN(n15981) );
  AND2_X1 U13454 ( .A1(n15774), .A2(n15981), .ZN(n10638) );
  INV_X1 U13455 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n13103) );
  AND2_X1 U13456 ( .A1(n11197), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10641) );
  XNOR2_X1 U13457 ( .A(n10642), .B(n10641), .ZN(n19277) );
  NAND2_X1 U13458 ( .A1(n19277), .A2(n10626), .ZN(n10652) );
  INV_X1 U13459 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16580) );
  NAND2_X1 U13460 ( .A1(n11197), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10643) );
  INV_X1 U13461 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13107) );
  MUX2_X1 U13462 ( .A(P2_EBX_REG_10__SCAN_IN), .B(n10643), .S(n10645), .Z(
        n10644) );
  NAND2_X1 U13463 ( .A1(n10644), .A2(n10725), .ZN(n19264) );
  OR2_X1 U13464 ( .A1(n19264), .A2(n11020), .ZN(n10653) );
  INV_X1 U13465 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16599) );
  NAND2_X1 U13466 ( .A1(n10653), .A2(n16599), .ZN(n15764) );
  NAND2_X1 U13467 ( .A1(n11197), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10646) );
  OR2_X1 U13468 ( .A1(n10647), .A2(n10646), .ZN(n10649) );
  INV_X1 U13469 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13272) );
  INV_X1 U13470 ( .A(n10654), .ZN(n10648) );
  NAND2_X1 U13471 ( .A1(n10649), .A2(n10648), .ZN(n13544) );
  INV_X1 U13472 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16594) );
  OR2_X1 U13473 ( .A1(n10651), .A2(n16594), .ZN(n16503) );
  NOR2_X1 U13474 ( .A1(n10652), .A2(n16580), .ZN(n15969) );
  NOR2_X1 U13475 ( .A1(n16599), .A2(n10653), .ZN(n15762) );
  NOR2_X1 U13476 ( .A1(n15969), .A2(n15762), .ZN(n16502) );
  AND2_X1 U13477 ( .A1(n16503), .A2(n16502), .ZN(n15646) );
  NAND2_X1 U13478 ( .A1(n11197), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10655) );
  NAND2_X1 U13479 ( .A1(n9942), .A2(n10656), .ZN(n10657) );
  INV_X1 U13480 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16571) );
  OR2_X1 U13481 ( .A1(n19248), .A2(n11020), .ZN(n10658) );
  AND2_X1 U13482 ( .A1(n11197), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13483 ( .A1(n11197), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10659) );
  INV_X1 U13484 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10660) );
  INV_X1 U13485 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n14074) );
  NAND2_X1 U13486 ( .A1(n10660), .A2(n14074), .ZN(n10661) );
  AND2_X1 U13487 ( .A1(n11197), .A2(n10661), .ZN(n10662) );
  INV_X1 U13488 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19202) );
  INV_X1 U13489 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10663) );
  NAND2_X1 U13490 ( .A1(n19202), .A2(n10663), .ZN(n10664) );
  INV_X1 U13491 ( .A(n10666), .ZN(n10667) );
  INV_X1 U13492 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10665) );
  AOI21_X1 U13493 ( .B1(n10668), .B2(n10667), .A(n10709), .ZN(n15437) );
  AOI21_X1 U13494 ( .B1(n15437), .B2(n10626), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15660) );
  NAND2_X1 U13495 ( .A1(n10681), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10669) );
  MUX2_X1 U13496 ( .A(n10681), .B(n10669), .S(n11197), .Z(n10670) );
  OR2_X1 U13497 ( .A1(n10681), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10672) );
  NAND2_X1 U13498 ( .A1(n19201), .A2(n10626), .ZN(n10671) );
  INV_X1 U13499 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15900) );
  NAND2_X1 U13500 ( .A1(n10671), .A2(n15900), .ZN(n15696) );
  NAND3_X1 U13501 ( .A1(n10672), .A2(P2_EBX_REG_19__SCAN_IN), .A3(n11197), 
        .ZN(n10673) );
  AND2_X1 U13502 ( .A1(n10673), .A2(n10675), .ZN(n19191) );
  NAND2_X1 U13503 ( .A1(n19191), .A2(n10626), .ZN(n10696) );
  INV_X1 U13504 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15891) );
  NAND2_X1 U13505 ( .A1(n10696), .A2(n15891), .ZN(n15686) );
  AND2_X1 U13506 ( .A1(n15696), .A2(n15686), .ZN(n15676) );
  AND2_X1 U13507 ( .A1(n11197), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10674) );
  XNOR2_X1 U13508 ( .A(n10675), .B(n10674), .ZN(n10704) );
  INV_X1 U13509 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15879) );
  OAI21_X1 U13510 ( .B1(n10704), .B2(n11020), .A(n15879), .ZN(n15675) );
  NAND2_X1 U13511 ( .A1(n15676), .A2(n15675), .ZN(n15656) );
  OR2_X1 U13512 ( .A1(n10690), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10680) );
  NAND3_X1 U13513 ( .A1(n10690), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n11197), 
        .ZN(n10676) );
  NAND3_X1 U13514 ( .A1(n10680), .A2(n10725), .A3(n10676), .ZN(n19214) );
  NOR2_X1 U13515 ( .A1(n19214), .A2(n11020), .ZN(n10678) );
  NAND2_X1 U13516 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10677) );
  OAI21_X1 U13517 ( .B1(n10678), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15651), .ZN(n15713) );
  AND2_X1 U13518 ( .A1(n11197), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13519 ( .A1(n10680), .A2(n10679), .ZN(n10682) );
  NAND2_X1 U13520 ( .A1(n10682), .A2(n10681), .ZN(n14203) );
  OR2_X1 U13521 ( .A1(n14203), .A2(n11020), .ZN(n10683) );
  INV_X1 U13522 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10852) );
  NAND2_X1 U13523 ( .A1(n10683), .A2(n10852), .ZN(n15654) );
  INV_X1 U13524 ( .A(n10684), .ZN(n10685) );
  XNOR2_X1 U13525 ( .A(n10693), .B(n10685), .ZN(n19237) );
  NAND2_X1 U13526 ( .A1(n19237), .A2(n10626), .ZN(n10686) );
  INV_X1 U13527 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15958) );
  NAND2_X1 U13528 ( .A1(n10686), .A2(n15958), .ZN(n15730) );
  INV_X1 U13529 ( .A(n10687), .ZN(n10688) );
  NAND3_X1 U13530 ( .A1(n10688), .A2(n11197), .A3(P2_EBX_REG_15__SCAN_IN), 
        .ZN(n10689) );
  NAND2_X1 U13531 ( .A1(n10690), .A2(n10689), .ZN(n19229) );
  INV_X1 U13532 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15944) );
  OAI21_X1 U13533 ( .B1(n19229), .B2(n11020), .A(n15944), .ZN(n15722) );
  NAND2_X1 U13534 ( .A1(n10693), .A2(n10692), .ZN(n13563) );
  OR2_X1 U13535 ( .A1(n13563), .A2(n11020), .ZN(n10694) );
  INV_X1 U13536 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15742) );
  NAND2_X1 U13537 ( .A1(n10694), .A2(n15742), .ZN(n15740) );
  NAND4_X1 U13538 ( .A1(n15654), .A2(n15730), .A3(n15722), .A4(n15740), .ZN(
        n10695) );
  NOR4_X1 U13539 ( .A1(n15660), .A2(n15656), .A3(n15713), .A4(n10695), .ZN(
        n10707) );
  NAND3_X1 U13540 ( .A1(n15437), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n10626), .ZN(n15658) );
  NOR2_X1 U13541 ( .A1(n10696), .A2(n15891), .ZN(n15655) );
  INV_X1 U13542 ( .A(n15651), .ZN(n10703) );
  NAND2_X1 U13543 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10697) );
  NOR2_X1 U13544 ( .A1(n14203), .A2(n10697), .ZN(n15652) );
  INV_X1 U13545 ( .A(n19229), .ZN(n10699) );
  AND2_X1 U13546 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10698) );
  NAND2_X1 U13547 ( .A1(n10699), .A2(n10698), .ZN(n15721) );
  AND2_X1 U13548 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10700) );
  NAND2_X1 U13549 ( .A1(n19237), .A2(n10700), .ZN(n15729) );
  NAND2_X1 U13550 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10701) );
  OR2_X1 U13551 ( .A1(n13563), .A2(n10701), .ZN(n15739) );
  NAND3_X1 U13552 ( .A1(n15721), .A2(n15729), .A3(n15739), .ZN(n10702) );
  NOR4_X1 U13553 ( .A1(n15655), .A2(n10703), .A3(n15652), .A4(n10702), .ZN(
        n10706) );
  INV_X1 U13554 ( .A(n10704), .ZN(n19177) );
  AND2_X1 U13555 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10705) );
  NAND2_X1 U13556 ( .A1(n19177), .A2(n10705), .ZN(n15674) );
  NAND3_X1 U13557 ( .A1(n19201), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n10626), .ZN(n15695) );
  NAND2_X1 U13558 ( .A1(n11197), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10708) );
  INV_X1 U13559 ( .A(n10708), .ZN(n10712) );
  AOI21_X1 U13560 ( .B1(n10712), .B2(n10711), .A(n10710), .ZN(n15424) );
  AOI21_X1 U13561 ( .B1(n15424), .B2(n10626), .A(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15851) );
  NAND3_X1 U13562 ( .A1(n15424), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n10626), .ZN(n15852) );
  NAND2_X1 U13563 ( .A1(n10717), .A2(n10713), .ZN(n15423) );
  XNOR2_X1 U13564 ( .A(n10714), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n16481) );
  NAND2_X1 U13565 ( .A1(n16480), .A2(n16481), .ZN(n10716) );
  INV_X1 U13566 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10715) );
  INV_X1 U13567 ( .A(n10717), .ZN(n10719) );
  NAND2_X1 U13568 ( .A1(n11197), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10718) );
  OAI211_X1 U13569 ( .C1(n10719), .C2(n10718), .A(n10725), .B(n10724), .ZN(
        n16455) );
  NOR2_X1 U13570 ( .A1(n16455), .A2(n11020), .ZN(n15637) );
  INV_X1 U13571 ( .A(n15637), .ZN(n10720) );
  NAND2_X1 U13572 ( .A1(n11197), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10721) );
  OR2_X1 U13573 ( .A1(n10728), .A2(n10721), .ZN(n10723) );
  INV_X1 U13574 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U13575 ( .A1(n10722), .A2(n10728), .ZN(n10735) );
  INV_X1 U13576 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10929) );
  NAND3_X1 U13577 ( .A1(n10724), .A2(P2_EBX_REG_25__SCAN_IN), .A3(n11197), 
        .ZN(n10726) );
  NAND2_X1 U13578 ( .A1(n10726), .A2(n10725), .ZN(n10727) );
  NOR2_X1 U13579 ( .A1(n10728), .A2(n10727), .ZN(n15395) );
  NAND2_X1 U13580 ( .A1(n15395), .A2(n10626), .ZN(n10730) );
  INV_X1 U13581 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15634) );
  INV_X1 U13582 ( .A(n10729), .ZN(n16447) );
  NAND2_X1 U13583 ( .A1(n10626), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10732) );
  INV_X1 U13584 ( .A(n10730), .ZN(n10731) );
  NAND2_X1 U13585 ( .A1(n10731), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15624) );
  OAI21_X1 U13586 ( .B1(n16447), .B2(n10732), .A(n15624), .ZN(n11186) );
  INV_X1 U13587 ( .A(n14424), .ZN(n10733) );
  NAND2_X1 U13588 ( .A1(n11197), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10734) );
  INV_X1 U13589 ( .A(n10734), .ZN(n10736) );
  NAND2_X1 U13590 ( .A1(n10736), .A2(n10735), .ZN(n10737) );
  NAND2_X1 U13591 ( .A1(n11195), .A2(n10737), .ZN(n15385) );
  NOR2_X1 U13592 ( .A1(n15385), .A2(n11020), .ZN(n10740) );
  INV_X1 U13593 ( .A(n10738), .ZN(n10739) );
  NAND2_X1 U13594 ( .A1(n11197), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11193) );
  XNOR2_X1 U13595 ( .A(n11195), .B(n11193), .ZN(n16432) );
  NAND2_X1 U13596 ( .A1(n16432), .A2(n10626), .ZN(n11187) );
  XOR2_X1 U13597 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n11187), .Z(
        n10741) );
  XNOR2_X1 U13598 ( .A(n10742), .B(n10741), .ZN(n14373) );
  INV_X1 U13599 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16673) );
  NOR2_X1 U13600 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16673), .ZN(
        n10743) );
  NAND2_X1 U13601 ( .A1(n10754), .A2(n10747), .ZN(n10774) );
  NAND2_X1 U13602 ( .A1(n10748), .A2(n10774), .ZN(n10770) );
  INV_X1 U13603 ( .A(n10770), .ZN(n10749) );
  OAI21_X1 U13604 ( .B1(n19514), .B2(n10750), .A(n10749), .ZN(n10752) );
  NAND2_X1 U13605 ( .A1(n9740), .A2(n10769), .ZN(n10751) );
  NAND2_X1 U13606 ( .A1(n10752), .A2(n10751), .ZN(n10753) );
  NAND2_X1 U13607 ( .A1(n10753), .A2(n20179), .ZN(n10760) );
  OAI21_X1 U13608 ( .B1(n10789), .B2(n10754), .A(n10043), .ZN(n10759) );
  NAND2_X1 U13609 ( .A1(n10755), .A2(n19514), .ZN(n10757) );
  INV_X1 U13610 ( .A(n10769), .ZN(n10756) );
  NAND2_X1 U13611 ( .A1(n10757), .A2(n10756), .ZN(n10758) );
  AOI22_X1 U13612 ( .A1(n10760), .A2(n10759), .B1(n10758), .B2(n10775), .ZN(
        n10761) );
  NAND2_X1 U13613 ( .A1(n10777), .A2(n10761), .ZN(n10762) );
  OAI21_X1 U13614 ( .B1(n10777), .B2(n10502), .A(n10762), .ZN(n10763) );
  OR2_X1 U13615 ( .A1(n10781), .A2(n10763), .ZN(n10764) );
  MUX2_X1 U13616 ( .A(n10764), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19151), .Z(n10767) );
  NAND2_X1 U13617 ( .A1(n10781), .A2(n12725), .ZN(n10765) );
  NAND2_X1 U13618 ( .A1(n12859), .A2(n19514), .ZN(n12723) );
  NAND2_X1 U13619 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20061), .ZN(n20194) );
  INV_X2 U13620 ( .A(n20194), .ZN(n20193) );
  NAND2_X1 U13621 ( .A1(n20193), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20119) );
  NOR2_X1 U13622 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20062) );
  INV_X1 U13623 ( .A(n20062), .ZN(n20074) );
  NAND3_X1 U13624 ( .A1(n20061), .A2(n20115), .A3(n20074), .ZN(n20068) );
  NAND2_X1 U13625 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20190) );
  INV_X1 U13626 ( .A(n20190), .ZN(n20183) );
  NOR2_X1 U13627 ( .A1(n20068), .A2(n20183), .ZN(n12688) );
  NAND2_X1 U13628 ( .A1(n10766), .A2(n12688), .ZN(n10812) );
  AOI21_X1 U13629 ( .B1(n10767), .B2(n20179), .A(n10267), .ZN(n10768) );
  NAND2_X1 U13630 ( .A1(n12723), .A2(n10768), .ZN(n10811) );
  NAND2_X1 U13631 ( .A1(n10777), .A2(n10769), .ZN(n10788) );
  NOR2_X1 U13632 ( .A1(n10770), .A2(n10788), .ZN(n10771) );
  OR2_X1 U13633 ( .A1(n10781), .A2(n10771), .ZN(n16657) );
  MUX2_X1 U13634 ( .A(n10794), .B(n10766), .S(n9739), .Z(n10772) );
  NAND2_X1 U13635 ( .A1(n10772), .A2(n20190), .ZN(n10793) );
  NAND3_X1 U13636 ( .A1(n10777), .A2(n10774), .A3(n10773), .ZN(n10779) );
  INV_X1 U13637 ( .A(n10775), .ZN(n10776) );
  NAND2_X1 U13638 ( .A1(n10777), .A2(n10776), .ZN(n10778) );
  NAND2_X1 U13639 ( .A1(n10779), .A2(n10778), .ZN(n10780) );
  OR2_X1 U13640 ( .A1(n10781), .A2(n10780), .ZN(n20172) );
  INV_X1 U13641 ( .A(n20172), .ZN(n10782) );
  NAND2_X1 U13642 ( .A1(n9740), .A2(n19503), .ZN(n10797) );
  NOR2_X1 U13643 ( .A1(n10814), .A2(n10797), .ZN(n20171) );
  NAND2_X1 U13644 ( .A1(n10782), .A2(n20171), .ZN(n12664) );
  INV_X1 U13645 ( .A(n10814), .ZN(n16652) );
  NAND2_X1 U13646 ( .A1(n10784), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13647 ( .A1(n10785), .A2(n12700), .ZN(n16650) );
  INV_X1 U13648 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n20943) );
  OAI21_X1 U13649 ( .B1(n10456), .B2(n16650), .A(n20943), .ZN(n10786) );
  AND2_X1 U13650 ( .A1(n10786), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20163) );
  NOR2_X1 U13651 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n16657), .ZN(n10787) );
  OAI21_X1 U13652 ( .B1(n10789), .B2(n10788), .A(n10787), .ZN(n10790) );
  INV_X1 U13653 ( .A(n10790), .ZN(n10791) );
  NOR2_X1 U13654 ( .A1(n20163), .A2(n10791), .ZN(n20169) );
  INV_X1 U13655 ( .A(n20169), .ZN(n12662) );
  NAND3_X1 U13656 ( .A1(n16652), .A2(n19514), .A3(n12662), .ZN(n10792) );
  OAI211_X1 U13657 ( .C1(n16657), .C2(n10793), .A(n12664), .B(n10792), .ZN(
        n10809) );
  NAND2_X1 U13658 ( .A1(n10794), .A2(n12688), .ZN(n10795) );
  OR2_X1 U13659 ( .A1(n16657), .A2(n10795), .ZN(n10808) );
  INV_X1 U13660 ( .A(n10797), .ZN(n10798) );
  OAI21_X1 U13661 ( .B1(n10796), .B2(n13430), .A(n10798), .ZN(n10944) );
  NAND2_X1 U13662 ( .A1(n10800), .A2(n10941), .ZN(n10801) );
  NAND2_X1 U13663 ( .A1(n16656), .A2(n10801), .ZN(n10806) );
  OAI21_X1 U13664 ( .B1(n10267), .B2(n19514), .A(n20179), .ZN(n10802) );
  NAND2_X1 U13665 ( .A1(n10802), .A2(n10973), .ZN(n10803) );
  AOI21_X1 U13666 ( .B1(n10803), .B2(n10941), .A(n10298), .ZN(n10805) );
  AND4_X1 U13667 ( .A1(n10944), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10807) );
  NAND2_X1 U13668 ( .A1(n10808), .A2(n10807), .ZN(n12691) );
  NOR2_X1 U13669 ( .A1(n10809), .A2(n12691), .ZN(n10810) );
  OAI211_X1 U13670 ( .C1(n12723), .C2(n10812), .A(n10811), .B(n10810), .ZN(
        n10813) );
  NAND2_X1 U13671 ( .A1(n16011), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20059) );
  NOR2_X1 U13672 ( .A1(n10814), .A2(n10502), .ZN(n20170) );
  XNOR2_X1 U13673 ( .A(n10815), .B(n11010), .ZN(n13791) );
  NAND2_X1 U13674 ( .A1(n13791), .A2(n13797), .ZN(n10832) );
  INV_X1 U13675 ( .A(n10817), .ZN(n12960) );
  NAND3_X1 U13676 ( .A1(n12960), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n10818), .ZN(n10820) );
  NOR2_X1 U13677 ( .A1(n10817), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10819) );
  INV_X1 U13678 ( .A(n10818), .ZN(n10990) );
  XOR2_X1 U13679 ( .A(n10819), .B(n10990), .Z(n12912) );
  NAND2_X1 U13680 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12912), .ZN(
        n12911) );
  NAND2_X1 U13681 ( .A1(n10820), .A2(n12911), .ZN(n10826) );
  XNOR2_X1 U13682 ( .A(n10329), .B(n10826), .ZN(n12806) );
  INV_X1 U13683 ( .A(n10821), .ZN(n10822) );
  NAND2_X1 U13684 ( .A1(n10823), .A2(n10822), .ZN(n10824) );
  NAND2_X1 U13685 ( .A1(n10825), .A2(n10824), .ZN(n12807) );
  NAND2_X1 U13686 ( .A1(n12806), .A2(n12807), .ZN(n10828) );
  NAND2_X1 U13687 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10826), .ZN(
        n10827) );
  NAND2_X1 U13688 ( .A1(n10828), .A2(n10827), .ZN(n10829) );
  XNOR2_X1 U13689 ( .A(n10829), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13451) );
  NAND2_X1 U13690 ( .A1(n10829), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10830) );
  NAND2_X1 U13691 ( .A1(n10831), .A2(n10830), .ZN(n13790) );
  NAND2_X1 U13692 ( .A1(n10832), .A2(n13790), .ZN(n10835) );
  INV_X1 U13693 ( .A(n13791), .ZN(n10833) );
  NAND2_X1 U13694 ( .A1(n10833), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10834) );
  INV_X1 U13695 ( .A(n10836), .ZN(n10837) );
  NAND2_X1 U13696 ( .A1(n10837), .A2(n10961), .ZN(n16531) );
  NAND2_X1 U13697 ( .A1(n16533), .A2(n16531), .ZN(n10842) );
  NAND2_X1 U13698 ( .A1(n10842), .A2(n16532), .ZN(n10844) );
  INV_X1 U13699 ( .A(n10838), .ZN(n10843) );
  NAND2_X1 U13700 ( .A1(n10844), .A2(n10843), .ZN(n10845) );
  NAND2_X1 U13701 ( .A1(n10846), .A2(n11020), .ZN(n10847) );
  NAND2_X1 U13702 ( .A1(n10850), .A2(n10847), .ZN(n15985) );
  XNOR2_X1 U13703 ( .A(n10850), .B(n16609), .ZN(n15777) );
  AND2_X1 U13704 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16582) );
  AND2_X1 U13705 ( .A1(n16582), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15915) );
  NAND2_X1 U13706 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15957) );
  NOR2_X1 U13707 ( .A1(n15957), .A2(n15958), .ZN(n15916) );
  AND2_X1 U13708 ( .A1(n15915), .A2(n15916), .ZN(n15896) );
  NAND2_X1 U13709 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15919) );
  NOR2_X1 U13710 ( .A1(n15919), .A2(n10852), .ZN(n15899) );
  AND2_X1 U13711 ( .A1(n15896), .A2(n15899), .ZN(n15901) );
  NAND2_X1 U13712 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15861) );
  INV_X1 U13713 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10853) );
  NOR2_X1 U13714 ( .A1(n15861), .A2(n10853), .ZN(n11181) );
  NAND2_X1 U13715 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16543) );
  INV_X1 U13716 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15810) );
  NAND2_X1 U13717 ( .A1(n14371), .A2(n16624), .ZN(n11185) );
  INV_X1 U13718 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10858) );
  NAND2_X1 U13719 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10857) );
  NAND2_X1 U13720 ( .A1(n10339), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10856) );
  OAI211_X1 U13721 ( .C1(n14432), .C2(n10858), .A(n10857), .B(n10856), .ZN(
        n10859) );
  INV_X1 U13722 ( .A(n10859), .ZN(n10860) );
  OAI21_X1 U13723 ( .B1(n11210), .B2(n15984), .A(n10860), .ZN(n13091) );
  INV_X1 U13724 ( .A(n10862), .ZN(n10864) );
  NAND2_X1 U13725 ( .A1(n10864), .A2(n10863), .ZN(n10865) );
  INV_X1 U13726 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U13727 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10867) );
  NAND2_X1 U13728 ( .A1(n10339), .A2(P2_EBX_REG_4__SCAN_IN), .ZN(n10866) );
  OAI211_X1 U13729 ( .C1(n14432), .C2(n10868), .A(n10867), .B(n10866), .ZN(
        n10869) );
  AOI21_X1 U13730 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n10869), .ZN(n13014) );
  AOI22_X1 U13731 ( .A1(n10339), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10871) );
  INV_X1 U13732 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13523) );
  OR2_X1 U13733 ( .A1(n14432), .A2(n13523), .ZN(n10870) );
  OAI211_X1 U13734 ( .C1(n11210), .C2(n10961), .A(n10871), .B(n10870), .ZN(
        n13020) );
  INV_X1 U13735 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n14014) );
  NAND2_X1 U13736 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10873) );
  NAND2_X1 U13737 ( .A1(n10339), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10872) );
  OAI211_X1 U13738 ( .C1(n14432), .C2(n14014), .A(n10873), .B(n10872), .ZN(
        n10874) );
  AOI21_X1 U13739 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10874), .ZN(n13069) );
  AOI22_X1 U13740 ( .A1(n10339), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10876) );
  NAND2_X1 U13741 ( .A1(n11205), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10875) );
  OAI211_X1 U13742 ( .C1(n11210), .C2(n16609), .A(n10876), .B(n10875), .ZN(
        n13098) );
  AOI22_X1 U13743 ( .A1(n10339), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10878) );
  NAND2_X1 U13744 ( .A1(n11205), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10877) );
  OAI211_X1 U13745 ( .C1(n11210), .C2(n16580), .A(n10878), .B(n10877), .ZN(
        n13104) );
  INV_X1 U13746 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U13747 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10880) );
  NAND2_X1 U13748 ( .A1(n10339), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10879) );
  OAI211_X1 U13749 ( .C1(n14432), .C2(n11067), .A(n10880), .B(n10879), .ZN(
        n10881) );
  AOI21_X1 U13750 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10881), .ZN(n13111) );
  NOR2_X2 U13751 ( .A1(n13110), .A2(n13111), .ZN(n13268) );
  INV_X1 U13752 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U13753 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10883) );
  NAND2_X1 U13754 ( .A1(n9725), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10882) );
  OAI211_X1 U13755 ( .C1(n14432), .C2(n11083), .A(n10883), .B(n10882), .ZN(
        n10884) );
  INV_X1 U13756 ( .A(n10884), .ZN(n10885) );
  OAI21_X1 U13757 ( .B1(n11210), .B2(n16594), .A(n10885), .ZN(n13269) );
  NAND2_X1 U13758 ( .A1(n13268), .A2(n13269), .ZN(n13271) );
  INV_X1 U13759 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U13760 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U13761 ( .A1(n10339), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10886) );
  OAI211_X1 U13762 ( .C1(n14432), .C2(n11097), .A(n10887), .B(n10886), .ZN(
        n10888) );
  AOI21_X1 U13763 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10888), .ZN(n13187) );
  INV_X1 U13764 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13765 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10890) );
  NAND2_X1 U13766 ( .A1(n9725), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10889) );
  OAI211_X1 U13767 ( .C1(n14432), .C2(n10891), .A(n10890), .B(n10889), .ZN(
        n10892) );
  AOI21_X1 U13768 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10892), .ZN(n13398) );
  INV_X1 U13769 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11129) );
  NAND2_X1 U13770 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U13771 ( .A1(n10339), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10893) );
  OAI211_X1 U13772 ( .C1(n14432), .C2(n11129), .A(n10894), .B(n10893), .ZN(
        n10895) );
  AOI21_X1 U13773 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10895), .ZN(n13462) );
  NOR2_X4 U13774 ( .A1(n13461), .A2(n13462), .ZN(n13820) );
  AOI22_X1 U13775 ( .A1(n9725), .A2(P2_EBX_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10897) );
  INV_X1 U13776 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20910) );
  OR2_X1 U13777 ( .A1(n14432), .A2(n20910), .ZN(n10896) );
  OAI211_X1 U13778 ( .C1(n11210), .C2(n15944), .A(n10897), .B(n10896), .ZN(
        n13819) );
  INV_X1 U13779 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n20808) );
  NAND2_X1 U13780 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10899) );
  NAND2_X1 U13781 ( .A1(n10339), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10898) );
  OAI211_X1 U13782 ( .C1(n14432), .C2(n20808), .A(n10899), .B(n10898), .ZN(
        n10900) );
  AOI21_X1 U13783 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10900), .ZN(n13878) );
  INV_X1 U13784 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20097) );
  NAND2_X1 U13785 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10902) );
  NAND2_X1 U13786 ( .A1(n9725), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10901) );
  OAI211_X1 U13787 ( .C1(n14432), .C2(n20097), .A(n10902), .B(n10901), .ZN(
        n10903) );
  AOI21_X1 U13788 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10903), .ZN(n14071) );
  AOI22_X1 U13789 ( .A1(n9725), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10905) );
  INV_X1 U13790 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20099) );
  OR2_X1 U13791 ( .A1(n14432), .A2(n20099), .ZN(n10904) );
  OAI211_X1 U13792 ( .C1(n11210), .C2(n15900), .A(n10905), .B(n10904), .ZN(
        n14199) );
  AOI22_X1 U13793 ( .A1(n9725), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10907) );
  NAND2_X1 U13794 ( .A1(n11205), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10906) );
  OAI211_X1 U13795 ( .C1(n11210), .C2(n15891), .A(n10907), .B(n10906), .ZN(
        n14222) );
  NAND2_X1 U13796 ( .A1(n14198), .A2(n14222), .ZN(n14221) );
  INV_X1 U13797 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20103) );
  NAND2_X1 U13798 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10909) );
  NAND2_X1 U13799 ( .A1(n9725), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10908) );
  OAI211_X1 U13800 ( .C1(n14432), .C2(n20103), .A(n10909), .B(n10908), .ZN(
        n10910) );
  AOI21_X1 U13801 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10910), .ZN(n15532) );
  OR2_X2 U13802 ( .A1(n14221), .A2(n15532), .ZN(n15535) );
  INV_X1 U13803 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n15663) );
  NAND2_X1 U13804 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U13805 ( .A1(n10339), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10911) );
  OAI211_X1 U13806 ( .C1(n14432), .C2(n15663), .A(n10912), .B(n10911), .ZN(
        n10913) );
  AOI21_X1 U13807 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10913), .ZN(n15440) );
  INV_X1 U13808 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16546) );
  AOI22_X1 U13809 ( .A1(n9725), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10915) );
  NAND2_X1 U13810 ( .A1(n11205), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10914) );
  OAI211_X1 U13811 ( .C1(n11210), .C2(n16546), .A(n10915), .B(n10914), .ZN(
        n15427) );
  INV_X1 U13812 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n11157) );
  NAND2_X1 U13813 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10917) );
  NAND2_X1 U13814 ( .A1(n9725), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10916) );
  OAI211_X1 U13815 ( .C1(n14432), .C2(n11157), .A(n10917), .B(n10916), .ZN(
        n10918) );
  AOI21_X1 U13816 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10918), .ZN(n15413) );
  INV_X1 U13817 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20109) );
  NAND2_X1 U13818 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10920) );
  NAND2_X1 U13819 ( .A1(n10339), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10919) );
  OAI211_X1 U13820 ( .C1(n14432), .C2(n20109), .A(n10920), .B(n10919), .ZN(
        n10921) );
  AOI21_X1 U13821 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10921), .ZN(n15516) );
  INV_X1 U13822 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n10925) );
  NAND2_X1 U13823 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10924) );
  NAND2_X1 U13824 ( .A1(n9725), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10923) );
  OAI211_X1 U13825 ( .C1(n14432), .C2(n10925), .A(n10924), .B(n10923), .ZN(
        n10926) );
  AOI21_X1 U13826 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10926), .ZN(n15399) );
  AOI22_X1 U13827 ( .A1(n10339), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10928) );
  INV_X1 U13828 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20111) );
  OR2_X1 U13829 ( .A1(n14432), .A2(n20111), .ZN(n10927) );
  OAI211_X1 U13830 ( .C1(n11210), .C2(n10929), .A(n10928), .B(n10927), .ZN(
        n15499) );
  NAND2_X1 U13831 ( .A1(n15398), .A2(n15499), .ZN(n15379) );
  INV_X1 U13832 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n15608) );
  NAND2_X1 U13833 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10931) );
  NAND2_X1 U13834 ( .A1(n9725), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10930) );
  OAI211_X1 U13835 ( .C1(n14432), .C2(n15608), .A(n10931), .B(n10930), .ZN(
        n10932) );
  AOI21_X1 U13836 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10932), .ZN(n15380) );
  INV_X1 U13837 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n20113) );
  NAND2_X1 U13838 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U13839 ( .A1(n9725), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10933) );
  OAI211_X1 U13840 ( .C1(n14432), .C2(n20113), .A(n10934), .B(n10933), .ZN(
        n10935) );
  AOI21_X1 U13841 ( .B1(n10936), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10935), .ZN(n10937) );
  AND2_X1 U13842 ( .A1(n15382), .A2(n10937), .ZN(n10938) );
  OR2_X1 U13843 ( .A1(n10938), .A2(n15344), .ZN(n15488) );
  INV_X1 U13844 ( .A(n15488), .ZN(n16434) );
  NAND2_X1 U13845 ( .A1(n11173), .A2(n10939), .ZN(n19491) );
  AND3_X1 U13846 ( .A1(n9740), .A2(n10941), .A3(n10212), .ZN(n10942) );
  AND2_X1 U13847 ( .A1(n10940), .A2(n10942), .ZN(n16658) );
  INV_X1 U13848 ( .A(n15924), .ZN(n10957) );
  NAND2_X1 U13849 ( .A1(n10943), .A2(n19514), .ZN(n15999) );
  NAND2_X1 U13850 ( .A1(n15999), .A2(n10944), .ZN(n10952) );
  NAND2_X1 U13851 ( .A1(n10947), .A2(n10946), .ZN(n13423) );
  NAND2_X1 U13852 ( .A1(n19503), .A2(n10766), .ZN(n10949) );
  INV_X1 U13853 ( .A(n12660), .ZN(n20181) );
  OAI21_X1 U13854 ( .B1(n10298), .B2(n10287), .A(n20181), .ZN(n10948) );
  NAND4_X1 U13855 ( .A1(n10950), .A2(n13423), .A3(n10949), .A4(n10948), .ZN(
        n10951) );
  AOI21_X1 U13856 ( .B1(n10952), .B2(n13890), .A(n10951), .ZN(n10953) );
  OAI21_X1 U13857 ( .B1(n10955), .B2(n10954), .A(n10953), .ZN(n16043) );
  OR2_X1 U13858 ( .A1(n16043), .A2(n16018), .ZN(n10956) );
  NAND2_X1 U13859 ( .A1(n11173), .A2(n10956), .ZN(n15925) );
  AND2_X1 U13860 ( .A1(n15901), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11180) );
  INV_X1 U13861 ( .A(n11180), .ZN(n10965) );
  INV_X1 U13862 ( .A(n11173), .ZN(n10959) );
  NAND2_X1 U13863 ( .A1(n16011), .A2(n19670), .ZN(n20133) );
  NOR2_X1 U13864 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20133), .ZN(n10958) );
  AND2_X1 U13865 ( .A1(n10958), .A2(n20182), .ZN(n19461) );
  INV_X2 U13866 ( .A(n19461), .ZN(n19304) );
  NAND2_X1 U13867 ( .A1(n10959), .A2(n19304), .ZN(n19494) );
  INV_X1 U13868 ( .A(n19494), .ZN(n10960) );
  OR2_X1 U13869 ( .A1(n15952), .A2(n10960), .ZN(n16578) );
  NOR2_X1 U13870 ( .A1(n13797), .A2(n10961), .ZN(n11178) );
  INV_X1 U13871 ( .A(n11178), .ZN(n16626) );
  INV_X1 U13872 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19493) );
  NOR2_X1 U13873 ( .A1(n19493), .A2(n12964), .ZN(n19486) );
  INV_X1 U13874 ( .A(n19486), .ZN(n12819) );
  NAND3_X1 U13875 ( .A1(n15924), .A2(n10329), .A3(n12819), .ZN(n12815) );
  INV_X1 U13876 ( .A(n15925), .ZN(n10962) );
  OAI21_X1 U13877 ( .B1(n10329), .B2(n12819), .A(n10962), .ZN(n10963) );
  NAND4_X1 U13878 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12815), .A3(
        n19494), .A4(n10963), .ZN(n13795) );
  NOR2_X1 U13879 ( .A1(n16626), .A2(n13795), .ZN(n13996) );
  AND3_X1 U13880 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10964) );
  NAND2_X1 U13881 ( .A1(n13996), .A2(n10964), .ZN(n16579) );
  AND2_X1 U13882 ( .A1(n16578), .A2(n16579), .ZN(n15972) );
  AOI21_X1 U13883 ( .B1(n15952), .B2(n10965), .A(n15972), .ZN(n15886) );
  INV_X1 U13884 ( .A(n11181), .ZN(n10966) );
  NAND2_X1 U13885 ( .A1(n15952), .A2(n10966), .ZN(n10967) );
  AND2_X1 U13886 ( .A1(n15886), .A2(n10967), .ZN(n16555) );
  NAND2_X1 U13887 ( .A1(n15952), .A2(n16543), .ZN(n10968) );
  NAND2_X1 U13888 ( .A1(n16555), .A2(n10968), .ZN(n15813) );
  INV_X1 U13889 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15840) );
  NAND2_X1 U13890 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10969) );
  NOR2_X1 U13891 ( .A1(n15840), .A2(n10969), .ZN(n11182) );
  INV_X1 U13892 ( .A(n11182), .ZN(n10970) );
  AND2_X1 U13893 ( .A1(n15952), .A2(n10970), .ZN(n10971) );
  OR2_X1 U13894 ( .A1(n15813), .A2(n10971), .ZN(n15806) );
  AND2_X1 U13895 ( .A1(n15952), .A2(n15810), .ZN(n10972) );
  NOR2_X1 U13896 ( .A1(n15806), .A2(n10972), .ZN(n15787) );
  INV_X1 U13897 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11175) );
  NAND2_X1 U13898 ( .A1(n19326), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n14368) );
  INV_X1 U13899 ( .A(n10272), .ZN(n13429) );
  NAND2_X1 U13900 ( .A1(n13429), .A2(n9727), .ZN(n10994) );
  NOR2_X1 U13901 ( .A1(n10973), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10996) );
  AND2_X1 U13902 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10974) );
  NOR2_X1 U13903 ( .A1(n10996), .A2(n10974), .ZN(n10975) );
  NAND2_X1 U13904 ( .A1(n10994), .A2(n10975), .ZN(n10978) );
  NOR2_X1 U13905 ( .A1(n10278), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10976) );
  NOR2_X1 U13906 ( .A1(n12960), .A2(n11140), .ZN(n10977) );
  INV_X1 U13907 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U13908 ( .A1(n10980), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10981) );
  OAI211_X1 U13909 ( .C1(n10973), .C2(n10982), .A(n10981), .B(n19670), .ZN(
        n10983) );
  INV_X1 U13910 ( .A(n10983), .ZN(n10984) );
  OAI21_X1 U13911 ( .B1(n14444), .B2(n10985), .A(n10984), .ZN(n12957) );
  INV_X1 U13912 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13913 ( .A1(n10996), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n9727), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13914 ( .A1(n10272), .A2(n10973), .ZN(n10988) );
  MUX2_X1 U13915 ( .A(n10988), .B(n20159), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10989) );
  NAND2_X1 U13916 ( .A1(n10991), .A2(n12956), .ZN(n10992) );
  OR2_X1 U13917 ( .A1(n11140), .A2(n10993), .ZN(n10995) );
  OAI211_X1 U13918 ( .C1(n19670), .C2(n20149), .A(n10995), .B(n10994), .ZN(
        n10999) );
  XNOR2_X1 U13919 ( .A(n11000), .B(n10999), .ZN(n12811) );
  NAND2_X1 U13920 ( .A1(n11211), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U13921 ( .A1(n14442), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11215), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10997) );
  INV_X1 U13922 ( .A(n10999), .ZN(n11001) );
  NAND2_X1 U13923 ( .A1(n11001), .A2(n11000), .ZN(n11002) );
  NAND2_X1 U13924 ( .A1(n12812), .A2(n11002), .ZN(n13415) );
  INV_X1 U13925 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13926 ( .A1(n11215), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11003) );
  OAI21_X1 U13927 ( .B1(n14444), .B2(n11004), .A(n11003), .ZN(n11008) );
  NAND2_X1 U13928 ( .A1(n14442), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n11005) );
  OAI21_X1 U13929 ( .B1(n11140), .B2(n11006), .A(n11005), .ZN(n11007) );
  AOI22_X1 U13930 ( .A1(n11211), .A2(P2_REIP_REG_4__SCAN_IN), .B1(n14442), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11013) );
  OAI22_X1 U13931 ( .A1(n11140), .A2(n11010), .B1(n11038), .B2(n13797), .ZN(
        n11011) );
  INV_X1 U13932 ( .A(n11011), .ZN(n11012) );
  NAND2_X1 U13933 ( .A1(n11013), .A2(n11012), .ZN(n13421) );
  AOI22_X1 U13934 ( .A1(n14442), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11215), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11016) );
  OR2_X1 U13935 ( .A1(n11140), .A2(n11014), .ZN(n11015) );
  OAI211_X1 U13936 ( .C1(n14444), .C2(n13523), .A(n11016), .B(n11015), .ZN(
        n13509) );
  NAND2_X1 U13937 ( .A1(n13419), .A2(n13509), .ZN(n13508) );
  OR2_X1 U13938 ( .A1(n11140), .A2(n11017), .ZN(n11018) );
  AOI22_X1 U13939 ( .A1(n14442), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n11215), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n11019) );
  OAI21_X1 U13940 ( .B1(n14444), .B2(n14014), .A(n11019), .ZN(n14000) );
  NAND2_X1 U13941 ( .A1(n13998), .A2(n14000), .ZN(n13999) );
  OR2_X1 U13942 ( .A1(n11140), .A2(n11020), .ZN(n11021) );
  NAND2_X1 U13943 ( .A1(n11211), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U13944 ( .A1(n14442), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n11215), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n11022) );
  INV_X1 U13945 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11037) );
  INV_X1 U13946 ( .A(n11140), .ZN(n11126) );
  AOI22_X1 U13947 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13948 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U13949 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11026) );
  AOI22_X1 U13950 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11025) );
  NAND4_X1 U13951 ( .A1(n11028), .A2(n11027), .A3(n11026), .A4(n11025), .ZN(
        n11034) );
  AOI22_X1 U13952 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U13953 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10456), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U13954 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11030) );
  AOI22_X1 U13955 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14508), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11029) );
  NAND4_X1 U13956 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11033) );
  NAND2_X1 U13957 ( .A1(n11126), .A2(n13115), .ZN(n11036) );
  AOI22_X1 U13958 ( .A1(n14442), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11215), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11035) );
  OAI211_X1 U13959 ( .C1(n11037), .C2(n14444), .A(n11036), .B(n11035), .ZN(
        n16608) );
  INV_X1 U13960 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U13961 ( .A1(n14442), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n11215), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11053) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11040) );
  INV_X1 U13963 ( .A(n14503), .ZN(n11101) );
  INV_X1 U13964 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11039) );
  OAI22_X1 U13965 ( .A1(n11040), .A2(n11101), .B1(n11099), .B2(n11039), .ZN(
        n11041) );
  INV_X1 U13966 ( .A(n11041), .ZN(n11045) );
  AOI22_X1 U13967 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U13968 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10528), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U13969 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11042) );
  NAND4_X1 U13970 ( .A1(n11045), .A2(n11044), .A3(n11043), .A4(n11042), .ZN(
        n11051) );
  AOI22_X1 U13971 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U13972 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U13973 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13974 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14508), .ZN(n11046) );
  NAND4_X1 U13975 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n11050) );
  NOR2_X1 U13976 ( .A1(n11051), .A2(n11050), .ZN(n13119) );
  OR2_X1 U13977 ( .A1(n11140), .A2(n13119), .ZN(n11052) );
  OAI211_X1 U13978 ( .C1(n14444), .C2(n11054), .A(n11053), .B(n11052), .ZN(
        n15975) );
  AOI22_X1 U13979 ( .A1(n14442), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11066) );
  AOI22_X1 U13980 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14503), .B1(
        n10438), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11058) );
  AOI22_X1 U13981 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11057) );
  AOI22_X1 U13982 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11056) );
  AOI22_X1 U13983 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10528), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11055) );
  NAND4_X1 U13984 ( .A1(n11058), .A2(n11057), .A3(n11056), .A4(n11055), .ZN(
        n11064) );
  AOI22_X1 U13985 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10455), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11062) );
  AOI22_X1 U13986 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n13847), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11061) );
  AOI22_X1 U13987 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10472), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U13988 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14508), .ZN(n11059) );
  NAND4_X1 U13989 ( .A1(n11062), .A2(n11061), .A3(n11060), .A4(n11059), .ZN(
        n11063) );
  NOR2_X1 U13990 ( .A1(n11064), .A2(n11063), .ZN(n13120) );
  OR2_X1 U13991 ( .A1(n11140), .A2(n13120), .ZN(n11065) );
  OAI211_X1 U13992 ( .C1(n14444), .C2(n11067), .A(n11066), .B(n11065), .ZN(
        n16596) );
  NAND2_X1 U13993 ( .A1(n16595), .A2(n16596), .ZN(n13537) );
  AOI22_X1 U13994 ( .A1(n14442), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11082) );
  OAI22_X1 U13995 ( .A1(n11069), .A2(n11101), .B1(n11099), .B2(n11068), .ZN(
        n11070) );
  INV_X1 U13996 ( .A(n11070), .ZN(n11074) );
  AOI22_X1 U13997 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10528), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U13999 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U14000 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11080) );
  AOI22_X1 U14001 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14002 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14003 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14004 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14508), .ZN(n11075) );
  NAND4_X1 U14005 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11079) );
  INV_X1 U14006 ( .A(n13267), .ZN(n13189) );
  OR2_X1 U14007 ( .A1(n11140), .A2(n13189), .ZN(n11081) );
  OAI211_X1 U14008 ( .C1(n14444), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        n11084) );
  INV_X1 U14009 ( .A(n11084), .ZN(n13538) );
  AOI22_X1 U14010 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14011 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11087) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10528), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11086) );
  AOI22_X1 U14013 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10563), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11085) );
  NAND4_X1 U14014 ( .A1(n11088), .A2(n11087), .A3(n11086), .A4(n11085), .ZN(
        n11094) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10456), .B1(
        n10444), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U14016 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14017 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14018 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14508), .ZN(n11089) );
  NAND4_X1 U14019 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n11093) );
  OR2_X1 U14020 ( .A1(n11094), .A2(n11093), .ZN(n13193) );
  NAND2_X1 U14021 ( .A1(n11126), .A2(n13193), .ZN(n11096) );
  AOI22_X1 U14022 ( .A1(n14442), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11095) );
  OAI211_X1 U14023 ( .C1(n14444), .C2(n11097), .A(n11096), .B(n11095), .ZN(
        n16567) );
  NAND2_X1 U14024 ( .A1(n13536), .A2(n16567), .ZN(n13553) );
  AOI22_X1 U14025 ( .A1(n14442), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11114) );
  OAI22_X1 U14026 ( .A1(n11101), .A2(n11100), .B1(n11099), .B2(n11098), .ZN(
        n11102) );
  INV_X1 U14027 ( .A(n11102), .ZN(n11106) );
  AOI22_X1 U14028 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14029 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14030 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11103) );
  NAND4_X1 U14031 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11112) );
  AOI22_X1 U14032 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14033 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14034 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11108) );
  AOI22_X1 U14035 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14508), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11107) );
  NAND4_X1 U14036 ( .A1(n11110), .A2(n11109), .A3(n11108), .A4(n11107), .ZN(
        n11111) );
  INV_X1 U14037 ( .A(n13465), .ZN(n13463) );
  OR2_X1 U14038 ( .A1(n11140), .A2(n13463), .ZN(n11113) );
  OAI211_X1 U14039 ( .C1(n14444), .C2(n10891), .A(n11114), .B(n11113), .ZN(
        n11115) );
  INV_X1 U14040 ( .A(n11115), .ZN(n13555) );
  AOI22_X1 U14041 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14503), .B1(
        n10438), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14042 ( .A1(n10437), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14043 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10528), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11116) );
  NAND4_X1 U14045 ( .A1(n11119), .A2(n11118), .A3(n11117), .A4(n11116), .ZN(
        n11125) );
  AOI22_X1 U14046 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10456), .B1(
        n13847), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14047 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n13848), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14048 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11121) );
  AOI22_X1 U14049 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n13846), .ZN(n11120) );
  NAND4_X1 U14050 ( .A1(n11123), .A2(n11122), .A3(n11121), .A4(n11120), .ZN(
        n11124) );
  OR2_X1 U14051 ( .A1(n11125), .A2(n11124), .ZN(n13468) );
  NAND2_X1 U14052 ( .A1(n11126), .A2(n13468), .ZN(n11128) );
  AOI22_X1 U14053 ( .A1(n14442), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11127) );
  OAI211_X1 U14054 ( .C1(n14444), .C2(n11129), .A(n11128), .B(n11127), .ZN(
        n15956) );
  AOI22_X1 U14055 ( .A1(n14442), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11142) );
  AOI22_X1 U14056 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11133) );
  AOI22_X1 U14057 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14058 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10477), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14059 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10528), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11130) );
  NAND4_X1 U14060 ( .A1(n11133), .A2(n11132), .A3(n11131), .A4(n11130), .ZN(
        n11139) );
  AOI22_X1 U14061 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11137) );
  AOI22_X1 U14062 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11136) );
  AOI22_X1 U14063 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11135) );
  AOI22_X1 U14064 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n13846), .ZN(n11134) );
  NAND4_X1 U14065 ( .A1(n11137), .A2(n11136), .A3(n11135), .A4(n11134), .ZN(
        n11138) );
  NOR2_X1 U14066 ( .A1(n11139), .A2(n11138), .ZN(n13816) );
  OR2_X1 U14067 ( .A1(n11140), .A2(n13816), .ZN(n11141) );
  OAI211_X1 U14068 ( .C1(n14444), .C2(n20910), .A(n11142), .B(n11141), .ZN(
        n15938) );
  AOI22_X1 U14069 ( .A1(n14442), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11143) );
  OAI21_X1 U14070 ( .B1(n14444), .B2(n20808), .A(n11143), .ZN(n13712) );
  AOI22_X1 U14071 ( .A1(n14442), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11145) );
  OAI21_X1 U14072 ( .B1(n14444), .B2(n20097), .A(n11145), .ZN(n13864) );
  NAND2_X1 U14073 ( .A1(n11211), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11147) );
  AOI22_X1 U14074 ( .A1(n14442), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11146) );
  AND2_X1 U14075 ( .A1(n11147), .A2(n11146), .ZN(n13910) );
  NAND2_X1 U14076 ( .A1(n11211), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14077 ( .A1(n14442), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11148) );
  AND2_X1 U14078 ( .A1(n11149), .A2(n11148), .ZN(n13981) );
  AOI22_X1 U14079 ( .A1(n14442), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11150) );
  OAI21_X1 U14080 ( .B1(n14444), .B2(n20103), .A(n11150), .ZN(n14091) );
  NAND2_X1 U14081 ( .A1(n14092), .A2(n14091), .ZN(n14090) );
  NAND2_X1 U14082 ( .A1(n11211), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11152) );
  AOI22_X1 U14083 ( .A1(n14442), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11151) );
  AND2_X1 U14084 ( .A1(n11152), .A2(n11151), .ZN(n15444) );
  NOR2_X2 U14085 ( .A1(n14090), .A2(n15444), .ZN(n15430) );
  NAND2_X1 U14086 ( .A1(n11211), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11154) );
  AOI22_X1 U14087 ( .A1(n14442), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11153) );
  AND2_X1 U14088 ( .A1(n11154), .A2(n11153), .ZN(n15431) );
  AOI22_X1 U14089 ( .A1(n14442), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11156) );
  OAI21_X1 U14090 ( .B1(n14444), .B2(n11157), .A(n11156), .ZN(n15416) );
  AOI22_X1 U14091 ( .A1(n14442), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11158) );
  OAI21_X1 U14092 ( .B1(n14444), .B2(n20109), .A(n11158), .ZN(n15569) );
  NAND2_X1 U14093 ( .A1(n11211), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11160) );
  AOI22_X1 U14094 ( .A1(n14442), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11159) );
  AND2_X1 U14095 ( .A1(n11160), .A2(n11159), .ZN(n15401) );
  NAND2_X1 U14096 ( .A1(n11211), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11162) );
  AOI22_X1 U14097 ( .A1(n14442), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11161) );
  AND2_X1 U14098 ( .A1(n11162), .A2(n11161), .ZN(n15556) );
  AOI22_X1 U14099 ( .A1(n14442), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11163) );
  OAI21_X1 U14100 ( .B1(n14444), .B2(n15608), .A(n11163), .ZN(n15387) );
  NAND2_X1 U14101 ( .A1(n15558), .A2(n15387), .ZN(n11166) );
  NAND2_X1 U14102 ( .A1(n11211), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14103 ( .A1(n14442), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11164) );
  AND2_X1 U14104 ( .A1(n11165), .A2(n11164), .ZN(n11167) );
  NAND2_X1 U14105 ( .A1(n11166), .A2(n11167), .ZN(n11168) );
  AND2_X2 U14106 ( .A1(n9784), .A2(n11168), .ZN(n16433) );
  INV_X1 U14107 ( .A(n11169), .ZN(n12659) );
  INV_X1 U14108 ( .A(n11170), .ZN(n11171) );
  AND2_X1 U14109 ( .A1(n10940), .A2(n11171), .ZN(n16021) );
  INV_X1 U14110 ( .A(n16021), .ZN(n16660) );
  OAI21_X1 U14111 ( .B1(n9739), .B2(n12659), .A(n16660), .ZN(n11172) );
  NAND2_X1 U14112 ( .A1(n16433), .A2(n16621), .ZN(n11174) );
  OAI211_X1 U14113 ( .C1(n15787), .C2(n11175), .A(n14368), .B(n11174), .ZN(
        n11183) );
  NOR2_X1 U14114 ( .A1(n10329), .A2(n12819), .ZN(n11177) );
  NAND2_X1 U14115 ( .A1(n10329), .A2(n12819), .ZN(n11176) );
  OAI211_X1 U14116 ( .C1(n15924), .C2(n11177), .A(n11176), .B(n15952), .ZN(
        n16642) );
  NOR2_X1 U14117 ( .A1(n10522), .A2(n16642), .ZN(n16627) );
  NAND2_X1 U14118 ( .A1(n16627), .A2(n11178), .ZN(n15988) );
  NAND3_X1 U14119 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n11179) );
  NAND2_X1 U14120 ( .A1(n15892), .A2(n11181), .ZN(n16544) );
  NOR2_X1 U14121 ( .A1(n16544), .A2(n16543), .ZN(n15829) );
  NAND2_X1 U14122 ( .A1(n15829), .A2(n11182), .ZN(n15789) );
  NOR3_X1 U14123 ( .A1(n15789), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15810), .ZN(n15786) );
  AOI211_X1 U14124 ( .C1(n16434), .C2(n16635), .A(n11183), .B(n15786), .ZN(
        n11184) );
  OAI21_X1 U14125 ( .B1(n14373), .B2(n19500), .A(n10155), .ZN(P2_U3018) );
  AND2_X1 U14126 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15791) );
  AOI21_X1 U14127 ( .B1(n11190), .B2(n15791), .A(n11186), .ZN(n11192) );
  NAND2_X1 U14128 ( .A1(n15810), .A2(n11175), .ZN(n11189) );
  INV_X1 U14129 ( .A(n11187), .ZN(n11188) );
  OAI21_X1 U14130 ( .B1(n11190), .B2(n11189), .A(n11188), .ZN(n11191) );
  NAND2_X1 U14131 ( .A1(n11192), .A2(n11191), .ZN(n15595) );
  INV_X1 U14132 ( .A(n11193), .ZN(n11194) );
  NAND2_X1 U14133 ( .A1(n11197), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11196) );
  XNOR2_X1 U14134 ( .A(n11198), .B(n11196), .ZN(n15375) );
  INV_X1 U14135 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15790) );
  OAI21_X1 U14136 ( .B1(n15375), .B2(n11020), .A(n15790), .ZN(n15596) );
  NOR3_X1 U14137 ( .A1(n15375), .A2(n11020), .A3(n15790), .ZN(n15598) );
  AOI21_X1 U14138 ( .B1(n15595), .B2(n15596), .A(n15598), .ZN(n14421) );
  NAND2_X1 U14139 ( .A1(n11197), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11200) );
  INV_X1 U14140 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n15371) );
  OAI21_X1 U14141 ( .B1(n15371), .B2(n11199), .A(n11198), .ZN(n14422) );
  XOR2_X1 U14142 ( .A(n11200), .B(n14422), .Z(n16420) );
  NOR2_X1 U14143 ( .A1(n16420), .A2(n11020), .ZN(n11201) );
  NOR2_X1 U14144 ( .A1(n11201), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14420) );
  INV_X1 U14145 ( .A(n14420), .ZN(n11202) );
  NAND2_X1 U14146 ( .A1(n11201), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14419) );
  NAND2_X1 U14147 ( .A1(n11202), .A2(n14419), .ZN(n11203) );
  XNOR2_X1 U14148 ( .A(n14421), .B(n11203), .ZN(n15594) );
  NAND2_X1 U14149 ( .A1(n15791), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14456) );
  XOR2_X1 U14150 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n15600), .Z(
        n15592) );
  NOR3_X1 U14151 ( .A1(n15789), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14456), .ZN(n11204) );
  AOI22_X1 U14152 ( .A1(n9725), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n11207) );
  NAND2_X1 U14153 ( .A1(n11205), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11206) );
  OAI211_X1 U14154 ( .C1(n11210), .C2(n15790), .A(n11207), .B(n11206), .ZN(
        n15343) );
  INV_X1 U14155 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14457) );
  AOI22_X1 U14156 ( .A1(n9725), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n11209) );
  INV_X1 U14157 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20743) );
  OR2_X1 U14158 ( .A1(n14432), .A2(n20743), .ZN(n11208) );
  OAI211_X1 U14159 ( .C1(n11210), .C2(n14457), .A(n11209), .B(n11208), .ZN(
        n14428) );
  NAND2_X1 U14160 ( .A1(n11211), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14161 ( .A1(n14442), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11212) );
  AND2_X1 U14162 ( .A1(n11213), .A2(n11212), .ZN(n15370) );
  INV_X1 U14163 ( .A(n15370), .ZN(n11214) );
  AOI22_X1 U14164 ( .A1(n14442), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11216) );
  OAI21_X1 U14165 ( .B1(n14444), .B2(n20743), .A(n11216), .ZN(n14441) );
  INV_X1 U14166 ( .A(n14441), .ZN(n11217) );
  AOI21_X1 U14167 ( .B1(n15952), .B2(n14456), .A(n15806), .ZN(n14447) );
  NOR2_X1 U14168 ( .A1(n14447), .A2(n14457), .ZN(n11218) );
  NOR2_X1 U14169 ( .A1(n19304), .A2(n20743), .ZN(n15589) );
  OAI21_X1 U14170 ( .B1(n16422), .B2(n19491), .A(n11219), .ZN(n11220) );
  INV_X1 U14171 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11223) );
  INV_X1 U14172 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11224) );
  AND2_X2 U14173 ( .A1(n11230), .A2(n11234), .ZN(n11286) );
  AOI22_X1 U14174 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14175 ( .A1(n11552), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11455), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11227) );
  AOI22_X1 U14176 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11226) );
  AND2_X2 U14177 ( .A1(n13231), .A2(n11232), .ZN(n11297) );
  AOI22_X1 U14178 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11225) );
  AND2_X2 U14179 ( .A1(n11231), .A2(n11233), .ZN(n11394) );
  AND2_X2 U14180 ( .A1(n11231), .A2(n11230), .ZN(n11306) );
  AOI22_X1 U14181 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11238) );
  AND2_X2 U14182 ( .A1(n11231), .A2(n13231), .ZN(n12049) );
  AOI22_X1 U14183 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11237) );
  AND2_X2 U14184 ( .A1(n12903), .A2(n13231), .ZN(n11299) );
  AND2_X2 U14185 ( .A1(n11233), .A2(n11234), .ZN(n11298) );
  AOI22_X1 U14186 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11236) );
  AND2_X2 U14187 ( .A1(n11234), .A2(n13231), .ZN(n11701) );
  AOI22_X1 U14188 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14189 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14190 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14191 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11552), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14192 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14193 ( .A1(n11306), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11261), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14194 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11508), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14195 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11246) );
  AOI22_X1 U14196 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11245) );
  AOI22_X1 U14197 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11254) );
  AOI22_X1 U14198 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14199 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14200 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11251) );
  NAND4_X1 U14201 ( .A1(n11254), .A2(n11253), .A3(n11252), .A4(n11251), .ZN(
        n11260) );
  AOI22_X1 U14202 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11552), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14203 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11257) );
  AOI22_X1 U14204 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11256) );
  AOI22_X1 U14205 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11255) );
  NAND4_X1 U14206 ( .A1(n11258), .A2(n11257), .A3(n11256), .A4(n11255), .ZN(
        n11259) );
  NAND2_X1 U14207 ( .A1(n11306), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11265) );
  NAND2_X1 U14208 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11264) );
  NAND2_X1 U14209 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11263) );
  NAND2_X1 U14210 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11262) );
  NAND2_X1 U14211 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11269) );
  NAND2_X1 U14212 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11268) );
  NAND2_X1 U14213 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11267) );
  NAND2_X1 U14214 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11266) );
  NAND2_X1 U14215 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11273) );
  NAND2_X1 U14216 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11272) );
  NAND2_X1 U14217 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14218 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11270) );
  NAND2_X1 U14219 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14220 ( .A1(n11552), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11276) );
  NAND2_X1 U14221 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11275) );
  NAND2_X1 U14222 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11274) );
  NAND4_X4 U14223 ( .A1(n11281), .A2(n11280), .A3(n11279), .A4(n11278), .ZN(
        n11348) );
  AOI22_X1 U14224 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11552), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14225 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11284) );
  AOI22_X1 U14226 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11283) );
  AOI22_X1 U14227 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14228 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14229 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11289) );
  AOI22_X1 U14230 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14231 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11287) );
  NAND2_X2 U14232 ( .A1(n10172), .A2(n10169), .ZN(n11428) );
  AOI22_X1 U14233 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11296) );
  AOI22_X1 U14234 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14235 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11294) );
  AOI22_X1 U14236 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11293) );
  NAND4_X1 U14237 ( .A1(n11296), .A2(n11295), .A3(n11294), .A4(n11293), .ZN(
        n11305) );
  AOI22_X1 U14238 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11552), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14239 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14240 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11300) );
  NAND4_X1 U14241 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11304) );
  NAND2_X1 U14242 ( .A1(n11306), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11310) );
  NAND2_X1 U14243 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11309) );
  NAND2_X1 U14244 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11308) );
  NAND2_X1 U14245 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U14246 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11314) );
  NAND2_X1 U14247 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U14248 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11312) );
  NAND2_X1 U14249 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11311) );
  NAND2_X1 U14250 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11318) );
  NAND2_X1 U14251 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11317) );
  NAND2_X1 U14252 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11316) );
  NAND2_X1 U14253 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11315) );
  NAND2_X1 U14254 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U14255 ( .A1(n11552), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11321) );
  NAND2_X1 U14256 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11320) );
  NAND2_X1 U14257 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11319) );
  NAND4_X4 U14258 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n13472) );
  NAND2_X1 U14259 ( .A1(n11718), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11331) );
  NAND2_X1 U14260 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11330) );
  NAND2_X1 U14261 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11329) );
  NAND2_X1 U14262 ( .A1(n11286), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11328) );
  NAND2_X1 U14263 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14264 ( .A1(n11306), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11334) );
  NAND2_X1 U14265 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14266 ( .A1(n11386), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11332) );
  NAND2_X1 U14267 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11339) );
  NAND2_X1 U14268 ( .A1(n11508), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11338) );
  NAND2_X1 U14269 ( .A1(n11455), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11337) );
  NAND2_X1 U14270 ( .A1(n12489), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11336) );
  NAND2_X1 U14271 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11343) );
  NAND2_X1 U14272 ( .A1(n11552), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U14273 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11341) );
  NAND2_X1 U14274 ( .A1(n11701), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11340) );
  NAND4_X4 U14275 ( .A1(n11347), .A2(n11346), .A3(n11345), .A4(n11344), .ZN(
        n13479) );
  NAND2_X1 U14276 ( .A1(n12720), .A2(n13292), .ZN(n12517) );
  AND2_X2 U14277 ( .A1(n13034), .A2(n11428), .ZN(n11358) );
  NAND2_X1 U14278 ( .A1(n12786), .A2(n13472), .ZN(n12792) );
  INV_X1 U14279 ( .A(n12515), .ZN(n11350) );
  NAND2_X1 U14280 ( .A1(n11350), .A2(n13479), .ZN(n11351) );
  XNOR2_X1 U14281 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12769) );
  NAND2_X1 U14282 ( .A1(n13282), .A2(n13479), .ZN(n13481) );
  NAND2_X1 U14283 ( .A1(n11356), .A2(n13472), .ZN(n12777) );
  OAI211_X1 U14284 ( .C1(n13577), .C2(n20700), .A(n13052), .B(n11357), .ZN(
        n11375) );
  INV_X1 U14285 ( .A(n11428), .ZN(n13311) );
  NAND2_X1 U14286 ( .A1(n13311), .A2(n13472), .ZN(n13438) );
  NOR2_X1 U14287 ( .A1(n11375), .A2(n12779), .ZN(n11363) );
  OAI21_X1 U14288 ( .B1(n11348), .B2(n11360), .A(n9862), .ZN(n11361) );
  NAND2_X1 U14289 ( .A1(n13077), .A2(n11361), .ZN(n12782) );
  NAND2_X1 U14290 ( .A1(n12782), .A2(n15329), .ZN(n11362) );
  NAND3_X1 U14291 ( .A1(n11364), .A2(n11363), .A3(n11362), .ZN(n11365) );
  NAND2_X1 U14292 ( .A1(n15334), .A2(n10118), .ZN(n12136) );
  NAND2_X1 U14293 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11443) );
  OAI21_X1 U14294 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11443), .ZN(n13919) );
  NAND2_X1 U14295 ( .A1(n20614), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16183) );
  NAND2_X1 U14296 ( .A1(n16183), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11436) );
  OAI21_X1 U14297 ( .B1(n12136), .B2(n13919), .A(n11436), .ZN(n11366) );
  INV_X1 U14298 ( .A(n16183), .ZN(n11368) );
  MUX2_X1 U14299 ( .A(n11368), .B(n12136), .S(n20549), .Z(n11369) );
  INV_X1 U14300 ( .A(n12782), .ZN(n11379) );
  NAND2_X1 U14301 ( .A1(n15329), .A2(n13479), .ZN(n11378) );
  INV_X1 U14302 ( .A(n13495), .ZN(n12772) );
  NAND3_X1 U14303 ( .A1(n11359), .A2(n12772), .A3(n11428), .ZN(n11370) );
  NAND2_X1 U14304 ( .A1(n11355), .A2(n11370), .ZN(n11377) );
  NAND2_X1 U14305 ( .A1(n13135), .A2(n11371), .ZN(n13050) );
  NAND2_X1 U14306 ( .A1(n13297), .A2(n11360), .ZN(n11372) );
  INV_X1 U14307 ( .A(n20700), .ZN(n11582) );
  NAND2_X1 U14308 ( .A1(n11675), .A2(n11582), .ZN(n11373) );
  NAND4_X1 U14309 ( .A1(n13050), .A2(n11373), .A3(n15334), .A4(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n11374) );
  NOR2_X1 U14310 ( .A1(n11375), .A2(n11374), .ZN(n11376) );
  INV_X1 U14311 ( .A(n12612), .ZN(n11381) );
  INV_X1 U14312 ( .A(n11450), .ZN(n11468) );
  AOI22_X1 U14313 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14314 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11384) );
  AOI22_X1 U14315 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14316 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11382) );
  NAND4_X1 U14317 ( .A1(n11385), .A2(n11384), .A3(n11383), .A4(n11382), .ZN(
        n11392) );
  AOI22_X1 U14319 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11390) );
  AOI22_X1 U14320 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11389) );
  BUF_X1 U14321 ( .A(n11386), .Z(n11690) );
  AOI22_X1 U14322 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14323 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11387) );
  NAND4_X1 U14324 ( .A1(n11390), .A2(n11389), .A3(n11388), .A4(n11387), .ZN(
        n11391) );
  NAND2_X1 U14325 ( .A1(n11468), .A2(n11464), .ZN(n11393) );
  AOI22_X1 U14326 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11398) );
  BUF_X1 U14327 ( .A(n11394), .Z(n12048) );
  AOI22_X1 U14328 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12048), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14329 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n12057), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11396) );
  AOI22_X1 U14330 ( .A1(n12056), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11395) );
  NAND4_X1 U14331 ( .A1(n11398), .A2(n11397), .A3(n11396), .A4(n11395), .ZN(
        n11404) );
  AOI22_X1 U14332 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14333 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12051), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14334 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14335 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U14336 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11403) );
  OR2_X1 U14337 ( .A1(n11404), .A2(n11403), .ZN(n11429) );
  NAND2_X1 U14338 ( .A1(n11429), .A2(n11464), .ZN(n11497) );
  OAI21_X1 U14339 ( .B1(n11429), .B2(n11464), .A(n11497), .ZN(n11405) );
  OAI211_X1 U14340 ( .C1(n11405), .C2(n20700), .A(n11358), .B(n11352), .ZN(
        n11406) );
  INV_X1 U14341 ( .A(n11406), .ZN(n11407) );
  INV_X1 U14342 ( .A(n11408), .ZN(n11409) );
  INV_X1 U14343 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13836) );
  AOI21_X1 U14344 ( .B1(n13282), .B2(n11429), .A(n10118), .ZN(n11421) );
  AOI22_X1 U14345 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14346 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14347 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14348 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11411) );
  NAND4_X1 U14349 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11420) );
  AOI22_X1 U14350 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14351 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14352 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14353 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11415) );
  NAND4_X1 U14354 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11419) );
  NAND2_X1 U14355 ( .A1(n13577), .A2(n11581), .ZN(n11588) );
  OAI211_X1 U14356 ( .C1(n11662), .C2(n13836), .A(n11421), .B(n11588), .ZN(
        n11424) );
  INV_X1 U14357 ( .A(n11581), .ZN(n11590) );
  XNOR2_X1 U14358 ( .A(n11590), .B(n11429), .ZN(n11422) );
  NAND2_X1 U14359 ( .A1(n11422), .A2(n11468), .ZN(n11425) );
  AND2_X1 U14360 ( .A1(n11424), .A2(n11425), .ZN(n11423) );
  NAND2_X1 U14361 ( .A1(n11467), .A2(n11423), .ZN(n11427) );
  OR2_X1 U14362 ( .A1(n11425), .A2(n11424), .ZN(n11426) );
  NAND2_X1 U14363 ( .A1(n11352), .A2(n13479), .ZN(n11622) );
  INV_X1 U14364 ( .A(n11622), .ZN(n11577) );
  NAND2_X1 U14365 ( .A1(n13282), .A2(n11428), .ZN(n11470) );
  OAI21_X1 U14366 ( .B1(n20700), .B2(n11429), .A(n11470), .ZN(n11430) );
  INV_X1 U14367 ( .A(n11430), .ZN(n11431) );
  INV_X1 U14368 ( .A(n11432), .ZN(n13024) );
  NAND2_X1 U14369 ( .A1(n13024), .A2(n11433), .ZN(n11434) );
  INV_X1 U14370 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20962) );
  INV_X1 U14371 ( .A(n11435), .ZN(n11438) );
  NAND2_X1 U14372 ( .A1(n11436), .A2(n11223), .ZN(n11437) );
  NAND2_X1 U14373 ( .A1(n11438), .A2(n11437), .ZN(n11439) );
  INV_X1 U14374 ( .A(n12136), .ZN(n11481) );
  INV_X1 U14375 ( .A(n11443), .ZN(n11442) );
  NAND2_X1 U14376 ( .A1(n11442), .A2(n20788), .ZN(n13631) );
  NAND2_X1 U14377 ( .A1(n11443), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11444) );
  NAND2_X1 U14378 ( .A1(n13631), .A2(n11444), .ZN(n12619) );
  AOI22_X1 U14379 ( .A1(n11481), .A2(n12619), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16183), .ZN(n11445) );
  NAND2_X1 U14380 ( .A1(n11448), .A2(n12952), .ZN(n11449) );
  AOI22_X1 U14381 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14382 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11453) );
  AOI22_X1 U14383 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11452) );
  AOI22_X1 U14384 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11451) );
  NAND4_X1 U14385 ( .A1(n11454), .A2(n11453), .A3(n11452), .A4(n11451), .ZN(
        n11461) );
  AOI22_X1 U14386 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14387 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14388 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11457) );
  AOI22_X1 U14389 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11456) );
  NAND4_X1 U14390 ( .A1(n11459), .A2(n11458), .A3(n11457), .A4(n11456), .ZN(
        n11460) );
  OR2_X1 U14391 ( .A1(n11461), .A2(n11460), .ZN(n11469) );
  AOI22_X1 U14392 ( .A1(n11651), .A2(n11469), .B1(n11665), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11462) );
  INV_X1 U14393 ( .A(n11463), .ZN(n11465) );
  AOI22_X1 U14394 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11465), .B2(n11464), .ZN(n11466) );
  NAND2_X1 U14395 ( .A1(n9748), .A2(n11577), .ZN(n11474) );
  INV_X1 U14396 ( .A(n11469), .ZN(n11496) );
  XNOR2_X1 U14397 ( .A(n11497), .B(n11496), .ZN(n11472) );
  INV_X1 U14398 ( .A(n11470), .ZN(n11471) );
  AOI21_X1 U14399 ( .B1(n11472), .B2(n11582), .A(n11471), .ZN(n11473) );
  NAND2_X1 U14400 ( .A1(n11475), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11476) );
  INV_X1 U14401 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20380) );
  XNOR2_X1 U14402 ( .A(n11502), .B(n20380), .ZN(n13405) );
  NAND3_X1 U14403 ( .A1(n16172), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13921) );
  INV_X1 U14404 ( .A(n13921), .ZN(n13377) );
  NAND2_X1 U14405 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13377), .ZN(
        n13581) );
  NAND2_X1 U14406 ( .A1(n16172), .A2(n13581), .ZN(n11480) );
  NOR3_X1 U14407 ( .A1(n16172), .A2(n20788), .A3(n16166), .ZN(n14100) );
  NAND2_X1 U14408 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14100), .ZN(
        n13594) );
  AOI22_X1 U14409 ( .A1(n11481), .A2(n13826), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16183), .ZN(n11482) );
  AOI22_X1 U14410 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14411 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14412 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14413 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11483) );
  NAND4_X1 U14414 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11492) );
  AOI22_X1 U14415 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14416 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14417 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14418 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11487) );
  NAND4_X1 U14419 ( .A1(n11490), .A2(n11489), .A3(n11488), .A4(n11487), .ZN(
        n11491) );
  AOI22_X1 U14420 ( .A1(n11651), .A2(n11539), .B1(n11665), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U14421 ( .A1(n11523), .A2(n11495), .ZN(n11797) );
  OR2_X1 U14422 ( .A1(n11797), .A2(n11622), .ZN(n11501) );
  NAND2_X1 U14423 ( .A1(n11497), .A2(n11496), .ZN(n11541) );
  INV_X1 U14424 ( .A(n11539), .ZN(n11498) );
  XNOR2_X1 U14425 ( .A(n11541), .B(n11498), .ZN(n11499) );
  NAND2_X1 U14426 ( .A1(n11499), .A2(n11582), .ZN(n11500) );
  NAND2_X1 U14427 ( .A1(n11501), .A2(n11500), .ZN(n13404) );
  NAND2_X1 U14428 ( .A1(n11502), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11503) );
  AOI22_X1 U14429 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14430 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U14431 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14432 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U14433 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11514) );
  AOI22_X1 U14434 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14435 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14436 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14437 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14438 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  NAND2_X1 U14439 ( .A1(n11651), .A2(n11538), .ZN(n11516) );
  NAND2_X1 U14440 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11515) );
  NAND2_X1 U14441 ( .A1(n11516), .A2(n11515), .ZN(n11524) );
  XNOR2_X1 U14442 ( .A(n11523), .B(n11524), .ZN(n11813) );
  NAND2_X1 U14443 ( .A1(n11813), .A2(n11577), .ZN(n11520) );
  NAND2_X1 U14444 ( .A1(n11541), .A2(n11539), .ZN(n11517) );
  XNOR2_X1 U14445 ( .A(n11517), .B(n11538), .ZN(n11518) );
  NAND2_X1 U14446 ( .A1(n11518), .A2(n11582), .ZN(n11519) );
  NAND2_X1 U14447 ( .A1(n11520), .A2(n11519), .ZN(n11521) );
  INV_X1 U14448 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20963) );
  XNOR2_X1 U14449 ( .A(n11521), .B(n20963), .ZN(n20351) );
  NAND2_X1 U14450 ( .A1(n11521), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11522) );
  AOI22_X1 U14451 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14452 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11528) );
  AOI22_X1 U14453 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14454 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U14455 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11535) );
  AOI22_X1 U14456 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14457 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14458 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11531) );
  INV_X1 U14459 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20979) );
  AOI22_X1 U14460 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14461 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11534) );
  NAND2_X1 U14462 ( .A1(n11651), .A2(n11566), .ZN(n11537) );
  NAND2_X1 U14463 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U14464 ( .A1(n11537), .A2(n11536), .ZN(n11547) );
  NAND2_X1 U14465 ( .A1(n11814), .A2(n11577), .ZN(n11544) );
  AND2_X1 U14466 ( .A1(n11539), .A2(n11538), .ZN(n11540) );
  NAND2_X1 U14467 ( .A1(n11541), .A2(n11540), .ZN(n11565) );
  XNOR2_X1 U14468 ( .A(n11565), .B(n11566), .ZN(n11542) );
  NAND2_X1 U14469 ( .A1(n11542), .A2(n11582), .ZN(n11543) );
  NAND2_X1 U14470 ( .A1(n11544), .A2(n11543), .ZN(n11545) );
  INV_X1 U14471 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16388) );
  XNOR2_X1 U14472 ( .A(n11545), .B(n16388), .ZN(n16321) );
  NAND2_X1 U14473 ( .A1(n11545), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11546) );
  AOI22_X1 U14474 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14475 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14476 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14477 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14478 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11558) );
  AOI22_X1 U14479 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14480 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14481 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14482 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11553) );
  NAND4_X1 U14483 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n11557) );
  NAND2_X1 U14484 ( .A1(n11651), .A2(n11579), .ZN(n11560) );
  NAND2_X1 U14485 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11559) );
  NAND2_X1 U14486 ( .A1(n11564), .A2(n11563), .ZN(n11828) );
  NAND3_X1 U14487 ( .A1(n11576), .A2(n11828), .A3(n11577), .ZN(n11570) );
  INV_X1 U14488 ( .A(n11565), .ZN(n11567) );
  NAND2_X1 U14489 ( .A1(n11567), .A2(n11566), .ZN(n11578) );
  XNOR2_X1 U14490 ( .A(n11578), .B(n11579), .ZN(n11568) );
  NAND2_X1 U14491 ( .A1(n11568), .A2(n11582), .ZN(n11569) );
  NAND2_X1 U14492 ( .A1(n11570), .A2(n11569), .ZN(n13724) );
  OR2_X1 U14493 ( .A1(n13724), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11571) );
  NAND2_X1 U14494 ( .A1(n13724), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11572) );
  NAND2_X1 U14495 ( .A1(n11651), .A2(n11581), .ZN(n11574) );
  NAND2_X1 U14496 ( .A1(n11665), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14497 ( .A1(n11574), .A2(n11573), .ZN(n11575) );
  NAND2_X1 U14498 ( .A1(n11835), .A2(n11577), .ZN(n11585) );
  INV_X1 U14499 ( .A(n11578), .ZN(n11580) );
  NAND2_X1 U14500 ( .A1(n11580), .A2(n11579), .ZN(n11591) );
  XNOR2_X1 U14501 ( .A(n11591), .B(n11581), .ZN(n11583) );
  NAND2_X1 U14502 ( .A1(n11583), .A2(n11582), .ZN(n11584) );
  NAND2_X1 U14503 ( .A1(n11585), .A2(n11584), .ZN(n11586) );
  OR2_X1 U14504 ( .A1(n11586), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16316) );
  NAND2_X1 U14505 ( .A1(n11586), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16315) );
  NOR3_X1 U14506 ( .A1(n11588), .A2(n11622), .A3(n10118), .ZN(n11589) );
  NAND2_X4 U14507 ( .A1(n11576), .A2(n11589), .ZN(n11601) );
  OR3_X1 U14508 ( .A1(n11591), .A2(n11590), .A3(n20700), .ZN(n11592) );
  NAND2_X1 U14509 ( .A1(n11601), .A2(n11592), .ZN(n14006) );
  OR2_X1 U14510 ( .A1(n14006), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11593) );
  NAND2_X1 U14511 ( .A1(n14006), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11594) );
  INV_X1 U14512 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14053) );
  NAND2_X1 U14513 ( .A1(n11601), .A2(n14053), .ZN(n11595) );
  INV_X1 U14514 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15231) );
  NAND2_X1 U14515 ( .A1(n11601), .A2(n15231), .ZN(n11596) );
  NAND2_X1 U14516 ( .A1(n16298), .A2(n11596), .ZN(n15124) );
  INV_X1 U14517 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15313) );
  NAND2_X1 U14518 ( .A1(n11601), .A2(n15313), .ZN(n15122) );
  NAND2_X1 U14519 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11597) );
  NAND2_X1 U14520 ( .A1(n11601), .A2(n11597), .ZN(n15120) );
  NAND2_X1 U14521 ( .A1(n15122), .A2(n15120), .ZN(n11598) );
  NOR2_X1 U14522 ( .A1(n15124), .A2(n11598), .ZN(n16295) );
  INV_X1 U14523 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20883) );
  NAND2_X1 U14524 ( .A1(n11601), .A2(n20883), .ZN(n11599) );
  NAND2_X1 U14525 ( .A1(n16295), .A2(n11599), .ZN(n15108) );
  OR2_X1 U14526 ( .A1(n11601), .A2(n20883), .ZN(n11600) );
  NAND2_X1 U14527 ( .A1(n16298), .A2(n11600), .ZN(n15109) );
  INV_X1 U14528 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11602) );
  NAND2_X1 U14529 ( .A1(n15108), .A2(n11606), .ZN(n11604) );
  XNOR2_X1 U14530 ( .A(n11601), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15282) );
  NAND2_X1 U14531 ( .A1(n11601), .A2(n11602), .ZN(n15279) );
  AND2_X1 U14532 ( .A1(n15282), .A2(n15279), .ZN(n11603) );
  NAND2_X1 U14533 ( .A1(n11604), .A2(n11603), .ZN(n15096) );
  INV_X1 U14534 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n20797) );
  NAND2_X1 U14535 ( .A1(n11601), .A2(n20797), .ZN(n11605) );
  INV_X1 U14536 ( .A(n11606), .ZN(n11608) );
  NOR2_X1 U14537 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11607) );
  INV_X1 U14538 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15238) );
  OAI21_X2 U14539 ( .B1(n15061), .B2(n11609), .A(n11601), .ZN(n15053) );
  NAND2_X1 U14540 ( .A1(n15053), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14375) );
  INV_X1 U14541 ( .A(n15089), .ZN(n11611) );
  NOR2_X1 U14542 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11610) );
  AND2_X1 U14543 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U14544 ( .A1(n15188), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15186) );
  NOR2_X1 U14545 ( .A1(n9782), .A2(n15010), .ZN(n11613) );
  NAND2_X1 U14546 ( .A1(n9801), .A2(n11612), .ZN(n11614) );
  INV_X1 U14547 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15202) );
  INV_X1 U14548 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20816) );
  INV_X1 U14549 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15209) );
  NAND3_X1 U14550 ( .A1(n15202), .A2(n20816), .A3(n15209), .ZN(n14374) );
  XNOR2_X1 U14551 ( .A(n11615), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15177) );
  XNOR2_X1 U14552 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11630) );
  NAND2_X1 U14553 ( .A1(n11636), .A2(n11630), .ZN(n11617) );
  NAND2_X1 U14554 ( .A1(n16166), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11616) );
  NAND2_X1 U14555 ( .A1(n20788), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11621) );
  NAND2_X1 U14556 ( .A1(n12894), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11618) );
  NAND2_X1 U14557 ( .A1(n11621), .A2(n11618), .ZN(n11647) );
  INV_X1 U14558 ( .A(n11647), .ZN(n11619) );
  NAND2_X1 U14559 ( .A1(n11620), .A2(n11619), .ZN(n11649) );
  XNOR2_X1 U14560 ( .A(n11229), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11625) );
  AOI222_X1 U14561 ( .A1(n11660), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n11660), .B2(n20961), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n20961), .ZN(n12522) );
  NAND2_X1 U14562 ( .A1(n12522), .A2(n11659), .ZN(n11673) );
  NAND2_X1 U14563 ( .A1(n11651), .A2(n12522), .ZN(n11671) );
  AOI21_X1 U14564 ( .B1(n11625), .B2(n11624), .A(n11623), .ZN(n11626) );
  INV_X1 U14565 ( .A(n11626), .ZN(n12520) );
  NAND2_X1 U14566 ( .A1(n13297), .A2(n13472), .ZN(n11627) );
  NAND2_X1 U14567 ( .A1(n11627), .A2(n13292), .ZN(n11639) );
  INV_X1 U14568 ( .A(n11639), .ZN(n11655) );
  INV_X1 U14569 ( .A(n11651), .ZN(n11629) );
  NAND2_X1 U14570 ( .A1(n13297), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11631) );
  AND2_X1 U14571 ( .A1(n11631), .A2(n13479), .ZN(n11628) );
  NAND2_X1 U14572 ( .A1(n11629), .A2(n11628), .ZN(n11663) );
  XNOR2_X1 U14573 ( .A(n11630), .B(n11636), .ZN(n12518) );
  NAND2_X1 U14574 ( .A1(n11663), .A2(n12518), .ZN(n11634) );
  INV_X1 U14575 ( .A(n12518), .ZN(n11633) );
  NAND2_X1 U14576 ( .A1(n11651), .A2(n13479), .ZN(n11632) );
  OAI211_X1 U14577 ( .C1(n11633), .C2(n11662), .A(n11632), .B(n11631), .ZN(
        n11643) );
  NAND2_X1 U14578 ( .A1(n11634), .A2(n11643), .ZN(n11646) );
  AND2_X1 U14579 ( .A1(n11224), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11635) );
  NOR2_X1 U14580 ( .A1(n11636), .A2(n11635), .ZN(n11637) );
  AND2_X1 U14581 ( .A1(n11651), .A2(n11637), .ZN(n11642) );
  NAND2_X1 U14582 ( .A1(n11348), .A2(n11637), .ZN(n11638) );
  NAND2_X1 U14583 ( .A1(n11638), .A2(n13472), .ZN(n11640) );
  OAI21_X1 U14584 ( .B1(n13136), .B2(n11640), .A(n11639), .ZN(n11641) );
  OAI21_X1 U14585 ( .B1(n11659), .B2(n11642), .A(n11641), .ZN(n11645) );
  INV_X1 U14586 ( .A(n11643), .ZN(n11644) );
  AOI22_X1 U14587 ( .A1(n11646), .A2(n11645), .B1(n11644), .B2(n12518), .ZN(
        n11653) );
  NAND2_X1 U14588 ( .A1(n11648), .A2(n11647), .ZN(n11650) );
  NAND2_X1 U14589 ( .A1(n11650), .A2(n11649), .ZN(n12519) );
  INV_X1 U14590 ( .A(n12519), .ZN(n11652) );
  OAI211_X1 U14591 ( .C1(n11655), .C2(n11653), .A(n11652), .B(n11651), .ZN(
        n11657) );
  NOR2_X1 U14592 ( .A1(n11652), .A2(n11662), .ZN(n11654) );
  OAI21_X1 U14593 ( .B1(n11655), .B2(n11654), .A(n11653), .ZN(n11656) );
  AOI22_X1 U14594 ( .A1(n11662), .A2(n12520), .B1(n11657), .B2(n11656), .ZN(
        n11658) );
  AOI21_X1 U14595 ( .B1(n11659), .B2(n12520), .A(n11658), .ZN(n11668) );
  NAND2_X1 U14596 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11660), .ZN(
        n11661) );
  AND2_X1 U14597 ( .A1(n12521), .A2(n11662), .ZN(n11667) );
  INV_X1 U14598 ( .A(n11663), .ZN(n11664) );
  NAND3_X1 U14599 ( .A1(n11665), .A2(n11664), .A3(n12521), .ZN(n11666) );
  OAI21_X1 U14600 ( .B1(n11668), .B2(n11667), .A(n11666), .ZN(n11669) );
  AOI21_X1 U14601 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10118), .A(
        n11669), .ZN(n11670) );
  NAND2_X1 U14602 ( .A1(n11671), .A2(n11670), .ZN(n11672) );
  OR2_X1 U14603 ( .A1(n16183), .A2(n10118), .ZN(n20197) );
  AOI21_X1 U14604 ( .B1(n15329), .B2(n13282), .A(n11674), .ZN(n12516) );
  INV_X1 U14605 ( .A(n11675), .ZN(n11677) );
  OR2_X1 U14606 ( .A1(n11359), .A2(n11348), .ZN(n11676) );
  AND2_X1 U14607 ( .A1(n11677), .A2(n11676), .ZN(n12775) );
  AND2_X1 U14608 ( .A1(n12516), .A2(n12775), .ZN(n12882) );
  NAND2_X1 U14609 ( .A1(n12882), .A2(n11678), .ZN(n16175) );
  INV_X1 U14610 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16250) );
  INV_X1 U14611 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15102) );
  INV_X1 U14612 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14815) );
  INV_X1 U14613 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14787) );
  INV_X1 U14614 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14763) );
  AND2_X1 U14615 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11683) );
  INV_X1 U14616 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14748) );
  INV_X1 U14617 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14732) );
  OAI21_X1 U14618 ( .B1(n12127), .B2(n14748), .A(n14732), .ZN(n11685) );
  NAND2_X1 U14619 ( .A1(n12484), .A2(n11685), .ZN(n14731) );
  INV_X1 U14620 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U14621 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14622 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14623 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14624 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U14625 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11696) );
  AOI22_X1 U14626 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14627 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14628 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11692) );
  AOI22_X1 U14629 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11691) );
  NAND4_X1 U14630 ( .A1(n11694), .A2(n11693), .A3(n11692), .A4(n11691), .ZN(
        n11695) );
  NOR2_X1 U14631 ( .A1(n11696), .A2(n11695), .ZN(n12123) );
  AOI22_X1 U14632 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14633 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14634 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11698) );
  AOI22_X1 U14635 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11697) );
  NAND4_X1 U14636 ( .A1(n11700), .A2(n11699), .A3(n11698), .A4(n11697), .ZN(
        n11707) );
  AOI22_X1 U14637 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14638 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11298), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14639 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14640 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U14641 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  NOR2_X1 U14642 ( .A1(n11707), .A2(n11706), .ZN(n12107) );
  AOI22_X1 U14643 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14644 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14645 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11709) );
  AOI22_X1 U14646 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11708) );
  NAND4_X1 U14647 ( .A1(n11711), .A2(n11710), .A3(n11709), .A4(n11708), .ZN(
        n11717) );
  AOI22_X1 U14648 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11715) );
  AOI22_X1 U14649 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11714) );
  AOI22_X1 U14650 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11713) );
  AOI22_X1 U14651 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11712) );
  NAND4_X1 U14652 ( .A1(n11715), .A2(n11714), .A3(n11713), .A4(n11712), .ZN(
        n11716) );
  NOR2_X1 U14653 ( .A1(n11717), .A2(n11716), .ZN(n12092) );
  AOI22_X1 U14654 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11722) );
  AOI22_X1 U14655 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14656 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14657 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11719) );
  NAND4_X1 U14658 ( .A1(n11722), .A2(n11721), .A3(n11720), .A4(n11719), .ZN(
        n11728) );
  AOI22_X1 U14659 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n9730), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11726) );
  AOI22_X1 U14660 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14661 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n12494), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14662 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11723) );
  NAND4_X1 U14663 ( .A1(n11726), .A2(n11725), .A3(n11724), .A4(n11723), .ZN(
        n11727) );
  NOR2_X1 U14664 ( .A1(n11728), .A2(n11727), .ZN(n12093) );
  NOR2_X1 U14665 ( .A1(n12092), .A2(n12093), .ZN(n12102) );
  AOI22_X1 U14666 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11732) );
  AOI22_X1 U14667 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11731) );
  AOI22_X1 U14668 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11730) );
  AOI22_X1 U14669 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14670 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n11738) );
  AOI22_X1 U14671 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11736) );
  AOI22_X1 U14672 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11735) );
  INV_X1 U14673 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20725) );
  AOI22_X1 U14674 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11734) );
  AOI22_X1 U14675 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11733) );
  NAND4_X1 U14676 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11737) );
  OR2_X1 U14677 ( .A1(n11738), .A2(n11737), .ZN(n12101) );
  NAND2_X1 U14678 ( .A1(n12102), .A2(n12101), .ZN(n12108) );
  NOR2_X1 U14679 ( .A1(n12107), .A2(n12108), .ZN(n12118) );
  AOI22_X1 U14680 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11743) );
  AOI22_X1 U14681 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14682 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14683 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11740) );
  NAND4_X1 U14684 ( .A1(n11743), .A2(n11742), .A3(n11741), .A4(n11740), .ZN(
        n11749) );
  AOI22_X1 U14685 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14686 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U14687 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11745) );
  AOI22_X1 U14688 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11744) );
  NAND4_X1 U14689 ( .A1(n11747), .A2(n11746), .A3(n11745), .A4(n11744), .ZN(
        n11748) );
  OR2_X1 U14690 ( .A1(n11749), .A2(n11748), .ZN(n12117) );
  NAND2_X1 U14691 ( .A1(n12118), .A2(n12117), .ZN(n12124) );
  NOR2_X1 U14692 ( .A1(n12123), .A2(n12124), .ZN(n11761) );
  AOI22_X1 U14693 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U14694 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11752) );
  AOI22_X1 U14695 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U14696 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11750) );
  NAND4_X1 U14697 ( .A1(n11753), .A2(n11752), .A3(n11751), .A4(n11750), .ZN(
        n11759) );
  AOI22_X1 U14698 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14699 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11756) );
  AOI22_X1 U14700 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U14701 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11754) );
  NAND4_X1 U14702 ( .A1(n11757), .A2(n11756), .A3(n11755), .A4(n11754), .ZN(
        n11758) );
  OR2_X1 U14703 ( .A1(n11759), .A2(n11758), .ZN(n11760) );
  NAND2_X1 U14704 ( .A1(n11761), .A2(n11760), .ZN(n12502) );
  INV_X1 U14705 ( .A(n15329), .ZN(n14359) );
  OAI211_X1 U14706 ( .C1(n11761), .C2(n11760), .A(n12502), .B(n12482), .ZN(
        n11763) );
  INV_X1 U14707 ( .A(n13475), .ZN(n12506) );
  AOI21_X1 U14708 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20616), .A(
        n12506), .ZN(n11762) );
  OAI211_X1 U14709 ( .C1(n11821), .C2(n12969), .A(n11763), .B(n11762), .ZN(
        n11764) );
  NAND2_X1 U14710 ( .A1(n11765), .A2(n11955), .ZN(n11771) );
  NAND2_X1 U14711 ( .A1(n11353), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11803) );
  XNOR2_X1 U14712 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13565) );
  AOI21_X1 U14713 ( .B1(n12506), .B2(n13565), .A(n12512), .ZN(n11768) );
  INV_X1 U14714 ( .A(n11766), .ZN(n11821) );
  NAND2_X1 U14715 ( .A1(n12513), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11767) );
  OAI211_X1 U14716 ( .C1(n11803), .C2(n12894), .A(n11768), .B(n11767), .ZN(
        n11769) );
  INV_X1 U14717 ( .A(n11769), .ZN(n11770) );
  NAND2_X1 U14718 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  NAND2_X1 U14719 ( .A1(n12512), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11796) );
  NAND2_X1 U14720 ( .A1(n11772), .A2(n11796), .ZN(n13185) );
  INV_X1 U14721 ( .A(n11773), .ZN(n11775) );
  NAND2_X1 U14722 ( .A1(n11775), .A2(n11774), .ZN(n11781) );
  INV_X1 U14723 ( .A(n11776), .ZN(n11779) );
  INV_X1 U14724 ( .A(n11777), .ZN(n11778) );
  NAND2_X1 U14725 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  NAND2_X1 U14726 ( .A1(n12607), .A2(n11955), .ZN(n11785) );
  AOI22_X1 U14727 ( .A1(n12513), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20616), .ZN(n11783) );
  INV_X1 U14728 ( .A(n11803), .ZN(n11806) );
  NAND2_X1 U14729 ( .A1(n11806), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11782) );
  AND2_X1 U14730 ( .A1(n11783), .A2(n11782), .ZN(n11784) );
  NAND2_X1 U14731 ( .A1(n11785), .A2(n11784), .ZN(n13081) );
  OR2_X1 U14732 ( .A1(n13659), .A2(n11360), .ZN(n11786) );
  NAND2_X1 U14733 ( .A1(n11786), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U14734 ( .A1(n11787), .A2(n11955), .ZN(n11789) );
  AOI22_X1 U14735 ( .A1(n11806), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n12513), .B2(P1_EAX_REG_0__SCAN_IN), .ZN(n11788) );
  NAND2_X1 U14736 ( .A1(n11789), .A2(n11788), .ZN(n13075) );
  AND2_X1 U14737 ( .A1(n20616), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U14738 ( .A1(n13076), .A2(n11791), .ZN(n13074) );
  INV_X1 U14739 ( .A(n11791), .ZN(n11792) );
  NAND2_X1 U14740 ( .A1(n11792), .A2(n13475), .ZN(n11793) );
  NAND2_X1 U14741 ( .A1(n13081), .A2(n13080), .ZN(n13184) );
  INV_X1 U14742 ( .A(n13184), .ZN(n11794) );
  NAND2_X1 U14743 ( .A1(n11795), .A2(n11794), .ZN(n13182) );
  INV_X1 U14744 ( .A(n11798), .ZN(n11800) );
  INV_X1 U14745 ( .A(n11816), .ZN(n11799) );
  OAI21_X1 U14746 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11800), .A(
        n11799), .ZN(n14879) );
  AOI22_X1 U14747 ( .A1(n12506), .A2(n14879), .B1(n12512), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14748 ( .A1(n12513), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11801) );
  OAI211_X1 U14749 ( .C1(n11803), .C2(n11229), .A(n11802), .B(n11801), .ZN(
        n11804) );
  INV_X1 U14750 ( .A(n11804), .ZN(n11805) );
  NAND2_X1 U14751 ( .A1(n13145), .A2(n13144), .ZN(n13143) );
  NAND2_X1 U14752 ( .A1(n11806), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11811) );
  INV_X1 U14753 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11807) );
  AOI21_X1 U14754 ( .B1(n11807), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11808) );
  AOI21_X1 U14755 ( .B1(n12513), .B2(P1_EAX_REG_4__SCAN_IN), .A(n11808), .ZN(
        n11810) );
  XNOR2_X1 U14756 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B(n11816), .ZN(
        n20360) );
  NOR2_X1 U14757 ( .A1(n20360), .A2(n13475), .ZN(n11809) );
  AOI21_X1 U14758 ( .B1(n11811), .B2(n11810), .A(n11809), .ZN(n11812) );
  NOR2_X2 U14759 ( .A1(n13143), .A2(n13347), .ZN(n13354) );
  INV_X1 U14760 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13356) );
  NAND2_X1 U14761 ( .A1(n11814), .A2(n11955), .ZN(n11820) );
  INV_X1 U14762 ( .A(n11815), .ZN(n11823) );
  INV_X1 U14763 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20256) );
  NAND2_X1 U14764 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11816), .ZN(
        n11817) );
  NAND2_X1 U14765 ( .A1(n20256), .A2(n11817), .ZN(n11818) );
  NAND2_X1 U14766 ( .A1(n11823), .A2(n11818), .ZN(n20261) );
  AOI22_X1 U14767 ( .A1(n20261), .A2(n12506), .B1(n12512), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n11819) );
  OAI211_X1 U14768 ( .C1(n11821), .C2(n13356), .A(n11820), .B(n11819), .ZN(
        n13353) );
  NAND2_X1 U14769 ( .A1(n13354), .A2(n13353), .ZN(n13351) );
  INV_X1 U14770 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20307) );
  INV_X1 U14771 ( .A(n11831), .ZN(n11825) );
  INV_X1 U14772 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11822) );
  NAND2_X1 U14773 ( .A1(n11823), .A2(n11822), .ZN(n11824) );
  NAND2_X1 U14774 ( .A1(n11825), .A2(n11824), .ZN(n20248) );
  AOI22_X1 U14775 ( .A1(n20248), .A2(n12506), .B1(n12512), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11826) );
  OAI21_X1 U14776 ( .B1(n11821), .B2(n20307), .A(n11826), .ZN(n11827) );
  INV_X1 U14777 ( .A(n13437), .ZN(n11829) );
  NAND2_X1 U14778 ( .A1(n11830), .A2(n11829), .ZN(n13436) );
  INV_X1 U14779 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11833) );
  OAI21_X1 U14780 ( .B1(n11831), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11848), .ZN(n20237) );
  AOI22_X1 U14781 ( .A1(n20237), .A2(n12506), .B1(n12512), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11832) );
  OAI21_X1 U14782 ( .B1(n11821), .B2(n11833), .A(n11832), .ZN(n11834) );
  NAND2_X1 U14783 ( .A1(n11837), .A2(n11836), .ZN(n13612) );
  NAND2_X1 U14784 ( .A1(n12513), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U14785 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U14786 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12057), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11840) );
  AOI22_X1 U14787 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14788 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11838) );
  NAND4_X1 U14789 ( .A1(n11841), .A2(n11840), .A3(n11839), .A4(n11838), .ZN(
        n11847) );
  AOI22_X1 U14790 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n12032), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11845) );
  AOI22_X1 U14791 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n12051), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14792 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14793 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11842) );
  NAND4_X1 U14794 ( .A1(n11845), .A2(n11844), .A3(n11843), .A4(n11842), .ZN(
        n11846) );
  OAI21_X1 U14795 ( .B1(n11847), .B2(n11846), .A(n11955), .ZN(n11851) );
  INV_X1 U14796 ( .A(n11848), .ZN(n11849) );
  OAI21_X1 U14797 ( .B1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11849), .A(
        n11853), .ZN(n14009) );
  AOI22_X1 U14798 ( .A1(n12506), .A2(n14009), .B1(n12512), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11850) );
  NOR2_X2 U14799 ( .A1(n13612), .A2(n13788), .ZN(n13786) );
  AOI21_X1 U14800 ( .B1(n11853), .B2(n20969), .A(n11878), .ZN(n20220) );
  OR2_X1 U14801 ( .A1(n20220), .A2(n13475), .ZN(n11867) );
  AOI22_X1 U14802 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11857) );
  AOI22_X1 U14803 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14804 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14805 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11854) );
  NAND4_X1 U14806 ( .A1(n11857), .A2(n11856), .A3(n11855), .A4(n11854), .ZN(
        n11863) );
  AOI22_X1 U14807 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14808 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14809 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14810 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11858) );
  NAND4_X1 U14811 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11862) );
  NOR2_X1 U14812 ( .A1(n11863), .A2(n11862), .ZN(n11864) );
  INV_X1 U14813 ( .A(n12512), .ZN(n11992) );
  OAI22_X1 U14814 ( .A1(n11943), .A2(n11864), .B1(n11992), .B2(n20969), .ZN(
        n11865) );
  AOI21_X1 U14815 ( .B1(n12513), .B2(P1_EAX_REG_9__SCAN_IN), .A(n11865), .ZN(
        n11866) );
  NAND2_X1 U14816 ( .A1(n11867), .A2(n11866), .ZN(n13873) );
  AOI22_X1 U14817 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14818 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14819 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U14820 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11868) );
  NAND4_X1 U14821 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11877) );
  AOI22_X1 U14822 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11875) );
  AOI22_X1 U14823 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11874) );
  AOI22_X1 U14824 ( .A1(n12056), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14825 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11872) );
  NAND4_X1 U14826 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n11876) );
  NOR2_X1 U14827 ( .A1(n11877), .A2(n11876), .ZN(n11881) );
  XNOR2_X1 U14828 ( .A(n11878), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15142) );
  NAND2_X1 U14829 ( .A1(n15142), .A2(n12506), .ZN(n11880) );
  AOI22_X1 U14830 ( .A1(n12513), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12512), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11879) );
  OAI211_X1 U14831 ( .C1(n11881), .C2(n11943), .A(n11880), .B(n11879), .ZN(
        n13956) );
  INV_X1 U14832 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11885) );
  OAI21_X1 U14833 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11883), .A(
        n11882), .ZN(n16313) );
  NAND2_X1 U14834 ( .A1(n16313), .A2(n12506), .ZN(n11884) );
  OAI21_X1 U14835 ( .B1(n11885), .B2(n11992), .A(n11884), .ZN(n11886) );
  AOI21_X1 U14836 ( .B1(n12513), .B2(P1_EAX_REG_11__SCAN_IN), .A(n11886), .ZN(
        n14226) );
  AOI22_X1 U14837 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14838 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14839 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14840 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U14841 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11897) );
  AOI22_X1 U14842 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11895) );
  AOI22_X1 U14843 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11894) );
  AOI22_X1 U14844 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11893) );
  AOI22_X1 U14845 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11892) );
  NAND4_X1 U14846 ( .A1(n11895), .A2(n11894), .A3(n11893), .A4(n11892), .ZN(
        n11896) );
  OR2_X1 U14847 ( .A1(n11897), .A2(n11896), .ZN(n11898) );
  NAND2_X1 U14848 ( .A1(n11955), .A2(n11898), .ZN(n14254) );
  AOI22_X1 U14849 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14850 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14851 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11901) );
  AOI22_X1 U14852 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11900) );
  NAND4_X1 U14853 ( .A1(n11903), .A2(n11902), .A3(n11901), .A4(n11900), .ZN(
        n11909) );
  AOI22_X1 U14854 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14855 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14856 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11905) );
  AOI22_X1 U14857 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11904) );
  NAND4_X1 U14858 ( .A1(n11907), .A2(n11906), .A3(n11905), .A4(n11904), .ZN(
        n11908) );
  NOR2_X1 U14859 ( .A1(n11909), .A2(n11908), .ZN(n11915) );
  INV_X1 U14860 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14291) );
  OR2_X1 U14861 ( .A1(n11821), .A2(n14291), .ZN(n11914) );
  NOR2_X1 U14862 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n11910), .ZN(
        n11911) );
  NOR2_X1 U14863 ( .A1(n11926), .A2(n11911), .ZN(n16266) );
  INV_X1 U14864 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20960) );
  OAI22_X1 U14865 ( .A1(n16266), .A2(n13475), .B1(n11992), .B2(n20960), .ZN(
        n11912) );
  INV_X1 U14866 ( .A(n11912), .ZN(n11913) );
  OAI211_X1 U14867 ( .C1(n11915), .C2(n11943), .A(n11914), .B(n11913), .ZN(
        n14286) );
  AOI22_X1 U14868 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U14869 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U14870 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11917) );
  AOI22_X1 U14871 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11916) );
  NAND4_X1 U14872 ( .A1(n11919), .A2(n11918), .A3(n11917), .A4(n11916), .ZN(
        n11925) );
  AOI22_X1 U14873 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U14874 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U14875 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11921) );
  AOI22_X1 U14876 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11920) );
  NAND4_X1 U14877 ( .A1(n11923), .A2(n11922), .A3(n11921), .A4(n11920), .ZN(
        n11924) );
  NOR2_X1 U14878 ( .A1(n11925), .A2(n11924), .ZN(n11929) );
  INV_X1 U14879 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14280) );
  OR2_X1 U14880 ( .A1(n11821), .A2(n14280), .ZN(n11928) );
  XNOR2_X1 U14881 ( .A(n11926), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15125) );
  AOI22_X1 U14882 ( .A1(n15125), .A2(n12506), .B1(n12512), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11927) );
  OAI211_X1 U14883 ( .C1(n11929), .C2(n11943), .A(n11928), .B(n11927), .ZN(
        n14257) );
  XOR2_X1 U14884 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11930), .Z(
        n16302) );
  AOI22_X1 U14885 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U14886 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U14887 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U14888 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U14889 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11940) );
  AOI22_X1 U14890 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U14891 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U14892 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U14893 ( .A1(n12056), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U14894 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11939) );
  NOR2_X1 U14895 ( .A1(n11940), .A2(n11939), .ZN(n11942) );
  INV_X1 U14896 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11941) );
  OAI22_X1 U14897 ( .A1(n11943), .A2(n11942), .B1(n11992), .B2(n11941), .ZN(
        n11944) );
  AOI21_X1 U14898 ( .B1(n11766), .B2(P1_EAX_REG_14__SCAN_IN), .A(n11944), .ZN(
        n11945) );
  OAI21_X1 U14899 ( .B1(n16302), .B2(n13475), .A(n11945), .ZN(n14229) );
  XNOR2_X1 U14900 ( .A(n11946), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16255) );
  INV_X1 U14901 ( .A(n16255), .ZN(n11961) );
  AOI22_X1 U14902 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U14903 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U14904 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14905 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U14906 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11957) );
  AOI22_X1 U14907 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U14908 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14909 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14910 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U14911 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11956) );
  OAI21_X1 U14912 ( .B1(n11957), .B2(n11956), .A(n11955), .ZN(n11959) );
  NAND2_X1 U14913 ( .A1(n12513), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n11958) );
  OAI211_X1 U14914 ( .C1(n11992), .C2(n16250), .A(n11959), .B(n11958), .ZN(
        n11960) );
  AOI21_X1 U14915 ( .B1(n11961), .B2(n12506), .A(n11960), .ZN(n14270) );
  AOI22_X1 U14916 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U14917 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n12051), .B1(
        n12475), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U14918 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n12032), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U14919 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11963) );
  NAND4_X1 U14920 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n11972) );
  AOI22_X1 U14921 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11970) );
  AOI22_X1 U14922 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n12470), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11969) );
  AOI22_X1 U14923 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12494), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11968) );
  AOI22_X1 U14924 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11967) );
  NAND4_X1 U14925 ( .A1(n11970), .A2(n11969), .A3(n11968), .A4(n11967), .ZN(
        n11971) );
  NOR2_X1 U14926 ( .A1(n11972), .A2(n11971), .ZN(n11976) );
  NAND2_X1 U14927 ( .A1(n20616), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11973) );
  NAND2_X1 U14928 ( .A1(n13475), .A2(n11973), .ZN(n11974) );
  AOI21_X1 U14929 ( .B1(n11766), .B2(P1_EAX_REG_16__SCAN_IN), .A(n11974), .ZN(
        n11975) );
  OAI21_X1 U14930 ( .B1(n12509), .B2(n11976), .A(n11975), .ZN(n11979) );
  OAI21_X1 U14931 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11977), .A(
        n11991), .ZN(n16294) );
  OR2_X1 U14932 ( .A1(n13475), .A2(n16294), .ZN(n11978) );
  NAND2_X1 U14933 ( .A1(n11979), .A2(n11978), .ZN(n14931) );
  AOI22_X1 U14934 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U14935 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U14936 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U14937 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11980) );
  NAND4_X1 U14938 ( .A1(n11983), .A2(n11982), .A3(n11981), .A4(n11980), .ZN(
        n11989) );
  AOI22_X1 U14939 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U14940 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U14941 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U14942 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11984) );
  NAND4_X1 U14943 ( .A1(n11987), .A2(n11986), .A3(n11985), .A4(n11984), .ZN(
        n11988) );
  OR2_X1 U14944 ( .A1(n11989), .A2(n11988), .ZN(n11990) );
  NAND2_X1 U14945 ( .A1(n12482), .A2(n11990), .ZN(n11995) );
  XNOR2_X1 U14946 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11991), .ZN(
        n15104) );
  OAI22_X1 U14947 ( .A1(n13475), .A2(n15104), .B1(n11992), .B2(n15102), .ZN(
        n11993) );
  AOI21_X1 U14948 ( .B1(n11766), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11993), .ZN(
        n11994) );
  NAND2_X1 U14949 ( .A1(n11995), .A2(n11994), .ZN(n14859) );
  AOI22_X1 U14950 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U14951 ( .A1(n9743), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U14952 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U14953 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U14954 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12005) );
  AOI22_X1 U14955 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U14956 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U14957 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U14958 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12000) );
  NAND4_X1 U14959 ( .A1(n12003), .A2(n12002), .A3(n12001), .A4(n12000), .ZN(
        n12004) );
  NOR2_X1 U14960 ( .A1(n12005), .A2(n12004), .ZN(n12008) );
  INV_X1 U14961 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20998) );
  AOI21_X1 U14962 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n20998), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12006) );
  AOI21_X1 U14963 ( .B1(n11766), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12006), .ZN(
        n12007) );
  OAI21_X1 U14964 ( .B1(n12509), .B2(n12008), .A(n12007), .ZN(n12011) );
  NAND2_X1 U14965 ( .A1(n12029), .A2(n20998), .ZN(n12009) );
  NAND2_X1 U14966 ( .A1(n12074), .A2(n12009), .ZN(n15068) );
  OR2_X1 U14967 ( .A1(n15068), .A2(n13475), .ZN(n12010) );
  AOI22_X1 U14968 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12051), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U14969 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U14970 ( .A1(n12076), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U14971 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U14972 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12021) );
  AOI22_X1 U14973 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U14974 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U14975 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U14976 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U14977 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  NOR2_X1 U14978 ( .A1(n12021), .A2(n12020), .ZN(n12025) );
  NAND2_X1 U14979 ( .A1(n20616), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12022) );
  NAND2_X1 U14980 ( .A1(n13475), .A2(n12022), .ZN(n12023) );
  AOI21_X1 U14981 ( .B1(n11766), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12023), .ZN(
        n12024) );
  OAI21_X1 U14982 ( .B1(n12509), .B2(n12025), .A(n12024), .ZN(n12031) );
  INV_X1 U14983 ( .A(n12026), .ZN(n12027) );
  INV_X1 U14984 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15073) );
  NAND2_X1 U14985 ( .A1(n12027), .A2(n15073), .ZN(n12028) );
  AND2_X1 U14986 ( .A1(n12029), .A2(n12028), .ZN(n16222) );
  NAND2_X1 U14987 ( .A1(n16222), .A2(n12506), .ZN(n12030) );
  NAND2_X1 U14988 ( .A1(n12031), .A2(n12030), .ZN(n14917) );
  AOI22_X1 U14989 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U14990 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12032), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12035) );
  AOI22_X1 U14991 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U14992 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12033) );
  NAND4_X1 U14993 ( .A1(n12036), .A2(n12035), .A3(n12034), .A4(n12033), .ZN(
        n12042) );
  AOI22_X1 U14994 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12040) );
  AOI22_X1 U14995 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12039) );
  AOI22_X1 U14996 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U14997 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12037) );
  NAND4_X1 U14998 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        n12041) );
  NOR2_X1 U14999 ( .A1(n12042), .A2(n12041), .ZN(n12045) );
  INV_X1 U15000 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15083) );
  AOI21_X1 U15001 ( .B1(n15083), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12043) );
  AOI21_X1 U15002 ( .B1(n11766), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12043), .ZN(
        n12044) );
  OAI21_X1 U15003 ( .B1(n12509), .B2(n12045), .A(n12044), .ZN(n12047) );
  XNOR2_X1 U15004 ( .A(n12068), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15085) );
  NAND2_X1 U15005 ( .A1(n15085), .A2(n12506), .ZN(n12046) );
  NAND2_X1 U15006 ( .A1(n12047), .A2(n12046), .ZN(n14839) );
  NOR2_X1 U15007 ( .A1(n14917), .A2(n14839), .ZN(n14825) );
  AOI22_X1 U15008 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11739), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12055) );
  AOI22_X1 U15009 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15010 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12049), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15011 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12050), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12052) );
  NAND4_X1 U15012 ( .A1(n12055), .A2(n12054), .A3(n12053), .A4(n12052), .ZN(
        n12063) );
  AOI22_X1 U15013 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U15014 ( .A1(n12081), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U15015 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12059) );
  AOI22_X1 U15016 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12058) );
  NAND4_X1 U15017 ( .A1(n12061), .A2(n12060), .A3(n12059), .A4(n12058), .ZN(
        n12062) );
  NOR2_X1 U15018 ( .A1(n12063), .A2(n12062), .ZN(n12067) );
  NAND2_X1 U15019 ( .A1(n20616), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12064) );
  NAND2_X1 U15020 ( .A1(n13475), .A2(n12064), .ZN(n12065) );
  AOI21_X1 U15021 ( .B1(n11766), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12065), .ZN(
        n12066) );
  OAI21_X1 U15022 ( .B1(n12509), .B2(n12067), .A(n12066), .ZN(n12071) );
  OAI21_X1 U15023 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12069), .A(
        n12068), .ZN(n15092) );
  INV_X1 U15024 ( .A(n15092), .ZN(n16232) );
  NAND2_X1 U15025 ( .A1(n16232), .A2(n12506), .ZN(n12070) );
  NAND2_X1 U15026 ( .A1(n12074), .A2(n14815), .ZN(n12075) );
  NAND2_X1 U15027 ( .A1(n12096), .A2(n12075), .ZN(n15057) );
  INV_X1 U15028 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U15029 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15030 ( .A1(n12051), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15031 ( .A1(n9730), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12056), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12078) );
  AOI22_X1 U15032 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12077) );
  NAND4_X1 U15033 ( .A1(n12080), .A2(n12079), .A3(n12078), .A4(n12077), .ZN(
        n12087) );
  AOI22_X1 U15034 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12081), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15035 ( .A1(n9737), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15036 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15037 ( .A1(n12048), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12082) );
  NAND4_X1 U15038 ( .A1(n12085), .A2(n12084), .A3(n12083), .A4(n12082), .ZN(
        n12086) );
  OAI21_X1 U15039 ( .B1(n12087), .B2(n12086), .A(n12482), .ZN(n12089) );
  AOI21_X1 U15040 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20616), .A(
        n12506), .ZN(n12088) );
  OAI211_X1 U15041 ( .C1(n11821), .C2(n12090), .A(n12089), .B(n12088), .ZN(
        n12091) );
  OAI21_X1 U15042 ( .B1(n13475), .B2(n15057), .A(n12091), .ZN(n14809) );
  XOR2_X1 U15043 ( .A(n12093), .B(n12092), .Z(n12094) );
  NAND2_X1 U15044 ( .A1(n12482), .A2(n12094), .ZN(n12098) );
  INV_X1 U15045 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14800) );
  NOR2_X1 U15046 ( .A1(n14800), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12095) );
  AOI211_X1 U15047 ( .C1(n11766), .C2(P1_EAX_REG_23__SCAN_IN), .A(n12506), .B(
        n12095), .ZN(n12097) );
  XNOR2_X1 U15048 ( .A(n12096), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14799) );
  AOI22_X1 U15049 ( .A1(n12098), .A2(n12097), .B1(n12506), .B2(n14799), .ZN(
        n14798) );
  NAND2_X1 U15050 ( .A1(n12099), .A2(n14787), .ZN(n12100) );
  NAND2_X1 U15051 ( .A1(n12112), .A2(n12100), .ZN(n15041) );
  XNOR2_X1 U15052 ( .A(n12102), .B(n12101), .ZN(n12105) );
  INV_X1 U15053 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20818) );
  OAI21_X1 U15054 ( .B1(n20818), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n20616), .ZN(n12104) );
  NAND2_X1 U15055 ( .A1(n12513), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n12103) );
  OAI211_X1 U15056 ( .C1(n12105), .C2(n12509), .A(n12104), .B(n12103), .ZN(
        n12106) );
  OAI21_X1 U15057 ( .B1(n13475), .B2(n15041), .A(n12106), .ZN(n14783) );
  XOR2_X1 U15058 ( .A(n12108), .B(n12107), .Z(n12109) );
  NAND2_X1 U15059 ( .A1(n12109), .A2(n12482), .ZN(n12114) );
  INV_X1 U15060 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12110) );
  NOR2_X1 U15061 ( .A1(n12110), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12111) );
  AOI211_X1 U15062 ( .C1(n12513), .C2(P1_EAX_REG_25__SCAN_IN), .A(n12506), .B(
        n12111), .ZN(n12113) );
  XNOR2_X1 U15063 ( .A(n12112), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15030) );
  AOI22_X1 U15064 ( .A1(n12114), .A2(n12113), .B1(n12506), .B2(n15030), .ZN(
        n14775) );
  NAND2_X1 U15065 ( .A1(n12115), .A2(n14763), .ZN(n12116) );
  NAND2_X1 U15066 ( .A1(n12127), .A2(n12116), .ZN(n15022) );
  XNOR2_X1 U15067 ( .A(n12118), .B(n12117), .ZN(n12121) );
  AOI21_X1 U15068 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n20616), .A(
        n12506), .ZN(n12120) );
  NAND2_X1 U15069 ( .A1(n12513), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n12119) );
  OAI211_X1 U15070 ( .C1(n12121), .C2(n12509), .A(n12120), .B(n12119), .ZN(
        n12122) );
  XOR2_X1 U15071 ( .A(n12124), .B(n12123), .Z(n12125) );
  NAND2_X1 U15072 ( .A1(n12125), .A2(n12482), .ZN(n12129) );
  NOR2_X1 U15073 ( .A1(n14748), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12126) );
  AOI211_X1 U15074 ( .C1(n11766), .C2(P1_EAX_REG_27__SCAN_IN), .A(n12506), .B(
        n12126), .ZN(n12128) );
  XNOR2_X1 U15075 ( .A(n12127), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14747) );
  AOI22_X1 U15076 ( .A1(n12129), .A2(n12128), .B1(n12506), .B2(n14747), .ZN(
        n14742) );
  AOI21_X1 U15077 ( .B1(n12131), .B2(n12130), .A(n12488), .ZN(n14728) );
  NAND3_X1 U15078 ( .A1(n10118), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16395) );
  INV_X1 U15079 ( .A(n16395), .ZN(n12132) );
  NOR2_X1 U15080 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n13917) );
  AND2_X1 U15081 ( .A1(n12132), .A2(n13917), .ZN(n14067) );
  INV_X1 U15082 ( .A(n13917), .ZN(n20559) );
  NAND2_X1 U15083 ( .A1(n20559), .A2(n12136), .ZN(n20694) );
  NAND2_X1 U15084 ( .A1(n20694), .A2(n10118), .ZN(n12133) );
  NAND2_X1 U15085 ( .A1(n10118), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U15086 ( .A1(n20818), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12134) );
  AND2_X1 U15087 ( .A1(n12135), .A2(n12134), .ZN(n13085) );
  OR2_X2 U15088 ( .A1(n20350), .A2(n13085), .ZN(n20361) );
  OR2_X2 U15089 ( .A1(n12136), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20254) );
  INV_X1 U15090 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14736) );
  NOR2_X1 U15091 ( .A1(n20254), .A2(n14736), .ZN(n15173) );
  AOI21_X1 U15092 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15173), .ZN(n12137) );
  OAI21_X1 U15093 ( .B1(n20361), .B2(n14731), .A(n12137), .ZN(n12138) );
  AOI21_X1 U15094 ( .B1(n14728), .B2(n14067), .A(n12138), .ZN(n12139) );
  OAI21_X1 U15095 ( .B1(n15177), .B2(n20203), .A(n12139), .ZN(P1_U2971) );
  NAND2_X1 U15096 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12441) );
  NAND2_X1 U15097 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n18179) );
  NOR2_X1 U15098 ( .A1(n12441), .A2(n18179), .ZN(n12454) );
  INV_X1 U15099 ( .A(n12454), .ZN(n12577) );
  NAND2_X1 U15100 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18220) );
  INV_X1 U15101 ( .A(n18220), .ZN(n18235) );
  NAND3_X1 U15102 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18235), .ZN(n17888) );
  INV_X2 U15103 ( .A(n9786), .ZN(n17472) );
  INV_X4 U15104 ( .A(n9776), .ZN(n17480) );
  AOI22_X1 U15105 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n17472), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15106 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12154) );
  BUF_X2 U15107 ( .A(n12315), .Z(n17227) );
  INV_X1 U15108 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20854) );
  AOI22_X1 U15109 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12141) );
  OAI21_X1 U15110 ( .B1(n20854), .B2(n9778), .A(n12141), .ZN(n12152) );
  AOI22_X1 U15111 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12150) );
  NOR2_X2 U15112 ( .A1(n12146), .A2(n12143), .ZN(n12188) );
  AOI22_X1 U15113 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15114 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15115 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12147) );
  NAND4_X1 U15116 ( .A1(n12150), .A2(n12149), .A3(n12148), .A4(n12147), .ZN(
        n12151) );
  AOI211_X1 U15117 ( .C1(n17227), .C2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A(
        n12152), .B(n12151), .ZN(n12153) );
  NAND3_X1 U15118 ( .A1(n12155), .A2(n12154), .A3(n12153), .ZN(n12386) );
  INV_X1 U15119 ( .A(n12386), .ZN(n17652) );
  AOI22_X1 U15120 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12166) );
  INV_X2 U15121 ( .A(n9786), .ZN(n17453) );
  AOI22_X1 U15122 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12165) );
  INV_X1 U15123 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U15124 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12157) );
  OAI21_X1 U15125 ( .B1(n9777), .B2(n17507), .A(n12157), .ZN(n12163) );
  AOI22_X1 U15126 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12161) );
  INV_X2 U15127 ( .A(n10166), .ZN(n17474) );
  AOI22_X1 U15128 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15129 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12159) );
  INV_X2 U15130 ( .A(n9778), .ZN(n16122) );
  AOI22_X1 U15131 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12158) );
  NAND4_X1 U15132 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12162) );
  AOI211_X1 U15133 ( .C1(n12316), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n12163), .B(n12162), .ZN(n12164) );
  NAND3_X1 U15134 ( .A1(n12166), .A2(n12165), .A3(n12164), .ZN(n12376) );
  AOI22_X1 U15135 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15136 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12176) );
  INV_X1 U15137 ( .A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U15138 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12189), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12167) );
  OAI21_X1 U15139 ( .B1(n20936), .B2(n10166), .A(n12167), .ZN(n12174) );
  INV_X4 U15140 ( .A(n17267), .ZN(n16109) );
  AOI22_X1 U15141 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15142 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12171) );
  INV_X2 U15143 ( .A(n12253), .ZN(n16120) );
  AOI22_X1 U15144 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12168), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12170) );
  AOI22_X1 U15145 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12169) );
  NAND4_X1 U15146 ( .A1(n12172), .A2(n12171), .A3(n12170), .A4(n12169), .ZN(
        n12173) );
  AOI211_X1 U15147 ( .C1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .C2(n9729), .A(
        n12174), .B(n12173), .ZN(n12175) );
  NAND3_X1 U15148 ( .A1(n12177), .A2(n12176), .A3(n12175), .ZN(n12368) );
  AOI22_X1 U15149 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12168), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15150 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15151 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15152 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12178) );
  NAND4_X1 U15153 ( .A1(n12181), .A2(n12180), .A3(n12179), .A4(n12178), .ZN(
        n12187) );
  AOI22_X1 U15154 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15155 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12184) );
  AOI22_X1 U15156 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n12189), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12183) );
  AOI22_X1 U15157 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12182) );
  NAND4_X1 U15158 ( .A1(n12185), .A2(n12184), .A3(n12183), .A4(n12182), .ZN(
        n12186) );
  AOI22_X1 U15159 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17454), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17409), .ZN(n12198) );
  AOI22_X1 U15160 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17355), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12197) );
  INV_X1 U15161 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n20821) );
  AOI22_X1 U15162 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n12189), .ZN(n12190) );
  OAI21_X1 U15163 ( .B1(n20821), .B2(n10151), .A(n12190), .ZN(n12196) );
  AOI22_X1 U15164 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n16109), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15165 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12168), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17461), .ZN(n12194) );
  AOI22_X1 U15166 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15167 ( .A1(n12315), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15168 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12202) );
  AOI22_X1 U15169 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n17461), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12201) );
  AOI22_X1 U15170 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17311), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15171 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12199) );
  NAND4_X1 U15172 ( .A1(n12202), .A2(n12201), .A3(n12200), .A4(n12199), .ZN(
        n12208) );
  AOI22_X1 U15173 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15174 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15175 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15176 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12203) );
  NAND4_X1 U15177 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(
        n12207) );
  NAND2_X1 U15178 ( .A1(n12229), .A2(n12373), .ZN(n12237) );
  AOI22_X1 U15179 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15180 ( .A1(n16109), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15181 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15182 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n17355), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15183 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12218) );
  AOI22_X1 U15184 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15185 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15186 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15187 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12213) );
  NAND4_X1 U15188 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12217) );
  INV_X1 U15189 ( .A(n17655), .ZN(n12378) );
  NAND2_X1 U15190 ( .A1(n12239), .A2(n12378), .ZN(n12241) );
  NOR2_X1 U15191 ( .A1(n17652), .A2(n12241), .ZN(n12245) );
  AOI22_X1 U15192 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15193 ( .A1(n12189), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15194 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15195 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n17473), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12219) );
  NAND4_X1 U15196 ( .A1(n12222), .A2(n12221), .A3(n12220), .A4(n12219), .ZN(
        n12228) );
  AOI22_X1 U15197 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15198 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15199 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15200 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12223) );
  NAND4_X1 U15201 ( .A1(n12226), .A2(n12225), .A3(n12224), .A4(n12223), .ZN(
        n12227) );
  INV_X1 U15202 ( .A(n17648), .ZN(n12557) );
  NAND2_X1 U15203 ( .A1(n12245), .A2(n12557), .ZN(n12246) );
  XNOR2_X1 U15204 ( .A(n12229), .B(n12373), .ZN(n12235) );
  INV_X1 U15205 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n12392) );
  XNOR2_X1 U15206 ( .A(n12230), .B(n17665), .ZN(n12231) );
  INV_X1 U15207 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18436) );
  NOR2_X1 U15208 ( .A1(n12231), .A2(n18436), .ZN(n12234) );
  XOR2_X1 U15209 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12231), .Z(
        n18142) );
  INV_X1 U15210 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19106) );
  NOR2_X1 U15211 ( .A1(n12367), .A2(n19106), .ZN(n12233) );
  NAND3_X1 U15212 ( .A1(n18161), .A2(n12367), .A3(n19106), .ZN(n12232) );
  OAI221_X1 U15213 ( .B1(n12233), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18161), .C2(n12367), .A(n12232), .ZN(n18141) );
  NOR2_X1 U15214 ( .A1(n18142), .A2(n18141), .ZN(n18140) );
  NOR2_X1 U15215 ( .A1(n12234), .A2(n18140), .ZN(n18134) );
  XOR2_X1 U15216 ( .A(n12235), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18133) );
  INV_X1 U15217 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18417) );
  NOR2_X1 U15218 ( .A1(n12236), .A2(n18417), .ZN(n12238) );
  XOR2_X1 U15219 ( .A(n12376), .B(n12237), .Z(n18116) );
  XOR2_X1 U15220 ( .A(n12239), .B(n17655), .Z(n18105) );
  XOR2_X1 U15221 ( .A(n12386), .B(n12241), .Z(n12243) );
  NOR2_X1 U15222 ( .A1(n12242), .A2(n12243), .ZN(n12244) );
  INV_X1 U15223 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18386) );
  NOR2_X1 U15224 ( .A1(n18386), .A2(n18094), .ZN(n18093) );
  NOR2_X1 U15225 ( .A1(n12244), .A2(n18093), .ZN(n12247) );
  XOR2_X1 U15226 ( .A(n12245), .B(n17648), .Z(n12248) );
  NAND2_X1 U15227 ( .A1(n12247), .A2(n12248), .ZN(n18084) );
  NAND2_X1 U15228 ( .A1(n18084), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12250) );
  INV_X1 U15229 ( .A(n12246), .ZN(n12251) );
  OR2_X1 U15230 ( .A1(n12248), .A2(n12247), .ZN(n18085) );
  OAI21_X1 U15231 ( .B1(n12251), .B2(n12250), .A(n18085), .ZN(n12249) );
  AOI21_X1 U15232 ( .B1(n12251), .B2(n12250), .A(n12249), .ZN(n18074) );
  INV_X1 U15233 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n20850) );
  NOR2_X1 U15234 ( .A1(n12252), .A2(n18073), .ZN(n18340) );
  AOI22_X1 U15235 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15236 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15237 ( .A1(n16109), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15238 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n16120), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12254) );
  NAND4_X1 U15239 ( .A1(n12257), .A2(n12256), .A3(n12255), .A4(n12254), .ZN(
        n12263) );
  AOI22_X1 U15240 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15241 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17481), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15242 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15243 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15244 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  AOI22_X1 U15245 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15246 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15247 ( .A1(n17473), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12264) );
  OAI21_X1 U15248 ( .B1(n20937), .B2(n9786), .A(n12264), .ZN(n12271) );
  AOI22_X1 U15249 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12168), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15250 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15251 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15252 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12266) );
  NAND4_X1 U15253 ( .A1(n12269), .A2(n12268), .A3(n12267), .A4(n12266), .ZN(
        n12270) );
  AOI211_X1 U15254 ( .C1(n9729), .C2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A(
        n12271), .B(n12270), .ZN(n12272) );
  NAND3_X1 U15255 ( .A1(n12274), .A2(n12273), .A3(n12272), .ZN(n16211) );
  NAND2_X1 U15256 ( .A1(n18485), .A2(n17729), .ZN(n12346) );
  AOI22_X1 U15257 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15258 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15259 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15260 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12275) );
  NAND4_X1 U15261 ( .A1(n12278), .A2(n12277), .A3(n12276), .A4(n12275), .ZN(
        n12284) );
  AOI22_X1 U15262 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15263 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15264 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15265 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12279) );
  NAND4_X1 U15266 ( .A1(n12282), .A2(n12281), .A3(n12280), .A4(n12279), .ZN(
        n12283) );
  AOI22_X1 U15267 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12294) );
  AOI22_X1 U15268 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12293) );
  INV_X1 U15269 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n20726) );
  AOI22_X1 U15270 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12285) );
  OAI21_X1 U15271 ( .B1(n20726), .B2(n17267), .A(n12285), .ZN(n12291) );
  AOI22_X1 U15272 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15273 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15274 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12287) );
  AOI22_X1 U15275 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12286) );
  NAND4_X1 U15276 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n12286), .ZN(
        n12290) );
  AOI211_X1 U15277 ( .C1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n17454), .A(
        n12291), .B(n12290), .ZN(n12292) );
  NAND3_X1 U15278 ( .A1(n12294), .A2(n12293), .A3(n12292), .ZN(n12343) );
  NAND2_X1 U15279 ( .A1(n16052), .A2(n18510), .ZN(n18920) );
  AOI22_X1 U15280 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15281 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12303) );
  INV_X1 U15282 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20789) );
  AOI22_X1 U15283 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12295) );
  OAI21_X1 U15284 ( .B1(n20789), .B2(n10151), .A(n12295), .ZN(n12301) );
  AOI22_X1 U15285 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15286 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15287 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12168), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15288 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15289 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12300) );
  AOI211_X2 U15290 ( .C1(n17460), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n12301), .B(n12300), .ZN(n12302) );
  NAND3_X2 U15291 ( .A1(n12304), .A2(n12303), .A3(n12302), .ZN(n17533) );
  NOR2_X2 U15292 ( .A1(n18510), .A2(n17533), .ZN(n12366) );
  INV_X1 U15293 ( .A(n12366), .ZN(n12337) );
  AOI22_X1 U15294 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15295 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12313) );
  INV_X1 U15296 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n20777) );
  AOI22_X1 U15297 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12305) );
  OAI21_X1 U15298 ( .B1(n20777), .B2(n10152), .A(n12305), .ZN(n12311) );
  AOI22_X1 U15299 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15300 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15301 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n17355), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12307) );
  AOI22_X1 U15302 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12306) );
  NAND4_X1 U15303 ( .A1(n12309), .A2(n12308), .A3(n12307), .A4(n12306), .ZN(
        n12310) );
  AOI211_X1 U15304 ( .C1(n12316), .C2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A(
        n12311), .B(n12310), .ZN(n12312) );
  NAND3_X1 U15305 ( .A1(n12314), .A2(n12313), .A3(n12312), .ZN(n12340) );
  NAND3_X1 U15306 ( .A1(n18920), .A2(n12337), .A3(n18491), .ZN(n12351) );
  NAND2_X1 U15307 ( .A1(n17533), .A2(n18491), .ZN(n12425) );
  NAND2_X1 U15308 ( .A1(n12351), .A2(n12425), .ZN(n12353) );
  AOI22_X1 U15309 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12326) );
  INV_X2 U15310 ( .A(n12156), .ZN(n17460) );
  AOI22_X1 U15311 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12325) );
  INV_X1 U15312 ( .A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n20718) );
  AOI22_X1 U15313 ( .A1(n16122), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12168), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12317) );
  OAI21_X1 U15314 ( .B1(n20718), .B2(n9777), .A(n12317), .ZN(n12324) );
  AOI22_X1 U15315 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15316 ( .A1(n12189), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U15317 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12320) );
  AOI22_X1 U15318 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12319) );
  NAND4_X1 U15319 ( .A1(n12322), .A2(n12321), .A3(n12320), .A4(n12319), .ZN(
        n12323) );
  AOI22_X1 U15320 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U15321 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12335) );
  INV_X1 U15322 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20836) );
  AOI22_X1 U15323 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12327) );
  OAI21_X1 U15324 ( .B1(n20836), .B2(n9776), .A(n12327), .ZN(n12333) );
  AOI22_X1 U15325 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15326 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17227), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15327 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9724), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15328 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12328) );
  NAND4_X1 U15329 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12328), .ZN(
        n12332) );
  AOI211_X1 U15330 ( .C1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .C2(n9722), .A(
        n12333), .B(n12332), .ZN(n12334) );
  NAND3_X1 U15331 ( .A1(n12336), .A2(n12335), .A3(n12334), .ZN(n12339) );
  NOR2_X2 U15332 ( .A1(n19145), .A2(n16054), .ZN(n18963) );
  NAND2_X1 U15333 ( .A1(n18491), .A2(n18496), .ZN(n18919) );
  NOR2_X1 U15334 ( .A1(n12345), .A2(n16053), .ZN(n12342) );
  AND2_X2 U15335 ( .A1(n17725), .A2(n16211), .ZN(n12341) );
  NAND2_X1 U15336 ( .A1(n12343), .A2(n17533), .ZN(n12348) );
  NOR4_X2 U15337 ( .A1(n16052), .A2(n12339), .A3(n12345), .A4(n12348), .ZN(
        n12355) );
  NOR2_X2 U15338 ( .A1(n12341), .A2(n12417), .ZN(n16818) );
  INV_X2 U15339 ( .A(n12632), .ZN(n17678) );
  XNOR2_X1 U15340 ( .A(n17729), .B(n18491), .ZN(n12422) );
  INV_X1 U15341 ( .A(n17533), .ZN(n18506) );
  NOR2_X1 U15342 ( .A1(n18506), .A2(n12343), .ZN(n18929) );
  NOR2_X1 U15343 ( .A1(n18516), .A2(n18929), .ZN(n16216) );
  AOI22_X1 U15344 ( .A1(n18501), .A2(n18929), .B1(n18496), .B2(n12345), .ZN(
        n12350) );
  NAND2_X1 U15345 ( .A1(n18491), .A2(n12346), .ZN(n12362) );
  AOI21_X1 U15346 ( .B1(n17647), .B2(n12348), .A(n18501), .ZN(n12347) );
  AOI21_X1 U15347 ( .B1(n12348), .B2(n12362), .A(n12347), .ZN(n12349) );
  OAI211_X1 U15348 ( .C1(n16211), .C2(n12351), .A(n12350), .B(n12349), .ZN(
        n12352) );
  INV_X1 U15349 ( .A(n12352), .ZN(n12415) );
  OAI211_X1 U15350 ( .C1(n12353), .C2(n18496), .A(n12414), .B(n12415), .ZN(
        n12358) );
  INV_X1 U15351 ( .A(n12358), .ZN(n12354) );
  NAND2_X1 U15352 ( .A1(n12355), .A2(n12354), .ZN(n18923) );
  NOR2_X1 U15353 ( .A1(n19132), .A2(n12364), .ZN(n12360) );
  INV_X1 U15354 ( .A(n12357), .ZN(n12359) );
  NAND2_X1 U15355 ( .A1(n18491), .A2(n17729), .ZN(n12361) );
  NOR2_X1 U15356 ( .A1(n18510), .A2(n12361), .ZN(n12427) );
  INV_X1 U15357 ( .A(n12362), .ZN(n12363) );
  OAI211_X1 U15358 ( .C1(n18501), .C2(n18929), .A(n12364), .B(n12363), .ZN(
        n12365) );
  NOR2_X1 U15359 ( .A1(n12366), .A2(n12365), .ZN(n12416) );
  NAND2_X1 U15360 ( .A1(n12427), .A2(n12416), .ZN(n18956) );
  NOR2_X1 U15361 ( .A1(n12557), .A2(n18956), .ZN(n18339) );
  XOR2_X1 U15362 ( .A(n12373), .B(n12372), .Z(n18129) );
  XNOR2_X1 U15363 ( .A(n12368), .B(n12367), .ZN(n12370) );
  NAND2_X1 U15364 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12370), .ZN(
        n12371) );
  NAND2_X1 U15365 ( .A1(n12367), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12369) );
  INV_X1 U15366 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19090) );
  NOR2_X1 U15367 ( .A1(n18161), .A2(n19106), .ZN(n18160) );
  NAND2_X1 U15368 ( .A1(n12369), .A2(n18151), .ZN(n18144) );
  NAND2_X1 U15369 ( .A1(n12371), .A2(n18143), .ZN(n18128) );
  NAND2_X1 U15370 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12374), .ZN(
        n12375) );
  XNOR2_X1 U15371 ( .A(n12378), .B(n12383), .ZN(n12381) );
  NAND2_X1 U15372 ( .A1(n12381), .A2(n12380), .ZN(n12382) );
  XOR2_X1 U15373 ( .A(n12386), .B(n12387), .Z(n12384) );
  XOR2_X1 U15374 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12384), .Z(
        n18092) );
  NAND2_X1 U15375 ( .A1(n18091), .A2(n18092), .ZN(n18090) );
  NAND2_X1 U15376 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12384), .ZN(
        n12385) );
  AOI21_X1 U15377 ( .B1(n17648), .B2(n12451), .A(n18075), .ZN(n12390) );
  XNOR2_X1 U15378 ( .A(n12389), .B(n12388), .ZN(n18081) );
  NAND2_X1 U15379 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  NAND2_X1 U15380 ( .A1(n12429), .A2(n17997), .ZN(n18035) );
  OAI22_X1 U15381 ( .A1(n18340), .A2(n18193), .B1(n18376), .B2(n18338), .ZN(
        n18264) );
  NAND2_X1 U15382 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18393) );
  NOR2_X1 U15383 ( .A1(n12392), .A2(n18393), .ZN(n18262) );
  AOI21_X1 U15384 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18410) );
  INV_X1 U15385 ( .A(n18410), .ZN(n18428) );
  NAND2_X1 U15386 ( .A1(n18262), .A2(n18428), .ZN(n18368) );
  NAND3_X1 U15387 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18263) );
  NOR2_X1 U15388 ( .A1(n18368), .A2(n18263), .ZN(n12395) );
  INV_X1 U15389 ( .A(n12395), .ZN(n18276) );
  NAND3_X1 U15390 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18262), .ZN(n18367) );
  OR2_X1 U15391 ( .A1(n18263), .A2(n18367), .ZN(n18275) );
  NAND2_X1 U15392 ( .A1(n18930), .A2(n19106), .ZN(n18445) );
  NAND2_X1 U15393 ( .A1(n18930), .A2(n18916), .ZN(n18426) );
  NAND2_X1 U15394 ( .A1(n18445), .A2(n18426), .ZN(n18429) );
  OAI22_X1 U15395 ( .A1(n18943), .A2(n18276), .B1(n18275), .B2(n18429), .ZN(
        n12393) );
  NAND2_X1 U15396 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17939) );
  INV_X1 U15397 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18304) );
  INV_X1 U15398 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18352) );
  NOR2_X1 U15399 ( .A1(n18365), .A2(n18352), .ZN(n18344) );
  NAND2_X1 U15400 ( .A1(n18344), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18330) );
  INV_X1 U15401 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18336) );
  NOR2_X1 U15402 ( .A1(n18330), .A2(n18336), .ZN(n18329) );
  INV_X1 U15403 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18299) );
  NOR3_X1 U15404 ( .A1(n18304), .A2(n18319), .A3(n18299), .ZN(n18289) );
  NAND2_X1 U15405 ( .A1(n18289), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18265) );
  NOR2_X1 U15406 ( .A1(n17939), .A2(n18265), .ZN(n12394) );
  OAI21_X1 U15407 ( .B1(n18264), .B2(n12393), .A(n12394), .ZN(n18229) );
  NOR2_X1 U15408 ( .A1(n17888), .A2(n18229), .ZN(n18225) );
  NAND2_X1 U15409 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18225), .ZN(
        n18206) );
  NOR2_X1 U15410 ( .A1(n12577), .A2(n18206), .ZN(n12398) );
  INV_X1 U15411 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18228) );
  NOR2_X1 U15412 ( .A1(n17888), .A2(n18228), .ZN(n12396) );
  INV_X1 U15413 ( .A(n12396), .ZN(n17867) );
  NAND2_X1 U15414 ( .A1(n12395), .A2(n12394), .ZN(n18213) );
  NOR2_X1 U15415 ( .A1(n17867), .A2(n18213), .ZN(n18177) );
  AOI21_X1 U15416 ( .B1(n18177), .B2(n12454), .A(n18943), .ZN(n12452) );
  INV_X1 U15417 ( .A(n18289), .ZN(n18303) );
  NAND2_X1 U15418 ( .A1(n12396), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n18200) );
  NOR2_X1 U15419 ( .A1(n17939), .A2(n18200), .ZN(n12437) );
  INV_X1 U15420 ( .A(n12437), .ZN(n17851) );
  INV_X1 U15421 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n18191) );
  NOR2_X1 U15422 ( .A1(n17844), .A2(n18191), .ZN(n17843) );
  NAND2_X1 U15423 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18321), .ZN(
        n17994) );
  NAND2_X1 U15424 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18192), .ZN(
        n17846) );
  NAND2_X1 U15425 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17845), .ZN(
        n17804) );
  NOR2_X1 U15426 ( .A1(n18265), .A2(n18275), .ZN(n18256) );
  INV_X1 U15427 ( .A(n18256), .ZN(n18215) );
  INV_X1 U15428 ( .A(n17939), .ZN(n18260) );
  NAND2_X1 U15429 ( .A1(n18260), .A2(n12396), .ZN(n17870) );
  NOR2_X1 U15430 ( .A1(n18215), .A2(n17870), .ZN(n12576) );
  NAND2_X1 U15431 ( .A1(n18928), .A2(n19106), .ZN(n18434) );
  NAND2_X1 U15432 ( .A1(n12576), .A2(n18434), .ZN(n18195) );
  OAI21_X1 U15433 ( .B1(n18179), .B2(n18195), .A(n18426), .ZN(n18176) );
  INV_X1 U15434 ( .A(n18168), .ZN(n12397) );
  MUX2_X1 U15435 ( .A(n12398), .B(n12397), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n12448) );
  NAND2_X1 U15436 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18932), .ZN(
        n12407) );
  OAI22_X1 U15437 ( .A1(n19096), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18938), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12400) );
  XNOR2_X1 U15438 ( .A(n12401), .B(n12400), .ZN(n12413) );
  NOR2_X1 U15439 ( .A1(n12401), .A2(n12400), .ZN(n12402) );
  AOI21_X1 U15440 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18938), .A(
        n12402), .ZN(n12403) );
  AOI22_X1 U15441 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16143), .B1(
        n12403), .B2(n19085), .ZN(n12408) );
  INV_X1 U15442 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18479) );
  NOR2_X1 U15443 ( .A1(n12403), .A2(n19085), .ZN(n12409) );
  NAND2_X1 U15444 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16143), .ZN(
        n12404) );
  OAI22_X1 U15445 ( .A1(n12408), .A2(n18479), .B1(n12409), .B2(n12404), .ZN(
        n12406) );
  INV_X1 U15446 ( .A(n12406), .ZN(n12405) );
  OAI211_X1 U15447 ( .C1(n18932), .C2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12407), .B(n12405), .ZN(n12420) );
  XNOR2_X1 U15448 ( .A(n12407), .B(n12421), .ZN(n12412) );
  OAI21_X1 U15449 ( .B1(n18479), .B2(n12409), .A(n12408), .ZN(n12410) );
  OAI21_X1 U15450 ( .B1(n16143), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n12410), .ZN(n12411) );
  INV_X1 U15451 ( .A(n12411), .ZN(n12419) );
  OAI21_X1 U15452 ( .B1(n12413), .B2(n12420), .A(n18959), .ZN(n12556) );
  INV_X1 U15453 ( .A(n12556), .ZN(n18957) );
  OAI211_X1 U15454 ( .C1(n12417), .C2(n12416), .A(n12415), .B(n12414), .ZN(
        n16136) );
  INV_X1 U15455 ( .A(n12422), .ZN(n12423) );
  NAND2_X1 U15456 ( .A1(n19012), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19141) );
  INV_X2 U15457 ( .A(n19141), .ZN(n19069) );
  NAND2_X2 U15458 ( .A1(n19069), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19067) );
  OAI211_X1 U15459 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19012), .B(n19067), .ZN(n19130) );
  NAND2_X1 U15460 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19133) );
  INV_X1 U15461 ( .A(n19133), .ZN(n19004) );
  AOI21_X1 U15462 ( .B1(n12423), .B2(n19130), .A(n19004), .ZN(n16817) );
  NAND2_X1 U15463 ( .A1(n12425), .A2(n16817), .ZN(n12424) );
  OAI22_X1 U15464 ( .A1(n12425), .A2(n18962), .B1(n16816), .B2(n12424), .ZN(
        n12426) );
  INV_X1 U15465 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19143) );
  NAND2_X1 U15466 ( .A1(n19088), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18989) );
  NOR2_X1 U15467 ( .A1(n19143), .A2(n18989), .ZN(n19128) );
  INV_X1 U15468 ( .A(n19128), .ZN(n18983) );
  NOR2_X1 U15469 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17992) );
  INV_X1 U15470 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18298) );
  NAND3_X1 U15471 ( .A1(n17992), .A2(n18336), .A3(n18298), .ZN(n12432) );
  NAND3_X1 U15472 ( .A1(n12430), .A2(n18365), .A3(n18352), .ZN(n12431) );
  NOR2_X2 U15473 ( .A1(n12434), .A2(n18265), .ZN(n17956) );
  INV_X1 U15474 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18280) );
  NAND2_X1 U15475 ( .A1(n17955), .A2(n12436), .ZN(n17947) );
  NAND2_X1 U15476 ( .A1(n18260), .A2(n17956), .ZN(n17900) );
  NAND2_X1 U15477 ( .A1(n17956), .A2(n12437), .ZN(n12439) );
  NOR2_X1 U15478 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18075), .ZN(
        n17936) );
  INV_X1 U15479 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17925) );
  NAND2_X1 U15480 ( .A1(n17936), .A2(n17925), .ZN(n12438) );
  NOR2_X1 U15481 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12438), .ZN(
        n17901) );
  INV_X1 U15482 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n18219) );
  NAND2_X1 U15483 ( .A1(n17901), .A2(n18219), .ZN(n17887) );
  OR2_X1 U15484 ( .A1(n18075), .A2(n17849), .ZN(n17832) );
  OAI221_X1 U15485 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17997), 
        .C1(n18191), .C2(n17833), .A(n17832), .ZN(n17821) );
  NAND2_X1 U15486 ( .A1(n18075), .A2(n12441), .ZN(n12442) );
  NAND2_X1 U15487 ( .A1(n10157), .A2(n12442), .ZN(n12443) );
  NOR2_X2 U15488 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10149), .ZN(
        n12549) );
  INV_X1 U15489 ( .A(n12549), .ZN(n12444) );
  NAND2_X1 U15490 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10149), .ZN(
        n16151) );
  AOI21_X1 U15491 ( .B1(n17997), .B2(n12445), .A(n12450), .ZN(n17819) );
  INV_X1 U15492 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18986) );
  NOR2_X1 U15493 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19144) );
  NAND2_X1 U15494 ( .A1(n18455), .A2(n18461), .ZN(n18454) );
  INV_X1 U15495 ( .A(n18455), .ZN(n18444) );
  INV_X1 U15496 ( .A(n12449), .ZN(P3_U2835) );
  NAND2_X1 U15497 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18075), .ZN(
        n16150) );
  OAI21_X1 U15498 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18075), .A(
        n16150), .ZN(n17794) );
  NAND3_X1 U15499 ( .A1(n12462), .A2(n12557), .A3(n10165), .ZN(n12458) );
  NAND2_X1 U15500 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12576), .ZN(
        n18221) );
  NAND2_X1 U15501 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n12454), .ZN(
        n12463) );
  AOI221_X1 U15502 ( .B1(n18221), .B2(n18928), .C1(n12463), .C2(n18928), .A(
        n12452), .ZN(n12453) );
  OAI221_X1 U15503 ( .B1(n18930), .B2(n12454), .C1(n18930), .C2(n12576), .A(
        n12453), .ZN(n16144) );
  NOR2_X1 U15504 ( .A1(n18439), .A2(n16144), .ZN(n12580) );
  NAND2_X1 U15505 ( .A1(n12458), .A2(n12457), .ZN(n12461) );
  INV_X1 U15506 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17790) );
  NOR2_X1 U15507 ( .A1(n17790), .A2(n12455), .ZN(n16154) );
  INV_X1 U15508 ( .A(n16154), .ZN(n12459) );
  NOR2_X1 U15509 ( .A1(n17803), .A2(n12459), .ZN(n16708) );
  NOR2_X1 U15510 ( .A1(n12459), .A2(n17804), .ZN(n16711) );
  OAI22_X1 U15511 ( .A1(n16708), .A2(n18193), .B1(n16711), .B2(n18376), .ZN(
        n12460) );
  OAI211_X1 U15512 ( .C1(n12461), .C2(n12460), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18455), .ZN(n12469) );
  INV_X1 U15513 ( .A(n12462), .ZN(n12464) );
  OAI22_X1 U15514 ( .A1(n17997), .A2(n12464), .B1(n12463), .B2(n18206), .ZN(
        n12465) );
  NAND3_X1 U15515 ( .A1(n12465), .A2(n18438), .A3(n17790), .ZN(n12468) );
  NAND2_X1 U15516 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n9731), .ZN(n17799) );
  NAND3_X1 U15517 ( .A1(n12469), .A2(n12468), .A3(n12467), .ZN(P3_U2834) );
  AOI22_X1 U15518 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11306), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15519 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9737), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15520 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12494), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15521 ( .A1(n12050), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12471) );
  NAND4_X1 U15522 ( .A1(n12474), .A2(n12473), .A3(n12472), .A4(n12471), .ZN(
        n12481) );
  AOI22_X1 U15523 ( .A1(n12057), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15524 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15525 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15526 ( .A1(n12032), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U15527 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  OR2_X1 U15528 ( .A1(n12481), .A2(n12480), .ZN(n12501) );
  XNOR2_X1 U15529 ( .A(n12502), .B(n12501), .ZN(n12483) );
  NAND2_X1 U15530 ( .A1(n12483), .A2(n12482), .ZN(n12487) );
  INV_X1 U15531 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20939) );
  NAND2_X1 U15532 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n20939), .ZN(n20976) );
  AOI22_X1 U15533 ( .A1(n12513), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20976), 
        .B2(n20616), .ZN(n12486) );
  NAND2_X1 U15534 ( .A1(n12484), .A2(n20939), .ZN(n12485) );
  AOI22_X1 U15535 ( .A1(n12487), .A2(n12486), .B1(n12506), .B2(n15003), .ZN(
        n14720) );
  INV_X1 U15536 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14711) );
  XNOR2_X1 U15537 ( .A(n13487), .B(n14711), .ZN(n14995) );
  AOI22_X1 U15538 ( .A1(n11394), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12076), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15539 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11286), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15540 ( .A1(n12049), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11386), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15541 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12489), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12490) );
  NAND4_X1 U15542 ( .A1(n12493), .A2(n12492), .A3(n12491), .A4(n12490), .ZN(
        n12500) );
  AOI22_X1 U15543 ( .A1(n11739), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12057), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15544 ( .A1(n12475), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9730), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15545 ( .A1(n11298), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15546 ( .A1(n12494), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11701), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12495) );
  NAND4_X1 U15547 ( .A1(n12498), .A2(n12497), .A3(n12496), .A4(n12495), .ZN(
        n12499) );
  NOR2_X1 U15548 ( .A1(n12500), .A2(n12499), .ZN(n12505) );
  INV_X1 U15549 ( .A(n12501), .ZN(n12503) );
  NOR2_X1 U15550 ( .A1(n12503), .A2(n12502), .ZN(n12504) );
  XOR2_X1 U15551 ( .A(n12505), .B(n12504), .Z(n12510) );
  AOI21_X1 U15552 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20616), .A(
        n12506), .ZN(n12508) );
  NAND2_X1 U15553 ( .A1(n12513), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12507) );
  OAI211_X1 U15554 ( .C1(n12510), .C2(n12509), .A(n12508), .B(n12507), .ZN(
        n12511) );
  OAI21_X1 U15555 ( .B1(n13475), .B2(n14995), .A(n12511), .ZN(n14710) );
  AOI22_X1 U15556 ( .A1(n12513), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12512), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12514) );
  XNOR2_X2 U15557 ( .A(n14709), .B(n12514), .ZN(n14416) );
  NAND2_X1 U15558 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n16398) );
  NAND2_X1 U15559 ( .A1(n13479), .A2(n16398), .ZN(n12529) );
  NAND2_X1 U15560 ( .A1(n12516), .A2(n13495), .ZN(n12878) );
  NOR4_X1 U15561 ( .A1(n12521), .A2(n12520), .A3(n12519), .A4(n12518), .ZN(
        n12523) );
  NOR2_X1 U15562 ( .A1(n12523), .A2(n12522), .ZN(n12796) );
  NAND2_X1 U15563 ( .A1(n12796), .A2(n16398), .ZN(n12885) );
  NOR2_X1 U15564 ( .A1(n20197), .A2(n12885), .ZN(n12525) );
  INV_X1 U15565 ( .A(n20197), .ZN(n13132) );
  NAND3_X1 U15566 ( .A1(n14940), .A2(n13132), .A3(n11360), .ZN(n13134) );
  NOR2_X1 U15567 ( .A1(n13134), .A2(n11348), .ZN(n12524) );
  AOI22_X1 U15568 ( .A1(n13233), .A2(n12525), .B1(n12787), .B2(n12524), .ZN(
        n12526) );
  OAI21_X1 U15569 ( .B1(n13037), .B2(n12878), .A(n12526), .ZN(n12527) );
  INV_X1 U15570 ( .A(n12527), .ZN(n12528) );
  AND2_X1 U15571 ( .A1(n14290), .A2(n14940), .ZN(n12530) );
  NAND2_X1 U15572 ( .A1(n14416), .A2(n12530), .ZN(n12548) );
  NOR4_X1 U15573 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12534) );
  NOR4_X1 U15574 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n12533) );
  NOR4_X1 U15575 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12532) );
  NOR4_X1 U15576 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12531) );
  AND4_X1 U15577 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n12540) );
  NOR4_X1 U15578 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n12538) );
  NOR4_X1 U15579 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n12537) );
  NOR4_X1 U15580 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n12536) );
  INV_X1 U15581 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12535) );
  AND4_X1 U15582 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12539) );
  NAND2_X1 U15583 ( .A1(n12540), .A2(n12539), .ZN(n12541) );
  NOR2_X1 U15584 ( .A1(n12791), .A2(n13197), .ZN(n12542) );
  NAND2_X1 U15585 ( .A1(n14290), .A2(n12542), .ZN(n16289) );
  INV_X1 U15586 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16727) );
  NOR2_X1 U15587 ( .A1(n16289), .A2(n16727), .ZN(n12546) );
  NOR3_X1 U15588 ( .A1(n16280), .A2(n14279), .A3(n12791), .ZN(n12543) );
  AOI22_X1 U15589 ( .A1(n16284), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n16280), .ZN(n12544) );
  INV_X1 U15590 ( .A(n12544), .ZN(n12545) );
  NOR2_X1 U15591 ( .A1(n12546), .A2(n12545), .ZN(n12547) );
  NAND2_X1 U15592 ( .A1(n12548), .A2(n12547), .ZN(P1_U2873) );
  INV_X1 U15593 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19089) );
  NOR2_X1 U15594 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19089), .ZN(
        n12584) );
  INV_X1 U15595 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16713) );
  NAND3_X1 U15596 ( .A1(n12549), .A2(n17790), .A3(n17997), .ZN(n16149) );
  NOR2_X1 U15597 ( .A1(n18075), .A2(n16198), .ZN(n12551) );
  AOI211_X1 U15598 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n19089), .A(
        n16199), .B(n12551), .ZN(n12550) );
  AOI22_X1 U15599 ( .A1(n18075), .A2(n19089), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17997), .ZN(n12552) );
  OAI21_X1 U15600 ( .B1(n12584), .B2(n12550), .A(n12552), .ZN(n12555) );
  AOI221_X1 U15601 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C1(n16199), .C2(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(n12551), .ZN(n12553) );
  OR2_X1 U15602 ( .A1(n12553), .A2(n12552), .ZN(n12554) );
  NAND2_X1 U15603 ( .A1(n12555), .A2(n12554), .ZN(n12573) );
  NAND2_X1 U15604 ( .A1(n12573), .A2(n18076), .ZN(n12572) );
  NAND2_X1 U15605 ( .A1(n16154), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16201) );
  NAND2_X1 U15606 ( .A1(n16709), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12558) );
  XNOR2_X1 U15607 ( .A(n19089), .B(n12558), .ZN(n12589) );
  NAND2_X1 U15608 ( .A1(n16712), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12559) );
  XOR2_X1 U15609 ( .A(n12559), .B(n19089), .Z(n12574) );
  OAI21_X1 U15610 ( .B1(n19088), .B2(n19143), .A(n19079), .ZN(n19127) );
  INV_X1 U15611 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19131) );
  NOR2_X1 U15612 ( .A1(n19088), .A2(n19131), .ZN(n18121) );
  INV_X1 U15613 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16846) );
  INV_X1 U15614 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18155) );
  NAND3_X1 U15615 ( .A1(n18067), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17046) );
  NAND2_X1 U15616 ( .A1(n18066), .A2(n18030), .ZN(n18004) );
  NAND2_X1 U15617 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18006) );
  NAND2_X1 U15618 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17960) );
  NAND2_X1 U15619 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17919) );
  INV_X1 U15620 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17898) );
  INV_X1 U15621 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17884) );
  NOR2_X1 U15622 ( .A1(n17898), .A2(n17884), .ZN(n17883) );
  INV_X1 U15623 ( .A(n17883), .ZN(n12560) );
  NAND2_X1 U15624 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17838) );
  NAND2_X1 U15625 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17823), .ZN(
        n17796) );
  NAND2_X1 U15626 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17797) );
  INV_X1 U15627 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19071) );
  NOR2_X1 U15628 ( .A1(n18455), .A2(n19071), .ZN(n12582) );
  NAND2_X1 U15629 ( .A1(n18986), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18163) );
  NAND3_X1 U15630 ( .A1(n19079), .A2(n19143), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18722) );
  NOR2_X1 U15631 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19079), .ZN(
        n19104) );
  AOI221_X1 U15632 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n19088), .C1(n19143), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n19104), .ZN(n12561) );
  INV_X1 U15633 ( .A(n12561), .ZN(n18483) );
  INV_X2 U15634 ( .A(n18826), .ZN(n18862) );
  OR2_X1 U15635 ( .A1(n12562), .A2(n18005), .ZN(n16701) );
  XNOR2_X1 U15636 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n12565) );
  INV_X1 U15637 ( .A(n12562), .ZN(n12564) );
  INV_X1 U15638 ( .A(n18163), .ZN(n18002) );
  INV_X1 U15639 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12639) );
  NOR2_X1 U15640 ( .A1(n18155), .A2(n17837), .ZN(n12642) );
  INV_X1 U15641 ( .A(n12642), .ZN(n12641) );
  NOR2_X1 U15642 ( .A1(n17838), .A2(n12641), .ZN(n17791) );
  INV_X1 U15643 ( .A(n17791), .ZN(n12638) );
  NOR2_X1 U15644 ( .A1(n12639), .A2(n12638), .ZN(n16838) );
  NAND2_X1 U15645 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16838), .ZN(
        n16837) );
  INV_X1 U15646 ( .A(n16837), .ZN(n16836) );
  NAND2_X1 U15647 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16836), .ZN(
        n16835) );
  AOI21_X1 U15648 ( .B1(n18002), .B2(n16835), .A(n18119), .ZN(n12563) );
  OAI21_X1 U15649 ( .B1(n12564), .B2(n18826), .A(n12563), .ZN(n16718) );
  AOI21_X1 U15650 ( .B1(n17944), .B2(n9992), .A(n16718), .ZN(n16700) );
  OAI22_X1 U15651 ( .A1(n16701), .A2(n12565), .B1(n16700), .B2(n16846), .ZN(
        n12566) );
  AOI211_X1 U15652 ( .C1(n17943), .C2(n17171), .A(n12582), .B(n12566), .ZN(
        n12567) );
  NAND2_X1 U15653 ( .A1(n12572), .A2(n12571), .ZN(P3_U2799) );
  NAND2_X1 U15654 ( .A1(n12573), .A2(n18378), .ZN(n12592) );
  INV_X1 U15655 ( .A(n18460), .ZN(n16147) );
  INV_X1 U15656 ( .A(n12574), .ZN(n12579) );
  INV_X1 U15657 ( .A(n18429), .ZN(n12575) );
  AOI22_X1 U15658 ( .A1(n18963), .A2(n18177), .B1(n12576), .B2(n12575), .ZN(
        n18175) );
  NOR2_X1 U15659 ( .A1(n18175), .A2(n12577), .ZN(n16153) );
  NAND3_X1 U15660 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16153), .A3(
        n19089), .ZN(n12578) );
  OAI22_X1 U15661 ( .A1(n18376), .A2(n12579), .B1(n16201), .B2(n12578), .ZN(
        n12587) );
  NOR2_X1 U15662 ( .A1(n9886), .A2(n18461), .ZN(n18446) );
  INV_X1 U15663 ( .A(n12580), .ZN(n12581) );
  AOI21_X1 U15664 ( .B1(n18370), .B2(n16201), .A(n12581), .ZN(n16195) );
  NOR3_X1 U15665 ( .A1(n9731), .A2(n16195), .A3(n19089), .ZN(n12583) );
  AOI211_X1 U15666 ( .C1(n12584), .C2(n18446), .A(n12583), .B(n12582), .ZN(
        n12585) );
  INV_X1 U15667 ( .A(n12585), .ZN(n12586) );
  INV_X1 U15668 ( .A(n12590), .ZN(n12591) );
  NAND2_X1 U15669 ( .A1(n12592), .A2(n12591), .ZN(P3_U2831) );
  INV_X1 U15670 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20692) );
  NOR3_X1 U15671 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20692), .ZN(n12594) );
  NOR4_X1 U15672 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12593) );
  NAND4_X1 U15673 ( .A1(n14279), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12594), .A4(
        n12593), .ZN(U214) );
  NOR4_X1 U15674 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12598) );
  NOR4_X1 U15675 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12597) );
  NOR4_X1 U15676 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12596) );
  NOR4_X1 U15677 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12595) );
  NAND4_X1 U15678 ( .A1(n12598), .A2(n12597), .A3(n12596), .A4(n12595), .ZN(
        n12603) );
  NOR4_X1 U15679 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n12601) );
  NOR4_X1 U15680 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12600) );
  NOR4_X1 U15681 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12599) );
  INV_X1 U15682 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20083) );
  NAND4_X1 U15683 ( .A1(n12601), .A2(n12600), .A3(n12599), .A4(n20083), .ZN(
        n12602) );
  OAI21_X2 U15684 ( .B1(n12603), .B2(n12602), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13715) );
  NOR2_X1 U15685 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12605) );
  NOR4_X1 U15686 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12604) );
  NAND4_X1 U15687 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12605), .A4(n12604), .ZN(n12606) );
  NOR2_X1 U15688 ( .A1(n13715), .A2(n12606), .ZN(n16726) );
  NAND2_X1 U15689 ( .A1(n16726), .A2(U214), .ZN(U212) );
  NOR2_X1 U15690 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12606), .ZN(n16806)
         );
  INV_X1 U15691 ( .A(n13639), .ZN(n12608) );
  INV_X1 U15692 ( .A(n20559), .ZN(n20561) );
  NAND2_X1 U15693 ( .A1(n14048), .A2(n20561), .ZN(n12609) );
  NAND2_X1 U15694 ( .A1(n20561), .A2(n20818), .ZN(n14150) );
  OAI21_X1 U15695 ( .B1(n12609), .B2(n20544), .A(n14150), .ZN(n12623) );
  INV_X1 U15696 ( .A(n12611), .ZN(n13568) );
  NAND2_X1 U15697 ( .A1(n13629), .A2(n13568), .ZN(n20520) );
  NOR2_X1 U15698 ( .A1(n20520), .A2(n12613), .ZN(n12618) );
  NOR2_X1 U15699 ( .A1(n12619), .A2(n20616), .ZN(n14154) );
  OR2_X1 U15700 ( .A1(n13919), .A2(n16172), .ZN(n12620) );
  INV_X1 U15701 ( .A(n12620), .ZN(n14104) );
  INV_X1 U15702 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n16406) );
  NAND2_X1 U15703 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16397) );
  INV_X1 U15704 ( .A(n16397), .ZN(n13243) );
  OAI21_X1 U15705 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_2__SCAN_IN), .A(n10118), .ZN(n20702) );
  INV_X1 U15706 ( .A(DATAI_6_), .ZN(n12615) );
  NAND2_X1 U15707 ( .A1(n14279), .A2(BUF1_REG_6__SCAN_IN), .ZN(n12614) );
  OAI21_X1 U15708 ( .B1(n14279), .B2(n12615), .A(n12614), .ZN(n14968) );
  INV_X1 U15709 ( .A(n14968), .ZN(n13445) );
  NOR2_X1 U15710 ( .A1(n14051), .A2(n14165), .ZN(n12631) );
  NOR2_X2 U15711 ( .A1(n15147), .A2(n13197), .ZN(n13576) );
  NOR2_X2 U15712 ( .A1(n14279), .A2(n15147), .ZN(n13575) );
  AOI22_X1 U15713 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13576), .B1(DATAI_30_), 
        .B2(n13575), .ZN(n20602) );
  INV_X1 U15714 ( .A(n20602), .ZN(n20481) );
  AND2_X1 U15715 ( .A1(n20544), .A2(n20481), .ZN(n12630) );
  AOI22_X1 U15716 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13576), .B1(DATAI_22_), 
        .B2(n13575), .ZN(n20484) );
  NOR2_X1 U15717 ( .A1(n14048), .A2(n20484), .ZN(n12629) );
  INV_X1 U15718 ( .A(n13578), .ZN(n12616) );
  NAND2_X1 U15719 ( .A1(n12616), .A2(n11360), .ZN(n13780) );
  NOR3_X1 U15720 ( .A1(n16172), .A2(n16166), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13320) );
  INV_X1 U15721 ( .A(n13320), .ZN(n12617) );
  NOR2_X1 U15722 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12617), .ZN(
        n14046) );
  INV_X1 U15723 ( .A(n14046), .ZN(n12627) );
  INV_X1 U15724 ( .A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12626) );
  INV_X1 U15725 ( .A(n12618), .ZN(n12622) );
  NAND2_X1 U15726 ( .A1(n12619), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20451) );
  NAND2_X1 U15727 ( .A1(n13239), .A2(n20451), .ZN(n14158) );
  NAND2_X1 U15728 ( .A1(n12620), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14109) );
  INV_X1 U15729 ( .A(n14109), .ZN(n12621) );
  AOI211_X1 U15730 ( .C1(n12623), .C2(n12622), .A(n14158), .B(n12621), .ZN(
        n12624) );
  INV_X1 U15731 ( .A(n14045), .ZN(n12625) );
  OAI22_X1 U15732 ( .A1(n13780), .A2(n12627), .B1(n12626), .B2(n12625), .ZN(
        n12628) );
  OR4_X1 U15733 ( .A1(n12631), .A2(n12630), .A3(n12629), .A4(n12628), .ZN(
        P1_U3119) );
  NOR3_X1 U15734 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17166) );
  INV_X1 U15735 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17164) );
  NAND2_X1 U15736 ( .A1(n17166), .A2(n17164), .ZN(n17160) );
  NOR2_X1 U15737 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17160), .ZN(n17134) );
  INV_X1 U15738 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17499) );
  NAND2_X1 U15739 ( .A1(n17134), .A2(n17499), .ZN(n17129) );
  NOR2_X1 U15740 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17129), .ZN(n17113) );
  INV_X1 U15741 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17435) );
  NAND2_X1 U15742 ( .A1(n17113), .A2(n17435), .ZN(n17110) );
  INV_X1 U15743 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17082) );
  NAND2_X1 U15744 ( .A1(n17079), .A2(n17082), .ZN(n17062) );
  INV_X1 U15745 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17060) );
  NAND2_X1 U15746 ( .A1(n17061), .A2(n17060), .ZN(n17052) );
  INV_X1 U15747 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17405) );
  NAND2_X1 U15748 ( .A1(n17034), .A2(n17405), .ZN(n17030) );
  INV_X1 U15749 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20865) );
  NAND2_X1 U15750 ( .A1(n17016), .A2(n20865), .ZN(n17006) );
  INV_X1 U15751 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17348) );
  NAND2_X1 U15752 ( .A1(n16987), .A2(n17348), .ZN(n16981) );
  NOR2_X1 U15753 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16981), .ZN(n16965) );
  INV_X1 U15754 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17319) );
  NAND2_X1 U15755 ( .A1(n16965), .A2(n17319), .ZN(n16960) );
  NOR2_X1 U15756 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16960), .ZN(n16941) );
  INV_X1 U15757 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17292) );
  NAND2_X1 U15758 ( .A1(n16941), .A2(n17292), .ZN(n16938) );
  NOR2_X1 U15759 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16938), .ZN(n16925) );
  INV_X1 U15760 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16921) );
  NAND2_X1 U15761 ( .A1(n16925), .A2(n16921), .ZN(n16918) );
  NOR2_X1 U15762 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16918), .ZN(n16890) );
  INV_X1 U15763 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16892) );
  NAND2_X1 U15764 ( .A1(n16890), .A2(n16892), .ZN(n12634) );
  NOR2_X1 U15765 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n12634), .ZN(n16886) );
  OAI21_X2 U15766 ( .B1(n18923), .B2(n18922), .A(n17728), .ZN(n16135) );
  NOR2_X1 U15767 ( .A1(n12632), .A2(n16135), .ZN(n18958) );
  NAND2_X1 U15768 ( .A1(n19146), .A2(n16211), .ZN(n12648) );
  NAND2_X1 U15769 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17729), .ZN(n12633) );
  AOI211_X4 U15770 ( .C1(n19133), .C2(n19131), .A(n12648), .B(n12633), .ZN(
        n17196) );
  AOI211_X1 U15771 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n12634), .A(n16886), .B(
        n17165), .ZN(n12654) );
  INV_X1 U15772 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19060) );
  AOI211_X1 U15773 ( .C1(n19132), .C2(n19130), .A(n19004), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n12649) );
  INV_X1 U15774 ( .A(n12649), .ZN(n18977) );
  INV_X1 U15775 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19055) );
  INV_X1 U15776 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19051) );
  INV_X1 U15777 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19036) );
  INV_X1 U15778 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20772) );
  INV_X1 U15779 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19022) );
  INV_X1 U15780 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19019) );
  NAND2_X1 U15781 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n17150) );
  NOR2_X1 U15782 ( .A1(n19019), .A2(n17150), .ZN(n17145) );
  NAND2_X1 U15783 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n17145), .ZN(n17089) );
  NOR2_X1 U15784 ( .A1(n19022), .A2(n17089), .ZN(n17104) );
  NAND4_X1 U15785 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n17104), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n17063) );
  NAND2_X1 U15786 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n17064) );
  NOR3_X1 U15787 ( .A1(n20772), .A2(n17063), .A3(n17064), .ZN(n17041) );
  NAND2_X1 U15788 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17041), .ZN(n17024) );
  NOR2_X1 U15789 ( .A1(n19036), .A2(n17024), .ZN(n17009) );
  NAND2_X1 U15790 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n17009), .ZN(n17010) );
  NAND3_X1 U15791 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16944) );
  NAND3_X1 U15792 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16935) );
  NOR4_X1 U15793 ( .A1(n19051), .A2(n17010), .A3(n16944), .A4(n16935), .ZN(
        n16922) );
  NAND2_X1 U15794 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16922), .ZN(n16914) );
  NOR2_X1 U15795 ( .A1(n19055), .A2(n16914), .ZN(n16912) );
  NAND2_X1 U15796 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16912), .ZN(n12635) );
  NOR2_X1 U15797 ( .A1(n17173), .A2(n12635), .ZN(n16897) );
  NAND2_X1 U15798 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16897), .ZN(n16833) );
  INV_X1 U15799 ( .A(n19146), .ZN(n19126) );
  NAND3_X1 U15800 ( .A1(n18986), .A2(n19143), .A3(n19131), .ZN(n18994) );
  NOR2_X1 U15801 ( .A1(n19088), .A2(n18994), .ZN(n17184) );
  NAND2_X1 U15802 ( .A1(n19143), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18856) );
  OR2_X1 U15803 ( .A1(n18989), .A2(n18856), .ZN(n18981) );
  INV_X1 U15804 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19058) );
  NOR3_X1 U15805 ( .A1(n17185), .A2(n12635), .A3(n19058), .ZN(n12636) );
  NOR2_X1 U15806 ( .A1(n17178), .A2(n17185), .ZN(n16957) );
  AOI21_X1 U15807 ( .B1(P3_REIP_REG_26__SCAN_IN), .B2(n12636), .A(n16957), 
        .ZN(n16883) );
  INV_X1 U15808 ( .A(n16883), .ZN(n12637) );
  AOI21_X1 U15809 ( .B1(n19060), .B2(n16833), .A(n12637), .ZN(n12653) );
  AOI21_X1 U15810 ( .B1(n12639), .B2(n12638), .A(n16838), .ZN(n17824) );
  INV_X1 U15811 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17840) );
  NAND2_X1 U15812 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12642), .ZN(
        n12640) );
  AOI21_X1 U15813 ( .B1(n17840), .B2(n12640), .A(n17791), .ZN(n17842) );
  INV_X1 U15814 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17855) );
  AOI22_X1 U15815 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12642), .B1(
        n12641), .B2(n17855), .ZN(n17853) );
  INV_X1 U15816 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17836) );
  NOR2_X1 U15817 ( .A1(n18155), .A2(n17882), .ZN(n12645) );
  NAND2_X1 U15818 ( .A1(n17883), .A2(n12645), .ZN(n12643) );
  AOI21_X1 U15819 ( .B1(n17836), .B2(n12643), .A(n12642), .ZN(n17874) );
  NAND2_X1 U15820 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12645), .ZN(
        n12644) );
  INV_X1 U15821 ( .A(n12643), .ZN(n17835) );
  AOI21_X1 U15822 ( .B1(n17884), .B2(n12644), .A(n17835), .ZN(n17881) );
  XNOR2_X1 U15823 ( .A(n17898), .B(n12645), .ZN(n17894) );
  INV_X1 U15824 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12646) );
  NOR2_X1 U15825 ( .A1(n18155), .A2(n17918), .ZN(n17917) );
  NAND2_X1 U15826 ( .A1(n9981), .A2(n17917), .ZN(n17880) );
  AOI21_X1 U15827 ( .B1(n12646), .B2(n17880), .A(n12645), .ZN(n17911) );
  INV_X1 U15828 ( .A(n17917), .ZN(n16953) );
  NOR2_X1 U15829 ( .A1(n18155), .A2(n17959), .ZN(n17958) );
  NAND2_X1 U15830 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17958), .ZN(
        n17000) );
  NOR2_X1 U15831 ( .A1(n17000), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16978) );
  INV_X1 U15832 ( .A(n16978), .ZN(n17001) );
  NOR2_X1 U15833 ( .A1(n16953), .A2(n17001), .ZN(n16966) );
  AOI21_X1 U15834 ( .B1(n9981), .B2(n16966), .A(n9816), .ZN(n16947) );
  NOR2_X1 U15835 ( .A1(n17911), .A2(n16947), .ZN(n16946) );
  NOR2_X1 U15836 ( .A1(n16946), .A2(n9816), .ZN(n16933) );
  NOR2_X1 U15837 ( .A1(n17894), .A2(n16933), .ZN(n16932) );
  NOR2_X1 U15838 ( .A1(n16932), .A2(n9816), .ZN(n16924) );
  NOR2_X1 U15839 ( .A1(n17881), .A2(n16924), .ZN(n16923) );
  NOR2_X1 U15840 ( .A1(n16923), .A2(n9816), .ZN(n16911) );
  NOR2_X1 U15841 ( .A1(n17874), .A2(n16911), .ZN(n16910) );
  NOR2_X1 U15842 ( .A1(n16894), .A2(n9816), .ZN(n12647) );
  NOR2_X1 U15843 ( .A1(n17824), .A2(n12647), .ZN(n16839) );
  AOI211_X1 U15844 ( .C1(n17824), .C2(n12647), .A(n16839), .B(n18992), .ZN(
        n12652) );
  AOI211_X4 U15845 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17729), .A(n12649), .B(
        n12648), .ZN(n17197) );
  AOI22_X1 U15846 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17182), .B1(
        n17197), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n12650) );
  INV_X1 U15847 ( .A(n12650), .ZN(n12651) );
  OR4_X1 U15848 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        P3_U2645) );
  OR2_X1 U15849 ( .A1(n16656), .A2(n12667), .ZN(n12722) );
  NOR2_X1 U15850 ( .A1(n16657), .A2(n12722), .ZN(n19349) );
  INV_X1 U15851 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12658) );
  NAND2_X1 U15852 ( .A1(n12655), .A2(n16682), .ZN(n12656) );
  NOR2_X2 U15853 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20152) );
  INV_X1 U15854 ( .A(n20152), .ZN(n20129) );
  NOR2_X1 U15855 ( .A1(n20129), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12668) );
  INV_X1 U15856 ( .A(n12668), .ZN(n12657) );
  OAI211_X1 U15857 ( .C1(n19349), .C2(n12658), .A(n12670), .B(n12657), .ZN(
        P2_U2814) );
  OR2_X1 U15858 ( .A1(n16657), .A2(n12659), .ZN(n12690) );
  AND2_X1 U15859 ( .A1(n12660), .A2(n20190), .ZN(n13426) );
  OR2_X1 U15860 ( .A1(n13426), .A2(n12688), .ZN(n12661) );
  NOR2_X1 U15861 ( .A1(n12690), .A2(n12661), .ZN(n16651) );
  OR2_X1 U15862 ( .A1(n16651), .A2(n12667), .ZN(n20176) );
  INV_X1 U15863 ( .A(n20176), .ZN(n12666) );
  NAND2_X1 U15864 ( .A1(n20170), .A2(n12662), .ZN(n12663) );
  NAND2_X1 U15865 ( .A1(n12664), .A2(n12663), .ZN(n12665) );
  NAND2_X1 U15866 ( .A1(n12665), .A2(n16682), .ZN(n12871) );
  OAI21_X1 U15867 ( .B1(n12666), .B2(n20943), .A(n12871), .ZN(P2_U2819) );
  INV_X1 U15868 ( .A(n20188), .ZN(n19152) );
  OAI21_X1 U15869 ( .B1(n12668), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19152), 
        .ZN(n12669) );
  OAI21_X1 U15870 ( .B1(n20181), .B2(n19152), .A(n12669), .ZN(P2_U3612) );
  INV_X1 U15871 ( .A(n12670), .ZN(n13516) );
  OAI21_X1 U15872 ( .B1(n9740), .B2(n20190), .A(n13516), .ZN(n12740) );
  AOI22_X1 U15873 ( .A1(P2_UWORD_REG_8__SCAN_IN), .A2(n12740), .B1(n12717), 
        .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12675) );
  NOR3_X1 U15874 ( .A1(n12670), .A2(n9740), .A3(n20183), .ZN(n12671) );
  INV_X1 U15875 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n12672) );
  NOR2_X1 U15876 ( .A1(n13716), .A2(n12672), .ZN(n12673) );
  AOI21_X1 U15877 ( .B1(BUF1_REG_8__SCAN_IN), .B2(n13716), .A(n12673), .ZN(
        n19380) );
  INV_X1 U15878 ( .A(n19380), .ZN(n12674) );
  NAND2_X1 U15879 ( .A1(n12750), .A2(n12674), .ZN(n12763) );
  NAND2_X1 U15880 ( .A1(n12675), .A2(n12763), .ZN(P2_U2960) );
  AOI22_X1 U15881 ( .A1(P2_UWORD_REG_10__SCAN_IN), .A2(n12740), .B1(n12717), 
        .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12679) );
  INV_X1 U15882 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n12676) );
  NOR2_X1 U15883 ( .A1(n13716), .A2(n12676), .ZN(n12677) );
  AOI21_X1 U15884 ( .B1(BUF1_REG_10__SCAN_IN), .B2(n13716), .A(n12677), .ZN(
        n19374) );
  INV_X1 U15885 ( .A(n19374), .ZN(n12678) );
  NAND2_X1 U15886 ( .A1(n12750), .A2(n12678), .ZN(n12745) );
  NAND2_X1 U15887 ( .A1(n12679), .A2(n12745), .ZN(P2_U2962) );
  AOI22_X1 U15888 ( .A1(P2_UWORD_REG_3__SCAN_IN), .A2(n12740), .B1(n12717), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U15889 ( .A1(n13716), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13715), .ZN(n19403) );
  INV_X1 U15890 ( .A(n19403), .ZN(n12680) );
  NAND2_X1 U15891 ( .A1(n12750), .A2(n12680), .ZN(n12760) );
  NAND2_X1 U15892 ( .A1(n12681), .A2(n12760), .ZN(P2_U2955) );
  AOI22_X1 U15893 ( .A1(P2_UWORD_REG_7__SCAN_IN), .A2(n12740), .B1(n12717), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12682) );
  OAI22_X1 U15894 ( .A1(n13715), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13716), .ZN(n19382) );
  INV_X1 U15895 ( .A(n19382), .ZN(n16466) );
  NAND2_X1 U15896 ( .A1(n12750), .A2(n16466), .ZN(n12758) );
  NAND2_X1 U15897 ( .A1(n12682), .A2(n12758), .ZN(P2_U2959) );
  AOI22_X1 U15898 ( .A1(P2_UWORD_REG_5__SCAN_IN), .A2(n12762), .B1(n12717), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15899 ( .A1(n13716), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13715), .ZN(n19395) );
  INV_X1 U15900 ( .A(n19395), .ZN(n12683) );
  NAND2_X1 U15901 ( .A1(n12750), .A2(n12683), .ZN(n12754) );
  NAND2_X1 U15902 ( .A1(n12684), .A2(n12754), .ZN(P2_U2957) );
  AOI22_X1 U15903 ( .A1(P2_UWORD_REG_4__SCAN_IN), .A2(n12762), .B1(n12717), 
        .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12686) );
  AOI22_X1 U15904 ( .A1(n13716), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13715), .ZN(n19526) );
  INV_X1 U15905 ( .A(n19526), .ZN(n12685) );
  NAND2_X1 U15906 ( .A1(n12750), .A2(n12685), .ZN(n12747) );
  NAND2_X1 U15907 ( .A1(n12686), .A2(n12747), .ZN(P2_U2956) );
  AOI22_X1 U15908 ( .A1(P2_UWORD_REG_6__SCAN_IN), .A2(n12740), .B1(n12717), 
        .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n12687) );
  INV_X1 U15909 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16765) );
  INV_X1 U15910 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18509) );
  AOI22_X1 U15911 ( .A1(n13716), .A2(n16765), .B1(n18509), .B2(n13715), .ZN(
        n19384) );
  NAND2_X1 U15912 ( .A1(n12750), .A2(n19384), .ZN(n12743) );
  NAND2_X1 U15913 ( .A1(n12687), .A2(n12743), .ZN(P2_U2958) );
  INV_X1 U15914 ( .A(n12688), .ZN(n12689) );
  OR2_X1 U15915 ( .A1(n16656), .A2(n12689), .ZN(n12695) );
  INV_X1 U15916 ( .A(n12690), .ZN(n12692) );
  AOI21_X1 U15917 ( .B1(n12692), .B2(n13426), .A(n12691), .ZN(n12693) );
  NAND2_X1 U15918 ( .A1(n12859), .A2(n16658), .ZN(n13424) );
  AND2_X1 U15919 ( .A1(n12693), .A2(n13424), .ZN(n12694) );
  INV_X1 U15920 ( .A(n12859), .ZN(n16661) );
  NAND2_X1 U15921 ( .A1(n16661), .A2(n16021), .ZN(n12835) );
  OAI211_X1 U15922 ( .C1(n12723), .C2(n12695), .A(n12694), .B(n12835), .ZN(
        n16646) );
  NAND2_X1 U15923 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n12860) );
  NOR2_X1 U15924 ( .A1(n19151), .A2(n12860), .ZN(n16210) );
  INV_X1 U15925 ( .A(n16210), .ZN(n16696) );
  OAI22_X1 U15926 ( .A1(n16696), .A2(n20943), .B1(P2_STATE2_REG_0__SCAN_IN), 
        .B2(n19670), .ZN(n12696) );
  AOI21_X1 U15927 ( .B1(n16646), .B2(n16682), .A(n12696), .ZN(n16045) );
  INV_X1 U15928 ( .A(n16045), .ZN(n12701) );
  INV_X1 U15929 ( .A(n16650), .ZN(n12697) );
  NOR4_X1 U15930 ( .A1(n16656), .A2(n12697), .A3(n20133), .A4(n19514), .ZN(
        n12698) );
  NAND2_X1 U15931 ( .A1(n12701), .A2(n12698), .ZN(n12699) );
  OAI21_X1 U15932 ( .B1(n12701), .B2(n12700), .A(n12699), .ZN(P2_U3595) );
  INV_X1 U15933 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12848) );
  NAND2_X1 U15934 ( .A1(n13715), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12703) );
  INV_X1 U15935 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16760) );
  OR2_X1 U15936 ( .A1(n13715), .A2(n16760), .ZN(n12702) );
  NAND2_X1 U15937 ( .A1(n12703), .A2(n12702), .ZN(n19377) );
  NAND2_X1 U15938 ( .A1(n12750), .A2(n19377), .ZN(n12709) );
  NAND2_X1 U15939 ( .A1(n12762), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12704) );
  OAI211_X1 U15940 ( .C1(n12848), .C2(n12727), .A(n12709), .B(n12704), .ZN(
        P2_U2961) );
  INV_X1 U15941 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n12857) );
  NAND2_X1 U15942 ( .A1(n13715), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12706) );
  INV_X1 U15943 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16754) );
  OR2_X1 U15944 ( .A1(n13715), .A2(n16754), .ZN(n12705) );
  NAND2_X1 U15945 ( .A1(n12706), .A2(n12705), .ZN(n19365) );
  NAND2_X1 U15946 ( .A1(n12750), .A2(n19365), .ZN(n12716) );
  NAND2_X1 U15947 ( .A1(n12762), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12707) );
  OAI211_X1 U15948 ( .C1(n12857), .C2(n12727), .A(n12716), .B(n12707), .ZN(
        P2_U2965) );
  INV_X1 U15949 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19439) );
  NAND2_X1 U15950 ( .A1(n12762), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12708) );
  OAI211_X1 U15951 ( .C1(n19439), .C2(n12727), .A(n12709), .B(n12708), .ZN(
        P2_U2976) );
  INV_X1 U15952 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n12855) );
  NAND2_X1 U15953 ( .A1(n13715), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12711) );
  INV_X1 U15954 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16756) );
  OR2_X1 U15955 ( .A1(n13715), .A2(n16756), .ZN(n12710) );
  NAND2_X1 U15956 ( .A1(n12711), .A2(n12710), .ZN(n19371) );
  NAND2_X1 U15957 ( .A1(n12750), .A2(n19371), .ZN(n12714) );
  NAND2_X1 U15958 ( .A1(n12762), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12712) );
  OAI211_X1 U15959 ( .C1(n12855), .C2(n12727), .A(n12714), .B(n12712), .ZN(
        P2_U2963) );
  INV_X1 U15960 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19436) );
  NAND2_X1 U15961 ( .A1(n12762), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12713) );
  OAI211_X1 U15962 ( .C1(n19436), .C2(n12727), .A(n12714), .B(n12713), .ZN(
        P2_U2978) );
  INV_X1 U15963 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n20804) );
  NAND2_X1 U15964 ( .A1(n12762), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12715) );
  OAI211_X1 U15965 ( .C1(n20804), .C2(n12727), .A(n12716), .B(n12715), .ZN(
        P2_U2980) );
  INV_X1 U15966 ( .A(n12750), .ZN(n12719) );
  AOI22_X1 U15967 ( .A1(n13716), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13715), .ZN(n19361) );
  AOI22_X1 U15968 ( .A1(P2_LWORD_REG_15__SCAN_IN), .A2(n12762), .B1(n12717), 
        .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12718) );
  OAI21_X1 U15969 ( .B1(n12719), .B2(n19361), .A(n12718), .ZN(P2_U2982) );
  AND2_X1 U15970 ( .A1(n12796), .A2(n12720), .ZN(n12765) );
  NAND2_X1 U15971 ( .A1(n12765), .A2(n13132), .ZN(n12802) );
  NAND2_X1 U15972 ( .A1(n20561), .A2(n20614), .ZN(n20200) );
  INV_X1 U15973 ( .A(n20200), .ZN(n12803) );
  AOI21_X1 U15974 ( .B1(n12802), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12803), 
        .ZN(n12721) );
  NAND2_X1 U15975 ( .A1(n13149), .A2(n12721), .ZN(P1_U2801) );
  OAI21_X1 U15976 ( .B1(n12723), .B2(n12722), .A(n12727), .ZN(n12724) );
  INV_X1 U15977 ( .A(n20068), .ZN(n20178) );
  NAND2_X1 U15978 ( .A1(n19458), .A2(n12725), .ZN(n19425) );
  INV_X1 U15979 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15576) );
  INV_X1 U15980 ( .A(n12860), .ZN(n12726) );
  NAND2_X1 U15981 ( .A1(n19151), .A2(n12726), .ZN(n19428) );
  INV_X1 U15982 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16795) );
  INV_X1 U15983 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n20835) );
  OAI222_X1 U15984 ( .A1(n19425), .A2(n15576), .B1(n19424), .B2(n16795), .C1(
        n19428), .C2(n20835), .ZN(P2_U2930) );
  AOI22_X1 U15985 ( .A1(P2_LWORD_REG_2__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15986 ( .A1(n13716), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13715), .ZN(n19518) );
  INV_X1 U15987 ( .A(n19518), .ZN(n12728) );
  NAND2_X1 U15988 ( .A1(n12750), .A2(n12728), .ZN(n12730) );
  NAND2_X1 U15989 ( .A1(n12729), .A2(n12730), .ZN(P2_U2969) );
  AOI22_X1 U15990 ( .A1(P2_UWORD_REG_2__SCAN_IN), .A2(n12740), .B1(n16411), 
        .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12731) );
  NAND2_X1 U15991 ( .A1(n12731), .A2(n12730), .ZN(P2_U2954) );
  AOI22_X1 U15992 ( .A1(P2_UWORD_REG_12__SCAN_IN), .A2(n12740), .B1(n16411), 
        .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15993 ( .A1(n13716), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13715), .ZN(n19368) );
  INV_X1 U15994 ( .A(n19368), .ZN(n12732) );
  NAND2_X1 U15995 ( .A1(n12750), .A2(n12732), .ZN(n12741) );
  NAND2_X1 U15996 ( .A1(n12733), .A2(n12741), .ZN(P2_U2964) );
  AOI22_X1 U15997 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12735) );
  AOI22_X1 U15998 ( .A1(n13716), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n13715), .ZN(n19363) );
  INV_X1 U15999 ( .A(n19363), .ZN(n12734) );
  NAND2_X1 U16000 ( .A1(n12750), .A2(n12734), .ZN(n12736) );
  NAND2_X1 U16001 ( .A1(n12735), .A2(n12736), .ZN(P2_U2981) );
  AOI22_X1 U16002 ( .A1(P2_UWORD_REG_14__SCAN_IN), .A2(n12740), .B1(n16411), 
        .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U16003 ( .A1(n12737), .A2(n12736), .ZN(P2_U2966) );
  AOI22_X1 U16004 ( .A1(P2_LWORD_REG_0__SCAN_IN), .A2(n12740), .B1(n16411), 
        .B2(P2_EAX_REG_0__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U16005 ( .A1(n13716), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13715), .ZN(n19508) );
  INV_X1 U16006 ( .A(n19508), .ZN(n12738) );
  NAND2_X1 U16007 ( .A1(n12750), .A2(n12738), .ZN(n12752) );
  NAND2_X1 U16008 ( .A1(n12739), .A2(n12752), .ZN(P2_U2967) );
  AOI22_X1 U16009 ( .A1(P2_LWORD_REG_12__SCAN_IN), .A2(n12740), .B1(n16411), 
        .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12742) );
  NAND2_X1 U16010 ( .A1(n12742), .A2(n12741), .ZN(P2_U2979) );
  AOI22_X1 U16011 ( .A1(P2_LWORD_REG_6__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12744) );
  NAND2_X1 U16012 ( .A1(n12744), .A2(n12743), .ZN(P2_U2973) );
  AOI22_X1 U16013 ( .A1(P2_LWORD_REG_10__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12746) );
  NAND2_X1 U16014 ( .A1(n12746), .A2(n12745), .ZN(P2_U2977) );
  AOI22_X1 U16015 ( .A1(P2_LWORD_REG_4__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12748) );
  NAND2_X1 U16016 ( .A1(n12748), .A2(n12747), .ZN(P2_U2971) );
  AOI22_X1 U16017 ( .A1(P2_UWORD_REG_1__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12751) );
  AOI22_X1 U16018 ( .A1(n13716), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13715), .ZN(n19515) );
  INV_X1 U16019 ( .A(n19515), .ZN(n12749) );
  NAND2_X1 U16020 ( .A1(n12750), .A2(n12749), .ZN(n12756) );
  NAND2_X1 U16021 ( .A1(n12751), .A2(n12756), .ZN(P2_U2953) );
  AOI22_X1 U16022 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U16023 ( .A1(n12753), .A2(n12752), .ZN(P2_U2952) );
  AOI22_X1 U16024 ( .A1(P2_LWORD_REG_5__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U16025 ( .A1(n12755), .A2(n12754), .ZN(P2_U2972) );
  AOI22_X1 U16026 ( .A1(P2_LWORD_REG_1__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U16027 ( .A1(n12757), .A2(n12756), .ZN(P2_U2968) );
  AOI22_X1 U16028 ( .A1(P2_LWORD_REG_7__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U16029 ( .A1(n12759), .A2(n12758), .ZN(P2_U2974) );
  AOI22_X1 U16030 ( .A1(P2_LWORD_REG_3__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_3__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U16031 ( .A1(n12761), .A2(n12760), .ZN(P2_U2970) );
  AOI22_X1 U16032 ( .A1(P2_LWORD_REG_8__SCAN_IN), .A2(n12762), .B1(n16411), 
        .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U16033 ( .A1(n12764), .A2(n12763), .ZN(P2_U2975) );
  NAND2_X1 U16034 ( .A1(n16187), .A2(n12772), .ZN(n12768) );
  INV_X1 U16035 ( .A(n12765), .ZN(n12766) );
  NAND2_X1 U16036 ( .A1(n12766), .A2(n12515), .ZN(n12767) );
  NAND2_X1 U16037 ( .A1(n12768), .A2(n12767), .ZN(n20198) );
  INV_X1 U16038 ( .A(n12769), .ZN(n12771) );
  INV_X1 U16039 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12770) );
  NAND2_X1 U16040 ( .A1(n12771), .A2(n12770), .ZN(n16208) );
  AND2_X4 U16041 ( .A1(n13472), .A2(n13479), .ZN(n14308) );
  NAND3_X1 U16042 ( .A1(n12772), .A2(n16208), .A3(n14341), .ZN(n12773) );
  AND2_X1 U16043 ( .A1(n12773), .A2(n16398), .ZN(n20699) );
  NOR2_X1 U16044 ( .A1(n20198), .A2(n20699), .ZN(n16173) );
  OR2_X1 U16045 ( .A1(n16173), .A2(n20197), .ZN(n12799) );
  INV_X1 U16046 ( .A(n12799), .ZN(n20205) );
  INV_X1 U16047 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12801) );
  NAND2_X1 U16048 ( .A1(n11355), .A2(n13495), .ZN(n12785) );
  AOI21_X1 U16049 ( .B1(n9862), .B2(n13282), .A(n13135), .ZN(n12774) );
  NAND2_X1 U16050 ( .A1(n12775), .A2(n12774), .ZN(n12776) );
  NAND2_X1 U16051 ( .A1(n12776), .A2(n13479), .ZN(n12784) );
  INV_X1 U16052 ( .A(n12777), .ZN(n12778) );
  NOR2_X1 U16053 ( .A1(n12779), .A2(n12778), .ZN(n12783) );
  NAND2_X1 U16054 ( .A1(n11359), .A2(n13472), .ZN(n12780) );
  NAND2_X1 U16055 ( .A1(n12780), .A2(n20700), .ZN(n12781) );
  NAND2_X1 U16056 ( .A1(n12782), .A2(n12781), .ZN(n12883) );
  INV_X1 U16057 ( .A(n12786), .ZN(n12877) );
  INV_X1 U16058 ( .A(n12787), .ZN(n12788) );
  AND3_X1 U16059 ( .A1(n12877), .A2(n12788), .A3(n13052), .ZN(n12789) );
  NAND2_X1 U16060 ( .A1(n13051), .A2(n12789), .ZN(n12790) );
  NOR2_X1 U16061 ( .A1(n12790), .A2(n13233), .ZN(n12924) );
  AND2_X1 U16062 ( .A1(n12791), .A2(n13472), .ZN(n13032) );
  NAND2_X1 U16063 ( .A1(n16175), .A2(n12878), .ZN(n13042) );
  INV_X1 U16064 ( .A(n13042), .ZN(n12793) );
  NAND2_X1 U16065 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  MUX2_X1 U16066 ( .A(n13133), .B(n12794), .S(n16187), .Z(n12798) );
  INV_X1 U16067 ( .A(n12720), .ZN(n12795) );
  NOR2_X1 U16068 ( .A1(n12796), .A2(n12795), .ZN(n12797) );
  OR2_X1 U16069 ( .A1(n12799), .A2(n16176), .ZN(n12800) );
  OAI21_X1 U16070 ( .B1(n20205), .B2(n12801), .A(n12800), .ZN(P1_U3484) );
  INV_X2 U16071 ( .A(n13172), .ZN(n14705) );
  NOR2_X1 U16072 ( .A1(n13495), .A2(n14705), .ZN(n12805) );
  OAI21_X1 U16073 ( .B1(n12803), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20696), 
        .ZN(n12804) );
  OAI21_X1 U16074 ( .B1(n20696), .B2(n12805), .A(n12804), .ZN(P1_U3487) );
  XOR2_X1 U16075 ( .A(n12807), .B(n12806), .Z(n12870) );
  NAND2_X1 U16076 ( .A1(n12809), .A2(n12808), .ZN(n12872) );
  AND3_X1 U16077 ( .A1(n12872), .A2(n16639), .A3(n12873), .ZN(n12818) );
  OR2_X1 U16078 ( .A1(n12811), .A2(n12810), .ZN(n12813) );
  NAND2_X1 U16079 ( .A1(n12813), .A2(n12812), .ZN(n20147) );
  INV_X1 U16080 ( .A(n20147), .ZN(n12816) );
  NAND2_X1 U16081 ( .A1(n19326), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12814) );
  OAI211_X1 U16082 ( .C1(n12816), .C2(n19487), .A(n12815), .B(n12814), .ZN(
        n12817) );
  AOI211_X1 U16083 ( .C1(n16624), .C2(n12870), .A(n12818), .B(n12817), .ZN(
        n12825) );
  NOR2_X1 U16084 ( .A1(n15925), .A2(n12819), .ZN(n12822) );
  NAND2_X1 U16085 ( .A1(n15924), .A2(n19486), .ZN(n12820) );
  OAI211_X1 U16086 ( .C1(n19486), .C2(n15925), .A(n12820), .B(n19494), .ZN(
        n12821) );
  MUX2_X1 U16087 ( .A(n12822), .B(n12821), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n12823) );
  INV_X1 U16088 ( .A(n12823), .ZN(n12824) );
  OAI211_X1 U16089 ( .C1(n19491), .C2(n10013), .A(n12825), .B(n12824), .ZN(
        P2_U3044) );
  AND2_X1 U16090 ( .A1(n19151), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U16091 ( .A1(n13008), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12826) );
  AOI22_X1 U16092 ( .A1(n12998), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n20152), .B2(n20166), .ZN(n12827) );
  NAND2_X1 U16093 ( .A1(n14570), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12944) );
  XNOR2_X1 U16094 ( .A(n12943), .B(n12944), .ZN(n12833) );
  NAND2_X1 U16095 ( .A1(n12998), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12829) );
  NAND2_X1 U16096 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20159), .ZN(
        n19819) );
  NAND2_X1 U16097 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20166), .ZN(
        n19848) );
  NAND2_X1 U16098 ( .A1(n19819), .A2(n19848), .ZN(n19631) );
  NAND2_X1 U16099 ( .A1(n20152), .A2(n19631), .ZN(n19850) );
  NAND2_X1 U16100 ( .A1(n12829), .A2(n19850), .ZN(n12830) );
  NAND2_X1 U16101 ( .A1(n12833), .A2(n12832), .ZN(n12946) );
  OR2_X1 U16102 ( .A1(n12833), .A2(n12832), .ZN(n12834) );
  NAND2_X1 U16103 ( .A1(n12835), .A2(n10041), .ZN(n12836) );
  INV_X1 U16104 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n15476) );
  MUX2_X1 U16105 ( .A(n15476), .B(n19492), .S(n15537), .Z(n12837) );
  OAI21_X1 U16106 ( .B1(n20153), .B2(n15539), .A(n12837), .ZN(P2_U2886) );
  NAND2_X1 U16107 ( .A1(n19514), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12838) );
  AND4_X1 U16108 ( .A1(n10305), .A2(n12838), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19670), .ZN(n12839) );
  MUX2_X1 U16109 ( .A(n19347), .B(n12840), .S(n9726), .Z(n12841) );
  OAI21_X1 U16110 ( .B1(n20161), .B2(n15539), .A(n12841), .ZN(P2_U2887) );
  INV_X1 U16111 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12843) );
  INV_X2 U16112 ( .A(n19424), .ZN(n19459) );
  AOI22_X1 U16113 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n19459), .B1(n19454), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n12842) );
  OAI21_X1 U16114 ( .B1(n12843), .B2(n19425), .A(n12842), .ZN(P2_U2929) );
  INV_X1 U16115 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U16116 ( .A1(n19454), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U16117 ( .B1(n15546), .B2(n19425), .A(n12844), .ZN(P2_U2923) );
  INV_X1 U16118 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U16119 ( .A1(n19454), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12845) );
  OAI21_X1 U16120 ( .B1(n13912), .B2(n19425), .A(n12845), .ZN(P2_U2933) );
  INV_X1 U16121 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U16122 ( .A1(n19454), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12846) );
  OAI21_X1 U16123 ( .B1(n20871), .B2(n19425), .A(n12846), .ZN(P2_U2925) );
  AOI22_X1 U16124 ( .A1(n19454), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12847) );
  OAI21_X1 U16125 ( .B1(n12848), .B2(n19425), .A(n12847), .ZN(P2_U2926) );
  INV_X1 U16126 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20897) );
  AOI22_X1 U16127 ( .A1(n19454), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12849) );
  OAI21_X1 U16128 ( .B1(n20897), .B2(n19425), .A(n12849), .ZN(P2_U2931) );
  INV_X1 U16129 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U16130 ( .A1(n19454), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12850) );
  OAI21_X1 U16131 ( .B1(n13984), .B2(n19425), .A(n12850), .ZN(P2_U2932) );
  INV_X1 U16132 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U16133 ( .A1(n19454), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12851) );
  OAI21_X1 U16134 ( .B1(n14695), .B2(n19425), .A(n12851), .ZN(P2_U2921) );
  INV_X1 U16135 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13714) );
  AOI22_X1 U16136 ( .A1(n19454), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U16137 ( .B1(n13714), .B2(n19425), .A(n12852), .ZN(P2_U2935) );
  INV_X1 U16138 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n15571) );
  AOI22_X1 U16139 ( .A1(n19454), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12853) );
  OAI21_X1 U16140 ( .B1(n15571), .B2(n19425), .A(n12853), .ZN(P2_U2927) );
  AOI22_X1 U16141 ( .A1(n19454), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U16142 ( .B1(n12855), .B2(n19425), .A(n12854), .ZN(P2_U2924) );
  AOI22_X1 U16143 ( .A1(n19454), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12856) );
  OAI21_X1 U16144 ( .B1(n12857), .B2(n19425), .A(n12856), .ZN(P2_U2922) );
  INV_X1 U16145 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13866) );
  AOI22_X1 U16146 ( .A1(n19454), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12858) );
  OAI21_X1 U16147 ( .B1(n13866), .B2(n19425), .A(n12858), .ZN(P2_U2934) );
  NOR2_X1 U16148 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20184) );
  INV_X1 U16149 ( .A(n20184), .ZN(n12861) );
  NAND2_X1 U16150 ( .A1(n12861), .A2(n12860), .ZN(n12862) );
  INV_X1 U16151 ( .A(n13256), .ZN(n19480) );
  INV_X1 U16152 ( .A(n12871), .ZN(n12864) );
  INV_X1 U16153 ( .A(n20133), .ZN(n19153) );
  OR2_X1 U16154 ( .A1(n20152), .A2(n19153), .ZN(n20150) );
  NAND2_X1 U16155 ( .A1(n20150), .A2(n19151), .ZN(n12865) );
  INV_X1 U16156 ( .A(n12994), .ZN(n12867) );
  INV_X1 U16157 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n13249) );
  NAND2_X1 U16158 ( .A1(n13249), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12866) );
  NAND2_X1 U16159 ( .A1(n12867), .A2(n12866), .ZN(n19472) );
  OAI21_X1 U16160 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n13449), .ZN(n15461) );
  AOI22_X1 U16161 ( .A1(n19473), .A2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n19326), .B2(P2_REIP_REG_2__SCAN_IN), .ZN(n12868) );
  OAI21_X1 U16162 ( .B1(n19471), .B2(n15461), .A(n12868), .ZN(n12869) );
  AOI21_X1 U16163 ( .B1(n12870), .B2(n19475), .A(n12869), .ZN(n12875) );
  OR2_X2 U16164 ( .A1(n12871), .A2(n9739), .ZN(n16514) );
  INV_X1 U16165 ( .A(n16514), .ZN(n16538) );
  NAND3_X1 U16166 ( .A1(n12873), .A2(n16538), .A3(n12872), .ZN(n12874) );
  OAI211_X1 U16167 ( .C1(n13256), .C2(n10013), .A(n12875), .B(n12874), .ZN(
        P2_U3012) );
  INV_X1 U16168 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n20204) );
  NAND2_X1 U16169 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13243), .ZN(n16404) );
  AND2_X1 U16170 ( .A1(n12720), .A2(n13479), .ZN(n16159) );
  INV_X1 U16171 ( .A(n16208), .ZN(n13031) );
  OAI21_X1 U16172 ( .B1(n16159), .B2(n12786), .A(n13031), .ZN(n12876) );
  OAI21_X1 U16173 ( .B1(n14341), .B2(n12877), .A(n12876), .ZN(n12879) );
  INV_X1 U16174 ( .A(n12878), .ZN(n12892) );
  AOI21_X1 U16175 ( .B1(n12879), .B2(n16398), .A(n12892), .ZN(n12881) );
  INV_X1 U16176 ( .A(n13133), .ZN(n12880) );
  MUX2_X1 U16177 ( .A(n12881), .B(n12880), .S(n16187), .Z(n12889) );
  OR2_X1 U16178 ( .A1(n12882), .A2(n12720), .ZN(n12884) );
  INV_X1 U16179 ( .A(n12885), .ZN(n13025) );
  NAND2_X1 U16180 ( .A1(n13233), .A2(n13025), .ZN(n12886) );
  OAI211_X1 U16181 ( .C1(n13481), .C2(n11356), .A(n13028), .B(n12886), .ZN(
        n12887) );
  INV_X1 U16182 ( .A(n12887), .ZN(n12888) );
  NAND2_X1 U16183 ( .A1(n12889), .A2(n12888), .ZN(n13236) );
  AOI22_X1 U16184 ( .A1(n10118), .A2(P1_STATE2_REG_3__SCAN_IN), .B1(n13236), 
        .B2(n13132), .ZN(n12890) );
  OAI21_X1 U16185 ( .B1(n20204), .B2(n16404), .A(n12890), .ZN(n15341) );
  INV_X1 U16186 ( .A(n15341), .ZN(n14363) );
  INV_X1 U16187 ( .A(n12924), .ZN(n15332) );
  NAND2_X1 U16188 ( .A1(n13629), .A2(n15332), .ZN(n12907) );
  AND2_X1 U16189 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12895) );
  INV_X1 U16190 ( .A(n12895), .ZN(n12891) );
  NAND2_X1 U16191 ( .A1(n16159), .A2(n12891), .ZN(n12898) );
  OR2_X1 U16192 ( .A1(n13133), .A2(n12892), .ZN(n12922) );
  INV_X1 U16193 ( .A(n12893), .ZN(n12902) );
  NAND2_X1 U16194 ( .A1(n12902), .A2(n12894), .ZN(n12896) );
  AOI22_X1 U16195 ( .A1(n12922), .A2(n12896), .B1(n16159), .B2(n12895), .ZN(
        n12897) );
  MUX2_X1 U16196 ( .A(n12898), .B(n12897), .S(n11229), .Z(n12906) );
  NAND2_X1 U16197 ( .A1(n12893), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12899) );
  NAND2_X1 U16198 ( .A1(n12899), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12900) );
  NAND2_X1 U16199 ( .A1(n12901), .A2(n12900), .ZN(n12908) );
  NAND3_X1 U16200 ( .A1(n12924), .A2(n13135), .A3(n12908), .ZN(n12905) );
  NAND3_X1 U16201 ( .A1(n12922), .A2(n12903), .A3(n12902), .ZN(n12904) );
  NAND4_X1 U16202 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n13227) );
  AOI22_X1 U16203 ( .A1(n13227), .A2(n15334), .B1(n12930), .B2(n12908), .ZN(
        n12910) );
  NAND2_X1 U16204 ( .A1(n14363), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12909) );
  OAI21_X1 U16205 ( .B1(n14363), .B2(n12910), .A(n12909), .ZN(P1_U3469) );
  INV_X1 U16206 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15471) );
  OAI21_X1 U16207 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12912), .A(
        n12911), .ZN(n19489) );
  INV_X1 U16208 ( .A(n19489), .ZN(n12913) );
  NAND2_X1 U16209 ( .A1(n19475), .A2(n12913), .ZN(n12914) );
  NAND2_X1 U16210 ( .A1(n19326), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n19498) );
  OAI211_X1 U16211 ( .C1(n15471), .C2(n16541), .A(n12914), .B(n19498), .ZN(
        n12918) );
  OAI21_X1 U16212 ( .B1(n12955), .B2(n15469), .A(n12915), .ZN(n12916) );
  XOR2_X1 U16213 ( .A(n12916), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n19501) );
  NOR2_X1 U16214 ( .A1(n19501), .A2(n16514), .ZN(n12917) );
  AOI211_X1 U16215 ( .C1(n16530), .C2(n15471), .A(n12918), .B(n12917), .ZN(
        n12919) );
  OAI21_X1 U16216 ( .B1(n19492), .B2(n13256), .A(n12919), .ZN(P2_U3013) );
  NAND2_X1 U16217 ( .A1(n12611), .A2(n15332), .ZN(n12928) );
  NAND2_X1 U16218 ( .A1(n16159), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12921) );
  AND2_X1 U16219 ( .A1(n16159), .A2(n11223), .ZN(n15331) );
  INV_X1 U16220 ( .A(n15331), .ZN(n12920) );
  MUX2_X1 U16221 ( .A(n12921), .B(n12920), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12927) );
  XNOR2_X1 U16222 ( .A(n12893), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12923) );
  NAND2_X1 U16223 ( .A1(n12922), .A2(n12923), .ZN(n12926) );
  INV_X1 U16224 ( .A(n12923), .ZN(n12929) );
  NAND3_X1 U16225 ( .A1(n12924), .A2(n13135), .A3(n12929), .ZN(n12925) );
  NAND4_X1 U16226 ( .A1(n12928), .A2(n12927), .A3(n12926), .A4(n12925), .ZN(
        n13226) );
  INV_X1 U16227 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13732) );
  NOR2_X1 U16228 ( .A1(n20614), .A2(n13732), .ZN(n15337) );
  INV_X1 U16229 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14401) );
  INV_X1 U16230 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13731) );
  OAI22_X1 U16231 ( .A1(n14401), .A2(n13731), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15338) );
  INV_X1 U16232 ( .A(n15338), .ZN(n12931) );
  AOI222_X1 U16233 ( .A1(n13226), .A2(n15334), .B1(n15337), .B2(n12931), .C1(
        n12930), .C2(n12929), .ZN(n12933) );
  NAND2_X1 U16234 ( .A1(n14363), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12932) );
  OAI21_X1 U16235 ( .B1(n14363), .B2(n12933), .A(n12932), .ZN(P1_U3472) );
  NAND2_X1 U16236 ( .A1(n9750), .A2(n12994), .ZN(n12939) );
  NAND2_X1 U16237 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19989) );
  INV_X1 U16238 ( .A(n19989), .ZN(n12934) );
  AND2_X1 U16239 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12934), .ZN(
        n12995) );
  INV_X1 U16240 ( .A(n12995), .ZN(n12936) );
  NAND2_X1 U16241 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19879) );
  NAND2_X1 U16242 ( .A1(n19879), .A2(n20149), .ZN(n12935) );
  NAND2_X1 U16243 ( .A1(n12936), .A2(n12935), .ZN(n19632) );
  NOR2_X1 U16244 ( .A1(n20129), .A2(n19632), .ZN(n12937) );
  AOI21_X1 U16245 ( .B1(n12998), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12937), .ZN(n12938) );
  NAND2_X1 U16246 ( .A1(n12939), .A2(n12938), .ZN(n12941) );
  INV_X1 U16247 ( .A(n14570), .ZN(n14623) );
  INV_X1 U16248 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n14553) );
  NOR2_X1 U16249 ( .A1(n14623), .A2(n14553), .ZN(n12940) );
  NAND2_X1 U16250 ( .A1(n12941), .A2(n12940), .ZN(n13003) );
  OR2_X1 U16251 ( .A1(n12941), .A2(n12940), .ZN(n12942) );
  NAND2_X1 U16252 ( .A1(n13003), .A2(n12942), .ZN(n12948) );
  INV_X1 U16253 ( .A(n12943), .ZN(n16002) );
  NAND2_X1 U16254 ( .A1(n16002), .A2(n12944), .ZN(n12945) );
  NAND2_X1 U16255 ( .A1(n12946), .A2(n12945), .ZN(n12947) );
  NAND2_X1 U16256 ( .A1(n12948), .A2(n12947), .ZN(n12949) );
  NOR2_X1 U16257 ( .A1(n10013), .A2(n9726), .ZN(n12950) );
  AOI21_X1 U16258 ( .B1(P2_EBX_REG_2__SCAN_IN), .B2(n9726), .A(n12950), .ZN(
        n12951) );
  OAI21_X1 U16259 ( .B1(n20145), .B2(n15539), .A(n12951), .ZN(P2_U2885) );
  INV_X1 U16260 ( .A(n13283), .ZN(n13370) );
  NOR2_X1 U16261 ( .A1(n12952), .A2(n13370), .ZN(n12953) );
  XOR2_X1 U16262 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12953), .Z(
        n20265) );
  NAND4_X1 U16263 ( .A1(n15341), .A2(n13233), .A3(n15334), .A4(n20265), .ZN(
        n12954) );
  OAI21_X1 U16264 ( .B1(n15341), .B2(n20961), .A(n12954), .ZN(P1_U3468) );
  OAI21_X1 U16265 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19340), .A(
        n12955), .ZN(n19478) );
  OAI22_X1 U16266 ( .A1(n19500), .A2(n19478), .B1(n19494), .B2(n12964), .ZN(
        n12963) );
  OAI21_X1 U16267 ( .B1(n12958), .B2(n12957), .A(n12956), .ZN(n12959) );
  INV_X1 U16268 ( .A(n12959), .ZN(n19419) );
  AOI22_X1 U16269 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n12960), .B1(
        n10817), .B2(n12964), .ZN(n19474) );
  AOI22_X1 U16270 ( .A1(n16621), .A2(n19419), .B1(n16624), .B2(n19474), .ZN(
        n12961) );
  NAND2_X1 U16271 ( .A1(n19326), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n19476) );
  OAI211_X1 U16272 ( .C1(n19491), .C2(n19347), .A(n12961), .B(n19476), .ZN(
        n12962) );
  AOI211_X1 U16273 ( .C1(n12964), .C2(n15952), .A(n12963), .B(n12962), .ZN(
        n12965) );
  INV_X1 U16274 ( .A(n12965), .ZN(P2_U3046) );
  NAND2_X1 U16275 ( .A1(n13292), .A2(n13031), .ZN(n12966) );
  NOR2_X1 U16276 ( .A1(n12515), .A2(n12966), .ZN(n16185) );
  AOI21_X1 U16277 ( .B1(n16159), .B2(n13031), .A(n16185), .ZN(n12967) );
  NAND2_X1 U16278 ( .A1(n20297), .A2(n13472), .ZN(n20287) );
  NAND2_X1 U16279 ( .A1(n10118), .A2(n13243), .ZN(n20698) );
  INV_X1 U16280 ( .A(n20698), .ZN(n20296) );
  AOI22_X1 U16281 ( .A1(n20319), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n20318), .ZN(n12968) );
  OAI21_X1 U16282 ( .B1(n20287), .B2(n12969), .A(n12968), .ZN(P1_U2908) );
  INV_X1 U16283 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n20862) );
  AOI22_X1 U16284 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n12970) );
  OAI21_X1 U16285 ( .B1(n20862), .B2(n20287), .A(n12970), .ZN(P1_U2920) );
  INV_X1 U16286 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16287 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12971) );
  OAI21_X1 U16288 ( .B1(n12972), .B2(n20287), .A(n12971), .ZN(P1_U2909) );
  INV_X1 U16289 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16290 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n12973) );
  OAI21_X1 U16291 ( .B1(n12974), .B2(n20287), .A(n12973), .ZN(P1_U2919) );
  INV_X1 U16292 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U16293 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n12975) );
  OAI21_X1 U16294 ( .B1(n12976), .B2(n20287), .A(n12975), .ZN(P1_U2916) );
  INV_X1 U16295 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U16296 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U16297 ( .B1(n12978), .B2(n20287), .A(n12977), .ZN(P1_U2907) );
  INV_X1 U16298 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n12980) );
  AOI22_X1 U16299 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n12979) );
  OAI21_X1 U16300 ( .B1(n12980), .B2(n20287), .A(n12979), .ZN(P1_U2915) );
  INV_X1 U16301 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12982) );
  AOI22_X1 U16302 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12981) );
  OAI21_X1 U16303 ( .B1(n12982), .B2(n20287), .A(n12981), .ZN(P1_U2906) );
  INV_X1 U16304 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16305 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n12983) );
  OAI21_X1 U16306 ( .B1(n12984), .B2(n20287), .A(n12983), .ZN(P1_U2917) );
  AOI22_X1 U16307 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20296), .B1(n20318), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n12985) );
  OAI21_X1 U16308 ( .B1(n12090), .B2(n20287), .A(n12985), .ZN(P1_U2914) );
  INV_X1 U16309 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16310 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20296), .B1(n20318), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12986) );
  OAI21_X1 U16311 ( .B1(n12987), .B2(n20287), .A(n12986), .ZN(P1_U2911) );
  INV_X1 U16312 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U16313 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20296), .B1(n20318), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12988) );
  OAI21_X1 U16314 ( .B1(n12989), .B2(n20287), .A(n12988), .ZN(P1_U2912) );
  INV_X1 U16315 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12991) );
  AOI22_X1 U16316 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20296), .B1(n20318), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12990) );
  OAI21_X1 U16317 ( .B1(n12991), .B2(n20287), .A(n12990), .ZN(P1_U2910) );
  INV_X1 U16318 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16319 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20296), .B1(n20318), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n12992) );
  OAI21_X1 U16320 ( .B1(n12993), .B2(n20287), .A(n12992), .ZN(P1_U2913) );
  NAND2_X1 U16321 ( .A1(n13064), .A2(n12994), .ZN(n13000) );
  OAI21_X1 U16322 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12995), .A(
        n20152), .ZN(n12996) );
  AND2_X1 U16323 ( .A1(n12995), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20042) );
  NOR2_X1 U16324 ( .A1(n12996), .A2(n20042), .ZN(n12997) );
  AOI21_X1 U16325 ( .B1(n12998), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12997), .ZN(n12999) );
  INV_X1 U16326 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n14581) );
  NOR2_X1 U16327 ( .A1(n14623), .A2(n14581), .ZN(n13001) );
  NAND2_X1 U16328 ( .A1(n13005), .A2(n13001), .ZN(n13011) );
  NAND2_X1 U16329 ( .A1(n13005), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13006) );
  INV_X1 U16330 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14606) );
  NOR2_X1 U16331 ( .A1(n14623), .A2(n14606), .ZN(n13117) );
  NAND2_X1 U16332 ( .A1(n13123), .A2(n13117), .ZN(n13095) );
  NAND2_X1 U16333 ( .A1(n13008), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13009) );
  AND2_X1 U16334 ( .A1(n13007), .A2(n13009), .ZN(n13012) );
  INV_X1 U16335 ( .A(n13117), .ZN(n13010) );
  NAND3_X1 U16336 ( .A1(n13012), .A2(n13011), .A3(n13010), .ZN(n13013) );
  NAND2_X1 U16337 ( .A1(n13095), .A2(n13013), .ZN(n19391) );
  NAND2_X1 U16338 ( .A1(n13015), .A2(n13014), .ZN(n13017) );
  INV_X1 U16339 ( .A(n13019), .ZN(n13016) );
  AND2_X1 U16340 ( .A1(n13017), .A2(n13016), .ZN(n19467) );
  INV_X1 U16341 ( .A(n19467), .ZN(n19327) );
  MUX2_X1 U16342 ( .A(n10525), .B(n19327), .S(n15537), .Z(n13018) );
  OAI21_X1 U16343 ( .B1(n19391), .B2(n15539), .A(n13018), .ZN(P2_U2883) );
  XOR2_X1 U16344 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13095), .Z(n13023)
         );
  OR2_X1 U16345 ( .A1(n13020), .A2(n13019), .ZN(n13021) );
  NAND2_X1 U16346 ( .A1(n13021), .A2(n13068), .ZN(n16535) );
  MUX2_X1 U16347 ( .A(n16535), .B(n10576), .S(n9726), .Z(n13022) );
  OAI21_X1 U16348 ( .B1(n13023), .B2(n15539), .A(n13022), .ZN(P2_U2882) );
  AOI21_X1 U16349 ( .B1(n9828), .B2(n13732), .A(n13024), .ZN(n13088) );
  INV_X1 U16350 ( .A(n13088), .ZN(n13061) );
  NAND3_X1 U16351 ( .A1(n16187), .A2(n14359), .A3(n13479), .ZN(n13029) );
  NAND2_X1 U16352 ( .A1(n13479), .A2(n16208), .ZN(n13026) );
  NAND3_X1 U16353 ( .A1(n13026), .A2(n11356), .A3(n13025), .ZN(n13027) );
  NAND3_X1 U16354 ( .A1(n13029), .A2(n13028), .A3(n13027), .ZN(n13030) );
  NAND2_X1 U16355 ( .A1(n13030), .A2(n13132), .ZN(n13039) );
  OR2_X1 U16356 ( .A1(n13479), .A2(n13031), .ZN(n13473) );
  NAND3_X1 U16357 ( .A1(n12786), .A2(n16398), .A3(n13473), .ZN(n13033) );
  NAND2_X1 U16358 ( .A1(n13033), .A2(n13032), .ZN(n13035) );
  NAND2_X1 U16359 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NOR2_X1 U16360 ( .A1(n13044), .A2(n13577), .ZN(n13040) );
  OR3_X1 U16361 ( .A1(n13042), .A2(n13041), .A3(n13040), .ZN(n13043) );
  OAI22_X1 U16362 ( .A1(n12515), .A2(n13479), .B1(n11348), .B2(n13044), .ZN(
        n13045) );
  INV_X1 U16363 ( .A(n14342), .ZN(n14339) );
  NAND2_X1 U16364 ( .A1(n13438), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13047) );
  INV_X1 U16365 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U16366 ( .A1(n13172), .A2(n13141), .ZN(n13046) );
  NAND2_X1 U16367 ( .A1(n13047), .A2(n13046), .ZN(n13131) );
  INV_X1 U16368 ( .A(n13131), .ZN(n13048) );
  AOI21_X1 U16369 ( .B1(n14339), .B2(n13732), .A(n13048), .ZN(n13494) );
  INV_X1 U16370 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13049) );
  NOR2_X1 U16371 ( .A1(n20254), .A2(n13049), .ZN(n13087) );
  INV_X1 U16372 ( .A(n15293), .ZN(n13058) );
  NAND2_X1 U16373 ( .A1(n13054), .A2(n13133), .ZN(n20363) );
  INV_X1 U16374 ( .A(n20363), .ZN(n20389) );
  OR2_X1 U16375 ( .A1(n13054), .A2(n20349), .ZN(n13056) );
  OAI211_X1 U16376 ( .C1(n13052), .C2(n13472), .A(n13051), .B(n13050), .ZN(
        n13053) );
  NAND2_X1 U16377 ( .A1(n13732), .A2(n15232), .ZN(n13055) );
  NAND2_X1 U16378 ( .A1(n13056), .A2(n13055), .ZN(n20383) );
  AOI21_X1 U16379 ( .B1(n20389), .B2(n13732), .A(n20383), .ZN(n15319) );
  NOR3_X1 U16380 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20389), .A3(
        n15232), .ZN(n13057) );
  AOI21_X1 U16381 ( .B1(n13058), .B2(n15319), .A(n13057), .ZN(n13059) );
  AOI211_X1 U16382 ( .C1(n20374), .C2(n13494), .A(n13087), .B(n13059), .ZN(
        n13060) );
  OAI21_X1 U16383 ( .B1(n13061), .B2(n20385), .A(n13060), .ZN(P1_U3031) );
  INV_X1 U16384 ( .A(n19549), .ZN(n20137) );
  MUX2_X1 U16385 ( .A(P2_EBX_REG_3__SCAN_IN), .B(n13064), .S(n15537), .Z(
        n13065) );
  AOI21_X1 U16386 ( .B1(n20137), .B2(n15527), .A(n13065), .ZN(n13066) );
  INV_X1 U16387 ( .A(n13066), .ZN(P2_U2884) );
  AOI21_X1 U16388 ( .B1(n13069), .B2(n13068), .A(n13067), .ZN(n19314) );
  INV_X1 U16389 ( .A(n19314), .ZN(n14015) );
  INV_X1 U16390 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14632) );
  NOR2_X1 U16391 ( .A1(n13095), .A2(n14632), .ZN(n13070) );
  NAND2_X1 U16392 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13116) );
  OR2_X1 U16393 ( .A1(n13095), .A2(n13116), .ZN(n13090) );
  OAI211_X1 U16394 ( .C1(n13070), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n15527), .B(n13090), .ZN(n13072) );
  NAND2_X1 U16395 ( .A1(n9726), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n13071) );
  OAI211_X1 U16396 ( .C1(n14015), .C2(n9726), .A(n13072), .B(n13071), .ZN(
        P2_U2881) );
  INV_X1 U16397 ( .A(n13077), .ZN(n13073) );
  NAND2_X2 U16398 ( .A1(n14290), .A2(n13073), .ZN(n16283) );
  OAI21_X1 U16399 ( .B1(n13076), .B2(n13075), .A(n13074), .ZN(n13499) );
  INV_X1 U16400 ( .A(n13499), .ZN(n13140) );
  NAND2_X1 U16401 ( .A1(n14290), .A2(n13077), .ZN(n14293) );
  NAND2_X1 U16402 ( .A1(n13197), .A2(DATAI_0_), .ZN(n13079) );
  NAND2_X1 U16403 ( .A1(n14279), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13078) );
  AND2_X1 U16404 ( .A1(n13079), .A2(n13078), .ZN(n13286) );
  INV_X1 U16405 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20322) );
  OAI222_X1 U16406 ( .A1(n16283), .A2(n13140), .B1(n14293), .B2(n13286), .C1(
        n14290), .C2(n20322), .ZN(P1_U2904) );
  OAI21_X1 U16407 ( .B1(n13081), .B2(n13080), .A(n13184), .ZN(n14899) );
  NAND2_X1 U16408 ( .A1(n13197), .A2(DATAI_1_), .ZN(n13083) );
  NAND2_X1 U16409 ( .A1(n14279), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13082) );
  AND2_X1 U16410 ( .A1(n13083), .A2(n13082), .ZN(n13293) );
  INV_X1 U16411 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20317) );
  OAI222_X1 U16412 ( .A1(n14899), .A2(n16283), .B1(n14293), .B2(n13293), .C1(
        n14290), .C2(n20317), .ZN(P1_U2903) );
  INV_X1 U16413 ( .A(n20350), .ZN(n15134) );
  INV_X1 U16414 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13084) );
  AOI21_X1 U16415 ( .B1(n15134), .B2(n13085), .A(n13084), .ZN(n13086) );
  AOI211_X1 U16416 ( .C1(n13088), .C2(n20356), .A(n13087), .B(n13086), .ZN(
        n13089) );
  OAI21_X1 U16417 ( .B1(n13140), .B2(n15147), .A(n13089), .ZN(P1_U2999) );
  XOR2_X1 U16418 ( .A(n13090), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13094)
         );
  NOR2_X1 U16419 ( .A1(n13091), .A2(n13067), .ZN(n13092) );
  OR2_X1 U16420 ( .A1(n13099), .A2(n13092), .ZN(n19299) );
  MUX2_X1 U16421 ( .A(n19299), .B(n10630), .S(n9726), .Z(n13093) );
  OAI21_X1 U16422 ( .B1(n13094), .B2(n15539), .A(n13093), .ZN(P2_U2880) );
  NOR2_X1 U16423 ( .A1(n13095), .A2(n13116), .ZN(n13096) );
  AND2_X1 U16424 ( .A1(n13096), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n13097) );
  NAND2_X1 U16425 ( .A1(n13097), .A2(n13115), .ZN(n13114) );
  OAI211_X1 U16426 ( .C1(n13097), .C2(n13115), .A(n13114), .B(n15527), .ZN(
        n13102) );
  NOR2_X1 U16427 ( .A1(n13099), .A2(n13098), .ZN(n13100) );
  NOR2_X1 U16428 ( .A1(n13105), .A2(n13100), .ZN(n19290) );
  NAND2_X1 U16429 ( .A1(n19290), .A2(n15537), .ZN(n13101) );
  OAI211_X1 U16430 ( .C1(n15537), .C2(n13103), .A(n13102), .B(n13101), .ZN(
        P2_U2879) );
  XNOR2_X1 U16431 ( .A(n13114), .B(n13119), .ZN(n13109) );
  OR2_X1 U16432 ( .A1(n13105), .A2(n13104), .ZN(n13106) );
  NAND2_X1 U16433 ( .A1(n13106), .A2(n13110), .ZN(n19279) );
  MUX2_X1 U16434 ( .A(n19279), .B(n13107), .S(n9726), .Z(n13108) );
  OAI21_X1 U16435 ( .B1(n13109), .B2(n15539), .A(n13108), .ZN(P2_U2878) );
  NAND2_X1 U16436 ( .A1(n13111), .A2(n13110), .ZN(n13113) );
  INV_X1 U16437 ( .A(n13268), .ZN(n13112) );
  NAND2_X1 U16438 ( .A1(n13113), .A2(n13112), .ZN(n19268) );
  NOR2_X1 U16439 ( .A1(n13114), .A2(n13119), .ZN(n13125) );
  INV_X1 U16440 ( .A(n13120), .ZN(n13124) );
  NOR2_X1 U16441 ( .A1(n10167), .A2(n13116), .ZN(n13118) );
  AND2_X1 U16442 ( .A1(n13118), .A2(n13117), .ZN(n13121) );
  INV_X1 U16443 ( .A(n13192), .ZN(n13190) );
  OAI211_X1 U16444 ( .C1(n13125), .C2(n13124), .A(n13190), .B(n15527), .ZN(
        n13127) );
  NAND2_X1 U16445 ( .A1(n9726), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13126) );
  OAI211_X1 U16446 ( .C1(n19268), .C2(n9726), .A(n13127), .B(n13126), .ZN(
        P2_U2877) );
  OAI21_X1 U16447 ( .B1(n14308), .B2(n13731), .A(n14238), .ZN(n13128) );
  INV_X1 U16448 ( .A(n13128), .ZN(n13130) );
  MUX2_X1 U16449 ( .A(n13168), .B(n13438), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n13129) );
  NAND2_X1 U16450 ( .A1(n13130), .A2(n13129), .ZN(n13165) );
  XNOR2_X1 U16451 ( .A(n13165), .B(n13131), .ZN(n13167) );
  XNOR2_X1 U16452 ( .A(n13167), .B(n14341), .ZN(n15320) );
  NAND3_X1 U16453 ( .A1(n13133), .A2(n13132), .A3(n16187), .ZN(n13139) );
  INV_X1 U16454 ( .A(n13134), .ZN(n13137) );
  NAND4_X1 U16455 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n14308), .ZN(
        n13138) );
  INV_X1 U16456 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20820) );
  OAI222_X1 U16457 ( .A1(n15320), .A2(n14936), .B1(n20282), .B2(n20820), .C1(
        n14939), .C2(n14899), .ZN(P1_U2871) );
  INV_X1 U16458 ( .A(n13494), .ZN(n13142) );
  OAI222_X1 U16459 ( .A1(n13142), .A2(n14936), .B1(n20282), .B2(n13141), .C1(
        n14939), .C2(n13140), .ZN(P1_U2872) );
  OAI21_X1 U16460 ( .B1(n13145), .B2(n13144), .A(n13143), .ZN(n13407) );
  NAND2_X1 U16461 ( .A1(n13197), .A2(DATAI_3_), .ZN(n13147) );
  NAND2_X1 U16462 ( .A1(n14279), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13146) );
  AND2_X1 U16463 ( .A1(n13147), .A2(n13146), .ZN(n13312) );
  INV_X1 U16464 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20313) );
  OAI222_X1 U16465 ( .A1(n13407), .A2(n16283), .B1(n14293), .B2(n13312), .C1(
        n14290), .C2(n20313), .ZN(P1_U2901) );
  INV_X1 U16466 ( .A(n16398), .ZN(n20697) );
  AND2_X1 U16467 ( .A1(n20700), .A2(n20697), .ZN(n13148) );
  NOR2_X2 U16468 ( .A1(n20345), .A2(n13292), .ZN(n20333) );
  NAND2_X1 U16469 ( .A1(n13197), .A2(DATAI_7_), .ZN(n13151) );
  NAND2_X1 U16470 ( .A1(n14279), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13150) );
  AND2_X1 U16471 ( .A1(n13151), .A2(n13150), .ZN(n13615) );
  INV_X1 U16472 ( .A(n13615), .ZN(n14964) );
  NAND2_X1 U16473 ( .A1(n20333), .A2(n14964), .ZN(n13203) );
  AOI22_X1 U16474 ( .A1(n20346), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13152) );
  NAND2_X1 U16475 ( .A1(n13203), .A2(n13152), .ZN(P1_U2959) );
  INV_X1 U16476 ( .A(n13293), .ZN(n14982) );
  NAND2_X1 U16477 ( .A1(n20333), .A2(n14982), .ZN(n13216) );
  AOI22_X1 U16478 ( .A1(n20346), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13153) );
  NAND2_X1 U16479 ( .A1(n13216), .A2(n13153), .ZN(P1_U2938) );
  NAND2_X1 U16480 ( .A1(n13197), .A2(DATAI_4_), .ZN(n13155) );
  NAND2_X1 U16481 ( .A1(n14279), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13154) );
  AND2_X1 U16482 ( .A1(n13155), .A2(n13154), .ZN(n13579) );
  INV_X1 U16483 ( .A(n13579), .ZN(n16281) );
  NAND2_X1 U16484 ( .A1(n20333), .A2(n16281), .ZN(n13220) );
  AOI22_X1 U16485 ( .A1(n20346), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13156) );
  NAND2_X1 U16486 ( .A1(n13220), .A2(n13156), .ZN(P1_U2941) );
  NAND2_X1 U16487 ( .A1(n13197), .A2(DATAI_2_), .ZN(n13158) );
  NAND2_X1 U16488 ( .A1(n14279), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13157) );
  AND2_X1 U16489 ( .A1(n13158), .A2(n13157), .ZN(n13307) );
  INV_X1 U16490 ( .A(n13307), .ZN(n14978) );
  NAND2_X1 U16491 ( .A1(n20333), .A2(n14978), .ZN(n13218) );
  AOI22_X1 U16492 ( .A1(n20346), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13159) );
  NAND2_X1 U16493 ( .A1(n13218), .A2(n13159), .ZN(P1_U2939) );
  INV_X1 U16494 ( .A(n13312), .ZN(n14975) );
  NAND2_X1 U16495 ( .A1(n20333), .A2(n14975), .ZN(n13210) );
  AOI22_X1 U16496 ( .A1(n20346), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13160) );
  NAND2_X1 U16497 ( .A1(n13210), .A2(n13160), .ZN(P1_U2940) );
  INV_X1 U16498 ( .A(n13286), .ZN(n14986) );
  NAND2_X1 U16499 ( .A1(n20333), .A2(n14986), .ZN(n13214) );
  AOI22_X1 U16500 ( .A1(n20346), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U16501 ( .A1(n13214), .A2(n13161), .ZN(P1_U2937) );
  INV_X1 U16502 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n14283) );
  INV_X1 U16503 ( .A(n20333), .ZN(n13164) );
  INV_X1 U16504 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13162) );
  NOR2_X1 U16505 ( .A1(n13197), .A2(n13162), .ZN(n13163) );
  AOI21_X1 U16506 ( .B1(DATAI_15_), .B2(n13197), .A(n13163), .ZN(n14284) );
  INV_X1 U16507 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20291) );
  OAI222_X1 U16508 ( .A1(n13200), .A2(n14283), .B1(n13164), .B2(n14284), .C1(
        n13181), .C2(n20291), .ZN(P1_U2967) );
  INV_X1 U16509 ( .A(n13165), .ZN(n13166) );
  AOI21_X2 U16510 ( .B1(n13167), .B2(n14308), .A(n13166), .ZN(n13222) );
  MUX2_X1 U16511 ( .A(n13168), .B(n14335), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13171) );
  NAND2_X1 U16512 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14341), .ZN(
        n13169) );
  AND2_X1 U16513 ( .A1(n14238), .A2(n13169), .ZN(n13170) );
  NAND2_X1 U16514 ( .A1(n13171), .A2(n13170), .ZN(n13221) );
  NAND2_X1 U16515 ( .A1(n13222), .A2(n13221), .ZN(n13174) );
  MUX2_X1 U16516 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13173) );
  OAI21_X1 U16517 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14342), .A(
        n13173), .ZN(n13178) );
  INV_X1 U16518 ( .A(n13174), .ZN(n13176) );
  NAND2_X1 U16519 ( .A1(n13176), .A2(n13175), .ZN(n13345) );
  INV_X1 U16520 ( .A(n13345), .ZN(n13177) );
  AOI21_X1 U16521 ( .B1(n13174), .B2(n13178), .A(n13177), .ZN(n20373) );
  INV_X1 U16522 ( .A(n20373), .ZN(n13179) );
  INV_X1 U16523 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n14880) );
  OAI222_X1 U16524 ( .A1(n13179), .A2(n14936), .B1(n20282), .B2(n14880), .C1(
        n14939), .C2(n13407), .ZN(P1_U2869) );
  INV_X1 U16525 ( .A(P1_UWORD_REG_12__SCAN_IN), .ZN(n20783) );
  MUX2_X1 U16526 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n14279), .Z(
        n14948) );
  NAND2_X1 U16527 ( .A1(n20333), .A2(n14948), .ZN(n20341) );
  NAND2_X1 U16528 ( .A1(n20346), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13180) );
  OAI211_X1 U16529 ( .C1(n13181), .C2(n20783), .A(n20341), .B(n13180), .ZN(
        P1_U2949) );
  INV_X1 U16530 ( .A(n13182), .ZN(n13183) );
  AOI21_X1 U16531 ( .B1(n13185), .B2(n13184), .A(n13183), .ZN(n13571) );
  INV_X1 U16532 ( .A(n13571), .ZN(n13224) );
  INV_X1 U16533 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20315) );
  OAI222_X1 U16534 ( .A1(n13224), .A2(n16283), .B1(n14293), .B2(n13307), .C1(
        n14290), .C2(n20315), .ZN(P1_U2902) );
  INV_X1 U16535 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20304) );
  MUX2_X1 U16536 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n14279), .Z(
        n14960) );
  NAND2_X1 U16537 ( .A1(n20333), .A2(n14960), .ZN(n13208) );
  NAND2_X1 U16538 ( .A1(n20345), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13186) );
  OAI211_X1 U16539 ( .C1(n20304), .C2(n13200), .A(n13208), .B(n13186), .ZN(
        P1_U2960) );
  NAND2_X1 U16540 ( .A1(n13271), .A2(n13187), .ZN(n13188) );
  NAND2_X1 U16541 ( .A1(n13399), .A2(n13188), .ZN(n19255) );
  NOR2_X1 U16542 ( .A1(n13190), .A2(n13189), .ZN(n13194) );
  AND2_X1 U16543 ( .A1(n13267), .A2(n13193), .ZN(n13191) );
  INV_X1 U16544 ( .A(n13467), .ZN(n13464) );
  OAI211_X1 U16545 ( .C1(n13194), .C2(n13193), .A(n13464), .B(n15527), .ZN(
        n13196) );
  NAND2_X1 U16546 ( .A1(n9726), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13195) );
  OAI211_X1 U16547 ( .C1(n19255), .C2(n9726), .A(n13196), .B(n13195), .ZN(
        P2_U2875) );
  NAND2_X1 U16548 ( .A1(n13197), .A2(DATAI_5_), .ZN(n13199) );
  NAND2_X1 U16549 ( .A1(n14279), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13198) );
  AND2_X1 U16550 ( .A1(n13199), .A2(n13198), .ZN(n13357) );
  INV_X1 U16551 ( .A(n13357), .ZN(n14972) );
  NAND2_X1 U16552 ( .A1(n20333), .A2(n14972), .ZN(n13212) );
  AOI22_X1 U16553 ( .A1(n20323), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13201) );
  NAND2_X1 U16554 ( .A1(n13212), .A2(n13201), .ZN(P1_U2942) );
  AOI22_X1 U16555 ( .A1(n20323), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13202) );
  NAND2_X1 U16556 ( .A1(n13203), .A2(n13202), .ZN(P1_U2944) );
  NAND2_X1 U16557 ( .A1(n20333), .A2(n14968), .ZN(n13206) );
  AOI22_X1 U16558 ( .A1(n20323), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16559 ( .A1(n13206), .A2(n13204), .ZN(P1_U2943) );
  AOI22_X1 U16560 ( .A1(n20323), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U16561 ( .A1(n13206), .A2(n13205), .ZN(P1_U2958) );
  AOI22_X1 U16562 ( .A1(n20323), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13207) );
  NAND2_X1 U16563 ( .A1(n13208), .A2(n13207), .ZN(P1_U2945) );
  AOI22_X1 U16564 ( .A1(n20323), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16565 ( .A1(n13210), .A2(n13209), .ZN(P1_U2955) );
  AOI22_X1 U16566 ( .A1(n20323), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U16567 ( .A1(n13212), .A2(n13211), .ZN(P1_U2957) );
  AOI22_X1 U16568 ( .A1(n20323), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13213) );
  NAND2_X1 U16569 ( .A1(n13214), .A2(n13213), .ZN(P1_U2952) );
  AOI22_X1 U16570 ( .A1(n20323), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13215) );
  NAND2_X1 U16571 ( .A1(n13216), .A2(n13215), .ZN(P1_U2953) );
  AOI22_X1 U16572 ( .A1(n20323), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13217) );
  NAND2_X1 U16573 ( .A1(n13218), .A2(n13217), .ZN(P1_U2954) );
  AOI22_X1 U16574 ( .A1(n20323), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13219) );
  NAND2_X1 U16575 ( .A1(n13220), .A2(n13219), .ZN(P1_U2956) );
  OR2_X1 U16576 ( .A1(n13222), .A2(n13221), .ZN(n13223) );
  NAND2_X1 U16577 ( .A1(n13174), .A2(n13223), .ZN(n20391) );
  INV_X1 U16578 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13225) );
  OAI222_X1 U16579 ( .A1(n20391), .A2(n14936), .B1(n20282), .B2(n13225), .C1(
        n14939), .C2(n13224), .ZN(P1_U2870) );
  NAND2_X1 U16580 ( .A1(n20204), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13238) );
  INV_X1 U16581 ( .A(n13238), .ZN(n13228) );
  MUX2_X1 U16582 ( .A(n13226), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16163), .Z(n16158) );
  AOI22_X1 U16583 ( .A1(n13228), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n16158), .B2(n20614), .ZN(n13230) );
  MUX2_X1 U16584 ( .A(n13227), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16163), .Z(n16171) );
  AOI22_X1 U16585 ( .A1(n13228), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20614), .B2(n16171), .ZN(n13229) );
  NOR2_X1 U16586 ( .A1(n13230), .A2(n13229), .ZN(n16181) );
  INV_X1 U16587 ( .A(n13231), .ZN(n13232) );
  NAND2_X1 U16588 ( .A1(n16181), .A2(n13232), .ZN(n13244) );
  AOI21_X1 U16589 ( .B1(n20265), .B2(n13233), .A(n16163), .ZN(n13234) );
  NOR2_X1 U16590 ( .A1(n13234), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13235) );
  OAI21_X1 U16591 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13236), .A(
        n13235), .ZN(n13237) );
  OAI21_X1 U16592 ( .B1(n13238), .B2(n20961), .A(n13237), .ZN(n16180) );
  INV_X1 U16593 ( .A(n16180), .ZN(n13242) );
  NAND3_X1 U16594 ( .A1(n13244), .A2(n20204), .A3(n13242), .ZN(n13241) );
  INV_X1 U16595 ( .A(n16404), .ZN(n13240) );
  AOI21_X1 U16596 ( .B1(n13241), .B2(n13240), .A(n13239), .ZN(n20400) );
  AND3_X1 U16597 ( .A1(n13244), .A2(n13243), .A3(n13242), .ZN(n16189) );
  INV_X1 U16598 ( .A(n11787), .ZN(n13492) );
  NAND2_X1 U16599 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n16406), .ZN(n13265) );
  INV_X1 U16600 ( .A(n13265), .ZN(n13245) );
  OAI22_X1 U16601 ( .A1(n13246), .A2(n20559), .B1(n13492), .B2(n13245), .ZN(
        n13247) );
  OAI21_X1 U16602 ( .B1(n16189), .B2(n13247), .A(n13349), .ZN(n13248) );
  OAI21_X1 U16603 ( .B1(n13349), .B2(n20549), .A(n13248), .ZN(P1_U3478) );
  OR2_X1 U16604 ( .A1(n19549), .A2(n13249), .ZN(n19882) );
  NAND3_X1 U16605 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20159), .ZN(n19909) );
  OAI21_X1 U16606 ( .B1(n19882), .B2(n19672), .A(n19909), .ZN(n13255) );
  NOR2_X1 U16607 ( .A1(n20166), .A2(n19909), .ZN(n19961) );
  INV_X1 U16608 ( .A(n19961), .ZN(n13250) );
  AND2_X1 U16609 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13250), .ZN(n13251) );
  NAND2_X1 U16610 ( .A1(n13252), .A2(n13251), .ZN(n13258) );
  OAI211_X1 U16611 ( .C1(n19961), .C2(n19670), .A(n13258), .B(n19999), .ZN(
        n13253) );
  INV_X1 U16612 ( .A(n13253), .ZN(n13254) );
  INV_X1 U16613 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13261) );
  NOR2_X2 U16614 ( .A1(n19851), .A2(n19672), .ZN(n19963) );
  AOI22_X1 U16615 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19531), .ZN(n19946) );
  NOR2_X2 U16616 ( .A1(n19877), .A2(n19672), .ZN(n19984) );
  AOI22_X1 U16617 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19531), .ZN(n20051) );
  AOI22_X1 U16618 ( .A1(n19963), .A2(n20045), .B1(n19984), .B2(n19941), .ZN(
        n13260) );
  OAI21_X1 U16619 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19909), .A(n20182), 
        .ZN(n13257) );
  AND2_X1 U16620 ( .A1(n13258), .A2(n13257), .ZN(n19962) );
  NOR2_X2 U16621 ( .A1(n19382), .A2(n19913), .ZN(n20043) );
  NAND2_X1 U16622 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19999), .ZN(n19533) );
  AND2_X1 U16623 ( .A1(n10973), .A2(n19525), .ZN(n20041) );
  AOI22_X1 U16624 ( .A1(n19962), .A2(n20043), .B1(n19961), .B2(n20041), .ZN(
        n13259) );
  OAI211_X1 U16625 ( .C1(n19966), .C2(n13261), .A(n13260), .B(n13259), .ZN(
        P2_U3159) );
  AOI22_X1 U16626 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19531), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19532), .ZN(n19935) );
  AOI22_X1 U16627 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19531), .ZN(n20034) );
  AOI22_X1 U16628 ( .A1(n19963), .A2(n20031), .B1(n19984), .B2(n19979), .ZN(
        n13263) );
  NOR2_X2 U16629 ( .A1(n19395), .A2(n19913), .ZN(n20030) );
  NOR2_X2 U16630 ( .A1(n11197), .A2(n19533), .ZN(n20029) );
  AOI22_X1 U16631 ( .A1(n19962), .A2(n20030), .B1(n19961), .B2(n20029), .ZN(
        n13262) );
  OAI211_X1 U16632 ( .C1(n19966), .C2(n13264), .A(n13263), .B(n13262), .ZN(
        P2_U3157) );
  NAND2_X1 U16633 ( .A1(n13349), .A2(n13265), .ZN(n13368) );
  NAND2_X1 U16634 ( .A1(n13349), .A2(n20561), .ZN(n13360) );
  NAND2_X1 U16635 ( .A1(n12607), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13633) );
  XOR2_X1 U16636 ( .A(n9748), .B(n13633), .Z(n13266) );
  OAI222_X1 U16637 ( .A1(n13368), .A2(n13568), .B1(n13360), .B2(n13266), .C1(
        n20788), .C2(n13349), .ZN(P1_U3476) );
  XNOR2_X1 U16638 ( .A(n13192), .B(n13267), .ZN(n13274) );
  OR2_X1 U16639 ( .A1(n13269), .A2(n13268), .ZN(n13270) );
  AND2_X1 U16640 ( .A1(n13271), .A2(n13270), .ZN(n16500) );
  INV_X1 U16641 ( .A(n16500), .ZN(n16588) );
  MUX2_X1 U16642 ( .A(n16588), .B(n13272), .S(n9726), .Z(n13273) );
  OAI21_X1 U16643 ( .B1(n13274), .B2(n15539), .A(n13273), .ZN(P2_U2876) );
  INV_X1 U16644 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13275) );
  NOR2_X1 U16645 ( .A1(n20254), .A2(n13275), .ZN(n15322) );
  AOI21_X1 U16646 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n15322), .ZN(n13276) );
  OAI21_X1 U16647 ( .B1(n20361), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13276), .ZN(n13277) );
  INV_X1 U16648 ( .A(n13277), .ZN(n13281) );
  OR2_X1 U16649 ( .A1(n13278), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n15318) );
  NAND3_X1 U16650 ( .A1(n15318), .A2(n20356), .A3(n13279), .ZN(n13280) );
  OAI211_X1 U16651 ( .C1(n14899), .C2(n15147), .A(n13281), .B(n13280), .ZN(
        P1_U2998) );
  AOI22_X1 U16652 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13576), .B1(DATAI_24_), 
        .B2(n13575), .ZN(n20566) );
  NAND2_X1 U16653 ( .A1(n9748), .A2(n13361), .ZN(n14099) );
  NAND2_X1 U16654 ( .A1(n12607), .A2(n13659), .ZN(n13369) );
  OR2_X1 U16655 ( .A1(n14099), .A2(n13369), .ZN(n13830) );
  AOI22_X1 U16656 ( .A1(DATAI_16_), .A2(n13575), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n13576), .ZN(n20460) );
  INV_X1 U16657 ( .A(n20460), .ZN(n20563) );
  NOR2_X1 U16658 ( .A1(n13578), .A2(n13282), .ZN(n20554) );
  INV_X1 U16659 ( .A(n20554), .ZN(n14137) );
  NAND2_X1 U16660 ( .A1(n12611), .A2(n13283), .ZN(n14105) );
  NAND2_X1 U16661 ( .A1(n11787), .A2(n13284), .ZN(n13630) );
  OAI21_X1 U16662 ( .B1(n14105), .B2(n13630), .A(n13594), .ZN(n13285) );
  AOI22_X1 U16663 ( .A1(n13285), .A2(n13917), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14100), .ZN(n13593) );
  OAI22_X1 U16664 ( .A1(n14137), .A2(n13594), .B1(n13593), .B2(n14169), .ZN(
        n13287) );
  AOI21_X1 U16665 ( .B1(n20414), .B2(n20563), .A(n13287), .ZN(n13291) );
  INV_X1 U16666 ( .A(n13633), .ZN(n13288) );
  NAND2_X1 U16667 ( .A1(n13288), .A2(n20561), .ZN(n13319) );
  NOR2_X1 U16668 ( .A1(n14099), .A2(n13319), .ZN(n13289) );
  OAI21_X1 U16669 ( .B1(n13289), .B2(n14100), .A(n20557), .ZN(n13596) );
  NAND2_X1 U16670 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13290) );
  OAI211_X1 U16671 ( .C1(n20566), .C2(n14106), .A(n13291), .B(n13290), .ZN(
        P1_U3153) );
  AOI22_X1 U16672 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n13576), .B1(DATAI_25_), 
        .B2(n13575), .ZN(n20572) );
  AOI22_X1 U16673 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n13576), .B1(DATAI_17_), 
        .B2(n13575), .ZN(n20464) );
  INV_X1 U16674 ( .A(n20464), .ZN(n20569) );
  NOR2_X1 U16675 ( .A1(n13578), .A2(n13292), .ZN(n20568) );
  INV_X1 U16676 ( .A(n20568), .ZN(n14116) );
  OAI22_X1 U16677 ( .A1(n14116), .A2(n13594), .B1(n13593), .B2(n14173), .ZN(
        n13294) );
  AOI21_X1 U16678 ( .B1(n20414), .B2(n20569), .A(n13294), .ZN(n13296) );
  NAND2_X1 U16679 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13295) );
  OAI211_X1 U16680 ( .C1(n20572), .C2(n14106), .A(n13296), .B(n13295), .ZN(
        P1_U3154) );
  AOI22_X1 U16681 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13576), .B1(DATAI_29_), 
        .B2(n13575), .ZN(n20596) );
  AOI22_X1 U16682 ( .A1(DATAI_21_), .A2(n13575), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13576), .ZN(n20480) );
  INV_X1 U16683 ( .A(n20480), .ZN(n20593) );
  NOR2_X1 U16684 ( .A1(n13578), .A2(n13297), .ZN(n20592) );
  INV_X1 U16685 ( .A(n20592), .ZN(n14120) );
  OAI22_X1 U16686 ( .A1(n14120), .A2(n13594), .B1(n13593), .B2(n14189), .ZN(
        n13298) );
  AOI21_X1 U16687 ( .B1(n20414), .B2(n20593), .A(n13298), .ZN(n13300) );
  NAND2_X1 U16688 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n13299) );
  OAI211_X1 U16689 ( .C1(n20596), .C2(n14106), .A(n13300), .B(n13299), .ZN(
        P1_U3158) );
  INV_X1 U16690 ( .A(n20484), .ZN(n20599) );
  OAI22_X1 U16691 ( .A1(n14165), .A2(n13593), .B1(n13594), .B2(n13780), .ZN(
        n13301) );
  AOI21_X1 U16692 ( .B1(n20414), .B2(n20599), .A(n13301), .ZN(n13303) );
  NAND2_X1 U16693 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n13302) );
  OAI211_X1 U16694 ( .C1(n20602), .C2(n14106), .A(n13303), .B(n13302), .ZN(
        P1_U3159) );
  AOI22_X1 U16695 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n13576), .B1(DATAI_31_), 
        .B2(n13575), .ZN(n20613) );
  AOI22_X1 U16696 ( .A1(DATAI_23_), .A2(n13575), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n13576), .ZN(n20492) );
  INV_X1 U16697 ( .A(n20492), .ZN(n20607) );
  NOR2_X1 U16698 ( .A1(n13578), .A2(n14940), .ZN(n20606) );
  INV_X1 U16699 ( .A(n20606), .ZN(n14128) );
  OAI22_X1 U16700 ( .A1(n14128), .A2(n13594), .B1(n13593), .B2(n14181), .ZN(
        n13304) );
  AOI21_X1 U16701 ( .B1(n20414), .B2(n20607), .A(n13304), .ZN(n13306) );
  NAND2_X1 U16702 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n13305) );
  OAI211_X1 U16703 ( .C1(n20613), .C2(n14106), .A(n13306), .B(n13305), .ZN(
        P1_U3160) );
  AOI22_X1 U16704 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13576), .B1(DATAI_26_), 
        .B2(n13575), .ZN(n20578) );
  AOI22_X1 U16705 ( .A1(DATAI_18_), .A2(n13575), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n13576), .ZN(n20468) );
  INV_X1 U16706 ( .A(n20468), .ZN(n20575) );
  INV_X1 U16707 ( .A(n20574), .ZN(n14124) );
  OAI22_X1 U16708 ( .A1(n14124), .A2(n13594), .B1(n13593), .B2(n14185), .ZN(
        n13308) );
  AOI21_X1 U16709 ( .B1(n20414), .B2(n20575), .A(n13308), .ZN(n13310) );
  NAND2_X1 U16710 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n13309) );
  OAI211_X1 U16711 ( .C1(n20578), .C2(n14106), .A(n13310), .B(n13309), .ZN(
        P1_U3155) );
  AOI22_X1 U16712 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13576), .B1(DATAI_27_), 
        .B2(n13575), .ZN(n20584) );
  AOI22_X1 U16713 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n13576), .B1(DATAI_19_), 
        .B2(n13575), .ZN(n20472) );
  INV_X1 U16714 ( .A(n20472), .ZN(n20581) );
  NOR2_X1 U16715 ( .A1(n13578), .A2(n13311), .ZN(n20580) );
  INV_X1 U16716 ( .A(n20580), .ZN(n14112) );
  OAI22_X1 U16717 ( .A1(n14112), .A2(n13594), .B1(n13593), .B2(n14177), .ZN(
        n13313) );
  AOI21_X1 U16718 ( .B1(n20414), .B2(n20581), .A(n13313), .ZN(n13315) );
  NAND2_X1 U16719 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n13314) );
  OAI211_X1 U16720 ( .C1(n20584), .C2(n14106), .A(n13315), .B(n13314), .ZN(
        P1_U3156) );
  INV_X1 U16721 ( .A(n13369), .ZN(n13627) );
  NAND2_X1 U16722 ( .A1(n13660), .A2(n13627), .ZN(n13741) );
  INV_X1 U16723 ( .A(n13631), .ZN(n13316) );
  NAND2_X1 U16724 ( .A1(n13316), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13588) );
  OAI21_X1 U16725 ( .B1(n20520), .B2(n13630), .A(n13588), .ZN(n13317) );
  AOI22_X1 U16726 ( .A1(n13317), .A2(n20561), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13320), .ZN(n13587) );
  OAI22_X1 U16727 ( .A1(n14128), .A2(n13588), .B1(n13587), .B2(n14181), .ZN(
        n13318) );
  AOI21_X1 U16728 ( .B1(n13773), .B2(n20607), .A(n13318), .ZN(n13323) );
  NOR2_X1 U16729 ( .A1(n20525), .A2(n13319), .ZN(n13321) );
  OAI21_X1 U16730 ( .B1(n13321), .B2(n13320), .A(n20557), .ZN(n13590) );
  NAND2_X1 U16731 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n13322) );
  OAI211_X1 U16732 ( .C1(n20613), .C2(n14048), .A(n13323), .B(n13322), .ZN(
        P1_U3128) );
  OAI22_X1 U16733 ( .A1(n14165), .A2(n13587), .B1(n13780), .B2(n13588), .ZN(
        n13324) );
  AOI21_X1 U16734 ( .B1(n13773), .B2(n20599), .A(n13324), .ZN(n13326) );
  NAND2_X1 U16735 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n13325) );
  OAI211_X1 U16736 ( .C1(n20602), .C2(n14048), .A(n13326), .B(n13325), .ZN(
        P1_U3127) );
  OAI22_X1 U16737 ( .A1(n14120), .A2(n13588), .B1(n13587), .B2(n14189), .ZN(
        n13327) );
  AOI21_X1 U16738 ( .B1(n13773), .B2(n20593), .A(n13327), .ZN(n13329) );
  NAND2_X1 U16739 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n13328) );
  OAI211_X1 U16740 ( .C1(n20596), .C2(n14048), .A(n13329), .B(n13328), .ZN(
        P1_U3126) );
  OAI22_X1 U16741 ( .A1(n14112), .A2(n13588), .B1(n13587), .B2(n14177), .ZN(
        n13330) );
  AOI21_X1 U16742 ( .B1(n13773), .B2(n20581), .A(n13330), .ZN(n13332) );
  NAND2_X1 U16743 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n13331) );
  OAI211_X1 U16744 ( .C1(n20584), .C2(n14048), .A(n13332), .B(n13331), .ZN(
        P1_U3124) );
  OAI22_X1 U16745 ( .A1(n14124), .A2(n13588), .B1(n13587), .B2(n14185), .ZN(
        n13333) );
  AOI21_X1 U16746 ( .B1(n13773), .B2(n20575), .A(n13333), .ZN(n13335) );
  NAND2_X1 U16747 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n13334) );
  OAI211_X1 U16748 ( .C1(n20578), .C2(n14048), .A(n13335), .B(n13334), .ZN(
        P1_U3123) );
  OAI22_X1 U16749 ( .A1(n14116), .A2(n13588), .B1(n13587), .B2(n14173), .ZN(
        n13336) );
  AOI21_X1 U16750 ( .B1(n13773), .B2(n20569), .A(n13336), .ZN(n13338) );
  NAND2_X1 U16751 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13337) );
  OAI211_X1 U16752 ( .C1(n20572), .C2(n14048), .A(n13338), .B(n13337), .ZN(
        P1_U3122) );
  OAI22_X1 U16753 ( .A1(n14137), .A2(n13588), .B1(n13587), .B2(n14169), .ZN(
        n13339) );
  AOI21_X1 U16754 ( .B1(n13773), .B2(n20563), .A(n13339), .ZN(n13341) );
  NAND2_X1 U16755 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13340) );
  OAI211_X1 U16756 ( .C1(n20566), .C2(n14048), .A(n13341), .B(n13340), .ZN(
        P1_U3121) );
  MUX2_X1 U16757 ( .A(n13168), .B(n14335), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13343) );
  NAND2_X1 U16758 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n14341), .ZN(
        n13342) );
  AND2_X1 U16759 ( .A1(n13345), .A2(n13344), .ZN(n13346) );
  OR2_X1 U16760 ( .A1(n13346), .A2(n9824), .ZN(n20367) );
  XOR2_X1 U16761 ( .A(n13143), .B(n13347), .Z(n20355) );
  INV_X1 U16762 ( .A(n20355), .ZN(n13359) );
  INV_X1 U16763 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13348) );
  OAI222_X1 U16764 ( .A1(n20367), .A2(n14936), .B1(n14939), .B2(n13359), .C1(
        n20282), .C2(n13348), .ZN(P1_U2868) );
  NOR2_X1 U16765 ( .A1(n12607), .A2(n20818), .ZN(n13363) );
  AOI21_X1 U16766 ( .B1(n20818), .B2(n12607), .A(n13363), .ZN(n13350) );
  OAI222_X1 U16767 ( .A1(n13368), .A2(n12613), .B1(n13360), .B2(n13350), .C1(
        n16166), .C2(n13349), .ZN(P1_U3477) );
  OR2_X1 U16768 ( .A1(n13354), .A2(n13353), .ZN(n13355) );
  AND2_X1 U16769 ( .A1(n13352), .A2(n13355), .ZN(n20284) );
  INV_X1 U16770 ( .A(n20284), .ZN(n13358) );
  OAI222_X1 U16771 ( .A1(n13358), .A2(n16283), .B1(n14293), .B2(n13357), .C1(
        n13356), .C2(n14290), .ZN(P1_U2899) );
  INV_X1 U16772 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20311) );
  OAI222_X1 U16773 ( .A1(n14290), .A2(n20311), .B1(n14293), .B2(n13579), .C1(
        n16283), .C2(n13359), .ZN(P1_U2900) );
  INV_X1 U16774 ( .A(n13629), .ZN(n14884) );
  INV_X1 U16775 ( .A(n13360), .ZN(n13366) );
  INV_X1 U16776 ( .A(n13361), .ZN(n13362) );
  OR2_X1 U16777 ( .A1(n20496), .A2(n13633), .ZN(n13375) );
  INV_X1 U16778 ( .A(n13363), .ZN(n20524) );
  OR2_X1 U16779 ( .A1(n14099), .A2(n20524), .ZN(n20556) );
  OR2_X1 U16780 ( .A1(n11797), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13364) );
  NAND4_X1 U16781 ( .A1(n13375), .A2(n20556), .A3(n20525), .A4(n13364), .ZN(
        n13365) );
  AOI22_X1 U16782 ( .A1(n13366), .A2(n13365), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20400), .ZN(n13367) );
  OAI21_X1 U16783 ( .B1(n14884), .B2(n13368), .A(n13367), .ZN(P1_U3475) );
  INV_X1 U16784 ( .A(n20584), .ZN(n20469) );
  INV_X1 U16785 ( .A(n20493), .ZN(n13371) );
  OAI21_X1 U16786 ( .B1(n13371), .B2(n13630), .A(n13581), .ZN(n13373) );
  AOI22_X1 U16787 ( .A1(n13373), .A2(n20561), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13377), .ZN(n13580) );
  OAI22_X1 U16788 ( .A1(n14112), .A2(n13581), .B1(n13580), .B2(n14177), .ZN(
        n13372) );
  AOI21_X1 U16789 ( .B1(n13583), .B2(n20469), .A(n13372), .ZN(n13379) );
  INV_X1 U16790 ( .A(n13373), .ZN(n13374) );
  NAND3_X1 U16791 ( .A1(n13375), .A2(n20561), .A3(n13374), .ZN(n13376) );
  OAI211_X1 U16792 ( .C1(n13917), .C2(n13377), .A(n13376), .B(n20557), .ZN(
        n13584) );
  NAND2_X1 U16793 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n13378) );
  OAI211_X1 U16794 ( .C1(n20472), .C2(n13668), .A(n13379), .B(n13378), .ZN(
        P1_U3092) );
  INV_X1 U16795 ( .A(n20613), .ZN(n20487) );
  OAI22_X1 U16796 ( .A1(n14128), .A2(n13581), .B1(n13580), .B2(n14181), .ZN(
        n13380) );
  AOI21_X1 U16797 ( .B1(n13583), .B2(n20487), .A(n13380), .ZN(n13382) );
  NAND2_X1 U16798 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n13381) );
  OAI211_X1 U16799 ( .C1(n20492), .C2(n13668), .A(n13382), .B(n13381), .ZN(
        P1_U3096) );
  INV_X1 U16800 ( .A(n20578), .ZN(n20465) );
  OAI22_X1 U16801 ( .A1(n14124), .A2(n13581), .B1(n13580), .B2(n14185), .ZN(
        n13383) );
  AOI21_X1 U16802 ( .B1(n13583), .B2(n20465), .A(n13383), .ZN(n13385) );
  NAND2_X1 U16803 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n13384) );
  OAI211_X1 U16804 ( .C1(n20468), .C2(n13668), .A(n13385), .B(n13384), .ZN(
        P1_U3091) );
  INV_X1 U16805 ( .A(n20572), .ZN(n20461) );
  OAI22_X1 U16806 ( .A1(n14116), .A2(n13581), .B1(n13580), .B2(n14173), .ZN(
        n13386) );
  AOI21_X1 U16807 ( .B1(n13583), .B2(n20461), .A(n13386), .ZN(n13388) );
  NAND2_X1 U16808 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13387) );
  OAI211_X1 U16809 ( .C1(n20464), .C2(n13668), .A(n13388), .B(n13387), .ZN(
        P1_U3090) );
  INV_X1 U16810 ( .A(n20596), .ZN(n20477) );
  OAI22_X1 U16811 ( .A1(n14120), .A2(n13581), .B1(n13580), .B2(n14189), .ZN(
        n13389) );
  AOI21_X1 U16812 ( .B1(n13583), .B2(n20477), .A(n13389), .ZN(n13391) );
  NAND2_X1 U16813 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n13390) );
  OAI211_X1 U16814 ( .C1(n20480), .C2(n13668), .A(n13391), .B(n13390), .ZN(
        P1_U3094) );
  OAI22_X1 U16815 ( .A1(n14165), .A2(n13580), .B1(n13581), .B2(n13780), .ZN(
        n13392) );
  AOI21_X1 U16816 ( .B1(n13583), .B2(n20481), .A(n13392), .ZN(n13394) );
  NAND2_X1 U16817 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n13393) );
  OAI211_X1 U16818 ( .C1(n20484), .C2(n13668), .A(n13394), .B(n13393), .ZN(
        P1_U3095) );
  INV_X1 U16819 ( .A(n20566), .ZN(n20457) );
  OAI22_X1 U16820 ( .A1(n14137), .A2(n13581), .B1(n13580), .B2(n14169), .ZN(
        n13395) );
  AOI21_X1 U16821 ( .B1(n13583), .B2(n20457), .A(n13395), .ZN(n13397) );
  NAND2_X1 U16822 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13396) );
  OAI211_X1 U16823 ( .C1(n20460), .C2(n13668), .A(n13397), .B(n13396), .ZN(
        P1_U3089) );
  XNOR2_X1 U16824 ( .A(n13467), .B(n13465), .ZN(n13402) );
  NAND2_X1 U16825 ( .A1(n13399), .A2(n13398), .ZN(n13400) );
  NAND2_X1 U16826 ( .A1(n13461), .A2(n13400), .ZN(n16558) );
  INV_X1 U16827 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13558) );
  MUX2_X1 U16828 ( .A(n16558), .B(n13558), .S(n9726), .Z(n13401) );
  OAI21_X1 U16829 ( .B1(n13402), .B2(n15539), .A(n13401), .ZN(P2_U2874) );
  OR2_X1 U16830 ( .A1(n13405), .A2(n13404), .ZN(n13406) );
  NAND2_X1 U16831 ( .A1(n13403), .A2(n13406), .ZN(n20376) );
  INV_X1 U16832 ( .A(n13407), .ZN(n14888) );
  INV_X1 U16833 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14890) );
  NOR2_X1 U16834 ( .A1(n20254), .A2(n14890), .ZN(n20372) );
  AOI21_X1 U16835 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20372), .ZN(n13408) );
  OAI21_X1 U16836 ( .B1(n20361), .B2(n14879), .A(n13408), .ZN(n13409) );
  AOI21_X1 U16837 ( .B1(n14888), .B2(n14067), .A(n13409), .ZN(n13410) );
  OAI21_X1 U16838 ( .B1(n20376), .B2(n20203), .A(n13410), .ZN(P1_U2996) );
  XOR2_X1 U16839 ( .A(n20147), .B(n15465), .Z(n19406) );
  NAND2_X1 U16840 ( .A1(n13412), .A2(n13411), .ZN(n13413) );
  NAND2_X1 U16841 ( .A1(n13414), .A2(n13413), .ZN(n20157) );
  XNOR2_X1 U16842 ( .A(n20153), .B(n20157), .ZN(n19411) );
  NAND2_X1 U16843 ( .A1(n19548), .A2(n19419), .ZN(n19418) );
  NAND2_X1 U16844 ( .A1(n19411), .A2(n19418), .ZN(n19410) );
  OAI21_X1 U16845 ( .B1(n20157), .B2(n19573), .A(n19410), .ZN(n19405) );
  NAND2_X1 U16846 ( .A1(n19406), .A2(n19405), .ZN(n19404) );
  OAI21_X1 U16847 ( .B1(n15465), .B2(n20147), .A(n19404), .ZN(n19398) );
  INV_X1 U16848 ( .A(n13415), .ZN(n13416) );
  XNOR2_X1 U16849 ( .A(n13417), .B(n13416), .ZN(n20135) );
  XOR2_X1 U16850 ( .A(n20135), .B(n19549), .Z(n19399) );
  NAND2_X1 U16851 ( .A1(n19398), .A2(n19399), .ZN(n19397) );
  NAND2_X1 U16852 ( .A1(n19549), .A2(n20135), .ZN(n13422) );
  INV_X1 U16853 ( .A(n13419), .ZN(n13420) );
  OAI21_X1 U16854 ( .B1(n13418), .B2(n13421), .A(n13420), .ZN(n19322) );
  INV_X1 U16855 ( .A(n19322), .ZN(n13433) );
  AOI21_X1 U16856 ( .B1(n19397), .B2(n13422), .A(n13433), .ZN(n19392) );
  XNOR2_X1 U16857 ( .A(n19392), .B(n19391), .ZN(n13435) );
  NAND2_X1 U16858 ( .A1(n13424), .A2(n13423), .ZN(n13425) );
  NAND2_X1 U16859 ( .A1(n13425), .A2(n16682), .ZN(n13428) );
  NAND2_X1 U16860 ( .A1(n20188), .A2(n13426), .ZN(n13427) );
  NAND2_X1 U16861 ( .A1(n19387), .A2(n10300), .ZN(n15577) );
  NOR2_X1 U16862 ( .A1(n13430), .A2(n10305), .ZN(n13431) );
  INV_X1 U16863 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19449) );
  OAI22_X1 U16864 ( .A1(n19422), .A2(n19526), .B1(n19449), .B2(n19387), .ZN(
        n13432) );
  AOI21_X1 U16865 ( .B1(n13433), .B2(n19416), .A(n13432), .ZN(n13434) );
  OAI21_X1 U16866 ( .B1(n13435), .B2(n19390), .A(n13434), .ZN(P2_U2915) );
  AOI21_X1 U16867 ( .B1(n13437), .B2(n13352), .A(n11837), .ZN(n13729) );
  INV_X1 U16868 ( .A(n13729), .ZN(n20243) );
  INV_X1 U16869 ( .A(n14332), .ZN(n14326) );
  INV_X1 U16870 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20286) );
  NAND2_X1 U16871 ( .A1(n14326), .A2(n20286), .ZN(n13441) );
  NAND2_X1 U16872 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13439) );
  OAI211_X1 U16873 ( .C1(n14341), .C2(P1_EBX_REG_5__SCAN_IN), .A(n14335), .B(
        n13439), .ZN(n13440) );
  MUX2_X1 U16874 ( .A(n13168), .B(n14335), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13443) );
  NAND2_X1 U16875 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14341), .ZN(
        n13442) );
  XOR2_X1 U16876 ( .A(n16386), .B(n13617), .Z(n20246) );
  INV_X1 U16877 ( .A(n20282), .ZN(n20707) );
  AOI22_X1 U16878 ( .A1(n20246), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13444) );
  OAI21_X1 U16879 ( .B1(n20243), .B2(n14939), .A(n13444), .ZN(P1_U2866) );
  OAI222_X1 U16880 ( .A1(n20243), .A2(n16283), .B1(n14293), .B2(n13445), .C1(
        n20307), .C2(n14290), .ZN(P1_U2898) );
  XNOR2_X1 U16881 ( .A(n13448), .B(n13447), .ZN(n16632) );
  AOI21_X1 U16882 ( .B1(n13603), .B2(n13449), .A(n13505), .ZN(n13601) );
  NAND2_X1 U16883 ( .A1(n16530), .A2(n13601), .ZN(n13450) );
  NAND2_X1 U16884 ( .A1(n19326), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16633) );
  OAI211_X1 U16885 ( .C1(n13603), .C2(n16541), .A(n13450), .B(n16633), .ZN(
        n13453) );
  XNOR2_X1 U16886 ( .A(n10816), .B(n13451), .ZN(n16637) );
  NOR2_X1 U16887 ( .A1(n16637), .A2(n19464), .ZN(n13452) );
  AOI211_X1 U16888 ( .C1(n19480), .C2(n13064), .A(n13453), .B(n13452), .ZN(
        n13454) );
  OAI21_X1 U16889 ( .B1(n16632), .B2(n16514), .A(n13454), .ZN(P2_U3011) );
  NAND2_X1 U16890 ( .A1(n20349), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20390) );
  NAND2_X1 U16891 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13455) );
  OAI211_X1 U16892 ( .C1(n20361), .C2(n13565), .A(n20390), .B(n13455), .ZN(
        n13459) );
  INV_X1 U16893 ( .A(n13457), .ZN(n20386) );
  NOR3_X1 U16894 ( .A1(n20387), .A2(n20386), .A3(n20203), .ZN(n13458) );
  AOI211_X1 U16895 ( .C1(n13571), .C2(n14067), .A(n13459), .B(n13458), .ZN(
        n13460) );
  INV_X1 U16896 ( .A(n13460), .ZN(P1_U2997) );
  AOI21_X1 U16897 ( .B1(n13462), .B2(n13461), .A(n13820), .ZN(n19243) );
  INV_X1 U16898 ( .A(n19243), .ZN(n15734) );
  NOR2_X1 U16899 ( .A1(n13464), .A2(n13463), .ZN(n13469) );
  AND2_X1 U16900 ( .A1(n13468), .A2(n13465), .ZN(n13466) );
  AND2_X2 U16901 ( .A1(n13467), .A2(n13466), .ZN(n13907) );
  INV_X1 U16902 ( .A(n13907), .ZN(n13817) );
  OAI211_X1 U16903 ( .C1(n13469), .C2(n13468), .A(n15527), .B(n13817), .ZN(
        n13471) );
  NAND2_X1 U16904 ( .A1(n9726), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n13470) );
  OAI211_X1 U16905 ( .C1(n15734), .C2(n9726), .A(n13471), .B(n13470), .ZN(
        P2_U2873) );
  AND2_X1 U16906 ( .A1(n13496), .A2(n13472), .ZN(n13486) );
  AND2_X1 U16907 ( .A1(n16398), .A2(n20818), .ZN(n16184) );
  NAND2_X1 U16908 ( .A1(n13473), .A2(n16184), .ZN(n13484) );
  INV_X1 U16909 ( .A(n13484), .ZN(n13474) );
  NOR3_X1 U16910 ( .A1(n16406), .A2(P1_STATE2_REG_1__SCAN_IN), .A3(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n16403) );
  NAND2_X1 U16911 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n10118), .ZN(n13476) );
  OAI21_X1 U16912 ( .B1(n13476), .B2(n13475), .A(n20254), .ZN(n13477) );
  AOI21_X1 U16913 ( .B1(n16403), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n13477), 
        .ZN(n13478) );
  INV_X1 U16914 ( .A(n14892), .ZN(n14845) );
  NAND2_X1 U16915 ( .A1(n20271), .A2(n14845), .ZN(n14847) );
  INV_X1 U16916 ( .A(n14847), .ZN(n20252) );
  NAND2_X1 U16917 ( .A1(n13479), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13483) );
  NOR2_X1 U16918 ( .A1(n13483), .A2(n16184), .ZN(n13480) );
  INV_X1 U16919 ( .A(n13481), .ZN(n13482) );
  NAND2_X1 U16920 ( .A1(n13496), .A2(n13482), .ZN(n20262) );
  AND2_X1 U16921 ( .A1(n13484), .A2(n13483), .ZN(n13485) );
  NAND2_X1 U16922 ( .A1(n20263), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13491) );
  NOR2_X2 U16923 ( .A1(n14892), .A2(n16406), .ZN(n20269) );
  XNOR2_X1 U16924 ( .A(n13488), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14414) );
  NAND2_X1 U16925 ( .A1(n14414), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13489) );
  OAI21_X1 U16926 ( .B1(n20269), .B2(n20221), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13490) );
  OAI211_X1 U16927 ( .C1(n20262), .C2(n13492), .A(n13491), .B(n13490), .ZN(
        n13493) );
  AOI21_X1 U16928 ( .B1(n20253), .B2(n13494), .A(n13493), .ZN(n13501) );
  AND2_X1 U16929 ( .A1(n13496), .A2(n13495), .ZN(n13498) );
  NAND2_X1 U16930 ( .A1(n13499), .A2(n20272), .ZN(n13500) );
  OAI211_X1 U16931 ( .C1(n20252), .C2(n13049), .A(n13501), .B(n13500), .ZN(
        P1_U2840) );
  AOI21_X1 U16932 ( .B1(n16542), .B2(n13504), .A(n13530), .ZN(n16529) );
  INV_X1 U16933 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15443) );
  INV_X1 U16934 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15705) );
  INV_X1 U16935 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15745) );
  INV_X1 U16936 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16511) );
  INV_X1 U16937 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n19228) );
  INV_X1 U16938 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15690) );
  INV_X1 U16939 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16487) );
  INV_X1 U16940 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15630) );
  INV_X1 U16941 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15386) );
  INV_X1 U16942 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U16943 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14429) );
  OAI22_X1 U16944 ( .A1(n19151), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n19355) );
  OAI22_X1 U16945 ( .A1(n19151), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15471), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15468) );
  AND2_X1 U16946 ( .A1(n19355), .A2(n15468), .ZN(n15459) );
  NAND2_X1 U16947 ( .A1(n15459), .A2(n15461), .ZN(n13599) );
  NOR2_X1 U16948 ( .A1(n13601), .A2(n13599), .ZN(n19330) );
  OAI21_X1 U16949 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13505), .A(
        n13504), .ZN(n19470) );
  NAND2_X1 U16950 ( .A1(n19330), .A2(n19470), .ZN(n13528) );
  NAND2_X1 U16951 ( .A1(n15347), .A2(n13528), .ZN(n13506) );
  XNOR2_X1 U16952 ( .A(n16529), .B(n13506), .ZN(n13507) );
  NAND4_X1 U16953 ( .A1(n20182), .A2(n19151), .A3(n13249), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20056) );
  INV_X1 U16954 ( .A(n20056), .ZN(n19316) );
  NAND2_X1 U16955 ( .A1(n13507), .A2(n19316), .ZN(n13527) );
  OAI21_X1 U16956 ( .B1(n13419), .B2(n13509), .A(n13508), .ZN(n13510) );
  INV_X1 U16957 ( .A(n13510), .ZN(n19389) );
  NOR2_X1 U16958 ( .A1(n20183), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n13521) );
  INV_X1 U16959 ( .A(n13521), .ZN(n13511) );
  NOR2_X1 U16960 ( .A1(n20068), .A2(n13511), .ZN(n16684) );
  AND3_X1 U16961 ( .A1(n10043), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n13511), .ZN(
        n13512) );
  NAND2_X1 U16962 ( .A1(n20188), .A2(n13512), .ZN(n19308) );
  NOR2_X1 U16963 ( .A1(n19670), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19704) );
  INV_X1 U16964 ( .A(n19704), .ZN(n20052) );
  NOR2_X1 U16965 ( .A1(n20059), .A2(n20052), .ZN(n16681) );
  NAND2_X1 U16966 ( .A1(n19304), .A2(n20056), .ZN(n13513) );
  OR2_X1 U16967 ( .A1(n16681), .A2(n13513), .ZN(n13514) );
  NAND2_X1 U16968 ( .A1(n19305), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19306) );
  INV_X1 U16969 ( .A(n16684), .ZN(n16410) );
  NAND2_X1 U16970 ( .A1(n16411), .A2(n16410), .ZN(n13518) );
  NOR2_X1 U16971 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13521), .ZN(n13515) );
  NAND2_X1 U16972 ( .A1(n13516), .A2(n13515), .ZN(n13517) );
  AOI22_X1 U16973 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19351), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19342), .ZN(n13519) );
  OAI211_X1 U16974 ( .C1(n19308), .C2(n13520), .A(n13519), .B(n19304), .ZN(
        n13525) );
  AND2_X1 U16975 ( .A1(n10043), .A2(n13521), .ZN(n13522) );
  NAND2_X1 U16976 ( .A1(n20188), .A2(n13522), .ZN(n19346) );
  OAI22_X1 U16977 ( .A1(n19346), .A2(n16535), .B1(n19305), .B2(n13523), .ZN(
        n13524) );
  AOI211_X1 U16978 ( .C1(n19389), .C2(n19339), .A(n13525), .B(n13524), .ZN(
        n13526) );
  NAND2_X1 U16979 ( .A1(n13527), .A2(n13526), .ZN(P2_U2850) );
  AOI21_X1 U16980 ( .B1(n16511), .B2(n13533), .A(n9807), .ZN(n16495) );
  AOI21_X1 U16981 ( .B1(n16520), .B2(n13531), .A(n13534), .ZN(n19275) );
  AOI21_X1 U16982 ( .B1(n16528), .B2(n13529), .A(n13532), .ZN(n19295) );
  NOR2_X1 U16983 ( .A1(n16529), .A2(n13528), .ZN(n19311) );
  OAI21_X1 U16984 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13530), .A(
        n13529), .ZN(n19312) );
  NAND2_X1 U16985 ( .A1(n19311), .A2(n19312), .ZN(n19294) );
  NOR2_X1 U16986 ( .A1(n19295), .A2(n19294), .ZN(n19287) );
  OAI21_X1 U16987 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13532), .A(
        n13531), .ZN(n19288) );
  NAND2_X1 U16988 ( .A1(n19287), .A2(n19288), .ZN(n19274) );
  NOR2_X1 U16989 ( .A1(n19275), .A2(n19274), .ZN(n19260) );
  OAI21_X1 U16990 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13534), .A(
        n13533), .ZN(n19261) );
  NAND2_X1 U16991 ( .A1(n19260), .A2(n19261), .ZN(n13548) );
  NAND2_X1 U16992 ( .A1(n15347), .A2(n13548), .ZN(n13535) );
  XNOR2_X1 U16993 ( .A(n16495), .B(n13535), .ZN(n13546) );
  AOI21_X1 U16994 ( .B1(n13538), .B2(n13537), .A(n13536), .ZN(n19372) );
  INV_X1 U16995 ( .A(n19372), .ZN(n16586) );
  OAI21_X1 U16996 ( .B1(n11083), .B2(n19305), .A(n19304), .ZN(n13539) );
  AOI21_X1 U16997 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19351), .A(
        n13539), .ZN(n13540) );
  OAI21_X1 U16998 ( .B1(n19323), .B2(n16586), .A(n13540), .ZN(n13541) );
  INV_X1 U16999 ( .A(n13541), .ZN(n13543) );
  AOI22_X1 U17000 ( .A1(n19315), .A2(n16500), .B1(n19342), .B2(
        P2_EBX_REG_11__SCAN_IN), .ZN(n13542) );
  OAI211_X1 U17001 ( .C1(n13544), .C2(n19308), .A(n13543), .B(n13542), .ZN(
        n13545) );
  AOI21_X1 U17002 ( .B1(n13546), .B2(n19316), .A(n13545), .ZN(n13547) );
  INV_X1 U17003 ( .A(n13547), .ZN(P2_U2844) );
  AOI21_X1 U17004 ( .B1(n15745), .B2(n13549), .A(n14213), .ZN(n15746) );
  NOR2_X1 U17005 ( .A1(n16495), .A2(n13548), .ZN(n19252) );
  OAI21_X1 U17006 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9807), .A(
        n13549), .ZN(n19253) );
  NAND2_X1 U17007 ( .A1(n19252), .A2(n19253), .ZN(n14211) );
  NAND2_X1 U17008 ( .A1(n15347), .A2(n14211), .ZN(n13550) );
  XNOR2_X1 U17009 ( .A(n15746), .B(n13550), .ZN(n13551) );
  NAND2_X1 U17010 ( .A1(n13551), .A2(n19316), .ZN(n13562) );
  INV_X1 U17011 ( .A(n16558), .ZN(n13560) );
  OAI21_X1 U17012 ( .B1(n10891), .B2(n19305), .A(n19304), .ZN(n13552) );
  AOI21_X1 U17013 ( .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19351), .A(
        n13552), .ZN(n13557) );
  AOI21_X1 U17014 ( .B1(n13555), .B2(n13553), .A(n13554), .ZN(n19366) );
  NAND2_X1 U17015 ( .A1(n19339), .A2(n19366), .ZN(n13556) );
  OAI211_X1 U17016 ( .C1(n19324), .C2(n13558), .A(n13557), .B(n13556), .ZN(
        n13559) );
  AOI21_X1 U17017 ( .B1(n13560), .B2(n19315), .A(n13559), .ZN(n13561) );
  OAI211_X1 U17018 ( .C1(n19308), .C2(n13563), .A(n13562), .B(n13561), .ZN(
        P2_U2842) );
  NAND2_X1 U17019 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n14885) );
  NAND2_X1 U17020 ( .A1(n16239), .A2(n14885), .ZN(n13574) );
  AND2_X1 U17021 ( .A1(n13574), .A2(n14845), .ZN(n14891) );
  INV_X1 U17022 ( .A(n14891), .ZN(n13564) );
  NAND2_X1 U17023 ( .A1(n13564), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13573) );
  INV_X1 U17024 ( .A(n13565), .ZN(n13566) );
  AOI22_X1 U17025 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20269), .B1(
        n20221), .B2(n13566), .ZN(n13567) );
  OAI21_X1 U17026 ( .B1(n16272), .B2(n13225), .A(n13567), .ZN(n13570) );
  OAI22_X1 U17027 ( .A1(n20267), .A2(n20391), .B1(n13568), .B2(n20262), .ZN(
        n13569) );
  AOI211_X1 U17028 ( .C1(n13571), .C2(n20272), .A(n13570), .B(n13569), .ZN(
        n13572) );
  OAI211_X1 U17029 ( .C1(n13574), .C2(n13275), .A(n13573), .B(n13572), .ZN(
        P1_U2838) );
  AOI22_X1 U17030 ( .A1(DATAI_20_), .A2(n13575), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n13576), .ZN(n20476) );
  AOI22_X1 U17031 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13576), .B1(DATAI_28_), 
        .B2(n13575), .ZN(n20590) );
  INV_X1 U17032 ( .A(n20590), .ZN(n20473) );
  NOR2_X1 U17033 ( .A1(n13578), .A2(n13577), .ZN(n20586) );
  INV_X1 U17034 ( .A(n20586), .ZN(n14144) );
  OAI22_X1 U17035 ( .A1(n14144), .A2(n13581), .B1(n13580), .B2(n14196), .ZN(
        n13582) );
  AOI21_X1 U17036 ( .B1(n13583), .B2(n20473), .A(n13582), .ZN(n13586) );
  NAND2_X1 U17037 ( .A1(n13584), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n13585) );
  OAI211_X1 U17038 ( .C1(n20476), .C2(n13668), .A(n13586), .B(n13585), .ZN(
        P1_U3093) );
  INV_X1 U17039 ( .A(n20476), .ZN(n20587) );
  OAI22_X1 U17040 ( .A1(n14144), .A2(n13588), .B1(n13587), .B2(n14196), .ZN(
        n13589) );
  AOI21_X1 U17041 ( .B1(n13773), .B2(n20587), .A(n13589), .ZN(n13592) );
  NAND2_X1 U17042 ( .A1(n13590), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n13591) );
  OAI211_X1 U17043 ( .C1(n20590), .C2(n14048), .A(n13592), .B(n13591), .ZN(
        P1_U3125) );
  OAI22_X1 U17044 ( .A1(n14144), .A2(n13594), .B1(n13593), .B2(n14196), .ZN(
        n13595) );
  AOI21_X1 U17045 ( .B1(n20414), .B2(n20587), .A(n13595), .ZN(n13598) );
  NAND2_X1 U17046 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n13597) );
  OAI211_X1 U17047 ( .C1(n20590), .C2(n14106), .A(n13598), .B(n13597), .ZN(
        P1_U3157) );
  INV_X1 U17048 ( .A(n19349), .ZN(n19328) );
  NAND2_X1 U17049 ( .A1(n15347), .A2(n13599), .ZN(n13600) );
  XNOR2_X1 U17050 ( .A(n13601), .B(n13600), .ZN(n13602) );
  NAND2_X1 U17051 ( .A1(n13602), .A2(n19316), .ZN(n13611) );
  INV_X1 U17052 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13604) );
  OAI22_X1 U17053 ( .A1(n19324), .A2(n13604), .B1(n13603), .B2(n19306), .ZN(
        n13605) );
  INV_X1 U17054 ( .A(n13605), .ZN(n13606) );
  OAI21_X1 U17055 ( .B1(n19308), .B2(n13607), .A(n13606), .ZN(n13609) );
  OAI22_X1 U17056 ( .A1(n11004), .A2(n19305), .B1(n19323), .B2(n20135), .ZN(
        n13608) );
  AOI211_X1 U17057 ( .C1(n13064), .C2(n19315), .A(n13609), .B(n13608), .ZN(
        n13610) );
  OAI211_X1 U17058 ( .C1(n19549), .C2(n19328), .A(n13611), .B(n13610), .ZN(
        P2_U2852) );
  NAND2_X1 U17059 ( .A1(n13436), .A2(n13613), .ZN(n13614) );
  AND2_X1 U17060 ( .A1(n13612), .A2(n13614), .ZN(n20234) );
  INV_X1 U17061 ( .A(n20234), .ZN(n13616) );
  OAI222_X1 U17062 ( .A1(n13616), .A2(n16283), .B1(n14293), .B2(n13615), .C1(
        n14290), .C2(n11833), .ZN(P1_U2897) );
  INV_X1 U17063 ( .A(n14939), .ZN(n20708) );
  NAND2_X1 U17064 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13618) );
  OAI211_X1 U17065 ( .C1(n14341), .C2(P1_EBX_REG_7__SCAN_IN), .A(n13438), .B(
        n13618), .ZN(n13619) );
  OAI21_X1 U17066 ( .B1(n14332), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13619), .ZN(
        n13620) );
  NAND2_X1 U17067 ( .A1(n13621), .A2(n13620), .ZN(n13622) );
  NAND2_X1 U17068 ( .A1(n13809), .A2(n13622), .ZN(n20229) );
  INV_X1 U17069 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13623) );
  OAI22_X1 U17070 ( .A1(n20229), .A2(n14936), .B1(n13623), .B2(n20282), .ZN(
        n13624) );
  AOI21_X1 U17071 ( .B1(n20234), .B2(n20708), .A(n13624), .ZN(n13625) );
  INV_X1 U17072 ( .A(n13625), .ZN(P1_U2865) );
  INV_X1 U17073 ( .A(n9748), .ZN(n13626) );
  INV_X1 U17074 ( .A(n20424), .ZN(n13628) );
  OR2_X1 U17075 ( .A1(n12611), .A2(n13629), .ZN(n14152) );
  INV_X1 U17076 ( .A(n13630), .ZN(n13632) );
  NOR2_X1 U17077 ( .A1(n13631), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13656) );
  AOI21_X1 U17078 ( .B1(n20421), .B2(n13632), .A(n13656), .ZN(n13638) );
  OR2_X1 U17079 ( .A1(n20424), .A2(n13633), .ZN(n13634) );
  AND2_X1 U17080 ( .A1(n13634), .A2(n13917), .ZN(n13636) );
  NAND3_X1 U17081 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16172), .A3(
        n20788), .ZN(n14155) );
  AOI22_X1 U17082 ( .A1(n13638), .A2(n13636), .B1(n20559), .B2(n14155), .ZN(
        n13635) );
  NAND2_X1 U17083 ( .A1(n20557), .A2(n13635), .ZN(n13655) );
  INV_X1 U17084 ( .A(n13636), .ZN(n13637) );
  OAI22_X1 U17085 ( .A1(n13638), .A2(n13637), .B1(n20616), .B2(n14155), .ZN(
        n13654) );
  AOI22_X1 U17086 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n13655), .B1(
        n20579), .B2(n13654), .ZN(n13641) );
  AOI22_X1 U17087 ( .A1(n14148), .A2(n20469), .B1(n20580), .B2(n13656), .ZN(
        n13640) );
  OAI211_X1 U17088 ( .C1(n20472), .C2(n20456), .A(n13641), .B(n13640), .ZN(
        P1_U3060) );
  AOI22_X1 U17089 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n13655), .B1(
        n20597), .B2(n13654), .ZN(n13643) );
  AOI22_X1 U17090 ( .A1(n20598), .A2(n13656), .B1(n14148), .B2(n20481), .ZN(
        n13642) );
  OAI211_X1 U17091 ( .C1(n20484), .C2(n20456), .A(n13643), .B(n13642), .ZN(
        P1_U3063) );
  AOI22_X1 U17092 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n13655), .B1(
        n20573), .B2(n13654), .ZN(n13645) );
  AOI22_X1 U17093 ( .A1(n14148), .A2(n20465), .B1(n20574), .B2(n13656), .ZN(
        n13644) );
  OAI211_X1 U17094 ( .C1(n20468), .C2(n20456), .A(n13645), .B(n13644), .ZN(
        P1_U3059) );
  AOI22_X1 U17095 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n13655), .B1(
        n20604), .B2(n13654), .ZN(n13647) );
  AOI22_X1 U17096 ( .A1(n14148), .A2(n20487), .B1(n20606), .B2(n13656), .ZN(
        n13646) );
  OAI211_X1 U17097 ( .C1(n20492), .C2(n20456), .A(n13647), .B(n13646), .ZN(
        P1_U3064) );
  AOI22_X1 U17098 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n13655), .B1(
        n20591), .B2(n13654), .ZN(n13649) );
  AOI22_X1 U17099 ( .A1(n14148), .A2(n20477), .B1(n20592), .B2(n13656), .ZN(
        n13648) );
  OAI211_X1 U17100 ( .C1(n20480), .C2(n20456), .A(n13649), .B(n13648), .ZN(
        P1_U3062) );
  AOI22_X1 U17101 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n13655), .B1(
        n20553), .B2(n13654), .ZN(n13651) );
  AOI22_X1 U17102 ( .A1(n14148), .A2(n20457), .B1(n20554), .B2(n13656), .ZN(
        n13650) );
  OAI211_X1 U17103 ( .C1(n20460), .C2(n20456), .A(n13651), .B(n13650), .ZN(
        P1_U3057) );
  AOI22_X1 U17104 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n13655), .B1(
        n20567), .B2(n13654), .ZN(n13653) );
  AOI22_X1 U17105 ( .A1(n14148), .A2(n20461), .B1(n9857), .B2(n13656), .ZN(
        n13652) );
  OAI211_X1 U17106 ( .C1(n20464), .C2(n20456), .A(n13653), .B(n13652), .ZN(
        P1_U3058) );
  AOI22_X1 U17107 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n13655), .B1(
        n20585), .B2(n13654), .ZN(n13658) );
  AOI22_X1 U17108 ( .A1(n14148), .A2(n20473), .B1(n20586), .B2(n13656), .ZN(
        n13657) );
  OAI211_X1 U17109 ( .C1(n20476), .C2(n20456), .A(n13658), .B(n13657), .ZN(
        P1_U3061) );
  NOR3_X1 U17110 ( .A1(n16172), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20527) );
  INV_X1 U17111 ( .A(n20527), .ZN(n20522) );
  NOR2_X1 U17112 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20522), .ZN(
        n13694) );
  INV_X1 U17113 ( .A(n14158), .ZN(n13664) );
  AOI21_X1 U17114 ( .B1(n20548), .B2(n13668), .A(n20818), .ZN(n13662) );
  INV_X1 U17115 ( .A(n12613), .ZN(n15333) );
  OR2_X1 U17116 ( .A1(n20520), .A2(n15333), .ZN(n13661) );
  INV_X1 U17117 ( .A(n13694), .ZN(n13779) );
  NAND2_X1 U17118 ( .A1(n13661), .A2(n13779), .ZN(n13665) );
  OR2_X1 U17119 ( .A1(n13662), .A2(n13665), .ZN(n13663) );
  OAI211_X1 U17120 ( .C1(n13694), .C2(n16406), .A(n13664), .B(n13663), .ZN(
        n13778) );
  NAND2_X1 U17121 ( .A1(n13665), .A2(n20561), .ZN(n13667) );
  NAND2_X1 U17122 ( .A1(n13826), .A2(n13919), .ZN(n13747) );
  INV_X1 U17123 ( .A(n13747), .ZN(n13743) );
  NAND2_X1 U17124 ( .A1(n14154), .A2(n13743), .ZN(n13666) );
  AND2_X1 U17125 ( .A1(n13667), .A2(n13666), .ZN(n13781) );
  INV_X1 U17126 ( .A(n13781), .ZN(n13693) );
  AOI22_X1 U17127 ( .A1(n20568), .A2(n13694), .B1(n20567), .B2(n13693), .ZN(
        n13670) );
  NAND2_X1 U17128 ( .A1(n13783), .A2(n20461), .ZN(n13669) );
  OAI211_X1 U17129 ( .C1(n20464), .C2(n20548), .A(n13670), .B(n13669), .ZN(
        n13671) );
  AOI21_X1 U17130 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n13671), .ZN(n13672) );
  INV_X1 U17131 ( .A(n13672), .ZN(P1_U3098) );
  AOI22_X1 U17132 ( .A1(n20574), .A2(n13694), .B1(n20573), .B2(n13693), .ZN(
        n13674) );
  NAND2_X1 U17133 ( .A1(n13783), .A2(n20465), .ZN(n13673) );
  OAI211_X1 U17134 ( .C1(n20468), .C2(n20548), .A(n13674), .B(n13673), .ZN(
        n13675) );
  AOI21_X1 U17135 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n13675), .ZN(n13676) );
  INV_X1 U17136 ( .A(n13676), .ZN(P1_U3099) );
  AOI22_X1 U17137 ( .A1(n20592), .A2(n13694), .B1(n20591), .B2(n13693), .ZN(
        n13678) );
  NAND2_X1 U17138 ( .A1(n13783), .A2(n20477), .ZN(n13677) );
  OAI211_X1 U17139 ( .C1(n20480), .C2(n20548), .A(n13678), .B(n13677), .ZN(
        n13679) );
  AOI21_X1 U17140 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n13679), .ZN(n13680) );
  INV_X1 U17141 ( .A(n13680), .ZN(P1_U3102) );
  AOI22_X1 U17142 ( .A1(n20554), .A2(n13694), .B1(n20553), .B2(n13693), .ZN(
        n13682) );
  NAND2_X1 U17143 ( .A1(n13783), .A2(n20457), .ZN(n13681) );
  OAI211_X1 U17144 ( .C1(n20460), .C2(n20548), .A(n13682), .B(n13681), .ZN(
        n13683) );
  AOI21_X1 U17145 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n13683), .ZN(n13684) );
  INV_X1 U17146 ( .A(n13684), .ZN(P1_U3097) );
  AOI22_X1 U17147 ( .A1(n20606), .A2(n13694), .B1(n20604), .B2(n13693), .ZN(
        n13686) );
  NAND2_X1 U17148 ( .A1(n13783), .A2(n20487), .ZN(n13685) );
  OAI211_X1 U17149 ( .C1(n20492), .C2(n20548), .A(n13686), .B(n13685), .ZN(
        n13687) );
  AOI21_X1 U17150 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n13687), .ZN(n13688) );
  INV_X1 U17151 ( .A(n13688), .ZN(P1_U3104) );
  AOI22_X1 U17152 ( .A1(n20586), .A2(n13694), .B1(n20585), .B2(n13693), .ZN(
        n13690) );
  NAND2_X1 U17153 ( .A1(n13783), .A2(n20473), .ZN(n13689) );
  OAI211_X1 U17154 ( .C1(n20476), .C2(n20548), .A(n13690), .B(n13689), .ZN(
        n13691) );
  AOI21_X1 U17155 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n13691), .ZN(n13692) );
  INV_X1 U17156 ( .A(n13692), .ZN(P1_U3101) );
  AOI22_X1 U17157 ( .A1(n20580), .A2(n13694), .B1(n20579), .B2(n13693), .ZN(
        n13696) );
  NAND2_X1 U17158 ( .A1(n13783), .A2(n20469), .ZN(n13695) );
  OAI211_X1 U17159 ( .C1(n20472), .C2(n20548), .A(n13696), .B(n13695), .ZN(
        n13697) );
  AOI21_X1 U17160 ( .B1(n13778), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n13697), .ZN(n13698) );
  INV_X1 U17161 ( .A(n13698), .ZN(P1_U3100) );
  AOI22_X1 U17162 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13702) );
  AOI22_X1 U17163 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13701) );
  AOI22_X1 U17164 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13700) );
  AOI22_X1 U17165 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13699) );
  NAND4_X1 U17166 ( .A1(n13702), .A2(n13701), .A3(n13700), .A4(n13699), .ZN(
        n13708) );
  AOI22_X1 U17167 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13706) );
  AOI22_X1 U17168 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13705) );
  AOI22_X1 U17169 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13704) );
  AOI22_X1 U17170 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14508), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13703) );
  NAND4_X1 U17171 ( .A1(n13706), .A2(n13705), .A3(n13704), .A4(n13703), .ZN(
        n13707) );
  NOR2_X1 U17172 ( .A1(n13708), .A2(n13707), .ZN(n13710) );
  OR2_X1 U17173 ( .A1(n13817), .A2(n13816), .ZN(n13709) );
  OR2_X1 U17174 ( .A1(n13710), .A2(n13816), .ZN(n13858) );
  NOR2_X1 U17175 ( .A1(n13817), .A2(n13858), .ZN(n13862) );
  AOI21_X1 U17176 ( .B1(n13710), .B2(n13709), .A(n13862), .ZN(n13711) );
  INV_X1 U17177 ( .A(n13711), .ZN(n13882) );
  AOI21_X1 U17178 ( .B1(n15938), .B2(n15954), .A(n13712), .ZN(n13713) );
  OR2_X1 U17179 ( .A1(n13865), .A2(n13713), .ZN(n19224) );
  INV_X1 U17180 ( .A(n19224), .ZN(n13721) );
  OAI22_X1 U17181 ( .A1(n15577), .A2(n19508), .B1(n13714), .B2(n19387), .ZN(
        n13720) );
  INV_X1 U17182 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n13718) );
  INV_X1 U17183 ( .A(n19356), .ZN(n15579) );
  OAI22_X1 U17184 ( .A1(n15581), .A2(n13718), .B1(n15579), .B2(n16749), .ZN(
        n13719) );
  AOI211_X1 U17185 ( .C1(n19416), .C2(n13721), .A(n13720), .B(n13719), .ZN(
        n13722) );
  OAI21_X1 U17186 ( .B1(n13882), .B2(n19390), .A(n13722), .ZN(P2_U2903) );
  XOR2_X1 U17187 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13724), .Z(
        n13725) );
  XNOR2_X1 U17188 ( .A(n13723), .B(n13725), .ZN(n13739) );
  INV_X1 U17189 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13726) );
  NOR2_X1 U17190 ( .A1(n20254), .A2(n13726), .ZN(n13736) );
  AOI21_X1 U17191 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13736), .ZN(n13727) );
  OAI21_X1 U17192 ( .B1(n20361), .B2(n20248), .A(n13727), .ZN(n13728) );
  AOI21_X1 U17193 ( .B1(n13729), .B2(n14067), .A(n13728), .ZN(n13730) );
  OAI21_X1 U17194 ( .B1(n13739), .B2(n20203), .A(n13730), .ZN(P1_U2993) );
  NOR2_X1 U17195 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15293), .ZN(
        n15324) );
  NAND3_X1 U17196 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n20382), .ZN(n13734) );
  NOR2_X1 U17197 ( .A1(n20963), .A2(n20380), .ZN(n20364) );
  NAND2_X1 U17198 ( .A1(n20364), .A2(n16388), .ZN(n16393) );
  INV_X1 U17199 ( .A(n20364), .ZN(n13733) );
  NOR2_X1 U17200 ( .A1(n20962), .A2(n13731), .ZN(n20388) );
  NOR2_X1 U17201 ( .A1(n15304), .A2(n20388), .ZN(n20384) );
  NOR2_X1 U17202 ( .A1(n16388), .A2(n13733), .ZN(n14055) );
  OAI21_X1 U17203 ( .B1(n13732), .B2(n13731), .A(n20962), .ZN(n20362) );
  NAND2_X1 U17204 ( .A1(n14055), .A2(n20362), .ZN(n14388) );
  AOI21_X1 U17205 ( .B1(n20389), .B2(n14388), .A(n20383), .ZN(n15302) );
  INV_X1 U17206 ( .A(n15302), .ZN(n14056) );
  AOI211_X1 U17207 ( .C1(n14387), .C2(n13733), .A(n20384), .B(n14056), .ZN(
        n16389) );
  OAI21_X1 U17208 ( .B1(n13734), .B2(n16393), .A(n16389), .ZN(n16367) );
  NAND2_X1 U17209 ( .A1(n20363), .A2(n13734), .ZN(n16344) );
  NAND2_X1 U17210 ( .A1(n20362), .A2(n16344), .ZN(n20375) );
  INV_X1 U17211 ( .A(n20375), .ZN(n13735) );
  INV_X1 U17212 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16369) );
  AOI22_X1 U17213 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16367), .B1(
        n16370), .B2(n16369), .ZN(n13738) );
  AOI21_X1 U17214 ( .B1(n20246), .B2(n20374), .A(n13736), .ZN(n13737) );
  OAI211_X1 U17215 ( .C1(n13739), .C2(n20385), .A(n13738), .B(n13737), .ZN(
        P1_U3025) );
  AOI21_X1 U17216 ( .B1(n13741), .B2(n20612), .A(n20818), .ZN(n13742) );
  NOR2_X1 U17217 ( .A1(n13742), .A2(n20559), .ZN(n13745) );
  NOR2_X1 U17218 ( .A1(n14105), .A2(n15333), .ZN(n13749) );
  INV_X1 U17219 ( .A(n20451), .ZN(n14103) );
  AOI22_X1 U17220 ( .A1(n13745), .A2(n13749), .B1(n13743), .B2(n14103), .ZN(
        n13777) );
  NOR3_X1 U17221 ( .A1(n20788), .A2(n16172), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20560) );
  NAND2_X1 U17222 ( .A1(n20549), .A2(n20560), .ZN(n13771) );
  OAI22_X1 U17223 ( .A1(n14128), .A2(n13771), .B1(n20492), .B2(n20612), .ZN(
        n13744) );
  AOI21_X1 U17224 ( .B1(n13773), .B2(n20487), .A(n13744), .ZN(n13752) );
  INV_X1 U17225 ( .A(n13745), .ZN(n13750) );
  AOI22_X1 U17226 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n13747), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n13771), .ZN(n13748) );
  NAND2_X1 U17227 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n13751) );
  OAI211_X1 U17228 ( .C1(n13777), .C2(n14181), .A(n13752), .B(n13751), .ZN(
        P1_U3136) );
  OAI22_X1 U17229 ( .A1(n14137), .A2(n13771), .B1(n20460), .B2(n20612), .ZN(
        n13753) );
  AOI21_X1 U17230 ( .B1(n13773), .B2(n20457), .A(n13753), .ZN(n13755) );
  NAND2_X1 U17231 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n13754) );
  OAI211_X1 U17232 ( .C1(n13777), .C2(n14169), .A(n13755), .B(n13754), .ZN(
        P1_U3129) );
  OAI22_X1 U17233 ( .A1(n14120), .A2(n13771), .B1(n20480), .B2(n20612), .ZN(
        n13756) );
  AOI21_X1 U17234 ( .B1(n13773), .B2(n20477), .A(n13756), .ZN(n13758) );
  NAND2_X1 U17235 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n13757) );
  OAI211_X1 U17236 ( .C1(n13777), .C2(n14189), .A(n13758), .B(n13757), .ZN(
        P1_U3134) );
  OAI22_X1 U17237 ( .A1(n14144), .A2(n13771), .B1(n20476), .B2(n20612), .ZN(
        n13759) );
  AOI21_X1 U17238 ( .B1(n13773), .B2(n20473), .A(n13759), .ZN(n13761) );
  NAND2_X1 U17239 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13760) );
  OAI211_X1 U17240 ( .C1(n13777), .C2(n14196), .A(n13761), .B(n13760), .ZN(
        P1_U3133) );
  OAI22_X1 U17241 ( .A1(n14112), .A2(n13771), .B1(n20472), .B2(n20612), .ZN(
        n13762) );
  AOI21_X1 U17242 ( .B1(n13773), .B2(n20469), .A(n13762), .ZN(n13764) );
  NAND2_X1 U17243 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n13763) );
  OAI211_X1 U17244 ( .C1(n13777), .C2(n14177), .A(n13764), .B(n13763), .ZN(
        P1_U3132) );
  OAI22_X1 U17245 ( .A1(n14124), .A2(n13771), .B1(n20468), .B2(n20612), .ZN(
        n13765) );
  AOI21_X1 U17246 ( .B1(n13773), .B2(n20465), .A(n13765), .ZN(n13767) );
  NAND2_X1 U17247 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13766) );
  OAI211_X1 U17248 ( .C1(n13777), .C2(n14185), .A(n13767), .B(n13766), .ZN(
        P1_U3131) );
  OAI22_X1 U17249 ( .A1(n13780), .A2(n13771), .B1(n20484), .B2(n20612), .ZN(
        n13768) );
  AOI21_X1 U17250 ( .B1(n13773), .B2(n20481), .A(n13768), .ZN(n13770) );
  NAND2_X1 U17251 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n13769) );
  OAI211_X1 U17252 ( .C1(n13777), .C2(n14165), .A(n13770), .B(n13769), .ZN(
        P1_U3135) );
  OAI22_X1 U17253 ( .A1(n14116), .A2(n13771), .B1(n20464), .B2(n20612), .ZN(
        n13772) );
  AOI21_X1 U17254 ( .B1(n13773), .B2(n20461), .A(n13772), .ZN(n13776) );
  NAND2_X1 U17255 ( .A1(n13774), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n13775) );
  OAI211_X1 U17256 ( .C1(n13777), .C2(n14173), .A(n13776), .B(n13775), .ZN(
        P1_U3130) );
  NAND2_X1 U17257 ( .A1(n13778), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n13785) );
  OAI22_X1 U17258 ( .A1(n14165), .A2(n13781), .B1(n13780), .B2(n13779), .ZN(
        n13782) );
  AOI21_X1 U17259 ( .B1(n13783), .B2(n20481), .A(n13782), .ZN(n13784) );
  OAI211_X1 U17260 ( .C1(n20484), .C2(n20548), .A(n13785), .B(n13784), .ZN(
        P1_U3103) );
  AOI21_X1 U17261 ( .B1(n13788), .B2(n13612), .A(n13787), .ZN(n14011) );
  INV_X1 U17262 ( .A(n14011), .ZN(n13876) );
  INV_X1 U17263 ( .A(n14293), .ZN(n14232) );
  AOI22_X1 U17264 ( .A1(n14232), .A2(n14960), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n16280), .ZN(n13789) );
  OAI21_X1 U17265 ( .B1(n13876), .B2(n16283), .A(n13789), .ZN(P1_U2896) );
  XNOR2_X1 U17266 ( .A(n13790), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13792) );
  XNOR2_X1 U17267 ( .A(n13792), .B(n13791), .ZN(n19463) );
  XOR2_X1 U17268 ( .A(n13794), .B(n13793), .Z(n19462) );
  INV_X1 U17269 ( .A(n16578), .ZN(n13995) );
  INV_X1 U17270 ( .A(n13795), .ZN(n16643) );
  NOR2_X1 U17271 ( .A1(n13995), .A2(n16643), .ZN(n16620) );
  NOR2_X1 U17272 ( .A1(n10868), .A2(n19304), .ZN(n13796) );
  AOI221_X1 U17273 ( .B1(n16620), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n16627), .C2(n13797), .A(n13796), .ZN(n13799) );
  NAND2_X1 U17274 ( .A1(n19467), .A2(n16635), .ZN(n13798) );
  OAI211_X1 U17275 ( .C1(n19322), .C2(n19487), .A(n13799), .B(n13798), .ZN(
        n13800) );
  AOI21_X1 U17276 ( .B1(n19462), .B2(n16639), .A(n13800), .ZN(n13801) );
  OAI21_X1 U17277 ( .B1(n19490), .B2(n19463), .A(n13801), .ZN(P2_U3042) );
  INV_X1 U17278 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n16371) );
  NAND4_X1 U17279 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20249)
         );
  NAND2_X1 U17280 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n13802) );
  NOR3_X1 U17281 ( .A1(n20271), .A2(n20249), .A3(n13802), .ZN(n20232) );
  NAND2_X1 U17282 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20232), .ZN(n14262) );
  NAND2_X1 U17283 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .ZN(n13804) );
  INV_X1 U17284 ( .A(n13802), .ZN(n13803) );
  NOR2_X1 U17285 ( .A1(n14892), .A2(n20249), .ZN(n20251) );
  AOI21_X1 U17286 ( .B1(n13803), .B2(n20251), .A(n20252), .ZN(n20239) );
  AOI21_X1 U17287 ( .B1(n13804), .B2(n14847), .A(n20239), .ZN(n20227) );
  AOI21_X1 U17288 ( .B1(n16371), .B2(n14262), .A(n20227), .ZN(n13805) );
  INV_X1 U17289 ( .A(n13805), .ZN(n13815) );
  INV_X1 U17290 ( .A(n14009), .ZN(n13813) );
  MUX2_X1 U17291 ( .A(n13168), .B(n14335), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13807) );
  NAND2_X1 U17292 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n14341), .ZN(
        n13806) );
  AND2_X1 U17293 ( .A1(n13809), .A2(n13808), .ZN(n13810) );
  OR2_X1 U17294 ( .A1(n13810), .A2(n9821), .ZN(n16372) );
  AOI22_X1 U17295 ( .A1(P1_EBX_REG_8__SCAN_IN), .A2(n20263), .B1(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n20269), .ZN(n13811) );
  OAI211_X1 U17296 ( .C1(n20267), .C2(n16372), .A(n13811), .B(n20254), .ZN(
        n13812) );
  AOI21_X1 U17297 ( .B1(n20221), .B2(n13813), .A(n13812), .ZN(n13814) );
  OAI211_X1 U17298 ( .C1(n13876), .C2(n20242), .A(n13815), .B(n13814), .ZN(
        P1_U2832) );
  XNOR2_X1 U17299 ( .A(n13817), .B(n13816), .ZN(n13824) );
  OR2_X1 U17300 ( .A1(n13820), .A2(n13819), .ZN(n13821) );
  NAND2_X1 U17301 ( .A1(n13818), .A2(n13821), .ZN(n19232) );
  INV_X1 U17302 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13822) );
  MUX2_X1 U17303 ( .A(n19232), .B(n13822), .S(n9726), .Z(n13823) );
  OAI21_X1 U17304 ( .B1(n13824), .B2(n15539), .A(n13823), .ZN(P2_U2872) );
  INV_X1 U17305 ( .A(n20447), .ZN(n13839) );
  OAI21_X1 U17306 ( .B1(n13839), .B2(n20414), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13825) );
  NAND2_X1 U17307 ( .A1(n13825), .A2(n20561), .ZN(n13831) );
  NAND2_X1 U17308 ( .A1(n20421), .A2(n12613), .ZN(n13834) );
  INV_X1 U17309 ( .A(n14154), .ZN(n13828) );
  INV_X1 U17310 ( .A(n13826), .ZN(n13827) );
  NAND2_X1 U17311 ( .A1(n13827), .A2(n13919), .ZN(n20450) );
  INV_X1 U17312 ( .A(n20416), .ZN(n13841) );
  NOR3_X1 U17313 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20426) );
  INV_X1 U17314 ( .A(n20426), .ZN(n20422) );
  NOR2_X1 U17315 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20422), .ZN(
        n20415) );
  NAND2_X1 U17316 ( .A1(n20554), .A2(n20415), .ZN(n13829) );
  OAI21_X1 U17317 ( .B1(n20566), .B2(n13830), .A(n13829), .ZN(n13838) );
  INV_X1 U17318 ( .A(n13831), .ZN(n13835) );
  INV_X1 U17319 ( .A(n20450), .ZN(n13832) );
  OAI22_X1 U17320 ( .A1(n13832), .A2(n20616), .B1(n20415), .B2(n16406), .ZN(
        n13833) );
  AOI211_X1 U17321 ( .C1(n13835), .C2(n13834), .A(n14158), .B(n13833), .ZN(
        n20401) );
  NOR2_X1 U17322 ( .A1(n20401), .A2(n13836), .ZN(n13837) );
  AOI211_X1 U17323 ( .C1(n13839), .C2(n20563), .A(n13838), .B(n13837), .ZN(
        n13840) );
  OAI21_X1 U17324 ( .B1(n13841), .B2(n14169), .A(n13840), .ZN(P1_U3033) );
  AOI22_X1 U17325 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13845) );
  AOI22_X1 U17326 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17327 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U17328 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13842) );
  NAND4_X1 U17329 ( .A1(n13845), .A2(n13844), .A3(n13843), .A4(n13842), .ZN(
        n13857) );
  AOI22_X1 U17330 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13855) );
  AOI22_X1 U17331 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13854) );
  AOI22_X1 U17332 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n13846), .ZN(n13853) );
  INV_X1 U17333 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14531) );
  INV_X1 U17334 ( .A(n13847), .ZN(n13850) );
  INV_X1 U17335 ( .A(n13848), .ZN(n13849) );
  INV_X1 U17336 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20925) );
  OAI22_X1 U17337 ( .A1(n14531), .A2(n13850), .B1(n13849), .B2(n20925), .ZN(
        n13851) );
  INV_X1 U17338 ( .A(n13851), .ZN(n13852) );
  NAND4_X1 U17339 ( .A1(n13855), .A2(n13854), .A3(n13853), .A4(n13852), .ZN(
        n13856) );
  OR2_X1 U17340 ( .A1(n13857), .A2(n13856), .ZN(n13861) );
  INV_X1 U17341 ( .A(n13861), .ZN(n13859) );
  NOR2_X1 U17342 ( .A1(n13859), .A2(n13858), .ZN(n13905) );
  AND2_X1 U17343 ( .A1(n13907), .A2(n13905), .ZN(n13909) );
  INV_X1 U17344 ( .A(n13909), .ZN(n13860) );
  OAI21_X1 U17345 ( .B1(n13862), .B2(n13861), .A(n13860), .ZN(n14076) );
  OAI21_X1 U17346 ( .B1(n13865), .B2(n13864), .A(n13863), .ZN(n15914) );
  INV_X1 U17347 ( .A(n15914), .ZN(n14204) );
  OAI22_X1 U17348 ( .A1(n15577), .A2(n19515), .B1(n13866), .B2(n19387), .ZN(
        n13870) );
  INV_X1 U17349 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13868) );
  INV_X1 U17350 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n13867) );
  OAI22_X1 U17351 ( .A1(n15581), .A2(n13868), .B1(n15579), .B2(n13867), .ZN(
        n13869) );
  AOI211_X1 U17352 ( .C1(n19416), .C2(n14204), .A(n13870), .B(n13869), .ZN(
        n13871) );
  OAI21_X1 U17353 ( .B1(n14076), .B2(n19390), .A(n13871), .ZN(P2_U2902) );
  NOR2_X1 U17354 ( .A1(n13787), .A2(n13873), .ZN(n13874) );
  OR2_X1 U17355 ( .A1(n13872), .A2(n13874), .ZN(n14066) );
  MUX2_X1 U17356 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n14279), .Z(
        n20324) );
  AOI22_X1 U17357 ( .A1(n14232), .A2(n20324), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n16280), .ZN(n13875) );
  OAI21_X1 U17358 ( .B1(n14066), .B2(n16283), .A(n13875), .ZN(P1_U2895) );
  INV_X1 U17359 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13877) );
  OAI222_X1 U17360 ( .A1(n16372), .A2(n14936), .B1(n20282), .B2(n13877), .C1(
        n14939), .C2(n13876), .ZN(P1_U2864) );
  NAND2_X1 U17361 ( .A1(n13818), .A2(n13878), .ZN(n13879) );
  AND2_X1 U17362 ( .A1(n14072), .A2(n13879), .ZN(n19220) );
  NOR2_X1 U17363 ( .A1(n15537), .A2(n10660), .ZN(n13880) );
  AOI21_X1 U17364 ( .B1(n19220), .B2(n15537), .A(n13880), .ZN(n13881) );
  OAI21_X1 U17365 ( .B1(n13882), .B2(n15539), .A(n13881), .ZN(P2_U2871) );
  NOR2_X2 U17366 ( .A1(n19403), .A2(n19913), .ZN(n20018) );
  OAI21_X1 U17367 ( .B1(n19984), .B2(n20046), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13883) );
  NAND2_X1 U17368 ( .A1(n13883), .A2(n20152), .ZN(n13885) );
  NOR3_X2 U17369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20142), .A3(
        n19989), .ZN(n19982) );
  NOR2_X1 U17370 ( .A1(n19982), .A2(n19961), .ZN(n13888) );
  OAI21_X1 U17371 ( .B1(n13886), .B2(n19982), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13884) );
  OAI21_X1 U17372 ( .B1(n13885), .B2(n13888), .A(n13884), .ZN(n19985) );
  INV_X1 U17373 ( .A(n13885), .ZN(n13889) );
  AOI211_X1 U17374 ( .C1(n13886), .C2(n19670), .A(n19982), .B(n20152), .ZN(
        n13887) );
  AOI211_X2 U17375 ( .C1(n13889), .C2(n13888), .A(n13887), .B(n19913), .ZN(
        n19988) );
  INV_X1 U17376 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14587) );
  AOI22_X1 U17377 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19531), .ZN(n20022) );
  AND2_X1 U17378 ( .A1(n13890), .A2(n19525), .ZN(n20017) );
  AOI22_X1 U17379 ( .A1(n19955), .A2(n20046), .B1(n19982), .B2(n20017), .ZN(
        n13892) );
  AOI22_X1 U17380 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19531), .ZN(n19929) );
  INV_X1 U17381 ( .A(n19929), .ZN(n20019) );
  NAND2_X1 U17382 ( .A1(n20019), .A2(n19984), .ZN(n13891) );
  OAI211_X1 U17383 ( .C1(n19988), .C2(n14587), .A(n13892), .B(n13891), .ZN(
        n13893) );
  AOI21_X1 U17384 ( .B1(n20018), .B2(n19985), .A(n13893), .ZN(n13894) );
  INV_X1 U17385 ( .A(n13894), .ZN(P2_U3163) );
  AOI22_X1 U17386 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U17387 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13897) );
  AOI22_X1 U17388 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U17389 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13895) );
  NAND4_X1 U17390 ( .A1(n13898), .A2(n13897), .A3(n13896), .A4(n13895), .ZN(
        n13904) );
  AOI22_X1 U17391 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13902) );
  AOI22_X1 U17392 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U17393 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17394 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__2__SCAN_IN), .B2(n14508), .ZN(n13899) );
  NAND4_X1 U17395 ( .A1(n13902), .A2(n13901), .A3(n13900), .A4(n13899), .ZN(
        n13903) );
  OR2_X1 U17396 ( .A1(n13904), .A2(n13903), .ZN(n13908) );
  AND2_X1 U17397 ( .A1(n13908), .A2(n13905), .ZN(n13906) );
  OAI21_X1 U17398 ( .B1(n13909), .B2(n13908), .A(n13979), .ZN(n14202) );
  NAND2_X1 U17399 ( .A1(n13863), .A2(n13910), .ZN(n13911) );
  NAND2_X1 U17400 ( .A1(n13982), .A2(n13911), .ZN(n19213) );
  INV_X1 U17401 ( .A(n19213), .ZN(n15903) );
  OAI22_X1 U17402 ( .A1(n15577), .A2(n19518), .B1(n13912), .B2(n19387), .ZN(
        n13915) );
  INV_X1 U17403 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n13913) );
  OAI22_X1 U17404 ( .A1(n15581), .A2(n13913), .B1(n15579), .B2(n16746), .ZN(
        n13914) );
  AOI211_X1 U17405 ( .C1(n19416), .C2(n15903), .A(n13915), .B(n13914), .ZN(
        n13916) );
  OAI21_X1 U17406 ( .B1(n14202), .B2(n19390), .A(n13916), .ZN(P2_U2901) );
  NAND3_X1 U17407 ( .A1(n13920), .A2(n13951), .A3(n13917), .ZN(n13918) );
  NAND2_X1 U17408 ( .A1(n13918), .A2(n14150), .ZN(n13925) );
  OR2_X1 U17409 ( .A1(n13919), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13923) );
  INV_X1 U17410 ( .A(n13923), .ZN(n14153) );
  NOR2_X1 U17411 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13921), .ZN(
        n13949) );
  INV_X1 U17412 ( .A(n13922), .ZN(n13924) );
  AND2_X1 U17413 ( .A1(n13923), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14157) );
  AOI21_X1 U17414 ( .B1(n13925), .B2(n13924), .A(n14157), .ZN(n13926) );
  OAI211_X1 U17415 ( .C1(n13949), .C2(n16406), .A(n20454), .B(n13926), .ZN(
        n13948) );
  AOI22_X1 U17416 ( .A1(n20554), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n13948), .ZN(n13927) );
  OAI21_X1 U17417 ( .B1(n20460), .B2(n13951), .A(n13927), .ZN(n13928) );
  AOI21_X1 U17418 ( .B1(n20515), .B2(n20457), .A(n13928), .ZN(n13929) );
  OAI21_X1 U17419 ( .B1(n13954), .B2(n14169), .A(n13929), .ZN(P1_U3081) );
  AOI22_X1 U17420 ( .A1(n20586), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n13948), .ZN(n13930) );
  OAI21_X1 U17421 ( .B1(n20476), .B2(n13951), .A(n13930), .ZN(n13931) );
  AOI21_X1 U17422 ( .B1(n20515), .B2(n20473), .A(n13931), .ZN(n13932) );
  OAI21_X1 U17423 ( .B1(n13954), .B2(n14196), .A(n13932), .ZN(P1_U3085) );
  AOI22_X1 U17424 ( .A1(n20598), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n13948), .ZN(n13933) );
  OAI21_X1 U17425 ( .B1(n20484), .B2(n13951), .A(n13933), .ZN(n13934) );
  AOI21_X1 U17426 ( .B1(n20515), .B2(n20481), .A(n13934), .ZN(n13935) );
  OAI21_X1 U17427 ( .B1(n13954), .B2(n14165), .A(n13935), .ZN(P1_U3087) );
  AOI22_X1 U17428 ( .A1(n20592), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n13948), .ZN(n13936) );
  OAI21_X1 U17429 ( .B1(n20480), .B2(n13951), .A(n13936), .ZN(n13937) );
  AOI21_X1 U17430 ( .B1(n20515), .B2(n20477), .A(n13937), .ZN(n13938) );
  OAI21_X1 U17431 ( .B1(n13954), .B2(n14189), .A(n13938), .ZN(P1_U3086) );
  AOI22_X1 U17432 ( .A1(n20574), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n13948), .ZN(n13939) );
  OAI21_X1 U17433 ( .B1(n20468), .B2(n13951), .A(n13939), .ZN(n13940) );
  AOI21_X1 U17434 ( .B1(n20515), .B2(n20465), .A(n13940), .ZN(n13941) );
  OAI21_X1 U17435 ( .B1(n13954), .B2(n14185), .A(n13941), .ZN(P1_U3083) );
  AOI22_X1 U17436 ( .A1(n20580), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n13948), .ZN(n13942) );
  OAI21_X1 U17437 ( .B1(n20472), .B2(n13951), .A(n13942), .ZN(n13943) );
  AOI21_X1 U17438 ( .B1(n20515), .B2(n20469), .A(n13943), .ZN(n13944) );
  OAI21_X1 U17439 ( .B1(n13954), .B2(n14177), .A(n13944), .ZN(P1_U3084) );
  AOI22_X1 U17440 ( .A1(n20606), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n13948), .ZN(n13945) );
  OAI21_X1 U17441 ( .B1(n20492), .B2(n13951), .A(n13945), .ZN(n13946) );
  AOI21_X1 U17442 ( .B1(n20515), .B2(n20487), .A(n13946), .ZN(n13947) );
  OAI21_X1 U17443 ( .B1(n13954), .B2(n14181), .A(n13947), .ZN(P1_U3088) );
  AOI22_X1 U17444 ( .A1(n20568), .A2(n13949), .B1(
        P1_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n13948), .ZN(n13950) );
  OAI21_X1 U17445 ( .B1(n20464), .B2(n13951), .A(n13950), .ZN(n13952) );
  AOI21_X1 U17446 ( .B1(n20515), .B2(n20461), .A(n13952), .ZN(n13953) );
  OAI21_X1 U17447 ( .B1(n13954), .B2(n14173), .A(n13953), .ZN(P1_U3082) );
  OAI21_X1 U17448 ( .B1(n13872), .B2(n13956), .A(n13955), .ZN(n15146) );
  OR2_X1 U17449 ( .A1(n13168), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n13961) );
  INV_X1 U17450 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13957) );
  NAND2_X1 U17451 ( .A1(n14335), .A2(n13957), .ZN(n13959) );
  INV_X1 U17452 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14875) );
  NAND2_X1 U17453 ( .A1(n14308), .A2(n14875), .ZN(n13958) );
  NAND3_X1 U17454 ( .A1(n13959), .A2(n14313), .A3(n13958), .ZN(n13960) );
  INV_X1 U17455 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n20281) );
  NAND2_X1 U17456 ( .A1(n14326), .A2(n20281), .ZN(n13964) );
  NAND2_X1 U17457 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13962) );
  OAI211_X1 U17458 ( .C1(n14341), .C2(P1_EBX_REG_9__SCAN_IN), .A(n14335), .B(
        n13962), .ZN(n13963) );
  INV_X1 U17459 ( .A(n14237), .ZN(n14295) );
  AOI21_X1 U17460 ( .B1(n13966), .B2(n13965), .A(n14237), .ZN(n16360) );
  AOI22_X1 U17461 ( .A1(n16360), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n13967) );
  OAI21_X1 U17462 ( .B1(n15146), .B2(n14939), .A(n13967), .ZN(P1_U2862) );
  MUX2_X1 U17463 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n14279), .Z(
        n20326) );
  AOI22_X1 U17464 ( .A1(n14232), .A2(n20326), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n16280), .ZN(n13968) );
  OAI21_X1 U17465 ( .B1(n15146), .B2(n16283), .A(n13968), .ZN(P1_U2894) );
  INV_X1 U17466 ( .A(n13979), .ZN(n13980) );
  AOI22_X1 U17467 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13972) );
  AOI22_X1 U17468 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13971) );
  AOI22_X1 U17469 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13970) );
  AOI22_X1 U17470 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13969) );
  NAND4_X1 U17471 ( .A1(n13972), .A2(n13971), .A3(n13970), .A4(n13969), .ZN(
        n13978) );
  AOI22_X1 U17472 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13976) );
  AOI22_X1 U17473 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17474 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17475 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__3__SCAN_IN), .B2(n14508), .ZN(n13973) );
  NAND4_X1 U17476 ( .A1(n13976), .A2(n13975), .A3(n13974), .A4(n13973), .ZN(
        n13977) );
  OAI21_X1 U17477 ( .B1(n13980), .B2(n9846), .A(n14087), .ZN(n14225) );
  AND2_X1 U17478 ( .A1(n13982), .A2(n13981), .ZN(n13983) );
  NOR2_X1 U17479 ( .A1(n14092), .A2(n13983), .ZN(n19196) );
  OAI22_X1 U17480 ( .A1(n15577), .A2(n19403), .B1(n13984), .B2(n19387), .ZN(
        n13988) );
  INV_X1 U17481 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n13986) );
  INV_X1 U17482 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n13985) );
  OAI22_X1 U17483 ( .A1(n15581), .A2(n13986), .B1(n15579), .B2(n13985), .ZN(
        n13987) );
  AOI211_X1 U17484 ( .C1(n19416), .C2(n19196), .A(n13988), .B(n13987), .ZN(
        n13989) );
  OAI21_X1 U17485 ( .B1(n14225), .B2(n19390), .A(n13989), .ZN(P2_U2900) );
  XNOR2_X1 U17486 ( .A(n13990), .B(n13991), .ZN(n14020) );
  OAI21_X1 U17487 ( .B1(n13993), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13992), .ZN(n13994) );
  INV_X1 U17488 ( .A(n13994), .ZN(n14018) );
  NAND2_X1 U17489 ( .A1(n14018), .A2(n16624), .ZN(n14004) );
  INV_X1 U17490 ( .A(n15988), .ZN(n16610) );
  AOI21_X1 U17491 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n13996), .A(
        n13995), .ZN(n16615) );
  AOI22_X1 U17492 ( .A1(n19326), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16615), .ZN(n13997) );
  OAI21_X1 U17493 ( .B1(n19491), .B2(n14015), .A(n13997), .ZN(n14002) );
  OAI21_X1 U17494 ( .B1(n13998), .B2(n14000), .A(n13999), .ZN(n19386) );
  NOR2_X1 U17495 ( .A1(n19386), .A2(n19487), .ZN(n14001) );
  AOI211_X1 U17496 ( .C1(n16610), .C2(n15989), .A(n14002), .B(n14001), .ZN(
        n14003) );
  OAI211_X1 U17497 ( .C1(n14020), .C2(n19500), .A(n14004), .B(n14003), .ZN(
        P2_U3040) );
  XNOR2_X1 U17498 ( .A(n14006), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14007) );
  XNOR2_X1 U17499 ( .A(n14005), .B(n14007), .ZN(n16375) );
  INV_X1 U17500 ( .A(n16375), .ZN(n14013) );
  AOI22_X1 U17501 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n14008) );
  OAI21_X1 U17502 ( .B1(n20361), .B2(n14009), .A(n14008), .ZN(n14010) );
  AOI21_X1 U17503 ( .B1(n14011), .B2(n14067), .A(n14010), .ZN(n14012) );
  OAI21_X1 U17504 ( .B1(n14013), .B2(n20203), .A(n14012), .ZN(P1_U2991) );
  OAI22_X1 U17505 ( .A1(n10012), .A2(n16541), .B1(n19471), .B2(n19312), .ZN(
        n14017) );
  OAI22_X1 U17506 ( .A1(n13256), .A2(n14015), .B1(n19304), .B2(n14014), .ZN(
        n14016) );
  AOI211_X1 U17507 ( .C1(n14018), .C2(n19475), .A(n14017), .B(n14016), .ZN(
        n14019) );
  OAI21_X1 U17508 ( .B1(n16514), .B2(n14020), .A(n14019), .ZN(P2_U3008) );
  AOI22_X1 U17509 ( .A1(n9857), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n14045), .ZN(n14022) );
  NAND2_X1 U17510 ( .A1(n20544), .A2(n20461), .ZN(n14021) );
  OAI211_X1 U17511 ( .C1(n20464), .C2(n14048), .A(n14022), .B(n14021), .ZN(
        n14023) );
  INV_X1 U17512 ( .A(n14023), .ZN(n14024) );
  OAI21_X1 U17513 ( .B1(n14051), .B2(n14173), .A(n14024), .ZN(P1_U3114) );
  AOI22_X1 U17514 ( .A1(n20574), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__2__SCAN_IN), .B2(n14045), .ZN(n14026) );
  NAND2_X1 U17515 ( .A1(n20544), .A2(n20465), .ZN(n14025) );
  OAI211_X1 U17516 ( .C1(n20468), .C2(n14048), .A(n14026), .B(n14025), .ZN(
        n14027) );
  INV_X1 U17517 ( .A(n14027), .ZN(n14028) );
  OAI21_X1 U17518 ( .B1(n14051), .B2(n14185), .A(n14028), .ZN(P1_U3115) );
  AOI22_X1 U17519 ( .A1(n20606), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n14045), .ZN(n14030) );
  NAND2_X1 U17520 ( .A1(n20544), .A2(n20487), .ZN(n14029) );
  OAI211_X1 U17521 ( .C1(n20492), .C2(n14048), .A(n14030), .B(n14029), .ZN(
        n14031) );
  INV_X1 U17522 ( .A(n14031), .ZN(n14032) );
  OAI21_X1 U17523 ( .B1(n14051), .B2(n14181), .A(n14032), .ZN(P1_U3120) );
  AOI22_X1 U17524 ( .A1(n20580), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n14045), .ZN(n14034) );
  NAND2_X1 U17525 ( .A1(n20544), .A2(n20469), .ZN(n14033) );
  OAI211_X1 U17526 ( .C1(n20472), .C2(n14048), .A(n14034), .B(n14033), .ZN(
        n14035) );
  INV_X1 U17527 ( .A(n14035), .ZN(n14036) );
  OAI21_X1 U17528 ( .B1(n14051), .B2(n14177), .A(n14036), .ZN(P1_U3116) );
  AOI22_X1 U17529 ( .A1(n20592), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__5__SCAN_IN), .B2(n14045), .ZN(n14038) );
  NAND2_X1 U17530 ( .A1(n20544), .A2(n20477), .ZN(n14037) );
  OAI211_X1 U17531 ( .C1(n20480), .C2(n14048), .A(n14038), .B(n14037), .ZN(
        n14039) );
  INV_X1 U17532 ( .A(n14039), .ZN(n14040) );
  OAI21_X1 U17533 ( .B1(n14051), .B2(n14189), .A(n14040), .ZN(P1_U3118) );
  AOI22_X1 U17534 ( .A1(n20586), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n14045), .ZN(n14042) );
  NAND2_X1 U17535 ( .A1(n20544), .A2(n20473), .ZN(n14041) );
  OAI211_X1 U17536 ( .C1(n20476), .C2(n14048), .A(n14042), .B(n14041), .ZN(
        n14043) );
  INV_X1 U17537 ( .A(n14043), .ZN(n14044) );
  OAI21_X1 U17538 ( .B1(n14051), .B2(n14196), .A(n14044), .ZN(P1_U3117) );
  AOI22_X1 U17539 ( .A1(n20554), .A2(n14046), .B1(
        P1_INSTQUEUE_REG_10__0__SCAN_IN), .B2(n14045), .ZN(n14047) );
  OAI21_X1 U17540 ( .B1(n20460), .B2(n14048), .A(n14047), .ZN(n14049) );
  AOI21_X1 U17541 ( .B1(n20544), .B2(n20457), .A(n14049), .ZN(n14050) );
  OAI21_X1 U17542 ( .B1(n14051), .B2(n14169), .A(n14050), .ZN(P1_U3113) );
  MUX2_X1 U17543 ( .A(n14053), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .S(
        n11601), .Z(n14054) );
  XNOR2_X1 U17544 ( .A(n14052), .B(n14054), .ZN(n14070) );
  INV_X1 U17545 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16377) );
  INV_X1 U17546 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20964) );
  NOR3_X1 U17547 ( .A1(n16377), .A2(n20964), .A3(n16369), .ZN(n16358) );
  NAND2_X1 U17548 ( .A1(n20388), .A2(n14055), .ZN(n14385) );
  AOI21_X1 U17549 ( .B1(n14387), .B2(n14385), .A(n14056), .ZN(n14057) );
  NAND2_X1 U17550 ( .A1(n15304), .A2(n20363), .ZN(n16368) );
  NOR2_X1 U17551 ( .A1(n16368), .A2(n20383), .ZN(n14395) );
  AOI21_X1 U17552 ( .B1(n16358), .B2(n14057), .A(n14395), .ZN(n16362) );
  AND2_X1 U17553 ( .A1(n16358), .A2(n16370), .ZN(n14058) );
  AOI22_X1 U17554 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16362), .B1(
        n14058), .B2(n14053), .ZN(n14063) );
  OAI21_X1 U17555 ( .B1(n9821), .B2(n14059), .A(n13965), .ZN(n14060) );
  INV_X1 U17556 ( .A(n14060), .ZN(n20278) );
  INV_X1 U17557 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14061) );
  NOR2_X1 U17558 ( .A1(n20254), .A2(n14061), .ZN(n14065) );
  AOI21_X1 U17559 ( .B1(n20278), .B2(n20374), .A(n14065), .ZN(n14062) );
  OAI211_X1 U17560 ( .C1(n14070), .C2(n20385), .A(n14063), .B(n14062), .ZN(
        P1_U3022) );
  NOR2_X1 U17561 ( .A1(n15134), .A2(n20969), .ZN(n14064) );
  AOI211_X1 U17562 ( .C1(n16303), .C2(n20220), .A(n14065), .B(n14064), .ZN(
        n14069) );
  NAND2_X1 U17563 ( .A1(n20279), .A2(n14067), .ZN(n14068) );
  OAI211_X1 U17564 ( .C1(n14070), .C2(n20203), .A(n14069), .B(n14068), .ZN(
        P1_U2990) );
  AND2_X1 U17565 ( .A1(n14072), .A2(n14071), .ZN(n14073) );
  OR2_X1 U17566 ( .A1(n14073), .A2(n9809), .ZN(n15912) );
  MUX2_X1 U17567 ( .A(n15912), .B(n14074), .S(n9726), .Z(n14075) );
  OAI21_X1 U17568 ( .B1(n14076), .B2(n15539), .A(n14075), .ZN(P2_U2870) );
  AOI22_X1 U17569 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14080) );
  AOI22_X1 U17570 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14079) );
  AOI22_X1 U17571 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17572 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14077) );
  NAND4_X1 U17573 ( .A1(n14080), .A2(n14079), .A3(n14078), .A4(n14077), .ZN(
        n14086) );
  AOI22_X1 U17574 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14084) );
  AOI22_X1 U17575 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17576 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17577 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__4__SCAN_IN), .B2(n14508), .ZN(n14081) );
  NAND4_X1 U17578 ( .A1(n14084), .A2(n14083), .A3(n14082), .A4(n14081), .ZN(
        n14085) );
  NOR2_X1 U17579 ( .A1(n14086), .A2(n14085), .ZN(n14088) );
  AOI21_X1 U17580 ( .B1(n14088), .B2(n14087), .A(n9827), .ZN(n14089) );
  INV_X1 U17581 ( .A(n14089), .ZN(n15540) );
  OR2_X1 U17582 ( .A1(n14092), .A2(n14091), .ZN(n14093) );
  NAND2_X1 U17583 ( .A1(n14090), .A2(n14093), .ZN(n19187) );
  INV_X1 U17584 ( .A(n19187), .ZN(n15875) );
  OAI22_X1 U17585 ( .A1(n15577), .A2(n19526), .B1(n20897), .B2(n19387), .ZN(
        n14097) );
  INV_X1 U17586 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n14095) );
  INV_X1 U17587 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14094) );
  OAI22_X1 U17588 ( .A1(n15581), .A2(n14095), .B1(n15579), .B2(n14094), .ZN(
        n14096) );
  AOI211_X1 U17589 ( .C1(n19416), .C2(n15875), .A(n14097), .B(n14096), .ZN(
        n14098) );
  OAI21_X1 U17590 ( .B1(n15540), .B2(n19390), .A(n14098), .ZN(P2_U2899) );
  INV_X1 U17591 ( .A(n14100), .ZN(n14101) );
  NOR2_X1 U17592 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14101), .ZN(
        n14131) );
  INV_X1 U17593 ( .A(n14131), .ZN(n14143) );
  NOR3_X1 U17594 ( .A1(n14105), .A2(n12613), .A3(n20559), .ZN(n14102) );
  AOI21_X1 U17595 ( .B1(n14104), .B2(n14103), .A(n14102), .ZN(n14133) );
  INV_X1 U17596 ( .A(n14105), .ZN(n20551) );
  AOI21_X1 U17597 ( .B1(n20562), .B2(n14106), .A(n20818), .ZN(n14107) );
  AOI21_X1 U17598 ( .B1(n20551), .B2(n15333), .A(n14107), .ZN(n14108) );
  NOR2_X1 U17599 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n14108), .ZN(n14110) );
  OAI211_X1 U17600 ( .C1(n14131), .C2(n14110), .A(n20454), .B(n14109), .ZN(
        n14140) );
  AOI22_X1 U17601 ( .A1(n14141), .A2(n20579), .B1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .B2(n14140), .ZN(n14111) );
  OAI21_X1 U17602 ( .B1(n14112), .B2(n14143), .A(n14111), .ZN(n14113) );
  AOI21_X1 U17603 ( .B1(n14146), .B2(n20581), .A(n14113), .ZN(n14114) );
  OAI21_X1 U17604 ( .B1(n20584), .B2(n20562), .A(n14114), .ZN(P1_U3148) );
  AOI22_X1 U17605 ( .A1(n14141), .A2(n20567), .B1(
        P1_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n14140), .ZN(n14115) );
  OAI21_X1 U17606 ( .B1(n14116), .B2(n14143), .A(n14115), .ZN(n14117) );
  AOI21_X1 U17607 ( .B1(n14146), .B2(n20569), .A(n14117), .ZN(n14118) );
  OAI21_X1 U17608 ( .B1(n20572), .B2(n20562), .A(n14118), .ZN(P1_U3146) );
  AOI22_X1 U17609 ( .A1(n14141), .A2(n20591), .B1(
        P1_INSTQUEUE_REG_14__5__SCAN_IN), .B2(n14140), .ZN(n14119) );
  OAI21_X1 U17610 ( .B1(n14120), .B2(n14143), .A(n14119), .ZN(n14121) );
  AOI21_X1 U17611 ( .B1(n14146), .B2(n20593), .A(n14121), .ZN(n14122) );
  OAI21_X1 U17612 ( .B1(n20596), .B2(n20562), .A(n14122), .ZN(P1_U3150) );
  AOI22_X1 U17613 ( .A1(n14141), .A2(n20573), .B1(
        P1_INSTQUEUE_REG_14__2__SCAN_IN), .B2(n14140), .ZN(n14123) );
  OAI21_X1 U17614 ( .B1(n14124), .B2(n14143), .A(n14123), .ZN(n14125) );
  AOI21_X1 U17615 ( .B1(n14146), .B2(n20575), .A(n14125), .ZN(n14126) );
  OAI21_X1 U17616 ( .B1(n20578), .B2(n20562), .A(n14126), .ZN(P1_U3147) );
  AOI22_X1 U17617 ( .A1(n14141), .A2(n20604), .B1(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .B2(n14140), .ZN(n14127) );
  OAI21_X1 U17618 ( .B1(n14128), .B2(n14143), .A(n14127), .ZN(n14129) );
  AOI21_X1 U17619 ( .B1(n14146), .B2(n20607), .A(n14129), .ZN(n14130) );
  OAI21_X1 U17620 ( .B1(n20613), .B2(n20562), .A(n14130), .ZN(P1_U3152) );
  AOI22_X1 U17621 ( .A1(n20598), .A2(n14131), .B1(
        P1_INSTQUEUE_REG_14__6__SCAN_IN), .B2(n14140), .ZN(n14132) );
  OAI21_X1 U17622 ( .B1(n14133), .B2(n14165), .A(n14132), .ZN(n14134) );
  AOI21_X1 U17623 ( .B1(n14146), .B2(n20599), .A(n14134), .ZN(n14135) );
  OAI21_X1 U17624 ( .B1(n20602), .B2(n20562), .A(n14135), .ZN(P1_U3151) );
  AOI22_X1 U17625 ( .A1(n14141), .A2(n20553), .B1(
        P1_INSTQUEUE_REG_14__0__SCAN_IN), .B2(n14140), .ZN(n14136) );
  OAI21_X1 U17626 ( .B1(n14137), .B2(n14143), .A(n14136), .ZN(n14138) );
  AOI21_X1 U17627 ( .B1(n14146), .B2(n20563), .A(n14138), .ZN(n14139) );
  OAI21_X1 U17628 ( .B1(n20566), .B2(n20562), .A(n14139), .ZN(P1_U3145) );
  AOI22_X1 U17629 ( .A1(n14141), .A2(n20585), .B1(
        P1_INSTQUEUE_REG_14__4__SCAN_IN), .B2(n14140), .ZN(n14142) );
  OAI21_X1 U17630 ( .B1(n14144), .B2(n14143), .A(n14142), .ZN(n14145) );
  AOI21_X1 U17631 ( .B1(n14146), .B2(n20587), .A(n14145), .ZN(n14147) );
  OAI21_X1 U17632 ( .B1(n20590), .B2(n20562), .A(n14147), .ZN(P1_U3149) );
  NAND2_X1 U17633 ( .A1(n14193), .A2(n20561), .ZN(n14151) );
  OAI21_X1 U17634 ( .B1(n14151), .B2(n20443), .A(n14150), .ZN(n14160) );
  NOR2_X1 U17635 ( .A1(n14152), .A2(n12613), .ZN(n14156) );
  NOR2_X1 U17636 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14155), .ZN(
        n14191) );
  INV_X1 U17637 ( .A(n14156), .ZN(n14159) );
  AOI211_X1 U17638 ( .C1(n14160), .C2(n14159), .A(n14158), .B(n14157), .ZN(
        n14161) );
  AOI22_X1 U17639 ( .A1(n20598), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n14190), .ZN(n14162) );
  OAI21_X1 U17640 ( .B1(n20484), .B2(n14193), .A(n14162), .ZN(n14163) );
  AOI21_X1 U17641 ( .B1(n20443), .B2(n20481), .A(n14163), .ZN(n14164) );
  OAI21_X1 U17642 ( .B1(n14197), .B2(n14165), .A(n14164), .ZN(P1_U3055) );
  AOI22_X1 U17643 ( .A1(n20554), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__0__SCAN_IN), .B2(n14190), .ZN(n14166) );
  OAI21_X1 U17644 ( .B1(n14193), .B2(n20460), .A(n14166), .ZN(n14167) );
  AOI21_X1 U17645 ( .B1(n20443), .B2(n20457), .A(n14167), .ZN(n14168) );
  OAI21_X1 U17646 ( .B1(n14197), .B2(n14169), .A(n14168), .ZN(P1_U3049) );
  AOI22_X1 U17647 ( .A1(n20568), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n14190), .ZN(n14170) );
  OAI21_X1 U17648 ( .B1(n14193), .B2(n20464), .A(n14170), .ZN(n14171) );
  AOI21_X1 U17649 ( .B1(n20443), .B2(n20461), .A(n14171), .ZN(n14172) );
  OAI21_X1 U17650 ( .B1(n14197), .B2(n14173), .A(n14172), .ZN(P1_U3050) );
  AOI22_X1 U17651 ( .A1(n20580), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n14190), .ZN(n14174) );
  OAI21_X1 U17652 ( .B1(n14193), .B2(n20472), .A(n14174), .ZN(n14175) );
  AOI21_X1 U17653 ( .B1(n20443), .B2(n20469), .A(n14175), .ZN(n14176) );
  OAI21_X1 U17654 ( .B1(n14197), .B2(n14177), .A(n14176), .ZN(P1_U3052) );
  AOI22_X1 U17655 ( .A1(n20606), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14190), .ZN(n14178) );
  OAI21_X1 U17656 ( .B1(n14193), .B2(n20492), .A(n14178), .ZN(n14179) );
  AOI21_X1 U17657 ( .B1(n20443), .B2(n20487), .A(n14179), .ZN(n14180) );
  OAI21_X1 U17658 ( .B1(n14197), .B2(n14181), .A(n14180), .ZN(P1_U3056) );
  AOI22_X1 U17659 ( .A1(n20574), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n14190), .ZN(n14182) );
  OAI21_X1 U17660 ( .B1(n14193), .B2(n20468), .A(n14182), .ZN(n14183) );
  AOI21_X1 U17661 ( .B1(n20443), .B2(n20465), .A(n14183), .ZN(n14184) );
  OAI21_X1 U17662 ( .B1(n14197), .B2(n14185), .A(n14184), .ZN(P1_U3051) );
  AOI22_X1 U17663 ( .A1(n20592), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n14190), .ZN(n14186) );
  OAI21_X1 U17664 ( .B1(n14193), .B2(n20480), .A(n14186), .ZN(n14187) );
  AOI21_X1 U17665 ( .B1(n20443), .B2(n20477), .A(n14187), .ZN(n14188) );
  OAI21_X1 U17666 ( .B1(n14197), .B2(n14189), .A(n14188), .ZN(P1_U3054) );
  AOI22_X1 U17667 ( .A1(n20586), .A2(n14191), .B1(
        P1_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n14190), .ZN(n14192) );
  OAI21_X1 U17668 ( .B1(n14193), .B2(n20476), .A(n14192), .ZN(n14194) );
  AOI21_X1 U17669 ( .B1(n20443), .B2(n20473), .A(n14194), .ZN(n14195) );
  OAI21_X1 U17670 ( .B1(n14197), .B2(n14196), .A(n14195), .ZN(P1_U3053) );
  NOR2_X1 U17671 ( .A1(n9809), .A2(n14199), .ZN(n14200) );
  OR2_X1 U17672 ( .A1(n14198), .A2(n14200), .ZN(n19206) );
  MUX2_X1 U17673 ( .A(n19206), .B(n19202), .S(n9726), .Z(n14201) );
  OAI21_X1 U17674 ( .B1(n14202), .B2(n15539), .A(n14201), .ZN(P2_U2869) );
  INV_X1 U17675 ( .A(n14203), .ZN(n14210) );
  AOI22_X1 U17676 ( .A1(n19339), .A2(n14204), .B1(n19342), .B2(
        P2_EBX_REG_17__SCAN_IN), .ZN(n14205) );
  OAI21_X1 U17677 ( .B1(n15912), .B2(n19346), .A(n14205), .ZN(n14209) );
  NAND2_X1 U17678 ( .A1(n15705), .A2(n14214), .ZN(n14206) );
  AND2_X1 U17679 ( .A1(n14206), .A2(n10009), .ZN(n15708) );
  INV_X1 U17680 ( .A(n15708), .ZN(n14217) );
  NAND2_X1 U17681 ( .A1(n19331), .A2(n19316), .ZN(n15470) );
  INV_X1 U17682 ( .A(n19305), .ZN(n19343) );
  AOI22_X1 U17683 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19343), .ZN(n14207) );
  OAI211_X1 U17684 ( .C1(n14217), .C2(n15470), .A(n14207), .B(n19304), .ZN(
        n14208) );
  AOI211_X1 U17685 ( .C1(n19341), .C2(n14210), .A(n14209), .B(n14208), .ZN(
        n14220) );
  AOI21_X1 U17686 ( .B1(n14212), .B2(n19228), .A(n14215), .ZN(n19226) );
  NOR2_X1 U17687 ( .A1(n15746), .A2(n14211), .ZN(n19240) );
  OAI21_X1 U17688 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n14213), .A(
        n14212), .ZN(n19241) );
  NAND2_X1 U17689 ( .A1(n19240), .A2(n19241), .ZN(n19225) );
  NOR2_X1 U17690 ( .A1(n19226), .A2(n19225), .ZN(n19217) );
  OAI21_X1 U17691 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n14215), .A(
        n14214), .ZN(n19218) );
  NAND2_X1 U17692 ( .A1(n19217), .A2(n19218), .ZN(n14216) );
  INV_X1 U17693 ( .A(n14216), .ZN(n14218) );
  NOR2_X1 U17694 ( .A1(n15708), .A2(n14216), .ZN(n15355) );
  NOR2_X1 U17695 ( .A1(n19331), .A2(n15355), .ZN(n19208) );
  OAI211_X1 U17696 ( .C1(n14218), .C2(n14217), .A(n19208), .B(n19316), .ZN(
        n14219) );
  NAND2_X1 U17697 ( .A1(n14220), .A2(n14219), .ZN(P2_U2838) );
  OAI21_X1 U17698 ( .B1(n14198), .B2(n14222), .A(n15533), .ZN(n19195) );
  NOR2_X1 U17699 ( .A1(n19195), .A2(n9726), .ZN(n14223) );
  AOI21_X1 U17700 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n9726), .A(n14223), .ZN(
        n14224) );
  OAI21_X1 U17701 ( .B1(n14225), .B2(n15539), .A(n14224), .ZN(P2_U2868) );
  INV_X1 U17702 ( .A(n13955), .ZN(n14227) );
  OAI21_X1 U17703 ( .B1(n14227), .B2(n11887), .A(n14253), .ZN(n14255) );
  XOR2_X1 U17704 ( .A(n14254), .B(n14255), .Z(n16310) );
  INV_X1 U17705 ( .A(n16310), .ZN(n14297) );
  MUX2_X1 U17706 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n14279), .Z(
        n20328) );
  AOI22_X1 U17707 ( .A1(n14232), .A2(n20328), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n16280), .ZN(n14228) );
  OAI21_X1 U17708 ( .B1(n14297), .B2(n16283), .A(n14228), .ZN(P1_U2893) );
  INV_X1 U17709 ( .A(n14229), .ZN(n14231) );
  INV_X1 U17710 ( .A(n14230), .ZN(n14256) );
  AOI21_X1 U17711 ( .B1(n14231), .B2(n14256), .A(n9800), .ZN(n16304) );
  INV_X1 U17712 ( .A(n16304), .ZN(n14234) );
  MUX2_X1 U17713 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n14279), .Z(
        n20332) );
  AOI22_X1 U17714 ( .A1(n14232), .A2(n20332), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n16280), .ZN(n14233) );
  OAI21_X1 U17715 ( .B1(n14234), .B2(n16283), .A(n14233), .ZN(P1_U2890) );
  MUX2_X1 U17716 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n14235) );
  OAI21_X1 U17717 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14342), .A(
        n14235), .ZN(n14294) );
  OAI21_X1 U17718 ( .B1(n14308), .B2(n15313), .A(n14238), .ZN(n14239) );
  INV_X1 U17719 ( .A(n14239), .ZN(n14241) );
  MUX2_X1 U17720 ( .A(n13168), .B(n14335), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n14240) );
  NAND2_X1 U17721 ( .A1(n14241), .A2(n14240), .ZN(n15306) );
  MUX2_X1 U17722 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n14243) );
  OR2_X1 U17723 ( .A1(n14342), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14242) );
  NAND2_X1 U17724 ( .A1(n15309), .A2(n14258), .ZN(n14248) );
  OR2_X1 U17725 ( .A1(n13168), .A2(P1_EBX_REG_14__SCAN_IN), .ZN(n14247) );
  NAND2_X1 U17726 ( .A1(n13438), .A2(n20883), .ZN(n14245) );
  INV_X1 U17727 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n20984) );
  NAND2_X1 U17728 ( .A1(n14308), .A2(n20984), .ZN(n14244) );
  NAND3_X1 U17729 ( .A1(n14245), .A2(n14313), .A3(n14244), .ZN(n14246) );
  OR2_X2 U17730 ( .A1(n14248), .A2(n14249), .ZN(n14275) );
  NAND2_X1 U17731 ( .A1(n14248), .A2(n14249), .ZN(n14250) );
  NAND2_X1 U17732 ( .A1(n14275), .A2(n14250), .ZN(n16341) );
  OAI22_X1 U17733 ( .A1(n16341), .A2(n14936), .B1(n20984), .B2(n20282), .ZN(
        n14251) );
  AOI21_X1 U17734 ( .B1(n16304), .B2(n20708), .A(n14251), .ZN(n14252) );
  INV_X1 U17735 ( .A(n14252), .ZN(P1_U2858) );
  OAI21_X1 U17736 ( .B1(n14255), .B2(n14254), .A(n14253), .ZN(n14285) );
  INV_X1 U17737 ( .A(n15125), .ZN(n14268) );
  INV_X1 U17738 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14261) );
  OAI21_X1 U17739 ( .B1(n15309), .B2(n14258), .A(n14248), .ZN(n15300) );
  INV_X1 U17740 ( .A(n15300), .ZN(n14259) );
  AOI22_X1 U17741 ( .A1(n14259), .A2(n20253), .B1(n20263), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14260) );
  OAI211_X1 U17742 ( .C1(n20257), .C2(n14261), .A(n14260), .B(n20254), .ZN(
        n14267) );
  NAND2_X1 U17743 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n14345) );
  NOR2_X1 U17744 ( .A1(n16371), .A2(n14262), .ZN(n20224) );
  NAND3_X1 U17745 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n20224), .ZN(n16279) );
  NOR2_X1 U17746 ( .A1(n14345), .A2(n16279), .ZN(n14265) );
  INV_X1 U17747 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20644) );
  NOR2_X1 U17748 ( .A1(n20644), .A2(n14061), .ZN(n14263) );
  OAI21_X1 U17749 ( .B1(n14263), .B2(n20271), .A(n20227), .ZN(n16276) );
  AOI21_X1 U17750 ( .B1(n16239), .B2(n14345), .A(n16276), .ZN(n16270) );
  INV_X1 U17751 ( .A(n16270), .ZN(n14264) );
  MUX2_X1 U17752 ( .A(n14265), .B(n14264), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14266) );
  AOI211_X1 U17753 ( .C1(n20221), .C2(n14268), .A(n14267), .B(n14266), .ZN(
        n14269) );
  OAI21_X1 U17754 ( .B1(n20242), .B2(n15129), .A(n14269), .ZN(P1_U2827) );
  OAI21_X1 U17755 ( .B1(n9800), .B2(n11962), .A(n14271), .ZN(n16252) );
  NAND2_X1 U17756 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14272) );
  OAI211_X1 U17757 ( .C1(n14341), .C2(P1_EBX_REG_15__SCAN_IN), .A(n14335), .B(
        n14272), .ZN(n14273) );
  OAI21_X1 U17758 ( .B1(n14332), .B2(P1_EBX_REG_15__SCAN_IN), .A(n14273), .ZN(
        n14274) );
  AND2_X1 U17759 ( .A1(n14275), .A2(n14274), .ZN(n14276) );
  NOR2_X1 U17760 ( .A1(n14934), .A2(n14276), .ZN(n16335) );
  INV_X1 U17761 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n20918) );
  NOR2_X1 U17762 ( .A1(n20282), .A2(n20918), .ZN(n14277) );
  AOI21_X1 U17763 ( .B1(n16335), .B2(n20706), .A(n14277), .ZN(n14278) );
  OAI21_X1 U17764 ( .B1(n16252), .B2(n14939), .A(n14278), .ZN(P1_U2857) );
  MUX2_X1 U17765 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n14279), .Z(
        n20330) );
  INV_X1 U17766 ( .A(n20330), .ZN(n14281) );
  OAI222_X1 U17767 ( .A1(n15129), .A2(n16283), .B1(n14293), .B2(n14281), .C1(
        n14280), .C2(n14290), .ZN(P1_U2891) );
  INV_X1 U17768 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14282) );
  OAI222_X1 U17769 ( .A1(n15300), .A2(n14936), .B1(n14282), .B2(n20282), .C1(
        n15129), .C2(n14939), .ZN(P1_U2859) );
  OAI222_X1 U17770 ( .A1(n16252), .A2(n16283), .B1(n14293), .B2(n14284), .C1(
        n14290), .C2(n14283), .ZN(P1_U2889) );
  INV_X1 U17771 ( .A(n14285), .ZN(n14289) );
  INV_X1 U17772 ( .A(n14286), .ZN(n14288) );
  INV_X1 U17773 ( .A(n20709), .ZN(n15138) );
  INV_X1 U17774 ( .A(n14948), .ZN(n14292) );
  OAI222_X1 U17775 ( .A1(n15138), .A2(n16283), .B1(n14293), .B2(n14292), .C1(
        n14291), .C2(n14290), .ZN(P1_U2892) );
  AND2_X1 U17776 ( .A1(n14295), .A2(n14294), .ZN(n14296) );
  OR2_X1 U17777 ( .A1(n14296), .A2(n15307), .ZN(n16350) );
  INV_X1 U17778 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n16271) );
  OAI222_X1 U17779 ( .A1(n16350), .A2(n14936), .B1(n16271), .B2(n20282), .C1(
        n14939), .C2(n14297), .ZN(P1_U2861) );
  OAI211_X1 U17780 ( .C1(n19085), .C2(n18948), .A(n12156), .B(n16143), .ZN(
        n18465) );
  NOR2_X1 U17781 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18465), .ZN(n14298) );
  NAND3_X1 U17782 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n19077)
         );
  OAI21_X1 U17783 ( .B1(n14298), .B2(n19077), .A(n18562), .ZN(n18471) );
  INV_X1 U17784 ( .A(n18471), .ZN(n18477) );
  NOR2_X1 U17785 ( .A1(n19127), .A2(n18121), .ZN(n18469) );
  AOI21_X1 U17786 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18469), .ZN(n18470) );
  NOR2_X1 U17787 ( .A1(n18477), .A2(n18470), .ZN(n14300) );
  INV_X1 U17788 ( .A(n18722), .ZN(n18482) );
  NOR2_X1 U17789 ( .A1(n19079), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18520) );
  OR2_X1 U17790 ( .A1(n18520), .A2(n18477), .ZN(n18468) );
  OR2_X1 U17791 ( .A1(n18482), .A2(n18468), .ZN(n14299) );
  MUX2_X1 U17792 ( .A(n14300), .B(n14299), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AND2_X1 U17793 ( .A1(n14341), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14301) );
  AOI21_X1 U17794 ( .B1(n14342), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14301), .ZN(
        n14706) );
  OR2_X1 U17795 ( .A1(n13168), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n14305) );
  INV_X1 U17796 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15285) );
  NAND2_X1 U17797 ( .A1(n14335), .A2(n15285), .ZN(n14303) );
  INV_X1 U17798 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16240) );
  NAND2_X1 U17799 ( .A1(n14308), .A2(n16240), .ZN(n14302) );
  NAND3_X1 U17800 ( .A1(n14303), .A2(n14313), .A3(n14302), .ZN(n14304) );
  NAND2_X1 U17801 ( .A1(n14305), .A2(n14304), .ZN(n14933) );
  MUX2_X1 U17802 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n14307) );
  OR2_X1 U17803 ( .A1(n14342), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14306) );
  AND2_X1 U17804 ( .A1(n14307), .A2(n14306), .ZN(n14864) );
  NAND2_X1 U17805 ( .A1(n14863), .A2(n14864), .ZN(n14862) );
  OR2_X1 U17806 ( .A1(n13168), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14312) );
  INV_X1 U17807 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15080) );
  NAND2_X1 U17808 ( .A1(n14335), .A2(n15080), .ZN(n14310) );
  INV_X1 U17809 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14927) );
  NAND2_X1 U17810 ( .A1(n14308), .A2(n14927), .ZN(n14309) );
  NAND3_X1 U17811 ( .A1(n14310), .A2(n14313), .A3(n14309), .ZN(n14311) );
  AND2_X1 U17812 ( .A1(n14312), .A2(n14311), .ZN(n14924) );
  NAND2_X1 U17813 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14314) );
  OAI211_X1 U17814 ( .C1(n14341), .C2(P1_EBX_REG_19__SCAN_IN), .A(n14335), .B(
        n14314), .ZN(n14315) );
  OAI21_X1 U17815 ( .B1(n14332), .B2(P1_EBX_REG_19__SCAN_IN), .A(n14315), .ZN(
        n14842) );
  MUX2_X1 U17816 ( .A(n13168), .B(n14335), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14317) );
  NAND2_X1 U17817 ( .A1(n14341), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14316) );
  NAND2_X1 U17818 ( .A1(n14317), .A2(n14316), .ZN(n14912) );
  MUX2_X1 U17819 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14318) );
  OAI21_X1 U17820 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14342), .A(
        n14318), .ZN(n14830) );
  OR2_X1 U17821 ( .A1(n13168), .A2(P1_EBX_REG_22__SCAN_IN), .ZN(n14321) );
  INV_X1 U17822 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15237) );
  NAND2_X1 U17823 ( .A1(n14335), .A2(n15237), .ZN(n14319) );
  OAI211_X1 U17824 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n14341), .A(n14319), .B(
        n14313), .ZN(n14320) );
  AND2_X1 U17825 ( .A1(n14321), .A2(n14320), .ZN(n14812) );
  MUX2_X1 U17826 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14322) );
  OAI21_X1 U17827 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14342), .A(
        n14322), .ZN(n14794) );
  OR2_X1 U17828 ( .A1(n13168), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14325) );
  NAND2_X1 U17829 ( .A1(n14335), .A2(n15209), .ZN(n14323) );
  OAI211_X1 U17830 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n14341), .A(n14323), .B(
        n14313), .ZN(n14324) );
  NAND2_X1 U17831 ( .A1(n14325), .A2(n14324), .ZN(n14784) );
  INV_X1 U17832 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14907) );
  NAND2_X1 U17833 ( .A1(n14326), .A2(n14907), .ZN(n14329) );
  NAND2_X1 U17834 ( .A1(n14313), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14327) );
  OAI211_X1 U17835 ( .C1(n14341), .C2(P1_EBX_REG_25__SCAN_IN), .A(n14335), .B(
        n14327), .ZN(n14328) );
  AND2_X1 U17836 ( .A1(n14329), .A2(n14328), .ZN(n14771) );
  MUX2_X1 U17837 ( .A(n13168), .B(n13438), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14331) );
  NAND2_X1 U17838 ( .A1(n14341), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14330) );
  AND2_X1 U17839 ( .A1(n14331), .A2(n14330), .ZN(n14760) );
  MUX2_X1 U17840 ( .A(n14332), .B(n14313), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14333) );
  OAI21_X1 U17841 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14342), .A(
        n14333), .ZN(n14745) );
  INV_X1 U17842 ( .A(n13168), .ZN(n14338) );
  INV_X1 U17843 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14337) );
  INV_X1 U17844 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14378) );
  NOR2_X1 U17845 ( .A1(n14341), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14334) );
  AOI211_X1 U17846 ( .C1(n14335), .C2(n14378), .A(n14705), .B(n14334), .ZN(
        n14336) );
  AOI21_X1 U17847 ( .B1(n14338), .B2(n14337), .A(n14336), .ZN(n14730) );
  NOR2_X1 U17848 ( .A1(n14341), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14340) );
  INV_X1 U17849 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15158) );
  AOI21_X1 U17850 ( .B1(n14339), .B2(n15158), .A(n14340), .ZN(n14704) );
  MUX2_X1 U17851 ( .A(n14340), .B(n14704), .S(n14313), .Z(n14719) );
  NAND2_X1 U17852 ( .A1(n14729), .A2(n14719), .ZN(n14718) );
  MUX2_X1 U17853 ( .A(n14706), .B(n14313), .S(n14718), .Z(n14344) );
  AOI22_X1 U17854 ( .A1(n14342), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14341), .ZN(n14343) );
  XNOR2_X2 U17855 ( .A(n14344), .B(n14343), .ZN(n14901) );
  NAND2_X1 U17856 ( .A1(n14416), .A2(n20233), .ZN(n14358) );
  NAND2_X1 U17857 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14354) );
  INV_X1 U17858 ( .A(n14354), .ZN(n14350) );
  NAND2_X1 U17859 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14349) );
  NAND3_X1 U17860 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .A3(P1_REIP_REG_24__SCAN_IN), .ZN(n14353) );
  INV_X1 U17861 ( .A(n14353), .ZN(n14348) );
  INV_X1 U17862 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20649) );
  NOR2_X1 U17863 ( .A1(n20649), .A2(n14345), .ZN(n16257) );
  NAND4_X1 U17864 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(n16257), .ZN(n16238) );
  NAND2_X1 U17865 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16243) );
  NAND4_X1 U17866 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(P1_REIP_REG_8__SCAN_IN), .A4(P1_REIP_REG_7__SCAN_IN), .ZN(n14346)
         );
  NOR4_X1 U17867 ( .A1(n20249), .A2(n16238), .A3(n16243), .A4(n14346), .ZN(
        n14857) );
  NAND2_X1 U17868 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n14857), .ZN(n16227) );
  NAND2_X1 U17869 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n14849) );
  NOR2_X1 U17870 ( .A1(n16227), .A2(n14849), .ZN(n14813) );
  INV_X1 U17871 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20661) );
  NAND2_X1 U17872 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n14816) );
  NOR2_X1 U17873 ( .A1(n20661), .A2(n14816), .ZN(n14801) );
  AND2_X1 U17874 ( .A1(n14801), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14352) );
  NAND3_X1 U17875 ( .A1(n14845), .A2(n14813), .A3(n14352), .ZN(n14347) );
  NAND2_X1 U17876 ( .A1(n14847), .A2(n14347), .ZN(n14802) );
  OAI21_X1 U17877 ( .B1(n20271), .B2(n14348), .A(n14802), .ZN(n14761) );
  AOI21_X1 U17878 ( .B1(n14349), .B2(n14847), .A(n14761), .ZN(n14737) );
  OAI21_X1 U17879 ( .B1(n20252), .B2(n14350), .A(n14737), .ZN(n14714) );
  INV_X1 U17880 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14900) );
  INV_X1 U17881 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14351) );
  OAI22_X1 U17882 ( .A1(n16272), .A2(n14900), .B1(n14351), .B2(n20257), .ZN(
        n14356) );
  NAND2_X1 U17883 ( .A1(n16219), .A2(n14352), .ZN(n14788) );
  NOR2_X1 U17884 ( .A1(n14788), .A2(n14353), .ZN(n14746) );
  NAND3_X1 U17885 ( .A1(n14746), .A2(P1_REIP_REG_28__SCAN_IN), .A3(
        P1_REIP_REG_27__SCAN_IN), .ZN(n14722) );
  NOR3_X1 U17886 ( .A1(n14722), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14354), 
        .ZN(n14355) );
  AOI211_X1 U17887 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14714), .A(n14356), 
        .B(n14355), .ZN(n14357) );
  OAI211_X1 U17888 ( .C1(n14901), .C2(n20267), .A(n14358), .B(n14357), .ZN(
        P1_U2809) );
  AOI21_X1 U17889 ( .B1(n15334), .B2(n16159), .A(n14363), .ZN(n14365) );
  NAND2_X1 U17890 ( .A1(n11787), .A2(n15332), .ZN(n14361) );
  NAND2_X1 U17891 ( .A1(n14359), .A2(n11224), .ZN(n14360) );
  NAND2_X1 U17892 ( .A1(n14361), .A2(n14360), .ZN(n16161) );
  OAI22_X1 U17893 ( .A1(n20614), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15335), .ZN(n14362) );
  AOI21_X1 U17894 ( .B1(n16161), .B2(n15334), .A(n14362), .ZN(n14364) );
  OAI22_X1 U17895 ( .A1(n14365), .A2(n11224), .B1(n14364), .B2(n14363), .ZN(
        P1_U3474) );
  NOR2_X1 U17896 ( .A1(n15488), .A2(n13256), .ZN(n14370) );
  INV_X1 U17897 ( .A(n15349), .ZN(n14366) );
  OAI21_X1 U17898 ( .B1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n14366), .A(
        n10000), .ZN(n16437) );
  NAND2_X1 U17899 ( .A1(n19473), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14367) );
  OAI211_X1 U17900 ( .C1(n16437), .C2(n19471), .A(n14368), .B(n14367), .ZN(
        n14369) );
  AOI211_X1 U17901 ( .C1(n14371), .C2(n19475), .A(n14370), .B(n14369), .ZN(
        n14372) );
  OAI21_X1 U17902 ( .B1(n14373), .B2(n16514), .A(n14372), .ZN(P2_U2986) );
  NAND2_X1 U17903 ( .A1(n14375), .A2(n11601), .ZN(n15026) );
  NAND3_X1 U17904 ( .A1(n14376), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15026), .ZN(n14377) );
  AND2_X1 U17905 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15171) );
  INV_X1 U17906 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14379) );
  NAND2_X1 U17907 ( .A1(n14379), .A2(n14378), .ZN(n15169) );
  OAI21_X1 U17908 ( .B1(n14989), .B2(n15169), .A(n15097), .ZN(n14380) );
  NAND2_X1 U17909 ( .A1(n14381), .A2(n14380), .ZN(n14999) );
  INV_X1 U17910 ( .A(n14999), .ZN(n14383) );
  NAND2_X1 U17911 ( .A1(n15097), .A2(n15158), .ZN(n15001) );
  NAND2_X1 U17912 ( .A1(n11601), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15000) );
  NOR2_X1 U17913 ( .A1(n14381), .A2(n15000), .ZN(n14990) );
  AOI22_X1 U17914 ( .A1(n14383), .A2(n14382), .B1(n14990), .B2(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14384) );
  XNOR2_X1 U17915 ( .A(n14384), .B(n14401), .ZN(n14418) );
  NOR2_X1 U17916 ( .A1(n14901), .A2(n20392), .ZN(n14410) );
  INV_X1 U17917 ( .A(n16368), .ZN(n15325) );
  NAND3_X1 U17918 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16358), .ZN(n16357) );
  NOR2_X1 U17919 ( .A1(n14385), .A2(n16357), .ZN(n15303) );
  NAND3_X1 U17920 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15303), .ZN(n15235) );
  NOR2_X1 U17921 ( .A1(n15231), .A2(n15235), .ZN(n14402) );
  INV_X1 U17922 ( .A(n14402), .ZN(n14386) );
  AOI21_X1 U17923 ( .B1(n14387), .B2(n14386), .A(n20383), .ZN(n14392) );
  INV_X1 U17924 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16349) );
  NOR4_X1 U17925 ( .A1(n15313), .A2(n16349), .A3(n16357), .A4(n14388), .ZN(
        n15229) );
  NAND2_X1 U17926 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15229), .ZN(
        n16340) );
  INV_X1 U17927 ( .A(n16340), .ZN(n14389) );
  OR2_X1 U17928 ( .A1(n20363), .A2(n14389), .ZN(n14390) );
  NOR2_X1 U17929 ( .A1(n11602), .A2(n15285), .ZN(n16327) );
  NAND4_X1 U17930 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(n16327), .ZN(n15230) );
  INV_X1 U17931 ( .A(n15230), .ZN(n14391) );
  NAND2_X1 U17932 ( .A1(n16348), .A2(n14391), .ZN(n14394) );
  NAND2_X1 U17933 ( .A1(n15325), .A2(n14392), .ZN(n14393) );
  NAND2_X1 U17934 ( .A1(n14394), .A2(n14393), .ZN(n15261) );
  NAND2_X1 U17935 ( .A1(n15261), .A2(n9856), .ZN(n14397) );
  INV_X1 U17936 ( .A(n14395), .ZN(n14396) );
  NAND2_X1 U17937 ( .A1(n14397), .A2(n14396), .ZN(n15228) );
  NAND2_X1 U17938 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14404) );
  NAND2_X1 U17939 ( .A1(n16368), .A2(n14404), .ZN(n14398) );
  NAND2_X1 U17940 ( .A1(n15228), .A2(n14398), .ZN(n15221) );
  AOI21_X1 U17941 ( .B1(n20389), .B2(n20816), .A(n15221), .ZN(n15211) );
  OAI21_X1 U17942 ( .B1(n15188), .B2(n15325), .A(n15211), .ZN(n15187) );
  INV_X1 U17943 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15190) );
  NOR3_X1 U17944 ( .A1(n15187), .A2(n15202), .A3(n15190), .ZN(n14399) );
  NOR2_X1 U17945 ( .A1(n15221), .A2(n16368), .ZN(n15161) );
  NOR2_X1 U17946 ( .A1(n14399), .A2(n15161), .ZN(n15181) );
  NOR2_X1 U17947 ( .A1(n15181), .A2(n15158), .ZN(n15160) );
  AOI21_X1 U17948 ( .B1(n15160), .B2(n15171), .A(n15161), .ZN(n14400) );
  INV_X1 U17949 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15151) );
  NOR2_X1 U17950 ( .A1(n14400), .A2(n15151), .ZN(n15149) );
  NOR3_X1 U17951 ( .A1(n15149), .A2(n15161), .A3(n14401), .ZN(n14409) );
  INV_X1 U17952 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20986) );
  NOR2_X1 U17953 ( .A1(n20254), .A2(n20986), .ZN(n14412) );
  OR2_X1 U17954 ( .A1(n20363), .A2(n16340), .ZN(n14403) );
  NAND2_X1 U17955 ( .A1(n14402), .A2(n20382), .ZN(n15208) );
  NAND2_X1 U17956 ( .A1(n14403), .A2(n15208), .ZN(n15269) );
  INV_X1 U17957 ( .A(n14404), .ZN(n15236) );
  NAND2_X1 U17958 ( .A1(n9856), .A2(n15236), .ZN(n14405) );
  NOR2_X1 U17959 ( .A1(n14405), .A2(n15230), .ZN(n14406) );
  NOR2_X1 U17960 ( .A1(n15186), .A2(n15190), .ZN(n14407) );
  NAND3_X1 U17961 ( .A1(n15157), .A2(n15171), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15150) );
  NOR3_X1 U17962 ( .A1(n15150), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15151), .ZN(n14408) );
  NOR4_X2 U17963 ( .A1(n14410), .A2(n14409), .A3(n14412), .A4(n14408), .ZN(
        n14411) );
  OAI21_X1 U17964 ( .B1(n14418), .B2(n20385), .A(n14411), .ZN(P1_U3000) );
  AOI21_X1 U17965 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14412), .ZN(n14413) );
  OAI21_X1 U17966 ( .B1(n20361), .B2(n14414), .A(n14413), .ZN(n14415) );
  AOI21_X1 U17967 ( .B1(n14416), .B2(n14067), .A(n14415), .ZN(n14417) );
  OAI21_X1 U17968 ( .B1(n14418), .B2(n20203), .A(n14417), .ZN(P1_U2968) );
  OAI21_X1 U17969 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14427) );
  NOR2_X1 U17970 ( .A1(n14422), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14423) );
  MUX2_X1 U17971 ( .A(n14424), .B(n14423), .S(n11197), .Z(n16409) );
  NAND2_X1 U17972 ( .A1(n16409), .A2(n10626), .ZN(n14425) );
  XNOR2_X1 U17973 ( .A(n14425), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14426) );
  XNOR2_X1 U17974 ( .A(n14427), .B(n14426), .ZN(n14461) );
  INV_X1 U17975 ( .A(n14429), .ZN(n14434) );
  INV_X1 U17976 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16414) );
  NAND2_X1 U17977 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U17978 ( .A1(n9725), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14430) );
  OAI211_X1 U17979 ( .C1(n14432), .C2(n16414), .A(n14431), .B(n14430), .ZN(
        n14433) );
  AOI21_X1 U17980 ( .B1(n10939), .B2(n14434), .A(n14433), .ZN(n14435) );
  NOR2_X1 U17981 ( .A1(n14462), .A2(n13256), .ZN(n14439) );
  NAND2_X1 U17982 ( .A1(n19326), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14448) );
  NAND2_X1 U17983 ( .A1(n19473), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14436) );
  OAI211_X1 U17984 ( .C1(n14437), .C2(n19471), .A(n14448), .B(n14436), .ZN(
        n14438) );
  OAI21_X1 U17985 ( .B1(n14461), .B2(n16514), .A(n14440), .ZN(P2_U2983) );
  AOI22_X1 U17986 ( .A1(n14442), .A2(P2_EAX_REG_31__SCAN_IN), .B1(n11215), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14443) );
  OAI21_X1 U17987 ( .B1(n14444), .B2(n16414), .A(n14443), .ZN(n14445) );
  INV_X1 U17988 ( .A(n14445), .ZN(n14446) );
  INV_X1 U17989 ( .A(n15952), .ZN(n19485) );
  OAI21_X1 U17990 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n19485), .A(
        n14447), .ZN(n14450) );
  INV_X1 U17991 ( .A(n14448), .ZN(n14449) );
  AOI21_X1 U17992 ( .B1(n14453), .B2(n16621), .A(n14452), .ZN(n14454) );
  OAI21_X1 U17993 ( .B1(n14462), .B2(n19491), .A(n14454), .ZN(n14455) );
  INV_X1 U17994 ( .A(n14455), .ZN(n14460) );
  NAND2_X1 U17995 ( .A1(n14458), .A2(n16624), .ZN(n14459) );
  OAI21_X1 U17996 ( .B1(n14461), .B2(n19500), .A(n10161), .ZN(P2_U3015) );
  NAND2_X1 U17997 ( .A1(n9726), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14463) );
  OAI21_X1 U17998 ( .B1(n14462), .B2(n9726), .A(n14463), .ZN(P2_U2856) );
  AOI22_X1 U17999 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14467) );
  AOI22_X1 U18000 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14466) );
  AOI22_X1 U18001 ( .A1(n10477), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14465) );
  AOI22_X1 U18002 ( .A1(n10528), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10563), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14464) );
  NAND4_X1 U18003 ( .A1(n14467), .A2(n14466), .A3(n14465), .A4(n14464), .ZN(
        n14473) );
  AOI22_X1 U18004 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14471) );
  AOI22_X1 U18005 ( .A1(n13847), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14470) );
  AOI22_X1 U18006 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14469) );
  AOI22_X1 U18007 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14508), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14468) );
  NAND4_X1 U18008 ( .A1(n14471), .A2(n14470), .A3(n14469), .A4(n14468), .ZN(
        n14472) );
  OR2_X1 U18009 ( .A1(n14473), .A2(n14472), .ZN(n15530) );
  AOI22_X1 U18010 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14503), .B1(
        n10437), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14477) );
  AOI22_X1 U18011 ( .A1(n10438), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14476) );
  AOI22_X1 U18012 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n10432), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14475) );
  AOI22_X1 U18013 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10563), .B1(
        n10528), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14474) );
  NAND4_X1 U18014 ( .A1(n14477), .A2(n14476), .A3(n14475), .A4(n14474), .ZN(
        n14483) );
  AOI22_X1 U18015 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n10456), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14481) );
  AOI22_X1 U18016 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14480) );
  AOI22_X1 U18017 ( .A1(n10472), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14479) );
  AOI22_X1 U18018 ( .A1(n10444), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__6__SCAN_IN), .B2(n14508), .ZN(n14478) );
  NAND4_X1 U18019 ( .A1(n14481), .A2(n14480), .A3(n14479), .A4(n14478), .ZN(
        n14482) );
  NOR2_X1 U18020 ( .A1(n14483), .A2(n14482), .ZN(n15526) );
  INV_X1 U18021 ( .A(n14686), .ZN(n14660) );
  INV_X1 U18022 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14485) );
  INV_X1 U18023 ( .A(n14685), .ZN(n14658) );
  INV_X1 U18024 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14484) );
  OAI22_X1 U18025 ( .A1(n14660), .A2(n14485), .B1(n14658), .B2(n14484), .ZN(
        n14489) );
  INV_X1 U18026 ( .A(n14684), .ZN(n14664) );
  INV_X1 U18027 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14487) );
  INV_X1 U18028 ( .A(n10240), .ZN(n14662) );
  INV_X1 U18029 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14486) );
  OAI22_X1 U18030 ( .A1(n14664), .A2(n14487), .B1(n14662), .B2(n14486), .ZN(
        n14488) );
  NOR2_X1 U18031 ( .A1(n14489), .A2(n14488), .ZN(n14492) );
  AOI22_X1 U18032 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14490) );
  XNOR2_X1 U18033 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14678) );
  NAND4_X1 U18034 ( .A1(n14492), .A2(n14491), .A3(n14490), .A4(n14678), .ZN(
        n14502) );
  INV_X1 U18035 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14493) );
  INV_X1 U18036 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n20807) );
  OAI22_X1 U18037 ( .A1(n14660), .A2(n14493), .B1(n14658), .B2(n20807), .ZN(
        n14497) );
  INV_X1 U18038 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14495) );
  INV_X1 U18039 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14494) );
  OAI22_X1 U18040 ( .A1(n14664), .A2(n14495), .B1(n14662), .B2(n14494), .ZN(
        n14496) );
  NOR2_X1 U18041 ( .A1(n14497), .A2(n14496), .ZN(n14500) );
  INV_X1 U18042 ( .A(n14678), .ZN(n14687) );
  AOI22_X1 U18043 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14498) );
  NAND4_X1 U18044 ( .A1(n14500), .A2(n14687), .A3(n14499), .A4(n14498), .ZN(
        n14501) );
  AND2_X1 U18045 ( .A1(n14502), .A2(n14501), .ZN(n14543) );
  NAND2_X1 U18046 ( .A1(n19514), .A2(n14543), .ZN(n14515) );
  AOI22_X1 U18047 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10437), .B1(
        n10438), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14507) );
  AOI22_X1 U18048 ( .A1(n14503), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10439), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14506) );
  AOI22_X1 U18049 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10528), .B1(
        n10477), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14505) );
  AOI22_X1 U18050 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10563), .B1(
        n10432), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14504) );
  NAND4_X1 U18051 ( .A1(n14507), .A2(n14506), .A3(n14505), .A4(n14504), .ZN(
        n14514) );
  AOI22_X1 U18052 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n10444), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14512) );
  AOI22_X1 U18053 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n13847), .B1(
        n13848), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14511) );
  AOI22_X1 U18054 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n10472), .B1(
        n10455), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U18055 ( .A1(n10456), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n14508), .ZN(n14509) );
  NAND4_X1 U18056 ( .A1(n14512), .A2(n14511), .A3(n14510), .A4(n14509), .ZN(
        n14513) );
  OR2_X1 U18057 ( .A1(n14514), .A2(n14513), .ZN(n14540) );
  XNOR2_X1 U18058 ( .A(n14515), .B(n14540), .ZN(n14546) );
  XNOR2_X1 U18059 ( .A(n14516), .B(n14546), .ZN(n15521) );
  NAND2_X1 U18060 ( .A1(n9740), .A2(n14543), .ZN(n15520) );
  NOR2_X1 U18061 ( .A1(n15521), .A2(n15520), .ZN(n15519) );
  INV_X1 U18062 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14518) );
  OAI22_X1 U18063 ( .A1(n14660), .A2(n14519), .B1(n14658), .B2(n14518), .ZN(
        n14523) );
  INV_X1 U18064 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n14521) );
  INV_X1 U18065 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14520) );
  OAI22_X1 U18066 ( .A1(n14664), .A2(n14521), .B1(n14662), .B2(n14520), .ZN(
        n14522) );
  NOR2_X1 U18067 ( .A1(n14523), .A2(n14522), .ZN(n14527) );
  AOI22_X1 U18068 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9736), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14526) );
  AOI22_X1 U18069 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14525) );
  NAND4_X1 U18070 ( .A1(n14527), .A2(n14526), .A3(n14525), .A4(n14678), .ZN(
        n14539) );
  INV_X1 U18071 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14529) );
  INV_X1 U18072 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14528) );
  OAI22_X1 U18073 ( .A1(n14660), .A2(n14529), .B1(n14658), .B2(n14528), .ZN(
        n14533) );
  INV_X1 U18074 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14530) );
  OAI22_X1 U18075 ( .A1(n14664), .A2(n14531), .B1(n14662), .B2(n14530), .ZN(
        n14532) );
  NOR2_X1 U18076 ( .A1(n14533), .A2(n14532), .ZN(n14537) );
  AOI22_X1 U18077 ( .A1(n9738), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14524), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14536) );
  AOI22_X1 U18078 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14535) );
  NAND4_X1 U18079 ( .A1(n14537), .A2(n14687), .A3(n14536), .A4(n14535), .ZN(
        n14538) );
  NAND2_X1 U18080 ( .A1(n14539), .A2(n14538), .ZN(n14548) );
  NAND2_X1 U18081 ( .A1(n14540), .A2(n14543), .ZN(n14549) );
  XOR2_X1 U18082 ( .A(n14548), .B(n14549), .Z(n14541) );
  NAND2_X1 U18083 ( .A1(n14541), .A2(n14570), .ZN(n15509) );
  INV_X1 U18084 ( .A(n14548), .ZN(n14542) );
  NAND2_X1 U18085 ( .A1(n9739), .A2(n14542), .ZN(n15512) );
  INV_X1 U18086 ( .A(n14543), .ZN(n14544) );
  NOR2_X1 U18087 ( .A1(n15512), .A2(n14544), .ZN(n14545) );
  NOR2_X1 U18088 ( .A1(n14549), .A2(n14548), .ZN(n14571) );
  INV_X1 U18089 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14551) );
  INV_X1 U18090 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14550) );
  OAI22_X1 U18091 ( .A1(n14660), .A2(n14551), .B1(n14658), .B2(n14550), .ZN(
        n14555) );
  INV_X1 U18092 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14552) );
  OAI22_X1 U18093 ( .A1(n14664), .A2(n14553), .B1(n14662), .B2(n14552), .ZN(
        n14554) );
  NOR2_X1 U18094 ( .A1(n14555), .A2(n14554), .ZN(n14558) );
  AOI22_X1 U18095 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14556) );
  NAND4_X1 U18096 ( .A1(n14558), .A2(n14557), .A3(n14556), .A4(n14678), .ZN(
        n14569) );
  INV_X1 U18097 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14560) );
  INV_X1 U18098 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14559) );
  OAI22_X1 U18099 ( .A1(n14660), .A2(n14560), .B1(n14658), .B2(n14559), .ZN(
        n14564) );
  INV_X1 U18100 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14562) );
  INV_X1 U18101 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14561) );
  OAI22_X1 U18102 ( .A1(n14664), .A2(n14562), .B1(n14662), .B2(n14561), .ZN(
        n14563) );
  NOR2_X1 U18103 ( .A1(n14564), .A2(n14563), .ZN(n14567) );
  AOI22_X1 U18104 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14565) );
  NAND4_X1 U18105 ( .A1(n14567), .A2(n14687), .A3(n14566), .A4(n14565), .ZN(
        n14568) );
  AND2_X1 U18106 ( .A1(n14569), .A2(n14568), .ZN(n14573) );
  NAND2_X1 U18107 ( .A1(n14571), .A2(n14573), .ZN(n14598) );
  OAI211_X1 U18108 ( .C1(n14571), .C2(n14573), .A(n14570), .B(n14598), .ZN(
        n14576) );
  INV_X1 U18109 ( .A(n14576), .ZN(n14572) );
  XNOR2_X1 U18110 ( .A(n14575), .B(n14572), .ZN(n15505) );
  INV_X1 U18111 ( .A(n14573), .ZN(n14574) );
  NOR2_X1 U18112 ( .A1(n19514), .A2(n14574), .ZN(n15504) );
  NAND2_X1 U18113 ( .A1(n15505), .A2(n15504), .ZN(n15503) );
  INV_X1 U18114 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14578) );
  OAI22_X1 U18115 ( .A1(n14660), .A2(n14579), .B1(n14658), .B2(n14578), .ZN(
        n14583) );
  OAI22_X1 U18116 ( .A1(n14664), .A2(n14581), .B1(n14662), .B2(n14580), .ZN(
        n14582) );
  NOR2_X1 U18117 ( .A1(n14583), .A2(n14582), .ZN(n14586) );
  AOI22_X1 U18118 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14584) );
  NAND4_X1 U18119 ( .A1(n14586), .A2(n14585), .A3(n14584), .A4(n14678), .ZN(
        n14597) );
  OAI22_X1 U18120 ( .A1(n14660), .A2(n14588), .B1(n14658), .B2(n14587), .ZN(
        n14592) );
  INV_X1 U18121 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14590) );
  OAI22_X1 U18122 ( .A1(n14664), .A2(n14590), .B1(n14662), .B2(n14589), .ZN(
        n14591) );
  NOR2_X1 U18123 ( .A1(n14592), .A2(n14591), .ZN(n14595) );
  AOI22_X1 U18124 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14593) );
  NAND4_X1 U18125 ( .A1(n14595), .A2(n14687), .A3(n14594), .A4(n14593), .ZN(
        n14596) );
  NAND2_X1 U18126 ( .A1(n14597), .A2(n14596), .ZN(n14600) );
  AOI21_X1 U18127 ( .B1(n14598), .B2(n14600), .A(n14623), .ZN(n14599) );
  OR2_X1 U18128 ( .A1(n14598), .A2(n14600), .ZN(n14624) );
  NAND2_X1 U18129 ( .A1(n14599), .A2(n14624), .ZN(n14602) );
  NOR2_X1 U18130 ( .A1(n19514), .A2(n14600), .ZN(n15497) );
  INV_X1 U18131 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14604) );
  INV_X1 U18132 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14603) );
  OAI22_X1 U18133 ( .A1(n14660), .A2(n14604), .B1(n14658), .B2(n14603), .ZN(
        n14608) );
  INV_X1 U18134 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14605) );
  OAI22_X1 U18135 ( .A1(n14664), .A2(n14606), .B1(n14662), .B2(n14605), .ZN(
        n14607) );
  NOR2_X1 U18136 ( .A1(n14608), .A2(n14607), .ZN(n14611) );
  AOI22_X1 U18137 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14609) );
  NAND4_X1 U18138 ( .A1(n14611), .A2(n14610), .A3(n14609), .A4(n14678), .ZN(
        n14622) );
  INV_X1 U18139 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14613) );
  INV_X1 U18140 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14612) );
  OAI22_X1 U18141 ( .A1(n14660), .A2(n14613), .B1(n14658), .B2(n14612), .ZN(
        n14617) );
  INV_X1 U18142 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14615) );
  INV_X1 U18143 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14614) );
  OAI22_X1 U18144 ( .A1(n14664), .A2(n14615), .B1(n14662), .B2(n14614), .ZN(
        n14616) );
  NOR2_X1 U18145 ( .A1(n14617), .A2(n14616), .ZN(n14620) );
  AOI22_X1 U18146 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14618) );
  NAND4_X1 U18147 ( .A1(n14620), .A2(n14687), .A3(n14619), .A4(n14618), .ZN(
        n14621) );
  NAND2_X1 U18148 ( .A1(n14622), .A2(n14621), .ZN(n14626) );
  NOR2_X1 U18149 ( .A1(n14624), .A2(n14626), .ZN(n15484) );
  AOI211_X1 U18150 ( .C1(n14626), .C2(n14624), .A(n14623), .B(n15484), .ZN(
        n14625) );
  INV_X1 U18151 ( .A(n14626), .ZN(n14627) );
  NAND2_X1 U18152 ( .A1(n9739), .A2(n14627), .ZN(n15492) );
  INV_X1 U18153 ( .A(n14628), .ZN(n15485) );
  INV_X1 U18154 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14629) );
  OAI22_X1 U18155 ( .A1(n14660), .A2(n14630), .B1(n14658), .B2(n14629), .ZN(
        n14634) );
  OAI22_X1 U18156 ( .A1(n14664), .A2(n14632), .B1(n14662), .B2(n14631), .ZN(
        n14633) );
  NOR2_X1 U18157 ( .A1(n14634), .A2(n14633), .ZN(n14637) );
  AOI22_X1 U18158 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14635) );
  NAND4_X1 U18159 ( .A1(n14637), .A2(n14636), .A3(n14635), .A4(n14678), .ZN(
        n14648) );
  INV_X1 U18160 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14638) );
  OAI22_X1 U18161 ( .A1(n14660), .A2(n14639), .B1(n14658), .B2(n14638), .ZN(
        n14643) );
  INV_X1 U18162 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14641) );
  OAI22_X1 U18163 ( .A1(n14664), .A2(n14641), .B1(n14662), .B2(n14640), .ZN(
        n14642) );
  NOR2_X1 U18164 ( .A1(n14643), .A2(n14642), .ZN(n14646) );
  AOI22_X1 U18165 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14644) );
  NAND4_X1 U18166 ( .A1(n14646), .A2(n14687), .A3(n14645), .A4(n14644), .ZN(
        n14647) );
  AND2_X1 U18167 ( .A1(n14648), .A2(n14647), .ZN(n15487) );
  OAI21_X2 U18168 ( .B1(n15491), .B2(n15485), .A(n15487), .ZN(n15481) );
  AND2_X1 U18169 ( .A1(n19514), .A2(n15487), .ZN(n14649) );
  AND2_X1 U18170 ( .A1(n15484), .A2(n14649), .ZN(n14673) );
  INV_X1 U18171 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n20844) );
  OAI22_X1 U18172 ( .A1(n10595), .A2(n14660), .B1(n14658), .B2(n20844), .ZN(
        n14653) );
  INV_X1 U18173 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n14651) );
  OAI22_X1 U18174 ( .A1(n14664), .A2(n14651), .B1(n14662), .B2(n14650), .ZN(
        n14652) );
  NOR2_X1 U18175 ( .A1(n14653), .A2(n14652), .ZN(n14656) );
  AOI22_X1 U18176 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14654) );
  NAND4_X1 U18177 ( .A1(n14656), .A2(n14655), .A3(n14654), .A4(n14678), .ZN(
        n14671) );
  INV_X1 U18178 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14657) );
  OAI22_X1 U18179 ( .A1(n14660), .A2(n14659), .B1(n14658), .B2(n14657), .ZN(
        n14666) );
  INV_X1 U18180 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14663) );
  OAI22_X1 U18181 ( .A1(n14664), .A2(n14663), .B1(n14662), .B2(n14661), .ZN(
        n14665) );
  NOR2_X1 U18182 ( .A1(n14666), .A2(n14665), .ZN(n14669) );
  AOI22_X1 U18183 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14667) );
  NAND4_X1 U18184 ( .A1(n14669), .A2(n14687), .A3(n14668), .A4(n14667), .ZN(
        n14670) );
  AND2_X1 U18185 ( .A1(n14671), .A2(n14670), .ZN(n14672) );
  NAND2_X1 U18186 ( .A1(n14673), .A2(n14672), .ZN(n14674) );
  OAI21_X1 U18187 ( .B1(n14673), .B2(n14672), .A(n14674), .ZN(n15480) );
  INV_X1 U18188 ( .A(n14674), .ZN(n14675) );
  AOI22_X1 U18189 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14676) );
  NAND2_X1 U18190 ( .A1(n14677), .A2(n14676), .ZN(n14693) );
  AOI22_X1 U18191 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14680) );
  AOI22_X1 U18192 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14679) );
  NAND3_X1 U18193 ( .A1(n14680), .A2(n14679), .A3(n14678), .ZN(n14692) );
  AOI22_X1 U18194 ( .A1(n16033), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14682) );
  NAND2_X1 U18195 ( .A1(n14683), .A2(n14682), .ZN(n14691) );
  AOI22_X1 U18196 ( .A1(n10240), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14684), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14689) );
  AOI22_X1 U18197 ( .A1(n14686), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14685), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14688) );
  NAND3_X1 U18198 ( .A1(n14689), .A2(n14688), .A3(n14687), .ZN(n14690) );
  OAI22_X1 U18199 ( .A1(n14693), .A2(n14692), .B1(n14691), .B2(n14690), .ZN(
        n14694) );
  INV_X1 U18200 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14698) );
  OAI22_X1 U18201 ( .A1(n15577), .A2(n19363), .B1(n19387), .B2(n14695), .ZN(
        n14696) );
  AOI21_X1 U18202 ( .B1(n19356), .B2(BUF1_REG_30__SCAN_IN), .A(n14696), .ZN(
        n14697) );
  OAI21_X1 U18203 ( .B1(n15581), .B2(n14698), .A(n14697), .ZN(n14699) );
  AOI21_X1 U18204 ( .B1(n16423), .B2(n19416), .A(n14699), .ZN(n14700) );
  OAI21_X1 U18205 ( .B1(n14703), .B2(n19390), .A(n14700), .ZN(P2_U2889) );
  NOR2_X1 U18206 ( .A1(n16422), .A2(n9726), .ZN(n14701) );
  AOI21_X1 U18207 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n9726), .A(n14701), .ZN(
        n14702) );
  AOI22_X1 U18208 ( .A1(n14718), .A2(n14705), .B1(n14729), .B2(n14704), .ZN(
        n14707) );
  XNOR2_X1 U18209 ( .A(n14707), .B(n14706), .ZN(n15148) );
  AOI21_X2 U18210 ( .B1(n14710), .B2(n14708), .A(n14709), .ZN(n14997) );
  NAND2_X1 U18211 ( .A1(n14997), .A2(n20233), .ZN(n14717) );
  INV_X1 U18212 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20672) );
  INV_X1 U18213 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14993) );
  OAI21_X1 U18214 ( .B1(n14722), .B2(n20672), .A(n14993), .ZN(n14715) );
  INV_X1 U18215 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14902) );
  NOR2_X1 U18216 ( .A1(n16272), .A2(n14902), .ZN(n14713) );
  OAI22_X1 U18217 ( .A1(n14711), .A2(n20257), .B1(n20277), .B2(n14995), .ZN(
        n14712) );
  AOI211_X1 U18218 ( .C1(n14715), .C2(n14714), .A(n14713), .B(n14712), .ZN(
        n14716) );
  OAI211_X1 U18219 ( .C1(n20267), .C2(n15148), .A(n14717), .B(n14716), .ZN(
        P1_U2810) );
  OAI21_X1 U18220 ( .B1(n14729), .B2(n14719), .A(n14718), .ZN(n15162) );
  INV_X1 U18221 ( .A(n14947), .ZN(n15007) );
  NAND2_X1 U18222 ( .A1(n15007), .A2(n20233), .ZN(n14727) );
  INV_X1 U18223 ( .A(n14737), .ZN(n14725) );
  INV_X1 U18224 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14903) );
  AOI22_X1 U18225 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20269), .B1(
        n20221), .B2(n15003), .ZN(n14721) );
  OAI21_X1 U18226 ( .B1(n16272), .B2(n14903), .A(n14721), .ZN(n14724) );
  NOR2_X1 U18227 ( .A1(n14722), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14723) );
  AOI211_X1 U18228 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14725), .A(n14724), 
        .B(n14723), .ZN(n14726) );
  OAI211_X1 U18229 ( .C1(n20267), .C2(n15162), .A(n14727), .B(n14726), .ZN(
        P1_U2811) );
  INV_X1 U18230 ( .A(n14728), .ZN(n14951) );
  AOI21_X1 U18231 ( .B1(n14730), .B2(n14743), .A(n14729), .ZN(n15174) );
  OAI22_X1 U18232 ( .A1(n14732), .A2(n20257), .B1(n20277), .B2(n14731), .ZN(
        n14733) );
  AOI21_X1 U18233 ( .B1(n20263), .B2(P1_EBX_REG_28__SCAN_IN), .A(n14733), .ZN(
        n14735) );
  NAND3_X1 U18234 ( .A1(n14746), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14736), 
        .ZN(n14734) );
  OAI211_X1 U18235 ( .C1(n14737), .C2(n14736), .A(n14735), .B(n14734), .ZN(
        n14738) );
  AOI21_X1 U18236 ( .B1(n15174), .B2(n20253), .A(n14738), .ZN(n14739) );
  OAI21_X1 U18237 ( .B1(n14951), .B2(n20242), .A(n14739), .ZN(P1_U2812) );
  OAI21_X1 U18239 ( .B1(n14741), .B2(n14742), .A(n12130), .ZN(n15012) );
  INV_X1 U18240 ( .A(n14743), .ZN(n14744) );
  AOI21_X1 U18241 ( .B1(n14745), .B2(n14758), .A(n14744), .ZN(n15182) );
  INV_X1 U18242 ( .A(n14746), .ZN(n14752) );
  INV_X1 U18243 ( .A(n14747), .ZN(n15015) );
  OAI22_X1 U18244 ( .A1(n14748), .A2(n20257), .B1(n20277), .B2(n15015), .ZN(
        n14749) );
  AOI21_X1 U18245 ( .B1(n20263), .B2(P1_EBX_REG_27__SCAN_IN), .A(n14749), .ZN(
        n14751) );
  NAND2_X1 U18246 ( .A1(n14761), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14750) );
  OAI211_X1 U18247 ( .C1(n14752), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14751), 
        .B(n14750), .ZN(n14753) );
  AOI21_X1 U18248 ( .B1(n15182), .B2(n20253), .A(n14753), .ZN(n14754) );
  OAI21_X1 U18249 ( .B1(n15012), .B2(n20242), .A(n14754), .ZN(P1_U2813) );
  AOI21_X1 U18250 ( .B1(n14756), .B2(n14755), .A(n14741), .ZN(n15024) );
  INV_X1 U18251 ( .A(n15024), .ZN(n14956) );
  INV_X1 U18252 ( .A(n14758), .ZN(n14759) );
  AOI21_X1 U18253 ( .B1(n14760), .B2(n14757), .A(n14759), .ZN(n15194) );
  INV_X1 U18254 ( .A(n14761), .ZN(n14767) );
  INV_X1 U18255 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15020) );
  INV_X1 U18256 ( .A(n14788), .ZN(n14762) );
  NAND4_X1 U18257 ( .A1(n14762), .A2(P1_REIP_REG_24__SCAN_IN), .A3(
        P1_REIP_REG_25__SCAN_IN), .A4(n15020), .ZN(n14766) );
  OAI22_X1 U18258 ( .A1(n14763), .A2(n20257), .B1(n20277), .B2(n15022), .ZN(
        n14764) );
  AOI21_X1 U18259 ( .B1(n20263), .B2(P1_EBX_REG_26__SCAN_IN), .A(n14764), .ZN(
        n14765) );
  OAI211_X1 U18260 ( .C1(n14767), .C2(n15020), .A(n14766), .B(n14765), .ZN(
        n14768) );
  AOI21_X1 U18261 ( .B1(n15194), .B2(n20253), .A(n14768), .ZN(n14769) );
  OAI21_X1 U18262 ( .B1(n14956), .B2(n20242), .A(n14769), .ZN(P1_U2814) );
  OR2_X1 U18263 ( .A1(n14770), .A2(n14771), .ZN(n14772) );
  NAND2_X1 U18264 ( .A1(n14757), .A2(n14772), .ZN(n15198) );
  OAI21_X1 U18265 ( .B1(n14774), .B2(n14775), .A(n14755), .ZN(n14959) );
  INV_X1 U18266 ( .A(n14959), .ZN(n15035) );
  NAND2_X1 U18267 ( .A1(n15035), .A2(n20233), .ZN(n14781) );
  OAI21_X1 U18268 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n20271), .A(n14802), 
        .ZN(n14779) );
  AOI22_X1 U18269 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n20269), .B1(
        n20221), .B2(n15030), .ZN(n14776) );
  OAI21_X1 U18270 ( .B1(n16272), .B2(n14907), .A(n14776), .ZN(n14778) );
  INV_X1 U18271 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20663) );
  NOR3_X1 U18272 ( .A1(n14788), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n20663), 
        .ZN(n14777) );
  AOI211_X1 U18273 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14779), .A(n14778), 
        .B(n14777), .ZN(n14780) );
  OAI211_X1 U18274 ( .C1(n20267), .C2(n15198), .A(n14781), .B(n14780), .ZN(
        P1_U2815) );
  AOI21_X1 U18275 ( .B1(n14783), .B2(n14782), .A(n14774), .ZN(n15043) );
  INV_X1 U18276 ( .A(n15043), .ZN(n14963) );
  INV_X1 U18277 ( .A(n14784), .ZN(n14786) );
  INV_X1 U18278 ( .A(n14795), .ZN(n14785) );
  AOI21_X1 U18279 ( .B1(n14786), .B2(n14785), .A(n14770), .ZN(n15215) );
  OAI22_X1 U18280 ( .A1(n14787), .A2(n20257), .B1(n20277), .B2(n15041), .ZN(
        n14790) );
  NOR2_X1 U18281 ( .A1(n14788), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14789) );
  AOI211_X1 U18282 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n20263), .A(n14790), .B(
        n14789), .ZN(n14791) );
  OAI21_X1 U18283 ( .B1(n20663), .B2(n14802), .A(n14791), .ZN(n14792) );
  AOI21_X1 U18284 ( .B1(n15215), .B2(n20253), .A(n14792), .ZN(n14793) );
  OAI21_X1 U18285 ( .B1(n14963), .B2(n20242), .A(n14793), .ZN(P1_U2816) );
  AND2_X1 U18286 ( .A1(n14810), .A2(n14794), .ZN(n14796) );
  OR2_X1 U18287 ( .A1(n14796), .A2(n14795), .ZN(n15224) );
  OAI21_X1 U18288 ( .B1(n14797), .B2(n14798), .A(n14782), .ZN(n14967) );
  INV_X1 U18289 ( .A(n14967), .ZN(n15051) );
  NAND2_X1 U18290 ( .A1(n15051), .A2(n20233), .ZN(n14807) );
  INV_X1 U18291 ( .A(n14799), .ZN(n15049) );
  OAI22_X1 U18292 ( .A1(n14800), .A2(n20257), .B1(n20277), .B2(n15049), .ZN(
        n14805) );
  AOI21_X1 U18293 ( .B1(n16219), .B2(n14801), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n14803) );
  NOR2_X1 U18294 ( .A1(n14803), .A2(n14802), .ZN(n14804) );
  AOI211_X1 U18295 ( .C1(P1_EBX_REG_23__SCAN_IN), .C2(n20263), .A(n14805), .B(
        n14804), .ZN(n14806) );
  OAI211_X1 U18296 ( .C1(n20267), .C2(n15224), .A(n14807), .B(n14806), .ZN(
        P1_U2817) );
  AOI21_X1 U18297 ( .B1(n14809), .B2(n14808), .A(n14797), .ZN(n15059) );
  INV_X1 U18298 ( .A(n15059), .ZN(n14971) );
  INV_X1 U18299 ( .A(n14810), .ZN(n14811) );
  AOI21_X1 U18300 ( .B1(n14812), .B2(n14828), .A(n14811), .ZN(n15241) );
  INV_X1 U18301 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15066) );
  NAND2_X1 U18302 ( .A1(n14813), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n14831) );
  OAI21_X1 U18303 ( .B1(n14892), .B2(n14831), .A(n14847), .ZN(n16226) );
  INV_X1 U18304 ( .A(n16226), .ZN(n14814) );
  AOI21_X1 U18305 ( .B1(n16239), .B2(n15066), .A(n14814), .ZN(n14821) );
  OAI22_X1 U18306 ( .A1(n14815), .A2(n20257), .B1(n20277), .B2(n15057), .ZN(
        n14819) );
  INV_X1 U18307 ( .A(n16219), .ZN(n14817) );
  NOR3_X1 U18308 ( .A1(n14817), .A2(P1_REIP_REG_22__SCAN_IN), .A3(n14816), 
        .ZN(n14818) );
  AOI211_X1 U18309 ( .C1(P1_EBX_REG_22__SCAN_IN), .C2(n20263), .A(n14819), .B(
        n14818), .ZN(n14820) );
  OAI21_X1 U18310 ( .B1(n14821), .B2(n20661), .A(n14820), .ZN(n14822) );
  AOI21_X1 U18311 ( .B1(n15241), .B2(n20253), .A(n14822), .ZN(n14823) );
  OAI21_X1 U18312 ( .B1(n14971), .B2(n20242), .A(n14823), .ZN(P1_U2818) );
  OAI21_X1 U18313 ( .B1(n14915), .B2(n14826), .A(n14808), .ZN(n15065) );
  INV_X1 U18314 ( .A(n14828), .ZN(n14829) );
  AOI21_X1 U18315 ( .B1(n14830), .B2(n14827), .A(n14829), .ZN(n15249) );
  NOR2_X1 U18316 ( .A1(n16226), .A2(n15066), .ZN(n14837) );
  INV_X1 U18317 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14835) );
  OR3_X1 U18318 ( .A1(n20271), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14831), .ZN(
        n14834) );
  INV_X1 U18319 ( .A(n15068), .ZN(n14832) );
  AOI22_X1 U18320 ( .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n20269), .B1(
        n20221), .B2(n14832), .ZN(n14833) );
  OAI211_X1 U18321 ( .C1(n16272), .C2(n14835), .A(n14834), .B(n14833), .ZN(
        n14836) );
  AOI211_X1 U18322 ( .C1(n15249), .C2(n20253), .A(n14837), .B(n14836), .ZN(
        n14838) );
  OAI21_X1 U18323 ( .B1(n15065), .B2(n20242), .A(n14838), .ZN(P1_U2819) );
  INV_X1 U18324 ( .A(n14839), .ZN(n14840) );
  AND2_X1 U18325 ( .A1(n14926), .A2(n14842), .ZN(n14843) );
  OR2_X1 U18326 ( .A1(n14913), .A2(n14843), .ZN(n15268) );
  INV_X1 U18327 ( .A(n15268), .ZN(n14919) );
  INV_X1 U18328 ( .A(n16227), .ZN(n14844) );
  NAND2_X1 U18329 ( .A1(n14845), .A2(n14844), .ZN(n14846) );
  NAND2_X1 U18330 ( .A1(n14847), .A2(n14846), .ZN(n16230) );
  INV_X1 U18331 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20657) );
  NOR2_X1 U18332 ( .A1(n16230), .A2(n20657), .ZN(n14855) );
  INV_X1 U18333 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14853) );
  INV_X1 U18334 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20654) );
  AOI211_X1 U18335 ( .C1(n20657), .C2(n20654), .A(n16227), .B(n20271), .ZN(
        n14850) );
  OAI21_X1 U18336 ( .B1(n20257), .B2(n15083), .A(n20254), .ZN(n14848) );
  AOI21_X1 U18337 ( .B1(n14850), .B2(n14849), .A(n14848), .ZN(n14852) );
  NAND2_X1 U18338 ( .A1(n20221), .A2(n15085), .ZN(n14851) );
  OAI211_X1 U18339 ( .C1(n16272), .C2(n14853), .A(n14852), .B(n14851), .ZN(
        n14854) );
  AOI211_X1 U18340 ( .C1(n14919), .C2(n20253), .A(n14855), .B(n14854), .ZN(
        n14856) );
  OAI21_X1 U18341 ( .B1(n15088), .B2(n20242), .A(n14856), .ZN(P1_U2821) );
  AOI21_X1 U18342 ( .B1(n16239), .B2(n14857), .A(P1_REIP_REG_17__SCAN_IN), 
        .ZN(n14872) );
  NOR2_X1 U18343 ( .A1(n14858), .A2(n14859), .ZN(n14860) );
  OR2_X1 U18344 ( .A1(n14824), .A2(n14860), .ZN(n15107) );
  INV_X1 U18345 ( .A(n15107), .ZN(n14861) );
  NAND2_X1 U18346 ( .A1(n14861), .A2(n20233), .ZN(n14871) );
  OR2_X1 U18347 ( .A1(n14863), .A2(n14864), .ZN(n14865) );
  AND2_X1 U18348 ( .A1(n14862), .A2(n14865), .ZN(n16328) );
  INV_X1 U18349 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14868) );
  AOI21_X1 U18350 ( .B1(n20269), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n20349), .ZN(n14867) );
  NAND2_X1 U18351 ( .A1(n20221), .A2(n15104), .ZN(n14866) );
  OAI211_X1 U18352 ( .C1(n16272), .C2(n14868), .A(n14867), .B(n14866), .ZN(
        n14869) );
  AOI21_X1 U18353 ( .B1(n16328), .B2(n20253), .A(n14869), .ZN(n14870) );
  OAI211_X1 U18354 ( .C1(n14872), .C2(n16230), .A(n14871), .B(n14870), .ZN(
        P1_U2823) );
  OAI221_X1 U18355 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n20224), .C1(
        P1_REIP_REG_10__SCAN_IN), .C2(P1_REIP_REG_9__SCAN_IN), .A(n16276), 
        .ZN(n14878) );
  NOR2_X1 U18356 ( .A1(n20277), .A2(n15142), .ZN(n14873) );
  AOI211_X1 U18357 ( .C1(n20269), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20349), .B(n14873), .ZN(n14874) );
  OAI21_X1 U18358 ( .B1(n14875), .B2(n16272), .A(n14874), .ZN(n14876) );
  AOI21_X1 U18359 ( .B1(n20253), .B2(n16360), .A(n14876), .ZN(n14877) );
  OAI211_X1 U18360 ( .C1(n20242), .C2(n15146), .A(n14878), .B(n14877), .ZN(
        P1_U2830) );
  OAI22_X1 U18361 ( .A1(n14879), .A2(n20277), .B1(n20257), .B2(n20834), .ZN(
        n14882) );
  NOR2_X1 U18362 ( .A1(n16272), .A2(n14880), .ZN(n14881) );
  AOI211_X1 U18363 ( .C1(n20373), .C2(n20253), .A(n14882), .B(n14881), .ZN(
        n14883) );
  OAI21_X1 U18364 ( .B1(n14884), .B2(n20262), .A(n14883), .ZN(n14887) );
  NOR3_X1 U18365 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(n20271), .A3(n14885), .ZN(
        n14886) );
  AOI211_X1 U18366 ( .C1(n14888), .C2(n20272), .A(n14887), .B(n14886), .ZN(
        n14889) );
  OAI21_X1 U18367 ( .B1(n14891), .B2(n14890), .A(n14889), .ZN(P1_U2837) );
  INV_X1 U18368 ( .A(n20272), .ZN(n14898) );
  AOI22_X1 U18369 ( .A1(n16239), .A2(n13275), .B1(n20263), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n14897) );
  NOR2_X1 U18370 ( .A1(n20262), .A2(n12613), .ZN(n14895) );
  AOI22_X1 U18371 ( .A1(n20269), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14892), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14893) );
  OAI21_X1 U18372 ( .B1(n20277), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14893), .ZN(n14894) );
  AOI211_X1 U18373 ( .C1(n20253), .C2(n13167), .A(n14895), .B(n14894), .ZN(
        n14896) );
  OAI211_X1 U18374 ( .C1(n14899), .C2(n14898), .A(n14897), .B(n14896), .ZN(
        P1_U2839) );
  OAI22_X1 U18375 ( .A1(n14901), .A2(n14936), .B1(n14900), .B2(n20282), .ZN(
        P1_U2841) );
  INV_X1 U18376 ( .A(n14997), .ZN(n14944) );
  OAI222_X1 U18377 ( .A1(n14939), .A2(n14944), .B1(n20282), .B2(n14902), .C1(
        n15148), .C2(n14936), .ZN(P1_U2842) );
  OAI222_X1 U18378 ( .A1(n14903), .A2(n20282), .B1(n14936), .B2(n15162), .C1(
        n14947), .C2(n14939), .ZN(P1_U2843) );
  AOI22_X1 U18379 ( .A1(n15174), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_28__SCAN_IN), .ZN(n14904) );
  OAI21_X1 U18380 ( .B1(n14951), .B2(n14939), .A(n14904), .ZN(P1_U2844) );
  AOI22_X1 U18381 ( .A1(n15182), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14905) );
  OAI21_X1 U18382 ( .B1(n15012), .B2(n14939), .A(n14905), .ZN(P1_U2845) );
  AOI22_X1 U18383 ( .A1(n15194), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14906) );
  OAI21_X1 U18384 ( .B1(n14956), .B2(n14939), .A(n14906), .ZN(P1_U2846) );
  OAI222_X1 U18385 ( .A1(n14907), .A2(n20282), .B1(n14936), .B2(n15198), .C1(
        n14959), .C2(n14939), .ZN(P1_U2847) );
  AOI22_X1 U18386 ( .A1(n15215), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14908) );
  OAI21_X1 U18387 ( .B1(n14963), .B2(n14939), .A(n14908), .ZN(P1_U2848) );
  INV_X1 U18388 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14909) );
  OAI222_X1 U18389 ( .A1(n14909), .A2(n20282), .B1(n14936), .B2(n15224), .C1(
        n14967), .C2(n14939), .ZN(P1_U2849) );
  AOI22_X1 U18390 ( .A1(n15241), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_22__SCAN_IN), .ZN(n14910) );
  OAI21_X1 U18391 ( .B1(n14971), .B2(n14939), .A(n14910), .ZN(P1_U2850) );
  AOI22_X1 U18392 ( .A1(n15249), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14911) );
  OAI21_X1 U18393 ( .B1(n15065), .B2(n14939), .A(n14911), .ZN(P1_U2851) );
  INV_X1 U18394 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14918) );
  OR2_X1 U18395 ( .A1(n14913), .A2(n14912), .ZN(n14914) );
  NAND2_X1 U18396 ( .A1(n14827), .A2(n14914), .ZN(n16220) );
  INV_X1 U18397 ( .A(n16286), .ZN(n15079) );
  OAI222_X1 U18398 ( .A1(n14918), .A2(n20282), .B1(n14936), .B2(n16220), .C1(
        n15079), .C2(n14939), .ZN(P1_U2852) );
  AOI22_X1 U18399 ( .A1(n14919), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n14920) );
  OAI21_X1 U18400 ( .B1(n15088), .B2(n14939), .A(n14920), .ZN(P1_U2853) );
  OR2_X1 U18401 ( .A1(n14824), .A2(n14921), .ZN(n14922) );
  NAND2_X1 U18402 ( .A1(n14862), .A2(n14924), .ZN(n14925) );
  NAND2_X1 U18403 ( .A1(n14926), .A2(n14925), .ZN(n16236) );
  OAI22_X1 U18404 ( .A1(n16236), .A2(n14936), .B1(n14927), .B2(n20282), .ZN(
        n14928) );
  INV_X1 U18405 ( .A(n14928), .ZN(n14929) );
  OAI21_X1 U18406 ( .B1(n14981), .B2(n14939), .A(n14929), .ZN(P1_U2854) );
  AOI22_X1 U18407 ( .A1(n16328), .A2(n20706), .B1(n20707), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n14930) );
  OAI21_X1 U18408 ( .B1(n15107), .B2(n14939), .A(n14930), .ZN(P1_U2855) );
  AND2_X1 U18409 ( .A1(n14271), .A2(n14931), .ZN(n14932) );
  OR2_X1 U18410 ( .A1(n14932), .A2(n14858), .ZN(n16242) );
  NOR2_X1 U18411 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  OR2_X1 U18412 ( .A1(n14863), .A2(n14935), .ZN(n16244) );
  OAI22_X1 U18413 ( .A1(n16244), .A2(n14936), .B1(n16240), .B2(n20282), .ZN(
        n14937) );
  INV_X1 U18414 ( .A(n14937), .ZN(n14938) );
  OAI21_X1 U18415 ( .B1(n16242), .B2(n14939), .A(n14938), .ZN(P1_U2856) );
  AOI22_X1 U18416 ( .A1(n16284), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n16280), .ZN(n14943) );
  NOR3_X1 U18417 ( .A1(n16280), .A2(n14940), .A3(n11352), .ZN(n14941) );
  AOI22_X1 U18418 ( .A1(n16282), .A2(n20332), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n14985), .ZN(n14942) );
  OAI211_X1 U18419 ( .C1(n14944), .C2(n16283), .A(n14943), .B(n14942), .ZN(
        P1_U2874) );
  AOI22_X1 U18420 ( .A1(n16284), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n16280), .ZN(n14946) );
  AOI22_X1 U18421 ( .A1(n16282), .A2(n20330), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n14985), .ZN(n14945) );
  OAI211_X1 U18422 ( .C1(n14947), .C2(n16283), .A(n14946), .B(n14945), .ZN(
        P1_U2875) );
  AOI22_X1 U18423 ( .A1(n16284), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n16280), .ZN(n14950) );
  AOI22_X1 U18424 ( .A1(n16282), .A2(n14948), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n14985), .ZN(n14949) );
  OAI211_X1 U18425 ( .C1(n14951), .C2(n16283), .A(n14950), .B(n14949), .ZN(
        P1_U2876) );
  AOI22_X1 U18426 ( .A1(n16284), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n16280), .ZN(n14953) );
  AOI22_X1 U18427 ( .A1(n16282), .A2(n20328), .B1(BUF1_REG_27__SCAN_IN), .B2(
        n14985), .ZN(n14952) );
  OAI211_X1 U18428 ( .C1(n15012), .C2(n16283), .A(n14953), .B(n14952), .ZN(
        P1_U2877) );
  AOI22_X1 U18429 ( .A1(n16284), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n16280), .ZN(n14955) );
  AOI22_X1 U18430 ( .A1(n16282), .A2(n20326), .B1(BUF1_REG_26__SCAN_IN), .B2(
        n14985), .ZN(n14954) );
  OAI211_X1 U18431 ( .C1(n14956), .C2(n16283), .A(n14955), .B(n14954), .ZN(
        P1_U2878) );
  AOI22_X1 U18432 ( .A1(n16284), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n16280), .ZN(n14958) );
  AOI22_X1 U18433 ( .A1(n16282), .A2(n20324), .B1(n14985), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14957) );
  OAI211_X1 U18434 ( .C1(n14959), .C2(n16283), .A(n14958), .B(n14957), .ZN(
        P1_U2879) );
  AOI22_X1 U18435 ( .A1(n16284), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n16280), .ZN(n14962) );
  AOI22_X1 U18436 ( .A1(n16282), .A2(n14960), .B1(n14985), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14961) );
  OAI211_X1 U18437 ( .C1(n14963), .C2(n16283), .A(n14962), .B(n14961), .ZN(
        P1_U2880) );
  AOI22_X1 U18438 ( .A1(n16284), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n16280), .ZN(n14966) );
  AOI22_X1 U18439 ( .A1(n16282), .A2(n14964), .B1(n14985), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14965) );
  OAI211_X1 U18440 ( .C1(n14967), .C2(n16283), .A(n14966), .B(n14965), .ZN(
        P1_U2881) );
  AOI22_X1 U18441 ( .A1(n16284), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n16280), .ZN(n14970) );
  AOI22_X1 U18442 ( .A1(n16282), .A2(n14968), .B1(n14985), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14969) );
  OAI211_X1 U18443 ( .C1(n14971), .C2(n16283), .A(n14970), .B(n14969), .ZN(
        P1_U2882) );
  AOI22_X1 U18444 ( .A1(n16284), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n16280), .ZN(n14974) );
  AOI22_X1 U18445 ( .A1(n16282), .A2(n14972), .B1(n14985), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14973) );
  OAI211_X1 U18446 ( .C1(n15065), .C2(n16283), .A(n14974), .B(n14973), .ZN(
        P1_U2883) );
  AOI22_X1 U18447 ( .A1(n16284), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n16280), .ZN(n14977) );
  AOI22_X1 U18448 ( .A1(n16282), .A2(n14975), .B1(n14985), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14976) );
  OAI211_X1 U18449 ( .C1(n15088), .C2(n16283), .A(n14977), .B(n14976), .ZN(
        P1_U2885) );
  AOI22_X1 U18450 ( .A1(n16284), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n16280), .ZN(n14980) );
  AOI22_X1 U18451 ( .A1(n16282), .A2(n14978), .B1(n14985), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n14979) );
  OAI211_X1 U18452 ( .C1(n14981), .C2(n16283), .A(n14980), .B(n14979), .ZN(
        P1_U2886) );
  AOI22_X1 U18453 ( .A1(n16282), .A2(n14982), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n16280), .ZN(n14984) );
  AOI22_X1 U18454 ( .A1(n16284), .A2(DATAI_17_), .B1(n14985), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14983) );
  OAI211_X1 U18455 ( .C1(n15107), .C2(n16283), .A(n14984), .B(n14983), .ZN(
        P1_U2887) );
  AOI22_X1 U18456 ( .A1(n16284), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n16280), .ZN(n14988) );
  AOI22_X1 U18457 ( .A1(n16282), .A2(n14986), .B1(n14985), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n14987) );
  OAI211_X1 U18458 ( .C1(n16242), .C2(n16283), .A(n14988), .B(n14987), .ZN(
        P1_U2888) );
  INV_X1 U18459 ( .A(n14990), .ZN(n14991) );
  NOR2_X1 U18460 ( .A1(n20254), .A2(n14993), .ZN(n15153) );
  AOI21_X1 U18461 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15153), .ZN(n14994) );
  OAI21_X1 U18462 ( .B1(n20361), .B2(n14995), .A(n14994), .ZN(n14996) );
  AOI21_X1 U18463 ( .B1(n14997), .B2(n14067), .A(n14996), .ZN(n14998) );
  OAI21_X1 U18464 ( .B1(n15156), .B2(n20203), .A(n14998), .ZN(P1_U2969) );
  NAND2_X1 U18465 ( .A1(n15001), .A2(n15000), .ZN(n15002) );
  XNOR2_X1 U18466 ( .A(n14999), .B(n15002), .ZN(n15168) );
  INV_X1 U18467 ( .A(n15003), .ZN(n15005) );
  NOR2_X1 U18468 ( .A1(n20254), .A2(n20672), .ZN(n15164) );
  AOI21_X1 U18469 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15164), .ZN(n15004) );
  OAI21_X1 U18470 ( .B1(n20361), .B2(n15005), .A(n15004), .ZN(n15006) );
  OAI21_X1 U18471 ( .B1(n20203), .B2(n15168), .A(n15008), .ZN(P1_U2970) );
  OAI21_X1 U18472 ( .B1(n15097), .B2(n15010), .A(n15009), .ZN(n15019) );
  INV_X1 U18473 ( .A(n15012), .ZN(n15017) );
  INV_X1 U18474 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15013) );
  NOR2_X1 U18475 ( .A1(n20254), .A2(n15013), .ZN(n15180) );
  AOI21_X1 U18476 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15180), .ZN(n15014) );
  OAI21_X1 U18477 ( .B1(n20361), .B2(n15015), .A(n15014), .ZN(n15016) );
  AOI21_X1 U18478 ( .B1(n15017), .B2(n14067), .A(n15016), .ZN(n15018) );
  OAI21_X1 U18479 ( .B1(n20203), .B2(n15185), .A(n15018), .ZN(P1_U2972) );
  XOR2_X1 U18480 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15019), .Z(
        n15197) );
  NOR2_X1 U18481 ( .A1(n20254), .A2(n15020), .ZN(n15192) );
  AOI21_X1 U18482 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15192), .ZN(n15021) );
  OAI21_X1 U18483 ( .B1(n20361), .B2(n15022), .A(n15021), .ZN(n15023) );
  AOI21_X1 U18484 ( .B1(n15024), .B2(n14067), .A(n15023), .ZN(n15025) );
  OAI21_X1 U18485 ( .B1(n20203), .B2(n15197), .A(n15025), .ZN(P1_U2973) );
  NAND2_X1 U18486 ( .A1(n15026), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15037) );
  NAND2_X1 U18487 ( .A1(n11601), .A2(n15209), .ZN(n15027) );
  OAI21_X1 U18488 ( .B1(n11601), .B2(n20816), .A(n15027), .ZN(n15028) );
  AOI211_X1 U18489 ( .C1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C2(n15037), .A(
        n15028), .B(n9782), .ZN(n15029) );
  XNOR2_X1 U18490 ( .A(n15029), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15207) );
  INV_X1 U18491 ( .A(n15030), .ZN(n15033) );
  INV_X1 U18492 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15031) );
  NOR2_X1 U18493 ( .A1(n20254), .A2(n15031), .ZN(n15199) );
  AOI21_X1 U18494 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n15199), .ZN(n15032) );
  OAI21_X1 U18495 ( .B1(n20361), .B2(n15033), .A(n15032), .ZN(n15034) );
  AOI21_X1 U18496 ( .B1(n15035), .B2(n14067), .A(n15034), .ZN(n15036) );
  OAI21_X1 U18497 ( .B1(n15207), .B2(n20203), .A(n15036), .ZN(P1_U2974) );
  NAND2_X1 U18498 ( .A1(n15046), .A2(n15037), .ZN(n15038) );
  MUX2_X1 U18499 ( .A(n15038), .B(n15037), .S(n11601), .Z(n15039) );
  XNOR2_X1 U18500 ( .A(n15039), .B(n15209), .ZN(n15218) );
  NOR2_X1 U18501 ( .A1(n20254), .A2(n20663), .ZN(n15213) );
  AOI21_X1 U18502 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15213), .ZN(n15040) );
  OAI21_X1 U18503 ( .B1(n20361), .B2(n15041), .A(n15040), .ZN(n15042) );
  AOI21_X1 U18504 ( .B1(n15043), .B2(n14067), .A(n15042), .ZN(n15044) );
  OAI21_X1 U18505 ( .B1(n20203), .B2(n15218), .A(n15044), .ZN(P1_U2975) );
  XNOR2_X1 U18506 ( .A(n11601), .B(n20816), .ZN(n15045) );
  XNOR2_X1 U18507 ( .A(n15046), .B(n15045), .ZN(n15227) );
  INV_X1 U18508 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n15047) );
  NOR2_X1 U18509 ( .A1(n20254), .A2(n15047), .ZN(n15219) );
  AOI21_X1 U18510 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15219), .ZN(n15048) );
  OAI21_X1 U18511 ( .B1(n20361), .B2(n15049), .A(n15048), .ZN(n15050) );
  AOI21_X1 U18512 ( .B1(n15051), .B2(n14067), .A(n15050), .ZN(n15052) );
  OAI21_X1 U18513 ( .B1(n15227), .B2(n20203), .A(n15052), .ZN(P1_U2976) );
  NAND2_X1 U18514 ( .A1(n15054), .A2(n15053), .ZN(n15055) );
  XNOR2_X1 U18515 ( .A(n15055), .B(n15237), .ZN(n15244) );
  NOR2_X1 U18516 ( .A1(n20254), .A2(n20661), .ZN(n15240) );
  AOI21_X1 U18517 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15240), .ZN(n15056) );
  OAI21_X1 U18518 ( .B1(n20361), .B2(n15057), .A(n15056), .ZN(n15058) );
  AOI21_X1 U18519 ( .B1(n15059), .B2(n14067), .A(n15058), .ZN(n15060) );
  OAI21_X1 U18520 ( .B1(n20203), .B2(n15244), .A(n15060), .ZN(P1_U2977) );
  INV_X1 U18521 ( .A(n15061), .ZN(n15062) );
  NAND3_X1 U18522 ( .A1(n15062), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n11601), .ZN(n15075) );
  INV_X1 U18523 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n20987) );
  AOI22_X1 U18524 ( .A1(n15075), .A2(n15063), .B1(n11601), .B2(n20987), .ZN(
        n15064) );
  XNOR2_X1 U18525 ( .A(n15064), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15252) );
  INV_X1 U18526 ( .A(n15065), .ZN(n15070) );
  NOR2_X1 U18527 ( .A1(n20254), .A2(n15066), .ZN(n15247) );
  AOI21_X1 U18528 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15247), .ZN(n15067) );
  OAI21_X1 U18529 ( .B1(n20361), .B2(n15068), .A(n15067), .ZN(n15069) );
  AOI21_X1 U18530 ( .B1(n15070), .B2(n14067), .A(n15069), .ZN(n15071) );
  OAI21_X1 U18531 ( .B1(n15252), .B2(n20203), .A(n15071), .ZN(P1_U2978) );
  INV_X1 U18532 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15072) );
  NOR2_X1 U18533 ( .A1(n20254), .A2(n15072), .ZN(n15256) );
  NOR2_X1 U18534 ( .A1(n15134), .A2(n15073), .ZN(n15074) );
  AOI211_X1 U18535 ( .C1(n16303), .C2(n16222), .A(n15256), .B(n15074), .ZN(
        n15078) );
  XNOR2_X1 U18536 ( .A(n15076), .B(n20987), .ZN(n15253) );
  NAND2_X1 U18537 ( .A1(n15253), .A2(n20356), .ZN(n15077) );
  OAI211_X1 U18538 ( .C1(n15079), .C2(n15147), .A(n15078), .B(n15077), .ZN(
        P1_U2979) );
  NAND2_X1 U18539 ( .A1(n15061), .A2(n15080), .ZN(n15081) );
  MUX2_X1 U18540 ( .A(n15061), .B(n15081), .S(n15097), .Z(n15082) );
  XNOR2_X1 U18541 ( .A(n15082), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15260) );
  NAND2_X1 U18542 ( .A1(n15260), .A2(n20356), .ZN(n15087) );
  NOR2_X1 U18543 ( .A1(n20254), .A2(n20657), .ZN(n15263) );
  NOR2_X1 U18544 ( .A1(n15134), .A2(n15083), .ZN(n15084) );
  AOI211_X1 U18545 ( .C1(n16303), .C2(n15085), .A(n15263), .B(n15084), .ZN(
        n15086) );
  OAI211_X1 U18546 ( .C1(n15147), .C2(n15088), .A(n15087), .B(n15086), .ZN(
        P1_U2980) );
  OAI21_X1 U18547 ( .B1(n10120), .B2(n15090), .A(n15061), .ZN(n15277) );
  NOR2_X1 U18548 ( .A1(n20254), .A2(n20654), .ZN(n15272) );
  AOI21_X1 U18549 ( .B1(n20350), .B2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15272), .ZN(n15091) );
  OAI21_X1 U18550 ( .B1(n20361), .B2(n15092), .A(n15091), .ZN(n15093) );
  AOI21_X1 U18551 ( .B1(n16233), .B2(n14067), .A(n15093), .ZN(n15094) );
  OAI21_X1 U18552 ( .B1(n20203), .B2(n15277), .A(n15094), .ZN(P1_U2981) );
  AOI21_X1 U18553 ( .B1(n15095), .B2(n15278), .A(n15096), .ZN(n15099) );
  NOR2_X1 U18554 ( .A1(n15099), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15098) );
  MUX2_X1 U18555 ( .A(n15099), .B(n15098), .S(n15097), .Z(n15100) );
  XNOR2_X1 U18556 ( .A(n15100), .B(n20797), .ZN(n16329) );
  NAND2_X1 U18557 ( .A1(n16329), .A2(n20356), .ZN(n15106) );
  INV_X1 U18558 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15101) );
  OAI22_X1 U18559 ( .A1(n15134), .A2(n15102), .B1(n20254), .B2(n15101), .ZN(
        n15103) );
  AOI21_X1 U18560 ( .B1(n16303), .B2(n15104), .A(n15103), .ZN(n15105) );
  OAI211_X1 U18561 ( .C1(n15147), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        P1_U2982) );
  NOR2_X1 U18562 ( .A1(n15095), .A2(n15108), .ZN(n15281) );
  NOR3_X1 U18563 ( .A1(n15281), .A2(n16296), .A3(n15109), .ZN(n15113) );
  INV_X1 U18564 ( .A(n15279), .ZN(n15110) );
  NOR2_X1 U18565 ( .A1(n15111), .A2(n15110), .ZN(n15112) );
  XNOR2_X1 U18566 ( .A(n15113), .B(n15112), .ZN(n16336) );
  NAND2_X1 U18567 ( .A1(n16336), .A2(n20356), .ZN(n15117) );
  INV_X1 U18568 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15114) );
  OAI22_X1 U18569 ( .A1(n15134), .A2(n16250), .B1(n20254), .B2(n15114), .ZN(
        n15115) );
  AOI21_X1 U18570 ( .B1(n16303), .B2(n16255), .A(n15115), .ZN(n15116) );
  OAI211_X1 U18571 ( .C1(n15147), .C2(n16252), .A(n15117), .B(n15116), .ZN(
        P1_U2984) );
  INV_X1 U18572 ( .A(n15095), .ZN(n16297) );
  INV_X1 U18573 ( .A(n15118), .ZN(n15119) );
  AOI21_X1 U18574 ( .B1(n16297), .B2(n15120), .A(n15119), .ZN(n15132) );
  AND2_X1 U18575 ( .A1(n15121), .A2(n15122), .ZN(n15131) );
  NAND2_X1 U18576 ( .A1(n15132), .A2(n15131), .ZN(n15130) );
  NAND2_X1 U18577 ( .A1(n15130), .A2(n15122), .ZN(n15123) );
  XOR2_X1 U18578 ( .A(n15124), .B(n15123), .Z(n15290) );
  NAND2_X1 U18579 ( .A1(n15290), .A2(n20356), .ZN(n15128) );
  NOR2_X1 U18580 ( .A1(n20254), .A2(n20649), .ZN(n15296) );
  NOR2_X1 U18581 ( .A1(n20361), .A2(n15125), .ZN(n15126) );
  AOI211_X1 U18582 ( .C1(n20350), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15296), .B(n15126), .ZN(n15127) );
  OAI211_X1 U18583 ( .C1(n15147), .C2(n15129), .A(n15128), .B(n15127), .ZN(
        P1_U2986) );
  OAI21_X1 U18584 ( .B1(n15132), .B2(n15131), .A(n15130), .ZN(n15316) );
  NAND2_X1 U18585 ( .A1(n15316), .A2(n20356), .ZN(n15137) );
  INV_X1 U18586 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15133) );
  NOR2_X1 U18587 ( .A1(n20254), .A2(n15133), .ZN(n15310) );
  NOR2_X1 U18588 ( .A1(n15134), .A2(n20960), .ZN(n15135) );
  AOI211_X1 U18589 ( .C1(n16303), .C2(n16266), .A(n15310), .B(n15135), .ZN(
        n15136) );
  OAI211_X1 U18590 ( .C1(n15147), .C2(n15138), .A(n15137), .B(n15136), .ZN(
        P1_U2987) );
  MUX2_X1 U18591 ( .A(n15140), .B(n15095), .S(n11601), .Z(n15141) );
  XOR2_X1 U18592 ( .A(n13957), .B(n15141), .Z(n16361) );
  NAND2_X1 U18593 ( .A1(n16361), .A2(n20356), .ZN(n15145) );
  NOR2_X1 U18594 ( .A1(n20254), .A2(n20644), .ZN(n16359) );
  NOR2_X1 U18595 ( .A1(n20361), .A2(n15142), .ZN(n15143) );
  AOI211_X1 U18596 ( .C1(n20350), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16359), .B(n15143), .ZN(n15144) );
  OAI211_X1 U18597 ( .C1(n15147), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        P1_U2989) );
  INV_X1 U18598 ( .A(n15148), .ZN(n15154) );
  AOI21_X1 U18599 ( .B1(n15151), .B2(n15150), .A(n15149), .ZN(n15152) );
  AOI211_X1 U18600 ( .C1(n15154), .C2(n20374), .A(n15153), .B(n15152), .ZN(
        n15155) );
  OAI21_X1 U18601 ( .B1(n15156), .B2(n20385), .A(n15155), .ZN(P1_U3001) );
  INV_X1 U18602 ( .A(n15157), .ZN(n15178) );
  INV_X1 U18603 ( .A(n15171), .ZN(n15159) );
  OAI21_X1 U18604 ( .B1(n15178), .B2(n15159), .A(n15158), .ZN(n15166) );
  OAI21_X1 U18605 ( .B1(n15171), .B2(n15161), .A(n15160), .ZN(n15165) );
  NOR2_X1 U18606 ( .A1(n15162), .A2(n20392), .ZN(n15163) );
  AOI211_X1 U18607 ( .C1(n15166), .C2(n15165), .A(n15164), .B(n15163), .ZN(
        n15167) );
  OAI21_X1 U18608 ( .B1(n15168), .B2(n20385), .A(n15167), .ZN(P1_U3002) );
  INV_X1 U18609 ( .A(n15169), .ZN(n15170) );
  NOR3_X1 U18610 ( .A1(n15178), .A2(n15171), .A3(n15170), .ZN(n15172) );
  AOI211_X1 U18611 ( .C1(n15181), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n15173), .B(n15172), .ZN(n15176) );
  NAND2_X1 U18612 ( .A1(n15174), .A2(n20374), .ZN(n15175) );
  OAI211_X1 U18613 ( .C1(n15177), .C2(n20385), .A(n15176), .B(n15175), .ZN(
        P1_U3003) );
  NOR2_X1 U18614 ( .A1(n15178), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15179) );
  AOI211_X1 U18615 ( .C1(n15181), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15180), .B(n15179), .ZN(n15184) );
  NAND2_X1 U18616 ( .A1(n15182), .A2(n20374), .ZN(n15183) );
  OAI211_X1 U18617 ( .C1(n15185), .C2(n20385), .A(n15184), .B(n15183), .ZN(
        P1_U3004) );
  NOR2_X1 U18618 ( .A1(n15186), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15193) );
  INV_X1 U18619 ( .A(n15187), .ZN(n15203) );
  AND2_X1 U18620 ( .A1(n15188), .A2(n15202), .ZN(n15189) );
  NAND2_X1 U18621 ( .A1(n15220), .A2(n15189), .ZN(n15201) );
  AOI21_X1 U18622 ( .B1(n15203), .B2(n15201), .A(n15190), .ZN(n15191) );
  AOI211_X1 U18623 ( .C1(n15220), .C2(n15193), .A(n15192), .B(n15191), .ZN(
        n15196) );
  NAND2_X1 U18624 ( .A1(n15194), .A2(n20374), .ZN(n15195) );
  OAI211_X1 U18625 ( .C1(n15197), .C2(n20385), .A(n15196), .B(n15195), .ZN(
        P1_U3005) );
  INV_X1 U18626 ( .A(n15198), .ZN(n15205) );
  INV_X1 U18627 ( .A(n15199), .ZN(n15200) );
  OAI211_X1 U18628 ( .C1(n15203), .C2(n15202), .A(n15201), .B(n15200), .ZN(
        n15204) );
  AOI21_X1 U18629 ( .B1(n15205), .B2(n20374), .A(n15204), .ZN(n15206) );
  OAI21_X1 U18630 ( .B1(n15207), .B2(n20385), .A(n15206), .ZN(P1_U3006) );
  NOR2_X1 U18631 ( .A1(n20816), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15214) );
  OR2_X1 U18632 ( .A1(n15208), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15210) );
  AOI21_X1 U18633 ( .B1(n15211), .B2(n15210), .A(n15209), .ZN(n15212) );
  AOI211_X1 U18634 ( .C1(n15220), .C2(n15214), .A(n15213), .B(n15212), .ZN(
        n15217) );
  NAND2_X1 U18635 ( .A1(n15215), .A2(n20374), .ZN(n15216) );
  OAI211_X1 U18636 ( .C1(n15218), .C2(n20385), .A(n15217), .B(n15216), .ZN(
        P1_U3007) );
  AOI21_X1 U18637 ( .B1(n15220), .B2(n20816), .A(n15219), .ZN(n15223) );
  NAND2_X1 U18638 ( .A1(n15221), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15222) );
  OAI211_X1 U18639 ( .C1(n15224), .C2(n20392), .A(n15223), .B(n15222), .ZN(
        n15225) );
  INV_X1 U18640 ( .A(n15225), .ZN(n15226) );
  OAI21_X1 U18641 ( .B1(n15227), .B2(n20385), .A(n15226), .ZN(P1_U3008) );
  INV_X1 U18642 ( .A(n15228), .ZN(n15248) );
  NAND2_X1 U18643 ( .A1(n20389), .A2(n15229), .ZN(n15234) );
  INV_X1 U18644 ( .A(n15235), .ZN(n15292) );
  NAND3_X1 U18645 ( .A1(n15232), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n15292), .ZN(n15233) );
  NAND2_X1 U18646 ( .A1(n15234), .A2(n15233), .ZN(n15291) );
  NOR2_X1 U18647 ( .A1(n15291), .A2(n15293), .ZN(n15254) );
  AOI211_X1 U18648 ( .C1(n15235), .C2(n15234), .A(n10164), .B(n15254), .ZN(
        n15265) );
  NAND2_X1 U18649 ( .A1(n15265), .A2(n9856), .ZN(n15245) );
  AOI211_X1 U18650 ( .C1(n15238), .C2(n15237), .A(n15236), .B(n15245), .ZN(
        n15239) );
  AOI211_X1 U18651 ( .C1(n15248), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15240), .B(n15239), .ZN(n15243) );
  NAND2_X1 U18652 ( .A1(n15241), .A2(n20374), .ZN(n15242) );
  OAI211_X1 U18653 ( .C1(n15244), .C2(n20385), .A(n15243), .B(n15242), .ZN(
        P1_U3009) );
  NOR2_X1 U18654 ( .A1(n15245), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15246) );
  AOI211_X1 U18655 ( .C1(n15248), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15247), .B(n15246), .ZN(n15251) );
  NAND2_X1 U18656 ( .A1(n15249), .A2(n20374), .ZN(n15250) );
  OAI211_X1 U18657 ( .C1(n15252), .C2(n20385), .A(n15251), .B(n15250), .ZN(
        P1_U3010) );
  NAND2_X1 U18658 ( .A1(n15253), .A2(n16379), .ZN(n15259) );
  OAI21_X1 U18659 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15254), .A(
        n15261), .ZN(n15257) );
  AND3_X1 U18660 ( .A1(n15265), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n20987), .ZN(n15255) );
  AOI211_X1 U18661 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15257), .A(
        n15256), .B(n15255), .ZN(n15258) );
  OAI211_X1 U18662 ( .C1(n20392), .C2(n16220), .A(n15259), .B(n15258), .ZN(
        P1_U3011) );
  NAND2_X1 U18663 ( .A1(n15260), .A2(n16379), .ZN(n15267) );
  INV_X1 U18664 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15264) );
  NOR2_X1 U18665 ( .A1(n15261), .A2(n15264), .ZN(n15262) );
  AOI211_X1 U18666 ( .C1(n15265), .C2(n15264), .A(n15263), .B(n15262), .ZN(
        n15266) );
  OAI211_X1 U18667 ( .C1(n20392), .C2(n15268), .A(n15267), .B(n15266), .ZN(
        P1_U3012) );
  NAND2_X1 U18668 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n16327), .ZN(
        n15270) );
  OAI21_X1 U18669 ( .B1(n15325), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16348), .ZN(n16334) );
  AOI21_X1 U18670 ( .B1(n16368), .B2(n15270), .A(n16334), .ZN(n16333) );
  INV_X1 U18671 ( .A(n16333), .ZN(n15273) );
  NAND2_X1 U18672 ( .A1(n15269), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16339) );
  NOR3_X1 U18673 ( .A1(n16339), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15270), .ZN(n15271) );
  AOI211_X1 U18674 ( .C1(n15273), .C2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15272), .B(n15271), .ZN(n15276) );
  INV_X1 U18675 ( .A(n16236), .ZN(n15274) );
  NAND2_X1 U18676 ( .A1(n15274), .A2(n20374), .ZN(n15275) );
  OAI211_X1 U18677 ( .C1(n15277), .C2(n20385), .A(n15276), .B(n15275), .ZN(
        P1_U3013) );
  INV_X1 U18678 ( .A(n15278), .ZN(n15280) );
  OAI21_X1 U18679 ( .B1(n15281), .B2(n15280), .A(n15279), .ZN(n15283) );
  XNOR2_X1 U18680 ( .A(n15283), .B(n15282), .ZN(n16291) );
  NAND2_X1 U18681 ( .A1(n16291), .A2(n16379), .ZN(n15289) );
  INV_X1 U18682 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15284) );
  NOR2_X1 U18683 ( .A1(n20254), .A2(n15284), .ZN(n15287) );
  AOI211_X1 U18684 ( .C1(n11602), .C2(n15285), .A(n16327), .B(n16339), .ZN(
        n15286) );
  AOI211_X1 U18685 ( .C1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n16334), .A(
        n15287), .B(n15286), .ZN(n15288) );
  OAI211_X1 U18686 ( .C1(n20392), .C2(n16244), .A(n15289), .B(n15288), .ZN(
        P1_U3015) );
  NAND2_X1 U18687 ( .A1(n15290), .A2(n16379), .ZN(n15299) );
  INV_X1 U18688 ( .A(n16348), .ZN(n15297) );
  AOI21_X1 U18689 ( .B1(n15293), .B2(n15292), .A(n15291), .ZN(n15294) );
  NOR2_X1 U18690 ( .A1(n15294), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15295) );
  AOI211_X1 U18691 ( .C1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n15297), .A(
        n15296), .B(n15295), .ZN(n15298) );
  OAI211_X1 U18692 ( .C1(n20392), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        P1_U3018) );
  OAI21_X1 U18693 ( .B1(n16349), .B2(n16357), .A(n20389), .ZN(n15301) );
  OAI211_X1 U18694 ( .C1(n15304), .C2(n15303), .A(n15302), .B(n15301), .ZN(
        n16353) );
  AOI21_X1 U18695 ( .B1(n20382), .B2(n16349), .A(n16353), .ZN(n15314) );
  NOR3_X1 U18696 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16349), .A3(
        n16357), .ZN(n15305) );
  NAND2_X1 U18697 ( .A1(n16370), .A2(n15305), .ZN(n15312) );
  NOR2_X1 U18698 ( .A1(n15307), .A2(n15306), .ZN(n15308) );
  AOI21_X1 U18699 ( .B1(n9820), .B2(n20374), .A(n15310), .ZN(n15311) );
  OAI211_X1 U18700 ( .C1(n15314), .C2(n15313), .A(n15312), .B(n15311), .ZN(
        n15315) );
  AOI21_X1 U18701 ( .B1(n15316), .B2(n16379), .A(n15315), .ZN(n15317) );
  INV_X1 U18702 ( .A(n15317), .ZN(P1_U3019) );
  NAND3_X1 U18703 ( .A1(n15318), .A2(n16379), .A3(n13279), .ZN(n15328) );
  INV_X1 U18704 ( .A(n15319), .ZN(n15323) );
  NOR2_X1 U18705 ( .A1(n20392), .A2(n15320), .ZN(n15321) );
  AOI211_X1 U18706 ( .C1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n15323), .A(
        n15322), .B(n15321), .ZN(n15327) );
  OR3_X1 U18707 ( .A1(n15325), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n15324), .ZN(n15326) );
  NAND3_X1 U18708 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(P1_U3030) );
  NOR3_X1 U18709 ( .A1(n15329), .A2(n12893), .A3(n13231), .ZN(n15330) );
  AOI211_X1 U18710 ( .C1(n15333), .C2(n15332), .A(n15331), .B(n15330), .ZN(
        n16164) );
  INV_X1 U18711 ( .A(n15334), .ZN(n15340) );
  NOR3_X1 U18712 ( .A1(n13231), .A2(n12893), .A3(n15335), .ZN(n15336) );
  AOI21_X1 U18713 ( .B1(n15338), .B2(n15337), .A(n15336), .ZN(n15339) );
  OAI21_X1 U18714 ( .B1(n16164), .B2(n15340), .A(n15339), .ZN(n15342) );
  MUX2_X1 U18715 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15342), .S(
        n15341), .Z(P1_U3473) );
  NOR2_X1 U18716 ( .A1(n15344), .A2(n15343), .ZN(n15345) );
  NAND2_X1 U18717 ( .A1(n15365), .A2(n15386), .ZN(n15348) );
  NAND2_X1 U18718 ( .A1(n15349), .A2(n15348), .ZN(n15610) );
  OAI21_X1 U18719 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15350), .A(
        n15360), .ZN(n16461) );
  AOI21_X1 U18720 ( .B1(n16487), .B2(n15358), .A(n15350), .ZN(n16479) );
  INV_X1 U18721 ( .A(n16479), .ZN(n15411) );
  INV_X1 U18722 ( .A(n15356), .ZN(n15352) );
  INV_X1 U18723 ( .A(n15359), .ZN(n15351) );
  OAI21_X1 U18724 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n15352), .A(
        n15351), .ZN(n15665) );
  AOI21_X1 U18725 ( .B1(n15690), .B2(n15353), .A(n15357), .ZN(n19190) );
  OAI21_X1 U18726 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n15354), .A(
        n15353), .ZN(n19207) );
  NAND2_X1 U18727 ( .A1(n15355), .A2(n19207), .ZN(n19188) );
  NOR2_X1 U18728 ( .A1(n19190), .A2(n19188), .ZN(n19180) );
  OAI21_X1 U18729 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15357), .A(
        n15356), .ZN(n19179) );
  NAND2_X1 U18730 ( .A1(n19180), .A2(n19179), .ZN(n19178) );
  NAND2_X1 U18731 ( .A1(n15347), .A2(n19178), .ZN(n15439) );
  NAND2_X1 U18732 ( .A1(n15665), .A2(n15439), .ZN(n15438) );
  NAND2_X1 U18733 ( .A1(n16408), .A2(n15438), .ZN(n15426) );
  OAI21_X1 U18734 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15359), .A(
        n15358), .ZN(n16494) );
  NAND2_X1 U18735 ( .A1(n16408), .A2(n15425), .ZN(n15410) );
  NAND2_X1 U18736 ( .A1(n15411), .A2(n15410), .ZN(n15409) );
  NAND2_X1 U18737 ( .A1(n16408), .A2(n15409), .ZN(n16460) );
  NAND2_X1 U18738 ( .A1(n16461), .A2(n16460), .ZN(n16459) );
  NAND2_X1 U18739 ( .A1(n16408), .A2(n16459), .ZN(n15397) );
  INV_X1 U18740 ( .A(n15360), .ZN(n15362) );
  INV_X1 U18741 ( .A(n15363), .ZN(n15361) );
  OAI21_X1 U18742 ( .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n15362), .A(
        n15361), .ZN(n15629) );
  NAND2_X1 U18743 ( .A1(n16408), .A2(n15396), .ZN(n16450) );
  OR2_X1 U18744 ( .A1(n15363), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15364) );
  NAND2_X1 U18745 ( .A1(n15365), .A2(n15364), .ZN(n16451) );
  NAND2_X1 U18746 ( .A1(n16408), .A2(n16449), .ZN(n15384) );
  NAND2_X1 U18747 ( .A1(n15610), .A2(n15384), .ZN(n15383) );
  NAND2_X1 U18748 ( .A1(n16408), .A2(n15383), .ZN(n16436) );
  NAND2_X1 U18749 ( .A1(n16437), .A2(n16436), .ZN(n16435) );
  NAND2_X1 U18750 ( .A1(n15347), .A2(n16435), .ZN(n15368) );
  NOR2_X1 U18751 ( .A1(n15366), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15367) );
  OR2_X1 U18752 ( .A1(n15587), .A2(n15367), .ZN(n15603) );
  OAI211_X1 U18753 ( .C1(n15368), .C2(n15603), .A(n19316), .B(n16407), .ZN(
        n15378) );
  AOI21_X1 U18754 ( .B1(n15370), .B2(n9784), .A(n15369), .ZN(n15794) );
  INV_X1 U18755 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20116) );
  OAI22_X1 U18756 ( .A1(n9999), .A2(n19306), .B1(n20116), .B2(n19305), .ZN(
        n15373) );
  NOR2_X1 U18757 ( .A1(n19324), .A2(n15371), .ZN(n15372) );
  AOI211_X1 U18758 ( .C1(n15794), .C2(n19339), .A(n15373), .B(n15372), .ZN(
        n15374) );
  OAI21_X1 U18759 ( .B1(n15375), .B2(n19308), .A(n15374), .ZN(n15376) );
  INV_X1 U18760 ( .A(n15376), .ZN(n15377) );
  OAI211_X1 U18761 ( .C1(n15797), .C2(n19346), .A(n15378), .B(n15377), .ZN(
        P2_U2826) );
  NAND2_X1 U18762 ( .A1(n15379), .A2(n15380), .ZN(n15381) );
  NAND2_X1 U18763 ( .A1(n15382), .A2(n15381), .ZN(n15807) );
  OAI211_X1 U18764 ( .C1(n15384), .C2(n15610), .A(n19316), .B(n15383), .ZN(
        n15394) );
  INV_X1 U18765 ( .A(n15385), .ZN(n15392) );
  OAI22_X1 U18766 ( .A1(n15386), .A2(n19306), .B1(n15608), .B2(n19305), .ZN(
        n15391) );
  OR2_X1 U18767 ( .A1(n15558), .A2(n15387), .ZN(n15388) );
  NAND2_X1 U18768 ( .A1(n11166), .A2(n15388), .ZN(n15803) );
  INV_X1 U18769 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n15389) );
  OAI22_X1 U18770 ( .A1(n15803), .A2(n19323), .B1(n19324), .B2(n15389), .ZN(
        n15390) );
  AOI211_X1 U18771 ( .C1(n19341), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15393) );
  OAI211_X1 U18772 ( .C1(n19346), .C2(n15807), .A(n15394), .B(n15393), .ZN(
        P2_U2828) );
  INV_X1 U18773 ( .A(n15395), .ZN(n15408) );
  OAI211_X1 U18774 ( .C1(n15397), .C2(n15629), .A(n19316), .B(n15396), .ZN(
        n15407) );
  AOI21_X1 U18775 ( .B1(n15399), .B2(n15513), .A(n15398), .ZN(n15825) );
  OAI22_X1 U18776 ( .A1(n15630), .A2(n19306), .B1(n10925), .B2(n19305), .ZN(
        n15405) );
  NAND2_X1 U18777 ( .A1(n15400), .A2(n15401), .ZN(n15402) );
  NAND2_X1 U18778 ( .A1(n15557), .A2(n15402), .ZN(n15828) );
  INV_X1 U18779 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n15403) );
  OAI22_X1 U18780 ( .A1(n15828), .A2(n19323), .B1(n19324), .B2(n15403), .ZN(
        n15404) );
  AOI211_X1 U18781 ( .C1(n15825), .C2(n19315), .A(n15405), .B(n15404), .ZN(
        n15406) );
  OAI211_X1 U18782 ( .C1(n19308), .C2(n15408), .A(n15407), .B(n15406), .ZN(
        P2_U2830) );
  OAI211_X1 U18783 ( .C1(n15411), .C2(n15410), .A(n19316), .B(n15409), .ZN(
        n15422) );
  NAND2_X1 U18784 ( .A1(n9810), .A2(n15413), .ZN(n15414) );
  AND2_X1 U18785 ( .A1(n15515), .A2(n15414), .ZN(n16551) );
  OAI22_X1 U18786 ( .A1(n16487), .A2(n19306), .B1(n11157), .B2(n19305), .ZN(
        n15420) );
  NOR2_X1 U18787 ( .A1(n10171), .A2(n15416), .ZN(n15417) );
  OR2_X1 U18788 ( .A1(n15415), .A2(n15417), .ZN(n16547) );
  INV_X1 U18789 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n15418) );
  OAI22_X1 U18790 ( .A1(n16547), .A2(n19323), .B1(n19324), .B2(n15418), .ZN(
        n15419) );
  AOI211_X1 U18791 ( .C1(n16551), .C2(n19315), .A(n15420), .B(n15419), .ZN(
        n15421) );
  OAI211_X1 U18792 ( .C1(n15423), .C2(n19308), .A(n15422), .B(n15421), .ZN(
        P2_U2832) );
  INV_X1 U18793 ( .A(n15424), .ZN(n15436) );
  OAI211_X1 U18794 ( .C1(n16494), .C2(n15426), .A(n19316), .B(n15425), .ZN(
        n15435) );
  OR2_X1 U18795 ( .A1(n15442), .A2(n15427), .ZN(n15428) );
  AND2_X1 U18796 ( .A1(n9810), .A2(n15428), .ZN(n16491) );
  AOI22_X1 U18797 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19343), .ZN(n15429) );
  INV_X1 U18798 ( .A(n15429), .ZN(n15433) );
  XNOR2_X1 U18799 ( .A(n15446), .B(n15431), .ZN(n16473) );
  INV_X1 U18800 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n20926) );
  OAI22_X1 U18801 ( .A1(n16473), .A2(n19323), .B1(n19324), .B2(n20926), .ZN(
        n15432) );
  AOI211_X1 U18802 ( .C1(n16491), .C2(n19315), .A(n15433), .B(n15432), .ZN(
        n15434) );
  OAI211_X1 U18803 ( .C1(n15436), .C2(n19308), .A(n15435), .B(n15434), .ZN(
        P2_U2833) );
  INV_X1 U18804 ( .A(n15437), .ZN(n15453) );
  OAI211_X1 U18805 ( .C1(n15439), .C2(n15665), .A(n19316), .B(n15438), .ZN(
        n15452) );
  AND2_X1 U18806 ( .A1(n15535), .A2(n15440), .ZN(n15441) );
  NOR2_X1 U18807 ( .A1(n15442), .A2(n15441), .ZN(n15671) );
  OAI22_X1 U18808 ( .A1(n15443), .A2(n19306), .B1(n15663), .B2(n19305), .ZN(
        n15449) );
  NAND2_X1 U18809 ( .A1(n14090), .A2(n15444), .ZN(n15445) );
  NAND2_X1 U18810 ( .A1(n15446), .A2(n15445), .ZN(n15862) );
  NAND2_X1 U18811 ( .A1(n19342), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n15447) );
  OAI21_X1 U18812 ( .B1(n15862), .B2(n19323), .A(n15447), .ZN(n15448) );
  OR2_X1 U18813 ( .A1(n15449), .A2(n15448), .ZN(n15450) );
  AOI21_X1 U18814 ( .B1(n15671), .B2(n19315), .A(n15450), .ZN(n15451) );
  OAI211_X1 U18815 ( .C1(n19308), .C2(n15453), .A(n15452), .B(n15451), .ZN(
        P2_U2834) );
  NAND2_X1 U18816 ( .A1(n19343), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18817 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n19342), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19351), .ZN(n15454) );
  OAI211_X1 U18818 ( .C1(n19308), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15457) );
  AOI21_X1 U18819 ( .B1(n19339), .B2(n20147), .A(n15457), .ZN(n15458) );
  OAI21_X1 U18820 ( .B1(n10013), .B2(n19346), .A(n15458), .ZN(n15464) );
  INV_X1 U18821 ( .A(n15461), .ZN(n15462) );
  NOR2_X1 U18822 ( .A1(n19331), .A2(n15459), .ZN(n15467) );
  INV_X1 U18823 ( .A(n15467), .ZN(n15460) );
  AOI221_X1 U18824 ( .B1(n15462), .B2(n15467), .C1(n15461), .C2(n15460), .A(
        n20056), .ZN(n15463) );
  AOI211_X1 U18825 ( .C1(n15465), .C2(n19349), .A(n15464), .B(n15463), .ZN(
        n15466) );
  INV_X1 U18826 ( .A(n15466), .ZN(P2_U2853) );
  OAI21_X1 U18827 ( .B1(n19355), .B2(n15468), .A(n15467), .ZN(n16009) );
  INV_X1 U18828 ( .A(n15469), .ZN(n15472) );
  INV_X1 U18829 ( .A(n15470), .ZN(n19350) );
  AOI22_X1 U18830 ( .A1(n19341), .A2(n15472), .B1(n15471), .B2(n19350), .ZN(
        n15474) );
  NAND2_X1 U18831 ( .A1(n19339), .A2(n20157), .ZN(n15473) );
  OAI211_X1 U18832 ( .C1(n19492), .C2(n19346), .A(n15474), .B(n15473), .ZN(
        n15478) );
  AOI22_X1 U18833 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19343), .ZN(n15475) );
  OAI21_X1 U18834 ( .B1(n19324), .B2(n15476), .A(n15475), .ZN(n15477) );
  AOI211_X1 U18835 ( .C1(n19349), .C2(n19573), .A(n15478), .B(n15477), .ZN(
        n15479) );
  OAI21_X1 U18836 ( .B1(n16009), .B2(n20056), .A(n15479), .ZN(P2_U2854) );
  NAND2_X1 U18837 ( .A1(n15481), .A2(n15480), .ZN(n15541) );
  NAND3_X1 U18838 ( .A1(n9785), .A2(n15527), .A3(n15541), .ZN(n15483) );
  NAND2_X1 U18839 ( .A1(n9726), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15482) );
  OAI211_X1 U18840 ( .C1(n9726), .C2(n15797), .A(n15483), .B(n15482), .ZN(
        P2_U2858) );
  NOR2_X1 U18841 ( .A1(n15485), .A2(n15484), .ZN(n15486) );
  XOR2_X1 U18842 ( .A(n15487), .B(n15486), .Z(n15550) );
  NOR2_X1 U18843 ( .A1(n15488), .A2(n9726), .ZN(n15489) );
  AOI21_X1 U18844 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n9726), .A(n15489), .ZN(
        n15490) );
  OAI21_X1 U18845 ( .B1(n15550), .B2(n15539), .A(n15490), .ZN(P2_U2859) );
  AOI21_X1 U18846 ( .B1(n15493), .B2(n15492), .A(n15491), .ZN(n15554) );
  NAND2_X1 U18847 ( .A1(n15554), .A2(n15527), .ZN(n15495) );
  NAND2_X1 U18848 ( .A1(n9726), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15494) );
  OAI211_X1 U18849 ( .C1(n15807), .C2(n9726), .A(n15495), .B(n15494), .ZN(
        P2_U2860) );
  OAI21_X1 U18850 ( .B1(n15498), .B2(n15497), .A(n15496), .ZN(n15563) );
  NAND2_X1 U18851 ( .A1(n9726), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n15502) );
  OR2_X1 U18852 ( .A1(n15398), .A2(n15499), .ZN(n15500) );
  AND2_X1 U18853 ( .A1(n15500), .A2(n15379), .ZN(n16442) );
  NAND2_X1 U18854 ( .A1(n16442), .A2(n15537), .ZN(n15501) );
  OAI211_X1 U18855 ( .C1(n15563), .C2(n15539), .A(n15502), .B(n15501), .ZN(
        P2_U2861) );
  OAI21_X1 U18856 ( .B1(n15505), .B2(n15504), .A(n15503), .ZN(n15568) );
  NAND2_X1 U18857 ( .A1(n9726), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n15507) );
  NAND2_X1 U18858 ( .A1(n15825), .A2(n15537), .ZN(n15506) );
  OAI211_X1 U18859 ( .C1(n15568), .C2(n15539), .A(n15507), .B(n15506), .ZN(
        P2_U2862) );
  AOI21_X1 U18860 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(n15511) );
  XOR2_X1 U18861 ( .A(n15512), .B(n15511), .Z(n15575) );
  NAND2_X1 U18862 ( .A1(n9726), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n15518) );
  INV_X1 U18863 ( .A(n15513), .ZN(n15514) );
  AOI21_X1 U18864 ( .B1(n15516), .B2(n15515), .A(n15514), .ZN(n16458) );
  NAND2_X1 U18865 ( .A1(n16458), .A2(n15537), .ZN(n15517) );
  OAI211_X1 U18866 ( .C1(n15575), .C2(n15539), .A(n15518), .B(n15517), .ZN(
        P2_U2863) );
  INV_X1 U18867 ( .A(n16551), .ZN(n15524) );
  AOI21_X1 U18868 ( .B1(n15521), .B2(n15520), .A(n15519), .ZN(n16468) );
  NAND2_X1 U18869 ( .A1(n16468), .A2(n15527), .ZN(n15523) );
  NAND2_X1 U18870 ( .A1(n9726), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15522) );
  OAI211_X1 U18871 ( .C1(n15524), .C2(n9726), .A(n15523), .B(n15522), .ZN(
        P2_U2864) );
  AOI21_X1 U18872 ( .B1(n15526), .B2(n15525), .A(n14516), .ZN(n16475) );
  NAND2_X1 U18873 ( .A1(n16475), .A2(n15527), .ZN(n15529) );
  NAND2_X1 U18874 ( .A1(n16491), .A2(n15537), .ZN(n15528) );
  OAI211_X1 U18875 ( .C1(n15537), .C2(n20926), .A(n15529), .B(n15528), .ZN(
        P2_U2865) );
  OAI21_X1 U18876 ( .B1(n9827), .B2(n15530), .A(n15525), .ZN(n15586) );
  INV_X1 U18877 ( .A(n15671), .ZN(n15867) );
  MUX2_X1 U18878 ( .A(n10665), .B(n15867), .S(n15537), .Z(n15531) );
  OAI21_X1 U18879 ( .B1(n15586), .B2(n15539), .A(n15531), .ZN(P2_U2866) );
  NAND2_X1 U18880 ( .A1(n15533), .A2(n15532), .ZN(n15534) );
  AND2_X1 U18881 ( .A1(n15535), .A2(n15534), .ZN(n19184) );
  INV_X1 U18882 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n20999) );
  NOR2_X1 U18883 ( .A1(n15537), .A2(n20999), .ZN(n15536) );
  AOI21_X1 U18884 ( .B1(n19184), .B2(n15537), .A(n15536), .ZN(n15538) );
  OAI21_X1 U18885 ( .B1(n15540), .B2(n15539), .A(n15538), .ZN(P2_U2867) );
  NAND3_X1 U18886 ( .A1(n9785), .A2(n19417), .A3(n15541), .ZN(n15545) );
  INV_X1 U18887 ( .A(n19387), .ZN(n19415) );
  AOI22_X1 U18888 ( .A1(n16472), .A2(n19365), .B1(n19415), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15544) );
  AOI22_X1 U18889 ( .A1(n15794), .A2(n19416), .B1(n19357), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n15543) );
  NAND2_X1 U18890 ( .A1(n19356), .A2(BUF1_REG_29__SCAN_IN), .ZN(n15542) );
  NAND4_X1 U18891 ( .A1(n15545), .A2(n15544), .A3(n15543), .A4(n15542), .ZN(
        P2_U2890) );
  OAI22_X1 U18892 ( .A1(n15577), .A2(n19368), .B1(n19387), .B2(n15546), .ZN(
        n15547) );
  AOI21_X1 U18893 ( .B1(n16433), .B2(n19416), .A(n15547), .ZN(n15549) );
  AOI22_X1 U18894 ( .A1(n19357), .A2(BUF2_REG_28__SCAN_IN), .B1(n19356), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15548) );
  OAI211_X1 U18895 ( .C1(n15550), .C2(n19390), .A(n15549), .B(n15548), .ZN(
        P2_U2891) );
  INV_X1 U18896 ( .A(n19416), .ZN(n19360) );
  AOI22_X1 U18897 ( .A1(n16472), .A2(n19371), .B1(n19415), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15552) );
  AOI22_X1 U18898 ( .A1(n19357), .A2(BUF2_REG_27__SCAN_IN), .B1(n19356), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15551) );
  OAI211_X1 U18899 ( .C1(n15803), .C2(n19360), .A(n15552), .B(n15551), .ZN(
        n15553) );
  AOI21_X1 U18900 ( .B1(n15554), .B2(n19417), .A(n15553), .ZN(n15555) );
  INV_X1 U18901 ( .A(n15555), .ZN(P2_U2892) );
  AND2_X1 U18902 ( .A1(n15557), .A2(n15556), .ZN(n15559) );
  OR2_X1 U18903 ( .A1(n15559), .A2(n15558), .ZN(n16454) );
  INV_X1 U18904 ( .A(n16454), .ZN(n15816) );
  OAI22_X1 U18905 ( .A1(n15577), .A2(n19374), .B1(n19387), .B2(n20871), .ZN(
        n15560) );
  AOI21_X1 U18906 ( .B1(n15816), .B2(n19416), .A(n15560), .ZN(n15562) );
  AOI22_X1 U18907 ( .A1(n19357), .A2(BUF2_REG_26__SCAN_IN), .B1(n19356), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15561) );
  OAI211_X1 U18908 ( .C1(n15563), .C2(n19390), .A(n15562), .B(n15561), .ZN(
        P2_U2893) );
  AOI22_X1 U18909 ( .A1(n19357), .A2(BUF2_REG_25__SCAN_IN), .B1(n19356), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15565) );
  AOI22_X1 U18910 ( .A1(n16472), .A2(n19377), .B1(n19415), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15564) );
  OAI211_X1 U18911 ( .C1(n19360), .C2(n15828), .A(n15565), .B(n15564), .ZN(
        n15566) );
  INV_X1 U18912 ( .A(n15566), .ZN(n15567) );
  OAI21_X1 U18913 ( .B1(n15568), .B2(n19390), .A(n15567), .ZN(P2_U2894) );
  OAI21_X1 U18914 ( .B1(n15415), .B2(n15569), .A(n15400), .ZN(n15570) );
  INV_X1 U18915 ( .A(n15570), .ZN(n16457) );
  OAI22_X1 U18916 ( .A1(n15577), .A2(n19380), .B1(n19387), .B2(n15571), .ZN(
        n15572) );
  AOI21_X1 U18917 ( .B1(n16457), .B2(n19416), .A(n15572), .ZN(n15574) );
  AOI22_X1 U18918 ( .A1(n19357), .A2(BUF2_REG_24__SCAN_IN), .B1(n19356), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15573) );
  OAI211_X1 U18919 ( .C1(n15575), .C2(n19390), .A(n15574), .B(n15573), .ZN(
        P2_U2895) );
  INV_X1 U18920 ( .A(n15862), .ZN(n15584) );
  OAI22_X1 U18921 ( .A1(n15577), .A2(n19395), .B1(n15576), .B2(n19387), .ZN(
        n15583) );
  INV_X1 U18922 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15580) );
  INV_X1 U18923 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15578) );
  OAI22_X1 U18924 ( .A1(n15581), .A2(n15580), .B1(n15579), .B2(n15578), .ZN(
        n15582) );
  AOI211_X1 U18925 ( .C1(n19416), .C2(n15584), .A(n15583), .B(n15582), .ZN(
        n15585) );
  OAI21_X1 U18926 ( .B1(n15586), .B2(n19390), .A(n15585), .ZN(P2_U2898) );
  XNOR2_X1 U18927 ( .A(n15587), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16427) );
  NOR2_X1 U18928 ( .A1(n16427), .A2(n19471), .ZN(n15588) );
  AOI211_X1 U18929 ( .C1(n19473), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15589), .B(n15588), .ZN(n15590) );
  OAI21_X1 U18930 ( .B1(n16422), .B2(n13256), .A(n15590), .ZN(n15591) );
  AOI21_X1 U18931 ( .B1(n15592), .B2(n19475), .A(n15591), .ZN(n15593) );
  OAI21_X1 U18932 ( .B1(n15594), .B2(n16514), .A(n15593), .ZN(P2_U2984) );
  INV_X1 U18933 ( .A(n15596), .ZN(n15597) );
  NOR2_X1 U18934 ( .A1(n15598), .A2(n15597), .ZN(n15599) );
  XNOR2_X1 U18935 ( .A(n15595), .B(n15599), .ZN(n15802) );
  AOI21_X1 U18936 ( .B1(n15808), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15601) );
  NOR2_X1 U18937 ( .A1(n15601), .A2(n15600), .ZN(n15800) );
  NOR2_X1 U18938 ( .A1(n15797), .A2(n13256), .ZN(n15605) );
  NAND2_X1 U18939 ( .A1(n19326), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15792) );
  NAND2_X1 U18940 ( .A1(n19473), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15602) );
  OAI211_X1 U18941 ( .C1(n15603), .C2(n19471), .A(n15792), .B(n15602), .ZN(
        n15604) );
  AOI211_X1 U18942 ( .C1(n15800), .C2(n19475), .A(n15605), .B(n15604), .ZN(
        n15606) );
  OAI21_X1 U18943 ( .B1(n15802), .B2(n16514), .A(n15606), .ZN(P2_U2985) );
  XNOR2_X1 U18944 ( .A(n15607), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15812) );
  INV_X1 U18945 ( .A(n15807), .ZN(n15614) );
  NOR2_X1 U18946 ( .A1(n19304), .A2(n15608), .ZN(n15805) );
  AOI21_X1 U18947 ( .B1(n19473), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15805), .ZN(n15609) );
  OAI21_X1 U18948 ( .B1(n15610), .B2(n19471), .A(n15609), .ZN(n15613) );
  INV_X1 U18949 ( .A(n15621), .ZN(n15611) );
  NOR3_X1 U18950 ( .A1(n15809), .A2(n15808), .A3(n19464), .ZN(n15612) );
  AOI211_X2 U18951 ( .C1(n19480), .C2(n15614), .A(n15613), .B(n15612), .ZN(
        n15615) );
  OAI21_X1 U18952 ( .B1(n15812), .B2(n16514), .A(n15615), .ZN(P2_U2987) );
  AND2_X1 U18953 ( .A1(n15616), .A2(n15624), .ZN(n15627) );
  NOR2_X1 U18954 ( .A1(n15627), .A2(n15623), .ZN(n15617) );
  XOR2_X1 U18955 ( .A(n15618), .B(n15617), .Z(n15824) );
  NOR2_X1 U18956 ( .A1(n19304), .A2(n20111), .ZN(n15815) );
  AOI21_X1 U18957 ( .B1(n19473), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15815), .ZN(n15619) );
  OAI21_X1 U18958 ( .B1(n16451), .B2(n19471), .A(n15619), .ZN(n15622) );
  INV_X1 U18959 ( .A(n15623), .ZN(n15625) );
  AOI21_X1 U18960 ( .B1(n15625), .B2(n15624), .A(n15616), .ZN(n15628) );
  INV_X1 U18961 ( .A(n15616), .ZN(n15626) );
  OAI22_X1 U18962 ( .A1(n15628), .A2(n15627), .B1(n15626), .B2(n15625), .ZN(
        n15837) );
  NOR2_X1 U18963 ( .A1(n15629), .A2(n19471), .ZN(n15632) );
  NAND2_X1 U18964 ( .A1(n19326), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15826) );
  OAI21_X1 U18965 ( .B1(n16541), .B2(n15630), .A(n15826), .ZN(n15631) );
  AOI211_X1 U18966 ( .C1(n15825), .C2(n19480), .A(n15632), .B(n15631), .ZN(
        n15636) );
  NAND2_X1 U18967 ( .A1(n15845), .A2(n15634), .ZN(n15834) );
  NAND3_X1 U18968 ( .A1(n9924), .A2(n19475), .A3(n15834), .ZN(n15635) );
  OAI211_X1 U18969 ( .C1(n15837), .C2(n16514), .A(n15636), .B(n15635), .ZN(
        P2_U2989) );
  XNOR2_X1 U18970 ( .A(n15637), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15638) );
  XNOR2_X1 U18971 ( .A(n9791), .B(n15638), .ZN(n15849) );
  NOR2_X1 U18972 ( .A1(n19304), .A2(n20109), .ZN(n15838) );
  AOI21_X1 U18973 ( .B1(n19473), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15838), .ZN(n15639) );
  OAI21_X1 U18974 ( .B1(n16461), .B2(n19471), .A(n15639), .ZN(n15640) );
  AOI21_X1 U18975 ( .B1(n16458), .B2(n19480), .A(n15640), .ZN(n15644) );
  INV_X1 U18976 ( .A(n15641), .ZN(n15642) );
  NAND2_X1 U18977 ( .A1(n15642), .A2(n15840), .ZN(n15846) );
  NAND3_X1 U18978 ( .A1(n15846), .A2(n19475), .A3(n15845), .ZN(n15643) );
  OAI211_X1 U18979 ( .C1(n15849), .C2(n16514), .A(n15644), .B(n15643), .ZN(
        P2_U2990) );
  NAND3_X1 U18980 ( .A1(n15646), .A2(n15754), .A3(n15739), .ZN(n15647) );
  OAI21_X1 U18981 ( .B1(n15648), .B2(n15647), .A(n15740), .ZN(n15732) );
  INV_X1 U18982 ( .A(n15730), .ZN(n15649) );
  INV_X1 U18983 ( .A(n15721), .ZN(n15650) );
  INV_X1 U18984 ( .A(n15652), .ZN(n15653) );
  NAND2_X1 U18985 ( .A1(n15653), .A2(n15654), .ZN(n15704) );
  INV_X1 U18986 ( .A(n15655), .ZN(n15687) );
  NAND3_X1 U18987 ( .A1(n15698), .A2(n15687), .A3(n15695), .ZN(n15677) );
  INV_X1 U18988 ( .A(n15656), .ZN(n15657) );
  NAND3_X1 U18989 ( .A1(n15677), .A2(n15657), .A3(n15674), .ZN(n15673) );
  NAND2_X1 U18990 ( .A1(n15673), .A2(n15674), .ZN(n15662) );
  INV_X1 U18991 ( .A(n15658), .ZN(n15659) );
  NOR2_X1 U18992 ( .A1(n15660), .A2(n15659), .ZN(n15661) );
  XNOR2_X1 U18993 ( .A(n15662), .B(n15661), .ZN(n15872) );
  NOR2_X1 U18994 ( .A1(n19304), .A2(n15663), .ZN(n15864) );
  AOI21_X1 U18995 ( .B1(n19473), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15864), .ZN(n15664) );
  OAI21_X1 U18996 ( .B1(n19471), .B2(n15665), .A(n15664), .ZN(n15670) );
  NAND2_X1 U18997 ( .A1(n15666), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15684) );
  NOR2_X1 U18998 ( .A1(n15684), .A2(n15879), .ZN(n15668) );
  OAI21_X1 U18999 ( .B1(n15668), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16482), .ZN(n15860) );
  NOR2_X1 U19000 ( .A1(n15860), .A2(n19464), .ZN(n15669) );
  AOI211_X1 U19001 ( .C1(n19480), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15672) );
  OAI21_X1 U19002 ( .B1(n15872), .B2(n16514), .A(n15672), .ZN(P2_U2993) );
  XNOR2_X1 U19003 ( .A(n15684), .B(n15879), .ZN(n15884) );
  INV_X1 U19004 ( .A(n15673), .ZN(n15679) );
  AOI22_X1 U19005 ( .A1(n15677), .A2(n15676), .B1(n15675), .B2(n15674), .ZN(
        n15678) );
  NAND2_X1 U19006 ( .A1(n15873), .A2(n16538), .ZN(n15683) );
  NOR2_X1 U19007 ( .A1(n19304), .A2(n20103), .ZN(n15874) );
  AOI21_X1 U19008 ( .B1(n19473), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15874), .ZN(n15680) );
  OAI21_X1 U19009 ( .B1(n19471), .B2(n19179), .A(n15680), .ZN(n15681) );
  AOI21_X1 U19010 ( .B1(n19184), .B2(n19480), .A(n15681), .ZN(n15682) );
  OAI211_X1 U19011 ( .C1(n19464), .C2(n15884), .A(n15683), .B(n15682), .ZN(
        P2_U2994) );
  OAI21_X1 U19012 ( .B1(n15666), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15684), .ZN(n15895) );
  INV_X1 U19013 ( .A(n15696), .ZN(n15685) );
  OAI21_X1 U19014 ( .B1(n15698), .B2(n15685), .A(n15695), .ZN(n15689) );
  NAND2_X1 U19015 ( .A1(n15687), .A2(n15686), .ZN(n15688) );
  XNOR2_X1 U19016 ( .A(n15689), .B(n15688), .ZN(n15885) );
  NAND2_X1 U19017 ( .A1(n15885), .A2(n16538), .ZN(n15694) );
  NAND2_X1 U19018 ( .A1(n19326), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15888) );
  OAI21_X1 U19019 ( .B1(n16541), .B2(n15690), .A(n15888), .ZN(n15692) );
  NOR2_X1 U19020 ( .A1(n19195), .A2(n13256), .ZN(n15691) );
  AOI211_X1 U19021 ( .C1(n16530), .C2(n19190), .A(n15692), .B(n15691), .ZN(
        n15693) );
  OAI211_X1 U19022 ( .C1(n19464), .C2(n15895), .A(n15694), .B(n15693), .ZN(
        P2_U2995) );
  NAND2_X1 U19023 ( .A1(n15696), .A2(n15695), .ZN(n15697) );
  XNOR2_X1 U19024 ( .A(n15698), .B(n15697), .ZN(n15911) );
  AOI21_X1 U19025 ( .B1(n15900), .B2(n9753), .A(n15666), .ZN(n15908) );
  NOR2_X1 U19026 ( .A1(n19304), .A2(n20099), .ZN(n15902) );
  NOR2_X1 U19027 ( .A1(n19471), .A2(n19207), .ZN(n15699) );
  AOI211_X1 U19028 ( .C1(n19473), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15902), .B(n15699), .ZN(n15700) );
  OAI21_X1 U19029 ( .B1(n19206), .B2(n13256), .A(n15700), .ZN(n15701) );
  AOI21_X1 U19030 ( .B1(n15908), .B2(n19475), .A(n15701), .ZN(n15702) );
  OAI21_X1 U19031 ( .B1(n15911), .B2(n16514), .A(n15702), .ZN(P2_U2996) );
  XOR2_X1 U19032 ( .A(n15704), .B(n15703), .Z(n15929) );
  NAND2_X1 U19033 ( .A1(n19326), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15913) );
  OAI21_X1 U19034 ( .B1(n16541), .B2(n15705), .A(n15913), .ZN(n15707) );
  NOR2_X1 U19035 ( .A1(n15912), .A2(n13256), .ZN(n15706) );
  AOI211_X1 U19036 ( .C1(n16530), .C2(n15708), .A(n15707), .B(n15706), .ZN(
        n15712) );
  AND2_X2 U19037 ( .A1(n15709), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16512) );
  AND2_X2 U19038 ( .A1(n16512), .A2(n16582), .ZN(n16496) );
  INV_X1 U19039 ( .A(n15957), .ZN(n15953) );
  NAND2_X2 U19040 ( .A1(n16496), .A2(n15953), .ZN(n15743) );
  NOR2_X2 U19041 ( .A1(n15743), .A2(n15958), .ZN(n15918) );
  NAND2_X1 U19042 ( .A1(n15918), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15717) );
  INV_X1 U19043 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15710) );
  OAI211_X1 U19044 ( .C1(n15923), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n19475), .B(n9753), .ZN(n15711) );
  OAI211_X1 U19045 ( .C1(n15929), .C2(n16514), .A(n15712), .B(n15711), .ZN(
        P2_U2997) );
  XNOR2_X1 U19046 ( .A(n15714), .B(n15713), .ZN(n15936) );
  NOR2_X1 U19047 ( .A1(n20808), .A2(n19304), .ZN(n15716) );
  OAI22_X1 U19048 ( .A1(n10007), .A2(n16541), .B1(n19471), .B2(n19218), .ZN(
        n15715) );
  AOI211_X1 U19049 ( .C1(n19480), .C2(n19220), .A(n15716), .B(n15715), .ZN(
        n15720) );
  XNOR2_X1 U19050 ( .A(n15717), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15718) );
  NAND2_X1 U19051 ( .A1(n15718), .A2(n19475), .ZN(n15719) );
  OAI211_X1 U19052 ( .C1(n15936), .C2(n16514), .A(n15720), .B(n15719), .ZN(
        P2_U2998) );
  NAND2_X1 U19053 ( .A1(n15722), .A2(n15721), .ZN(n15724) );
  XOR2_X1 U19054 ( .A(n15724), .B(n15723), .Z(n15949) );
  XNOR2_X1 U19055 ( .A(n15918), .B(n15944), .ZN(n15947) );
  NAND2_X1 U19056 ( .A1(n19326), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15939) );
  OAI21_X1 U19057 ( .B1(n16541), .B2(n19228), .A(n15939), .ZN(n15725) );
  AOI21_X1 U19058 ( .B1(n16530), .B2(n19226), .A(n15725), .ZN(n15726) );
  OAI21_X1 U19059 ( .B1(n19232), .B2(n13256), .A(n15726), .ZN(n15727) );
  AOI21_X1 U19060 ( .B1(n15947), .B2(n19475), .A(n15727), .ZN(n15728) );
  OAI21_X1 U19061 ( .B1(n15949), .B2(n16514), .A(n15728), .ZN(P2_U2999) );
  NAND2_X1 U19062 ( .A1(n15730), .A2(n15729), .ZN(n15731) );
  XNOR2_X1 U19063 ( .A(n15732), .B(n15731), .ZN(n15965) );
  AOI21_X1 U19064 ( .B1(n15958), .B2(n15743), .A(n15918), .ZN(n15950) );
  OAI22_X1 U19065 ( .A1(n11129), .A2(n19304), .B1(n19471), .B2(n19241), .ZN(
        n15736) );
  INV_X1 U19066 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15733) );
  OAI22_X1 U19067 ( .A1(n15734), .A2(n13256), .B1(n15733), .B2(n16541), .ZN(
        n15735) );
  AOI211_X1 U19068 ( .C1(n15950), .C2(n19475), .A(n15736), .B(n15735), .ZN(
        n15737) );
  OAI21_X1 U19069 ( .B1(n16514), .B2(n15965), .A(n15737), .ZN(P2_U3000) );
  NAND2_X1 U19070 ( .A1(n15740), .A2(n15739), .ZN(n15741) );
  XNOR2_X1 U19071 ( .A(n15738), .B(n15741), .ZN(n16561) );
  INV_X1 U19072 ( .A(n16561), .ZN(n15751) );
  NAND2_X1 U19073 ( .A1(n16496), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15756) );
  NAND2_X1 U19074 ( .A1(n15756), .A2(n15742), .ZN(n15744) );
  AND2_X1 U19075 ( .A1(n15744), .A2(n15743), .ZN(n16560) );
  OAI22_X1 U19076 ( .A1(n15745), .A2(n16541), .B1(n10891), .B2(n19304), .ZN(
        n15749) );
  INV_X1 U19077 ( .A(n15746), .ZN(n15747) );
  OAI22_X1 U19078 ( .A1(n13256), .A2(n16558), .B1(n19471), .B2(n15747), .ZN(
        n15748) );
  AOI211_X1 U19079 ( .C1(n16560), .C2(n19475), .A(n15749), .B(n15748), .ZN(
        n15750) );
  OAI21_X1 U19080 ( .B1(n15751), .B2(n16514), .A(n15750), .ZN(P2_U3001) );
  NAND2_X1 U19081 ( .A1(n10143), .A2(n15754), .ZN(n15755) );
  XNOR2_X1 U19082 ( .A(n15752), .B(n15755), .ZN(n16577) );
  OAI21_X1 U19083 ( .B1(n16496), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15756), .ZN(n16573) );
  INV_X1 U19084 ( .A(n16573), .ZN(n15759) );
  OAI22_X1 U19085 ( .A1(n11097), .A2(n19304), .B1(n19471), .B2(n19253), .ZN(
        n15758) );
  OAI22_X1 U19086 ( .A1(n13256), .A2(n19255), .B1(n10004), .B2(n16541), .ZN(
        n15757) );
  AOI211_X1 U19087 ( .C1(n15759), .C2(n19475), .A(n15758), .B(n15757), .ZN(
        n15760) );
  OAI21_X1 U19088 ( .B1(n16577), .B2(n16514), .A(n15760), .ZN(P2_U3002) );
  OR2_X1 U19089 ( .A1(n15761), .A2(n15969), .ZN(n15766) );
  INV_X1 U19090 ( .A(n15762), .ZN(n15763) );
  AND2_X1 U19091 ( .A1(n15764), .A2(n15763), .ZN(n15765) );
  XNOR2_X1 U19092 ( .A(n15766), .B(n15765), .ZN(n16606) );
  NAND2_X1 U19093 ( .A1(n16512), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16497) );
  OAI21_X1 U19094 ( .B1(n16512), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16497), .ZN(n16602) );
  INV_X1 U19095 ( .A(n16602), .ZN(n15769) );
  OAI22_X1 U19096 ( .A1(n11067), .A2(n19304), .B1(n19471), .B2(n19261), .ZN(
        n15768) );
  OAI22_X1 U19097 ( .A1(n13256), .A2(n19268), .B1(n16541), .B2(n10003), .ZN(
        n15767) );
  AOI211_X1 U19098 ( .C1(n15769), .C2(n19475), .A(n15768), .B(n15767), .ZN(
        n15770) );
  OAI21_X1 U19099 ( .B1(n16606), .B2(n16514), .A(n15770), .ZN(P2_U3004) );
  INV_X1 U19100 ( .A(n15982), .ZN(n15772) );
  AOI21_X1 U19101 ( .B1(n15771), .B2(n15981), .A(n15772), .ZN(n15776) );
  NAND2_X1 U19102 ( .A1(n15774), .A2(n15773), .ZN(n15775) );
  XNOR2_X1 U19103 ( .A(n15776), .B(n15775), .ZN(n16619) );
  NAND2_X1 U19104 ( .A1(n15778), .A2(n15777), .ZN(n15779) );
  AND2_X1 U19105 ( .A1(n15780), .A2(n15779), .ZN(n16616) );
  OAI22_X1 U19106 ( .A1(n11037), .A2(n19304), .B1(n19471), .B2(n19288), .ZN(
        n15784) );
  INV_X1 U19107 ( .A(n19290), .ZN(n15782) );
  INV_X1 U19108 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n15781) );
  OAI22_X1 U19109 ( .A1(n15782), .A2(n13256), .B1(n16541), .B2(n15781), .ZN(
        n15783) );
  AOI211_X1 U19110 ( .C1(n16616), .C2(n19475), .A(n15784), .B(n15783), .ZN(
        n15785) );
  OAI21_X1 U19111 ( .B1(n16619), .B2(n16514), .A(n15785), .ZN(P2_U3006) );
  INV_X1 U19112 ( .A(n15786), .ZN(n15788) );
  AOI21_X1 U19113 ( .B1(n15788), .B2(n15787), .A(n15790), .ZN(n15799) );
  INV_X1 U19114 ( .A(n15789), .ZN(n15811) );
  NAND3_X1 U19115 ( .A1(n15811), .A2(n15791), .A3(n15790), .ZN(n15796) );
  INV_X1 U19116 ( .A(n15792), .ZN(n15793) );
  AOI21_X1 U19117 ( .B1(n15794), .B2(n16621), .A(n15793), .ZN(n15795) );
  OAI211_X1 U19118 ( .C1(n19491), .C2(n15797), .A(n15796), .B(n15795), .ZN(
        n15798) );
  OAI21_X1 U19119 ( .B1(n15802), .B2(n19500), .A(n15801), .ZN(P2_U3017) );
  NOR2_X1 U19120 ( .A1(n15803), .A2(n19487), .ZN(n15804) );
  NAND2_X1 U19121 ( .A1(n15829), .A2(n15840), .ZN(n15842) );
  INV_X1 U19122 ( .A(n15813), .ZN(n15841) );
  NAND2_X1 U19123 ( .A1(n15842), .A2(n15841), .ZN(n15833) );
  INV_X1 U19124 ( .A(n16442), .ZN(n15819) );
  OAI21_X1 U19125 ( .B1(n15840), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15814) );
  OAI211_X1 U19126 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15829), .B(n15814), .ZN(
        n15818) );
  AOI21_X1 U19127 ( .B1(n15816), .B2(n16621), .A(n15815), .ZN(n15817) );
  OAI211_X1 U19128 ( .C1(n15819), .C2(n19491), .A(n15818), .B(n15817), .ZN(
        n15822) );
  NOR2_X1 U19129 ( .A1(n15820), .A2(n19490), .ZN(n15821) );
  OAI21_X1 U19130 ( .B1(n15824), .B2(n19500), .A(n15823), .ZN(P2_U3020) );
  NAND2_X1 U19131 ( .A1(n15825), .A2(n16635), .ZN(n15827) );
  OAI211_X1 U19132 ( .C1(n19487), .C2(n15828), .A(n15827), .B(n15826), .ZN(
        n15832) );
  INV_X1 U19133 ( .A(n15829), .ZN(n15830) );
  NOR3_X1 U19134 ( .A1(n15830), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n15840), .ZN(n15831) );
  AOI211_X1 U19135 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n15833), .A(
        n15832), .B(n15831), .ZN(n15836) );
  NAND3_X1 U19136 ( .A1(n9924), .A2(n16624), .A3(n15834), .ZN(n15835) );
  OAI211_X1 U19137 ( .C1(n15837), .C2(n19500), .A(n15836), .B(n15835), .ZN(
        P2_U3021) );
  AOI21_X1 U19138 ( .B1(n16457), .B2(n16621), .A(n15838), .ZN(n15839) );
  OAI21_X1 U19139 ( .B1(n15841), .B2(n15840), .A(n15839), .ZN(n15844) );
  INV_X1 U19140 ( .A(n15842), .ZN(n15843) );
  AOI211_X1 U19141 ( .C1(n16635), .C2(n16458), .A(n15844), .B(n15843), .ZN(
        n15848) );
  NAND3_X1 U19142 ( .A1(n15846), .A2(n16624), .A3(n15845), .ZN(n15847) );
  OAI211_X1 U19143 ( .C1(n15849), .C2(n19500), .A(n15848), .B(n15847), .ZN(
        P2_U3022) );
  NAND2_X1 U19144 ( .A1(n9913), .A2(n15852), .ZN(n15853) );
  XNOR2_X1 U19145 ( .A(n15850), .B(n15853), .ZN(n16489) );
  NAND2_X1 U19146 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19326), .ZN(n15854) );
  OAI221_X1 U19147 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16544), 
        .C1(n16546), .C2(n16555), .A(n15854), .ZN(n15857) );
  NAND2_X1 U19148 ( .A1(n16491), .A2(n16635), .ZN(n15855) );
  OAI21_X1 U19149 ( .B1(n16473), .B2(n19487), .A(n15855), .ZN(n15856) );
  NOR2_X1 U19150 ( .A1(n15857), .A2(n15856), .ZN(n15859) );
  XNOR2_X1 U19151 ( .A(n16482), .B(n16546), .ZN(n16488) );
  OR2_X1 U19152 ( .A1(n16488), .A2(n19490), .ZN(n15858) );
  OAI211_X1 U19153 ( .C1(n16489), .C2(n19500), .A(n15859), .B(n15858), .ZN(
        P2_U3024) );
  INV_X1 U19154 ( .A(n15860), .ZN(n15870) );
  INV_X1 U19155 ( .A(n15892), .ZN(n15877) );
  NOR3_X1 U19156 ( .A1(n15877), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15861), .ZN(n15869) );
  INV_X1 U19157 ( .A(n15861), .ZN(n15878) );
  OAI21_X1 U19158 ( .B1(n15878), .B2(n19485), .A(n15886), .ZN(n15865) );
  NOR2_X1 U19159 ( .A1(n19487), .A2(n15862), .ZN(n15863) );
  AOI211_X1 U19160 ( .C1(n15865), .C2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15864), .B(n15863), .ZN(n15866) );
  OAI21_X1 U19161 ( .B1(n15867), .B2(n19491), .A(n15866), .ZN(n15868) );
  AOI211_X1 U19162 ( .C1(n15870), .C2(n16624), .A(n15869), .B(n15868), .ZN(
        n15871) );
  OAI21_X1 U19163 ( .B1(n15872), .B2(n19500), .A(n15871), .ZN(P2_U3025) );
  NAND2_X1 U19164 ( .A1(n15873), .A2(n16639), .ZN(n15883) );
  AOI21_X1 U19165 ( .B1(n16621), .B2(n15875), .A(n15874), .ZN(n15876) );
  OAI21_X1 U19166 ( .B1(n15886), .B2(n15879), .A(n15876), .ZN(n15881) );
  AOI211_X1 U19167 ( .C1(n15879), .C2(n15891), .A(n15878), .B(n15877), .ZN(
        n15880) );
  AOI211_X1 U19168 ( .C1(n19184), .C2(n16635), .A(n15881), .B(n15880), .ZN(
        n15882) );
  OAI211_X1 U19169 ( .C1(n15884), .C2(n19490), .A(n15883), .B(n15882), .ZN(
        P2_U3026) );
  NAND2_X1 U19170 ( .A1(n15885), .A2(n16639), .ZN(n15894) );
  NOR2_X1 U19171 ( .A1(n15886), .A2(n15891), .ZN(n15890) );
  NAND2_X1 U19172 ( .A1(n16621), .A2(n19196), .ZN(n15887) );
  OAI211_X1 U19173 ( .C1(n19195), .C2(n19491), .A(n15888), .B(n15887), .ZN(
        n15889) );
  AOI211_X1 U19174 ( .C1(n15892), .C2(n15891), .A(n15890), .B(n15889), .ZN(
        n15893) );
  OAI211_X1 U19175 ( .C1(n15895), .C2(n19490), .A(n15894), .B(n15893), .ZN(
        P2_U3027) );
  INV_X1 U19176 ( .A(n15896), .ZN(n15897) );
  OR2_X1 U19177 ( .A1(n16579), .A2(n15897), .ZN(n15898) );
  NAND2_X1 U19178 ( .A1(n15898), .A2(n16578), .ZN(n15945) );
  OAI21_X1 U19179 ( .B1(n15899), .B2(n19485), .A(n15945), .ZN(n15907) );
  NAND3_X1 U19180 ( .A1(n16581), .A2(n15901), .A3(n15900), .ZN(n15905) );
  AOI21_X1 U19181 ( .B1(n16621), .B2(n15903), .A(n15902), .ZN(n15904) );
  OAI211_X1 U19182 ( .C1(n19206), .C2(n19491), .A(n15905), .B(n15904), .ZN(
        n15906) );
  AOI21_X1 U19183 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15907), .A(
        n15906), .ZN(n15910) );
  NAND2_X1 U19184 ( .A1(n15908), .A2(n16624), .ZN(n15909) );
  OAI211_X1 U19185 ( .C1(n15911), .C2(n19500), .A(n15910), .B(n15909), .ZN(
        P2_U3028) );
  INV_X1 U19186 ( .A(n15912), .ZN(n15922) );
  OAI21_X1 U19187 ( .B1(n19487), .B2(n15914), .A(n15913), .ZN(n15921) );
  NAND2_X1 U19188 ( .A1(n16581), .A2(n15915), .ZN(n16566) );
  INV_X1 U19189 ( .A(n15916), .ZN(n15917) );
  NOR2_X1 U19190 ( .A1(n16566), .A2(n15917), .ZN(n15937) );
  NOR3_X1 U19191 ( .A1(n15930), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15919), .ZN(n15920) );
  NOR2_X1 U19192 ( .A1(n19485), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15926) );
  OAI21_X1 U19193 ( .B1(n15933), .B2(n15926), .A(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15927) );
  OAI211_X1 U19194 ( .C1(n15929), .C2(n19500), .A(n15928), .B(n15927), .ZN(
        P2_U3029) );
  OAI22_X1 U19195 ( .A1(n19487), .A2(n19224), .B1(n20808), .B2(n19304), .ZN(
        n15932) );
  NOR3_X1 U19196 ( .A1(n15930), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15944), .ZN(n15931) );
  NAND2_X1 U19197 ( .A1(n15933), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15934) );
  OAI211_X1 U19198 ( .C1(n15936), .C2(n19500), .A(n15935), .B(n15934), .ZN(
        P2_U3030) );
  NAND2_X1 U19199 ( .A1(n15937), .A2(n15944), .ZN(n15943) );
  INV_X1 U19200 ( .A(n19232), .ZN(n15941) );
  XNOR2_X1 U19201 ( .A(n15938), .B(n15954), .ZN(n19362) );
  OAI21_X1 U19202 ( .B1(n19487), .B2(n19362), .A(n15939), .ZN(n15940) );
  AOI21_X1 U19203 ( .B1(n15941), .B2(n16635), .A(n15940), .ZN(n15942) );
  OAI211_X1 U19204 ( .C1(n15945), .C2(n15944), .A(n15943), .B(n15942), .ZN(
        n15946) );
  AOI21_X1 U19205 ( .B1(n15947), .B2(n16624), .A(n15946), .ZN(n15948) );
  OAI21_X1 U19206 ( .B1(n15949), .B2(n19500), .A(n15948), .ZN(P2_U3031) );
  NAND2_X1 U19207 ( .A1(n15950), .A2(n16624), .ZN(n15964) );
  NAND2_X1 U19208 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16582), .ZN(
        n15951) );
  AOI21_X1 U19209 ( .B1(n15952), .B2(n15951), .A(n15972), .ZN(n16568) );
  OAI21_X1 U19210 ( .B1(n16566), .B2(n15953), .A(n16568), .ZN(n16557) );
  INV_X1 U19211 ( .A(n15954), .ZN(n15955) );
  OAI21_X1 U19212 ( .B1(n15956), .B2(n13554), .A(n15955), .ZN(n19364) );
  NAND2_X1 U19213 ( .A1(n19243), .A2(n16635), .ZN(n15961) );
  NOR2_X1 U19214 ( .A1(n15957), .A2(n16566), .ZN(n15959) );
  AOI22_X1 U19215 ( .A1(n19326), .A2(P2_REIP_REG_14__SCAN_IN), .B1(n15959), 
        .B2(n15958), .ZN(n15960) );
  OAI211_X1 U19216 ( .C1(n19487), .C2(n19364), .A(n15961), .B(n15960), .ZN(
        n15962) );
  AOI21_X1 U19217 ( .B1(n16557), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15962), .ZN(n15963) );
  OAI211_X1 U19218 ( .C1(n15965), .C2(n19500), .A(n15964), .B(n15963), .ZN(
        P2_U3032) );
  NOR2_X1 U19219 ( .A1(n15709), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16513) );
  NOR3_X1 U19220 ( .A1(n16513), .A2(n16512), .A3(n19490), .ZN(n15980) );
  INV_X1 U19221 ( .A(n15761), .ZN(n15970) );
  OAI21_X1 U19222 ( .B1(n15967), .B2(n15969), .A(n15966), .ZN(n15968) );
  OAI21_X1 U19223 ( .B1(n15970), .B2(n15969), .A(n15968), .ZN(n16515) );
  NOR2_X1 U19224 ( .A1(n11054), .A2(n19304), .ZN(n15971) );
  AOI221_X1 U19225 ( .B1(n15972), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n16581), .C2(n16580), .A(n15971), .ZN(n15978) );
  INV_X1 U19226 ( .A(n15973), .ZN(n15974) );
  XNOR2_X1 U19227 ( .A(n15975), .B(n15974), .ZN(n19379) );
  OAI22_X1 U19228 ( .A1(n19491), .A2(n19279), .B1(n19487), .B2(n19379), .ZN(
        n15976) );
  INV_X1 U19229 ( .A(n15976), .ZN(n15977) );
  OAI211_X1 U19230 ( .C1(n16515), .C2(n19500), .A(n15978), .B(n15977), .ZN(
        n15979) );
  OR2_X1 U19231 ( .A1(n15980), .A2(n15979), .ZN(P2_U3037) );
  NAND2_X1 U19232 ( .A1(n15982), .A2(n15981), .ZN(n15983) );
  XNOR2_X1 U19233 ( .A(n15771), .B(n15983), .ZN(n16522) );
  INV_X1 U19234 ( .A(n16522), .ZN(n15998) );
  XNOR2_X1 U19235 ( .A(n15985), .B(n15984), .ZN(n15986) );
  XNOR2_X1 U19236 ( .A(n15987), .B(n15986), .ZN(n16521) );
  NOR3_X1 U19237 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n15989), .A3(
        n15988), .ZN(n16614) );
  NOR2_X1 U19238 ( .A1(n10858), .A2(n19304), .ZN(n15990) );
  AOI211_X1 U19239 ( .C1(n16615), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16614), .B(n15990), .ZN(n15991) );
  INV_X1 U19240 ( .A(n15991), .ZN(n15996) );
  INV_X1 U19241 ( .A(n15992), .ZN(n15994) );
  XNOR2_X1 U19242 ( .A(n15994), .B(n15993), .ZN(n19383) );
  OAI22_X1 U19243 ( .A1(n19383), .A2(n19487), .B1(n19491), .B2(n19299), .ZN(
        n15995) );
  AOI211_X1 U19244 ( .C1(n16521), .C2(n16624), .A(n15996), .B(n15995), .ZN(
        n15997) );
  OAI21_X1 U19245 ( .B1(n15998), .B2(n19500), .A(n15997), .ZN(P2_U3039) );
  OAI22_X1 U19246 ( .A1(n15347), .A2(n12964), .B1(n19355), .B2(n19331), .ZN(
        n16010) );
  INV_X1 U19247 ( .A(n16043), .ZN(n16027) );
  INV_X1 U19248 ( .A(n10320), .ZN(n16036) );
  INV_X1 U19249 ( .A(n15999), .ZN(n16000) );
  NOR2_X1 U19250 ( .A1(n16000), .A2(n10940), .ZN(n16006) );
  OAI21_X1 U19251 ( .B1(n19347), .B2(n16027), .A(n16001), .ZN(n16663) );
  AOI22_X1 U19252 ( .A1(n16663), .A2(n19153), .B1(n16002), .B2(n16688), .ZN(
        n16003) );
  OAI21_X1 U19253 ( .B1(n16010), .B2(n16011), .A(n16003), .ZN(n16004) );
  MUX2_X1 U19254 ( .A(n16004), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n16045), .Z(P2_U3601) );
  XNOR2_X1 U19255 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16005) );
  OAI22_X1 U19256 ( .A1(n16006), .A2(n16005), .B1(n16036), .B2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16007) );
  AOI21_X1 U19257 ( .B1(n16008), .B2(n16043), .A(n16007), .ZN(n16664) );
  OAI21_X1 U19258 ( .B1(n15347), .B2(n19493), .A(n16009), .ZN(n16028) );
  INV_X1 U19259 ( .A(n16010), .ZN(n16012) );
  NOR2_X1 U19260 ( .A1(n16012), .A2(n16011), .ZN(n16029) );
  INV_X1 U19261 ( .A(n16029), .ZN(n16013) );
  OAI22_X1 U19262 ( .A1(n16664), .A2(n20133), .B1(n16028), .B2(n16013), .ZN(
        n16014) );
  AOI21_X1 U19263 ( .B1(n19573), .B2(n16688), .A(n16014), .ZN(n16016) );
  NAND2_X1 U19264 ( .A1(n16045), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n16015) );
  OAI21_X1 U19265 ( .B1(n16016), .B2(n16045), .A(n16015), .ZN(P2_U3600) );
  NOR2_X1 U19266 ( .A1(n16017), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16037) );
  NOR2_X1 U19267 ( .A1(n16037), .A2(n16033), .ZN(n16025) );
  NOR2_X1 U19268 ( .A1(n16019), .A2(n16018), .ZN(n16034) );
  INV_X1 U19269 ( .A(n16034), .ZN(n16024) );
  NOR3_X1 U19270 ( .A1(n16036), .A2(n16020), .A3(n10784), .ZN(n16023) );
  NOR2_X1 U19271 ( .A1(n16021), .A2(n16658), .ZN(n16038) );
  NOR2_X1 U19272 ( .A1(n16038), .A2(n16025), .ZN(n16022) );
  AOI211_X1 U19273 ( .C1(n16025), .C2(n16024), .A(n16023), .B(n16022), .ZN(
        n16026) );
  OAI21_X1 U19274 ( .B1(n10013), .B2(n16027), .A(n16026), .ZN(n16649) );
  AOI22_X1 U19275 ( .A1(n16649), .A2(n19153), .B1(n16029), .B2(n16028), .ZN(
        n16030) );
  OAI21_X1 U19276 ( .B1(n20145), .B2(n16044), .A(n16030), .ZN(n16031) );
  MUX2_X1 U19277 ( .A(n16031), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16045), .Z(P2_U3599) );
  INV_X1 U19278 ( .A(n10784), .ZN(n16035) );
  AOI21_X1 U19279 ( .B1(n10320), .B2(n16035), .A(n16037), .ZN(n16032) );
  OAI21_X1 U19280 ( .B1(n16034), .B2(n16033), .A(n16032), .ZN(n16041) );
  OAI22_X1 U19281 ( .A1(n16038), .A2(n16037), .B1(n16036), .B2(n16035), .ZN(
        n16040) );
  MUX2_X1 U19282 ( .A(n16041), .B(n16040), .S(n16039), .Z(n16042) );
  AOI211_X1 U19283 ( .C1(n13064), .C2(n16043), .A(n10432), .B(n16042), .ZN(
        n16644) );
  OAI22_X1 U19284 ( .A1(n19549), .A2(n16044), .B1(n20133), .B2(n16644), .ZN(
        n16046) );
  MUX2_X1 U19285 ( .A(n16046), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16045), .Z(P2_U3596) );
  INV_X1 U19286 ( .A(n19988), .ZN(n16047) );
  NAND2_X1 U19287 ( .A1(n16047), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n16051) );
  AOI22_X1 U19288 ( .A1(n19941), .A2(n20046), .B1(n20041), .B2(n19982), .ZN(
        n16050) );
  NAND2_X1 U19289 ( .A1(n19985), .A2(n20043), .ZN(n16049) );
  NAND2_X1 U19290 ( .A1(n20045), .A2(n19984), .ZN(n16048) );
  NAND4_X1 U19291 ( .A1(n16051), .A2(n16050), .A3(n16049), .A4(n16048), .ZN(
        P2_U3167) );
  INV_X1 U19292 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16885) );
  INV_X1 U19293 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16057) );
  NOR3_X1 U19294 ( .A1(n16053), .A2(n17647), .A3(n16052), .ZN(n16055) );
  NOR2_X2 U19295 ( .A1(n16054), .A2(n18962), .ZN(n16138) );
  INV_X1 U19296 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n17148) );
  NAND3_X1 U19297 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17504) );
  NOR3_X1 U19298 ( .A1(n17148), .A2(n17164), .A3(n17504), .ZN(n17379) );
  INV_X1 U19299 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17099) );
  INV_X1 U19300 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17497) );
  NOR4_X1 U19301 ( .A1(n17099), .A2(n17435), .A3(n17497), .A4(n17499), .ZN(
        n16056) );
  NAND4_X1 U19302 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(n16056), .ZN(n17380) );
  NAND2_X1 U19303 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17421), .ZN(n17406) );
  NAND3_X1 U19304 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(n17346), .ZN(n17318) );
  NAND2_X1 U19305 ( .A1(n18516), .A2(n17290), .ZN(n17291) );
  NAND2_X1 U19306 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17265), .ZN(n17259) );
  NAND2_X1 U19307 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17264), .ZN(n17249) );
  NAND2_X1 U19308 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n17253), .ZN(n17239) );
  NAND2_X1 U19309 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17243), .ZN(n17238) );
  INV_X2 U19310 ( .A(n17520), .ZN(n17508) );
  AOI21_X1 U19311 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n17508), .A(n17243), .ZN(
        n16058) );
  INV_X1 U19312 ( .A(n16058), .ZN(n16133) );
  AOI22_X1 U19313 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16062) );
  AOI22_X1 U19314 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16061) );
  AOI22_X1 U19315 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16060) );
  AOI22_X1 U19316 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16059) );
  NAND4_X1 U19317 ( .A1(n16062), .A2(n16061), .A3(n16060), .A4(n16059), .ZN(
        n16068) );
  AOI22_X1 U19318 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16066) );
  AOI22_X1 U19319 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n17479), .B1(
        n17439), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16065) );
  AOI22_X1 U19320 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n16064) );
  AOI22_X1 U19321 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16063) );
  NAND4_X1 U19322 ( .A1(n16066), .A2(n16065), .A3(n16064), .A4(n16063), .ZN(
        n16067) );
  NOR2_X1 U19323 ( .A1(n16068), .A2(n16067), .ZN(n16132) );
  AOI22_X1 U19324 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16072) );
  AOI22_X1 U19325 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n17454), .B1(
        n17227), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16071) );
  AOI22_X1 U19326 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17460), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16070) );
  AOI22_X1 U19327 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16069) );
  NAND4_X1 U19328 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        n16078) );
  AOI22_X1 U19329 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U19330 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16075) );
  AOI22_X1 U19331 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16074) );
  AOI22_X1 U19332 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16073) );
  NAND4_X1 U19333 ( .A1(n16076), .A2(n16075), .A3(n16074), .A4(n16073), .ZN(
        n16077) );
  NOR2_X1 U19334 ( .A1(n16078), .A2(n16077), .ZN(n17245) );
  AOI22_X1 U19335 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16082) );
  AOI22_X1 U19336 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9729), .ZN(n16081) );
  AOI22_X1 U19337 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n16120), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16080) );
  AOI22_X1 U19338 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n16122), .ZN(n16079) );
  NAND4_X1 U19339 ( .A1(n16082), .A2(n16081), .A3(n16080), .A4(n16079), .ZN(
        n16088) );
  AOI22_X1 U19340 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17480), .B1(
        n17311), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16086) );
  AOI22_X1 U19341 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n16109), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n16085) );
  AOI22_X1 U19342 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17474), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17454), .ZN(n16084) );
  AOI22_X1 U19343 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17479), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16083) );
  NAND4_X1 U19344 ( .A1(n16086), .A2(n16085), .A3(n16084), .A4(n16083), .ZN(
        n16087) );
  NOR2_X1 U19345 ( .A1(n16088), .A2(n16087), .ZN(n17255) );
  AOI22_X1 U19346 ( .A1(n12316), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16098) );
  AOI22_X1 U19347 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16097) );
  AOI22_X1 U19348 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16089) );
  OAI21_X1 U19349 ( .B1(n20937), .B2(n12253), .A(n16089), .ZN(n16095) );
  AOI22_X1 U19350 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16093) );
  AOI22_X1 U19351 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16092) );
  AOI22_X1 U19352 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16091) );
  AOI22_X1 U19353 ( .A1(n16122), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n16090) );
  NAND4_X1 U19354 ( .A1(n16093), .A2(n16092), .A3(n16091), .A4(n16090), .ZN(
        n16094) );
  AOI211_X1 U19355 ( .C1(n17480), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n16095), .B(n16094), .ZN(n16096) );
  NAND3_X1 U19356 ( .A1(n16098), .A2(n16097), .A3(n16096), .ZN(n17261) );
  AOI22_X1 U19357 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17311), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16108) );
  AOI22_X1 U19358 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16107) );
  AOI22_X1 U19359 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16099) );
  OAI21_X1 U19360 ( .B1(n20718), .B2(n17267), .A(n16099), .ZN(n16105) );
  AOI22_X1 U19361 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16103) );
  AOI22_X1 U19362 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16102) );
  AOI22_X1 U19363 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19364 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16100) );
  NAND4_X1 U19365 ( .A1(n16103), .A2(n16102), .A3(n16101), .A4(n16100), .ZN(
        n16104) );
  AOI211_X1 U19366 ( .C1(n9734), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n16105), .B(n16104), .ZN(n16106) );
  NAND3_X1 U19367 ( .A1(n16108), .A2(n16107), .A3(n16106), .ZN(n17262) );
  NAND2_X1 U19368 ( .A1(n17261), .A2(n17262), .ZN(n17260) );
  NOR2_X1 U19369 ( .A1(n17255), .A2(n17260), .ZN(n17254) );
  AOI22_X1 U19370 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16119) );
  AOI22_X1 U19371 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16118) );
  AOI22_X1 U19372 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16110) );
  OAI21_X1 U19373 ( .B1(n20777), .B2(n10151), .A(n16110), .ZN(n16116) );
  AOI22_X1 U19374 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16114) );
  AOI22_X1 U19375 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n9722), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16113) );
  AOI22_X1 U19376 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16112) );
  AOI22_X1 U19377 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n16111) );
  NAND4_X1 U19378 ( .A1(n16114), .A2(n16113), .A3(n16112), .A4(n16111), .ZN(
        n16115) );
  AOI211_X1 U19379 ( .C1(n17460), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n16116), .B(n16115), .ZN(n16117) );
  NAND3_X1 U19380 ( .A1(n16119), .A2(n16118), .A3(n16117), .ZN(n17251) );
  NAND2_X1 U19381 ( .A1(n17254), .A2(n17251), .ZN(n17250) );
  NOR2_X1 U19382 ( .A1(n17245), .A2(n17250), .ZN(n17244) );
  AOI22_X1 U19383 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16131) );
  AOI22_X1 U19384 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16130) );
  AOI22_X1 U19385 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16121) );
  OAI21_X1 U19386 ( .B1(n17267), .B2(n17507), .A(n16121), .ZN(n16128) );
  AOI22_X1 U19387 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16126) );
  AOI22_X1 U19388 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16125) );
  AOI22_X1 U19389 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16124) );
  AOI22_X1 U19390 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16122), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16123) );
  NAND4_X1 U19391 ( .A1(n16126), .A2(n16125), .A3(n16124), .A4(n16123), .ZN(
        n16127) );
  AOI211_X1 U19392 ( .C1(n17481), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n16128), .B(n16127), .ZN(n16129) );
  NAND3_X1 U19393 ( .A1(n16131), .A2(n16130), .A3(n16129), .ZN(n17241) );
  NAND2_X1 U19394 ( .A1(n17244), .A2(n17241), .ZN(n17240) );
  NOR2_X1 U19395 ( .A1(n16132), .A2(n17240), .ZN(n17236) );
  AOI21_X1 U19396 ( .B1(n16132), .B2(n17240), .A(n17236), .ZN(n17543) );
  AOI22_X1 U19397 ( .A1(n17238), .A2(n16133), .B1(n17543), .B2(n17520), .ZN(
        n16134) );
  INV_X1 U19398 ( .A(n16134), .ZN(P3_U2675) );
  NOR4_X1 U19399 ( .A1(n19004), .A2(n16816), .A3(n17678), .A4(n19130), .ZN(
        n16137) );
  INV_X1 U19400 ( .A(n18966), .ZN(n18945) );
  NOR2_X1 U19401 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19079), .ZN(n18484) );
  INV_X1 U19402 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18466) );
  NOR2_X1 U19403 ( .A1(n18466), .A2(n19077), .ZN(n16139) );
  INV_X1 U19404 ( .A(n19110), .ZN(n19107) );
  INV_X1 U19405 ( .A(n18948), .ZN(n16140) );
  AOI21_X1 U19406 ( .B1(n16140), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16141) );
  NOR3_X1 U19407 ( .A1(n16141), .A2(n18922), .A3(n18923), .ZN(n18965) );
  NAND3_X1 U19408 ( .A1(n19107), .A2(n19144), .A3(n18965), .ZN(n16142) );
  OAI21_X1 U19409 ( .B1(n19107), .B2(n16143), .A(n16142), .ZN(P3_U3284) );
  NOR2_X1 U19410 ( .A1(n16712), .A2(n18376), .ZN(n16145) );
  AOI211_X1 U19411 ( .C1(n17790), .C2(n18370), .A(n16145), .B(n16144), .ZN(
        n16146) );
  OAI211_X1 U19412 ( .C1(n18323), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18438), .B(n16146), .ZN(n16148) );
  NOR2_X1 U19413 ( .A1(n16709), .A2(n16147), .ZN(n16196) );
  AOI21_X1 U19414 ( .B1(n18455), .B2(n16148), .A(n16196), .ZN(n16157) );
  OAI21_X1 U19415 ( .B1(n16151), .B2(n16150), .A(n16149), .ZN(n16152) );
  XOR2_X1 U19416 ( .A(n16152), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16717) );
  AOI222_X1 U19417 ( .A1(n18961), .A2(n16708), .B1(n16154), .B2(n16153), .C1(
        n18339), .C2(n16711), .ZN(n16155) );
  NOR2_X1 U19418 ( .A1(n16155), .A2(n18461), .ZN(n16202) );
  AOI22_X1 U19419 ( .A1(n18378), .A2(n16717), .B1(n16202), .B2(n16713), .ZN(
        n16156) );
  NAND2_X1 U19420 ( .A1(n18444), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16722) );
  OAI211_X1 U19421 ( .C1(n16157), .C2(n16713), .A(n16156), .B(n16722), .ZN(
        P3_U2833) );
  INV_X1 U19422 ( .A(n16158), .ZN(n16169) );
  AND2_X1 U19423 ( .A1(n16159), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n16160) );
  OR3_X1 U19424 ( .A1(n16161), .A2(n16160), .A3(n20549), .ZN(n16167) );
  INV_X1 U19425 ( .A(n16167), .ZN(n16162) );
  OAI22_X1 U19426 ( .A1(n16164), .A2(n16163), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16162), .ZN(n16165) );
  OAI21_X1 U19427 ( .B1(n16167), .B2(n16166), .A(n16165), .ZN(n16168) );
  AOI222_X1 U19428 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16169), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16168), .C1(n16169), 
        .C2(n16168), .ZN(n16170) );
  AOI222_X1 U19429 ( .A1(n16172), .A2(n16171), .B1(n16172), .B2(n16170), .C1(
        n16171), .C2(n16170), .ZN(n16178) );
  OAI21_X1 U19430 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n16173), .ZN(n16174) );
  AND3_X1 U19431 ( .A1(n16176), .A2(n16175), .A3(n16174), .ZN(n16177) );
  OAI21_X1 U19432 ( .B1(n16178), .B2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n16177), .ZN(n16179) );
  NOR3_X1 U19433 ( .A1(n16181), .A2(n16180), .A3(n16179), .ZN(n16194) );
  NAND3_X1 U19434 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20697), .A3(n10118), 
        .ZN(n16182) );
  AOI22_X1 U19435 ( .A1(n16185), .A2(n16184), .B1(n16183), .B2(n16182), .ZN(
        n16396) );
  OAI221_X1 U19436 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n16194), 
        .A(n16396), .ZN(n16405) );
  INV_X1 U19437 ( .A(n16403), .ZN(n16186) );
  NOR2_X1 U19438 ( .A1(n16187), .A2(n16186), .ZN(n16188) );
  NOR2_X1 U19439 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16188), .ZN(n16192) );
  AOI211_X1 U19440 ( .C1(n20697), .C2(n20616), .A(n16189), .B(n16403), .ZN(
        n16190) );
  NAND2_X1 U19441 ( .A1(n16405), .A2(n16190), .ZN(n16191) );
  AOI22_X1 U19442 ( .A1(n16405), .A2(n16192), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16191), .ZN(n16193) );
  OAI21_X1 U19443 ( .B1(n16194), .B2(n20197), .A(n16193), .ZN(P1_U3161) );
  OAI21_X1 U19444 ( .B1(n16712), .B2(n18376), .A(n16195), .ZN(n16197) );
  AOI21_X1 U19445 ( .B1(n18455), .B2(n16197), .A(n16196), .ZN(n16205) );
  INV_X1 U19446 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16204) );
  NOR2_X1 U19447 ( .A1(n16199), .A2(n16198), .ZN(n16200) );
  XOR2_X1 U19448 ( .A(n16200), .B(n16204), .Z(n16703) );
  NOR2_X1 U19449 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16201), .ZN(
        n16698) );
  AOI22_X1 U19450 ( .A1(n18378), .A2(n16703), .B1(n16698), .B2(n16202), .ZN(
        n16203) );
  NAND2_X1 U19451 ( .A1(n18444), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16699) );
  OAI211_X1 U19452 ( .C1(n16205), .C2(n16204), .A(n16203), .B(n16699), .ZN(
        P3_U2832) );
  NAND2_X1 U19453 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20697), .ZN(n20623) );
  INV_X1 U19454 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20632) );
  NAND3_X1 U19455 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .A3(n20632), .ZN(
        n16207) );
  INV_X1 U19456 ( .A(HOLD), .ZN(n20624) );
  OAI211_X1 U19457 ( .C1(n20632), .C2(n20624), .A(P1_STATE_REG_0__SCAN_IN), 
        .B(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n16206) );
  NAND4_X1 U19458 ( .A1(n16208), .A2(n20623), .A3(n16207), .A4(n16206), .ZN(
        P1_U3195) );
  INV_X1 U19459 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16807) );
  NOR2_X1 U19460 ( .A1(n20310), .A2(n16807), .ZN(P1_U2905) );
  NOR3_X1 U19461 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19151), .A3(n20190), 
        .ZN(n16680) );
  NOR3_X1 U19462 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n16209) );
  NOR4_X1 U19463 ( .A1(n20184), .A2(n16210), .A3(n16680), .A4(n16209), .ZN(
        P2_U3178) );
  AOI221_X1 U19464 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16210), .C1(n20169), .C2(
        n16210), .A(n19999), .ZN(n20167) );
  INV_X1 U19465 ( .A(n20167), .ZN(n20164) );
  NOR2_X1 U19466 ( .A1(n16673), .A2(n20164), .ZN(P2_U3047) );
  NOR3_X1 U19467 ( .A1(n16212), .A2(n16211), .A3(n17729), .ZN(n16213) );
  INV_X1 U19468 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17759) );
  NOR2_X2 U19469 ( .A1(n16215), .A2(n17759), .ZN(n17675) );
  NAND2_X1 U19470 ( .A1(n18516), .A2(n17524), .ZN(n17577) );
  NAND2_X1 U19471 ( .A1(n16216), .A2(n17524), .ZN(n17669) );
  INV_X1 U19472 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18478) );
  OAI22_X1 U19473 ( .A1(n17669), .A2(n18478), .B1(n17666), .B2(n18161), .ZN(
        n16217) );
  INV_X1 U19474 ( .A(n16217), .ZN(n16218) );
  OAI221_X1 U19475 ( .B1(n17675), .B2(n17759), .C1(n17675), .C2(n17577), .A(
        n16218), .ZN(P3_U2735) );
  NOR2_X1 U19476 ( .A1(n16219), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n16225) );
  AOI22_X1 U19477 ( .A1(n20263), .A2(P1_EBX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20269), .ZN(n16224) );
  INV_X1 U19478 ( .A(n16220), .ZN(n16221) );
  AOI222_X1 U19479 ( .A1(n16286), .A2(n20233), .B1(n16222), .B2(n20221), .C1(
        n20253), .C2(n16221), .ZN(n16223) );
  OAI211_X1 U19480 ( .C1(n16226), .C2(n16225), .A(n16224), .B(n16223), .ZN(
        P1_U2820) );
  NOR3_X1 U19481 ( .A1(n20271), .A2(n16227), .A3(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n16228) );
  AOI21_X1 U19482 ( .B1(n20263), .B2(P1_EBX_REG_18__SCAN_IN), .A(n16228), .ZN(
        n16229) );
  OAI21_X1 U19483 ( .B1(n16230), .B2(n20654), .A(n16229), .ZN(n16231) );
  AOI211_X1 U19484 ( .C1(n20269), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20349), .B(n16231), .ZN(n16235) );
  AOI22_X1 U19485 ( .A1(n16233), .A2(n20233), .B1(n16232), .B2(n20221), .ZN(
        n16234) );
  OAI211_X1 U19486 ( .C1(n20267), .C2(n16236), .A(n16235), .B(n16234), .ZN(
        P1_U2822) );
  INV_X1 U19487 ( .A(n20227), .ZN(n16237) );
  AOI21_X1 U19488 ( .B1(n16239), .B2(n16238), .A(n16237), .ZN(n16262) );
  OAI22_X1 U19489 ( .A1(n16262), .A2(n15284), .B1(n16240), .B2(n16272), .ZN(
        n16241) );
  AOI211_X1 U19490 ( .C1(n20269), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20349), .B(n16241), .ZN(n16248) );
  INV_X1 U19491 ( .A(n16242), .ZN(n16290) );
  INV_X1 U19492 ( .A(n16279), .ZN(n16263) );
  NAND3_X1 U19493 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16257), .A3(n16263), 
        .ZN(n16251) );
  OAI21_X1 U19494 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n16243), .ZN(n16245) );
  OAI22_X1 U19495 ( .A1(n16251), .A2(n16245), .B1(n20267), .B2(n16244), .ZN(
        n16246) );
  AOI21_X1 U19496 ( .B1(n16290), .B2(n20233), .A(n16246), .ZN(n16247) );
  OAI211_X1 U19497 ( .C1(n16294), .C2(n20277), .A(n16248), .B(n16247), .ZN(
        P1_U2824) );
  AOI22_X1 U19498 ( .A1(n16335), .A2(n20253), .B1(n20263), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16249) );
  OAI211_X1 U19499 ( .C1(n20257), .C2(n16250), .A(n16249), .B(n20254), .ZN(
        n16254) );
  OAI22_X1 U19500 ( .A1(n16252), .A2(n20242), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n16251), .ZN(n16253) );
  AOI211_X1 U19501 ( .C1(n16255), .C2(n20221), .A(n16254), .B(n16253), .ZN(
        n16256) );
  OAI21_X1 U19502 ( .B1(n16262), .B2(n15114), .A(n16256), .ZN(P1_U2825) );
  AOI21_X1 U19503 ( .B1(n16257), .B2(n16263), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n16261) );
  OAI22_X1 U19504 ( .A1(n16341), .A2(n20267), .B1(n20984), .B2(n16272), .ZN(
        n16258) );
  AOI211_X1 U19505 ( .C1(n20269), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20349), .B(n16258), .ZN(n16260) );
  AOI22_X1 U19506 ( .A1(n16304), .A2(n20233), .B1(n20221), .B2(n16302), .ZN(
        n16259) );
  OAI211_X1 U19507 ( .C1(n16262), .C2(n16261), .A(n16260), .B(n16259), .ZN(
        P1_U2826) );
  AOI21_X1 U19508 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16263), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16269) );
  NAND2_X1 U19509 ( .A1(n20263), .A2(P1_EBX_REG_12__SCAN_IN), .ZN(n16264) );
  OAI211_X1 U19510 ( .C1(n20257), .C2(n20960), .A(n16264), .B(n20254), .ZN(
        n16265) );
  AOI21_X1 U19511 ( .B1(n9820), .B2(n20253), .A(n16265), .ZN(n16268) );
  AOI22_X1 U19512 ( .A1(n16266), .A2(n20221), .B1(n20233), .B2(n20709), .ZN(
        n16267) );
  OAI211_X1 U19513 ( .C1(n16270), .C2(n16269), .A(n16268), .B(n16267), .ZN(
        P1_U2828) );
  OAI22_X1 U19514 ( .A1(n16350), .A2(n20267), .B1(n16272), .B2(n16271), .ZN(
        n16273) );
  INV_X1 U19515 ( .A(n16273), .ZN(n16274) );
  OAI21_X1 U19516 ( .B1(n16313), .B2(n20277), .A(n16274), .ZN(n16275) );
  AOI211_X1 U19517 ( .C1(n20269), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n20349), .B(n16275), .ZN(n16278) );
  AOI22_X1 U19518 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16276), .B1(n20233), 
        .B2(n16310), .ZN(n16277) );
  OAI211_X1 U19519 ( .C1(P1_REIP_REG_11__SCAN_IN), .C2(n16279), .A(n16278), 
        .B(n16277), .ZN(P1_U2829) );
  AOI22_X1 U19520 ( .A1(n16282), .A2(n16281), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n16280), .ZN(n16288) );
  INV_X1 U19521 ( .A(n16283), .ZN(n16285) );
  AOI22_X1 U19522 ( .A1(n16286), .A2(n16285), .B1(n16284), .B2(DATAI_20_), 
        .ZN(n16287) );
  OAI211_X1 U19523 ( .C1(n16289), .C2(n14094), .A(n16288), .B(n16287), .ZN(
        P1_U2884) );
  AOI22_X1 U19524 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16293) );
  AOI22_X1 U19525 ( .A1(n16291), .A2(n20356), .B1(n14067), .B2(n16290), .ZN(
        n16292) );
  OAI211_X1 U19526 ( .C1(n20361), .C2(n16294), .A(n16293), .B(n16292), .ZN(
        P1_U2983) );
  OAI21_X1 U19527 ( .B1(n16297), .B2(n16296), .A(n16295), .ZN(n16299) );
  NAND2_X1 U19528 ( .A1(n16299), .A2(n16298), .ZN(n16301) );
  XNOR2_X1 U19529 ( .A(n11601), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16300) );
  XNOR2_X1 U19530 ( .A(n16301), .B(n16300), .ZN(n16342) );
  AOI22_X1 U19531 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16306) );
  AOI22_X1 U19532 ( .A1(n16304), .A2(n14067), .B1(n16303), .B2(n16302), .ZN(
        n16305) );
  OAI211_X1 U19533 ( .C1(n16342), .C2(n20203), .A(n16306), .B(n16305), .ZN(
        P1_U2985) );
  AOI22_X1 U19534 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16312) );
  NOR2_X1 U19535 ( .A1(n15140), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16308) );
  NOR2_X1 U19536 ( .A1(n15095), .A2(n13957), .ZN(n16307) );
  MUX2_X1 U19537 ( .A(n16308), .B(n16307), .S(n11601), .Z(n16309) );
  XOR2_X1 U19538 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16309), .Z(
        n16352) );
  AOI22_X1 U19539 ( .A1(n20356), .A2(n16352), .B1(n14067), .B2(n16310), .ZN(
        n16311) );
  OAI211_X1 U19540 ( .C1(n20361), .C2(n16313), .A(n16312), .B(n16311), .ZN(
        P1_U2988) );
  AOI22_X1 U19541 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16319) );
  NAND2_X1 U19542 ( .A1(n16316), .A2(n16315), .ZN(n16317) );
  XNOR2_X1 U19543 ( .A(n16314), .B(n16317), .ZN(n16380) );
  AOI22_X1 U19544 ( .A1(n16380), .A2(n20356), .B1(n14067), .B2(n20234), .ZN(
        n16318) );
  OAI211_X1 U19545 ( .C1(n20361), .C2(n20237), .A(n16319), .B(n16318), .ZN(
        P1_U2992) );
  AOI22_X1 U19546 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16325) );
  OAI21_X1 U19547 ( .B1(n16322), .B2(n16321), .A(n16320), .ZN(n16387) );
  INV_X1 U19548 ( .A(n16387), .ZN(n16323) );
  AOI22_X1 U19549 ( .A1(n16323), .A2(n20356), .B1(n14067), .B2(n20284), .ZN(
        n16324) );
  OAI211_X1 U19550 ( .C1(n20361), .C2(n20261), .A(n16325), .B(n16324), .ZN(
        P1_U2994) );
  INV_X1 U19551 ( .A(n16339), .ZN(n16326) );
  AOI21_X1 U19552 ( .B1(n16327), .B2(n16326), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16332) );
  AOI22_X1 U19553 ( .A1(n16329), .A2(n16379), .B1(n20374), .B2(n16328), .ZN(
        n16331) );
  NAND2_X1 U19554 ( .A1(n20349), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16330) );
  OAI211_X1 U19555 ( .C1(n16333), .C2(n16332), .A(n16331), .B(n16330), .ZN(
        P1_U3014) );
  AOI22_X1 U19556 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16334), .B1(
        n20349), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16338) );
  AOI22_X1 U19557 ( .A1(n16336), .A2(n16379), .B1(n20374), .B2(n16335), .ZN(
        n16337) );
  OAI211_X1 U19558 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16339), .A(
        n16338), .B(n16337), .ZN(P1_U3016) );
  NOR2_X1 U19559 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16340), .ZN(
        n16345) );
  OAI22_X1 U19560 ( .A1(n16342), .A2(n20385), .B1(n20392), .B2(n16341), .ZN(
        n16343) );
  AOI21_X1 U19561 ( .B1(n16345), .B2(n16344), .A(n16343), .ZN(n16347) );
  NAND2_X1 U19562 ( .A1(n20349), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n16346) );
  OAI211_X1 U19563 ( .C1(n16348), .C2(n20883), .A(n16347), .B(n16346), .ZN(
        P1_U3017) );
  NAND2_X1 U19564 ( .A1(n16370), .A2(n16349), .ZN(n16356) );
  OAI22_X1 U19565 ( .A1(n16350), .A2(n20392), .B1(n20254), .B2(n20646), .ZN(
        n16351) );
  INV_X1 U19566 ( .A(n16351), .ZN(n16355) );
  AOI22_X1 U19567 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16353), .B1(
        n16379), .B2(n16352), .ZN(n16354) );
  OAI211_X1 U19568 ( .C1(n16357), .C2(n16356), .A(n16355), .B(n16354), .ZN(
        P1_U3020) );
  NOR2_X1 U19569 ( .A1(n13957), .A2(n14053), .ZN(n16366) );
  OAI211_X1 U19570 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n16358), .B(n16370), .ZN(n16365) );
  AOI21_X1 U19571 ( .B1(n16360), .B2(n20374), .A(n16359), .ZN(n16364) );
  AOI22_X1 U19572 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16362), .B1(
        n16379), .B2(n16361), .ZN(n16363) );
  OAI211_X1 U19573 ( .C1(n16366), .C2(n16365), .A(n16364), .B(n16363), .ZN(
        P1_U3021) );
  AOI21_X1 U19574 ( .B1(n16369), .B2(n16368), .A(n16367), .ZN(n16382) );
  NAND2_X1 U19575 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16370), .ZN(
        n16383) );
  AOI221_X1 U19576 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16377), .C2(n20964), .A(
        n16383), .ZN(n16374) );
  OAI22_X1 U19577 ( .A1(n16372), .A2(n20392), .B1(n16371), .B2(n20254), .ZN(
        n16373) );
  AOI211_X1 U19578 ( .C1(n16375), .C2(n16379), .A(n16374), .B(n16373), .ZN(
        n16376) );
  OAI21_X1 U19579 ( .B1(n16382), .B2(n16377), .A(n16376), .ZN(P1_U3023) );
  INV_X1 U19580 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20231) );
  OAI22_X1 U19581 ( .A1(n20229), .A2(n20392), .B1(n20231), .B2(n20254), .ZN(
        n16378) );
  AOI21_X1 U19582 ( .B1(n16380), .B2(n16379), .A(n16378), .ZN(n16381) );
  OAI221_X1 U19583 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16383), .C1(
        n20964), .C2(n16382), .A(n16381), .ZN(P1_U3024) );
  OR2_X1 U19584 ( .A1(n9824), .A2(n16384), .ZN(n16385) );
  AND2_X1 U19585 ( .A1(n16386), .A2(n16385), .ZN(n20283) );
  AOI22_X1 U19586 ( .A1(n20374), .A2(n20283), .B1(n20349), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16392) );
  OAI22_X1 U19587 ( .A1(n16389), .A2(n16388), .B1(n16387), .B2(n20385), .ZN(
        n16390) );
  INV_X1 U19588 ( .A(n16390), .ZN(n16391) );
  OAI211_X1 U19589 ( .C1(n20375), .C2(n16393), .A(n16392), .B(n16391), .ZN(
        P1_U3026) );
  NAND4_X1 U19590 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_0__SCAN_IN), .A3(n20616), .A4(n16398), .ZN(n16394) );
  AND2_X1 U19591 ( .A1(n16395), .A2(n16394), .ZN(n20615) );
  AOI21_X1 U19592 ( .B1(n20615), .B2(n16397), .A(n16396), .ZN(n16402) );
  NOR2_X1 U19593 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n16398), .ZN(n16399) );
  NOR2_X1 U19594 ( .A1(n10118), .A2(n16399), .ZN(n16400) );
  AOI21_X1 U19595 ( .B1(n16400), .B2(n16405), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n16401) );
  NOR3_X1 U19596 ( .A1(n16403), .A2(n16402), .A3(n16401), .ZN(P1_U3162) );
  OAI221_X1 U19597 ( .B1(n16406), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n16406), 
        .C2(n16405), .A(n16404), .ZN(P1_U3466) );
  NAND2_X1 U19598 ( .A1(n19316), .A2(n15347), .ZN(n19354) );
  NAND2_X1 U19599 ( .A1(n15347), .A2(n16407), .ZN(n16426) );
  NAND2_X1 U19600 ( .A1(n16409), .A2(n19341), .ZN(n16413) );
  NAND3_X1 U19601 ( .A1(n16411), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16410), 
        .ZN(n16412) );
  OAI211_X1 U19602 ( .C1(n19305), .C2(n16414), .A(n16413), .B(n16412), .ZN(
        n16415) );
  AOI21_X1 U19603 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19351), .A(
        n16415), .ZN(n16419) );
  OAI22_X1 U19604 ( .A1(n14462), .A2(n19346), .B1(n16416), .B2(n19323), .ZN(
        n16417) );
  INV_X1 U19605 ( .A(n16417), .ZN(n16418) );
  OAI211_X1 U19606 ( .C1(n19354), .C2(n16425), .A(n16419), .B(n16418), .ZN(
        P2_U2824) );
  AOI22_X1 U19607 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19343), .ZN(n16431) );
  INV_X1 U19608 ( .A(n16420), .ZN(n16421) );
  AOI22_X1 U19609 ( .A1(n16421), .A2(n19341), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n19342), .ZN(n16430) );
  INV_X1 U19610 ( .A(n16422), .ZN(n16424) );
  AOI22_X1 U19611 ( .A1(n16424), .A2(n19315), .B1(n19339), .B2(n16423), .ZN(
        n16429) );
  OAI211_X1 U19612 ( .C1(n16427), .C2(n16426), .A(n19316), .B(n16425), .ZN(
        n16428) );
  NAND4_X1 U19613 ( .A1(n16431), .A2(n16430), .A3(n16429), .A4(n16428), .ZN(
        P2_U2825) );
  AOI22_X1 U19614 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19343), .ZN(n16441) );
  AOI22_X1 U19615 ( .A1(n16432), .A2(n19341), .B1(P2_EBX_REG_28__SCAN_IN), 
        .B2(n19342), .ZN(n16440) );
  AOI22_X1 U19616 ( .A1(n16434), .A2(n19315), .B1(n16433), .B2(n19339), .ZN(
        n16439) );
  OAI211_X1 U19617 ( .C1(n16437), .C2(n16436), .A(n19316), .B(n16435), .ZN(
        n16438) );
  NAND4_X1 U19618 ( .A1(n16441), .A2(n16440), .A3(n16439), .A4(n16438), .ZN(
        P2_U2827) );
  NAND2_X1 U19619 ( .A1(n16442), .A2(n19315), .ZN(n16446) );
  AOI22_X1 U19620 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19343), .ZN(n16443) );
  INV_X1 U19621 ( .A(n16443), .ZN(n16444) );
  AOI21_X1 U19622 ( .B1(n19342), .B2(P2_EBX_REG_26__SCAN_IN), .A(n16444), .ZN(
        n16445) );
  OAI211_X1 U19623 ( .C1(n16447), .C2(n19308), .A(n16446), .B(n16445), .ZN(
        n16448) );
  INV_X1 U19624 ( .A(n16448), .ZN(n16453) );
  OAI211_X1 U19625 ( .C1(n16451), .C2(n16450), .A(n19316), .B(n16449), .ZN(
        n16452) );
  OAI211_X1 U19626 ( .C1(n19323), .C2(n16454), .A(n16453), .B(n16452), .ZN(
        P2_U2829) );
  AOI22_X1 U19627 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n19351), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19343), .ZN(n16465) );
  INV_X1 U19628 ( .A(n16455), .ZN(n16456) );
  AOI22_X1 U19629 ( .A1(n16456), .A2(n19341), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n19342), .ZN(n16464) );
  AOI22_X1 U19630 ( .A1(n16458), .A2(n19315), .B1(n16457), .B2(n19339), .ZN(
        n16463) );
  OAI211_X1 U19631 ( .C1(n16461), .C2(n16460), .A(n19316), .B(n16459), .ZN(
        n16462) );
  NAND4_X1 U19632 ( .A1(n16465), .A2(n16464), .A3(n16463), .A4(n16462), .ZN(
        P2_U2831) );
  AOI22_X1 U19633 ( .A1(n16472), .A2(n16466), .B1(n19415), .B2(
        P2_EAX_REG_23__SCAN_IN), .ZN(n16471) );
  AOI22_X1 U19634 ( .A1(n19356), .A2(BUF1_REG_23__SCAN_IN), .B1(n19357), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16470) );
  INV_X1 U19635 ( .A(n16547), .ZN(n16467) );
  AOI22_X1 U19636 ( .A1(n16468), .A2(n19417), .B1(n19416), .B2(n16467), .ZN(
        n16469) );
  NAND3_X1 U19637 ( .A1(n16471), .A2(n16470), .A3(n16469), .ZN(P2_U2896) );
  AOI22_X1 U19638 ( .A1(n16472), .A2(n19384), .B1(n19415), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U19639 ( .A1(n19356), .A2(BUF1_REG_22__SCAN_IN), .B1(n19357), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16477) );
  INV_X1 U19640 ( .A(n16473), .ZN(n16474) );
  AOI22_X1 U19641 ( .A1(n16475), .A2(n19417), .B1(n19416), .B2(n16474), .ZN(
        n16476) );
  NAND3_X1 U19642 ( .A1(n16478), .A2(n16477), .A3(n16476), .ZN(P2_U2897) );
  AOI22_X1 U19643 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19461), .B1(n16530), 
        .B2(n16479), .ZN(n16486) );
  XOR2_X1 U19644 ( .A(n16480), .B(n16481), .Z(n16552) );
  INV_X1 U19645 ( .A(n16482), .ZN(n16483) );
  NAND2_X1 U19646 ( .A1(n16483), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16484) );
  AOI21_X1 U19647 ( .B1(n10715), .B2(n16484), .A(n15641), .ZN(n16550) );
  AOI222_X1 U19648 ( .A1(n16552), .A2(n16538), .B1(n19480), .B2(n16551), .C1(
        n19475), .C2(n16550), .ZN(n16485) );
  OAI211_X1 U19649 ( .C1(n16487), .C2(n16541), .A(n16486), .B(n16485), .ZN(
        P2_U2991) );
  AOI22_X1 U19650 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19473), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19326), .ZN(n16493) );
  OAI22_X1 U19651 ( .A1(n16489), .A2(n16514), .B1(n19464), .B2(n16488), .ZN(
        n16490) );
  AOI21_X1 U19652 ( .B1(n19480), .B2(n16491), .A(n16490), .ZN(n16492) );
  OAI211_X1 U19653 ( .C1(n19471), .C2(n16494), .A(n16493), .B(n16492), .ZN(
        P2_U2992) );
  AOI22_X1 U19654 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19461), .B1(n16530), 
        .B2(n16495), .ZN(n16510) );
  INV_X1 U19655 ( .A(n16496), .ZN(n16499) );
  NAND2_X1 U19656 ( .A1(n16497), .A2(n16594), .ZN(n16498) );
  NAND2_X1 U19657 ( .A1(n16499), .A2(n16498), .ZN(n16589) );
  NAND2_X1 U19658 ( .A1(n19480), .A2(n16500), .ZN(n16507) );
  NAND2_X1 U19659 ( .A1(n16501), .A2(n16502), .ZN(n16505) );
  NAND2_X1 U19660 ( .A1(n9830), .A2(n16503), .ZN(n16504) );
  XNOR2_X1 U19661 ( .A(n16505), .B(n16504), .ZN(n16591) );
  NAND2_X1 U19662 ( .A1(n16591), .A2(n16538), .ZN(n16506) );
  OAI211_X1 U19663 ( .C1(n16589), .C2(n19464), .A(n16507), .B(n16506), .ZN(
        n16508) );
  INV_X1 U19664 ( .A(n16508), .ZN(n16509) );
  OAI211_X1 U19665 ( .C1(n16511), .C2(n16541), .A(n16510), .B(n16509), .ZN(
        P2_U3003) );
  AOI22_X1 U19666 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19326), .B1(n16530), 
        .B2(n19275), .ZN(n16519) );
  NOR3_X1 U19667 ( .A1(n16513), .A2(n16512), .A3(n19464), .ZN(n16517) );
  OAI22_X1 U19668 ( .A1(n16515), .A2(n16514), .B1(n13256), .B2(n19279), .ZN(
        n16516) );
  NOR2_X1 U19669 ( .A1(n16517), .A2(n16516), .ZN(n16518) );
  OAI211_X1 U19670 ( .C1(n16520), .C2(n16541), .A(n16519), .B(n16518), .ZN(
        P2_U3005) );
  AOI22_X1 U19671 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19326), .B1(n16530), 
        .B2(n19295), .ZN(n16527) );
  NAND2_X1 U19672 ( .A1(n16521), .A2(n19475), .ZN(n16524) );
  NAND2_X1 U19673 ( .A1(n16522), .A2(n16538), .ZN(n16523) );
  OAI211_X1 U19674 ( .C1(n13256), .C2(n19299), .A(n16524), .B(n16523), .ZN(
        n16525) );
  INV_X1 U19675 ( .A(n16525), .ZN(n16526) );
  OAI211_X1 U19676 ( .C1(n16528), .C2(n16541), .A(n16527), .B(n16526), .ZN(
        P2_U3007) );
  AOI22_X1 U19677 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19461), .B1(n16530), 
        .B2(n16529), .ZN(n16540) );
  NAND2_X1 U19678 ( .A1(n16532), .A2(n16531), .ZN(n16534) );
  XNOR2_X1 U19679 ( .A(n16534), .B(n16533), .ZN(n16625) );
  INV_X1 U19680 ( .A(n16535), .ZN(n16623) );
  XOR2_X1 U19681 ( .A(n16537), .B(n16536), .Z(n16622) );
  AOI222_X1 U19682 ( .A1(n16625), .A2(n19475), .B1(n19480), .B2(n16623), .C1(
        n16538), .C2(n16622), .ZN(n16539) );
  OAI211_X1 U19683 ( .C1(n16542), .C2(n16541), .A(n16540), .B(n16539), .ZN(
        P2_U3009) );
  INV_X1 U19684 ( .A(n16543), .ZN(n16545) );
  AOI211_X1 U19685 ( .C1(n16546), .C2(n10715), .A(n16545), .B(n16544), .ZN(
        n16549) );
  OAI22_X1 U19686 ( .A1(n16547), .A2(n19487), .B1(n11157), .B2(n19304), .ZN(
        n16548) );
  NOR2_X1 U19687 ( .A1(n16549), .A2(n16548), .ZN(n16554) );
  AOI222_X1 U19688 ( .A1(n16552), .A2(n16639), .B1(n16635), .B2(n16551), .C1(
        n16624), .C2(n16550), .ZN(n16553) );
  OAI211_X1 U19689 ( .C1(n16555), .C2(n10715), .A(n16554), .B(n16553), .ZN(
        P2_U3023) );
  OAI21_X1 U19690 ( .B1(n16566), .B2(n16571), .A(n15742), .ZN(n16556) );
  AOI22_X1 U19691 ( .A1(n16557), .A2(n16556), .B1(n16621), .B2(n19366), .ZN(
        n16565) );
  NOR2_X1 U19692 ( .A1(n19491), .A2(n16558), .ZN(n16559) );
  AOI21_X1 U19693 ( .B1(n16560), .B2(n16624), .A(n16559), .ZN(n16563) );
  NAND2_X1 U19694 ( .A1(n16561), .A2(n16639), .ZN(n16562) );
  AND2_X1 U19695 ( .A1(n16563), .A2(n16562), .ZN(n16564) );
  OAI211_X1 U19696 ( .C1(n10891), .C2(n19304), .A(n16565), .B(n16564), .ZN(
        P2_U3033) );
  INV_X1 U19697 ( .A(n16566), .ZN(n16572) );
  NOR2_X1 U19698 ( .A1(n11097), .A2(n19304), .ZN(n16570) );
  OAI21_X1 U19699 ( .B1(n16567), .B2(n13536), .A(n13553), .ZN(n19369) );
  OAI22_X1 U19700 ( .A1(n16568), .A2(n16571), .B1(n19487), .B2(n19369), .ZN(
        n16569) );
  AOI211_X1 U19701 ( .C1(n16572), .C2(n16571), .A(n16570), .B(n16569), .ZN(
        n16576) );
  OAI22_X1 U19702 ( .A1(n16573), .A2(n19490), .B1(n19491), .B2(n19255), .ZN(
        n16574) );
  INV_X1 U19703 ( .A(n16574), .ZN(n16575) );
  OAI211_X1 U19704 ( .C1(n16577), .C2(n19500), .A(n16576), .B(n16575), .ZN(
        P2_U3034) );
  OAI21_X1 U19705 ( .B1(n16580), .B2(n16579), .A(n16578), .ZN(n16598) );
  NAND2_X1 U19706 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16581), .ZN(
        n16600) );
  AOI21_X1 U19707 ( .B1(n16599), .B2(n16594), .A(n16600), .ZN(n16584) );
  INV_X1 U19708 ( .A(n16582), .ZN(n16583) );
  AOI22_X1 U19709 ( .A1(n16584), .A2(n16583), .B1(n19326), .B2(
        P2_REIP_REG_11__SCAN_IN), .ZN(n16585) );
  OAI21_X1 U19710 ( .B1(n19487), .B2(n16586), .A(n16585), .ZN(n16587) );
  INV_X1 U19711 ( .A(n16587), .ZN(n16593) );
  OAI22_X1 U19712 ( .A1(n16589), .A2(n19490), .B1(n19491), .B2(n16588), .ZN(
        n16590) );
  AOI21_X1 U19713 ( .B1(n16639), .B2(n16591), .A(n16590), .ZN(n16592) );
  OAI211_X1 U19714 ( .C1(n16594), .C2(n16598), .A(n16593), .B(n16592), .ZN(
        P2_U3035) );
  XNOR2_X1 U19715 ( .A(n16596), .B(n16595), .ZN(n19375) );
  INV_X1 U19716 ( .A(n19375), .ZN(n19269) );
  NAND2_X1 U19717 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19326), .ZN(n16597) );
  OAI221_X1 U19718 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16600), 
        .C1(n16599), .C2(n16598), .A(n16597), .ZN(n16601) );
  AOI21_X1 U19719 ( .B1(n16621), .B2(n19269), .A(n16601), .ZN(n16605) );
  OAI22_X1 U19720 ( .A1(n16602), .A2(n19490), .B1(n19491), .B2(n19268), .ZN(
        n16603) );
  INV_X1 U19721 ( .A(n16603), .ZN(n16604) );
  OAI211_X1 U19722 ( .C1(n16606), .C2(n19500), .A(n16605), .B(n16604), .ZN(
        P2_U3036) );
  OAI21_X1 U19723 ( .B1(n16608), .B2(n16607), .A(n15973), .ZN(n19381) );
  NAND4_X1 U19724 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n16610), .A4(n16609), .ZN(
        n16612) );
  NAND2_X1 U19725 ( .A1(n19326), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n16611) );
  OAI211_X1 U19726 ( .C1(n19487), .C2(n19381), .A(n16612), .B(n16611), .ZN(
        n16613) );
  AOI221_X1 U19727 ( .B1(n16615), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(
        n16614), .C2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16613), .ZN(
        n16618) );
  AOI22_X1 U19728 ( .A1(n16616), .A2(n16624), .B1(n16635), .B2(n19290), .ZN(
        n16617) );
  OAI211_X1 U19729 ( .C1(n16619), .C2(n19500), .A(n16618), .B(n16617), .ZN(
        P2_U3038) );
  AOI22_X1 U19730 ( .A1(n19389), .A2(n16621), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n16620), .ZN(n16631) );
  AOI222_X1 U19731 ( .A1(n16625), .A2(n16624), .B1(n16635), .B2(n16623), .C1(
        n16639), .C2(n16622), .ZN(n16630) );
  NAND2_X1 U19732 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19326), .ZN(n16629) );
  OAI211_X1 U19733 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n16627), .B(n16626), .ZN(n16628) );
  NAND4_X1 U19734 ( .A1(n16631), .A2(n16630), .A3(n16629), .A4(n16628), .ZN(
        P2_U3041) );
  INV_X1 U19735 ( .A(n16632), .ZN(n16640) );
  OAI21_X1 U19736 ( .B1(n19487), .B2(n20135), .A(n16633), .ZN(n16634) );
  AOI21_X1 U19737 ( .B1(n13064), .B2(n16635), .A(n16634), .ZN(n16636) );
  OAI21_X1 U19738 ( .B1(n16637), .B2(n19490), .A(n16636), .ZN(n16638) );
  AOI21_X1 U19739 ( .B1(n16640), .B2(n16639), .A(n16638), .ZN(n16641) );
  OAI221_X1 U19740 ( .B1(n16643), .B2(n10522), .C1(n16643), .C2(n16642), .A(
        n16641), .ZN(P2_U3043) );
  NAND2_X1 U19741 ( .A1(n16644), .A2(n16646), .ZN(n16645) );
  OAI21_X1 U19742 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16646), .A(
        n16645), .ZN(n16679) );
  INV_X1 U19743 ( .A(n16646), .ZN(n16669) );
  NAND2_X1 U19744 ( .A1(n16669), .A2(n16647), .ZN(n16648) );
  OAI21_X1 U19745 ( .B1(n16649), .B2(n16669), .A(n16648), .ZN(n16678) );
  NAND2_X1 U19746 ( .A1(n9740), .A2(n16650), .ZN(n16655) );
  OAI21_X1 U19747 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16651), .ZN(n16654) );
  NAND2_X1 U19748 ( .A1(n16652), .A2(n19503), .ZN(n16653) );
  OAI211_X1 U19749 ( .C1(n16656), .C2(n16655), .A(n16654), .B(n16653), .ZN(
        n16662) );
  AOI22_X1 U19750 ( .A1(n16661), .A2(n16658), .B1(n11169), .B2(n16657), .ZN(
        n16659) );
  OAI21_X1 U19751 ( .B1(n16661), .B2(n16660), .A(n16659), .ZN(n20173) );
  AOI211_X1 U19752 ( .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16669), .A(
        n16662), .B(n20173), .ZN(n16677) );
  NOR2_X1 U19753 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n16678), .ZN(
        n16674) );
  INV_X1 U19754 ( .A(n16664), .ZN(n16668) );
  NOR2_X1 U19755 ( .A1(n16663), .A2(n20166), .ZN(n16665) );
  INV_X1 U19756 ( .A(n16665), .ZN(n16667) );
  AOI21_X1 U19757 ( .B1(n16665), .B2(n16664), .A(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16666) );
  AOI21_X1 U19758 ( .B1(n16668), .B2(n16667), .A(n16666), .ZN(n16670) );
  NOR2_X1 U19759 ( .A1(n16670), .A2(n16669), .ZN(n16671) );
  OAI21_X1 U19760 ( .B1(n16674), .B2(n20149), .A(n16671), .ZN(n16672) );
  AOI222_X1 U19761 ( .A1(n16679), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .B1(n16679), .B2(n16672), .C1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .C2(n16672), .ZN(n16675) );
  OAI221_X1 U19762 ( .B1(n16675), .B2(n16674), .C1(n16675), .C2(n20149), .A(
        n16673), .ZN(n16676) );
  OAI211_X1 U19763 ( .C1(n16679), .C2(n16678), .A(n16677), .B(n16676), .ZN(
        n16691) );
  AOI211_X1 U19764 ( .C1(n16682), .C2(n16691), .A(n16681), .B(n16680), .ZN(
        n16695) );
  NAND2_X1 U19765 ( .A1(n16684), .A2(n9740), .ZN(n16685) );
  OR2_X1 U19766 ( .A1(n16686), .A2(n16685), .ZN(n16687) );
  AND3_X1 U19767 ( .A1(n16687), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20187), 
        .ZN(n16689) );
  AOI22_X1 U19768 ( .A1(n20183), .A2(n16689), .B1(n20184), .B2(n16688), .ZN(
        n16693) );
  INV_X1 U19769 ( .A(n16689), .ZN(n16690) );
  AOI221_X1 U19770 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16691), .C1(
        P2_STATE2_REG_0__SCAN_IN), .C2(P2_STATE2_REG_1__SCAN_IN), .A(n16690), 
        .ZN(n20055) );
  NOR2_X1 U19771 ( .A1(n19151), .A2(n20055), .ZN(n16697) );
  INV_X1 U19772 ( .A(n16697), .ZN(n16692) );
  OAI21_X1 U19773 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16693), .A(n16692), 
        .ZN(n16694) );
  OAI211_X1 U19774 ( .C1(n20169), .C2(n16696), .A(n16695), .B(n16694), .ZN(
        P2_U3176) );
  OAI21_X1 U19775 ( .B1(n16697), .B2(n19670), .A(n16696), .ZN(P2_U3593) );
  INV_X1 U19776 ( .A(n16698), .ZN(n16707) );
  XNOR2_X1 U19777 ( .A(n9993), .B(n9834), .ZN(n16849) );
  OAI221_X1 U19778 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16701), .C1(
        n9993), .C2(n16700), .A(n16699), .ZN(n16702) );
  AOI21_X1 U19779 ( .B1(n17943), .B2(n16849), .A(n16702), .ZN(n16706) );
  OAI22_X1 U19780 ( .A1(n16709), .A2(n18167), .B1(n16712), .B2(n18079), .ZN(
        n16704) );
  AOI22_X1 U19781 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16704), .B1(
        n18076), .B2(n16703), .ZN(n16705) );
  OAI211_X1 U19782 ( .C1(n17814), .C2(n16707), .A(n16706), .B(n16705), .ZN(
        P3_U2800) );
  INV_X1 U19783 ( .A(n16708), .ZN(n16710) );
  AOI211_X1 U19784 ( .C1(n16710), .C2(n16713), .A(n16709), .B(n18167), .ZN(
        n16716) );
  INV_X1 U19785 ( .A(n16711), .ZN(n16714) );
  AOI211_X1 U19786 ( .C1(n16714), .C2(n16713), .A(n16712), .B(n18079), .ZN(
        n16715) );
  AOI211_X1 U19787 ( .C1(n18076), .C2(n16717), .A(n16716), .B(n16715), .ZN(
        n16723) );
  INV_X1 U19788 ( .A(n17944), .ZN(n17906) );
  AOI21_X1 U19789 ( .B1(n9992), .B2(n16835), .A(n9834), .ZN(n16859) );
  OAI21_X1 U19790 ( .B1(n17944), .B2(n17943), .A(n16859), .ZN(n16721) );
  OAI221_X1 U19791 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18862), .C1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16719), .A(n16718), .ZN(
        n16720) );
  NAND4_X1 U19792 ( .A1(n16723), .A2(n16722), .A3(n16721), .A4(n16720), .ZN(
        P3_U2801) );
  NOR3_X1 U19793 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16725) );
  NOR4_X1 U19794 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16724) );
  NAND4_X1 U19795 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16725), .A3(n16724), .A4(
        U215), .ZN(U213) );
  INV_X1 U19796 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19423) );
  INV_X2 U19797 ( .A(U214), .ZN(n16774) );
  NOR2_X2 U19798 ( .A1(n16774), .A2(n16726), .ZN(n16775) );
  OAI222_X1 U19799 ( .A1(U212), .A2(n19423), .B1(n16772), .B2(n16727), .C1(
        U214), .C2(n16807), .ZN(U216) );
  INV_X1 U19800 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U19801 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16770), .ZN(n16728) );
  OAI21_X1 U19802 ( .B1(n20719), .B2(n16772), .A(n16728), .ZN(U217) );
  INV_X1 U19803 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16730) );
  AOI22_X1 U19804 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16770), .ZN(n16729) );
  OAI21_X1 U19805 ( .B1(n16730), .B2(n16772), .A(n16729), .ZN(U218) );
  AOI222_X1 U19806 ( .A1(n16770), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(n16775), 
        .B2(BUF1_REG_28__SCAN_IN), .C1(n16774), .C2(P1_DATAO_REG_28__SCAN_IN), 
        .ZN(n16731) );
  INV_X1 U19807 ( .A(n16731), .ZN(U219) );
  INV_X1 U19808 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16733) );
  AOI22_X1 U19809 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16770), .ZN(n16732) );
  OAI21_X1 U19810 ( .B1(n16733), .B2(n16772), .A(n16732), .ZN(U220) );
  INV_X1 U19811 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U19812 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16770), .ZN(n16734) );
  OAI21_X1 U19813 ( .B1(n20881), .B2(n16772), .A(n16734), .ZN(U221) );
  INV_X1 U19814 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16736) );
  AOI22_X1 U19815 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16770), .ZN(n16735) );
  OAI21_X1 U19816 ( .B1(n16736), .B2(n16772), .A(n16735), .ZN(U222) );
  INV_X1 U19817 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16738) );
  AOI22_X1 U19818 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16770), .ZN(n16737) );
  OAI21_X1 U19819 ( .B1(n16738), .B2(n16772), .A(n16737), .ZN(U223) );
  INV_X1 U19820 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16740) );
  AOI22_X1 U19821 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16770), .ZN(n16739) );
  OAI21_X1 U19822 ( .B1(n16740), .B2(n16772), .A(n16739), .ZN(U224) );
  INV_X1 U19823 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U19824 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16774), .ZN(n16741) );
  OAI21_X1 U19825 ( .B1(n20912), .B2(U212), .A(n16741), .ZN(U225) );
  AOI22_X1 U19826 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16774), .ZN(n16742) );
  OAI21_X1 U19827 ( .B1(n16795), .B2(U212), .A(n16742), .ZN(U226) );
  AOI22_X1 U19828 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16770), .ZN(n16743) );
  OAI21_X1 U19829 ( .B1(n14094), .B2(n16772), .A(n16743), .ZN(U227) );
  AOI22_X1 U19830 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16770), .ZN(n16744) );
  OAI21_X1 U19831 ( .B1(n13985), .B2(n16772), .A(n16744), .ZN(U228) );
  INV_X1 U19832 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16746) );
  AOI22_X1 U19833 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16770), .ZN(n16745) );
  OAI21_X1 U19834 ( .B1(n16746), .B2(n16772), .A(n16745), .ZN(U229) );
  AOI22_X1 U19835 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16770), .ZN(n16747) );
  OAI21_X1 U19836 ( .B1(n13867), .B2(n16772), .A(n16747), .ZN(U230) );
  INV_X1 U19837 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16749) );
  AOI22_X1 U19838 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16770), .ZN(n16748) );
  OAI21_X1 U19839 ( .B1(n16749), .B2(n16772), .A(n16748), .ZN(U231) );
  INV_X1 U19840 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16751) );
  AOI22_X1 U19841 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16774), .ZN(n16750) );
  OAI21_X1 U19842 ( .B1(n16751), .B2(U212), .A(n16750), .ZN(U232) );
  INV_X1 U19843 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16753) );
  AOI22_X1 U19844 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16774), .ZN(n16752) );
  OAI21_X1 U19845 ( .B1(n16753), .B2(U212), .A(n16752), .ZN(U233) );
  INV_X1 U19846 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n20791) );
  INV_X1 U19847 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n20758) );
  OAI222_X1 U19848 ( .A1(U214), .A2(n20791), .B1(n16772), .B2(n16754), .C1(
        U212), .C2(n20758), .ZN(U234) );
  INV_X1 U19849 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n20769) );
  AOI22_X1 U19850 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16774), .ZN(n16755) );
  OAI21_X1 U19851 ( .B1(n20769), .B2(U212), .A(n16755), .ZN(U235) );
  INV_X1 U19852 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16787) );
  INV_X1 U19853 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n20733) );
  OAI222_X1 U19854 ( .A1(U212), .A2(n16787), .B1(n16772), .B2(n16756), .C1(
        U214), .C2(n20733), .ZN(U236) );
  INV_X1 U19855 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16758) );
  AOI22_X1 U19856 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16774), .ZN(n16757) );
  OAI21_X1 U19857 ( .B1(n16758), .B2(U212), .A(n16757), .ZN(U237) );
  AOI22_X1 U19858 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16770), .ZN(n16759) );
  OAI21_X1 U19859 ( .B1(n16760), .B2(n16772), .A(n16759), .ZN(U238) );
  INV_X1 U19860 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16762) );
  AOI22_X1 U19861 ( .A1(BUF1_REG_8__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16774), .ZN(n16761) );
  OAI21_X1 U19862 ( .B1(n16762), .B2(U212), .A(n16761), .ZN(U239) );
  AOI222_X1 U19863 ( .A1(n16770), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n16775), 
        .B2(BUF1_REG_7__SCAN_IN), .C1(n16774), .C2(P1_DATAO_REG_7__SCAN_IN), 
        .ZN(n16763) );
  INV_X1 U19864 ( .A(n16763), .ZN(U240) );
  AOI22_X1 U19865 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16770), .ZN(n16764) );
  OAI21_X1 U19866 ( .B1(n16765), .B2(n16772), .A(n16764), .ZN(U241) );
  INV_X1 U19867 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16781) );
  AOI22_X1 U19868 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16774), .ZN(n16766) );
  OAI21_X1 U19869 ( .B1(n16781), .B2(U212), .A(n16766), .ZN(U242) );
  INV_X1 U19870 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n20309) );
  AOI22_X1 U19871 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16775), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16770), .ZN(n16767) );
  OAI21_X1 U19872 ( .B1(n20309), .B2(U214), .A(n16767), .ZN(U243) );
  INV_X1 U19873 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16779) );
  AOI22_X1 U19874 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16774), .ZN(n16768) );
  OAI21_X1 U19875 ( .B1(n16779), .B2(U212), .A(n16768), .ZN(U244) );
  INV_X1 U19876 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16778) );
  AOI22_X1 U19877 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16774), .ZN(n16769) );
  OAI21_X1 U19878 ( .B1(n16778), .B2(U212), .A(n16769), .ZN(U245) );
  INV_X1 U19879 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16773) );
  AOI22_X1 U19880 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16774), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16770), .ZN(n16771) );
  OAI21_X1 U19881 ( .B1(n16773), .B2(n16772), .A(n16771), .ZN(U246) );
  INV_X1 U19882 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n20870) );
  AOI22_X1 U19883 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16775), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16774), .ZN(n16776) );
  OAI21_X1 U19884 ( .B1(n20870), .B2(U212), .A(n16776), .ZN(U247) );
  AOI22_X1 U19885 ( .A1(n16804), .A2(n20870), .B1(n18478), .B2(U215), .ZN(U251) );
  OAI22_X1 U19886 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16804), .ZN(n16777) );
  INV_X1 U19887 ( .A(n16777), .ZN(U252) );
  INV_X1 U19888 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18490) );
  AOI22_X1 U19889 ( .A1(n16804), .A2(n16778), .B1(n18490), .B2(U215), .ZN(U253) );
  INV_X1 U19890 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18495) );
  AOI22_X1 U19891 ( .A1(n16804), .A2(n16779), .B1(n18495), .B2(U215), .ZN(U254) );
  OAI22_X1 U19892 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16804), .ZN(n16780) );
  INV_X1 U19893 ( .A(n16780), .ZN(U255) );
  INV_X1 U19894 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18505) );
  AOI22_X1 U19895 ( .A1(n16804), .A2(n16781), .B1(n18505), .B2(U215), .ZN(U256) );
  OAI22_X1 U19896 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16804), .ZN(n16782) );
  INV_X1 U19897 ( .A(n16782), .ZN(U257) );
  INV_X1 U19898 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16783) );
  INV_X1 U19899 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18513) );
  AOI22_X1 U19900 ( .A1(n16806), .A2(n16783), .B1(n18513), .B2(U215), .ZN(U258) );
  OAI22_X1 U19901 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16806), .ZN(n16784) );
  INV_X1 U19902 ( .A(n16784), .ZN(U259) );
  OAI22_X1 U19903 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16806), .ZN(n16785) );
  INV_X1 U19904 ( .A(n16785), .ZN(U260) );
  OAI22_X1 U19905 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16806), .ZN(n16786) );
  INV_X1 U19906 ( .A(n16786), .ZN(U261) );
  INV_X1 U19907 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17776) );
  AOI22_X1 U19908 ( .A1(n16804), .A2(n16787), .B1(n17776), .B2(U215), .ZN(U262) );
  INV_X1 U19909 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17778) );
  AOI22_X1 U19910 ( .A1(n16806), .A2(n20769), .B1(n17778), .B2(U215), .ZN(U263) );
  INV_X1 U19911 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17782) );
  AOI22_X1 U19912 ( .A1(n16804), .A2(n20758), .B1(n17782), .B2(U215), .ZN(U264) );
  OAI22_X1 U19913 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16806), .ZN(n16788) );
  INV_X1 U19914 ( .A(n16788), .ZN(U265) );
  OAI22_X1 U19915 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16806), .ZN(n16789) );
  INV_X1 U19916 ( .A(n16789), .ZN(U266) );
  OAI22_X1 U19917 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16804), .ZN(n16790) );
  INV_X1 U19918 ( .A(n16790), .ZN(U267) );
  OAI22_X1 U19919 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16806), .ZN(n16791) );
  INV_X1 U19920 ( .A(n16791), .ZN(U268) );
  OAI22_X1 U19921 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16804), .ZN(n16792) );
  INV_X1 U19922 ( .A(n16792), .ZN(U269) );
  OAI22_X1 U19923 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16804), .ZN(n16793) );
  INV_X1 U19924 ( .A(n16793), .ZN(U270) );
  OAI22_X1 U19925 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16804), .ZN(n16794) );
  INV_X1 U19926 ( .A(n16794), .ZN(U271) );
  AOI22_X1 U19927 ( .A1(n16804), .A2(n16795), .B1(n15580), .B2(U215), .ZN(U272) );
  INV_X1 U19928 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n16796) );
  AOI22_X1 U19929 ( .A1(n16806), .A2(n20912), .B1(n16796), .B2(U215), .ZN(U273) );
  OAI22_X1 U19930 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16804), .ZN(n16797) );
  INV_X1 U19931 ( .A(n16797), .ZN(U274) );
  OAI22_X1 U19932 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16804), .ZN(n16798) );
  INV_X1 U19933 ( .A(n16798), .ZN(U275) );
  OAI22_X1 U19934 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16804), .ZN(n16799) );
  INV_X1 U19935 ( .A(n16799), .ZN(U276) );
  OAI22_X1 U19936 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16804), .ZN(n16800) );
  INV_X1 U19937 ( .A(n16800), .ZN(U277) );
  OAI22_X1 U19938 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16804), .ZN(n16801) );
  INV_X1 U19939 ( .A(n16801), .ZN(U278) );
  INV_X1 U19940 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n16802) );
  INV_X1 U19941 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18499) );
  AOI22_X1 U19942 ( .A1(n16804), .A2(n16802), .B1(n18499), .B2(U215), .ZN(U279) );
  OAI22_X1 U19943 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16804), .ZN(n16803) );
  INV_X1 U19944 ( .A(n16803), .ZN(U280) );
  OAI22_X1 U19945 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16804), .ZN(n16805) );
  INV_X1 U19946 ( .A(n16805), .ZN(U281) );
  INV_X1 U19947 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U19948 ( .A1(n16806), .A2(n19423), .B1(n17532), .B2(U215), .ZN(U282) );
  INV_X1 U19949 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17679) );
  AOI222_X1 U19950 ( .A1(n16807), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19423), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17679), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16808) );
  INV_X1 U19951 ( .A(n16810), .ZN(n16809) );
  INV_X1 U19952 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19031) );
  INV_X1 U19953 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20090) );
  AOI22_X1 U19954 ( .A1(n16809), .A2(n19031), .B1(n20090), .B2(n16810), .ZN(
        U347) );
  INV_X1 U19955 ( .A(n16810), .ZN(n16811) );
  INV_X1 U19956 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19030) );
  INV_X1 U19957 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20089) );
  AOI22_X1 U19958 ( .A1(n16811), .A2(n19030), .B1(n20089), .B2(n16810), .ZN(
        U348) );
  INV_X1 U19959 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19027) );
  INV_X1 U19960 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20088) );
  AOI22_X1 U19961 ( .A1(n16809), .A2(n19027), .B1(n20088), .B2(n16810), .ZN(
        U349) );
  INV_X1 U19962 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19026) );
  INV_X1 U19963 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20087) );
  AOI22_X1 U19964 ( .A1(n16809), .A2(n19026), .B1(n20087), .B2(n16810), .ZN(
        U350) );
  INV_X1 U19965 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19024) );
  INV_X1 U19966 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20086) );
  AOI22_X1 U19967 ( .A1(n16809), .A2(n19024), .B1(n20086), .B2(n16810), .ZN(
        U351) );
  INV_X1 U19968 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19021) );
  INV_X1 U19969 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20085) );
  AOI22_X1 U19970 ( .A1(n16809), .A2(n19021), .B1(n20085), .B2(n16810), .ZN(
        U352) );
  INV_X1 U19971 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19020) );
  INV_X1 U19972 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U19973 ( .A1(n16811), .A2(n19020), .B1(n20084), .B2(n16810), .ZN(
        U353) );
  INV_X1 U19974 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19018) );
  AOI22_X1 U19975 ( .A1(n16809), .A2(n19018), .B1(n20083), .B2(n16810), .ZN(
        U354) );
  INV_X1 U19976 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19070) );
  INV_X1 U19977 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20120) );
  AOI22_X1 U19978 ( .A1(n16809), .A2(n19070), .B1(n20120), .B2(n16810), .ZN(
        U355) );
  INV_X1 U19979 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19066) );
  INV_X1 U19980 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20117) );
  AOI22_X1 U19981 ( .A1(n16809), .A2(n19066), .B1(n20117), .B2(n16810), .ZN(
        U356) );
  INV_X1 U19982 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19064) );
  INV_X1 U19983 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U19984 ( .A1(n16809), .A2(n19064), .B1(n20114), .B2(n16810), .ZN(
        U357) );
  INV_X1 U19985 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19061) );
  INV_X1 U19986 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U19987 ( .A1(n16809), .A2(n19061), .B1(n20901), .B2(n16810), .ZN(
        U358) );
  INV_X1 U19988 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20940) );
  INV_X1 U19989 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20112) );
  AOI22_X1 U19990 ( .A1(n16809), .A2(n20940), .B1(n20112), .B2(n16810), .ZN(
        U359) );
  INV_X1 U19991 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19059) );
  INV_X1 U19992 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U19993 ( .A1(n16809), .A2(n19059), .B1(n20110), .B2(n16810), .ZN(
        U360) );
  INV_X1 U19994 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19057) );
  INV_X1 U19995 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20842) );
  AOI22_X1 U19996 ( .A1(n16809), .A2(n19057), .B1(n20842), .B2(n16810), .ZN(
        U361) );
  INV_X1 U19997 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n20738) );
  INV_X1 U19998 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U19999 ( .A1(n16809), .A2(n20738), .B1(n20108), .B2(n16810), .ZN(
        U362) );
  INV_X1 U20000 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19054) );
  INV_X1 U20001 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U20002 ( .A1(n16809), .A2(n19054), .B1(n20107), .B2(n16810), .ZN(
        U363) );
  INV_X1 U20003 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19052) );
  INV_X1 U20004 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20105) );
  AOI22_X1 U20005 ( .A1(n16809), .A2(n19052), .B1(n20105), .B2(n16810), .ZN(
        U364) );
  INV_X1 U20006 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19017) );
  INV_X1 U20007 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20081) );
  AOI22_X1 U20008 ( .A1(n16809), .A2(n19017), .B1(n20081), .B2(n16810), .ZN(
        U365) );
  INV_X1 U20009 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19050) );
  INV_X1 U20010 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20104) );
  AOI22_X1 U20011 ( .A1(n16809), .A2(n19050), .B1(n20104), .B2(n16810), .ZN(
        U366) );
  INV_X1 U20012 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19048) );
  INV_X1 U20013 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20102) );
  AOI22_X1 U20014 ( .A1(n16809), .A2(n19048), .B1(n20102), .B2(n16810), .ZN(
        U367) );
  INV_X1 U20015 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19046) );
  INV_X1 U20016 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20100) );
  AOI22_X1 U20017 ( .A1(n16809), .A2(n19046), .B1(n20100), .B2(n16810), .ZN(
        U368) );
  INV_X1 U20018 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19043) );
  INV_X1 U20019 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20098) );
  AOI22_X1 U20020 ( .A1(n16809), .A2(n19043), .B1(n20098), .B2(n16810), .ZN(
        U369) );
  INV_X1 U20021 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19042) );
  INV_X1 U20022 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20096) );
  AOI22_X1 U20023 ( .A1(n16809), .A2(n19042), .B1(n20096), .B2(n16810), .ZN(
        U370) );
  INV_X1 U20024 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19040) );
  INV_X1 U20025 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20095) );
  AOI22_X1 U20026 ( .A1(n16811), .A2(n19040), .B1(n20095), .B2(n16810), .ZN(
        U371) );
  INV_X1 U20027 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20753) );
  INV_X1 U20028 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20094) );
  AOI22_X1 U20029 ( .A1(n16811), .A2(n20753), .B1(n20094), .B2(n16810), .ZN(
        U372) );
  INV_X1 U20030 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19037) );
  INV_X1 U20031 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20093) );
  AOI22_X1 U20032 ( .A1(n16811), .A2(n19037), .B1(n20093), .B2(n16810), .ZN(
        U373) );
  INV_X1 U20033 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19035) );
  INV_X1 U20034 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20092) );
  AOI22_X1 U20035 ( .A1(n16811), .A2(n19035), .B1(n20092), .B2(n16810), .ZN(
        U374) );
  INV_X1 U20036 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19033) );
  INV_X1 U20037 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20091) );
  AOI22_X1 U20038 ( .A1(n16811), .A2(n19033), .B1(n20091), .B2(n16810), .ZN(
        U375) );
  INV_X1 U20039 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19015) );
  INV_X1 U20040 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20080) );
  AOI22_X1 U20041 ( .A1(n16811), .A2(n19015), .B1(n20080), .B2(n16810), .ZN(
        U376) );
  INV_X1 U20042 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19014) );
  NAND2_X1 U20043 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19014), .ZN(n19001) );
  AOI22_X1 U20044 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19001), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19012), .ZN(n19076) );
  AOI21_X1 U20045 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19076), .ZN(n16812) );
  INV_X1 U20046 ( .A(n16812), .ZN(P3_U2633) );
  NAND2_X1 U20047 ( .A1(n19079), .A2(n19143), .ZN(n16814) );
  OAI21_X1 U20048 ( .B1(n16818), .B2(n17727), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16813) );
  OAI21_X1 U20049 ( .B1(n16814), .B2(n18989), .A(n16813), .ZN(P3_U2634) );
  AOI21_X1 U20050 ( .B1(n19012), .B2(n19014), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16815) );
  AOI22_X1 U20051 ( .A1(n19069), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16815), 
        .B2(n19141), .ZN(P3_U2635) );
  NOR2_X1 U20052 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18997) );
  OAI21_X1 U20053 ( .B1(n18997), .B2(BS16), .A(n19076), .ZN(n19074) );
  OAI21_X1 U20054 ( .B1(n19076), .B2(n19131), .A(n19074), .ZN(P3_U2636) );
  NOR3_X1 U20055 ( .A1(n16818), .A2(n16817), .A3(n16816), .ZN(n18967) );
  NOR2_X1 U20056 ( .A1(n18967), .A2(n18983), .ZN(n19122) );
  OAI21_X1 U20057 ( .B1(n19122), .B2(n18466), .A(n16819), .ZN(P3_U2637) );
  INV_X1 U20058 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19121) );
  NOR4_X1 U20059 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_10__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n16829) );
  NOR4_X1 U20060 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_6__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_8__SCAN_IN), .ZN(n16828) );
  NOR2_X1 U20061 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n20974) );
  AOI211_X1 U20062 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_3__SCAN_IN), .B(
        P3_DATAWIDTH_REG_4__SCAN_IN), .ZN(n16820) );
  NAND2_X1 U20063 ( .A1(n20974), .A2(n16820), .ZN(n16826) );
  NOR4_X1 U20064 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16824) );
  NOR4_X1 U20065 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_15__SCAN_IN), .A3(P3_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_17__SCAN_IN), .ZN(n16823) );
  NOR4_X1 U20066 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16822) );
  NOR4_X1 U20067 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16821) );
  NAND4_X1 U20068 ( .A1(n16824), .A2(n16823), .A3(n16822), .A4(n16821), .ZN(
        n16825) );
  NOR4_X1 U20069 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_2__SCAN_IN), .A3(n16826), .A4(n16825), .ZN(n16827) );
  NAND3_X1 U20070 ( .A1(n16829), .A2(n16828), .A3(n16827), .ZN(n19120) );
  INV_X1 U20071 ( .A(n19120), .ZN(n19118) );
  INV_X1 U20072 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n20771) );
  NAND2_X1 U20073 ( .A1(n19118), .A2(n20771), .ZN(n19117) );
  NOR3_X1 U20074 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(n19117), .ZN(n16831) );
  AOI21_X1 U20075 ( .B1(P3_BYTEENABLE_REG_1__SCAN_IN), .B2(n19120), .A(n16831), 
        .ZN(n16830) );
  OAI21_X1 U20076 ( .B1(n19121), .B2(n19120), .A(n16830), .ZN(P3_U2638) );
  NAND2_X1 U20077 ( .A1(n19118), .A2(n19121), .ZN(n19111) );
  AOI21_X1 U20078 ( .B1(P3_BYTEENABLE_REG_3__SCAN_IN), .B2(n19120), .A(n16831), 
        .ZN(n16832) );
  OAI21_X1 U20079 ( .B1(P3_DATAWIDTH_REG_1__SCAN_IN), .B2(n19111), .A(n16832), 
        .ZN(P3_U2639) );
  INV_X1 U20080 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19068) );
  NAND4_X1 U20081 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16877), .ZN(n16841) );
  NOR3_X1 U20082 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19068), .A3(n16841), 
        .ZN(n16834) );
  AOI21_X1 U20083 ( .B1(n17197), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16834), .ZN(
        n16845) );
  NAND2_X1 U20084 ( .A1(n16886), .A2(n16885), .ZN(n16884) );
  NOR2_X1 U20085 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16884), .ZN(n16867) );
  INV_X1 U20086 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16856) );
  NAND2_X1 U20087 ( .A1(n16867), .A2(n16856), .ZN(n16847) );
  NOR2_X1 U20088 ( .A1(n17165), .A2(n16847), .ZN(n16853) );
  INV_X1 U20089 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17208) );
  OAI21_X1 U20090 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16836), .A(
        n16835), .ZN(n17800) );
  INV_X1 U20091 ( .A(n17800), .ZN(n16870) );
  OAI21_X1 U20092 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n16838), .A(
        n16837), .ZN(n17809) );
  INV_X1 U20093 ( .A(n17809), .ZN(n16880) );
  NOR2_X1 U20094 ( .A1(n16839), .A2(n9816), .ZN(n16879) );
  NOR2_X1 U20095 ( .A1(n16880), .A2(n16879), .ZN(n16878) );
  NOR2_X1 U20096 ( .A1(n16878), .A2(n9816), .ZN(n16869) );
  NOR2_X1 U20097 ( .A1(n16870), .A2(n16869), .ZN(n16868) );
  NOR2_X1 U20098 ( .A1(n16868), .A2(n9816), .ZN(n16858) );
  NAND2_X1 U20099 ( .A1(n17171), .A2(n17184), .ZN(n17101) );
  NAND3_X1 U20100 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16840) );
  INV_X1 U20101 ( .A(n16957), .ZN(n17198) );
  AOI21_X1 U20102 ( .B1(n16840), .B2(n17198), .A(n16883), .ZN(n16860) );
  NOR2_X1 U20103 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16841), .ZN(n16851) );
  INV_X1 U20104 ( .A(n16851), .ZN(n16842) );
  AOI21_X1 U20105 ( .B1(n16860), .B2(n16842), .A(n19071), .ZN(n16843) );
  OAI211_X1 U20106 ( .C1(n16846), .C2(n17181), .A(n16845), .B(n16844), .ZN(
        P3_U2640) );
  NAND2_X1 U20107 ( .A1(n17196), .A2(n16847), .ZN(n16865) );
  XOR2_X1 U20108 ( .A(n16849), .B(n16848), .Z(n16852) );
  OAI22_X1 U20109 ( .A1(n16860), .A2(n19068), .B1(n9993), .B2(n17181), .ZN(
        n16850) );
  AOI211_X1 U20110 ( .C1(n16852), .C2(n17184), .A(n16851), .B(n16850), .ZN(
        n16855) );
  OAI21_X1 U20111 ( .B1(n17197), .B2(n16853), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16854) );
  OAI211_X1 U20112 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16865), .A(n16855), .B(
        n16854), .ZN(P3_U2641) );
  NOR2_X1 U20113 ( .A1(n16867), .A2(n16856), .ZN(n16866) );
  AOI211_X1 U20114 ( .C1(n16859), .C2(n16858), .A(n16857), .B(n18992), .ZN(
        n16862) );
  INV_X1 U20115 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19065) );
  OAI22_X1 U20116 ( .A1(n16860), .A2(n19065), .B1(n9992), .B2(n17181), .ZN(
        n16861) );
  AOI211_X1 U20117 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17197), .A(n16862), .B(
        n16861), .ZN(n16864) );
  NAND4_X1 U20118 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16877), .A4(n19065), .ZN(n16863) );
  OAI211_X1 U20119 ( .C1(n16866), .C2(n16865), .A(n16864), .B(n16863), .ZN(
        P3_U2642) );
  INV_X1 U20120 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16876) );
  AOI22_X1 U20121 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16883), .B1(n17197), 
        .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16875) );
  INV_X1 U20122 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19062) );
  INV_X1 U20123 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19063) );
  AOI22_X1 U20124 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .B1(n19062), .B2(n19063), .ZN(n16873) );
  AOI211_X1 U20125 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16884), .A(n16867), .B(
        n17165), .ZN(n16872) );
  AOI211_X1 U20126 ( .C1(n16870), .C2(n16869), .A(n16868), .B(n18992), .ZN(
        n16871) );
  AOI211_X1 U20127 ( .C1(n16877), .C2(n16873), .A(n16872), .B(n16871), .ZN(
        n16874) );
  OAI211_X1 U20128 ( .C1(n16876), .C2(n17181), .A(n16875), .B(n16874), .ZN(
        P3_U2643) );
  INV_X1 U20129 ( .A(n16877), .ZN(n16889) );
  AOI211_X1 U20130 ( .C1(n16880), .C2(n16879), .A(n16878), .B(n18992), .ZN(
        n16882) );
  INV_X1 U20131 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17812) );
  OAI22_X1 U20132 ( .A1(n17812), .A2(n17181), .B1(n17163), .B2(n16885), .ZN(
        n16881) );
  AOI211_X1 U20133 ( .C1(n16883), .C2(P3_REIP_REG_27__SCAN_IN), .A(n16882), 
        .B(n16881), .ZN(n16888) );
  OAI211_X1 U20134 ( .C1(n16886), .C2(n16885), .A(n17196), .B(n16884), .ZN(
        n16887) );
  OAI211_X1 U20135 ( .C1(P3_REIP_REG_27__SCAN_IN), .C2(n16889), .A(n16888), 
        .B(n16887), .ZN(P3_U2644) );
  INV_X1 U20136 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19056) );
  OAI21_X1 U20137 ( .B1(n16912), .B2(n17173), .A(n17199), .ZN(n16917) );
  AOI21_X1 U20138 ( .B1(n17178), .B2(n19056), .A(n16917), .ZN(n16900) );
  INV_X1 U20139 ( .A(n16890), .ZN(n16893) );
  NAND2_X1 U20140 ( .A1(n16893), .A2(n17196), .ZN(n16903) );
  OAI22_X1 U20141 ( .A1(n17840), .A2(n17181), .B1(n16903), .B2(
        P3_EBX_REG_25__SCAN_IN), .ZN(n16891) );
  INV_X1 U20142 ( .A(n16891), .ZN(n16899) );
  AOI221_X1 U20143 ( .B1(n17165), .B2(n17163), .C1(n16893), .C2(n17163), .A(
        n16892), .ZN(n16896) );
  AOI211_X1 U20144 ( .C1(n17842), .C2(n9773), .A(n16894), .B(n18992), .ZN(
        n16895) );
  AOI211_X1 U20145 ( .C1(n16897), .C2(n19058), .A(n16896), .B(n16895), .ZN(
        n16898) );
  OAI211_X1 U20146 ( .C1(n16900), .C2(n19058), .A(n16899), .B(n16898), .ZN(
        P3_U2646) );
  INV_X1 U20147 ( .A(n16917), .ZN(n16909) );
  AOI22_X1 U20148 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17182), .B1(
        n17197), .B2(P3_EBX_REG_24__SCAN_IN), .ZN(n16908) );
  NOR2_X1 U20149 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17173), .ZN(n16906) );
  AOI211_X1 U20150 ( .C1(n17853), .C2(n16902), .A(n16901), .B(n18992), .ZN(
        n16905) );
  AOI21_X1 U20151 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16918), .A(n16903), .ZN(
        n16904) );
  AOI211_X1 U20152 ( .C1(n16906), .C2(n16912), .A(n16905), .B(n16904), .ZN(
        n16907) );
  OAI211_X1 U20153 ( .C1(n16909), .C2(n19056), .A(n16908), .B(n16907), .ZN(
        P3_U2647) );
  AOI211_X1 U20154 ( .C1(n17874), .C2(n16911), .A(n16910), .B(n18992), .ZN(
        n16916) );
  OR2_X1 U20155 ( .A1(n17173), .A2(n16912), .ZN(n16913) );
  OAI22_X1 U20156 ( .A1(n17836), .A2(n17181), .B1(n16914), .B2(n16913), .ZN(
        n16915) );
  AOI211_X1 U20157 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16917), .A(n16916), 
        .B(n16915), .ZN(n16920) );
  OAI211_X1 U20158 ( .C1(n16925), .C2(n16921), .A(n17196), .B(n16918), .ZN(
        n16919) );
  OAI211_X1 U20159 ( .C1(n16921), .C2(n17163), .A(n16920), .B(n16919), .ZN(
        P3_U2648) );
  INV_X1 U20160 ( .A(n16922), .ZN(n16926) );
  AOI21_X1 U20161 ( .B1(n17178), .B2(n16926), .A(n17185), .ZN(n16934) );
  INV_X1 U20162 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19053) );
  AOI22_X1 U20163 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17182), .B1(
        n17197), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16931) );
  AOI211_X1 U20164 ( .C1(n17881), .C2(n16924), .A(n16923), .B(n18992), .ZN(
        n16929) );
  AOI211_X1 U20165 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16938), .A(n16925), .B(
        n17165), .ZN(n16928) );
  NOR3_X1 U20166 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n17173), .A3(n16926), 
        .ZN(n16927) );
  NOR3_X1 U20167 ( .A1(n16929), .A2(n16928), .A3(n16927), .ZN(n16930) );
  OAI211_X1 U20168 ( .C1(n16934), .C2(n19053), .A(n16931), .B(n16930), .ZN(
        P3_U2649) );
  AOI211_X1 U20169 ( .C1(n17894), .C2(n16933), .A(n16932), .B(n18992), .ZN(
        n16937) );
  INV_X1 U20170 ( .A(n17010), .ZN(n16985) );
  NAND2_X1 U20171 ( .A1(n17178), .A2(n16985), .ZN(n16999) );
  NOR2_X1 U20172 ( .A1(n16944), .A2(n16999), .ZN(n16959) );
  INV_X1 U20173 ( .A(n16959), .ZN(n16974) );
  AOI221_X1 U20174 ( .B1(n16935), .B2(n19051), .C1(n16974), .C2(n19051), .A(
        n16934), .ZN(n16936) );
  AOI211_X1 U20175 ( .C1(P3_EBX_REG_21__SCAN_IN), .C2(n17197), .A(n16937), .B(
        n16936), .ZN(n16940) );
  OAI211_X1 U20176 ( .C1(n16941), .C2(n17292), .A(n17196), .B(n16938), .ZN(
        n16939) );
  OAI211_X1 U20177 ( .C1(n17181), .C2(n17898), .A(n16940), .B(n16939), .ZN(
        P3_U2650) );
  INV_X1 U20178 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19049) );
  INV_X1 U20179 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19047) );
  INV_X1 U20180 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19045) );
  NOR2_X1 U20181 ( .A1(n19047), .A2(n19045), .ZN(n16945) );
  AND3_X1 U20182 ( .A1(n19049), .A2(n16945), .A3(n16959), .ZN(n16943) );
  AOI211_X1 U20183 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16960), .A(n16941), .B(
        n17165), .ZN(n16942) );
  AOI211_X1 U20184 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17197), .A(n16943), .B(
        n16942), .ZN(n16951) );
  NOR3_X1 U20185 ( .A1(n17185), .A2(n16944), .A3(n17010), .ZN(n16956) );
  AOI211_X1 U20186 ( .C1(n16945), .C2(n16956), .A(n16957), .B(n19049), .ZN(
        n16949) );
  AOI211_X1 U20187 ( .C1(n17911), .C2(n16947), .A(n16946), .B(n18992), .ZN(
        n16948) );
  AOI211_X1 U20188 ( .C1(n17182), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16949), .B(n16948), .ZN(n16950) );
  NAND2_X1 U20189 ( .A1(n16951), .A2(n16950), .ZN(P3_U2651) );
  AOI22_X1 U20190 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17182), .B1(
        n17197), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16964) );
  INV_X1 U20191 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17934) );
  NOR2_X1 U20192 ( .A1(n17934), .A2(n16953), .ZN(n16952) );
  OAI21_X1 U20193 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16952), .A(
        n17880), .ZN(n17921) );
  AOI22_X1 U20194 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16953), .B1(
        n17917), .B2(n17934), .ZN(n17931) );
  AOI21_X1 U20195 ( .B1(n16966), .B2(n17931), .A(n9816), .ZN(n16954) );
  XNOR2_X1 U20196 ( .A(n17921), .B(n16954), .ZN(n16955) );
  AOI21_X1 U20197 ( .B1(n16955), .B2(n17184), .A(n9731), .ZN(n16963) );
  NOR2_X1 U20198 ( .A1(n16957), .A2(n16956), .ZN(n16977) );
  XOR2_X1 U20199 ( .A(n19047), .B(n19045), .Z(n16958) );
  AOI22_X1 U20200 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16977), .B1(n16959), 
        .B2(n16958), .ZN(n16962) );
  OAI211_X1 U20201 ( .C1(n16965), .C2(n17319), .A(n17196), .B(n16960), .ZN(
        n16961) );
  NAND4_X1 U20202 ( .A1(n16964), .A2(n16963), .A3(n16962), .A4(n16961), .ZN(
        P3_U2652) );
  INV_X1 U20203 ( .A(n16977), .ZN(n16973) );
  AOI211_X1 U20204 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16981), .A(n16965), .B(
        n17165), .ZN(n16971) );
  INV_X1 U20205 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17332) );
  OR2_X1 U20206 ( .A1(n16966), .A2(n9816), .ZN(n16968) );
  OAI21_X1 U20207 ( .B1(n16966), .B2(n9816), .A(n17931), .ZN(n16967) );
  OAI211_X1 U20208 ( .C1(n17931), .C2(n16968), .A(n17184), .B(n16967), .ZN(
        n16969) );
  OAI211_X1 U20209 ( .C1(n17163), .C2(n17332), .A(n18455), .B(n16969), .ZN(
        n16970) );
  AOI211_X1 U20210 ( .C1(n17182), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16971), .B(n16970), .ZN(n16972) );
  OAI221_X1 U20211 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n16974), .C1(n19045), 
        .C2(n16973), .A(n16972), .ZN(P3_U2653) );
  INV_X1 U20212 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19041) );
  INV_X1 U20213 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19039) );
  NOR4_X1 U20214 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n19041), .A3(n19039), 
        .A4(n16999), .ZN(n16976) );
  OAI22_X1 U20215 ( .A1(n9984), .A2(n17181), .B1(n17163), .B2(n17348), .ZN(
        n16975) );
  AOI211_X1 U20216 ( .C1(n16977), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16976), 
        .B(n16975), .ZN(n16984) );
  NAND2_X1 U20217 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9845), .ZN(
        n16988) );
  AOI21_X1 U20218 ( .B1(n9984), .B2(n16988), .A(n17917), .ZN(n17945) );
  AOI21_X1 U20219 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16978), .A(
        n9816), .ZN(n16980) );
  AOI21_X1 U20220 ( .B1(n17945), .B2(n16980), .A(n18992), .ZN(n16979) );
  OAI21_X1 U20221 ( .B1(n17945), .B2(n16980), .A(n16979), .ZN(n16983) );
  OAI211_X1 U20222 ( .C1(n16987), .C2(n17348), .A(n17196), .B(n16981), .ZN(
        n16982) );
  NAND4_X1 U20223 ( .A1(n16984), .A2(n18455), .A3(n16983), .A4(n16982), .ZN(
        P3_U2654) );
  NAND2_X1 U20224 ( .A1(n16985), .A2(n17199), .ZN(n16986) );
  OAI21_X1 U20225 ( .B1(n19039), .B2(n16986), .A(n17198), .ZN(n16998) );
  AOI22_X1 U20226 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17182), .B1(
        n17197), .B2(P3_EBX_REG_16__SCAN_IN), .ZN(n16997) );
  NOR3_X1 U20227 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n19039), .A3(n16999), 
        .ZN(n16995) );
  AOI211_X1 U20228 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17006), .A(n16987), .B(
        n17165), .ZN(n16994) );
  INV_X1 U20229 ( .A(n17000), .ZN(n16989) );
  OAI21_X1 U20230 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16989), .A(
        n16988), .ZN(n17963) );
  INV_X1 U20231 ( .A(n17963), .ZN(n16992) );
  NAND2_X1 U20232 ( .A1(n17001), .A2(n17171), .ZN(n16990) );
  INV_X1 U20233 ( .A(n16990), .ZN(n16991) );
  AOI221_X1 U20234 ( .B1(n16992), .B2(n16991), .C1(n17963), .C2(n16990), .A(
        n18992), .ZN(n16993) );
  NOR4_X1 U20235 ( .A1(n9731), .A2(n16995), .A3(n16994), .A4(n16993), .ZN(
        n16996) );
  OAI211_X1 U20236 ( .C1(n16998), .C2(n19041), .A(n16997), .B(n16996), .ZN(
        P3_U2655) );
  AOI21_X1 U20237 ( .B1(n19039), .B2(n16999), .A(n16998), .ZN(n17005) );
  OAI21_X1 U20238 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17958), .A(
        n17000), .ZN(n17968) );
  INV_X1 U20239 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17154) );
  NOR2_X1 U20240 ( .A1(n9816), .A2(n17154), .ZN(n17183) );
  NOR2_X1 U20241 ( .A1(n18992), .A2(n17183), .ZN(n17115) );
  INV_X1 U20242 ( .A(n17115), .ZN(n17190) );
  AOI211_X1 U20243 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n17171), .A(
        n17968), .B(n17190), .ZN(n17004) );
  INV_X1 U20244 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17971) );
  NAND2_X1 U20245 ( .A1(n17001), .A2(n17968), .ZN(n17002) );
  OAI22_X1 U20246 ( .A1(n17971), .A2(n17181), .B1(n17101), .B2(n17002), .ZN(
        n17003) );
  NOR4_X1 U20247 ( .A1(n9731), .A2(n17005), .A3(n17004), .A4(n17003), .ZN(
        n17008) );
  OAI211_X1 U20248 ( .C1(n17016), .C2(n20865), .A(n17196), .B(n17006), .ZN(
        n17007) );
  OAI211_X1 U20249 ( .C1(n17163), .C2(n20865), .A(n17008), .B(n17007), .ZN(
        P3_U2656) );
  AOI21_X1 U20250 ( .B1(n17178), .B2(n17009), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n17021) );
  AOI21_X1 U20251 ( .B1(n17178), .B2(n17010), .A(n17185), .ZN(n17020) );
  INV_X1 U20252 ( .A(n18066), .ZN(n17048) );
  NOR2_X1 U20253 ( .A1(n18155), .A2(n17048), .ZN(n17045) );
  NAND2_X1 U20254 ( .A1(n18030), .A2(n17045), .ZN(n18001) );
  NOR2_X1 U20255 ( .A1(n18006), .A2(n18001), .ZN(n17012) );
  INV_X1 U20256 ( .A(n17958), .ZN(n17011) );
  OAI21_X1 U20257 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n17012), .A(
        n17011), .ZN(n17990) );
  INV_X1 U20258 ( .A(n17990), .ZN(n17014) );
  NOR2_X1 U20259 ( .A1(n18155), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17169) );
  INV_X1 U20260 ( .A(n17169), .ZN(n17138) );
  NOR2_X1 U20261 ( .A1(n17048), .A2(n17138), .ZN(n17102) );
  NAND2_X1 U20262 ( .A1(n18030), .A2(n17102), .ZN(n17037) );
  OAI21_X1 U20263 ( .B1(n18006), .B2(n17037), .A(n17171), .ZN(n17022) );
  INV_X1 U20264 ( .A(n17022), .ZN(n17013) );
  AOI221_X1 U20265 ( .B1(n17014), .B2(n17013), .C1(n17990), .C2(n17022), .A(
        n18992), .ZN(n17015) );
  AOI211_X1 U20266 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n17182), .A(
        n9731), .B(n17015), .ZN(n17019) );
  AOI211_X1 U20267 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17030), .A(n17016), .B(
        n17165), .ZN(n17017) );
  AOI21_X1 U20268 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17197), .A(n17017), .ZN(
        n17018) );
  OAI211_X1 U20269 ( .C1(n17021), .C2(n17020), .A(n17019), .B(n17018), .ZN(
        P3_U2657) );
  INV_X1 U20270 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17033) );
  OAI21_X1 U20271 ( .B1(n17041), .B2(n17173), .A(n17199), .ZN(n17058) );
  NOR2_X1 U20272 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17173), .ZN(n17040) );
  NOR2_X1 U20273 ( .A1(n18992), .A2(n17022), .ZN(n17027) );
  INV_X1 U20274 ( .A(n18001), .ZN(n17047) );
  NAND2_X1 U20275 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17047), .ZN(
        n17036) );
  INV_X1 U20276 ( .A(n17036), .ZN(n17023) );
  OAI22_X1 U20277 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17023), .B1(
        n18001), .B2(n18006), .ZN(n18009) );
  AOI211_X1 U20278 ( .C1(n17171), .C2(n17036), .A(n18009), .B(n17190), .ZN(
        n17026) );
  NOR3_X1 U20279 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17173), .A3(n17024), 
        .ZN(n17025) );
  AOI211_X1 U20280 ( .C1(n17027), .C2(n18009), .A(n17026), .B(n17025), .ZN(
        n17028) );
  OAI211_X1 U20281 ( .C1(n17163), .C2(n17405), .A(n17028), .B(n18455), .ZN(
        n17029) );
  AOI221_X1 U20282 ( .B1(n17058), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n17040), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n17029), .ZN(n17032) );
  OAI211_X1 U20283 ( .C1(n17034), .C2(n17405), .A(n17196), .B(n17030), .ZN(
        n17031) );
  OAI211_X1 U20284 ( .C1(n17181), .C2(n17033), .A(n17032), .B(n17031), .ZN(
        P3_U2658) );
  AOI211_X1 U20285 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17052), .A(n17034), .B(
        n17165), .ZN(n17035) );
  AOI21_X1 U20286 ( .B1(n17182), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n17035), .ZN(n17044) );
  OAI21_X1 U20287 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17047), .A(
        n17036), .ZN(n18015) );
  NAND2_X1 U20288 ( .A1(n17171), .A2(n17037), .ZN(n17038) );
  XOR2_X1 U20289 ( .A(n18015), .B(n17038), .Z(n17039) );
  AOI22_X1 U20290 ( .A1(n17197), .A2(P3_EBX_REG_12__SCAN_IN), .B1(n17184), 
        .B2(n17039), .ZN(n17043) );
  AOI22_X1 U20291 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n17058), .B1(n17041), 
        .B2(n17040), .ZN(n17042) );
  NAND4_X1 U20292 ( .A1(n17044), .A2(n17043), .A3(n17042), .A4(n18455), .ZN(
        P3_U2659) );
  OR2_X1 U20293 ( .A1(n17173), .A2(n17063), .ZN(n17080) );
  OAI21_X1 U20294 ( .B1(n17064), .B2(n17080), .A(n20772), .ZN(n17057) );
  INV_X1 U20295 ( .A(n17045), .ZN(n17114) );
  OR2_X1 U20296 ( .A1(n17046), .A2(n17114), .ZN(n17068) );
  AOI21_X1 U20297 ( .B1(n17055), .B2(n17068), .A(n17047), .ZN(n18033) );
  INV_X1 U20298 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18052) );
  NOR3_X1 U20299 ( .A1(n18155), .A2(n17048), .A3(n18083), .ZN(n17100) );
  NAND2_X1 U20300 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17100), .ZN(
        n17086) );
  NOR2_X1 U20301 ( .A1(n18052), .A2(n17086), .ZN(n17073) );
  INV_X1 U20302 ( .A(n17073), .ZN(n17049) );
  OAI21_X1 U20303 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17049), .A(
        n17171), .ZN(n17075) );
  OAI21_X1 U20304 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n9816), .A(
        n17075), .ZN(n17051) );
  AOI21_X1 U20305 ( .B1(n18033), .B2(n17051), .A(n18992), .ZN(n17050) );
  OAI21_X1 U20306 ( .B1(n18033), .B2(n17051), .A(n17050), .ZN(n17054) );
  OAI211_X1 U20307 ( .C1(n17061), .C2(n17060), .A(n17196), .B(n17052), .ZN(
        n17053) );
  OAI211_X1 U20308 ( .C1(n17181), .C2(n17055), .A(n17054), .B(n17053), .ZN(
        n17056) );
  AOI21_X1 U20309 ( .B1(n17058), .B2(n17057), .A(n17056), .ZN(n17059) );
  OAI211_X1 U20310 ( .C1(n17163), .C2(n17060), .A(n17059), .B(n18455), .ZN(
        P3_U2660) );
  INV_X1 U20311 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17072) );
  AOI211_X1 U20312 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17062), .A(n17061), .B(
        n17165), .ZN(n17067) );
  INV_X1 U20313 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19032) );
  AOI21_X1 U20314 ( .B1(n17178), .B2(n17063), .A(n17185), .ZN(n17090) );
  OAI21_X1 U20315 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(P3_REIP_REG_9__SCAN_IN), 
        .A(n17064), .ZN(n17065) );
  OAI22_X1 U20316 ( .A1(n19032), .A2(n17090), .B1(n17080), .B2(n17065), .ZN(
        n17066) );
  AOI211_X1 U20317 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17197), .A(n17067), .B(
        n17066), .ZN(n17071) );
  OAI21_X1 U20318 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17073), .A(
        n17068), .ZN(n18043) );
  XOR2_X1 U20319 ( .A(n18043), .B(n17075), .Z(n17069) );
  AOI21_X1 U20320 ( .B1(n17069), .B2(n17184), .A(n9731), .ZN(n17070) );
  OAI211_X1 U20321 ( .C1(n17181), .C2(n17072), .A(n17071), .B(n17070), .ZN(
        P3_U2661) );
  INV_X1 U20322 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19029) );
  AOI21_X1 U20323 ( .B1(n18067), .B2(n17102), .A(n9816), .ZN(n17076) );
  AOI21_X1 U20324 ( .B1(n18052), .B2(n17086), .A(n17073), .ZN(n18056) );
  INV_X1 U20325 ( .A(n18056), .ZN(n17074) );
  AOI221_X1 U20326 ( .B1(n17076), .B2(n18056), .C1(n17075), .C2(n17074), .A(
        n18992), .ZN(n17077) );
  AOI211_X1 U20327 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n17182), .A(
        n9731), .B(n17077), .ZN(n17085) );
  INV_X1 U20328 ( .A(n17079), .ZN(n17078) );
  OAI21_X1 U20329 ( .B1(n17165), .B2(n17078), .A(n17163), .ZN(n17083) );
  NOR2_X1 U20330 ( .A1(n17079), .A2(n17165), .ZN(n17095) );
  NOR2_X1 U20331 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17080), .ZN(n17081) );
  AOI221_X1 U20332 ( .B1(n17083), .B2(P3_EBX_REG_9__SCAN_IN), .C1(n17095), 
        .C2(n17082), .A(n17081), .ZN(n17084) );
  OAI211_X1 U20333 ( .C1(n19029), .C2(n17090), .A(n17085), .B(n17084), .ZN(
        P3_U2662) );
  AOI21_X1 U20334 ( .B1(n17100), .B2(n17154), .A(n9816), .ZN(n17087) );
  OAI21_X1 U20335 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17100), .A(
        n17086), .ZN(n18070) );
  XOR2_X1 U20336 ( .A(n17087), .B(n18070), .Z(n17088) );
  OAI22_X1 U20337 ( .A1(n18069), .A2(n17181), .B1(n18992), .B2(n17088), .ZN(
        n17094) );
  NAND2_X1 U20338 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n17106) );
  NOR2_X1 U20339 ( .A1(n17173), .A2(n17089), .ZN(n17124) );
  NAND2_X1 U20340 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17124), .ZN(n17123) );
  NOR2_X1 U20341 ( .A1(n17106), .A2(n17123), .ZN(n17092) );
  INV_X1 U20342 ( .A(n17090), .ZN(n17091) );
  MUX2_X1 U20343 ( .A(n17092), .B(n17091), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n17093) );
  NOR3_X1 U20344 ( .A1(n9731), .A2(n17094), .A3(n17093), .ZN(n17098) );
  INV_X1 U20345 ( .A(n17110), .ZN(n17096) );
  OAI21_X1 U20346 ( .B1(n17096), .B2(n17099), .A(n17095), .ZN(n17097) );
  OAI211_X1 U20347 ( .C1(n17099), .C2(n17163), .A(n17098), .B(n17097), .ZN(
        P3_U2663) );
  AOI21_X1 U20348 ( .B1(n18083), .B2(n17114), .A(n17100), .ZN(n18087) );
  OR2_X1 U20349 ( .A1(n17102), .A2(n17101), .ZN(n17118) );
  OAI211_X1 U20350 ( .C1(n17102), .C2(n9816), .A(n17184), .B(n18087), .ZN(
        n17103) );
  OAI211_X1 U20351 ( .C1(n18087), .C2(n17118), .A(n18455), .B(n17103), .ZN(
        n17109) );
  INV_X1 U20352 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19025) );
  OAI21_X1 U20353 ( .B1(n17173), .B2(n17104), .A(n17199), .ZN(n17105) );
  INV_X1 U20354 ( .A(n17105), .ZN(n17132) );
  OAI21_X1 U20355 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(P3_REIP_REG_6__SCAN_IN), 
        .A(n17106), .ZN(n17107) );
  OAI22_X1 U20356 ( .A1(n19025), .A2(n17132), .B1(n17123), .B2(n17107), .ZN(
        n17108) );
  AOI211_X1 U20357 ( .C1(n17197), .C2(P3_EBX_REG_7__SCAN_IN), .A(n17109), .B(
        n17108), .ZN(n17112) );
  OAI211_X1 U20358 ( .C1(n17113), .C2(n17435), .A(n17196), .B(n17110), .ZN(
        n17111) );
  OAI211_X1 U20359 ( .C1(n17181), .C2(n18083), .A(n17112), .B(n17111), .ZN(
        P3_U2664) );
  INV_X1 U20360 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19023) );
  AOI211_X1 U20361 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17129), .A(n17113), .B(
        n17165), .ZN(n17121) );
  NOR2_X1 U20362 ( .A1(n18155), .A2(n18095), .ZN(n17125) );
  OAI21_X1 U20363 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17125), .A(
        n17114), .ZN(n18096) );
  INV_X1 U20364 ( .A(n18096), .ZN(n17119) );
  OAI21_X1 U20365 ( .B1(n17125), .B2(n9816), .A(n17115), .ZN(n17117) );
  AOI21_X1 U20366 ( .B1(n17197), .B2(P3_EBX_REG_6__SCAN_IN), .A(n9731), .ZN(
        n17116) );
  OAI221_X1 U20367 ( .B1(n17119), .B2(n17118), .C1(n18096), .C2(n17117), .A(
        n17116), .ZN(n17120) );
  AOI211_X1 U20368 ( .C1(n17182), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n17121), .B(n17120), .ZN(n17122) );
  OAI221_X1 U20369 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17123), .C1(n19023), 
        .C2(n17132), .A(n17122), .ZN(P3_U2665) );
  NOR2_X1 U20370 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17124), .ZN(n17133) );
  INV_X1 U20371 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20716) );
  INV_X1 U20372 ( .A(n17137), .ZN(n18120) );
  NOR2_X1 U20373 ( .A1(n18155), .A2(n18120), .ZN(n17151) );
  NAND2_X1 U20374 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17151), .ZN(
        n17136) );
  AOI21_X1 U20375 ( .B1(n20716), .B2(n17136), .A(n17125), .ZN(n18109) );
  AOI21_X1 U20376 ( .B1(n17126), .B2(n17169), .A(n9816), .ZN(n17139) );
  XNOR2_X1 U20377 ( .A(n18109), .B(n17139), .ZN(n17127) );
  OAI22_X1 U20378 ( .A1(n17163), .A2(n17499), .B1(n18992), .B2(n17127), .ZN(
        n17128) );
  AOI211_X1 U20379 ( .C1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17182), .A(
        n9731), .B(n17128), .ZN(n17131) );
  OAI211_X1 U20380 ( .C1(n17134), .C2(n17499), .A(n17196), .B(n17129), .ZN(
        n17130) );
  OAI211_X1 U20381 ( .C1(n17133), .C2(n17132), .A(n17131), .B(n17130), .ZN(
        P3_U2666) );
  AOI211_X1 U20382 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17160), .A(n17134), .B(
        n17165), .ZN(n17144) );
  OAI21_X1 U20383 ( .B1(n17173), .B2(n17145), .A(n17199), .ZN(n17135) );
  INV_X1 U20384 ( .A(n17135), .ZN(n17149) );
  INV_X1 U20385 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20983) );
  NAND2_X1 U20386 ( .A1(n18485), .A2(n19146), .ZN(n17189) );
  INV_X1 U20387 ( .A(n17189), .ZN(n19147) );
  AOI221_X1 U20388 ( .B1(n17454), .B2(n19147), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n19147), .A(n9731), .ZN(
        n17142) );
  OAI21_X1 U20389 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17151), .A(
        n17136), .ZN(n18123) );
  INV_X1 U20390 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18122) );
  NAND2_X1 U20391 ( .A1(n17137), .A2(n18122), .ZN(n18118) );
  OAI22_X1 U20392 ( .A1(n17171), .A2(n18123), .B1(n17138), .B2(n18118), .ZN(
        n17140) );
  OAI221_X1 U20393 ( .B1(n17140), .B2(n17139), .C1(n17140), .C2(n18123), .A(
        n17184), .ZN(n17141) );
  OAI211_X1 U20394 ( .C1(n17149), .C2(n20983), .A(n17142), .B(n17141), .ZN(
        n17143) );
  AOI211_X1 U20395 ( .C1(n17182), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n17144), .B(n17143), .ZN(n17147) );
  NAND3_X1 U20396 ( .A1(n17178), .A2(n17145), .A3(n20983), .ZN(n17146) );
  OAI211_X1 U20397 ( .C1(n17148), .C2(n17163), .A(n17147), .B(n17146), .ZN(
        P3_U2667) );
  AOI221_X1 U20398 ( .B1(n17173), .B2(n19019), .C1(n17150), .C2(n19019), .A(
        n17149), .ZN(n17159) );
  NOR2_X1 U20399 ( .A1(n19109), .A2(n18948), .ZN(n18951) );
  OAI21_X1 U20400 ( .B1(n19085), .B2(n18951), .A(n12253), .ZN(n19083) );
  INV_X1 U20401 ( .A(n19083), .ZN(n17157) );
  NOR2_X1 U20402 ( .A1(n18155), .A2(n18150), .ZN(n17155) );
  INV_X1 U20403 ( .A(n17155), .ZN(n17167) );
  AOI21_X1 U20404 ( .B1(n17152), .B2(n17167), .A(n17151), .ZN(n18135) );
  AOI21_X1 U20405 ( .B1(n17155), .B2(n17154), .A(n9816), .ZN(n17168) );
  XNOR2_X1 U20406 ( .A(n18135), .B(n17168), .ZN(n17156) );
  OAI22_X1 U20407 ( .A1(n17157), .A2(n17189), .B1(n18992), .B2(n17156), .ZN(
        n17158) );
  AOI211_X1 U20408 ( .C1(n17182), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n17159), .B(n17158), .ZN(n17162) );
  OAI211_X1 U20409 ( .C1(n17166), .C2(n17164), .A(n17196), .B(n17160), .ZN(
        n17161) );
  OAI211_X1 U20410 ( .C1(n17164), .C2(n17163), .A(n17162), .B(n17161), .ZN(
        P3_U2668) );
  INV_X1 U20411 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17522) );
  INV_X1 U20412 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17518) );
  NAND2_X1 U20413 ( .A1(n17522), .A2(n17518), .ZN(n17186) );
  AOI211_X1 U20414 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17186), .A(n17166), .B(
        n17165), .ZN(n17177) );
  NAND2_X1 U20415 ( .A1(n19096), .A2(n18921), .ZN(n18949) );
  OAI21_X1 U20416 ( .B1(n18948), .B2(n19109), .A(n18949), .ZN(n19091) );
  OAI21_X1 U20417 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n17167), .ZN(n18145) );
  OAI21_X1 U20418 ( .B1(n17169), .B2(n18145), .A(n17168), .ZN(n17170) );
  OAI21_X1 U20419 ( .B1(n18145), .B2(n17171), .A(n17170), .ZN(n17172) );
  NAND2_X1 U20420 ( .A1(n17172), .A2(n17184), .ZN(n17175) );
  NOR2_X1 U20421 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17173), .ZN(n17192) );
  OAI21_X1 U20422 ( .B1(n17185), .B2(n17192), .A(P3_REIP_REG_2__SCAN_IN), .ZN(
        n17174) );
  OAI211_X1 U20423 ( .C1(n17189), .C2(n19091), .A(n17175), .B(n17174), .ZN(
        n17176) );
  AOI211_X1 U20424 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17197), .A(n17177), .B(
        n17176), .ZN(n17180) );
  INV_X1 U20425 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19016) );
  NAND3_X1 U20426 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17178), .A3(n19016), 
        .ZN(n17179) );
  OAI211_X1 U20427 ( .C1(n17181), .C2(n18150), .A(n17180), .B(n17179), .ZN(
        P3_U2669) );
  AOI21_X1 U20428 ( .B1(n17184), .B2(n17183), .A(n17182), .ZN(n17195) );
  AOI22_X1 U20429 ( .A1(n17197), .A2(P3_EBX_REG_1__SCAN_IN), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n17185), .ZN(n17194) );
  INV_X1 U20430 ( .A(n17186), .ZN(n17187) );
  AOI21_X1 U20431 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n17187), .ZN(n17516) );
  NAND2_X1 U20432 ( .A1(n17188), .A2(n18921), .ZN(n19097) );
  OAI22_X1 U20433 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17190), .B1(
        n17189), .B2(n19097), .ZN(n17191) );
  AOI211_X1 U20434 ( .C1(n17196), .C2(n17516), .A(n17192), .B(n17191), .ZN(
        n17193) );
  OAI211_X1 U20435 ( .C1(n17195), .C2(n18155), .A(n17194), .B(n17193), .ZN(
        P3_U2670) );
  NOR2_X1 U20436 ( .A1(n17197), .A2(n17196), .ZN(n17202) );
  AOI22_X1 U20437 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17198), .B1(n19147), 
        .B2(n19109), .ZN(n17201) );
  INV_X1 U20438 ( .A(n19144), .ZN(n19080) );
  NAND3_X1 U20439 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19080), .A3(
        n17199), .ZN(n17200) );
  OAI211_X1 U20440 ( .C1(n17202), .C2(n17522), .A(n17201), .B(n17200), .ZN(
        P3_U2671) );
  AND4_X1 U20441 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_24__SCAN_IN), .A4(P3_EBX_REG_23__SCAN_IN), .ZN(n17203)
         );
  AND4_X1 U20442 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n17203), .ZN(n17204) );
  NAND4_X1 U20443 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n17290), .A4(n17204), .ZN(n17207) );
  NOR2_X1 U20444 ( .A1(n17208), .A2(n17207), .ZN(n17233) );
  NAND2_X1 U20445 ( .A1(n17508), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17206) );
  NAND2_X1 U20446 ( .A1(n17233), .A2(n18516), .ZN(n17205) );
  OAI22_X1 U20447 ( .A1(n17233), .A2(n17206), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17205), .ZN(P3_U2672) );
  NAND2_X1 U20448 ( .A1(n17208), .A2(n17207), .ZN(n17209) );
  NAND2_X1 U20449 ( .A1(n17209), .A2(n17508), .ZN(n17232) );
  AOI22_X1 U20450 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n17453), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17213) );
  AOI22_X1 U20451 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U20452 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17211) );
  AOI22_X1 U20453 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17210) );
  NAND4_X1 U20454 ( .A1(n17213), .A2(n17212), .A3(n17211), .A4(n17210), .ZN(
        n17219) );
  AOI22_X1 U20455 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17217) );
  AOI22_X1 U20456 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U20457 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17215) );
  AOI22_X1 U20458 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17214) );
  NAND4_X1 U20459 ( .A1(n17217), .A2(n17216), .A3(n17215), .A4(n17214), .ZN(
        n17218) );
  NOR2_X1 U20460 ( .A1(n17219), .A2(n17218), .ZN(n17231) );
  AOI22_X1 U20461 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17230) );
  AOI22_X1 U20462 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17229) );
  AOI22_X1 U20463 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9734), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17220) );
  OAI21_X1 U20464 ( .B1(n20854), .B2(n9786), .A(n17220), .ZN(n17226) );
  AOI22_X1 U20465 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17224) );
  AOI22_X1 U20466 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17223) );
  AOI22_X1 U20467 ( .A1(n16122), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17222) );
  AOI22_X1 U20468 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17221) );
  NAND4_X1 U20469 ( .A1(n17224), .A2(n17223), .A3(n17222), .A4(n17221), .ZN(
        n17225) );
  AOI211_X1 U20470 ( .C1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .C2(n17227), .A(
        n17226), .B(n17225), .ZN(n17228) );
  NAND3_X1 U20471 ( .A1(n17230), .A2(n17229), .A3(n17228), .ZN(n17235) );
  NAND2_X1 U20472 ( .A1(n17236), .A2(n17235), .ZN(n17234) );
  XNOR2_X1 U20473 ( .A(n17231), .B(n17234), .ZN(n17534) );
  OAI22_X1 U20474 ( .A1(n17233), .A2(n17232), .B1(n17534), .B2(n17508), .ZN(
        P3_U2673) );
  OAI21_X1 U20475 ( .B1(n17236), .B2(n17235), .A(n17234), .ZN(n17542) );
  NAND3_X1 U20476 ( .A1(n17238), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17508), 
        .ZN(n17237) );
  OAI221_X1 U20477 ( .B1(n17238), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17508), 
        .C2(n17542), .A(n17237), .ZN(P3_U2674) );
  INV_X1 U20478 ( .A(n17239), .ZN(n17248) );
  AOI21_X1 U20479 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17508), .A(n17248), .ZN(
        n17242) );
  OAI21_X1 U20480 ( .B1(n17244), .B2(n17241), .A(n17240), .ZN(n17551) );
  OAI22_X1 U20481 ( .A1(n17243), .A2(n17242), .B1(n17551), .B2(n17508), .ZN(
        P3_U2676) );
  AOI21_X1 U20482 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17508), .A(n17253), .ZN(
        n17247) );
  AOI21_X1 U20483 ( .B1(n17245), .B2(n17250), .A(n17244), .ZN(n17552) );
  INV_X1 U20484 ( .A(n17552), .ZN(n17246) );
  OAI22_X1 U20485 ( .A1(n17248), .A2(n17247), .B1(n17508), .B2(n17246), .ZN(
        P3_U2677) );
  INV_X1 U20486 ( .A(n17249), .ZN(n17258) );
  AOI21_X1 U20487 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17508), .A(n17258), .ZN(
        n17252) );
  OAI21_X1 U20488 ( .B1(n17254), .B2(n17251), .A(n17250), .ZN(n17561) );
  OAI22_X1 U20489 ( .A1(n17253), .A2(n17252), .B1(n17508), .B2(n17561), .ZN(
        P3_U2678) );
  AOI21_X1 U20490 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17508), .A(n17264), .ZN(
        n17257) );
  AOI21_X1 U20491 ( .B1(n17255), .B2(n17260), .A(n17254), .ZN(n17562) );
  INV_X1 U20492 ( .A(n17562), .ZN(n17256) );
  OAI22_X1 U20493 ( .A1(n17258), .A2(n17257), .B1(n17508), .B2(n17256), .ZN(
        P3_U2679) );
  INV_X1 U20494 ( .A(n17259), .ZN(n17279) );
  AOI21_X1 U20495 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17508), .A(n17279), .ZN(
        n17263) );
  OAI21_X1 U20496 ( .B1(n17262), .B2(n17261), .A(n17260), .ZN(n17574) );
  OAI22_X1 U20497 ( .A1(n17264), .A2(n17263), .B1(n17508), .B2(n17574), .ZN(
        P3_U2680) );
  AOI21_X1 U20498 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17508), .A(n17265), .ZN(
        n17278) );
  AOI22_X1 U20499 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17276) );
  AOI22_X1 U20500 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n9729), .B1(
        n17311), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17275) );
  AOI22_X1 U20501 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17266) );
  OAI21_X1 U20502 ( .B1(n20854), .B2(n17267), .A(n17266), .ZN(n17273) );
  AOI22_X1 U20503 ( .A1(n17439), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17271) );
  AOI22_X1 U20504 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20505 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17269) );
  AOI22_X1 U20506 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17268) );
  NAND4_X1 U20507 ( .A1(n17271), .A2(n17270), .A3(n17269), .A4(n17268), .ZN(
        n17272) );
  AOI211_X1 U20508 ( .C1(n17460), .C2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n17273), .B(n17272), .ZN(n17274) );
  NAND3_X1 U20509 ( .A1(n17276), .A2(n17275), .A3(n17274), .ZN(n17576) );
  INV_X1 U20510 ( .A(n17576), .ZN(n17277) );
  OAI22_X1 U20511 ( .A1(n17279), .A2(n17278), .B1(n17277), .B2(n17508), .ZN(
        P3_U2681) );
  AOI22_X1 U20512 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17283) );
  AOI22_X1 U20513 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n17480), .B1(
        n17460), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20514 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17281) );
  AOI22_X1 U20515 ( .A1(n16122), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17280) );
  NAND4_X1 U20516 ( .A1(n17283), .A2(n17282), .A3(n17281), .A4(n17280), .ZN(
        n17289) );
  AOI22_X1 U20517 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17287) );
  AOI22_X1 U20518 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20519 ( .A1(n12189), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17285) );
  AOI22_X1 U20520 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17284) );
  NAND4_X1 U20521 ( .A1(n17287), .A2(n17286), .A3(n17285), .A4(n17284), .ZN(
        n17288) );
  NOR2_X1 U20522 ( .A1(n17289), .A2(n17288), .ZN(n17583) );
  NOR2_X1 U20523 ( .A1(n17520), .A2(n17290), .ZN(n17305) );
  INV_X1 U20524 ( .A(n17291), .ZN(n17293) );
  AOI22_X1 U20525 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17305), .B1(n17293), 
        .B2(n17292), .ZN(n17294) );
  OAI21_X1 U20526 ( .B1(n17583), .B2(n17508), .A(n17294), .ZN(P3_U2682) );
  AOI22_X1 U20527 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17298) );
  AOI22_X1 U20528 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17297) );
  AOI22_X1 U20529 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U20530 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17295) );
  NAND4_X1 U20531 ( .A1(n17298), .A2(n17297), .A3(n17296), .A4(n17295), .ZN(
        n17304) );
  AOI22_X1 U20532 ( .A1(n12188), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U20533 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20534 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U20535 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17299) );
  NAND4_X1 U20536 ( .A1(n17302), .A2(n17301), .A3(n17300), .A4(n17299), .ZN(
        n17303) );
  NOR2_X1 U20537 ( .A1(n17304), .A2(n17303), .ZN(n17590) );
  NAND2_X1 U20538 ( .A1(n18516), .A2(n17346), .ZN(n17347) );
  NOR3_X1 U20539 ( .A1(n17332), .A2(n17348), .A3(n17347), .ZN(n17320) );
  OAI221_X1 U20540 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(P3_EBX_REG_19__SCAN_IN), 
        .C1(P3_EBX_REG_20__SCAN_IN), .C2(n17320), .A(n17305), .ZN(n17306) );
  OAI21_X1 U20541 ( .B1(n17590), .B2(n17508), .A(n17306), .ZN(P3_U2683) );
  AOI22_X1 U20542 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U20543 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17309) );
  AOI22_X1 U20544 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17308) );
  AOI22_X1 U20545 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17473), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17307) );
  NAND4_X1 U20546 ( .A1(n17310), .A2(n17309), .A3(n17308), .A4(n17307), .ZN(
        n17317) );
  AOI22_X1 U20547 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n17311), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17315) );
  AOI22_X1 U20548 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17314) );
  AOI22_X1 U20549 ( .A1(n9729), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U20550 ( .A1(n12188), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17312) );
  NAND4_X1 U20551 ( .A1(n17315), .A2(n17314), .A3(n17313), .A4(n17312), .ZN(
        n17316) );
  NOR2_X1 U20552 ( .A1(n17317), .A2(n17316), .ZN(n17595) );
  AND2_X1 U20553 ( .A1(n17508), .A2(n17318), .ZN(n17333) );
  AOI22_X1 U20554 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17333), .B1(n17320), 
        .B2(n17319), .ZN(n17321) );
  OAI21_X1 U20555 ( .B1(n17595), .B2(n17508), .A(n17321), .ZN(P3_U2684) );
  AOI22_X1 U20556 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n16120), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U20557 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17324) );
  AOI22_X1 U20558 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n17461), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17323) );
  AOI22_X1 U20559 ( .A1(n16122), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17322) );
  NAND4_X1 U20560 ( .A1(n17325), .A2(n17324), .A3(n17323), .A4(n17322), .ZN(
        n17331) );
  AOI22_X1 U20561 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17329) );
  AOI22_X1 U20562 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20563 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20564 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17326) );
  NAND4_X1 U20565 ( .A1(n17329), .A2(n17328), .A3(n17327), .A4(n17326), .ZN(
        n17330) );
  NOR2_X1 U20566 ( .A1(n17331), .A2(n17330), .ZN(n17599) );
  OAI21_X1 U20567 ( .B1(n17348), .B2(n17347), .A(n17332), .ZN(n17334) );
  NAND2_X1 U20568 ( .A1(n17334), .A2(n17333), .ZN(n17335) );
  OAI21_X1 U20569 ( .B1(n17599), .B2(n17508), .A(n17335), .ZN(P3_U2685) );
  AOI22_X1 U20570 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17339) );
  AOI22_X1 U20571 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17338) );
  AOI22_X1 U20572 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17337) );
  AOI22_X1 U20573 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17474), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n16122), .ZN(n17336) );
  NAND4_X1 U20574 ( .A1(n17339), .A2(n17338), .A3(n17337), .A4(n17336), .ZN(
        n17345) );
  AOI22_X1 U20575 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17355), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17454), .ZN(n17343) );
  AOI22_X1 U20576 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17455), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n16120), .ZN(n17342) );
  AOI22_X1 U20577 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n17480), .ZN(n17341) );
  AOI22_X1 U20578 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17461), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17340) );
  NAND4_X1 U20579 ( .A1(n17343), .A2(n17342), .A3(n17341), .A4(n17340), .ZN(
        n17344) );
  NOR2_X1 U20580 ( .A1(n17345), .A2(n17344), .ZN(n17606) );
  NOR2_X1 U20581 ( .A1(n17520), .A2(n17346), .ZN(n17362) );
  INV_X1 U20582 ( .A(n17347), .ZN(n17349) );
  AOI22_X1 U20583 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17362), .B1(n17349), 
        .B2(n17348), .ZN(n17350) );
  OAI21_X1 U20584 ( .B1(n17606), .B2(n17508), .A(n17350), .ZN(P3_U2686) );
  AOI22_X1 U20585 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17354) );
  AOI22_X1 U20586 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U20587 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17352) );
  AOI22_X1 U20588 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17351) );
  NAND4_X1 U20589 ( .A1(n17354), .A2(n17353), .A3(n17352), .A4(n17351), .ZN(
        n17361) );
  AOI22_X1 U20590 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20591 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17355), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U20592 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20593 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n17439), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17356) );
  NAND4_X1 U20594 ( .A1(n17359), .A2(n17358), .A3(n17357), .A4(n17356), .ZN(
        n17360) );
  NOR2_X1 U20595 ( .A1(n17361), .A2(n17360), .ZN(n17613) );
  OAI21_X1 U20596 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17363), .A(n17362), .ZN(
        n17364) );
  OAI21_X1 U20597 ( .B1(n17613), .B2(n17508), .A(n17364), .ZN(P3_U2687) );
  AOI22_X1 U20598 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20599 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17373) );
  AOI22_X1 U20600 ( .A1(n17480), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U20601 ( .B1(n20718), .B2(n12156), .A(n17365), .ZN(n17371) );
  AOI22_X1 U20602 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20603 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17368) );
  AOI22_X1 U20604 ( .A1(n16120), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17367) );
  AOI22_X1 U20605 ( .A1(n17355), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17366) );
  NAND4_X1 U20606 ( .A1(n17369), .A2(n17368), .A3(n17367), .A4(n17366), .ZN(
        n17370) );
  AOI211_X1 U20607 ( .C1(n17481), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n17371), .B(n17370), .ZN(n17372) );
  NAND3_X1 U20608 ( .A1(n17374), .A2(n17373), .A3(n17372), .ZN(n17617) );
  INV_X1 U20609 ( .A(n17617), .ZN(n17378) );
  OAI21_X1 U20610 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17376), .A(n17375), .ZN(
        n17377) );
  AOI22_X1 U20611 ( .A1(n17520), .A2(n17378), .B1(n17377), .B2(n17508), .ZN(
        P3_U2688) );
  NAND2_X1 U20612 ( .A1(n18516), .A2(n17523), .ZN(n17503) );
  INV_X1 U20613 ( .A(n17503), .ZN(n17519) );
  NAND2_X1 U20614 ( .A1(n17379), .A2(n17519), .ZN(n17505) );
  NOR2_X1 U20615 ( .A1(n17380), .A2(n17505), .ZN(n17423) );
  NAND3_X1 U20616 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .A3(n17423), .ZN(n17393) );
  AOI22_X1 U20617 ( .A1(n16109), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20618 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20619 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20620 ( .B1(n20726), .B2(n10152), .A(n17381), .ZN(n17387) );
  AOI22_X1 U20621 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U20622 ( .A1(n17453), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17384) );
  AOI22_X1 U20623 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20624 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17382) );
  NAND4_X1 U20625 ( .A1(n17385), .A2(n17384), .A3(n17383), .A4(n17382), .ZN(
        n17386) );
  AOI211_X1 U20626 ( .C1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n17460), .A(
        n17387), .B(n17386), .ZN(n17388) );
  NAND3_X1 U20627 ( .A1(n17390), .A2(n17389), .A3(n17388), .ZN(n17620) );
  INV_X1 U20628 ( .A(n17620), .ZN(n17392) );
  NAND3_X1 U20629 ( .A1(n17393), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17508), 
        .ZN(n17391) );
  OAI221_X1 U20630 ( .B1(n17393), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17508), 
        .C2(n17392), .A(n17391), .ZN(P3_U2689) );
  AOI22_X1 U20631 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20632 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17396) );
  AOI22_X1 U20633 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U20634 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17394) );
  NAND4_X1 U20635 ( .A1(n17397), .A2(n17396), .A3(n17395), .A4(n17394), .ZN(
        n17403) );
  AOI22_X1 U20636 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20637 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U20638 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n17474), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20639 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9723), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17398) );
  NAND4_X1 U20640 ( .A1(n17401), .A2(n17400), .A3(n17399), .A4(n17398), .ZN(
        n17402) );
  NOR2_X1 U20641 ( .A1(n17403), .A2(n17402), .ZN(n17624) );
  OAI33_X1 U20642 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17647), .A3(n17406), 
        .B1(n17405), .B2(n17520), .B3(n17404), .ZN(n17407) );
  INV_X1 U20643 ( .A(n17407), .ZN(n17408) );
  OAI21_X1 U20644 ( .B1(n17624), .B2(n17508), .A(n17408), .ZN(P3_U2690) );
  AOI22_X1 U20645 ( .A1(n12188), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20646 ( .A1(n9723), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17409), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U20647 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17411) );
  AOI22_X1 U20648 ( .A1(n16122), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17410) );
  NAND4_X1 U20649 ( .A1(n17413), .A2(n17412), .A3(n17411), .A4(n17410), .ZN(
        n17420) );
  AOI22_X1 U20650 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17418) );
  AOI22_X1 U20651 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17417) );
  AOI22_X1 U20652 ( .A1(n17414), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17416) );
  AOI22_X1 U20653 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17461), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17415) );
  NAND4_X1 U20654 ( .A1(n17418), .A2(n17417), .A3(n17416), .A4(n17415), .ZN(
        n17419) );
  NOR2_X1 U20655 ( .A1(n17420), .A2(n17419), .ZN(n17628) );
  NOR2_X1 U20656 ( .A1(n17520), .A2(n17421), .ZN(n17437) );
  INV_X1 U20657 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U20658 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17437), .B1(n17423), 
        .B2(n17422), .ZN(n17424) );
  OAI21_X1 U20659 ( .B1(n17628), .B2(n17508), .A(n17424), .ZN(P3_U2691) );
  AOI22_X1 U20660 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n17454), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20661 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U20662 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20663 ( .A1(n9734), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17425) );
  NAND4_X1 U20664 ( .A1(n17428), .A2(n17427), .A3(n17426), .A4(n17425), .ZN(
        n17434) );
  AOI22_X1 U20665 ( .A1(n17462), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20666 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20667 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n9723), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20668 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17429) );
  NAND4_X1 U20669 ( .A1(n17432), .A2(n17431), .A3(n17430), .A4(n17429), .ZN(
        n17433) );
  NOR2_X1 U20670 ( .A1(n17434), .A2(n17433), .ZN(n17631) );
  INV_X1 U20671 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17436) );
  OR2_X1 U20672 ( .A1(n17499), .A2(n17498), .ZN(n17494) );
  NOR3_X1 U20673 ( .A1(n17435), .A2(n17497), .A3(n17494), .ZN(n17493) );
  AND2_X1 U20674 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17493), .ZN(n17488) );
  NAND2_X1 U20675 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17488), .ZN(n17450) );
  NOR2_X1 U20676 ( .A1(n17436), .A2(n17450), .ZN(n17452) );
  OAI21_X1 U20677 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17452), .A(n17437), .ZN(
        n17438) );
  OAI21_X1 U20678 ( .B1(n17631), .B2(n17508), .A(n17438), .ZN(P3_U2692) );
  AOI22_X1 U20679 ( .A1(n17472), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U20680 ( .A1(n17479), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20681 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n17480), .B1(
        n17471), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U20682 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n17439), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17440) );
  NAND4_X1 U20683 ( .A1(n17443), .A2(n17442), .A3(n17441), .A4(n17440), .ZN(
        n17449) );
  AOI22_X1 U20684 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17474), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U20685 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17462), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U20686 ( .A1(n9722), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U20687 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9729), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17444) );
  NAND4_X1 U20688 ( .A1(n17447), .A2(n17446), .A3(n17445), .A4(n17444), .ZN(
        n17448) );
  NOR2_X1 U20689 ( .A1(n17449), .A2(n17448), .ZN(n17638) );
  NOR2_X1 U20690 ( .A1(n17647), .A2(n17450), .ZN(n17470) );
  OAI21_X1 U20691 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17470), .A(n17508), .ZN(
        n17451) );
  OAI22_X1 U20692 ( .A1(n17638), .A2(n17508), .B1(n17452), .B2(n17451), .ZN(
        P3_U2693) );
  AOI22_X1 U20693 ( .A1(n17311), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9729), .ZN(n17459) );
  AOI22_X1 U20694 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17453), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20695 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17471), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17454), .ZN(n17457) );
  AOI22_X1 U20696 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17473), .B1(
        n17455), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17456) );
  NAND4_X1 U20697 ( .A1(n17459), .A2(n17458), .A3(n17457), .A4(n17456), .ZN(
        n17468) );
  AOI22_X1 U20698 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n16109), .ZN(n17466) );
  AOI22_X1 U20699 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n16120), .ZN(n17465) );
  AOI22_X1 U20700 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17474), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17461), .ZN(n17464) );
  AOI22_X1 U20701 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17462), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17480), .ZN(n17463) );
  NAND4_X1 U20702 ( .A1(n17466), .A2(n17465), .A3(n17464), .A4(n17463), .ZN(
        n17467) );
  NOR2_X1 U20703 ( .A1(n17468), .A2(n17467), .ZN(n17640) );
  NOR3_X1 U20704 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17520), .A3(n17488), .ZN(
        n17469) );
  AOI211_X1 U20705 ( .C1(n17640), .C2(n17520), .A(n17470), .B(n17469), .ZN(
        P3_U2694) );
  AOI22_X1 U20706 ( .A1(n17227), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n16109), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20707 ( .A1(n17471), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17454), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17477) );
  AOI22_X1 U20708 ( .A1(n12188), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17472), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20709 ( .A1(n17474), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17473), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17475) );
  NAND4_X1 U20710 ( .A1(n17478), .A2(n17477), .A3(n17476), .A4(n17475), .ZN(
        n17487) );
  AOI22_X1 U20711 ( .A1(n17460), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9722), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U20712 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n9729), .B1(
        n17479), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20713 ( .A1(n17481), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17480), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17483) );
  AOI22_X1 U20714 ( .A1(n17455), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n16120), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17482) );
  NAND4_X1 U20715 ( .A1(n17485), .A2(n17484), .A3(n17483), .A4(n17482), .ZN(
        n17486) );
  NOR2_X1 U20716 ( .A1(n17487), .A2(n17486), .ZN(n17646) );
  NOR2_X1 U20717 ( .A1(n17520), .A2(n17488), .ZN(n17489) );
  OAI21_X1 U20718 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17493), .A(n17489), .ZN(
        n17490) );
  OAI21_X1 U20719 ( .B1(n17646), .B2(n17508), .A(n17490), .ZN(P3_U2695) );
  NOR2_X1 U20720 ( .A1(n17647), .A2(n17494), .ZN(n17495) );
  AOI22_X1 U20721 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17508), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17495), .ZN(n17492) );
  INV_X1 U20722 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17491) );
  OAI22_X1 U20723 ( .A1(n17493), .A2(n17492), .B1(n17491), .B2(n17508), .ZN(
        P3_U2696) );
  NAND2_X1 U20724 ( .A1(n17508), .A2(n17494), .ZN(n17501) );
  AOI22_X1 U20725 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17520), .B1(
        n17495), .B2(n17497), .ZN(n17496) );
  OAI21_X1 U20726 ( .B1(n17497), .B2(n17501), .A(n17496), .ZN(P3_U2697) );
  AND2_X1 U20727 ( .A1(n17499), .A2(n17498), .ZN(n17502) );
  INV_X1 U20728 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17500) );
  OAI22_X1 U20729 ( .A1(n17502), .A2(n17501), .B1(n17500), .B2(n17508), .ZN(
        P3_U2698) );
  NOR2_X1 U20730 ( .A1(n17504), .A2(n17503), .ZN(n17513) );
  AND2_X1 U20731 ( .A1(P3_EBX_REG_3__SCAN_IN), .A2(n17513), .ZN(n17511) );
  OAI211_X1 U20732 ( .C1(n17511), .C2(P3_EBX_REG_4__SCAN_IN), .A(n17508), .B(
        n17505), .ZN(n17506) );
  OAI21_X1 U20733 ( .B1(n17508), .B2(n17507), .A(n17506), .ZN(P3_U2699) );
  AOI21_X1 U20734 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17508), .A(n17513), .ZN(
        n17510) );
  INV_X1 U20735 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17509) );
  OAI22_X1 U20736 ( .A1(n17511), .A2(n17510), .B1(n17509), .B2(n17508), .ZN(
        P3_U2700) );
  INV_X1 U20737 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17515) );
  NOR2_X1 U20738 ( .A1(n17522), .A2(n17518), .ZN(n17512) );
  AOI211_X1 U20739 ( .C1(n17520), .C2(n17515), .A(n17514), .B(n17513), .ZN(
        P3_U2701) );
  AOI22_X1 U20740 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17520), .B1(
        n17516), .B2(n17519), .ZN(n17517) );
  OAI21_X1 U20741 ( .B1(n17523), .B2(n17518), .A(n17517), .ZN(P3_U2702) );
  AOI22_X1 U20742 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17520), .B1(
        n17519), .B2(n17522), .ZN(n17521) );
  OAI21_X1 U20743 ( .B1(n17523), .B2(n17522), .A(n17521), .ZN(P3_U2703) );
  NAND2_X1 U20744 ( .A1(n17647), .A2(n17524), .ZN(n17673) );
  NOR2_X1 U20745 ( .A1(n17673), .A2(n18510), .ZN(n17607) );
  INV_X1 U20746 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17751) );
  INV_X1 U20747 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17747) );
  INV_X1 U20748 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17745) );
  INV_X1 U20749 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17743) );
  NAND4_X1 U20750 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17525) );
  NAND4_X1 U20751 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(n17526), .ZN(n17643) );
  AND4_X1 U20752 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .A3(P3_EAX_REG_10__SCAN_IN), .A4(P3_EAX_REG_9__SCAN_IN), .ZN(n17527)
         );
  NAND4_X1 U20753 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_14__SCAN_IN), 
        .A3(P3_EAX_REG_13__SCAN_IN), .A4(n17527), .ZN(n17614) );
  NOR2_X2 U20754 ( .A1(n17643), .A2(n17614), .ZN(n17616) );
  AND2_X2 U20755 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17616), .ZN(n17610) );
  AND4_X1 U20756 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17528)
         );
  NAND4_X1 U20757 ( .A1(n17575), .A2(P3_EAX_REG_21__SCAN_IN), .A3(
        P3_EAX_REG_20__SCAN_IN), .A4(n17528), .ZN(n17570) );
  NOR2_X2 U20758 ( .A1(n17743), .A2(n17570), .ZN(n17569) );
  NAND2_X1 U20759 ( .A1(n18516), .A2(n17569), .ZN(n17563) );
  OR2_X2 U20760 ( .A1(n17745), .A2(n17563), .ZN(n17564) );
  NOR2_X2 U20761 ( .A1(n17747), .A2(n17564), .ZN(n17557) );
  NAND2_X1 U20762 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17547), .ZN(n17544) );
  NAND2_X1 U20763 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17539), .ZN(n17538) );
  NOR2_X1 U20764 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17538), .ZN(n17530) );
  NAND2_X1 U20765 ( .A1(n17673), .A2(n17538), .ZN(n17537) );
  OAI21_X1 U20766 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17577), .A(n17537), .ZN(
        n17529) );
  AOI22_X1 U20767 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17530), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17529), .ZN(n17531) );
  OAI21_X1 U20768 ( .B1(n17532), .B2(n17582), .A(n17531), .ZN(P3_U2704) );
  INV_X1 U20769 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17757) );
  NOR2_X2 U20770 ( .A1(n17533), .A2(n17673), .ZN(n17608) );
  OAI22_X1 U20771 ( .A1(n17534), .A2(n17666), .B1(n14698), .B2(n17582), .ZN(
        n17535) );
  AOI21_X1 U20772 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17608), .A(n17535), .ZN(
        n17536) );
  OAI221_X1 U20773 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17538), .C1(n17757), 
        .C2(n17537), .A(n17536), .ZN(P3_U2705) );
  AOI22_X1 U20774 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17608), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17607), .ZN(n17541) );
  OAI211_X1 U20775 ( .C1(n17539), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17673), .B(
        n17538), .ZN(n17540) );
  OAI211_X1 U20776 ( .C1(n17542), .C2(n17666), .A(n17541), .B(n17540), .ZN(
        P3_U2706) );
  AOI22_X1 U20777 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17608), .B1(n17671), .B2(
        n17543), .ZN(n17546) );
  OAI211_X1 U20778 ( .C1(n17547), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17673), .B(
        n17544), .ZN(n17545) );
  OAI211_X1 U20779 ( .C1(n17582), .C2(n18499), .A(n17546), .B(n17545), .ZN(
        P3_U2707) );
  AOI22_X1 U20780 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17608), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17607), .ZN(n17550) );
  INV_X1 U20781 ( .A(n17673), .ZN(n17635) );
  AOI211_X1 U20782 ( .C1(n17751), .C2(n17553), .A(n17547), .B(n17635), .ZN(
        n17548) );
  INV_X1 U20783 ( .A(n17548), .ZN(n17549) );
  OAI211_X1 U20784 ( .C1(n17551), .C2(n17666), .A(n17550), .B(n17549), .ZN(
        P3_U2708) );
  INV_X1 U20785 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U20786 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17608), .B1(n17671), .B2(
        n17552), .ZN(n17555) );
  OAI211_X1 U20787 ( .C1(n17557), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17673), .B(
        n17553), .ZN(n17554) );
  OAI211_X1 U20788 ( .C1(n17582), .C2(n17556), .A(n17555), .B(n17554), .ZN(
        P3_U2709) );
  AOI22_X1 U20789 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17608), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17607), .ZN(n17560) );
  AOI211_X1 U20790 ( .C1(n17747), .C2(n17564), .A(n17557), .B(n17635), .ZN(
        n17558) );
  INV_X1 U20791 ( .A(n17558), .ZN(n17559) );
  OAI211_X1 U20792 ( .C1(n17561), .C2(n17666), .A(n17560), .B(n17559), .ZN(
        P3_U2710) );
  INV_X1 U20793 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U20794 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17608), .B1(n17671), .B2(
        n17562), .ZN(n17567) );
  OAI21_X1 U20795 ( .B1(n17745), .B2(n17635), .A(n17563), .ZN(n17565) );
  NAND2_X1 U20796 ( .A1(n17565), .A2(n17564), .ZN(n17566) );
  OAI211_X1 U20797 ( .C1(n17582), .C2(n17568), .A(n17567), .B(n17566), .ZN(
        P3_U2711) );
  AOI211_X1 U20798 ( .C1(n17743), .C2(n17570), .A(n17635), .B(n17569), .ZN(
        n17571) );
  AOI21_X1 U20799 ( .B1(n17607), .B2(BUF2_REG_23__SCAN_IN), .A(n17571), .ZN(
        n17573) );
  NAND2_X1 U20800 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17608), .ZN(n17572) );
  OAI211_X1 U20801 ( .C1(n17574), .C2(n17666), .A(n17573), .B(n17572), .ZN(
        P3_U2712) );
  INV_X1 U20802 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17736) );
  INV_X1 U20803 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17733) );
  NAND2_X1 U20804 ( .A1(n18516), .A2(n17575), .ZN(n17600) );
  NAND2_X1 U20805 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17601), .ZN(n17596) );
  NAND3_X1 U20806 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(n17591), .ZN(n17581) );
  AOI22_X1 U20807 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17607), .B1(n17671), .B2(
        n17576), .ZN(n17580) );
  NAND2_X1 U20808 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17591), .ZN(n17587) );
  NAND2_X1 U20809 ( .A1(n17673), .A2(n17587), .ZN(n17586) );
  OAI21_X1 U20810 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17577), .A(n17586), .ZN(
        n17578) );
  AOI22_X1 U20811 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17608), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17578), .ZN(n17579) );
  OAI211_X1 U20812 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17581), .A(n17580), .B(
        n17579), .ZN(P3_U2713) );
  INV_X1 U20813 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17739) );
  OAI22_X1 U20814 ( .A1(n17583), .A2(n17666), .B1(n15580), .B2(n17582), .ZN(
        n17584) );
  AOI21_X1 U20815 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17608), .A(n17584), .ZN(
        n17585) );
  OAI221_X1 U20816 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17587), .C1(n17739), 
        .C2(n17586), .A(n17585), .ZN(P3_U2714) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n17608), .ZN(n17589) );
  OAI211_X1 U20818 ( .C1(n17591), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17673), .B(
        n17587), .ZN(n17588) );
  OAI211_X1 U20819 ( .C1(n17590), .C2(n17666), .A(n17589), .B(n17588), .ZN(
        P3_U2715) );
  AOI22_X1 U20820 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17608), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17607), .ZN(n17594) );
  AOI211_X1 U20821 ( .C1(n17736), .C2(n17596), .A(n17591), .B(n17635), .ZN(
        n17592) );
  INV_X1 U20822 ( .A(n17592), .ZN(n17593) );
  OAI211_X1 U20823 ( .C1(n17595), .C2(n17666), .A(n17594), .B(n17593), .ZN(
        P3_U2716) );
  AOI22_X1 U20824 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17608), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17607), .ZN(n17598) );
  OAI211_X1 U20825 ( .C1(n17601), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17673), .B(
        n17596), .ZN(n17597) );
  OAI211_X1 U20826 ( .C1(n17599), .C2(n17666), .A(n17598), .B(n17597), .ZN(
        P3_U2717) );
  AOI22_X1 U20827 ( .A1(BUF2_REG_17__SCAN_IN), .A2(n17607), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n17608), .ZN(n17605) );
  OAI21_X1 U20828 ( .B1(n17733), .B2(n17635), .A(n17600), .ZN(n17603) );
  INV_X1 U20829 ( .A(n17601), .ZN(n17602) );
  NAND2_X1 U20830 ( .A1(n17603), .A2(n17602), .ZN(n17604) );
  OAI211_X1 U20831 ( .C1(n17606), .C2(n17666), .A(n17605), .B(n17604), .ZN(
        P3_U2718) );
  AOI22_X1 U20832 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17608), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17607), .ZN(n17612) );
  OAI211_X1 U20833 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17610), .A(n17673), .B(
        n17609), .ZN(n17611) );
  OAI211_X1 U20834 ( .C1(n17613), .C2(n17666), .A(n17612), .B(n17611), .ZN(
        P3_U2719) );
  INV_X1 U20835 ( .A(n17614), .ZN(n17615) );
  NOR2_X1 U20836 ( .A1(n17647), .A2(n17643), .ZN(n17650) );
  NAND2_X1 U20837 ( .A1(n17615), .A2(n17650), .ZN(n17619) );
  INV_X1 U20838 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17789) );
  OR2_X1 U20839 ( .A1(n17635), .A2(n17616), .ZN(n17622) );
  INV_X1 U20840 ( .A(n17669), .ZN(n17672) );
  AOI22_X1 U20841 ( .A1(n17671), .A2(n17617), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17672), .ZN(n17618) );
  OAI221_X1 U20842 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17619), .C1(n17789), 
        .C2(n17622), .A(n17618), .ZN(P3_U2720) );
  INV_X1 U20843 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17701) );
  INV_X1 U20844 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17774) );
  NAND3_X1 U20845 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17650), .ZN(n17639) );
  NAND2_X1 U20846 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17634), .ZN(n17627) );
  NOR2_X1 U20847 ( .A1(n17701), .A2(n17627), .ZN(n17630) );
  NAND2_X1 U20848 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17630), .ZN(n17623) );
  INV_X1 U20849 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17784) );
  AOI22_X1 U20850 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17672), .B1(n17671), .B2(
        n17620), .ZN(n17621) );
  OAI221_X1 U20851 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17623), .C1(n17784), 
        .C2(n17622), .A(n17621), .ZN(P3_U2721) );
  INV_X1 U20852 ( .A(n17623), .ZN(n17626) );
  AOI21_X1 U20853 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17673), .A(n17630), .ZN(
        n17625) );
  OAI222_X1 U20854 ( .A1(n17669), .A2(n17782), .B1(n17626), .B2(n17625), .C1(
        n17666), .C2(n17624), .ZN(P3_U2722) );
  INV_X1 U20855 ( .A(n17627), .ZN(n17633) );
  AOI21_X1 U20856 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17673), .A(n17633), .ZN(
        n17629) );
  OAI222_X1 U20857 ( .A1(n17669), .A2(n17778), .B1(n17630), .B2(n17629), .C1(
        n17666), .C2(n17628), .ZN(P3_U2723) );
  AOI21_X1 U20858 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17673), .A(n17634), .ZN(
        n17632) );
  OAI222_X1 U20859 ( .A1(n17669), .A2(n17776), .B1(n17633), .B2(n17632), .C1(
        n17666), .C2(n17631), .ZN(P3_U2724) );
  AOI211_X1 U20860 ( .C1(n17774), .C2(n17639), .A(n17635), .B(n17634), .ZN(
        n17636) );
  AOI21_X1 U20861 ( .B1(n17672), .B2(BUF2_REG_10__SCAN_IN), .A(n17636), .ZN(
        n17637) );
  OAI21_X1 U20862 ( .B1(n17638), .B2(n17666), .A(n17637), .ZN(P3_U2725) );
  INV_X1 U20863 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17772) );
  INV_X1 U20864 ( .A(n17639), .ZN(n17642) );
  AOI22_X1 U20865 ( .A1(n17650), .A2(P3_EAX_REG_8__SCAN_IN), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17673), .ZN(n17641) );
  OAI222_X1 U20866 ( .A1(n17669), .A2(n17772), .B1(n17642), .B2(n17641), .C1(
        n17666), .C2(n17640), .ZN(P3_U2726) );
  INV_X1 U20867 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17770) );
  AOI22_X1 U20868 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17672), .B1(n17650), .B2(
        n17770), .ZN(n17645) );
  NAND3_X1 U20869 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17673), .A3(n17643), .ZN(
        n17644) );
  OAI211_X1 U20870 ( .C1(n17646), .C2(n17666), .A(n17645), .B(n17644), .ZN(
        P3_U2727) );
  INV_X1 U20871 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17711) );
  INV_X1 U20872 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17716) );
  INV_X1 U20873 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17761) );
  NOR3_X1 U20874 ( .A1(n17647), .A2(n17674), .A3(n17761), .ZN(n17664) );
  AND2_X1 U20875 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17664), .ZN(n17668) );
  NAND2_X1 U20876 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17668), .ZN(n17658) );
  NOR2_X1 U20877 ( .A1(n17716), .A2(n17658), .ZN(n17659) );
  NAND2_X1 U20878 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17659), .ZN(n17651) );
  NOR2_X1 U20879 ( .A1(n17711), .A2(n17651), .ZN(n17653) );
  AOI21_X1 U20880 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17673), .A(n17653), .ZN(
        n17649) );
  OAI222_X1 U20881 ( .A1(n17669), .A2(n18513), .B1(n17650), .B2(n17649), .C1(
        n17666), .C2(n17648), .ZN(P3_U2728) );
  INV_X1 U20882 ( .A(n17651), .ZN(n17656) );
  AOI21_X1 U20883 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17673), .A(n17656), .ZN(
        n17654) );
  OAI222_X1 U20884 ( .A1(n17669), .A2(n18509), .B1(n17654), .B2(n17653), .C1(
        n17666), .C2(n17652), .ZN(P3_U2729) );
  AOI21_X1 U20885 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17673), .A(n17659), .ZN(
        n17657) );
  OAI222_X1 U20886 ( .A1(n17669), .A2(n18505), .B1(n17657), .B2(n17656), .C1(
        n17666), .C2(n17655), .ZN(P3_U2730) );
  INV_X1 U20887 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18500) );
  INV_X1 U20888 ( .A(n17658), .ZN(n17663) );
  AOI21_X1 U20889 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17673), .A(n17663), .ZN(
        n17660) );
  OAI222_X1 U20890 ( .A1(n17669), .A2(n18500), .B1(n17660), .B2(n17659), .C1(
        n17666), .C2(n9891), .ZN(P3_U2731) );
  AOI21_X1 U20891 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17673), .A(n17668), .ZN(
        n17662) );
  OAI222_X1 U20892 ( .A1(n18495), .A2(n17669), .B1(n17663), .B2(n17662), .C1(
        n17666), .C2(n17661), .ZN(P3_U2732) );
  AOI21_X1 U20893 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17673), .A(n17664), .ZN(
        n17667) );
  OAI222_X1 U20894 ( .A1(n18490), .A2(n17669), .B1(n17668), .B2(n17667), .C1(
        n17666), .C2(n17665), .ZN(P3_U2733) );
  AOI22_X1 U20895 ( .A1(n17672), .A2(BUF2_REG_1__SCAN_IN), .B1(n17671), .B2(
        n17670), .ZN(n17677) );
  OAI221_X1 U20896 ( .B1(n17675), .B2(P3_EAX_REG_1__SCAN_IN), .C1(n17674), 
        .C2(n17761), .A(n17673), .ZN(n17676) );
  NAND2_X1 U20897 ( .A1(n17677), .A2(n17676), .ZN(P3_U2734) );
  NAND2_X1 U20898 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18002), .ZN(n17714) );
  NAND2_X1 U20899 ( .A1(n17714), .A2(n17724), .ZN(n17703) );
  NOR2_X1 U20900 ( .A1(n17703), .A2(n17679), .ZN(P3_U2736) );
  NOR2_X1 U20901 ( .A1(n17724), .A2(n18485), .ZN(n17692) );
  AOI22_X1 U20902 ( .A1(n17722), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17680) );
  OAI21_X1 U20903 ( .B1(n17757), .B2(n17696), .A(n17680), .ZN(P3_U2737) );
  INV_X1 U20904 ( .A(P3_UWORD_REG_13__SCAN_IN), .ZN(n20754) );
  AOI22_X1 U20905 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17692), .B1(n17721), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17681) );
  OAI21_X1 U20906 ( .B1(n20754), .B2(n17714), .A(n17681), .ZN(P3_U2738) );
  INV_X1 U20907 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17753) );
  AOI22_X1 U20908 ( .A1(n17722), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17682) );
  OAI21_X1 U20909 ( .B1(n17753), .B2(n17696), .A(n17682), .ZN(P3_U2739) );
  AOI22_X1 U20910 ( .A1(n17722), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17683) );
  OAI21_X1 U20911 ( .B1(n17751), .B2(n17696), .A(n17683), .ZN(P3_U2740) );
  INV_X1 U20912 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17749) );
  AOI22_X1 U20913 ( .A1(n17722), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17684) );
  OAI21_X1 U20914 ( .B1(n17749), .B2(n17696), .A(n17684), .ZN(P3_U2741) );
  AOI22_X1 U20915 ( .A1(n17722), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17685) );
  OAI21_X1 U20916 ( .B1(n17747), .B2(n17696), .A(n17685), .ZN(P3_U2742) );
  AOI22_X1 U20917 ( .A1(n17722), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17686) );
  OAI21_X1 U20918 ( .B1(n17745), .B2(n17696), .A(n17686), .ZN(P3_U2743) );
  AOI22_X1 U20919 ( .A1(n17722), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17687) );
  OAI21_X1 U20920 ( .B1(n17743), .B2(n17696), .A(n17687), .ZN(P3_U2744) );
  INV_X1 U20921 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17741) );
  AOI22_X1 U20922 ( .A1(n17722), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17688) );
  OAI21_X1 U20923 ( .B1(n17741), .B2(n17696), .A(n17688), .ZN(P3_U2745) );
  AOI22_X1 U20924 ( .A1(n17722), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20925 ( .B1(n17739), .B2(n17696), .A(n17689), .ZN(P3_U2746) );
  INV_X1 U20926 ( .A(P3_UWORD_REG_4__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U20927 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17692), .B1(n17721), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17690) );
  OAI21_X1 U20928 ( .B1(n20942), .B2(n17714), .A(n17690), .ZN(P3_U2747) );
  AOI22_X1 U20929 ( .A1(n17722), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17691) );
  OAI21_X1 U20930 ( .B1(n17736), .B2(n17696), .A(n17691), .ZN(P3_U2748) );
  INV_X1 U20931 ( .A(P3_UWORD_REG_2__SCAN_IN), .ZN(n20845) );
  AOI22_X1 U20932 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17692), .B1(n17721), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17693) );
  OAI21_X1 U20933 ( .B1(n20845), .B2(n17714), .A(n17693), .ZN(P3_U2749) );
  AOI22_X1 U20934 ( .A1(n17722), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17694) );
  OAI21_X1 U20935 ( .B1(n17733), .B2(n17696), .A(n17694), .ZN(P3_U2750) );
  INV_X1 U20936 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17731) );
  AOI22_X1 U20937 ( .A1(n17722), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17695) );
  OAI21_X1 U20938 ( .B1(n17731), .B2(n17696), .A(n17695), .ZN(P3_U2751) );
  AOI22_X1 U20939 ( .A1(n17722), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17697) );
  OAI21_X1 U20940 ( .B1(n17789), .B2(n17724), .A(n17697), .ZN(P3_U2752) );
  AOI22_X1 U20941 ( .A1(n17722), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17698) );
  OAI21_X1 U20942 ( .B1(n17784), .B2(n17724), .A(n17698), .ZN(P3_U2753) );
  AOI222_X1 U20943 ( .A1(n17712), .A2(P3_EAX_REG_13__SCAN_IN), .B1(n17722), 
        .B2(P3_LWORD_REG_13__SCAN_IN), .C1(P3_DATAO_REG_13__SCAN_IN), .C2(
        n17721), .ZN(n17699) );
  INV_X1 U20944 ( .A(n17699), .ZN(P3_U2754) );
  AOI22_X1 U20945 ( .A1(n17722), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17700) );
  OAI21_X1 U20946 ( .B1(n17701), .B2(n17724), .A(n17700), .ZN(P3_U2755) );
  INV_X1 U20947 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n20923) );
  AOI22_X1 U20948 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17712), .B1(n17722), 
        .B2(P3_LWORD_REG_11__SCAN_IN), .ZN(n17702) );
  OAI21_X1 U20949 ( .B1(n20923), .B2(n17703), .A(n17702), .ZN(P3_U2756) );
  AOI22_X1 U20950 ( .A1(n17722), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17704) );
  OAI21_X1 U20951 ( .B1(n17774), .B2(n17724), .A(n17704), .ZN(P3_U2757) );
  INV_X1 U20952 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U20953 ( .A1(n17722), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17705) );
  OAI21_X1 U20954 ( .B1(n17706), .B2(n17724), .A(n17705), .ZN(P3_U2758) );
  AOI22_X1 U20955 ( .A1(n17722), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17707) );
  OAI21_X1 U20956 ( .B1(n17770), .B2(n17724), .A(n17707), .ZN(P3_U2759) );
  INV_X1 U20957 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17709) );
  AOI22_X1 U20958 ( .A1(n17722), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17708) );
  OAI21_X1 U20959 ( .B1(n17709), .B2(n17724), .A(n17708), .ZN(P3_U2760) );
  AOI22_X1 U20960 ( .A1(n17722), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17710) );
  OAI21_X1 U20961 ( .B1(n17711), .B2(n17724), .A(n17710), .ZN(P3_U2761) );
  INV_X1 U20962 ( .A(P3_LWORD_REG_5__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U20963 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17712), .B1(n17721), .B2(
        P3_DATAO_REG_5__SCAN_IN), .ZN(n17713) );
  OAI21_X1 U20964 ( .B1(n20930), .B2(n17714), .A(n17713), .ZN(P3_U2762) );
  AOI22_X1 U20965 ( .A1(n17722), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17715) );
  OAI21_X1 U20966 ( .B1(n17716), .B2(n17724), .A(n17715), .ZN(P3_U2763) );
  INV_X1 U20967 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U20968 ( .A1(n17722), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17717) );
  OAI21_X1 U20969 ( .B1(n17718), .B2(n17724), .A(n17717), .ZN(P3_U2764) );
  INV_X1 U20970 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17763) );
  AOI22_X1 U20971 ( .A1(P3_LWORD_REG_2__SCAN_IN), .A2(n17722), .B1(n17721), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17719) );
  OAI21_X1 U20972 ( .B1(n17763), .B2(n17724), .A(n17719), .ZN(P3_U2765) );
  AOI22_X1 U20973 ( .A1(n17722), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17720) );
  OAI21_X1 U20974 ( .B1(n17761), .B2(n17724), .A(n17720), .ZN(P3_U2766) );
  AOI22_X1 U20975 ( .A1(n17722), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17721), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17723) );
  OAI21_X1 U20976 ( .B1(n17759), .B2(n17724), .A(n17723), .ZN(P3_U2767) );
  NAND2_X1 U20977 ( .A1(n17726), .A2(n17725), .ZN(n18976) );
  INV_X2 U20978 ( .A(n17755), .ZN(n17785) );
  NOR2_X2 U20979 ( .A1(n17729), .A2(n17785), .ZN(n17779) );
  NAND2_X1 U20980 ( .A1(n17729), .A2(n17755), .ZN(n17781) );
  AOI22_X1 U20981 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17785), .ZN(n17730) );
  OAI21_X1 U20982 ( .B1(n17731), .B2(n17788), .A(n17730), .ZN(P3_U2768) );
  AOI22_X1 U20983 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17785), .ZN(n17732) );
  OAI21_X1 U20984 ( .B1(n17733), .B2(n17788), .A(n17732), .ZN(P3_U2769) );
  AOI22_X1 U20985 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17786), .B1(
        P3_EAX_REG_18__SCAN_IN), .B2(n17779), .ZN(n17734) );
  OAI21_X1 U20986 ( .B1(n17755), .B2(n20845), .A(n17734), .ZN(P3_U2770) );
  AOI22_X1 U20987 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17785), .ZN(n17735) );
  OAI21_X1 U20988 ( .B1(n17736), .B2(n17788), .A(n17735), .ZN(P3_U2771) );
  AOI22_X1 U20989 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17786), .B1(
        P3_EAX_REG_20__SCAN_IN), .B2(n17779), .ZN(n17737) );
  OAI21_X1 U20990 ( .B1(n17755), .B2(n20942), .A(n17737), .ZN(P3_U2772) );
  AOI22_X1 U20991 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17785), .ZN(n17738) );
  OAI21_X1 U20992 ( .B1(n17739), .B2(n17788), .A(n17738), .ZN(P3_U2773) );
  AOI22_X1 U20993 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17785), .ZN(n17740) );
  OAI21_X1 U20994 ( .B1(n17741), .B2(n17788), .A(n17740), .ZN(P3_U2774) );
  AOI22_X1 U20995 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17785), .ZN(n17742) );
  OAI21_X1 U20996 ( .B1(n17743), .B2(n17788), .A(n17742), .ZN(P3_U2775) );
  AOI22_X1 U20997 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17785), .ZN(n17744) );
  OAI21_X1 U20998 ( .B1(n17745), .B2(n17788), .A(n17744), .ZN(P3_U2776) );
  AOI22_X1 U20999 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17785), .ZN(n17746) );
  OAI21_X1 U21000 ( .B1(n17747), .B2(n17788), .A(n17746), .ZN(P3_U2777) );
  AOI22_X1 U21001 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17785), .ZN(n17748) );
  OAI21_X1 U21002 ( .B1(n17749), .B2(n17788), .A(n17748), .ZN(P3_U2778) );
  AOI22_X1 U21003 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17785), .ZN(n17750) );
  OAI21_X1 U21004 ( .B1(n17751), .B2(n17788), .A(n17750), .ZN(P3_U2779) );
  AOI22_X1 U21005 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17785), .ZN(n17752) );
  OAI21_X1 U21006 ( .B1(n17753), .B2(n17788), .A(n17752), .ZN(P3_U2780) );
  AOI22_X1 U21007 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17786), .B1(
        P3_EAX_REG_29__SCAN_IN), .B2(n17779), .ZN(n17754) );
  OAI21_X1 U21008 ( .B1(n17755), .B2(n20754), .A(n17754), .ZN(P3_U2781) );
  AOI22_X1 U21009 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17786), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17785), .ZN(n17756) );
  OAI21_X1 U21010 ( .B1(n17757), .B2(n17788), .A(n17756), .ZN(P3_U2782) );
  AOI22_X1 U21011 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17786), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17785), .ZN(n17758) );
  OAI21_X1 U21012 ( .B1(n17759), .B2(n17788), .A(n17758), .ZN(P3_U2783) );
  AOI22_X1 U21013 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17786), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17785), .ZN(n17760) );
  OAI21_X1 U21014 ( .B1(n17761), .B2(n17788), .A(n17760), .ZN(P3_U2784) );
  AOI22_X1 U21015 ( .A1(P3_LWORD_REG_2__SCAN_IN), .A2(n17785), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n17786), .ZN(n17762) );
  OAI21_X1 U21016 ( .B1(n17763), .B2(n17788), .A(n17762), .ZN(P3_U2785) );
  AOI22_X1 U21017 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17785), .ZN(n17764) );
  OAI21_X1 U21018 ( .B1(n18495), .B2(n17781), .A(n17764), .ZN(P3_U2786) );
  AOI22_X1 U21019 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17785), .ZN(n17765) );
  OAI21_X1 U21020 ( .B1(n18500), .B2(n17781), .A(n17765), .ZN(P3_U2787) );
  AOI22_X1 U21021 ( .A1(P3_LWORD_REG_5__SCAN_IN), .A2(n17785), .B1(
        P3_EAX_REG_5__SCAN_IN), .B2(n17779), .ZN(n17766) );
  OAI21_X1 U21022 ( .B1(n18505), .B2(n17781), .A(n17766), .ZN(P3_U2788) );
  AOI22_X1 U21023 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17785), .ZN(n17767) );
  OAI21_X1 U21024 ( .B1(n18509), .B2(n17781), .A(n17767), .ZN(P3_U2789) );
  AOI22_X1 U21025 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17785), .ZN(n17768) );
  OAI21_X1 U21026 ( .B1(n18513), .B2(n17781), .A(n17768), .ZN(P3_U2790) );
  AOI22_X1 U21027 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17786), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17785), .ZN(n17769) );
  OAI21_X1 U21028 ( .B1(n17770), .B2(n17788), .A(n17769), .ZN(P3_U2791) );
  AOI22_X1 U21029 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17785), .ZN(n17771) );
  OAI21_X1 U21030 ( .B1(n17772), .B2(n17781), .A(n17771), .ZN(P3_U2792) );
  AOI22_X1 U21031 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17786), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17785), .ZN(n17773) );
  OAI21_X1 U21032 ( .B1(n17774), .B2(n17788), .A(n17773), .ZN(P3_U2793) );
  AOI22_X1 U21033 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17785), .ZN(n17775) );
  OAI21_X1 U21034 ( .B1(n17776), .B2(n17781), .A(n17775), .ZN(P3_U2794) );
  AOI22_X1 U21035 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17779), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17785), .ZN(n17777) );
  OAI21_X1 U21036 ( .B1(n17778), .B2(n17781), .A(n17777), .ZN(P3_U2795) );
  AOI22_X1 U21037 ( .A1(P3_LWORD_REG_13__SCAN_IN), .A2(n17785), .B1(
        P3_EAX_REG_13__SCAN_IN), .B2(n17779), .ZN(n17780) );
  OAI21_X1 U21038 ( .B1(n17782), .B2(n17781), .A(n17780), .ZN(P3_U2796) );
  AOI22_X1 U21039 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17786), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17785), .ZN(n17783) );
  OAI21_X1 U21040 ( .B1(n17784), .B2(n17788), .A(n17783), .ZN(P3_U2797) );
  AOI22_X1 U21041 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17786), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17785), .ZN(n17787) );
  OAI21_X1 U21042 ( .B1(n17789), .B2(n17788), .A(n17787), .ZN(P3_U2798) );
  NAND2_X1 U21043 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17790), .ZN(
        n17808) );
  OAI21_X1 U21044 ( .B1(n17791), .B2(n18163), .A(n18162), .ZN(n17792) );
  AOI21_X1 U21045 ( .B1(n18121), .B2(n17796), .A(n17792), .ZN(n17827) );
  OAI21_X1 U21046 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17906), .A(
        n17827), .ZN(n17811) );
  AOI211_X1 U21047 ( .C1(n17795), .C2(n17794), .A(n17793), .B(n18042), .ZN(
        n17802) );
  NOR2_X1 U21048 ( .A1(n18005), .A2(n17796), .ZN(n17813) );
  OAI211_X1 U21049 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17813), .B(n17797), .ZN(n17798) );
  OAI211_X1 U21050 ( .C1(n18016), .C2(n17800), .A(n17799), .B(n17798), .ZN(
        n17801) );
  AOI211_X1 U21051 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17811), .A(
        n17802), .B(n17801), .ZN(n17807) );
  NOR2_X1 U21052 ( .A1(n18154), .A2(n18034), .ZN(n17912) );
  INV_X1 U21053 ( .A(n17912), .ZN(n17805) );
  AOI22_X1 U21054 ( .A1(n18034), .A2(n17804), .B1(n18154), .B2(n17803), .ZN(
        n17822) );
  NAND2_X1 U21055 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17822), .ZN(
        n17815) );
  NAND3_X1 U21056 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17805), .A3(
        n17815), .ZN(n17806) );
  OAI211_X1 U21057 ( .C1(n17814), .C2(n17808), .A(n17807), .B(n17806), .ZN(
        P3_U2802) );
  OAI22_X1 U21058 ( .A1(n18455), .A2(n19062), .B1(n18016), .B2(n17809), .ZN(
        n17810) );
  AOI221_X1 U21059 ( .B1(n17813), .B2(n17812), .C1(n17811), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17810), .ZN(n17818) );
  INV_X1 U21060 ( .A(n17814), .ZN(n17816) );
  OAI21_X1 U21061 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17816), .A(
        n17815), .ZN(n17817) );
  OAI211_X1 U21062 ( .C1(n17819), .C2(n18042), .A(n17818), .B(n17817), .ZN(
        P3_U2803) );
  AOI21_X1 U21063 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17821), .A(
        n17820), .ZN(n18174) );
  INV_X1 U21064 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18170) );
  INV_X1 U21065 ( .A(n17822), .ZN(n17829) );
  AOI21_X1 U21066 ( .B1(n18862), .B2(n17823), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17826) );
  OAI21_X1 U21067 ( .B1(n17943), .B2(n17944), .A(n17824), .ZN(n17825) );
  NAND2_X1 U21068 ( .A1(n9731), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18172) );
  OAI211_X1 U21069 ( .C1(n17827), .C2(n17826), .A(n17825), .B(n18172), .ZN(
        n17828) );
  AOI221_X1 U21070 ( .B1(n17830), .B2(n18170), .C1(n17829), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17828), .ZN(n17831) );
  OAI21_X1 U21071 ( .B1(n18174), .B2(n18042), .A(n17831), .ZN(P3_U2804) );
  OAI21_X1 U21072 ( .B1(n17997), .B2(n17833), .A(n17832), .ZN(n17834) );
  XOR2_X1 U21073 ( .A(n17834), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18185) );
  NAND2_X1 U21074 ( .A1(n18862), .A2(n17837), .ZN(n17860) );
  OAI211_X1 U21075 ( .C1(n17835), .C2(n18163), .A(n18162), .B(n17860), .ZN(
        n17863) );
  AOI21_X1 U21076 ( .B1(n17944), .B2(n17836), .A(n17863), .ZN(n17856) );
  NOR2_X1 U21077 ( .A1(n18005), .A2(n17837), .ZN(n17852) );
  OAI211_X1 U21078 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17852), .B(n17838), .ZN(n17839) );
  NAND2_X1 U21079 ( .A1(n9731), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n18189) );
  OAI211_X1 U21080 ( .C1(n17856), .C2(n17840), .A(n17839), .B(n18189), .ZN(
        n17841) );
  AOI21_X1 U21081 ( .B1(n17943), .B2(n17842), .A(n17841), .ZN(n17848) );
  AOI21_X1 U21082 ( .B1(n18191), .B2(n17844), .A(n17843), .ZN(n18188) );
  AOI21_X1 U21083 ( .B1(n18191), .B2(n17846), .A(n17845), .ZN(n18184) );
  AOI22_X1 U21084 ( .A1(n18154), .A2(n18188), .B1(n18034), .B2(n18184), .ZN(
        n17847) );
  OAI211_X1 U21085 ( .C1(n18042), .C2(n18185), .A(n17848), .B(n17847), .ZN(
        P3_U2805) );
  AOI21_X1 U21086 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17850), .A(
        n17849), .ZN(n18205) );
  NOR2_X1 U21087 ( .A1(n17851), .A2(n17967), .ZN(n17858) );
  OAI22_X1 U21088 ( .A1(n18192), .A2(n18079), .B1(n9790), .B2(n18167), .ZN(
        n17873) );
  AOI22_X1 U21089 ( .A1(n17853), .A2(n17943), .B1(n17852), .B2(n17855), .ZN(
        n17854) );
  NAND2_X1 U21090 ( .A1(n9731), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n18203) );
  OAI211_X1 U21091 ( .C1(n17856), .C2(n17855), .A(n17854), .B(n18203), .ZN(
        n17857) );
  AOI221_X1 U21092 ( .B1(n17858), .B2(n9895), .C1(n17873), .C2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n17857), .ZN(n17859) );
  OAI21_X1 U21093 ( .B1(n18205), .B2(n18042), .A(n17859), .ZN(P3_U2806) );
  INV_X1 U21094 ( .A(n17860), .ZN(n17861) );
  AOI22_X1 U21095 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17863), .B1(
        n17862), .B2(n17861), .ZN(n17877) );
  INV_X1 U21096 ( .A(n18285), .ZN(n17866) );
  NOR2_X1 U21097 ( .A1(n9790), .A2(n18167), .ZN(n17865) );
  INV_X1 U21098 ( .A(n18286), .ZN(n17977) );
  NOR2_X1 U21099 ( .A1(n18192), .A2(n18079), .ZN(n17864) );
  AOI22_X1 U21100 ( .A1(n17866), .A2(n17865), .B1(n17977), .B2(n17864), .ZN(
        n17871) );
  INV_X1 U21101 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18196) );
  OAI21_X1 U21102 ( .B1(n17938), .B2(n17867), .A(n17887), .ZN(n17868) );
  OAI211_X1 U21103 ( .C1(n18075), .C2(n18228), .A(n17913), .B(n17868), .ZN(
        n17869) );
  XNOR2_X1 U21104 ( .A(n18196), .B(n17869), .ZN(n18211) );
  OAI22_X1 U21105 ( .A1(n17871), .A2(n17870), .B1(n18042), .B2(n18211), .ZN(
        n17872) );
  AOI21_X1 U21106 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17873), .A(
        n17872), .ZN(n17876) );
  NAND2_X1 U21107 ( .A1(n18444), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18210) );
  OAI21_X1 U21108 ( .B1(n17943), .B2(n17944), .A(n17874), .ZN(n17875) );
  NAND4_X1 U21109 ( .A1(n17877), .A2(n17876), .A3(n18210), .A4(n17875), .ZN(
        P3_U2807) );
  AOI21_X1 U21110 ( .B1(n17882), .B2(n18121), .A(n18119), .ZN(n17878) );
  INV_X1 U21111 ( .A(n17878), .ZN(n17879) );
  AOI21_X1 U21112 ( .B1(n18002), .B2(n17880), .A(n17879), .ZN(n17909) );
  OAI21_X1 U21113 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17906), .A(
        n17909), .ZN(n17897) );
  AOI22_X1 U21114 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17897), .B1(
        n17943), .B2(n17881), .ZN(n17893) );
  NOR2_X1 U21115 ( .A1(n18005), .A2(n17882), .ZN(n17899) );
  AOI21_X1 U21116 ( .B1(n17898), .B2(n17884), .A(n17883), .ZN(n17885) );
  AOI22_X1 U21117 ( .A1(n9731), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n17899), 
        .B2(n17885), .ZN(n17892) );
  NOR2_X1 U21118 ( .A1(n17939), .A2(n17888), .ZN(n18217) );
  AOI22_X1 U21119 ( .A1(n18034), .A2(n18286), .B1(n18154), .B2(n18285), .ZN(
        n17966) );
  OAI21_X1 U21120 ( .B1(n17912), .B2(n18217), .A(n17966), .ZN(n17903) );
  AOI221_X1 U21121 ( .B1(n17888), .B2(n17887), .C1(n17900), .C2(n17887), .A(
        n17886), .ZN(n17889) );
  XOR2_X1 U21122 ( .A(n17889), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n18212) );
  AOI22_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17903), .B1(
        n18076), .B2(n18212), .ZN(n17891) );
  NAND3_X1 U21124 ( .A1(n17950), .A2(n18217), .A3(n18228), .ZN(n17890) );
  NAND4_X1 U21125 ( .A1(n17893), .A2(n17892), .A3(n17891), .A4(n17890), .ZN(
        P3_U2808) );
  NAND2_X1 U21126 ( .A1(n18235), .A2(n18219), .ZN(n18239) );
  NAND2_X1 U21127 ( .A1(n18260), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18233) );
  INV_X1 U21128 ( .A(n17894), .ZN(n17895) );
  OAI22_X1 U21129 ( .A1(n18455), .A2(n19051), .B1(n18016), .B2(n17895), .ZN(
        n17896) );
  AOI221_X1 U21130 ( .B1(n17899), .B2(n17898), .C1(n17897), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17896), .ZN(n17905) );
  INV_X1 U21131 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17942) );
  NOR3_X1 U21132 ( .A1(n17942), .A2(n17997), .A3(n17900), .ZN(n17923) );
  AOI22_X1 U21133 ( .A1(n18235), .A2(n17923), .B1(n17938), .B2(n17901), .ZN(
        n17902) );
  XOR2_X1 U21134 ( .A(n18219), .B(n17902), .Z(n18231) );
  AOI22_X1 U21135 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17903), .B1(
        n18076), .B2(n18231), .ZN(n17904) );
  OAI211_X1 U21136 ( .C1(n18239), .C2(n17929), .A(n17905), .B(n17904), .ZN(
        P3_U2809) );
  OR2_X1 U21137 ( .A1(n17925), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n18250) );
  AOI21_X1 U21138 ( .B1(n18862), .B2(n17907), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17908) );
  OAI22_X1 U21139 ( .A1(n17909), .A2(n17908), .B1(n18455), .B2(n19049), .ZN(
        n17910) );
  AOI221_X1 U21140 ( .B1(n17943), .B2(n17911), .C1(n17944), .C2(n17911), .A(
        n17910), .ZN(n17916) );
  NAND3_X1 U21141 ( .A1(n18260), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18214) );
  INV_X1 U21142 ( .A(n18214), .ZN(n18243) );
  OAI21_X1 U21143 ( .B1(n17912), .B2(n18243), .A(n17966), .ZN(n17926) );
  OAI221_X1 U21144 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17936), 
        .C1(n17925), .C2(n17923), .A(n17913), .ZN(n17914) );
  XNOR2_X1 U21145 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17914), .ZN(
        n18240) );
  AOI22_X1 U21146 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17926), .B1(
        n18076), .B2(n18240), .ZN(n17915) );
  OAI211_X1 U21147 ( .C1(n18250), .C2(n17929), .A(n17916), .B(n17915), .ZN(
        P3_U2810) );
  AOI21_X1 U21148 ( .B1(n18121), .B2(n17918), .A(n18119), .ZN(n17953) );
  OAI21_X1 U21149 ( .B1(n17917), .B2(n18163), .A(n17953), .ZN(n17933) );
  NOR2_X1 U21150 ( .A1(n18005), .A2(n17918), .ZN(n17935) );
  OAI211_X1 U21151 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17935), .B(n17919), .ZN(n17920) );
  NAND2_X1 U21152 ( .A1(n18444), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18253) );
  OAI211_X1 U21153 ( .C1(n18016), .C2(n17921), .A(n17920), .B(n18253), .ZN(
        n17922) );
  AOI21_X1 U21154 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17933), .A(
        n17922), .ZN(n17928) );
  AOI21_X1 U21155 ( .B1(n17936), .B2(n17938), .A(n17923), .ZN(n17924) );
  XOR2_X1 U21156 ( .A(n17925), .B(n17924), .Z(n18251) );
  AOI22_X1 U21157 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17926), .B1(
        n18076), .B2(n18251), .ZN(n17927) );
  OAI211_X1 U21158 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17929), .A(
        n17928), .B(n17927), .ZN(P3_U2811) );
  INV_X1 U21159 ( .A(n17966), .ZN(n17930) );
  AOI21_X1 U21160 ( .B1(n17950), .B2(n17939), .A(n17930), .ZN(n17948) );
  OAI22_X1 U21161 ( .A1(n18455), .A2(n19045), .B1(n18016), .B2(n17931), .ZN(
        n17932) );
  AOI221_X1 U21162 ( .B1(n17935), .B2(n17934), .C1(n17933), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17932), .ZN(n17941) );
  AOI21_X1 U21163 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18075), .A(
        n17936), .ZN(n17937) );
  XOR2_X1 U21164 ( .A(n17938), .B(n17937), .Z(n18267) );
  NOR2_X1 U21165 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17939), .ZN(
        n18266) );
  AOI22_X1 U21166 ( .A1(n18076), .A2(n18267), .B1(n17950), .B2(n18266), .ZN(
        n17940) );
  OAI211_X1 U21167 ( .C1(n17948), .C2(n17942), .A(n17941), .B(n17940), .ZN(
        P3_U2812) );
  AOI21_X1 U21168 ( .B1(n9845), .B2(n18862), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17954) );
  AOI22_X1 U21169 ( .A1(n9731), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n17945), 
        .B2(n18156), .ZN(n17952) );
  NOR2_X1 U21170 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18280), .ZN(
        n18270) );
  AOI21_X1 U21171 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17947), .A(
        n17946), .ZN(n18274) );
  INV_X1 U21172 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18261) );
  OAI22_X1 U21173 ( .A1(n18274), .A2(n18042), .B1(n17948), .B2(n18261), .ZN(
        n17949) );
  AOI21_X1 U21174 ( .B1(n17950), .B2(n18270), .A(n17949), .ZN(n17951) );
  OAI211_X1 U21175 ( .C1(n17954), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2813) );
  OAI21_X1 U21176 ( .B1(n17997), .B2(n17956), .A(n17955), .ZN(n17957) );
  XOR2_X1 U21177 ( .A(n17957), .B(n18280), .Z(n18282) );
  AOI21_X1 U21178 ( .B1(n18121), .B2(n17959), .A(n18119), .ZN(n17988) );
  OAI21_X1 U21179 ( .B1(n17958), .B2(n18163), .A(n17988), .ZN(n17970) );
  AOI22_X1 U21180 ( .A1(n9731), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17970), .ZN(n17962) );
  NOR2_X1 U21181 ( .A1(n18005), .A2(n17959), .ZN(n17972) );
  OAI211_X1 U21182 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17972), .B(n17960), .ZN(n17961) );
  OAI211_X1 U21183 ( .C1(n18016), .C2(n17963), .A(n17962), .B(n17961), .ZN(
        n17964) );
  AOI21_X1 U21184 ( .B1(n18076), .B2(n18282), .A(n17964), .ZN(n17965) );
  OAI221_X1 U21185 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17967), 
        .C1(n18280), .C2(n17966), .A(n17965), .ZN(P3_U2814) );
  NOR2_X1 U21186 ( .A1(n9783), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18293) );
  NAND2_X1 U21187 ( .A1(n18154), .A2(n18285), .ZN(n17982) );
  NAND2_X1 U21188 ( .A1(n9731), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18296) );
  OAI21_X1 U21189 ( .B1(n18016), .B2(n17968), .A(n18296), .ZN(n17969) );
  AOI221_X1 U21190 ( .B1(n17972), .B2(n17971), .C1(n17970), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17969), .ZN(n17981) );
  NOR2_X1 U21191 ( .A1(n17997), .A2(n12434), .ZN(n18057) );
  INV_X1 U21192 ( .A(n18057), .ZN(n18022) );
  NOR3_X1 U21193 ( .A1(n18330), .A2(n18336), .A3(n18022), .ZN(n17985) );
  INV_X1 U21194 ( .A(n17973), .ZN(n17974) );
  NAND2_X1 U21195 ( .A1(n17974), .A2(n17997), .ZN(n18021) );
  INV_X1 U21196 ( .A(n18021), .ZN(n17984) );
  AOI22_X1 U21197 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17985), .B1(
        n17992), .B2(n17984), .ZN(n17975) );
  NAND2_X1 U21198 ( .A1(n18299), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17983) );
  INV_X1 U21199 ( .A(n17983), .ZN(n18317) );
  NOR2_X1 U21200 ( .A1(n17975), .A2(n18317), .ZN(n17976) );
  XOR2_X1 U21201 ( .A(n17976), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n18294) );
  NOR2_X1 U21202 ( .A1(n17977), .A2(n18079), .ZN(n17979) );
  OR2_X1 U21203 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18287), .ZN(
        n17978) );
  AOI22_X1 U21204 ( .A1(n18076), .A2(n18294), .B1(n17979), .B2(n17978), .ZN(
        n17980) );
  OAI211_X1 U21205 ( .C1(n18293), .C2(n17982), .A(n17981), .B(n17980), .ZN(
        P3_U2815) );
  OAI221_X1 U21206 ( .B1(n17985), .B2(n17984), .C1(n17985), .C2(n18299), .A(
        n17983), .ZN(n17986) );
  XOR2_X1 U21207 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n17986), .Z(
        n18316) );
  AOI21_X1 U21208 ( .B1(n18862), .B2(n17987), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17989) );
  OAI22_X1 U21209 ( .A1(n18146), .A2(n17990), .B1(n17989), .B2(n17988), .ZN(
        n17991) );
  AOI21_X1 U21210 ( .B1(n18444), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17991), 
        .ZN(n17996) );
  NOR2_X1 U21211 ( .A1(n18340), .A2(n18319), .ZN(n18011) );
  INV_X1 U21212 ( .A(n18011), .ZN(n17993) );
  AOI211_X1 U21213 ( .C1(n18304), .C2(n17993), .A(n17992), .B(n9783), .ZN(
        n18312) );
  AOI21_X1 U21214 ( .B1(n18304), .B2(n17994), .A(n18287), .ZN(n18308) );
  AOI22_X1 U21215 ( .A1(n18154), .A2(n18312), .B1(n18034), .B2(n18308), .ZN(
        n17995) );
  OAI211_X1 U21216 ( .C1(n18042), .C2(n18316), .A(n17996), .B(n17995), .ZN(
        P3_U2816) );
  AOI22_X1 U21217 ( .A1(n17998), .A2(n18329), .B1(n18336), .B2(n17997), .ZN(
        n17999) );
  NOR2_X1 U21218 ( .A1(n17999), .A2(n10158), .ZN(n18000) );
  XOR2_X1 U21219 ( .A(n18000), .B(n18299), .Z(n18327) );
  AOI22_X1 U21220 ( .A1(n18002), .A2(n18001), .B1(n18121), .B2(n18004), .ZN(
        n18003) );
  NAND2_X1 U21221 ( .A1(n18003), .A2(n18162), .ZN(n18018) );
  NOR2_X1 U21222 ( .A1(n18005), .A2(n18004), .ZN(n18020) );
  OAI211_X1 U21223 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18020), .B(n18006), .ZN(n18008) );
  NAND2_X1 U21224 ( .A1(n18444), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n18007) );
  OAI211_X1 U21225 ( .C1(n18016), .C2(n18009), .A(n18008), .B(n18007), .ZN(
        n18010) );
  AOI21_X1 U21226 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18018), .A(
        n18010), .ZN(n18013) );
  OAI22_X1 U21227 ( .A1(n18321), .A2(n18079), .B1(n18011), .B2(n18167), .ZN(
        n18014) );
  NOR2_X1 U21228 ( .A1(n18040), .A2(n18330), .ZN(n18024) );
  AOI22_X1 U21229 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18014), .B1(
        n18317), .B2(n18024), .ZN(n18012) );
  OAI211_X1 U21230 ( .C1(n18042), .C2(n18327), .A(n18013), .B(n18012), .ZN(
        P3_U2817) );
  INV_X1 U21231 ( .A(n18014), .ZN(n18027) );
  INV_X1 U21232 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n18019) );
  INV_X1 U21233 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19034) );
  OAI22_X1 U21234 ( .A1(n18455), .A2(n19034), .B1(n18016), .B2(n18015), .ZN(
        n18017) );
  AOI221_X1 U21235 ( .B1(n18020), .B2(n18019), .C1(n18018), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n18017), .ZN(n18026) );
  OAI21_X1 U21236 ( .B1(n18330), .B2(n18022), .A(n18021), .ZN(n18023) );
  XOR2_X1 U21237 ( .A(n18023), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18328) );
  AOI22_X1 U21238 ( .A1(n18076), .A2(n18328), .B1(n18024), .B2(n18336), .ZN(
        n18025) );
  OAI211_X1 U21239 ( .C1(n18027), .C2(n18336), .A(n18026), .B(n18025), .ZN(
        P3_U2818) );
  NAND2_X1 U21240 ( .A1(n18344), .A2(n12430), .ZN(n18350) );
  NOR3_X1 U21241 ( .A1(n18826), .A2(n18095), .A3(n18028), .ZN(n18098) );
  NAND2_X1 U21242 ( .A1(n18067), .A2(n18098), .ZN(n18053) );
  NOR2_X1 U21243 ( .A1(n18052), .A2(n18053), .ZN(n18050) );
  NAND2_X1 U21244 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18050), .ZN(
        n18047) );
  INV_X1 U21245 ( .A(n18051), .ZN(n18157) );
  NAND2_X1 U21246 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18157), .ZN(
        n18029) );
  AOI22_X1 U21247 ( .A1(n18030), .A2(n18098), .B1(n18047), .B2(n18029), .ZN(
        n18032) );
  NOR2_X1 U21248 ( .A1(n20772), .A2(n18455), .ZN(n18031) );
  AOI211_X1 U21249 ( .C1(n18033), .C2(n18156), .A(n18032), .B(n18031), .ZN(
        n18039) );
  AOI22_X1 U21250 ( .A1(n18340), .A2(n18154), .B1(n18034), .B2(n18338), .ZN(
        n18063) );
  OAI21_X1 U21251 ( .B1(n18344), .B2(n18040), .A(n18063), .ZN(n18046) );
  NOR2_X1 U21252 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18036) );
  NOR2_X1 U21253 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18035), .ZN(
        n18058) );
  AOI22_X1 U21254 ( .A1(n18344), .A2(n18057), .B1(n18036), .B2(n18058), .ZN(
        n18037) );
  XOR2_X1 U21255 ( .A(n12430), .B(n18037), .Z(n18337) );
  AOI22_X1 U21256 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18046), .B1(
        n18076), .B2(n18337), .ZN(n18038) );
  OAI211_X1 U21257 ( .C1(n18040), .C2(n18350), .A(n18039), .B(n18038), .ZN(
        P3_U2819) );
  OAI21_X1 U21258 ( .B1(n18040), .B2(n18365), .A(n18352), .ZN(n18045) );
  AOI22_X1 U21259 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18057), .B1(
        n18058), .B2(n18365), .ZN(n18041) );
  XOR2_X1 U21260 ( .A(n18041), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18359) );
  OAI22_X1 U21261 ( .A1(n18146), .A2(n18043), .B1(n18359), .B2(n18042), .ZN(
        n18044) );
  AOI21_X1 U21262 ( .B1(n18046), .B2(n18045), .A(n18044), .ZN(n18049) );
  OAI211_X1 U21263 ( .C1(n18050), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n18157), .B(n18047), .ZN(n18048) );
  OAI211_X1 U21264 ( .C1(n19032), .C2(n18455), .A(n18049), .B(n18048), .ZN(
        P3_U2820) );
  AOI211_X1 U21265 ( .C1(n18053), .C2(n18052), .A(n18051), .B(n18050), .ZN(
        n18055) );
  NOR2_X1 U21266 ( .A1(n18455), .A2(n19029), .ZN(n18054) );
  AOI211_X1 U21267 ( .C1(n18056), .C2(n18156), .A(n18055), .B(n18054), .ZN(
        n18062) );
  NOR2_X1 U21268 ( .A1(n18058), .A2(n18057), .ZN(n18059) );
  XOR2_X1 U21269 ( .A(n18059), .B(n18365), .Z(n18362) );
  AOI22_X1 U21270 ( .A1(n18076), .A2(n18362), .B1(n18365), .B2(n18060), .ZN(
        n18061) );
  OAI211_X1 U21271 ( .C1(n18063), .C2(n18365), .A(n18062), .B(n18061), .ZN(
        P3_U2821) );
  NAND2_X1 U21272 ( .A1(n18064), .A2(n12434), .ZN(n18375) );
  INV_X1 U21273 ( .A(n18121), .ZN(n18065) );
  OAI21_X1 U21274 ( .B1(n18066), .B2(n18065), .A(n18162), .ZN(n18082) );
  NAND2_X1 U21275 ( .A1(n18066), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18068) );
  AOI211_X1 U21276 ( .C1(n18069), .C2(n18068), .A(n18067), .B(n18826), .ZN(
        n18072) );
  NAND2_X1 U21277 ( .A1(n18444), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18380) );
  OAI21_X1 U21278 ( .B1(n18146), .B2(n18070), .A(n18380), .ZN(n18071) );
  AOI211_X1 U21279 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18082), .A(
        n18072), .B(n18071), .ZN(n18078) );
  AOI21_X1 U21280 ( .B1(n18074), .B2(n20850), .A(n18073), .ZN(n18373) );
  XOR2_X1 U21281 ( .A(n18075), .B(n18375), .Z(n18377) );
  AOI22_X1 U21282 ( .A1(n18154), .A2(n18373), .B1(n18076), .B2(n18377), .ZN(
        n18077) );
  OAI211_X1 U21283 ( .C1(n18079), .C2(n18375), .A(n18078), .B(n18077), .ZN(
        P3_U2822) );
  INV_X1 U21284 ( .A(n18131), .ZN(n18166) );
  OAI21_X1 U21285 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18081), .A(
        n18080), .ZN(n18392) );
  NOR2_X1 U21286 ( .A1(n18455), .A2(n19025), .ZN(n18383) );
  AOI221_X1 U21287 ( .B1(n18098), .B2(n18083), .C1(n18082), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18383), .ZN(n18089) );
  NAND2_X1 U21288 ( .A1(n18085), .A2(n18084), .ZN(n18086) );
  INV_X1 U21289 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18385) );
  XOR2_X1 U21290 ( .A(n18086), .B(n18385), .Z(n18389) );
  AOI22_X1 U21291 ( .A1(n18154), .A2(n18389), .B1(n18087), .B2(n18156), .ZN(
        n18088) );
  OAI211_X1 U21292 ( .C1(n18166), .C2(n18392), .A(n18089), .B(n18088), .ZN(
        P3_U2823) );
  OAI21_X1 U21293 ( .B1(n18092), .B2(n18091), .A(n18090), .ZN(n18401) );
  AOI21_X1 U21294 ( .B1(n18386), .B2(n18094), .A(n18093), .ZN(n18398) );
  NOR2_X1 U21295 ( .A1(n18826), .A2(n18095), .ZN(n18106) );
  AOI21_X1 U21296 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18157), .A(
        n18106), .ZN(n18097) );
  OAI22_X1 U21297 ( .A1(n18098), .A2(n18097), .B1(n18146), .B2(n18096), .ZN(
        n18099) );
  AOI21_X1 U21298 ( .B1(n18154), .B2(n18398), .A(n18099), .ZN(n18100) );
  NAND2_X1 U21299 ( .A1(n18444), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18399) );
  OAI211_X1 U21300 ( .C1(n18166), .C2(n18401), .A(n18100), .B(n18399), .ZN(
        P3_U2824) );
  OAI21_X1 U21301 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n18102), .A(
        n18101), .ZN(n18408) );
  AOI21_X1 U21302 ( .B1(n18105), .B2(n18104), .A(n18103), .ZN(n18405) );
  AOI22_X1 U21303 ( .A1(n9731), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18154), .B2(
        n18405), .ZN(n18111) );
  AOI221_X1 U21304 ( .B1(n18119), .B2(n20716), .C1(n18107), .C2(n20716), .A(
        n18106), .ZN(n18108) );
  AOI22_X1 U21305 ( .A1(n18109), .A2(n18156), .B1(n18108), .B2(n18157), .ZN(
        n18110) );
  OAI211_X1 U21306 ( .C1(n18166), .C2(n18408), .A(n18111), .B(n18110), .ZN(
        P3_U2825) );
  OAI21_X1 U21307 ( .B1(n18114), .B2(n18113), .A(n18112), .ZN(n18412) );
  AOI21_X1 U21308 ( .B1(n18117), .B2(n18116), .A(n18115), .ZN(n18414) );
  OAI22_X1 U21309 ( .A1(n20983), .A2(n18455), .B1(n18826), .B2(n18118), .ZN(
        n18125) );
  AOI21_X1 U21310 ( .B1(n18121), .B2(n18120), .A(n18119), .ZN(n18138) );
  OAI22_X1 U21311 ( .A1(n18146), .A2(n18123), .B1(n18122), .B2(n18138), .ZN(
        n18124) );
  AOI211_X1 U21312 ( .C1(n18154), .C2(n18414), .A(n18125), .B(n18124), .ZN(
        n18126) );
  OAI21_X1 U21313 ( .B1(n18166), .B2(n18412), .A(n18126), .ZN(P3_U2826) );
  AOI21_X1 U21314 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18162), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18139) );
  AOI21_X1 U21315 ( .B1(n18129), .B2(n18128), .A(n18127), .ZN(n18130) );
  XOR2_X1 U21316 ( .A(n18130), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18419) );
  AOI22_X1 U21317 ( .A1(n18444), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18131), 
        .B2(n18419), .ZN(n18137) );
  AOI21_X1 U21318 ( .B1(n18134), .B2(n18133), .A(n18132), .ZN(n18420) );
  AOI22_X1 U21319 ( .A1(n18154), .A2(n18420), .B1(n18135), .B2(n18156), .ZN(
        n18136) );
  OAI211_X1 U21320 ( .C1(n18139), .C2(n18138), .A(n18137), .B(n18136), .ZN(
        P3_U2827) );
  AOI21_X1 U21321 ( .B1(n18142), .B2(n18141), .A(n18140), .ZN(n18432) );
  NAND2_X1 U21322 ( .A1(n18444), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18440) );
  INV_X1 U21323 ( .A(n18440), .ZN(n18148) );
  OAI22_X1 U21324 ( .A1(n18146), .A2(n18145), .B1(n18166), .B2(n18442), .ZN(
        n18147) );
  AOI211_X1 U21325 ( .C1(n18154), .C2(n18432), .A(n18148), .B(n18147), .ZN(
        n18149) );
  OAI221_X1 U21326 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18826), .C1(
        n18150), .C2(n18162), .A(n18149), .ZN(P3_U2828) );
  OAI21_X1 U21327 ( .B1(n18152), .B2(n18160), .A(n18151), .ZN(n18450) );
  NAND2_X1 U21328 ( .A1(n19106), .A2(n18161), .ZN(n18153) );
  XNOR2_X1 U21329 ( .A(n18153), .B(n18152), .ZN(n18452) );
  AOI22_X1 U21330 ( .A1(n9731), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18154), .B2(
        n18452), .ZN(n18159) );
  AOI22_X1 U21331 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18157), .B1(
        n18156), .B2(n18155), .ZN(n18158) );
  OAI211_X1 U21332 ( .C1(n18166), .C2(n18450), .A(n18159), .B(n18158), .ZN(
        P3_U2829) );
  AOI21_X1 U21333 ( .B1(n18161), .B2(n19106), .A(n18160), .ZN(n18457) );
  INV_X1 U21334 ( .A(n18457), .ZN(n18459) );
  NAND3_X1 U21335 ( .A1(n19088), .A2(n18163), .A3(n18162), .ZN(n18164) );
  AOI22_X1 U21336 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n9731), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18164), .ZN(n18165) );
  OAI221_X1 U21337 ( .B1(n18457), .B2(n18167), .C1(n18459), .C2(n18166), .A(
        n18165), .ZN(P3_U2830) );
  OR4_X1 U21338 ( .A1(n18191), .A2(n18200), .A3(n9895), .A4(n18229), .ZN(
        n18169) );
  AOI211_X1 U21339 ( .C1(n18170), .C2(n18169), .A(n18168), .B(n18461), .ZN(
        n18171) );
  AOI21_X1 U21340 ( .B1(n18439), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n18171), .ZN(n18173) );
  OAI211_X1 U21341 ( .C1(n18174), .C2(n18358), .A(n18173), .B(n18172), .ZN(
        P3_U2836) );
  NOR2_X1 U21342 ( .A1(n18175), .A2(n18179), .ZN(n18182) );
  INV_X1 U21343 ( .A(n18176), .ZN(n18178) );
  NOR2_X1 U21344 ( .A1(n18177), .A2(n18943), .ZN(n18197) );
  AOI211_X1 U21345 ( .C1(n18963), .C2(n18179), .A(n18178), .B(n18197), .ZN(
        n18180) );
  INV_X1 U21346 ( .A(n18180), .ZN(n18181) );
  MUX2_X1 U21347 ( .A(n18182), .B(n18181), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n18183) );
  AOI21_X1 U21348 ( .B1(n18339), .B2(n18184), .A(n18183), .ZN(n18186) );
  OAI22_X1 U21349 ( .A1(n18186), .A2(n18461), .B1(n18358), .B2(n18185), .ZN(
        n18187) );
  AOI21_X1 U21350 ( .B1(n18460), .B2(n18188), .A(n18187), .ZN(n18190) );
  OAI211_X1 U21351 ( .C1(n18454), .C2(n18191), .A(n18190), .B(n18189), .ZN(
        P3_U2837) );
  OAI22_X1 U21352 ( .A1(n9790), .A2(n18193), .B1(n18192), .B2(n18376), .ZN(
        n18194) );
  AOI211_X1 U21353 ( .C1(n18426), .C2(n18195), .A(n18439), .B(n18194), .ZN(
        n18199) );
  AOI21_X1 U21354 ( .B1(n9886), .B2(n18199), .A(n9895), .ZN(n18202) );
  NOR2_X1 U21355 ( .A1(n18197), .A2(n18196), .ZN(n18198) );
  AOI21_X1 U21356 ( .B1(n18199), .B2(n18198), .A(n9731), .ZN(n18207) );
  NOR4_X1 U21357 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18200), .A3(
        n18461), .A4(n18229), .ZN(n18201) );
  AOI21_X1 U21358 ( .B1(n18202), .B2(n18207), .A(n18201), .ZN(n18204) );
  OAI211_X1 U21359 ( .C1(n18205), .C2(n18358), .A(n18204), .B(n18203), .ZN(
        P3_U2838) );
  INV_X1 U21360 ( .A(n18206), .ZN(n18208) );
  OAI221_X1 U21361 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18208), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18454), .A(n18207), .ZN(
        n18209) );
  OAI211_X1 U21362 ( .C1(n18358), .C2(n18211), .A(n18210), .B(n18209), .ZN(
        P3_U2839) );
  AOI22_X1 U21363 ( .A1(n9731), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n18378), 
        .B2(n18212), .ZN(n18227) );
  NAND2_X1 U21364 ( .A1(n18963), .A2(n18213), .ZN(n18258) );
  OAI21_X1 U21365 ( .B1(n18215), .B2(n18214), .A(n18947), .ZN(n18216) );
  OAI211_X1 U21366 ( .C1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n18943), .A(
        n18258), .B(n18216), .ZN(n18244) );
  NOR2_X1 U21367 ( .A1(n18961), .A2(n18339), .ZN(n18343) );
  OAI22_X1 U21368 ( .A1(n18930), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18343), .B2(n18217), .ZN(n18218) );
  NOR2_X1 U21369 ( .A1(n18244), .A2(n18218), .ZN(n18234) );
  AOI22_X1 U21370 ( .A1(n18961), .A2(n18285), .B1(n18339), .B2(n18286), .ZN(
        n18242) );
  AOI22_X1 U21371 ( .A1(n18963), .A2(n18220), .B1(n18351), .B2(n18219), .ZN(
        n18223) );
  OAI21_X1 U21372 ( .B1(n18228), .B2(n18928), .A(n18221), .ZN(n18222) );
  NAND4_X1 U21373 ( .A1(n18234), .A2(n18242), .A3(n18223), .A4(n18222), .ZN(
        n18224) );
  OAI211_X1 U21374 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n18225), .A(
        n18438), .B(n18224), .ZN(n18226) );
  OAI211_X1 U21375 ( .C1(n18454), .C2(n18228), .A(n18227), .B(n18226), .ZN(
        P3_U2840) );
  NOR2_X1 U21376 ( .A1(n18461), .A2(n18229), .ZN(n18230) );
  NAND2_X1 U21377 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n18230), .ZN(
        n18255) );
  AOI22_X1 U21378 ( .A1(n18444), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18378), 
        .B2(n18231), .ZN(n18238) );
  NAND2_X1 U21379 ( .A1(n18438), .A2(n18242), .ZN(n18279) );
  NOR2_X1 U21380 ( .A1(n18963), .A2(n18928), .ZN(n18443) );
  INV_X1 U21381 ( .A(n18265), .ZN(n18232) );
  NOR2_X1 U21382 ( .A1(n19106), .A2(n18275), .ZN(n18342) );
  NAND2_X1 U21383 ( .A1(n18232), .A2(n18342), .ZN(n18277) );
  OAI21_X1 U21384 ( .B1(n18277), .B2(n18233), .A(n18928), .ZN(n18241) );
  OAI211_X1 U21385 ( .C1(n18235), .C2(n18443), .A(n18234), .B(n18241), .ZN(
        n18236) );
  OAI211_X1 U21386 ( .C1(n18279), .C2(n18236), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18455), .ZN(n18237) );
  OAI211_X1 U21387 ( .C1(n18255), .C2(n18239), .A(n18238), .B(n18237), .ZN(
        P3_U2841) );
  AOI22_X1 U21388 ( .A1(n9731), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18378), 
        .B2(n18240), .ZN(n18249) );
  OAI211_X1 U21389 ( .C1(n18243), .C2(n18343), .A(n18242), .B(n18241), .ZN(
        n18245) );
  NOR3_X1 U21390 ( .A1(n18245), .A2(n18461), .A3(n18244), .ZN(n18246) );
  NOR2_X1 U21391 ( .A1(n18246), .A2(n9731), .ZN(n18252) );
  NOR3_X1 U21392 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18443), .A3(
        n19143), .ZN(n18247) );
  OAI21_X1 U21393 ( .B1(n18252), .B2(n18247), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18248) );
  OAI211_X1 U21394 ( .C1(n18255), .C2(n18250), .A(n18249), .B(n18248), .ZN(
        P3_U2842) );
  AOI22_X1 U21395 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18252), .B1(
        n18378), .B2(n18251), .ZN(n18254) );
  OAI211_X1 U21396 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18255), .A(
        n18254), .B(n18253), .ZN(P3_U2843) );
  NAND3_X1 U21397 ( .A1(n18256), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18434), .ZN(n18257) );
  AOI21_X1 U21398 ( .B1(n18426), .B2(n18257), .A(n18279), .ZN(n18259) );
  OAI211_X1 U21399 ( .C1(n18260), .C2(n18343), .A(n18259), .B(n18258), .ZN(
        n18271) );
  OAI221_X1 U21400 ( .B1(n18271), .B2(n18261), .C1(n18271), .C2(n18426), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n18269) );
  NAND2_X1 U21401 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18409) );
  OAI22_X1 U21402 ( .A1(n18410), .A2(n18943), .B1(n18409), .B2(n18429), .ZN(
        n18422) );
  NAND2_X1 U21403 ( .A1(n18262), .A2(n18422), .ZN(n18384) );
  NOR2_X1 U21404 ( .A1(n18263), .A2(n18384), .ZN(n18300) );
  NOR2_X1 U21405 ( .A1(n18265), .A2(n18366), .ZN(n18281) );
  AOI22_X1 U21406 ( .A1(n18378), .A2(n18267), .B1(n18281), .B2(n18266), .ZN(
        n18268) );
  OAI221_X1 U21407 ( .B1(n18444), .B2(n18269), .C1(n18455), .C2(n19045), .A(
        n18268), .ZN(P3_U2844) );
  AOI22_X1 U21408 ( .A1(n9731), .A2(P3_REIP_REG_17__SCAN_IN), .B1(n18281), 
        .B2(n18270), .ZN(n18273) );
  NAND3_X1 U21409 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18455), .A3(
        n18271), .ZN(n18272) );
  OAI211_X1 U21410 ( .C1(n18274), .C2(n18358), .A(n18273), .B(n18272), .ZN(
        P3_U2845) );
  AOI22_X1 U21411 ( .A1(n18963), .A2(n18276), .B1(n18947), .B2(n18275), .ZN(
        n18302) );
  OAI21_X1 U21412 ( .B1(n18298), .B2(n18928), .A(n18277), .ZN(n18278) );
  OAI211_X1 U21413 ( .C1(n18323), .C2(n18289), .A(n18302), .B(n18278), .ZN(
        n18288) );
  OAI221_X1 U21414 ( .B1(n18279), .B2(n18370), .C1(n18279), .C2(n18288), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18284) );
  AOI22_X1 U21415 ( .A1(n18282), .A2(n18378), .B1(n18281), .B2(n18280), .ZN(
        n18283) );
  OAI221_X1 U21416 ( .B1(n9731), .B2(n18284), .C1(n18455), .C2(n19041), .A(
        n18283), .ZN(P3_U2846) );
  NAND2_X1 U21417 ( .A1(n18961), .A2(n18285), .ZN(n18292) );
  OAI211_X1 U21418 ( .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18287), .A(
        n18339), .B(n18286), .ZN(n18291) );
  OAI221_X1 U21419 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18289), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18300), .A(n18288), .ZN(
        n18290) );
  OAI211_X1 U21420 ( .C1(n18293), .C2(n18292), .A(n18291), .B(n18290), .ZN(
        n18295) );
  AOI22_X1 U21421 ( .A1(n18438), .A2(n18295), .B1(n18378), .B2(n18294), .ZN(
        n18297) );
  OAI211_X1 U21422 ( .C1(n18454), .C2(n18298), .A(n18297), .B(n18296), .ZN(
        P3_U2847) );
  AOI22_X1 U21423 ( .A1(n18444), .A2(P3_REIP_REG_14__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18439), .ZN(n18315) );
  NOR2_X1 U21424 ( .A1(n18319), .A2(n18299), .ZN(n18301) );
  AOI21_X1 U21425 ( .B1(n18301), .B2(n18300), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18311) );
  INV_X1 U21426 ( .A(n18302), .ZN(n18361) );
  OAI21_X1 U21427 ( .B1(n18304), .B2(n18947), .A(n18303), .ZN(n18306) );
  NAND2_X1 U21428 ( .A1(n18329), .A2(n18342), .ZN(n18305) );
  NAND2_X1 U21429 ( .A1(n18928), .A2(n18305), .ZN(n18322) );
  OAI211_X1 U21430 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18443), .A(
        n18306), .B(n18322), .ZN(n18307) );
  AOI211_X1 U21431 ( .C1(n18963), .C2(n18319), .A(n18361), .B(n18307), .ZN(
        n18310) );
  INV_X1 U21432 ( .A(n18308), .ZN(n18309) );
  OAI22_X1 U21433 ( .A1(n18311), .A2(n18310), .B1(n18376), .B2(n18309), .ZN(
        n18313) );
  AOI22_X1 U21434 ( .A1(n18438), .A2(n18313), .B1(n18460), .B2(n18312), .ZN(
        n18314) );
  OAI211_X1 U21435 ( .C1(n18358), .C2(n18316), .A(n18315), .B(n18314), .ZN(
        P3_U2848) );
  NOR2_X1 U21436 ( .A1(n18330), .A2(n18366), .ZN(n18318) );
  AOI22_X1 U21437 ( .A1(n18444), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18318), 
        .B2(n18317), .ZN(n18326) );
  AOI21_X1 U21438 ( .B1(n18351), .B2(n18330), .A(n18361), .ZN(n18346) );
  OAI21_X1 U21439 ( .B1(n18340), .B2(n18319), .A(n18961), .ZN(n18320) );
  OAI211_X1 U21440 ( .C1(n18321), .C2(n18376), .A(n18346), .B(n18320), .ZN(
        n18332) );
  OAI211_X1 U21441 ( .C1(n18323), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18322), .B(n18454), .ZN(n18324) );
  OAI211_X1 U21442 ( .C1(n18332), .C2(n18324), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18455), .ZN(n18325) );
  OAI211_X1 U21443 ( .C1(n18327), .C2(n18358), .A(n18326), .B(n18325), .ZN(
        P3_U2849) );
  AOI22_X1 U21444 ( .A1(n9731), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18378), 
        .B2(n18328), .ZN(n18335) );
  AOI22_X1 U21445 ( .A1(n18916), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n18329), .B2(n18342), .ZN(n18333) );
  OAI22_X1 U21446 ( .A1(n18330), .A2(n18366), .B1(n18336), .B2(n18461), .ZN(
        n18331) );
  OAI21_X1 U21447 ( .B1(n18333), .B2(n18332), .A(n18331), .ZN(n18334) );
  OAI211_X1 U21448 ( .C1(n18454), .C2(n18336), .A(n18335), .B(n18334), .ZN(
        P3_U2850) );
  AOI22_X1 U21449 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n9731), .B1(n18378), 
        .B2(n18337), .ZN(n18349) );
  AOI22_X1 U21450 ( .A1(n18961), .A2(n18340), .B1(n18339), .B2(n18338), .ZN(
        n18341) );
  OAI211_X1 U21451 ( .C1(n18916), .C2(n18342), .A(n18341), .B(n18454), .ZN(
        n18360) );
  OAI22_X1 U21452 ( .A1(n18916), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n18344), .B2(n18343), .ZN(n18345) );
  NOR2_X1 U21453 ( .A1(n18360), .A2(n18345), .ZN(n18354) );
  OAI211_X1 U21454 ( .C1(n18916), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18346), .B(n18354), .ZN(n18347) );
  NAND3_X1 U21455 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18455), .A3(
        n18347), .ZN(n18348) );
  OAI211_X1 U21456 ( .C1(n18350), .C2(n18366), .A(n18349), .B(n18348), .ZN(
        P3_U2851) );
  AOI21_X1 U21457 ( .B1(n18351), .B2(n18365), .A(n18361), .ZN(n18353) );
  AOI21_X1 U21458 ( .B1(n18354), .B2(n18353), .A(n18352), .ZN(n18356) );
  NOR3_X1 U21459 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18365), .A3(
        n18366), .ZN(n18355) );
  AOI221_X1 U21460 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9731), .C1(n18356), 
        .C2(n18455), .A(n18355), .ZN(n18357) );
  OAI21_X1 U21461 ( .B1(n18359), .B2(n18358), .A(n18357), .ZN(P3_U2852) );
  OAI21_X1 U21462 ( .B1(n18361), .B2(n18360), .A(n18455), .ZN(n18364) );
  AOI22_X1 U21463 ( .A1(n18444), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n18378), 
        .B2(n18362), .ZN(n18363) );
  OAI221_X1 U21464 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18366), .C1(
        n18365), .C2(n18364), .A(n18363), .ZN(P3_U2853) );
  AOI22_X1 U21465 ( .A1(n18963), .A2(n18368), .B1(n18367), .B2(n18426), .ZN(
        n18369) );
  NAND2_X1 U21466 ( .A1(n18369), .A2(n18434), .ZN(n18394) );
  AOI211_X1 U21467 ( .C1(n18370), .C2(n18386), .A(n18385), .B(n18394), .ZN(
        n18371) );
  INV_X1 U21468 ( .A(n18371), .ZN(n18387) );
  AOI21_X1 U21469 ( .B1(n18446), .B2(n18387), .A(n18439), .ZN(n18382) );
  NOR4_X1 U21470 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18385), .A3(
        n18386), .A4(n18384), .ZN(n18372) );
  AOI21_X1 U21471 ( .B1(n18373), .B2(n18961), .A(n18372), .ZN(n18374) );
  OAI21_X1 U21472 ( .B1(n18376), .B2(n18375), .A(n18374), .ZN(n18379) );
  AOI22_X1 U21473 ( .A1(n18438), .A2(n18379), .B1(n18378), .B2(n18377), .ZN(
        n18381) );
  OAI211_X1 U21474 ( .C1(n18382), .C2(n20850), .A(n18381), .B(n18380), .ZN(
        P3_U2854) );
  INV_X1 U21475 ( .A(n18458), .ZN(n18449) );
  AOI21_X1 U21476 ( .B1(n18439), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18383), .ZN(n18391) );
  AOI221_X1 U21477 ( .B1(n18386), .B2(n18385), .C1(n18384), .C2(n18385), .A(
        n18461), .ZN(n18388) );
  AOI22_X1 U21478 ( .A1(n18460), .A2(n18389), .B1(n18388), .B2(n18387), .ZN(
        n18390) );
  OAI211_X1 U21479 ( .C1(n18449), .C2(n18392), .A(n18391), .B(n18390), .ZN(
        P3_U2855) );
  NAND3_X1 U21480 ( .A1(n18438), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18422), .ZN(n18418) );
  NOR2_X1 U21481 ( .A1(n18393), .A2(n18418), .ZN(n18396) );
  OAI21_X1 U21482 ( .B1(n18461), .B2(n18394), .A(n18455), .ZN(n18395) );
  INV_X1 U21483 ( .A(n18395), .ZN(n18402) );
  MUX2_X1 U21484 ( .A(n18396), .B(n18402), .S(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Z(n18397) );
  AOI21_X1 U21485 ( .B1(n18460), .B2(n18398), .A(n18397), .ZN(n18400) );
  OAI211_X1 U21486 ( .C1(n18449), .C2(n18401), .A(n18400), .B(n18399), .ZN(
        P3_U2856) );
  NOR2_X1 U21487 ( .A1(n18417), .A2(n18418), .ZN(n18403) );
  MUX2_X1 U21488 ( .A(n18403), .B(n18402), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18404) );
  AOI21_X1 U21489 ( .B1(n18460), .B2(n18405), .A(n18404), .ZN(n18407) );
  NAND2_X1 U21490 ( .A1(n18444), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18406) );
  OAI211_X1 U21491 ( .C1(n18408), .C2(n18449), .A(n18407), .B(n18406), .ZN(
        P3_U2857) );
  AOI22_X1 U21492 ( .A1(n18963), .A2(n18410), .B1(n18409), .B2(n18426), .ZN(
        n18411) );
  NAND3_X1 U21493 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18411), .A3(
        n18434), .ZN(n18421) );
  AOI21_X1 U21494 ( .B1(n18446), .B2(n18421), .A(n18439), .ZN(n18416) );
  OAI22_X1 U21495 ( .A1(n20983), .A2(n18455), .B1(n18449), .B2(n18412), .ZN(
        n18413) );
  AOI21_X1 U21496 ( .B1(n18460), .B2(n18414), .A(n18413), .ZN(n18415) );
  OAI221_X1 U21497 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18418), .C1(
        n18417), .C2(n18416), .A(n18415), .ZN(P3_U2858) );
  AOI22_X1 U21498 ( .A1(n9731), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18458), .B2(
        n18419), .ZN(n18425) );
  AOI22_X1 U21499 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18439), .B1(
        n18460), .B2(n18420), .ZN(n18424) );
  OAI211_X1 U21500 ( .C1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n18422), .A(
        n18438), .B(n18421), .ZN(n18423) );
  NAND3_X1 U21501 ( .A1(n18425), .A2(n18424), .A3(n18423), .ZN(P3_U2859) );
  NOR2_X1 U21502 ( .A1(n19106), .A2(n19090), .ZN(n18427) );
  AOI22_X1 U21503 ( .A1(n18963), .A2(n18427), .B1(n19090), .B2(n18426), .ZN(
        n18435) );
  NOR2_X1 U21504 ( .A1(n18943), .A2(n18428), .ZN(n18431) );
  NOR3_X1 U21505 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n19090), .A3(
        n18429), .ZN(n18430) );
  AOI211_X1 U21506 ( .C1(n18432), .C2(n18961), .A(n18431), .B(n18430), .ZN(
        n18433) );
  OAI221_X1 U21507 ( .B1(n18436), .B2(n18435), .C1(n18436), .C2(n18434), .A(
        n18433), .ZN(n18437) );
  AOI22_X1 U21508 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18439), .B1(
        n18438), .B2(n18437), .ZN(n18441) );
  OAI211_X1 U21509 ( .C1(n18442), .C2(n18449), .A(n18441), .B(n18440), .ZN(
        P3_U2860) );
  OR3_X1 U21510 ( .A1(n18461), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18443), .ZN(n18463) );
  NAND2_X1 U21511 ( .A1(n18444), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18448) );
  NAND3_X1 U21512 ( .A1(n18446), .A2(n19090), .A3(n18445), .ZN(n18447) );
  OAI211_X1 U21513 ( .C1(n18450), .C2(n18449), .A(n18448), .B(n18447), .ZN(
        n18451) );
  AOI21_X1 U21514 ( .B1(n18460), .B2(n18452), .A(n18451), .ZN(n18453) );
  OAI221_X1 U21515 ( .B1(n19090), .B2(n18454), .C1(n19090), .C2(n18463), .A(
        n18453), .ZN(P3_U2861) );
  NOR2_X1 U21516 ( .A1(n20771), .A2(n18455), .ZN(n18456) );
  AOI221_X1 U21517 ( .B1(n18460), .B2(n18459), .C1(n18458), .C2(n18457), .A(
        n18456), .ZN(n18464) );
  OAI211_X1 U21518 ( .C1(n18947), .C2(n18461), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18455), .ZN(n18462) );
  NAND3_X1 U21519 ( .A1(n18464), .A2(n18463), .A3(n18462), .ZN(P3_U2862) );
  AOI211_X1 U21520 ( .C1(n18466), .C2(n18465), .A(n19143), .B(n19088), .ZN(
        n18978) );
  OAI21_X1 U21521 ( .B1(n18978), .B2(n18520), .A(n18471), .ZN(n18467) );
  OAI221_X1 U21522 ( .B1(n18932), .B2(n19127), .C1(n18932), .C2(n18471), .A(
        n18467), .ZN(P3_U2863) );
  NAND2_X1 U21523 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18653) );
  AOI221_X1 U21524 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18653), .C1(n18469), 
        .C2(n18653), .A(n18468), .ZN(n18476) );
  NOR2_X1 U21525 ( .A1(n18470), .A2(n18934), .ZN(n18472) );
  OAI21_X1 U21526 ( .B1(n18472), .B2(n18482), .A(n18471), .ZN(n18474) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18476), .B1(
        n18474), .B2(n18938), .ZN(P3_U2865) );
  NAND2_X1 U21528 ( .A1(n18479), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18609) );
  NAND2_X1 U21529 ( .A1(n18938), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18745) );
  INV_X1 U21530 ( .A(n18745), .ZN(n18473) );
  NAND2_X1 U21531 ( .A1(n18482), .A2(n18473), .ZN(n18768) );
  AND2_X1 U21532 ( .A1(n18609), .A2(n18768), .ZN(n18475) );
  OAI22_X1 U21533 ( .A1(n18476), .A2(n18479), .B1(n18475), .B2(n18474), .ZN(
        P3_U2866) );
  AND2_X1 U21534 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18477), .ZN(
        P3_U2867) );
  NAND2_X1 U21535 ( .A1(n18862), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18866) );
  NOR2_X1 U21536 ( .A1(n18938), .A2(n18479), .ZN(n18480) );
  NAND2_X1 U21537 ( .A1(n18932), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18721) );
  INV_X1 U21538 ( .A(n18721), .ZN(n18630) );
  NAND2_X1 U21539 ( .A1(n18480), .A2(n18630), .ZN(n18539) );
  NOR2_X2 U21540 ( .A1(n18562), .A2(n18478), .ZN(n18858) );
  INV_X1 U21541 ( .A(n18856), .ZN(n18987) );
  NOR2_X1 U21542 ( .A1(n18479), .A2(n18653), .ZN(n18860) );
  NAND2_X1 U21543 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18860), .ZN(
        n18556) );
  INV_X1 U21544 ( .A(n18556), .ZN(n18910) );
  NOR2_X1 U21545 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18584) );
  NOR2_X1 U21546 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18563) );
  NAND2_X1 U21547 ( .A1(n18584), .A2(n18563), .ZN(n18583) );
  INV_X1 U21548 ( .A(n18583), .ZN(n18574) );
  NOR2_X1 U21549 ( .A1(n18910), .A2(n18574), .ZN(n18540) );
  NOR2_X1 U21550 ( .A1(n18987), .A2(n18540), .ZN(n18514) );
  NAND2_X1 U21551 ( .A1(n18480), .A2(n18934), .ZN(n18798) );
  INV_X1 U21552 ( .A(n18798), .ZN(n18861) );
  NAND2_X1 U21553 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18861), .ZN(
        n18915) );
  INV_X1 U21554 ( .A(n18915), .ZN(n18899) );
  NAND2_X1 U21555 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18862), .ZN(n18832) );
  INV_X1 U21556 ( .A(n18832), .ZN(n18857) );
  AOI22_X1 U21557 ( .A1(n18858), .A2(n18514), .B1(n18899), .B2(n18857), .ZN(
        n18487) );
  NAND2_X1 U21558 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18934), .ZN(
        n18700) );
  NAND2_X1 U21559 ( .A1(n18721), .A2(n18700), .ZN(n18767) );
  NAND2_X1 U21560 ( .A1(n18480), .A2(n18767), .ZN(n18824) );
  NOR2_X1 U21561 ( .A1(n18562), .A2(n18824), .ZN(n18829) );
  INV_X1 U21562 ( .A(n18562), .ZN(n18771) );
  AOI21_X1 U21563 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18540), .ZN(n18481) );
  AOI22_X1 U21564 ( .A1(n18482), .A2(n18829), .B1(n18771), .B2(n18481), .ZN(
        n18517) );
  NAND2_X1 U21565 ( .A1(n18484), .A2(n18483), .ZN(n18515) );
  NOR2_X2 U21566 ( .A1(n18485), .A2(n18515), .ZN(n18863) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18863), .ZN(n18486) );
  OAI211_X1 U21568 ( .C1(n18866), .C2(n18539), .A(n18487), .B(n18486), .ZN(
        P3_U2868) );
  NOR2_X1 U21569 ( .A1(n13868), .A2(n18826), .ZN(n18868) );
  INV_X1 U21570 ( .A(n18868), .ZN(n18777) );
  AND2_X1 U21571 ( .A1(n18771), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18867) );
  NAND2_X1 U21572 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18862), .ZN(n18872) );
  INV_X1 U21573 ( .A(n18872), .ZN(n18774) );
  AOI22_X1 U21574 ( .A1(n18514), .A2(n18867), .B1(n18899), .B2(n18774), .ZN(
        n18489) );
  NOR2_X2 U21575 ( .A1(n19132), .A2(n18515), .ZN(n18869) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18869), .ZN(n18488) );
  OAI211_X1 U21577 ( .C1(n18539), .C2(n18777), .A(n18489), .B(n18488), .ZN(
        P3_U2869) );
  NAND2_X1 U21578 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n18862), .ZN(n18838) );
  NOR2_X2 U21579 ( .A1(n18490), .A2(n18562), .ZN(n18873) );
  NAND2_X1 U21580 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18862), .ZN(n18878) );
  INV_X1 U21581 ( .A(n18878), .ZN(n18835) );
  AOI22_X1 U21582 ( .A1(n18514), .A2(n18873), .B1(n18899), .B2(n18835), .ZN(
        n18493) );
  NOR2_X2 U21583 ( .A1(n18491), .A2(n18515), .ZN(n18875) );
  AOI22_X1 U21584 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18875), .ZN(n18492) );
  OAI211_X1 U21585 ( .C1(n18539), .C2(n18838), .A(n18493), .B(n18492), .ZN(
        P3_U2870) );
  INV_X1 U21586 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18494) );
  NOR2_X1 U21587 ( .A1(n18494), .A2(n18826), .ZN(n18880) );
  INV_X1 U21588 ( .A(n18880), .ZN(n18842) );
  INV_X1 U21589 ( .A(n18539), .ZN(n18852) );
  NAND2_X1 U21590 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n18862), .ZN(n18884) );
  INV_X1 U21591 ( .A(n18884), .ZN(n18839) );
  NOR2_X2 U21592 ( .A1(n18495), .A2(n18562), .ZN(n18879) );
  AOI22_X1 U21593 ( .A1(n18852), .A2(n18839), .B1(n18514), .B2(n18879), .ZN(
        n18498) );
  NOR2_X2 U21594 ( .A1(n18496), .A2(n18515), .ZN(n18881) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18881), .ZN(n18497) );
  OAI211_X1 U21596 ( .C1(n18915), .C2(n18842), .A(n18498), .B(n18497), .ZN(
        P3_U2871) );
  NOR2_X1 U21597 ( .A1(n18499), .A2(n18826), .ZN(n18886) );
  INV_X1 U21598 ( .A(n18886), .ZN(n18811) );
  NAND2_X1 U21599 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18862), .ZN(n18890) );
  INV_X1 U21600 ( .A(n18890), .ZN(n18808) );
  NOR2_X2 U21601 ( .A1(n18500), .A2(n18562), .ZN(n18885) );
  AOI22_X1 U21602 ( .A1(n18852), .A2(n18808), .B1(n18514), .B2(n18885), .ZN(
        n18503) );
  NOR2_X2 U21603 ( .A1(n18501), .A2(n18515), .ZN(n18887) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18887), .ZN(n18502) );
  OAI211_X1 U21605 ( .C1(n18915), .C2(n18811), .A(n18503), .B(n18502), .ZN(
        P3_U2872) );
  INV_X1 U21606 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18504) );
  NOR2_X1 U21607 ( .A1(n18504), .A2(n18826), .ZN(n18784) );
  INV_X1 U21608 ( .A(n18784), .ZN(n18896) );
  NAND2_X1 U21609 ( .A1(BUF2_REG_21__SCAN_IN), .A2(n18862), .ZN(n18787) );
  INV_X1 U21610 ( .A(n18787), .ZN(n18892) );
  NOR2_X2 U21611 ( .A1(n18505), .A2(n18562), .ZN(n18891) );
  AOI22_X1 U21612 ( .A1(n18852), .A2(n18892), .B1(n18514), .B2(n18891), .ZN(
        n18508) );
  NOR2_X2 U21613 ( .A1(n18506), .A2(n18515), .ZN(n18893) );
  AOI22_X1 U21614 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18893), .ZN(n18507) );
  OAI211_X1 U21615 ( .C1(n18915), .C2(n18896), .A(n18508), .B(n18507), .ZN(
        P3_U2873) );
  NAND2_X1 U21616 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n18862), .ZN(n18818) );
  NOR2_X2 U21617 ( .A1(n18509), .A2(n18562), .ZN(n18897) );
  NAND2_X1 U21618 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18862), .ZN(n18904) );
  INV_X1 U21619 ( .A(n18904), .ZN(n18815) );
  AOI22_X1 U21620 ( .A1(n18514), .A2(n18897), .B1(n18899), .B2(n18815), .ZN(
        n18512) );
  NOR2_X2 U21621 ( .A1(n18510), .A2(n18515), .ZN(n18900) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18900), .ZN(n18511) );
  OAI211_X1 U21623 ( .C1(n18539), .C2(n18818), .A(n18512), .B(n18511), .ZN(
        P3_U2874) );
  NAND2_X1 U21624 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18862), .ZN(n18914) );
  NOR2_X2 U21625 ( .A1(n18513), .A2(n18562), .ZN(n18906) );
  NAND2_X1 U21626 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n18862), .ZN(n18797) );
  INV_X1 U21627 ( .A(n18797), .ZN(n18908) );
  AOI22_X1 U21628 ( .A1(n18514), .A2(n18906), .B1(n18899), .B2(n18908), .ZN(
        n18519) );
  NOR2_X2 U21629 ( .A1(n18516), .A2(n18515), .ZN(n18909) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18517), .B1(
        n18574), .B2(n18909), .ZN(n18518) );
  OAI211_X1 U21631 ( .C1(n18539), .C2(n18914), .A(n18519), .B(n18518), .ZN(
        P3_U2875) );
  INV_X1 U21632 ( .A(n18866), .ZN(n18825) );
  INV_X1 U21633 ( .A(n18563), .ZN(n18561) );
  NAND2_X1 U21634 ( .A1(n18934), .A2(n18856), .ZN(n18698) );
  NOR2_X1 U21635 ( .A1(n18561), .A2(n18698), .ZN(n18535) );
  AOI22_X1 U21636 ( .A1(n18825), .A2(n18910), .B1(n18858), .B2(n18535), .ZN(
        n18522) );
  NOR2_X1 U21637 ( .A1(n18562), .A2(n18520), .ZN(n18859) );
  AND2_X1 U21638 ( .A1(n18934), .A2(n18859), .ZN(n18607) );
  AOI22_X1 U21639 ( .A1(n18862), .A2(n18860), .B1(n18563), .B2(n18607), .ZN(
        n18536) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18536), .B1(
        n18863), .B2(n9721), .ZN(n18521) );
  OAI211_X1 U21641 ( .C1(n18539), .C2(n18832), .A(n18522), .B(n18521), .ZN(
        P3_U2876) );
  AOI22_X1 U21642 ( .A1(n18852), .A2(n18774), .B1(n18867), .B2(n18535), .ZN(
        n18524) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18536), .B1(
        n18869), .B2(n9721), .ZN(n18523) );
  OAI211_X1 U21644 ( .C1(n18556), .C2(n18777), .A(n18524), .B(n18523), .ZN(
        P3_U2877) );
  INV_X1 U21645 ( .A(n18838), .ZN(n18874) );
  AOI22_X1 U21646 ( .A1(n18910), .A2(n18874), .B1(n18873), .B2(n18535), .ZN(
        n18526) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18536), .B1(
        n18875), .B2(n9721), .ZN(n18525) );
  OAI211_X1 U21648 ( .C1(n18539), .C2(n18878), .A(n18526), .B(n18525), .ZN(
        P3_U2878) );
  AOI22_X1 U21649 ( .A1(n18852), .A2(n18880), .B1(n18879), .B2(n18535), .ZN(
        n18528) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18536), .B1(
        n18881), .B2(n9721), .ZN(n18527) );
  OAI211_X1 U21651 ( .C1(n18556), .C2(n18884), .A(n18528), .B(n18527), .ZN(
        P3_U2879) );
  AOI22_X1 U21652 ( .A1(n18852), .A2(n18886), .B1(n18885), .B2(n18535), .ZN(
        n18530) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18536), .B1(
        n18887), .B2(n9721), .ZN(n18529) );
  OAI211_X1 U21654 ( .C1(n18556), .C2(n18890), .A(n18530), .B(n18529), .ZN(
        P3_U2880) );
  AOI22_X1 U21655 ( .A1(n18852), .A2(n18784), .B1(n18891), .B2(n18535), .ZN(
        n18532) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18536), .B1(
        n18893), .B2(n9721), .ZN(n18531) );
  OAI211_X1 U21657 ( .C1(n18556), .C2(n18787), .A(n18532), .B(n18531), .ZN(
        P3_U2881) );
  AOI22_X1 U21658 ( .A1(n18852), .A2(n18815), .B1(n18897), .B2(n18535), .ZN(
        n18534) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18536), .B1(
        n18900), .B2(n9721), .ZN(n18533) );
  OAI211_X1 U21660 ( .C1(n18556), .C2(n18818), .A(n18534), .B(n18533), .ZN(
        P3_U2882) );
  INV_X1 U21661 ( .A(n18914), .ZN(n18792) );
  AOI22_X1 U21662 ( .A1(n18910), .A2(n18792), .B1(n18906), .B2(n18535), .ZN(
        n18538) );
  AOI22_X1 U21663 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18536), .B1(
        n18909), .B2(n9721), .ZN(n18537) );
  OAI211_X1 U21664 ( .C1(n18539), .C2(n18797), .A(n18538), .B(n18537), .ZN(
        P3_U2883) );
  NAND2_X1 U21665 ( .A1(n18630), .A2(n18563), .ZN(n18629) );
  INV_X1 U21666 ( .A(n18629), .ZN(n18622) );
  NOR2_X1 U21667 ( .A1(n9721), .A2(n18622), .ZN(n18585) );
  NOR2_X1 U21668 ( .A1(n18987), .A2(n18585), .ZN(n18557) );
  AOI22_X1 U21669 ( .A1(n18910), .A2(n18857), .B1(n18858), .B2(n18557), .ZN(
        n18543) );
  OAI22_X1 U21670 ( .A1(n18540), .A2(n18826), .B1(n18585), .B2(n18562), .ZN(
        n18541) );
  OAI21_X1 U21671 ( .B1(n18622), .B2(n19079), .A(n18541), .ZN(n18558) );
  AOI22_X1 U21672 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18558), .B1(
        n18863), .B2(n18622), .ZN(n18542) );
  OAI211_X1 U21673 ( .C1(n18866), .C2(n18583), .A(n18543), .B(n18542), .ZN(
        P3_U2884) );
  AOI22_X1 U21674 ( .A1(n18574), .A2(n18868), .B1(n18867), .B2(n18557), .ZN(
        n18545) );
  AOI22_X1 U21675 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18558), .B1(
        n18869), .B2(n18622), .ZN(n18544) );
  OAI211_X1 U21676 ( .C1(n18556), .C2(n18872), .A(n18545), .B(n18544), .ZN(
        P3_U2885) );
  AOI22_X1 U21677 ( .A1(n18574), .A2(n18874), .B1(n18873), .B2(n18557), .ZN(
        n18547) );
  AOI22_X1 U21678 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18558), .B1(
        n18875), .B2(n18622), .ZN(n18546) );
  OAI211_X1 U21679 ( .C1(n18556), .C2(n18878), .A(n18547), .B(n18546), .ZN(
        P3_U2886) );
  AOI22_X1 U21680 ( .A1(n18574), .A2(n18839), .B1(n18879), .B2(n18557), .ZN(
        n18549) );
  AOI22_X1 U21681 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18558), .B1(
        n18881), .B2(n18622), .ZN(n18548) );
  OAI211_X1 U21682 ( .C1(n18556), .C2(n18842), .A(n18549), .B(n18548), .ZN(
        P3_U2887) );
  AOI22_X1 U21683 ( .A1(n18574), .A2(n18808), .B1(n18885), .B2(n18557), .ZN(
        n18551) );
  AOI22_X1 U21684 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18558), .B1(
        n18887), .B2(n18622), .ZN(n18550) );
  OAI211_X1 U21685 ( .C1(n18556), .C2(n18811), .A(n18551), .B(n18550), .ZN(
        P3_U2888) );
  AOI22_X1 U21686 ( .A1(n18574), .A2(n18892), .B1(n18891), .B2(n18557), .ZN(
        n18553) );
  AOI22_X1 U21687 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18558), .B1(
        n18893), .B2(n18622), .ZN(n18552) );
  OAI211_X1 U21688 ( .C1(n18556), .C2(n18896), .A(n18553), .B(n18552), .ZN(
        P3_U2889) );
  INV_X1 U21689 ( .A(n18818), .ZN(n18898) );
  AOI22_X1 U21690 ( .A1(n18574), .A2(n18898), .B1(n18897), .B2(n18557), .ZN(
        n18555) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18558), .B1(
        n18900), .B2(n18622), .ZN(n18554) );
  OAI211_X1 U21692 ( .C1(n18556), .C2(n18904), .A(n18555), .B(n18554), .ZN(
        P3_U2890) );
  AOI22_X1 U21693 ( .A1(n18910), .A2(n18908), .B1(n18906), .B2(n18557), .ZN(
        n18560) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18558), .B1(
        n18909), .B2(n18622), .ZN(n18559) );
  OAI211_X1 U21695 ( .C1(n18583), .C2(n18914), .A(n18560), .B(n18559), .ZN(
        P3_U2891) );
  NOR2_X1 U21696 ( .A1(n18934), .A2(n18561), .ZN(n18608) );
  NAND2_X1 U21697 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18608), .ZN(
        n18652) );
  INV_X1 U21698 ( .A(n18652), .ZN(n18645) );
  AOI21_X1 U21699 ( .B1(n18934), .B2(n18722), .A(n18562), .ZN(n18655) );
  OAI211_X1 U21700 ( .C1(n18645), .C2(n19079), .A(n18563), .B(n18655), .ZN(
        n18580) );
  AND2_X1 U21701 ( .A1(n18856), .A2(n18608), .ZN(n18579) );
  AOI22_X1 U21702 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18580), .B1(
        n18858), .B2(n18579), .ZN(n18565) );
  AOI22_X1 U21703 ( .A1(n18825), .A2(n9721), .B1(n18863), .B2(n18645), .ZN(
        n18564) );
  OAI211_X1 U21704 ( .C1(n18583), .C2(n18832), .A(n18565), .B(n18564), .ZN(
        P3_U2892) );
  AOI22_X1 U21705 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18580), .B1(
        n18867), .B2(n18579), .ZN(n18567) );
  AOI22_X1 U21706 ( .A1(n18868), .A2(n9721), .B1(n18869), .B2(n18645), .ZN(
        n18566) );
  OAI211_X1 U21707 ( .C1(n18583), .C2(n18872), .A(n18567), .B(n18566), .ZN(
        P3_U2893) );
  INV_X1 U21708 ( .A(n9721), .ZN(n18589) );
  AOI22_X1 U21709 ( .A1(n18574), .A2(n18835), .B1(n18873), .B2(n18579), .ZN(
        n18569) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18580), .B1(
        n18875), .B2(n18645), .ZN(n18568) );
  OAI211_X1 U21711 ( .C1(n18838), .C2(n18589), .A(n18569), .B(n18568), .ZN(
        P3_U2894) );
  AOI22_X1 U21712 ( .A1(n18839), .A2(n9721), .B1(n18879), .B2(n18579), .ZN(
        n18571) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18580), .B1(
        n18881), .B2(n18645), .ZN(n18570) );
  OAI211_X1 U21714 ( .C1(n18583), .C2(n18842), .A(n18571), .B(n18570), .ZN(
        P3_U2895) );
  AOI22_X1 U21715 ( .A1(n18574), .A2(n18886), .B1(n18885), .B2(n18579), .ZN(
        n18573) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18580), .B1(
        n18887), .B2(n18645), .ZN(n18572) );
  OAI211_X1 U21717 ( .C1(n18890), .C2(n18589), .A(n18573), .B(n18572), .ZN(
        P3_U2896) );
  AOI22_X1 U21718 ( .A1(n18574), .A2(n18784), .B1(n18891), .B2(n18579), .ZN(
        n18576) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18580), .B1(
        n18893), .B2(n18645), .ZN(n18575) );
  OAI211_X1 U21720 ( .C1(n18787), .C2(n18589), .A(n18576), .B(n18575), .ZN(
        P3_U2897) );
  AOI22_X1 U21721 ( .A1(n18898), .A2(n9721), .B1(n18897), .B2(n18579), .ZN(
        n18578) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18580), .B1(
        n18900), .B2(n18645), .ZN(n18577) );
  OAI211_X1 U21723 ( .C1(n18583), .C2(n18904), .A(n18578), .B(n18577), .ZN(
        P3_U2898) );
  AOI22_X1 U21724 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18580), .B1(
        n18906), .B2(n18579), .ZN(n18582) );
  AOI22_X1 U21725 ( .A1(n18792), .A2(n9721), .B1(n18909), .B2(n18645), .ZN(
        n18581) );
  OAI211_X1 U21726 ( .C1(n18583), .C2(n18797), .A(n18582), .B(n18581), .ZN(
        P3_U2899) );
  INV_X1 U21727 ( .A(n18584), .ZN(n18935) );
  NOR2_X2 U21728 ( .A1(n18935), .A2(n18609), .ZN(n18673) );
  INV_X1 U21729 ( .A(n18673), .ZN(n18666) );
  AOI21_X1 U21730 ( .B1(n18652), .B2(n18666), .A(n18987), .ZN(n18602) );
  AOI22_X1 U21731 ( .A1(n18825), .A2(n18622), .B1(n18858), .B2(n18602), .ZN(
        n18588) );
  AOI221_X1 U21732 ( .B1(n18585), .B2(n18652), .C1(n18722), .C2(n18652), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18586) );
  OAI21_X1 U21733 ( .B1(n18673), .B2(n18586), .A(n18771), .ZN(n18604) );
  AOI22_X1 U21734 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18604), .B1(
        n18863), .B2(n18673), .ZN(n18587) );
  OAI211_X1 U21735 ( .C1(n18832), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        P3_U2900) );
  AOI22_X1 U21736 ( .A1(n18774), .A2(n9721), .B1(n18867), .B2(n18602), .ZN(
        n18591) );
  AOI22_X1 U21737 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18604), .B1(
        n18869), .B2(n18673), .ZN(n18590) );
  OAI211_X1 U21738 ( .C1(n18777), .C2(n18629), .A(n18591), .B(n18590), .ZN(
        P3_U2901) );
  AOI22_X1 U21739 ( .A1(n18835), .A2(n9721), .B1(n18873), .B2(n18602), .ZN(
        n18593) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18604), .B1(
        n18875), .B2(n18673), .ZN(n18592) );
  OAI211_X1 U21741 ( .C1(n18838), .C2(n18629), .A(n18593), .B(n18592), .ZN(
        P3_U2902) );
  AOI22_X1 U21742 ( .A1(n18880), .A2(n9721), .B1(n18879), .B2(n18602), .ZN(
        n18595) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18604), .B1(
        n18881), .B2(n18673), .ZN(n18594) );
  OAI211_X1 U21744 ( .C1(n18884), .C2(n18629), .A(n18595), .B(n18594), .ZN(
        P3_U2903) );
  AOI22_X1 U21745 ( .A1(n18886), .A2(n9721), .B1(n18885), .B2(n18602), .ZN(
        n18597) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18604), .B1(
        n18887), .B2(n18673), .ZN(n18596) );
  OAI211_X1 U21747 ( .C1(n18890), .C2(n18629), .A(n18597), .B(n18596), .ZN(
        P3_U2904) );
  AOI22_X1 U21748 ( .A1(n18784), .A2(n9721), .B1(n18891), .B2(n18602), .ZN(
        n18599) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18604), .B1(
        n18893), .B2(n18673), .ZN(n18598) );
  OAI211_X1 U21750 ( .C1(n18787), .C2(n18629), .A(n18599), .B(n18598), .ZN(
        P3_U2905) );
  AOI22_X1 U21751 ( .A1(n18815), .A2(n9721), .B1(n18897), .B2(n18602), .ZN(
        n18601) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18604), .B1(
        n18900), .B2(n18673), .ZN(n18600) );
  OAI211_X1 U21753 ( .C1(n18818), .C2(n18629), .A(n18601), .B(n18600), .ZN(
        P3_U2906) );
  AOI22_X1 U21754 ( .A1(n18908), .A2(n9721), .B1(n18906), .B2(n18602), .ZN(
        n18606) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18604), .B1(
        n18909), .B2(n18673), .ZN(n18605) );
  OAI211_X1 U21756 ( .C1(n18914), .C2(n18629), .A(n18606), .B(n18605), .ZN(
        P3_U2907) );
  NOR2_X1 U21757 ( .A1(n18698), .A2(n18609), .ZN(n18625) );
  AOI22_X1 U21758 ( .A1(n18858), .A2(n18625), .B1(n18857), .B2(n18622), .ZN(
        n18611) );
  INV_X1 U21759 ( .A(n18609), .ZN(n18654) );
  AOI22_X1 U21760 ( .A1(n18862), .A2(n18608), .B1(n18607), .B2(n18654), .ZN(
        n18626) );
  NOR2_X2 U21761 ( .A1(n18700), .A2(n18609), .ZN(n18694) );
  AOI22_X1 U21762 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18626), .B1(
        n18863), .B2(n18694), .ZN(n18610) );
  OAI211_X1 U21763 ( .C1(n18866), .C2(n18652), .A(n18611), .B(n18610), .ZN(
        P3_U2908) );
  AOI22_X1 U21764 ( .A1(n18774), .A2(n18622), .B1(n18867), .B2(n18625), .ZN(
        n18613) );
  AOI22_X1 U21765 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18626), .B1(
        n18869), .B2(n18694), .ZN(n18612) );
  OAI211_X1 U21766 ( .C1(n18777), .C2(n18652), .A(n18613), .B(n18612), .ZN(
        P3_U2909) );
  AOI22_X1 U21767 ( .A1(n18835), .A2(n18622), .B1(n18873), .B2(n18625), .ZN(
        n18615) );
  AOI22_X1 U21768 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18626), .B1(
        n18875), .B2(n18694), .ZN(n18614) );
  OAI211_X1 U21769 ( .C1(n18838), .C2(n18652), .A(n18615), .B(n18614), .ZN(
        P3_U2910) );
  AOI22_X1 U21770 ( .A1(n18839), .A2(n18645), .B1(n18879), .B2(n18625), .ZN(
        n18617) );
  AOI22_X1 U21771 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18626), .B1(
        n18881), .B2(n18694), .ZN(n18616) );
  OAI211_X1 U21772 ( .C1(n18842), .C2(n18629), .A(n18617), .B(n18616), .ZN(
        P3_U2911) );
  AOI22_X1 U21773 ( .A1(n18808), .A2(n18645), .B1(n18885), .B2(n18625), .ZN(
        n18619) );
  AOI22_X1 U21774 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18626), .B1(
        n18887), .B2(n18694), .ZN(n18618) );
  OAI211_X1 U21775 ( .C1(n18811), .C2(n18629), .A(n18619), .B(n18618), .ZN(
        P3_U2912) );
  AOI22_X1 U21776 ( .A1(n18892), .A2(n18645), .B1(n18891), .B2(n18625), .ZN(
        n18621) );
  AOI22_X1 U21777 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18626), .B1(
        n18893), .B2(n18694), .ZN(n18620) );
  OAI211_X1 U21778 ( .C1(n18896), .C2(n18629), .A(n18621), .B(n18620), .ZN(
        P3_U2913) );
  AOI22_X1 U21779 ( .A1(n18815), .A2(n18622), .B1(n18897), .B2(n18625), .ZN(
        n18624) );
  AOI22_X1 U21780 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18626), .B1(
        n18900), .B2(n18694), .ZN(n18623) );
  OAI211_X1 U21781 ( .C1(n18818), .C2(n18652), .A(n18624), .B(n18623), .ZN(
        P3_U2914) );
  AOI22_X1 U21782 ( .A1(n18792), .A2(n18645), .B1(n18906), .B2(n18625), .ZN(
        n18628) );
  AOI22_X1 U21783 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18626), .B1(
        n18909), .B2(n18694), .ZN(n18627) );
  OAI211_X1 U21784 ( .C1(n18797), .C2(n18629), .A(n18628), .B(n18627), .ZN(
        P3_U2915) );
  NAND2_X1 U21785 ( .A1(n18630), .A2(n18654), .ZN(n18720) );
  INV_X1 U21786 ( .A(n18720), .ZN(n18709) );
  NOR2_X1 U21787 ( .A1(n18694), .A2(n18709), .ZN(n18676) );
  NOR2_X1 U21788 ( .A1(n18987), .A2(n18676), .ZN(n18648) );
  AOI22_X1 U21789 ( .A1(n18825), .A2(n18673), .B1(n18858), .B2(n18648), .ZN(
        n18634) );
  NOR2_X1 U21790 ( .A1(n18645), .A2(n18673), .ZN(n18631) );
  OAI21_X1 U21791 ( .B1(n18631), .B2(n18722), .A(n18676), .ZN(n18632) );
  OAI211_X1 U21792 ( .C1(n18709), .C2(n19079), .A(n18771), .B(n18632), .ZN(
        n18649) );
  AOI22_X1 U21793 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18649), .B1(
        n18863), .B2(n18709), .ZN(n18633) );
  OAI211_X1 U21794 ( .C1(n18832), .C2(n18652), .A(n18634), .B(n18633), .ZN(
        P3_U2916) );
  AOI22_X1 U21795 ( .A1(n18774), .A2(n18645), .B1(n18867), .B2(n18648), .ZN(
        n18636) );
  AOI22_X1 U21796 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18649), .B1(
        n18869), .B2(n18709), .ZN(n18635) );
  OAI211_X1 U21797 ( .C1(n18777), .C2(n18666), .A(n18636), .B(n18635), .ZN(
        P3_U2917) );
  AOI22_X1 U21798 ( .A1(n18835), .A2(n18645), .B1(n18873), .B2(n18648), .ZN(
        n18638) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18649), .B1(
        n18875), .B2(n18709), .ZN(n18637) );
  OAI211_X1 U21800 ( .C1(n18838), .C2(n18666), .A(n18638), .B(n18637), .ZN(
        P3_U2918) );
  AOI22_X1 U21801 ( .A1(n18880), .A2(n18645), .B1(n18879), .B2(n18648), .ZN(
        n18640) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18649), .B1(
        n18881), .B2(n18709), .ZN(n18639) );
  OAI211_X1 U21803 ( .C1(n18884), .C2(n18666), .A(n18640), .B(n18639), .ZN(
        P3_U2919) );
  AOI22_X1 U21804 ( .A1(n18808), .A2(n18673), .B1(n18885), .B2(n18648), .ZN(
        n18642) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18649), .B1(
        n18887), .B2(n18709), .ZN(n18641) );
  OAI211_X1 U21806 ( .C1(n18811), .C2(n18652), .A(n18642), .B(n18641), .ZN(
        P3_U2920) );
  AOI22_X1 U21807 ( .A1(n18784), .A2(n18645), .B1(n18891), .B2(n18648), .ZN(
        n18644) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18649), .B1(
        n18893), .B2(n18709), .ZN(n18643) );
  OAI211_X1 U21809 ( .C1(n18787), .C2(n18666), .A(n18644), .B(n18643), .ZN(
        P3_U2921) );
  AOI22_X1 U21810 ( .A1(n18815), .A2(n18645), .B1(n18897), .B2(n18648), .ZN(
        n18647) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18649), .B1(
        n18900), .B2(n18709), .ZN(n18646) );
  OAI211_X1 U21812 ( .C1(n18818), .C2(n18666), .A(n18647), .B(n18646), .ZN(
        P3_U2922) );
  AOI22_X1 U21813 ( .A1(n18792), .A2(n18673), .B1(n18906), .B2(n18648), .ZN(
        n18651) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18649), .B1(
        n18909), .B2(n18709), .ZN(n18650) );
  OAI211_X1 U21815 ( .C1(n18797), .C2(n18652), .A(n18651), .B(n18650), .ZN(
        P3_U2923) );
  NOR2_X1 U21816 ( .A1(n18653), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18699) );
  AND2_X1 U21817 ( .A1(n18856), .A2(n18699), .ZN(n18671) );
  AOI22_X1 U21818 ( .A1(n18825), .A2(n18694), .B1(n18858), .B2(n18671), .ZN(
        n18657) );
  NAND2_X1 U21819 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18699), .ZN(
        n18737) );
  INV_X1 U21820 ( .A(n18737), .ZN(n18741) );
  OAI211_X1 U21821 ( .C1(n18741), .C2(n19079), .A(n18655), .B(n18654), .ZN(
        n18672) );
  AOI22_X1 U21822 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18672), .B1(
        n18863), .B2(n18741), .ZN(n18656) );
  OAI211_X1 U21823 ( .C1(n18832), .C2(n18666), .A(n18657), .B(n18656), .ZN(
        P3_U2924) );
  AOI22_X1 U21824 ( .A1(n18868), .A2(n18694), .B1(n18867), .B2(n18671), .ZN(
        n18659) );
  AOI22_X1 U21825 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18672), .B1(
        n18869), .B2(n18741), .ZN(n18658) );
  OAI211_X1 U21826 ( .C1(n18872), .C2(n18666), .A(n18659), .B(n18658), .ZN(
        P3_U2925) );
  AOI22_X1 U21827 ( .A1(n18874), .A2(n18694), .B1(n18873), .B2(n18671), .ZN(
        n18661) );
  AOI22_X1 U21828 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18672), .B1(
        n18875), .B2(n18741), .ZN(n18660) );
  OAI211_X1 U21829 ( .C1(n18878), .C2(n18666), .A(n18661), .B(n18660), .ZN(
        P3_U2926) );
  AOI22_X1 U21830 ( .A1(n18839), .A2(n18694), .B1(n18879), .B2(n18671), .ZN(
        n18663) );
  AOI22_X1 U21831 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18672), .B1(
        n18881), .B2(n18741), .ZN(n18662) );
  OAI211_X1 U21832 ( .C1(n18842), .C2(n18666), .A(n18663), .B(n18662), .ZN(
        P3_U2927) );
  AOI22_X1 U21833 ( .A1(n18808), .A2(n18694), .B1(n18885), .B2(n18671), .ZN(
        n18665) );
  AOI22_X1 U21834 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18672), .B1(
        n18887), .B2(n18741), .ZN(n18664) );
  OAI211_X1 U21835 ( .C1(n18811), .C2(n18666), .A(n18665), .B(n18664), .ZN(
        P3_U2928) );
  INV_X1 U21836 ( .A(n18694), .ZN(n18690) );
  AOI22_X1 U21837 ( .A1(n18784), .A2(n18673), .B1(n18891), .B2(n18671), .ZN(
        n18668) );
  AOI22_X1 U21838 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18672), .B1(
        n18893), .B2(n18741), .ZN(n18667) );
  OAI211_X1 U21839 ( .C1(n18787), .C2(n18690), .A(n18668), .B(n18667), .ZN(
        P3_U2929) );
  AOI22_X1 U21840 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18672), .B1(
        n18897), .B2(n18671), .ZN(n18670) );
  AOI22_X1 U21841 ( .A1(n18900), .A2(n18741), .B1(n18815), .B2(n18673), .ZN(
        n18669) );
  OAI211_X1 U21842 ( .C1(n18818), .C2(n18690), .A(n18670), .B(n18669), .ZN(
        P3_U2930) );
  AOI22_X1 U21843 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18672), .B1(
        n18906), .B2(n18671), .ZN(n18675) );
  AOI22_X1 U21844 ( .A1(n18909), .A2(n18741), .B1(n18908), .B2(n18673), .ZN(
        n18674) );
  OAI211_X1 U21845 ( .C1(n18914), .C2(n18690), .A(n18675), .B(n18674), .ZN(
        P3_U2931) );
  NOR2_X2 U21846 ( .A1(n18935), .A2(n18745), .ZN(n18755) );
  INV_X1 U21847 ( .A(n18755), .ZN(n18766) );
  AOI21_X1 U21848 ( .B1(n18737), .B2(n18766), .A(n18987), .ZN(n18693) );
  AOI22_X1 U21849 ( .A1(n18858), .A2(n18693), .B1(n18857), .B2(n18694), .ZN(
        n18679) );
  AOI221_X1 U21850 ( .B1(n18676), .B2(n18737), .C1(n18722), .C2(n18737), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18677) );
  OAI21_X1 U21851 ( .B1(n18755), .B2(n18677), .A(n18771), .ZN(n18695) );
  AOI22_X1 U21852 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18695), .B1(
        n18863), .B2(n18755), .ZN(n18678) );
  OAI211_X1 U21853 ( .C1(n18866), .C2(n18720), .A(n18679), .B(n18678), .ZN(
        P3_U2932) );
  AOI22_X1 U21854 ( .A1(n18774), .A2(n18694), .B1(n18867), .B2(n18693), .ZN(
        n18681) );
  AOI22_X1 U21855 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18695), .B1(
        n18869), .B2(n18755), .ZN(n18680) );
  OAI211_X1 U21856 ( .C1(n18777), .C2(n18720), .A(n18681), .B(n18680), .ZN(
        P3_U2933) );
  AOI22_X1 U21857 ( .A1(n18874), .A2(n18709), .B1(n18873), .B2(n18693), .ZN(
        n18683) );
  AOI22_X1 U21858 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18695), .B1(
        n18875), .B2(n18755), .ZN(n18682) );
  OAI211_X1 U21859 ( .C1(n18878), .C2(n18690), .A(n18683), .B(n18682), .ZN(
        P3_U2934) );
  AOI22_X1 U21860 ( .A1(n18839), .A2(n18709), .B1(n18879), .B2(n18693), .ZN(
        n18685) );
  AOI22_X1 U21861 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18695), .B1(
        n18881), .B2(n18755), .ZN(n18684) );
  OAI211_X1 U21862 ( .C1(n18842), .C2(n18690), .A(n18685), .B(n18684), .ZN(
        P3_U2935) );
  AOI22_X1 U21863 ( .A1(n18808), .A2(n18709), .B1(n18885), .B2(n18693), .ZN(
        n18687) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18695), .B1(
        n18887), .B2(n18755), .ZN(n18686) );
  OAI211_X1 U21865 ( .C1(n18811), .C2(n18690), .A(n18687), .B(n18686), .ZN(
        P3_U2936) );
  AOI22_X1 U21866 ( .A1(n18892), .A2(n18709), .B1(n18891), .B2(n18693), .ZN(
        n18689) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18695), .B1(
        n18893), .B2(n18755), .ZN(n18688) );
  OAI211_X1 U21868 ( .C1(n18896), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        P3_U2937) );
  AOI22_X1 U21869 ( .A1(n18815), .A2(n18694), .B1(n18897), .B2(n18693), .ZN(
        n18692) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18695), .B1(
        n18900), .B2(n18755), .ZN(n18691) );
  OAI211_X1 U21871 ( .C1(n18818), .C2(n18720), .A(n18692), .B(n18691), .ZN(
        P3_U2938) );
  AOI22_X1 U21872 ( .A1(n18908), .A2(n18694), .B1(n18906), .B2(n18693), .ZN(
        n18697) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18695), .B1(
        n18909), .B2(n18755), .ZN(n18696) );
  OAI211_X1 U21874 ( .C1(n18914), .C2(n18720), .A(n18697), .B(n18696), .ZN(
        P3_U2939) );
  NOR2_X1 U21875 ( .A1(n18698), .A2(n18745), .ZN(n18716) );
  AOI22_X1 U21876 ( .A1(n18858), .A2(n18716), .B1(n18857), .B2(n18709), .ZN(
        n18702) );
  NOR2_X1 U21877 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18745), .ZN(
        n18746) );
  AOI22_X1 U21878 ( .A1(n18862), .A2(n18699), .B1(n18859), .B2(n18746), .ZN(
        n18717) );
  NOR2_X2 U21879 ( .A1(n18700), .A2(n18745), .ZN(n18788) );
  AOI22_X1 U21880 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18717), .B1(
        n18863), .B2(n18788), .ZN(n18701) );
  OAI211_X1 U21881 ( .C1(n18866), .C2(n18737), .A(n18702), .B(n18701), .ZN(
        P3_U2940) );
  AOI22_X1 U21882 ( .A1(n18774), .A2(n18709), .B1(n18867), .B2(n18716), .ZN(
        n18704) );
  AOI22_X1 U21883 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18717), .B1(
        n18869), .B2(n18788), .ZN(n18703) );
  OAI211_X1 U21884 ( .C1(n18777), .C2(n18737), .A(n18704), .B(n18703), .ZN(
        P3_U2941) );
  AOI22_X1 U21885 ( .A1(n18835), .A2(n18709), .B1(n18873), .B2(n18716), .ZN(
        n18706) );
  AOI22_X1 U21886 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18717), .B1(
        n18875), .B2(n18788), .ZN(n18705) );
  OAI211_X1 U21887 ( .C1(n18838), .C2(n18737), .A(n18706), .B(n18705), .ZN(
        P3_U2942) );
  AOI22_X1 U21888 ( .A1(n18839), .A2(n18741), .B1(n18879), .B2(n18716), .ZN(
        n18708) );
  AOI22_X1 U21889 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18717), .B1(
        n18881), .B2(n18788), .ZN(n18707) );
  OAI211_X1 U21890 ( .C1(n18842), .C2(n18720), .A(n18708), .B(n18707), .ZN(
        P3_U2943) );
  AOI22_X1 U21891 ( .A1(n18886), .A2(n18709), .B1(n18885), .B2(n18716), .ZN(
        n18711) );
  AOI22_X1 U21892 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18717), .B1(
        n18887), .B2(n18788), .ZN(n18710) );
  OAI211_X1 U21893 ( .C1(n18890), .C2(n18737), .A(n18711), .B(n18710), .ZN(
        P3_U2944) );
  AOI22_X1 U21894 ( .A1(n18892), .A2(n18741), .B1(n18891), .B2(n18716), .ZN(
        n18713) );
  AOI22_X1 U21895 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18717), .B1(
        n18893), .B2(n18788), .ZN(n18712) );
  OAI211_X1 U21896 ( .C1(n18896), .C2(n18720), .A(n18713), .B(n18712), .ZN(
        P3_U2945) );
  AOI22_X1 U21897 ( .A1(n18898), .A2(n18741), .B1(n18897), .B2(n18716), .ZN(
        n18715) );
  AOI22_X1 U21898 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18717), .B1(
        n18900), .B2(n18788), .ZN(n18714) );
  OAI211_X1 U21899 ( .C1(n18904), .C2(n18720), .A(n18715), .B(n18714), .ZN(
        P3_U2946) );
  AOI22_X1 U21900 ( .A1(n18792), .A2(n18741), .B1(n18906), .B2(n18716), .ZN(
        n18719) );
  AOI22_X1 U21901 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18717), .B1(
        n18909), .B2(n18788), .ZN(n18718) );
  OAI211_X1 U21902 ( .C1(n18797), .C2(n18720), .A(n18719), .B(n18718), .ZN(
        P3_U2947) );
  INV_X1 U21903 ( .A(n18788), .ZN(n18796) );
  NOR2_X2 U21904 ( .A1(n18721), .A2(n18745), .ZN(n18820) );
  INV_X1 U21905 ( .A(n18820), .ZN(n18814) );
  AOI21_X1 U21906 ( .B1(n18796), .B2(n18814), .A(n18987), .ZN(n18740) );
  AOI22_X1 U21907 ( .A1(n18858), .A2(n18740), .B1(n18857), .B2(n18741), .ZN(
        n18726) );
  NOR2_X1 U21908 ( .A1(n18741), .A2(n18755), .ZN(n18723) );
  OAI211_X1 U21909 ( .C1(n18723), .C2(n18722), .A(n18796), .B(n18814), .ZN(
        n18724) );
  OAI211_X1 U21910 ( .C1(n18820), .C2(n19079), .A(n18771), .B(n18724), .ZN(
        n18742) );
  AOI22_X1 U21911 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18742), .B1(
        n18863), .B2(n18820), .ZN(n18725) );
  OAI211_X1 U21912 ( .C1(n18866), .C2(n18766), .A(n18726), .B(n18725), .ZN(
        P3_U2948) );
  AOI22_X1 U21913 ( .A1(n18868), .A2(n18755), .B1(n18867), .B2(n18740), .ZN(
        n18728) );
  AOI22_X1 U21914 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18742), .B1(
        n18869), .B2(n18820), .ZN(n18727) );
  OAI211_X1 U21915 ( .C1(n18872), .C2(n18737), .A(n18728), .B(n18727), .ZN(
        P3_U2949) );
  AOI22_X1 U21916 ( .A1(n18835), .A2(n18741), .B1(n18873), .B2(n18740), .ZN(
        n18730) );
  AOI22_X1 U21917 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18742), .B1(
        n18875), .B2(n18820), .ZN(n18729) );
  OAI211_X1 U21918 ( .C1(n18838), .C2(n18766), .A(n18730), .B(n18729), .ZN(
        P3_U2950) );
  AOI22_X1 U21919 ( .A1(n18839), .A2(n18755), .B1(n18879), .B2(n18740), .ZN(
        n18732) );
  AOI22_X1 U21920 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18742), .B1(
        n18881), .B2(n18820), .ZN(n18731) );
  OAI211_X1 U21921 ( .C1(n18842), .C2(n18737), .A(n18732), .B(n18731), .ZN(
        P3_U2951) );
  AOI22_X1 U21922 ( .A1(n18808), .A2(n18755), .B1(n18885), .B2(n18740), .ZN(
        n18734) );
  AOI22_X1 U21923 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18742), .B1(
        n18887), .B2(n18820), .ZN(n18733) );
  OAI211_X1 U21924 ( .C1(n18811), .C2(n18737), .A(n18734), .B(n18733), .ZN(
        P3_U2952) );
  AOI22_X1 U21925 ( .A1(n18892), .A2(n18755), .B1(n18891), .B2(n18740), .ZN(
        n18736) );
  AOI22_X1 U21926 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18742), .B1(
        n18893), .B2(n18820), .ZN(n18735) );
  OAI211_X1 U21927 ( .C1(n18896), .C2(n18737), .A(n18736), .B(n18735), .ZN(
        P3_U2953) );
  AOI22_X1 U21928 ( .A1(n18815), .A2(n18741), .B1(n18897), .B2(n18740), .ZN(
        n18739) );
  AOI22_X1 U21929 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18742), .B1(
        n18900), .B2(n18820), .ZN(n18738) );
  OAI211_X1 U21930 ( .C1(n18818), .C2(n18766), .A(n18739), .B(n18738), .ZN(
        P3_U2954) );
  AOI22_X1 U21931 ( .A1(n18908), .A2(n18741), .B1(n18906), .B2(n18740), .ZN(
        n18744) );
  AOI22_X1 U21932 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18742), .B1(
        n18909), .B2(n18820), .ZN(n18743) );
  OAI211_X1 U21933 ( .C1(n18914), .C2(n18766), .A(n18744), .B(n18743), .ZN(
        P3_U2955) );
  NOR2_X1 U21934 ( .A1(n18934), .A2(n18745), .ZN(n18799) );
  AND2_X1 U21935 ( .A1(n18856), .A2(n18799), .ZN(n18762) );
  AOI22_X1 U21936 ( .A1(n18858), .A2(n18762), .B1(n18857), .B2(n18755), .ZN(
        n18748) );
  AOI22_X1 U21937 ( .A1(n18862), .A2(n18746), .B1(n18859), .B2(n18799), .ZN(
        n18763) );
  NAND2_X1 U21938 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18799), .ZN(
        n18849) );
  INV_X1 U21939 ( .A(n18849), .ZN(n18851) );
  AOI22_X1 U21940 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18763), .B1(
        n18863), .B2(n18851), .ZN(n18747) );
  OAI211_X1 U21941 ( .C1(n18866), .C2(n18796), .A(n18748), .B(n18747), .ZN(
        P3_U2956) );
  AOI22_X1 U21942 ( .A1(n18868), .A2(n18788), .B1(n18867), .B2(n18762), .ZN(
        n18750) );
  AOI22_X1 U21943 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18763), .B1(
        n18869), .B2(n18851), .ZN(n18749) );
  OAI211_X1 U21944 ( .C1(n18872), .C2(n18766), .A(n18750), .B(n18749), .ZN(
        P3_U2957) );
  AOI22_X1 U21945 ( .A1(n18874), .A2(n18788), .B1(n18873), .B2(n18762), .ZN(
        n18752) );
  AOI22_X1 U21946 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18763), .B1(
        n18875), .B2(n18851), .ZN(n18751) );
  OAI211_X1 U21947 ( .C1(n18878), .C2(n18766), .A(n18752), .B(n18751), .ZN(
        P3_U2958) );
  AOI22_X1 U21948 ( .A1(n18880), .A2(n18755), .B1(n18879), .B2(n18762), .ZN(
        n18754) );
  AOI22_X1 U21949 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18763), .B1(
        n18881), .B2(n18851), .ZN(n18753) );
  OAI211_X1 U21950 ( .C1(n18884), .C2(n18796), .A(n18754), .B(n18753), .ZN(
        P3_U2959) );
  AOI22_X1 U21951 ( .A1(n18886), .A2(n18755), .B1(n18885), .B2(n18762), .ZN(
        n18757) );
  AOI22_X1 U21952 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18763), .B1(
        n18887), .B2(n18851), .ZN(n18756) );
  OAI211_X1 U21953 ( .C1(n18890), .C2(n18796), .A(n18757), .B(n18756), .ZN(
        P3_U2960) );
  AOI22_X1 U21954 ( .A1(n18892), .A2(n18788), .B1(n18891), .B2(n18762), .ZN(
        n18759) );
  AOI22_X1 U21955 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18763), .B1(
        n18893), .B2(n18851), .ZN(n18758) );
  OAI211_X1 U21956 ( .C1(n18896), .C2(n18766), .A(n18759), .B(n18758), .ZN(
        P3_U2961) );
  AOI22_X1 U21957 ( .A1(n18898), .A2(n18788), .B1(n18897), .B2(n18762), .ZN(
        n18761) );
  AOI22_X1 U21958 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18763), .B1(
        n18900), .B2(n18851), .ZN(n18760) );
  OAI211_X1 U21959 ( .C1(n18904), .C2(n18766), .A(n18761), .B(n18760), .ZN(
        P3_U2962) );
  AOI22_X1 U21960 ( .A1(n18792), .A2(n18788), .B1(n18906), .B2(n18762), .ZN(
        n18765) );
  AOI22_X1 U21961 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18763), .B1(
        n18909), .B2(n18851), .ZN(n18764) );
  OAI211_X1 U21962 ( .C1(n18797), .C2(n18766), .A(n18765), .B(n18764), .ZN(
        P3_U2963) );
  NAND2_X1 U21963 ( .A1(n18932), .A2(n18861), .ZN(n18903) );
  INV_X1 U21964 ( .A(n18903), .ZN(n18907) );
  INV_X1 U21965 ( .A(n18767), .ZN(n18769) );
  NOR2_X1 U21966 ( .A1(n18851), .A2(n18907), .ZN(n18827) );
  OAI21_X1 U21967 ( .B1(n18769), .B2(n18768), .A(n18827), .ZN(n18770) );
  OAI211_X1 U21968 ( .C1(n18907), .C2(n19079), .A(n18771), .B(n18770), .ZN(
        n18793) );
  NOR2_X1 U21969 ( .A1(n18987), .A2(n18827), .ZN(n18791) );
  AOI22_X1 U21970 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18793), .B1(
        n18858), .B2(n18791), .ZN(n18773) );
  AOI22_X1 U21971 ( .A1(n18825), .A2(n18820), .B1(n18863), .B2(n18907), .ZN(
        n18772) );
  OAI211_X1 U21972 ( .C1(n18832), .C2(n18796), .A(n18773), .B(n18772), .ZN(
        P3_U2964) );
  AOI22_X1 U21973 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18793), .B1(
        n18867), .B2(n18791), .ZN(n18776) );
  AOI22_X1 U21974 ( .A1(n18869), .A2(n18907), .B1(n18774), .B2(n18788), .ZN(
        n18775) );
  OAI211_X1 U21975 ( .C1(n18777), .C2(n18814), .A(n18776), .B(n18775), .ZN(
        P3_U2965) );
  AOI22_X1 U21976 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18793), .B1(
        n18873), .B2(n18791), .ZN(n18779) );
  AOI22_X1 U21977 ( .A1(n18874), .A2(n18820), .B1(n18875), .B2(n18907), .ZN(
        n18778) );
  OAI211_X1 U21978 ( .C1(n18878), .C2(n18796), .A(n18779), .B(n18778), .ZN(
        P3_U2966) );
  AOI22_X1 U21979 ( .A1(n18880), .A2(n18788), .B1(n18879), .B2(n18791), .ZN(
        n18781) );
  AOI22_X1 U21980 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18793), .B1(
        n18881), .B2(n18907), .ZN(n18780) );
  OAI211_X1 U21981 ( .C1(n18884), .C2(n18814), .A(n18781), .B(n18780), .ZN(
        P3_U2967) );
  AOI22_X1 U21982 ( .A1(n18808), .A2(n18820), .B1(n18885), .B2(n18791), .ZN(
        n18783) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18793), .B1(
        n18887), .B2(n18907), .ZN(n18782) );
  OAI211_X1 U21984 ( .C1(n18811), .C2(n18796), .A(n18783), .B(n18782), .ZN(
        P3_U2968) );
  AOI22_X1 U21985 ( .A1(n18784), .A2(n18788), .B1(n18891), .B2(n18791), .ZN(
        n18786) );
  AOI22_X1 U21986 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18793), .B1(
        n18893), .B2(n18907), .ZN(n18785) );
  OAI211_X1 U21987 ( .C1(n18787), .C2(n18814), .A(n18786), .B(n18785), .ZN(
        P3_U2969) );
  AOI22_X1 U21988 ( .A1(n18815), .A2(n18788), .B1(n18897), .B2(n18791), .ZN(
        n18790) );
  AOI22_X1 U21989 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18793), .B1(
        n18900), .B2(n18907), .ZN(n18789) );
  OAI211_X1 U21990 ( .C1(n18818), .C2(n18814), .A(n18790), .B(n18789), .ZN(
        P3_U2970) );
  AOI22_X1 U21991 ( .A1(n18792), .A2(n18820), .B1(n18906), .B2(n18791), .ZN(
        n18795) );
  AOI22_X1 U21992 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18793), .B1(
        n18909), .B2(n18907), .ZN(n18794) );
  OAI211_X1 U21993 ( .C1(n18797), .C2(n18796), .A(n18795), .B(n18794), .ZN(
        P3_U2971) );
  NOR2_X1 U21994 ( .A1(n18987), .A2(n18798), .ZN(n18819) );
  AOI22_X1 U21995 ( .A1(n18858), .A2(n18819), .B1(n18857), .B2(n18820), .ZN(
        n18801) );
  AOI22_X1 U21996 ( .A1(n18862), .A2(n18799), .B1(n18861), .B2(n18859), .ZN(
        n18821) );
  AOI22_X1 U21997 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18821), .B1(
        n18863), .B2(n18899), .ZN(n18800) );
  OAI211_X1 U21998 ( .C1(n18866), .C2(n18849), .A(n18801), .B(n18800), .ZN(
        P3_U2972) );
  AOI22_X1 U21999 ( .A1(n18868), .A2(n18851), .B1(n18867), .B2(n18819), .ZN(
        n18803) );
  AOI22_X1 U22000 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18869), .ZN(n18802) );
  OAI211_X1 U22001 ( .C1(n18872), .C2(n18814), .A(n18803), .B(n18802), .ZN(
        P3_U2973) );
  AOI22_X1 U22002 ( .A1(n18874), .A2(n18851), .B1(n18873), .B2(n18819), .ZN(
        n18805) );
  AOI22_X1 U22003 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18875), .ZN(n18804) );
  OAI211_X1 U22004 ( .C1(n18878), .C2(n18814), .A(n18805), .B(n18804), .ZN(
        P3_U2974) );
  AOI22_X1 U22005 ( .A1(n18880), .A2(n18820), .B1(n18879), .B2(n18819), .ZN(
        n18807) );
  AOI22_X1 U22006 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18881), .ZN(n18806) );
  OAI211_X1 U22007 ( .C1(n18884), .C2(n18849), .A(n18807), .B(n18806), .ZN(
        P3_U2975) );
  AOI22_X1 U22008 ( .A1(n18808), .A2(n18851), .B1(n18885), .B2(n18819), .ZN(
        n18810) );
  AOI22_X1 U22009 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18887), .ZN(n18809) );
  OAI211_X1 U22010 ( .C1(n18811), .C2(n18814), .A(n18810), .B(n18809), .ZN(
        P3_U2976) );
  AOI22_X1 U22011 ( .A1(n18892), .A2(n18851), .B1(n18891), .B2(n18819), .ZN(
        n18813) );
  AOI22_X1 U22012 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18893), .ZN(n18812) );
  OAI211_X1 U22013 ( .C1(n18896), .C2(n18814), .A(n18813), .B(n18812), .ZN(
        P3_U2977) );
  AOI22_X1 U22014 ( .A1(n18815), .A2(n18820), .B1(n18897), .B2(n18819), .ZN(
        n18817) );
  AOI22_X1 U22015 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18900), .ZN(n18816) );
  OAI211_X1 U22016 ( .C1(n18818), .C2(n18849), .A(n18817), .B(n18816), .ZN(
        P3_U2978) );
  AOI22_X1 U22017 ( .A1(n18908), .A2(n18820), .B1(n18906), .B2(n18819), .ZN(
        n18823) );
  AOI22_X1 U22018 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18821), .B1(
        n18899), .B2(n18909), .ZN(n18822) );
  OAI211_X1 U22019 ( .C1(n18914), .C2(n18849), .A(n18823), .B(n18822), .ZN(
        P3_U2979) );
  NOR2_X1 U22020 ( .A1(n18987), .A2(n18824), .ZN(n18850) );
  AOI22_X1 U22021 ( .A1(n18825), .A2(n18907), .B1(n18858), .B2(n18850), .ZN(
        n18831) );
  NOR2_X1 U22022 ( .A1(n18827), .A2(n18826), .ZN(n18828) );
  OAI22_X1 U22023 ( .A1(n18852), .A2(n19079), .B1(n18829), .B2(n18828), .ZN(
        n18853) );
  AOI22_X1 U22024 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18863), .ZN(n18830) );
  OAI211_X1 U22025 ( .C1(n18832), .C2(n18849), .A(n18831), .B(n18830), .ZN(
        P3_U2980) );
  AOI22_X1 U22026 ( .A1(n18868), .A2(n18907), .B1(n18867), .B2(n18850), .ZN(
        n18834) );
  AOI22_X1 U22027 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18869), .ZN(n18833) );
  OAI211_X1 U22028 ( .C1(n18872), .C2(n18849), .A(n18834), .B(n18833), .ZN(
        P3_U2981) );
  AOI22_X1 U22029 ( .A1(n18835), .A2(n18851), .B1(n18873), .B2(n18850), .ZN(
        n18837) );
  AOI22_X1 U22030 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18875), .ZN(n18836) );
  OAI211_X1 U22031 ( .C1(n18838), .C2(n18903), .A(n18837), .B(n18836), .ZN(
        P3_U2982) );
  AOI22_X1 U22032 ( .A1(n18839), .A2(n18907), .B1(n18879), .B2(n18850), .ZN(
        n18841) );
  AOI22_X1 U22033 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18881), .ZN(n18840) );
  OAI211_X1 U22034 ( .C1(n18842), .C2(n18849), .A(n18841), .B(n18840), .ZN(
        P3_U2983) );
  AOI22_X1 U22035 ( .A1(n18886), .A2(n18851), .B1(n18885), .B2(n18850), .ZN(
        n18844) );
  AOI22_X1 U22036 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18887), .ZN(n18843) );
  OAI211_X1 U22037 ( .C1(n18890), .C2(n18903), .A(n18844), .B(n18843), .ZN(
        P3_U2984) );
  AOI22_X1 U22038 ( .A1(n18892), .A2(n18907), .B1(n18891), .B2(n18850), .ZN(
        n18846) );
  AOI22_X1 U22039 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18893), .ZN(n18845) );
  OAI211_X1 U22040 ( .C1(n18896), .C2(n18849), .A(n18846), .B(n18845), .ZN(
        P3_U2985) );
  AOI22_X1 U22041 ( .A1(n18898), .A2(n18907), .B1(n18897), .B2(n18850), .ZN(
        n18848) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18900), .ZN(n18847) );
  OAI211_X1 U22043 ( .C1(n18904), .C2(n18849), .A(n18848), .B(n18847), .ZN(
        P3_U2986) );
  AOI22_X1 U22044 ( .A1(n18908), .A2(n18851), .B1(n18906), .B2(n18850), .ZN(
        n18855) );
  AOI22_X1 U22045 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18853), .B1(
        n18852), .B2(n18909), .ZN(n18854) );
  OAI211_X1 U22046 ( .C1(n18914), .C2(n18903), .A(n18855), .B(n18854), .ZN(
        P3_U2987) );
  AND2_X1 U22047 ( .A1(n18856), .A2(n18860), .ZN(n18905) );
  AOI22_X1 U22048 ( .A1(n18858), .A2(n18905), .B1(n18857), .B2(n18907), .ZN(
        n18865) );
  AOI22_X1 U22049 ( .A1(n18862), .A2(n18861), .B1(n18860), .B2(n18859), .ZN(
        n18911) );
  AOI22_X1 U22050 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18863), .ZN(n18864) );
  OAI211_X1 U22051 ( .C1(n18866), .C2(n18915), .A(n18865), .B(n18864), .ZN(
        P3_U2988) );
  AOI22_X1 U22052 ( .A1(n18899), .A2(n18868), .B1(n18867), .B2(n18905), .ZN(
        n18871) );
  AOI22_X1 U22053 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18869), .ZN(n18870) );
  OAI211_X1 U22054 ( .C1(n18872), .C2(n18903), .A(n18871), .B(n18870), .ZN(
        P3_U2989) );
  AOI22_X1 U22055 ( .A1(n18899), .A2(n18874), .B1(n18873), .B2(n18905), .ZN(
        n18877) );
  AOI22_X1 U22056 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18875), .ZN(n18876) );
  OAI211_X1 U22057 ( .C1(n18878), .C2(n18903), .A(n18877), .B(n18876), .ZN(
        P3_U2990) );
  AOI22_X1 U22058 ( .A1(n18880), .A2(n18907), .B1(n18879), .B2(n18905), .ZN(
        n18883) );
  AOI22_X1 U22059 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18881), .ZN(n18882) );
  OAI211_X1 U22060 ( .C1(n18915), .C2(n18884), .A(n18883), .B(n18882), .ZN(
        P3_U2991) );
  AOI22_X1 U22061 ( .A1(n18886), .A2(n18907), .B1(n18885), .B2(n18905), .ZN(
        n18889) );
  AOI22_X1 U22062 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18887), .ZN(n18888) );
  OAI211_X1 U22063 ( .C1(n18915), .C2(n18890), .A(n18889), .B(n18888), .ZN(
        P3_U2992) );
  AOI22_X1 U22064 ( .A1(n18899), .A2(n18892), .B1(n18891), .B2(n18905), .ZN(
        n18895) );
  AOI22_X1 U22065 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18893), .ZN(n18894) );
  OAI211_X1 U22066 ( .C1(n18896), .C2(n18903), .A(n18895), .B(n18894), .ZN(
        P3_U2993) );
  AOI22_X1 U22067 ( .A1(n18899), .A2(n18898), .B1(n18897), .B2(n18905), .ZN(
        n18902) );
  AOI22_X1 U22068 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18900), .ZN(n18901) );
  OAI211_X1 U22069 ( .C1(n18904), .C2(n18903), .A(n18902), .B(n18901), .ZN(
        P3_U2994) );
  AOI22_X1 U22070 ( .A1(n18908), .A2(n18907), .B1(n18906), .B2(n18905), .ZN(
        n18913) );
  AOI22_X1 U22071 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18911), .B1(
        n18910), .B2(n18909), .ZN(n18912) );
  OAI211_X1 U22072 ( .C1(n18915), .C2(n18914), .A(n18913), .B(n18912), .ZN(
        P3_U2995) );
  NOR2_X1 U22073 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18974) );
  NOR2_X1 U22074 ( .A1(n18916), .A2(n19109), .ZN(n18917) );
  OAI21_X1 U22075 ( .B1(n18917), .B2(n18922), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18927) );
  OAI21_X1 U22076 ( .B1(n18920), .B2(n18919), .A(n18918), .ZN(n18946) );
  OAI221_X1 U22077 ( .B1(n18946), .B2(n19103), .C1(n18946), .C2(n18922), .A(
        n18921), .ZN(n18926) );
  AOI21_X1 U22078 ( .B1(n19096), .B2(n19103), .A(n18923), .ZN(n18924) );
  AOI22_X1 U22079 ( .A1(n18963), .A2(n19091), .B1(n18924), .B2(n18948), .ZN(
        n18925) );
  OAI221_X1 U22080 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18927), 
        .C1(n19096), .C2(n18926), .A(n18925), .ZN(n19094) );
  AOI22_X1 U22081 ( .A1(n18966), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19094), .B2(n18945), .ZN(n18955) );
  INV_X1 U22082 ( .A(n18955), .ZN(n18939) );
  NOR2_X1 U22083 ( .A1(n18929), .A2(n18928), .ZN(n18931) );
  AOI22_X1 U22084 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18930), .B1(
        n18931), .B2(n19109), .ZN(n19105) );
  NOR2_X1 U22085 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18947), .ZN(
        n18942) );
  OAI22_X1 U22086 ( .A1(n18931), .A2(n19097), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18942), .ZN(n19101) );
  OR3_X1 U22087 ( .A1(n19105), .A2(n18934), .A3(n18932), .ZN(n18933) );
  AOI22_X1 U22088 ( .A1(n19105), .A2(n18934), .B1(n19101), .B2(n18933), .ZN(
        n18936) );
  OAI21_X1 U22089 ( .B1(n18966), .B2(n18936), .A(n18935), .ZN(n18937) );
  OAI21_X1 U22090 ( .B1(n18939), .B2(n18938), .A(n18937), .ZN(n18940) );
  OAI21_X1 U22091 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18955), .A(
        n18940), .ZN(n18973) );
  AOI21_X1 U22092 ( .B1(n18940), .B2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18941) );
  INV_X1 U22093 ( .A(n18941), .ZN(n18954) );
  INV_X1 U22094 ( .A(n18949), .ZN(n18944) );
  OAI22_X1 U22095 ( .A1(n18944), .A2(n18943), .B1(n18942), .B2(n18948), .ZN(
        n19081) );
  AOI21_X1 U22096 ( .B1(n18945), .B2(n19081), .A(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18953) );
  AOI21_X1 U22097 ( .B1(n18948), .B2(n18947), .A(n18946), .ZN(n18950) );
  OAI21_X1 U22098 ( .B1(n18951), .B2(n18950), .A(n18949), .ZN(n19084) );
  NOR3_X1 U22099 ( .A1(n18966), .A2(n19085), .A3(n19084), .ZN(n18952) );
  AOI211_X1 U22100 ( .C1(n18955), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        n18972) );
  OAI22_X1 U22101 ( .A1(n18959), .A2(n18958), .B1(n18957), .B2(n18956), .ZN(
        n18960) );
  AOI221_X1 U22102 ( .B1(n18963), .B2(n18962), .C1(n18961), .C2(n18962), .A(
        n18960), .ZN(n19124) );
  INV_X1 U22103 ( .A(n18964), .ZN(n18970) );
  AOI21_X1 U22104 ( .B1(n18966), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18965), .ZN(n18969) );
  OAI21_X1 U22105 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18967), .ZN(n18968) );
  NAND4_X1 U22106 ( .A1(n19124), .A2(n18970), .A3(n18969), .A4(n18968), .ZN(
        n18971) );
  AOI211_X1 U22107 ( .C1(n18974), .C2(n18973), .A(n18972), .B(n18971), .ZN(
        n18984) );
  NAND2_X1 U22108 ( .A1(n19088), .A2(n19143), .ZN(n18995) );
  INV_X1 U22109 ( .A(n18995), .ZN(n19136) );
  AOI22_X1 U22110 ( .A1(n19004), .A2(n17722), .B1(n19104), .B2(n19136), .ZN(
        n18975) );
  INV_X1 U22111 ( .A(n18975), .ZN(n18980) );
  OAI211_X1 U22112 ( .C1(n18977), .C2(n18976), .A(n19128), .B(n18984), .ZN(
        n19078) );
  NAND2_X1 U22113 ( .A1(n19004), .A2(n19143), .ZN(n18985) );
  NAND2_X1 U22114 ( .A1(n19078), .A2(n18985), .ZN(n18988) );
  NOR2_X1 U22115 ( .A1(n18978), .A2(n18988), .ZN(n18979) );
  MUX2_X1 U22116 ( .A(n18980), .B(n18979), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18982) );
  OAI211_X1 U22117 ( .C1(n18984), .C2(n18983), .A(n18982), .B(n18981), .ZN(
        P3_U2996) );
  NAND2_X1 U22118 ( .A1(n19004), .A2(n17722), .ZN(n18991) );
  OR3_X1 U22119 ( .A1(n19088), .A2(n18986), .A3(n18985), .ZN(n18993) );
  NAND4_X1 U22120 ( .A1(n18992), .A2(n18991), .A3(n18993), .A4(n18990), .ZN(
        P3_U2997) );
  AND4_X1 U22121 ( .A1(n18995), .A2(n18994), .A3(n18993), .A4(n19077), .ZN(
        P3_U2998) );
  INV_X1 U22122 ( .A(n19076), .ZN(n18996) );
  AND2_X1 U22123 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18996), .ZN(
        P3_U2999) );
  AND2_X1 U22124 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18996), .ZN(
        P3_U3000) );
  INV_X1 U22125 ( .A(P3_DATAWIDTH_REG_29__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U22126 ( .A1(n20898), .A2(n19076), .ZN(P3_U3001) );
  AND2_X1 U22127 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18996), .ZN(
        P3_U3002) );
  AND2_X1 U22128 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18996), .ZN(
        P3_U3003) );
  AND2_X1 U22129 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18996), .ZN(
        P3_U3004) );
  AND2_X1 U22130 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18996), .ZN(
        P3_U3005) );
  AND2_X1 U22131 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18996), .ZN(
        P3_U3006) );
  AND2_X1 U22132 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18996), .ZN(
        P3_U3007) );
  AND2_X1 U22133 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18996), .ZN(
        P3_U3008) );
  AND2_X1 U22134 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18996), .ZN(
        P3_U3009) );
  AND2_X1 U22135 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18996), .ZN(
        P3_U3010) );
  AND2_X1 U22136 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18996), .ZN(
        P3_U3011) );
  INV_X1 U22137 ( .A(P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20895) );
  NOR2_X1 U22138 ( .A1(n20895), .A2(n19076), .ZN(P3_U3012) );
  AND2_X1 U22139 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18996), .ZN(
        P3_U3013) );
  AND2_X1 U22140 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18996), .ZN(
        P3_U3014) );
  AND2_X1 U22141 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18996), .ZN(
        P3_U3015) );
  AND2_X1 U22142 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18996), .ZN(
        P3_U3016) );
  INV_X1 U22143 ( .A(P3_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20841) );
  NOR2_X1 U22144 ( .A1(n20841), .A2(n19076), .ZN(P3_U3017) );
  AND2_X1 U22145 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18996), .ZN(
        P3_U3018) );
  AND2_X1 U22146 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18996), .ZN(
        P3_U3019) );
  AND2_X1 U22147 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18996), .ZN(
        P3_U3020) );
  AND2_X1 U22148 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18996), .ZN(P3_U3021) );
  AND2_X1 U22149 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18996), .ZN(P3_U3022) );
  AND2_X1 U22150 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18996), .ZN(P3_U3023) );
  AND2_X1 U22151 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18996), .ZN(P3_U3024) );
  AND2_X1 U22152 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18996), .ZN(P3_U3025) );
  AND2_X1 U22153 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18996), .ZN(P3_U3026) );
  AND2_X1 U22154 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18996), .ZN(P3_U3027) );
  AND2_X1 U22155 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18996), .ZN(P3_U3028) );
  OAI21_X1 U22156 ( .B1(n18997), .B2(n20624), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18998) );
  AOI22_X1 U22157 ( .A1(n19012), .A2(n19014), .B1(n19141), .B2(n18998), .ZN(
        n19000) );
  INV_X1 U22158 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18999) );
  NAND3_X1 U22159 ( .A1(NA), .A2(n19012), .A3(n18999), .ZN(n19007) );
  OAI211_X1 U22160 ( .C1(n19133), .C2(n19001), .A(n19000), .B(n19007), .ZN(
        P3_U3029) );
  NOR2_X1 U22161 ( .A1(n19014), .A2(n20624), .ZN(n19010) );
  INV_X1 U22162 ( .A(n19010), .ZN(n19003) );
  INV_X1 U22163 ( .A(n19001), .ZN(n19002) );
  AOI22_X1 U22164 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n19003), .B1(HOLD), 
        .B2(n19002), .ZN(n19005) );
  NAND2_X1 U22165 ( .A1(n19004), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19008) );
  OAI211_X1 U22166 ( .C1(n19005), .C2(n19012), .A(n19008), .B(n19130), .ZN(
        P3_U3030) );
  INV_X1 U22167 ( .A(n19008), .ZN(n19006) );
  AOI21_X1 U22168 ( .B1(n19012), .B2(n19007), .A(n19006), .ZN(n19013) );
  OAI22_X1 U22169 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n19008), .ZN(n19009) );
  OAI22_X1 U22170 ( .A1(n19010), .A2(n19009), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19011) );
  OAI22_X1 U22171 ( .A1(n19013), .A2(n19014), .B1(n19012), .B2(n19011), .ZN(
        P3_U3031) );
  OAI222_X1 U22172 ( .A1(n19121), .A2(n19067), .B1(n19015), .B2(n19069), .C1(
        n19016), .C2(n19072), .ZN(P3_U3032) );
  OAI222_X1 U22173 ( .A1(n19072), .A2(n19019), .B1(n19017), .B2(n19069), .C1(
        n19016), .C2(n19067), .ZN(P3_U3033) );
  OAI222_X1 U22174 ( .A1(n19067), .A2(n19019), .B1(n19018), .B2(n19069), .C1(
        n20983), .C2(n19072), .ZN(P3_U3034) );
  OAI222_X1 U22175 ( .A1(n19072), .A2(n19022), .B1(n19020), .B2(n19069), .C1(
        n20983), .C2(n19067), .ZN(P3_U3035) );
  OAI222_X1 U22176 ( .A1(n19022), .A2(n19067), .B1(n19021), .B2(n19069), .C1(
        n19023), .C2(n19072), .ZN(P3_U3036) );
  OAI222_X1 U22177 ( .A1(n19072), .A2(n19025), .B1(n19024), .B2(n19069), .C1(
        n19023), .C2(n19067), .ZN(P3_U3037) );
  INV_X1 U22178 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19028) );
  OAI222_X1 U22179 ( .A1(n19072), .A2(n19028), .B1(n19026), .B2(n19069), .C1(
        n19025), .C2(n19067), .ZN(P3_U3038) );
  OAI222_X1 U22180 ( .A1(n19028), .A2(n19067), .B1(n19027), .B2(n19069), .C1(
        n19029), .C2(n19072), .ZN(P3_U3039) );
  OAI222_X1 U22181 ( .A1(n19072), .A2(n19032), .B1(n19030), .B2(n19069), .C1(
        n19029), .C2(n19067), .ZN(P3_U3040) );
  OAI222_X1 U22182 ( .A1(n19067), .A2(n19032), .B1(n19031), .B2(n19069), .C1(
        n20772), .C2(n19072), .ZN(P3_U3041) );
  OAI222_X1 U22183 ( .A1(n19072), .A2(n19034), .B1(n19033), .B2(n19069), .C1(
        n20772), .C2(n19067), .ZN(P3_U3042) );
  OAI222_X1 U22184 ( .A1(n19072), .A2(n19036), .B1(n19035), .B2(n19069), .C1(
        n19034), .C2(n19067), .ZN(P3_U3043) );
  INV_X1 U22185 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19038) );
  OAI222_X1 U22186 ( .A1(n19072), .A2(n19038), .B1(n19037), .B2(n19069), .C1(
        n19036), .C2(n19067), .ZN(P3_U3044) );
  OAI222_X1 U22187 ( .A1(n19072), .A2(n19039), .B1(n20753), .B2(n19069), .C1(
        n19038), .C2(n19067), .ZN(P3_U3045) );
  OAI222_X1 U22188 ( .A1(n19072), .A2(n19041), .B1(n19040), .B2(n19069), .C1(
        n19039), .C2(n19067), .ZN(P3_U3046) );
  INV_X1 U22189 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19044) );
  OAI222_X1 U22190 ( .A1(n19072), .A2(n19044), .B1(n19042), .B2(n19069), .C1(
        n19041), .C2(n19067), .ZN(P3_U3047) );
  OAI222_X1 U22191 ( .A1(n19044), .A2(n19067), .B1(n19043), .B2(n19069), .C1(
        n19045), .C2(n19072), .ZN(P3_U3048) );
  OAI222_X1 U22192 ( .A1(n19072), .A2(n19047), .B1(n19046), .B2(n19069), .C1(
        n19045), .C2(n19067), .ZN(P3_U3049) );
  OAI222_X1 U22193 ( .A1(n19072), .A2(n19049), .B1(n19048), .B2(n19069), .C1(
        n19047), .C2(n19067), .ZN(P3_U3050) );
  OAI222_X1 U22194 ( .A1(n19072), .A2(n19051), .B1(n19050), .B2(n19069), .C1(
        n19049), .C2(n19067), .ZN(P3_U3051) );
  OAI222_X1 U22195 ( .A1(n19072), .A2(n19053), .B1(n19052), .B2(n19069), .C1(
        n19051), .C2(n19067), .ZN(P3_U3052) );
  OAI222_X1 U22196 ( .A1(n19072), .A2(n19055), .B1(n19054), .B2(n19069), .C1(
        n19053), .C2(n19067), .ZN(P3_U3053) );
  OAI222_X1 U22197 ( .A1(n19072), .A2(n19056), .B1(n20738), .B2(n19069), .C1(
        n19055), .C2(n19067), .ZN(P3_U3054) );
  OAI222_X1 U22198 ( .A1(n19072), .A2(n19058), .B1(n19057), .B2(n19069), .C1(
        n19056), .C2(n19067), .ZN(P3_U3055) );
  OAI222_X1 U22199 ( .A1(n19072), .A2(n19060), .B1(n19059), .B2(n19069), .C1(
        n19058), .C2(n19067), .ZN(P3_U3056) );
  OAI222_X1 U22200 ( .A1(n19060), .A2(n19067), .B1(n20940), .B2(n19069), .C1(
        n19062), .C2(n19072), .ZN(P3_U3057) );
  OAI222_X1 U22201 ( .A1(n19067), .A2(n19062), .B1(n19061), .B2(n19069), .C1(
        n19063), .C2(n19072), .ZN(P3_U3058) );
  OAI222_X1 U22202 ( .A1(n19072), .A2(n19065), .B1(n19064), .B2(n19069), .C1(
        n19063), .C2(n19067), .ZN(P3_U3059) );
  OAI222_X1 U22203 ( .A1(n19072), .A2(n19068), .B1(n19066), .B2(n19069), .C1(
        n19065), .C2(n19067), .ZN(P3_U3060) );
  OAI222_X1 U22204 ( .A1(n19072), .A2(n19071), .B1(n19070), .B2(n19069), .C1(
        n19068), .C2(n19067), .ZN(P3_U3061) );
  MUX2_X1 U22205 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n19141), .Z(P3_U3274) );
  MUX2_X1 U22206 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n19141), .Z(P3_U3275) );
  MUX2_X1 U22207 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(P3_BE_N_REG_1__SCAN_IN), .S(n19141), .Z(P3_U3276) );
  MUX2_X1 U22208 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .B(P3_BE_N_REG_0__SCAN_IN), .S(n19141), .Z(P3_U3277) );
  OAI21_X1 U22209 ( .B1(n19076), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19074), 
        .ZN(n19073) );
  INV_X1 U22210 ( .A(n19073), .ZN(P3_U3280) );
  INV_X1 U22211 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19075) );
  OAI21_X1 U22212 ( .B1(n19076), .B2(n19075), .A(n19074), .ZN(P3_U3281) );
  OAI221_X1 U22213 ( .B1(n19079), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19079), 
        .C2(n19078), .A(n19077), .ZN(P3_U3282) );
  NOR2_X1 U22214 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n19080), .ZN(
        n19082) );
  AOI22_X1 U22215 ( .A1(n19104), .A2(n19083), .B1(n19082), .B2(n19081), .ZN(
        n19087) );
  AOI21_X1 U22216 ( .B1(n19144), .B2(n19084), .A(n19110), .ZN(n19086) );
  OAI22_X1 U22217 ( .A1(n19110), .A2(n19087), .B1(n19086), .B2(n19085), .ZN(
        P3_U3285) );
  NOR2_X1 U22218 ( .A1(n19088), .A2(n19106), .ZN(n19098) );
  OAI22_X1 U22219 ( .A1(n19090), .A2(n19089), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19099) );
  INV_X1 U22220 ( .A(n19099), .ZN(n19093) );
  INV_X1 U22221 ( .A(n19091), .ZN(n19092) );
  AOI222_X1 U22222 ( .A1(n19094), .A2(n19144), .B1(n19098), .B2(n19093), .C1(
        n19104), .C2(n19092), .ZN(n19095) );
  AOI22_X1 U22223 ( .A1(n19110), .A2(n19096), .B1(n19095), .B2(n19107), .ZN(
        P3_U3288) );
  INV_X1 U22224 ( .A(n19097), .ZN(n19100) );
  AOI222_X1 U22225 ( .A1(n19101), .A2(n19144), .B1(n19104), .B2(n19100), .C1(
        n19099), .C2(n19098), .ZN(n19102) );
  AOI22_X1 U22226 ( .A1(n19110), .A2(n19103), .B1(n19102), .B2(n19107), .ZN(
        P3_U3289) );
  AOI222_X1 U22227 ( .A1(n19106), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19144), 
        .B2(n19105), .C1(n19109), .C2(n19104), .ZN(n19108) );
  AOI22_X1 U22228 ( .A1(n19110), .A2(n19109), .B1(n19108), .B2(n19107), .ZN(
        P3_U3290) );
  NOR2_X1 U22229 ( .A1(P3_DATAWIDTH_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19112) );
  AOI211_X1 U22230 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(n20771), .A(n19112), 
        .B(n19111), .ZN(n19116) );
  NOR2_X1 U22231 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n19121), .ZN(n19114) );
  INV_X1 U22232 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19113) );
  MUX2_X1 U22233 ( .A(n19114), .B(n19113), .S(n19120), .Z(n19115) );
  NOR2_X1 U22234 ( .A1(n19116), .A2(n19115), .ZN(P3_U3292) );
  OAI21_X1 U22235 ( .B1(n19118), .B2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n19117), 
        .ZN(n19119) );
  OAI21_X1 U22236 ( .B1(n19121), .B2(n19120), .A(n19119), .ZN(P3_U3293) );
  INV_X1 U22237 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n20751) );
  AOI22_X1 U22238 ( .A1(n19069), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n20751), 
        .B2(n19141), .ZN(P3_U3294) );
  INV_X1 U22239 ( .A(n19122), .ZN(n19125) );
  NAND2_X1 U22240 ( .A1(n19125), .A2(P3_MORE_REG_SCAN_IN), .ZN(n19123) );
  OAI21_X1 U22241 ( .B1(n19125), .B2(n19124), .A(n19123), .ZN(P3_U3295) );
  OAI21_X1 U22242 ( .B1(n19128), .B2(n19127), .A(n19126), .ZN(n19129) );
  AOI21_X1 U22243 ( .B1(n17722), .B2(n19133), .A(n19129), .ZN(n19140) );
  AOI21_X1 U22244 ( .B1(n19132), .B2(n19131), .A(n19130), .ZN(n19134) );
  OAI211_X1 U22245 ( .C1(n19135), .C2(n19134), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19133), .ZN(n19137) );
  AOI21_X1 U22246 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19137), .A(n19136), 
        .ZN(n19139) );
  NAND2_X1 U22247 ( .A1(n19140), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19138) );
  OAI21_X1 U22248 ( .B1(n19140), .B2(n19139), .A(n19138), .ZN(P3_U3296) );
  OAI22_X1 U22249 ( .A1(n19141), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n19069), .ZN(n19142) );
  INV_X1 U22250 ( .A(n19142), .ZN(P3_U3297) );
  AOI21_X1 U22251 ( .B1(n19144), .B2(n19143), .A(n19146), .ZN(n19149) );
  INV_X1 U22252 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n20851) );
  AOI22_X1 U22253 ( .A1(n19146), .A2(n19145), .B1(n19149), .B2(n20851), .ZN(
        P3_U3298) );
  INV_X1 U22254 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19148) );
  AOI21_X1 U22255 ( .B1(n19149), .B2(n19148), .A(n19147), .ZN(P3_U3299) );
  INV_X1 U22256 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20079) );
  NAND2_X1 U22257 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20079), .ZN(n20070) );
  AOI22_X1 U22258 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20070), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n20061), .ZN(n20128) );
  AOI21_X1 U22259 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20128), .ZN(n19150) );
  INV_X1 U22260 ( .A(n19150), .ZN(P2_U2815) );
  NOR2_X1 U22261 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19151), .ZN(n20054) );
  AOI22_X1 U22262 ( .A1(n19153), .A2(n20054), .B1(P2_CODEFETCH_REG_SCAN_IN), 
        .B2(n19152), .ZN(n19154) );
  INV_X1 U22263 ( .A(n19154), .ZN(P2_U2816) );
  AOI21_X1 U22264 ( .B1(n20061), .B2(n20079), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n19155) );
  AOI22_X1 U22265 ( .A1(n20193), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n19155), 
        .B2(n20194), .ZN(P2_U2817) );
  OAI21_X1 U22266 ( .B1(n20062), .B2(BS16), .A(n20128), .ZN(n20126) );
  OAI21_X1 U22267 ( .B1(n20128), .B2(n13249), .A(n20126), .ZN(P2_U2818) );
  NOR4_X1 U22268 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19165) );
  NOR4_X1 U22269 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_6__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19164) );
  AOI211_X1 U22270 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19156) );
  INV_X1 U22271 ( .A(P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20741) );
  INV_X1 U22272 ( .A(P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20731) );
  NAND3_X1 U22273 ( .A1(n19156), .A2(n20741), .A3(n20731), .ZN(n19162) );
  NOR4_X1 U22274 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19160) );
  NOR4_X1 U22275 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19159) );
  NOR4_X1 U22276 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19158) );
  NOR4_X1 U22277 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19157) );
  NAND4_X1 U22278 ( .A1(n19160), .A2(n19159), .A3(n19158), .A4(n19157), .ZN(
        n19161) );
  NOR4_X1 U22279 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(n19162), .A4(n19161), .ZN(n19163) );
  NAND3_X1 U22280 ( .A1(n19165), .A2(n19164), .A3(n19163), .ZN(n19173) );
  NOR2_X1 U22281 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19173), .ZN(n19168) );
  INV_X1 U22282 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19166) );
  AOI22_X1 U22283 ( .A1(n19168), .A2(n10985), .B1(n19173), .B2(n19166), .ZN(
        P2_U2820) );
  OR3_X1 U22284 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19172) );
  INV_X1 U22285 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19167) );
  AOI22_X1 U22286 ( .A1(n19168), .A2(n19172), .B1(n19173), .B2(n19167), .ZN(
        P2_U2821) );
  INV_X1 U22287 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20127) );
  NAND2_X1 U22288 ( .A1(n19168), .A2(n20127), .ZN(n19171) );
  INV_X1 U22289 ( .A(n19173), .ZN(n19175) );
  OAI21_X1 U22290 ( .B1(n10985), .B2(n10986), .A(n19175), .ZN(n19169) );
  OAI21_X1 U22291 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19175), .A(n19169), 
        .ZN(n19170) );
  OAI221_X1 U22292 ( .B1(n19171), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19171), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19170), .ZN(P2_U2822) );
  INV_X1 U22293 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19174) );
  OAI221_X1 U22294 ( .B1(n19175), .B2(n19174), .C1(n19173), .C2(n19172), .A(
        n19171), .ZN(P2_U2823) );
  INV_X1 U22295 ( .A(n19179), .ZN(n19176) );
  AOI22_X1 U22296 ( .A1(n19177), .A2(n19341), .B1(n19176), .B2(n19350), .ZN(
        n19186) );
  INV_X1 U22297 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n20868) );
  OAI22_X1 U22298 ( .A1(n20868), .A2(n19306), .B1(n20103), .B2(n19305), .ZN(
        n19183) );
  OAI21_X1 U22299 ( .B1(n19180), .B2(n19179), .A(n19178), .ZN(n19181) );
  OAI22_X1 U22300 ( .A1(n19324), .A2(n20999), .B1(n19354), .B2(n19181), .ZN(
        n19182) );
  AOI211_X1 U22301 ( .C1(n19315), .C2(n19184), .A(n19183), .B(n19182), .ZN(
        n19185) );
  OAI211_X1 U22302 ( .C1(n19187), .C2(n19323), .A(n19186), .B(n19185), .ZN(
        P2_U2835) );
  NAND2_X1 U22303 ( .A1(n15347), .A2(n19188), .ZN(n19189) );
  XOR2_X1 U22304 ( .A(n19190), .B(n19189), .Z(n19200) );
  INV_X1 U22305 ( .A(n19191), .ZN(n19193) );
  AOI22_X1 U22306 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19351), .B1(
        P2_EBX_REG_19__SCAN_IN), .B2(n19342), .ZN(n19192) );
  OAI21_X1 U22307 ( .B1(n19193), .B2(n19308), .A(n19192), .ZN(n19194) );
  AOI211_X1 U22308 ( .C1(P2_REIP_REG_19__SCAN_IN), .C2(n19343), .A(n19326), 
        .B(n19194), .ZN(n19199) );
  INV_X1 U22309 ( .A(n19195), .ZN(n19197) );
  AOI22_X1 U22310 ( .A1(n19197), .A2(n19315), .B1(n19196), .B2(n19339), .ZN(
        n19198) );
  OAI211_X1 U22311 ( .C1(n20056), .C2(n19200), .A(n19199), .B(n19198), .ZN(
        P2_U2836) );
  OAI21_X1 U22312 ( .B1(n20099), .B2(n19305), .A(n19304), .ZN(n19205) );
  INV_X1 U22313 ( .A(n19201), .ZN(n19203) );
  OAI22_X1 U22314 ( .A1(n19203), .A2(n19308), .B1(n19202), .B2(n19324), .ZN(
        n19204) );
  AOI211_X1 U22315 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19351), .A(
        n19205), .B(n19204), .ZN(n19212) );
  INV_X1 U22316 ( .A(n19206), .ZN(n19210) );
  XNOR2_X1 U22317 ( .A(n19208), .B(n19207), .ZN(n19209) );
  AOI22_X1 U22318 ( .A1(n19210), .A2(n19315), .B1(n19316), .B2(n19209), .ZN(
        n19211) );
  OAI211_X1 U22319 ( .C1(n19213), .C2(n19323), .A(n19212), .B(n19211), .ZN(
        P2_U2837) );
  OAI21_X1 U22320 ( .B1(n20808), .B2(n19305), .A(n19304), .ZN(n19216) );
  OAI22_X1 U22321 ( .A1(n19214), .A2(n19308), .B1(n19324), .B2(n10660), .ZN(
        n19215) );
  AOI211_X1 U22322 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19351), .A(
        n19216), .B(n19215), .ZN(n19223) );
  NOR2_X1 U22323 ( .A1(n19331), .A2(n19217), .ZN(n19219) );
  XNOR2_X1 U22324 ( .A(n19219), .B(n19218), .ZN(n19221) );
  AOI22_X1 U22325 ( .A1(n19221), .A2(n19316), .B1(n19220), .B2(n19315), .ZN(
        n19222) );
  OAI211_X1 U22326 ( .C1(n19224), .C2(n19323), .A(n19223), .B(n19222), .ZN(
        P2_U2839) );
  NAND2_X1 U22327 ( .A1(n15347), .A2(n19225), .ZN(n19227) );
  XOR2_X1 U22328 ( .A(n19227), .B(n19226), .Z(n19236) );
  OAI22_X1 U22329 ( .A1(n19229), .A2(n19308), .B1(n19306), .B2(n19228), .ZN(
        n19230) );
  INV_X1 U22330 ( .A(n19230), .ZN(n19231) );
  OAI211_X1 U22331 ( .C1(n20910), .C2(n19305), .A(n19231), .B(n19304), .ZN(
        n19234) );
  OAI22_X1 U22332 ( .A1(n19232), .A2(n19346), .B1(n19362), .B2(n19323), .ZN(
        n19233) );
  AOI211_X1 U22333 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19342), .A(n19234), .B(
        n19233), .ZN(n19235) );
  OAI21_X1 U22334 ( .B1(n19236), .B2(n20056), .A(n19235), .ZN(P2_U2840) );
  AOI22_X1 U22335 ( .A1(n19237), .A2(n19341), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19342), .ZN(n19238) );
  OAI211_X1 U22336 ( .C1(n11129), .C2(n19305), .A(n19238), .B(n19304), .ZN(
        n19239) );
  AOI21_X1 U22337 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19351), .A(
        n19239), .ZN(n19246) );
  NOR2_X1 U22338 ( .A1(n19331), .A2(n19240), .ZN(n19242) );
  XNOR2_X1 U22339 ( .A(n19242), .B(n19241), .ZN(n19244) );
  AOI22_X1 U22340 ( .A1(n19244), .A2(n19316), .B1(n19243), .B2(n19315), .ZN(
        n19245) );
  OAI211_X1 U22341 ( .C1(n19364), .C2(n19323), .A(n19246), .B(n19245), .ZN(
        P2_U2841) );
  INV_X1 U22342 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19247) );
  OAI22_X1 U22343 ( .A1(n19248), .A2(n19308), .B1(n19324), .B2(n19247), .ZN(
        n19249) );
  INV_X1 U22344 ( .A(n19249), .ZN(n19250) );
  OAI211_X1 U22345 ( .C1(n11097), .C2(n19305), .A(n19250), .B(n19304), .ZN(
        n19251) );
  AOI21_X1 U22346 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19351), .A(
        n19251), .ZN(n19259) );
  NOR2_X1 U22347 ( .A1(n19331), .A2(n19252), .ZN(n19254) );
  XNOR2_X1 U22348 ( .A(n19254), .B(n19253), .ZN(n19257) );
  INV_X1 U22349 ( .A(n19255), .ZN(n19256) );
  AOI22_X1 U22350 ( .A1(n19257), .A2(n19316), .B1(n19256), .B2(n19315), .ZN(
        n19258) );
  OAI211_X1 U22351 ( .C1(n19369), .C2(n19323), .A(n19259), .B(n19258), .ZN(
        P2_U2843) );
  NOR2_X1 U22352 ( .A1(n19331), .A2(n19260), .ZN(n19262) );
  XOR2_X1 U22353 ( .A(n19262), .B(n19261), .Z(n19273) );
  INV_X1 U22354 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n19263) );
  OAI22_X1 U22355 ( .A1(n19264), .A2(n19308), .B1(n19324), .B2(n19263), .ZN(
        n19265) );
  INV_X1 U22356 ( .A(n19265), .ZN(n19266) );
  OAI211_X1 U22357 ( .C1(n11067), .C2(n19305), .A(n19266), .B(n19304), .ZN(
        n19267) );
  AOI21_X1 U22358 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19351), .A(
        n19267), .ZN(n19272) );
  INV_X1 U22359 ( .A(n19268), .ZN(n19270) );
  AOI22_X1 U22360 ( .A1(n19270), .A2(n19315), .B1(n19339), .B2(n19269), .ZN(
        n19271) );
  OAI211_X1 U22361 ( .C1(n20056), .C2(n19273), .A(n19272), .B(n19271), .ZN(
        P2_U2845) );
  NAND2_X1 U22362 ( .A1(n15347), .A2(n19274), .ZN(n19276) );
  XOR2_X1 U22363 ( .A(n19276), .B(n19275), .Z(n19283) );
  AOI22_X1 U22364 ( .A1(n19277), .A2(n19341), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19351), .ZN(n19278) );
  OAI211_X1 U22365 ( .C1(n11054), .C2(n19305), .A(n19278), .B(n19304), .ZN(
        n19281) );
  OAI22_X1 U22366 ( .A1(n19279), .A2(n19346), .B1(n19323), .B2(n19379), .ZN(
        n19280) );
  AOI211_X1 U22367 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19342), .A(n19281), .B(
        n19280), .ZN(n19282) );
  OAI21_X1 U22368 ( .B1(n19283), .B2(n20056), .A(n19282), .ZN(P2_U2846) );
  AOI22_X1 U22369 ( .A1(n19284), .A2(n19341), .B1(n19342), .B2(
        P2_EBX_REG_8__SCAN_IN), .ZN(n19285) );
  OAI211_X1 U22370 ( .C1(n11037), .C2(n19305), .A(n19285), .B(n19304), .ZN(
        n19286) );
  AOI21_X1 U22371 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19351), .A(
        n19286), .ZN(n19293) );
  NOR2_X1 U22372 ( .A1(n19331), .A2(n19287), .ZN(n19289) );
  XNOR2_X1 U22373 ( .A(n19289), .B(n19288), .ZN(n19291) );
  AOI22_X1 U22374 ( .A1(n19291), .A2(n19316), .B1(n19315), .B2(n19290), .ZN(
        n19292) );
  OAI211_X1 U22375 ( .C1(n19323), .C2(n19381), .A(n19293), .B(n19292), .ZN(
        P2_U2847) );
  NAND2_X1 U22376 ( .A1(n15347), .A2(n19294), .ZN(n19296) );
  XOR2_X1 U22377 ( .A(n19296), .B(n19295), .Z(n19303) );
  AOI22_X1 U22378 ( .A1(n19341), .A2(n19297), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19351), .ZN(n19298) );
  OAI211_X1 U22379 ( .C1(n10858), .C2(n19305), .A(n19298), .B(n19304), .ZN(
        n19301) );
  OAI22_X1 U22380 ( .A1(n19383), .A2(n19323), .B1(n19346), .B2(n19299), .ZN(
        n19300) );
  AOI211_X1 U22381 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19342), .A(n19301), .B(
        n19300), .ZN(n19302) );
  OAI21_X1 U22382 ( .B1(n19303), .B2(n20056), .A(n19302), .ZN(P2_U2848) );
  OAI21_X1 U22383 ( .B1(n14014), .B2(n19305), .A(n19304), .ZN(n19310) );
  OAI22_X1 U22384 ( .A1(n19308), .A2(n19307), .B1(n19306), .B2(n10012), .ZN(
        n19309) );
  AOI211_X1 U22385 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19342), .A(n19310), .B(
        n19309), .ZN(n19319) );
  NOR2_X1 U22386 ( .A1(n19331), .A2(n19311), .ZN(n19313) );
  XNOR2_X1 U22387 ( .A(n19313), .B(n19312), .ZN(n19317) );
  AOI22_X1 U22388 ( .A1(n19317), .A2(n19316), .B1(n19315), .B2(n19314), .ZN(
        n19318) );
  OAI211_X1 U22389 ( .C1(n19323), .C2(n19386), .A(n19319), .B(n19318), .ZN(
        P2_U2849) );
  INV_X1 U22390 ( .A(n19320), .ZN(n19321) );
  AOI22_X1 U22391 ( .A1(n19341), .A2(n19321), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19351), .ZN(n19338) );
  OAI22_X1 U22392 ( .A1(n19324), .A2(n10525), .B1(n19323), .B2(n19322), .ZN(
        n19325) );
  AOI211_X1 U22393 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19343), .A(n19326), .B(
        n19325), .ZN(n19337) );
  OAI22_X1 U22394 ( .A1(n19391), .A2(n19328), .B1(n19346), .B2(n19327), .ZN(
        n19329) );
  INV_X1 U22395 ( .A(n19329), .ZN(n19336) );
  INV_X1 U22396 ( .A(n19470), .ZN(n19334) );
  NOR2_X1 U22397 ( .A1(n19331), .A2(n19330), .ZN(n19333) );
  AOI21_X1 U22398 ( .B1(n19334), .B2(n19333), .A(n20056), .ZN(n19332) );
  OAI21_X1 U22399 ( .B1(n19334), .B2(n19333), .A(n19332), .ZN(n19335) );
  NAND4_X1 U22400 ( .A1(n19338), .A2(n19337), .A3(n19336), .A4(n19335), .ZN(
        P2_U2851) );
  AOI22_X1 U22401 ( .A1(n19341), .A2(n19340), .B1(n19339), .B2(n19419), .ZN(
        n19345) );
  AOI22_X1 U22402 ( .A1(n19343), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19342), 
        .B2(P2_EBX_REG_0__SCAN_IN), .ZN(n19344) );
  OAI211_X1 U22403 ( .C1(n19347), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        n19348) );
  AOI21_X1 U22404 ( .B1(n19548), .B2(n19349), .A(n19348), .ZN(n19353) );
  OAI21_X1 U22405 ( .B1(n19351), .B2(n19350), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19352) );
  OAI211_X1 U22406 ( .C1(n19355), .C2(n19354), .A(n19353), .B(n19352), .ZN(
        P2_U2855) );
  AOI22_X1 U22407 ( .A1(n14453), .A2(n19416), .B1(n19356), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19359) );
  AOI22_X1 U22408 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n19357), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19415), .ZN(n19358) );
  NAND2_X1 U22409 ( .A1(n19359), .A2(n19358), .ZN(P2_U2888) );
  INV_X1 U22410 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19430) );
  OAI222_X1 U22411 ( .A1(n19430), .A2(n19387), .B1(n19362), .B2(n19385), .C1(
        n19361), .C2(n19422), .ZN(P2_U2904) );
  INV_X1 U22412 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19432) );
  OAI222_X1 U22413 ( .A1(n19432), .A2(n19387), .B1(n19364), .B2(n19385), .C1(
        n19422), .C2(n19363), .ZN(P2_U2905) );
  INV_X1 U22414 ( .A(n19385), .ZN(n19388) );
  AOI22_X1 U22415 ( .A1(n19366), .A2(n19388), .B1(n19365), .B2(n19376), .ZN(
        n19367) );
  OAI21_X1 U22416 ( .B1(n19387), .B2(n20804), .A(n19367), .ZN(P2_U2906) );
  INV_X1 U22417 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19370) );
  OAI222_X1 U22418 ( .A1(n19370), .A2(n19387), .B1(n19369), .B2(n19385), .C1(
        n19422), .C2(n19368), .ZN(P2_U2907) );
  AOI22_X1 U22419 ( .A1(n19372), .A2(n19388), .B1(n19371), .B2(n19376), .ZN(
        n19373) );
  OAI21_X1 U22420 ( .B1(n19387), .B2(n19436), .A(n19373), .ZN(P2_U2908) );
  INV_X1 U22421 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n20759) );
  OAI222_X1 U22422 ( .A1(n20759), .A2(n19387), .B1(n19375), .B2(n19385), .C1(
        n19422), .C2(n19374), .ZN(P2_U2909) );
  AOI22_X1 U22423 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n19415), .B1(n19377), .B2(
        n19376), .ZN(n19378) );
  OAI21_X1 U22424 ( .B1(n19385), .B2(n19379), .A(n19378), .ZN(P2_U2910) );
  INV_X1 U22425 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19441) );
  OAI222_X1 U22426 ( .A1(n19441), .A2(n19387), .B1(n19381), .B2(n19385), .C1(
        n19422), .C2(n19380), .ZN(P2_U2911) );
  INV_X1 U22427 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19443) );
  OAI222_X1 U22428 ( .A1(n19443), .A2(n19387), .B1(n19383), .B2(n19385), .C1(
        n19422), .C2(n19382), .ZN(P2_U2912) );
  INV_X1 U22429 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19445) );
  INV_X1 U22430 ( .A(n19384), .ZN(n19534) );
  OAI222_X1 U22431 ( .A1(n19445), .A2(n19387), .B1(n19386), .B2(n19385), .C1(
        n19422), .C2(n19534), .ZN(P2_U2913) );
  AOI22_X1 U22432 ( .A1(n19389), .A2(n19388), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19415), .ZN(n19394) );
  OR3_X1 U22433 ( .A1(n19392), .A2(n19391), .A3(n19390), .ZN(n19393) );
  OAI211_X1 U22434 ( .C1(n19395), .C2(n19422), .A(n19394), .B(n19393), .ZN(
        P2_U2914) );
  INV_X1 U22435 ( .A(n20135), .ZN(n19396) );
  AOI22_X1 U22436 ( .A1(n19416), .A2(n19396), .B1(n19415), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19402) );
  OAI21_X1 U22437 ( .B1(n19399), .B2(n19398), .A(n19397), .ZN(n19400) );
  NAND2_X1 U22438 ( .A1(n19400), .A2(n19417), .ZN(n19401) );
  OAI211_X1 U22439 ( .C1(n19403), .C2(n19422), .A(n19402), .B(n19401), .ZN(
        P2_U2916) );
  AOI22_X1 U22440 ( .A1(n19416), .A2(n20147), .B1(n19415), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n19409) );
  OAI21_X1 U22441 ( .B1(n19406), .B2(n19405), .A(n19404), .ZN(n19407) );
  NAND2_X1 U22442 ( .A1(n19407), .A2(n19417), .ZN(n19408) );
  OAI211_X1 U22443 ( .C1(n19518), .C2(n19422), .A(n19409), .B(n19408), .ZN(
        P2_U2917) );
  AOI22_X1 U22444 ( .A1(n19416), .A2(n20157), .B1(n19415), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19414) );
  OAI21_X1 U22445 ( .B1(n19411), .B2(n19418), .A(n19410), .ZN(n19412) );
  NAND2_X1 U22446 ( .A1(n19412), .A2(n19417), .ZN(n19413) );
  OAI211_X1 U22447 ( .C1(n19515), .C2(n19422), .A(n19414), .B(n19413), .ZN(
        P2_U2918) );
  AOI22_X1 U22448 ( .A1(n19416), .A2(n19419), .B1(n19415), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19421) );
  OAI211_X1 U22449 ( .C1(n19548), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        n19420) );
  OAI211_X1 U22450 ( .C1(n19508), .C2(n19422), .A(n19421), .B(n19420), .ZN(
        P2_U2919) );
  NOR2_X1 U22451 ( .A1(n19424), .A2(n19423), .ZN(P2_U2920) );
  INV_X1 U22452 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n20884) );
  INV_X1 U22453 ( .A(n19425), .ZN(n19426) );
  AOI22_X1 U22454 ( .A1(n19459), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(n19426), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n19427) );
  OAI21_X1 U22455 ( .B1(n20884), .B2(n19428), .A(n19427), .ZN(P2_U2928) );
  AOI22_X1 U22456 ( .A1(n19454), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19429) );
  OAI21_X1 U22457 ( .B1(n19430), .B2(n19456), .A(n19429), .ZN(P2_U2936) );
  AOI22_X1 U22458 ( .A1(n19454), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19431) );
  OAI21_X1 U22459 ( .B1(n19432), .B2(n19456), .A(n19431), .ZN(P2_U2937) );
  AOI222_X1 U22460 ( .A1(n19459), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n19458), 
        .B2(P2_EAX_REG_13__SCAN_IN), .C1(n19454), .C2(P2_LWORD_REG_13__SCAN_IN), .ZN(n19433) );
  INV_X1 U22461 ( .A(n19433), .ZN(P2_U2938) );
  AOI222_X1 U22462 ( .A1(n19459), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n19458), 
        .B2(P2_EAX_REG_12__SCAN_IN), .C1(n19454), .C2(P2_LWORD_REG_12__SCAN_IN), .ZN(n19434) );
  INV_X1 U22463 ( .A(n19434), .ZN(P2_U2939) );
  AOI22_X1 U22464 ( .A1(n19454), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19435) );
  OAI21_X1 U22465 ( .B1(n19436), .B2(n19456), .A(n19435), .ZN(P2_U2940) );
  AOI22_X1 U22466 ( .A1(n19454), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19437) );
  OAI21_X1 U22467 ( .B1(n20759), .B2(n19456), .A(n19437), .ZN(P2_U2941) );
  AOI22_X1 U22468 ( .A1(n19454), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19438) );
  OAI21_X1 U22469 ( .B1(n19439), .B2(n19456), .A(n19438), .ZN(P2_U2942) );
  AOI22_X1 U22470 ( .A1(n19454), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19440) );
  OAI21_X1 U22471 ( .B1(n19441), .B2(n19456), .A(n19440), .ZN(P2_U2943) );
  AOI22_X1 U22472 ( .A1(n19454), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19442) );
  OAI21_X1 U22473 ( .B1(n19443), .B2(n19456), .A(n19442), .ZN(P2_U2944) );
  AOI22_X1 U22474 ( .A1(n19454), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19444) );
  OAI21_X1 U22475 ( .B1(n19445), .B2(n19456), .A(n19444), .ZN(P2_U2945) );
  INV_X1 U22476 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19447) );
  AOI22_X1 U22477 ( .A1(n19454), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19446) );
  OAI21_X1 U22478 ( .B1(n19447), .B2(n19456), .A(n19446), .ZN(P2_U2946) );
  AOI22_X1 U22479 ( .A1(n19454), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19448) );
  OAI21_X1 U22480 ( .B1(n19449), .B2(n19456), .A(n19448), .ZN(P2_U2947) );
  INV_X1 U22481 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19451) );
  AOI22_X1 U22482 ( .A1(n19454), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19450) );
  OAI21_X1 U22483 ( .B1(n19451), .B2(n19456), .A(n19450), .ZN(P2_U2948) );
  INV_X1 U22484 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19453) );
  AOI22_X1 U22485 ( .A1(n19454), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19452) );
  OAI21_X1 U22486 ( .B1(n19453), .B2(n19456), .A(n19452), .ZN(P2_U2949) );
  INV_X1 U22487 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19457) );
  AOI22_X1 U22488 ( .A1(n19454), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19459), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19455) );
  OAI21_X1 U22489 ( .B1(n19457), .B2(n19456), .A(n19455), .ZN(P2_U2950) );
  AOI222_X1 U22490 ( .A1(n19459), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(n19458), 
        .B2(P2_EAX_REG_0__SCAN_IN), .C1(n19454), .C2(P2_LWORD_REG_0__SCAN_IN), 
        .ZN(n19460) );
  INV_X1 U22491 ( .A(n19460), .ZN(P2_U2951) );
  AOI22_X1 U22492 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19473), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19461), .ZN(n19469) );
  INV_X1 U22493 ( .A(n19462), .ZN(n19465) );
  OAI22_X1 U22494 ( .A1(n19465), .A2(n16514), .B1(n19464), .B2(n19463), .ZN(
        n19466) );
  AOI21_X1 U22495 ( .B1(n19480), .B2(n19467), .A(n19466), .ZN(n19468) );
  OAI211_X1 U22496 ( .C1(n19471), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U3010) );
  NOR2_X1 U22497 ( .A1(n19473), .A2(n19472), .ZN(n19484) );
  INV_X1 U22498 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19483) );
  NAND2_X1 U22499 ( .A1(n19475), .A2(n19474), .ZN(n19477) );
  OAI211_X1 U22500 ( .C1(n16514), .C2(n19478), .A(n19477), .B(n19476), .ZN(
        n19479) );
  AOI21_X1 U22501 ( .B1(n19481), .B2(n19480), .A(n19479), .ZN(n19482) );
  OAI21_X1 U22502 ( .B1(n19484), .B2(n19483), .A(n19482), .ZN(P2_U3014) );
  AOI211_X1 U22503 ( .C1(n12964), .C2(n19493), .A(n19486), .B(n19485), .ZN(
        n19497) );
  INV_X1 U22504 ( .A(n20157), .ZN(n19488) );
  OAI22_X1 U22505 ( .A1(n19490), .A2(n19489), .B1(n19488), .B2(n19487), .ZN(
        n19496) );
  OAI22_X1 U22506 ( .A1(n19494), .A2(n19493), .B1(n19492), .B2(n19491), .ZN(
        n19495) );
  NOR3_X1 U22507 ( .A1(n19497), .A2(n19496), .A3(n19495), .ZN(n19499) );
  OAI211_X1 U22508 ( .C1(n19501), .C2(n19500), .A(n19499), .B(n19498), .ZN(
        P2_U3045) );
  AOI22_X1 U22509 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19531), .ZN(n20004) );
  AOI22_X1 U22510 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19531), .ZN(n19920) );
  INV_X1 U22511 ( .A(n19920), .ZN(n20001) );
  INV_X1 U22512 ( .A(n19877), .ZN(n19502) );
  AND2_X1 U22513 ( .A1(n19503), .A2(n19525), .ZN(n19992) );
  NAND2_X1 U22514 ( .A1(n20142), .A2(n20149), .ZN(n19600) );
  OR2_X1 U22515 ( .A1(n19600), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19545) );
  NOR2_X1 U22516 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19545), .ZN(
        n19537) );
  AOI22_X1 U22517 ( .A1(n20001), .A2(n19538), .B1(n19992), .B2(n19537), .ZN(
        n19513) );
  AOI21_X1 U22518 ( .B1(n20050), .B2(n19569), .A(n13249), .ZN(n19504) );
  NOR2_X1 U22519 ( .A1(n19504), .A2(n20129), .ZN(n19509) );
  INV_X1 U22520 ( .A(n20042), .ZN(n19506) );
  AOI21_X1 U22521 ( .B1(n10546), .B2(n19670), .A(n20152), .ZN(n19505) );
  AOI21_X1 U22522 ( .B1(n19509), .B2(n19506), .A(n19505), .ZN(n19507) );
  NOR2_X2 U22523 ( .A1(n19508), .A2(n19913), .ZN(n19993) );
  OAI21_X1 U22524 ( .B1(n20042), .B2(n19537), .A(n19509), .ZN(n19511) );
  OAI21_X1 U22525 ( .B1(n10546), .B2(n19537), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19510) );
  NAND2_X1 U22526 ( .A1(n19511), .A2(n19510), .ZN(n19539) );
  AOI22_X1 U22527 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19540), .B1(
        n19993), .B2(n19539), .ZN(n19512) );
  OAI211_X1 U22528 ( .C1(n20004), .C2(n19569), .A(n19513), .B(n19512), .ZN(
        P2_U3048) );
  INV_X1 U22529 ( .A(n19531), .ZN(n19523) );
  INV_X1 U22530 ( .A(n19532), .ZN(n19524) );
  OAI22_X2 U22531 ( .A1(n13868), .A2(n19523), .B1(n13867), .B2(n19524), .ZN(
        n19970) );
  INV_X1 U22532 ( .A(n19970), .ZN(n20010) );
  AOI22_X1 U22533 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19531), .ZN(n19923) );
  INV_X1 U22534 ( .A(n19923), .ZN(n20007) );
  AOI22_X1 U22535 ( .A1(n20007), .A2(n19538), .B1(n20005), .B2(n19537), .ZN(
        n19517) );
  NOR2_X2 U22536 ( .A1(n19515), .A2(n19913), .ZN(n20006) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19540), .B1(
        n20006), .B2(n19539), .ZN(n19516) );
  OAI211_X1 U22538 ( .C1(n20010), .C2(n19569), .A(n19517), .B(n19516), .ZN(
        P2_U3049) );
  AOI22_X1 U22539 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19531), .ZN(n20016) );
  AOI22_X1 U22540 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19531), .ZN(n19926) );
  INV_X1 U22541 ( .A(n19926), .ZN(n20013) );
  AND2_X1 U22542 ( .A1(n10766), .A2(n19525), .ZN(n20011) );
  AOI22_X1 U22543 ( .A1(n20013), .A2(n19538), .B1(n20011), .B2(n19537), .ZN(
        n19520) );
  NOR2_X2 U22544 ( .A1(n19518), .A2(n19913), .ZN(n20012) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19540), .B1(
        n20012), .B2(n19539), .ZN(n19519) );
  OAI211_X1 U22546 ( .C1(n20016), .C2(n19569), .A(n19520), .B(n19519), .ZN(
        P2_U3050) );
  AOI22_X1 U22547 ( .A1(n20019), .A2(n19538), .B1(n20017), .B2(n19537), .ZN(
        n19522) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19540), .B1(
        n20018), .B2(n19539), .ZN(n19521) );
  OAI211_X1 U22549 ( .C1(n20022), .C2(n19569), .A(n19522), .B(n19521), .ZN(
        P2_U3051) );
  OAI22_X2 U22550 ( .A1(n14094), .A2(n19524), .B1(n14095), .B2(n19523), .ZN(
        n19976) );
  AOI22_X1 U22551 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19531), .ZN(n19932) );
  AND2_X1 U22552 ( .A1(n10287), .A2(n19525), .ZN(n20023) );
  AOI22_X1 U22553 ( .A1(n20025), .A2(n19538), .B1(n20023), .B2(n19537), .ZN(
        n19528) );
  NOR2_X2 U22554 ( .A1(n19526), .A2(n19913), .ZN(n20024) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19540), .B1(
        n20024), .B2(n19539), .ZN(n19527) );
  OAI211_X1 U22556 ( .C1(n20028), .C2(n19569), .A(n19528), .B(n19527), .ZN(
        P2_U3052) );
  AOI22_X1 U22557 ( .A1(n20031), .A2(n19538), .B1(n20029), .B2(n19537), .ZN(
        n19530) );
  AOI22_X1 U22558 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19540), .B1(
        n20030), .B2(n19539), .ZN(n19529) );
  OAI211_X1 U22559 ( .C1(n20034), .C2(n19569), .A(n19530), .B(n19529), .ZN(
        P2_U3053) );
  AOI22_X1 U22560 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19531), .ZN(n20040) );
  AOI22_X1 U22561 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19532), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19531), .ZN(n19938) );
  INV_X1 U22562 ( .A(n19938), .ZN(n20037) );
  NOR2_X2 U22563 ( .A1(n10305), .A2(n19533), .ZN(n20035) );
  AOI22_X1 U22564 ( .A1(n20037), .A2(n19538), .B1(n20035), .B2(n19537), .ZN(
        n19536) );
  NOR2_X2 U22565 ( .A1(n19534), .A2(n19913), .ZN(n20036) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19540), .B1(
        n20036), .B2(n19539), .ZN(n19535) );
  OAI211_X1 U22567 ( .C1(n20040), .C2(n19569), .A(n19536), .B(n19535), .ZN(
        P2_U3054) );
  AOI22_X1 U22568 ( .A1(n20045), .A2(n19538), .B1(n20041), .B2(n19537), .ZN(
        n19542) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19540), .B1(
        n20043), .B2(n19539), .ZN(n19541) );
  OAI211_X1 U22570 ( .C1(n20051), .C2(n19569), .A(n19542), .B(n19541), .ZN(
        P2_U3055) );
  NOR2_X1 U22571 ( .A1(n19819), .A2(n19600), .ZN(n19564) );
  OAI21_X1 U22572 ( .B1(n19543), .B2(n19564), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19544) );
  OAI21_X1 U22573 ( .B1(n19545), .B2(n20129), .A(n19544), .ZN(n19565) );
  AOI22_X1 U22574 ( .A1(n19565), .A2(n19993), .B1(n19992), .B2(n19564), .ZN(
        n19551) );
  AOI21_X1 U22575 ( .B1(n10543), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19547) );
  AND2_X1 U22576 ( .A1(n19549), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19762) );
  INV_X1 U22577 ( .A(n19762), .ZN(n19599) );
  OAI21_X1 U22578 ( .B1(n19599), .B2(n19820), .A(n19545), .ZN(n19546) );
  OAI211_X1 U22579 ( .C1(n19564), .C2(n19547), .A(n19546), .B(n19999), .ZN(
        n19566) );
  AOI22_X1 U22580 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19967), .ZN(n19550) );
  OAI211_X1 U22581 ( .C1(n19920), .C2(n19569), .A(n19551), .B(n19550), .ZN(
        P2_U3056) );
  AOI22_X1 U22582 ( .A1(n19565), .A2(n20006), .B1(n20005), .B2(n19564), .ZN(
        n19553) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19970), .ZN(n19552) );
  OAI211_X1 U22584 ( .C1(n19923), .C2(n19569), .A(n19553), .B(n19552), .ZN(
        P2_U3057) );
  AOI22_X1 U22585 ( .A1(n19565), .A2(n20012), .B1(n20011), .B2(n19564), .ZN(
        n19555) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19973), .ZN(n19554) );
  OAI211_X1 U22587 ( .C1(n19926), .C2(n19569), .A(n19555), .B(n19554), .ZN(
        P2_U3058) );
  AOI22_X1 U22588 ( .A1(n19565), .A2(n20018), .B1(n20017), .B2(n19564), .ZN(
        n19557) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19955), .ZN(n19556) );
  OAI211_X1 U22590 ( .C1(n19929), .C2(n19569), .A(n19557), .B(n19556), .ZN(
        P2_U3059) );
  AOI22_X1 U22591 ( .A1(n19565), .A2(n20024), .B1(n20023), .B2(n19564), .ZN(
        n19559) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19976), .ZN(n19558) );
  OAI211_X1 U22593 ( .C1(n19932), .C2(n19569), .A(n19559), .B(n19558), .ZN(
        P2_U3060) );
  AOI22_X1 U22594 ( .A1(n19565), .A2(n20030), .B1(n20029), .B2(n19564), .ZN(
        n19561) );
  AOI22_X1 U22595 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19979), .ZN(n19560) );
  OAI211_X1 U22596 ( .C1(n19935), .C2(n19569), .A(n19561), .B(n19560), .ZN(
        P2_U3061) );
  AOI22_X1 U22597 ( .A1(n19565), .A2(n20036), .B1(n20035), .B2(n19564), .ZN(
        n19563) );
  AOI22_X1 U22598 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19983), .ZN(n19562) );
  OAI211_X1 U22599 ( .C1(n19938), .C2(n19569), .A(n19563), .B(n19562), .ZN(
        P2_U3062) );
  AOI22_X1 U22600 ( .A1(n19565), .A2(n20043), .B1(n20041), .B2(n19564), .ZN(
        n19568) );
  AOI22_X1 U22601 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19566), .B1(
        n19574), .B2(n19941), .ZN(n19567) );
  OAI211_X1 U22602 ( .C1(n19946), .C2(n19569), .A(n19568), .B(n19567), .ZN(
        P2_U3063) );
  NOR2_X1 U22603 ( .A1(n19848), .A2(n19600), .ZN(n19593) );
  INV_X1 U22604 ( .A(n19593), .ZN(n19571) );
  AND2_X1 U22605 ( .A1(n19570), .A2(n19571), .ZN(n19572) );
  OR2_X1 U22606 ( .A1(n19850), .A2(n19600), .ZN(n19575) );
  OAI21_X1 U22607 ( .B1(n19572), .B2(n20182), .A(n19575), .ZN(n19594) );
  AOI22_X1 U22608 ( .A1(n19594), .A2(n19993), .B1(n19992), .B2(n19593), .ZN(
        n19580) );
  AOI21_X1 U22609 ( .B1(n19570), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19578) );
  NOR2_X2 U22610 ( .A1(n19700), .A2(n20132), .ZN(n19625) );
  OAI21_X1 U22611 ( .B1(n19574), .B2(n19625), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19576) );
  NAND3_X1 U22612 ( .A1(n19576), .A2(n20152), .A3(n19575), .ZN(n19577) );
  OAI211_X1 U22613 ( .C1(n19593), .C2(n19578), .A(n19577), .B(n19999), .ZN(
        n19595) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19967), .ZN(n19579) );
  OAI211_X1 U22615 ( .C1(n19920), .C2(n19598), .A(n19580), .B(n19579), .ZN(
        P2_U3064) );
  AOI22_X1 U22616 ( .A1(n19594), .A2(n20006), .B1(n20005), .B2(n19593), .ZN(
        n19582) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19970), .ZN(n19581) );
  OAI211_X1 U22618 ( .C1(n19923), .C2(n19598), .A(n19582), .B(n19581), .ZN(
        P2_U3065) );
  AOI22_X1 U22619 ( .A1(n19594), .A2(n20012), .B1(n20011), .B2(n19593), .ZN(
        n19584) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19973), .ZN(n19583) );
  OAI211_X1 U22621 ( .C1(n19926), .C2(n19598), .A(n19584), .B(n19583), .ZN(
        P2_U3066) );
  AOI22_X1 U22622 ( .A1(n19594), .A2(n20018), .B1(n20017), .B2(n19593), .ZN(
        n19586) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19955), .ZN(n19585) );
  OAI211_X1 U22624 ( .C1(n19929), .C2(n19598), .A(n19586), .B(n19585), .ZN(
        P2_U3067) );
  AOI22_X1 U22625 ( .A1(n19594), .A2(n20024), .B1(n20023), .B2(n19593), .ZN(
        n19588) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19976), .ZN(n19587) );
  OAI211_X1 U22627 ( .C1(n19932), .C2(n19598), .A(n19588), .B(n19587), .ZN(
        P2_U3068) );
  AOI22_X1 U22628 ( .A1(n19594), .A2(n20030), .B1(n20029), .B2(n19593), .ZN(
        n19590) );
  AOI22_X1 U22629 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19979), .ZN(n19589) );
  OAI211_X1 U22630 ( .C1(n19935), .C2(n19598), .A(n19590), .B(n19589), .ZN(
        P2_U3069) );
  AOI22_X1 U22631 ( .A1(n19594), .A2(n20036), .B1(n20035), .B2(n19593), .ZN(
        n19592) );
  AOI22_X1 U22632 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19983), .ZN(n19591) );
  OAI211_X1 U22633 ( .C1(n19938), .C2(n19598), .A(n19592), .B(n19591), .ZN(
        P2_U3070) );
  AOI22_X1 U22634 ( .A1(n19594), .A2(n20043), .B1(n20041), .B2(n19593), .ZN(
        n19597) );
  AOI22_X1 U22635 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19595), .B1(
        n19625), .B2(n19941), .ZN(n19596) );
  OAI211_X1 U22636 ( .C1(n19946), .C2(n19598), .A(n19597), .B(n19596), .ZN(
        P2_U3071) );
  INV_X1 U22637 ( .A(n19625), .ZN(n19619) );
  NOR2_X1 U22638 ( .A1(n19879), .A2(n19600), .ZN(n19624) );
  AOI22_X1 U22639 ( .A1(n19967), .A2(n19635), .B1(n19624), .B2(n19992), .ZN(
        n19610) );
  OAI21_X1 U22640 ( .B1(n19599), .B2(n20132), .A(n20152), .ZN(n19608) );
  NOR2_X1 U22641 ( .A1(n20159), .A2(n19600), .ZN(n19604) );
  INV_X1 U22642 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19670) );
  OAI21_X1 U22643 ( .B1(n19605), .B2(n20182), .A(n19670), .ZN(n19602) );
  INV_X1 U22644 ( .A(n19624), .ZN(n19601) );
  AOI21_X1 U22645 ( .B1(n19602), .B2(n19601), .A(n19913), .ZN(n19603) );
  OAI21_X1 U22646 ( .B1(n19608), .B2(n19604), .A(n19603), .ZN(n19627) );
  INV_X1 U22647 ( .A(n19604), .ZN(n19607) );
  OAI21_X1 U22648 ( .B1(n19605), .B2(n19624), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19606) );
  OAI21_X1 U22649 ( .B1(n19608), .B2(n19607), .A(n19606), .ZN(n19626) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19627), .B1(
        n19993), .B2(n19626), .ZN(n19609) );
  OAI211_X1 U22651 ( .C1(n19920), .C2(n19619), .A(n19610), .B(n19609), .ZN(
        P2_U3072) );
  AOI22_X1 U22652 ( .A1(n19970), .A2(n19635), .B1(n19624), .B2(n20005), .ZN(
        n19612) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19627), .B1(
        n20006), .B2(n19626), .ZN(n19611) );
  OAI211_X1 U22654 ( .C1(n19923), .C2(n19619), .A(n19612), .B(n19611), .ZN(
        P2_U3073) );
  AOI22_X1 U22655 ( .A1(n20013), .A2(n19625), .B1(n19624), .B2(n20011), .ZN(
        n19614) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19627), .B1(
        n20012), .B2(n19626), .ZN(n19613) );
  OAI211_X1 U22657 ( .C1(n20016), .C2(n19668), .A(n19614), .B(n19613), .ZN(
        P2_U3074) );
  AOI22_X1 U22658 ( .A1(n19955), .A2(n19635), .B1(n20017), .B2(n19624), .ZN(
        n19616) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19627), .B1(
        n20018), .B2(n19626), .ZN(n19615) );
  OAI211_X1 U22660 ( .C1(n19929), .C2(n19619), .A(n19616), .B(n19615), .ZN(
        P2_U3075) );
  AOI22_X1 U22661 ( .A1(n19976), .A2(n19635), .B1(n19624), .B2(n20023), .ZN(
        n19618) );
  AOI22_X1 U22662 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19627), .B1(
        n20024), .B2(n19626), .ZN(n19617) );
  OAI211_X1 U22663 ( .C1(n19932), .C2(n19619), .A(n19618), .B(n19617), .ZN(
        P2_U3076) );
  AOI22_X1 U22664 ( .A1(n20031), .A2(n19625), .B1(n20029), .B2(n19624), .ZN(
        n19621) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19627), .B1(
        n20030), .B2(n19626), .ZN(n19620) );
  OAI211_X1 U22666 ( .C1(n20034), .C2(n19668), .A(n19621), .B(n19620), .ZN(
        P2_U3077) );
  AOI22_X1 U22667 ( .A1(n20037), .A2(n19625), .B1(n19624), .B2(n20035), .ZN(
        n19623) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19627), .B1(
        n20036), .B2(n19626), .ZN(n19622) );
  OAI211_X1 U22669 ( .C1(n20040), .C2(n19668), .A(n19623), .B(n19622), .ZN(
        P2_U3078) );
  AOI22_X1 U22670 ( .A1(n20045), .A2(n19625), .B1(n20041), .B2(n19624), .ZN(
        n19629) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19627), .B1(
        n20043), .B2(n19626), .ZN(n19628) );
  OAI211_X1 U22672 ( .C1(n20051), .C2(n19668), .A(n19629), .B(n19628), .ZN(
        P2_U3079) );
  NAND3_X1 U22673 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20142), .A3(
        n20159), .ZN(n19676) );
  NOR2_X1 U22674 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19676), .ZN(
        n19641) );
  INV_X1 U22675 ( .A(n19641), .ZN(n19662) );
  NAND2_X1 U22676 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19662), .ZN(n19630) );
  OR2_X1 U22677 ( .A1(n10560), .A2(n19630), .ZN(n19639) );
  NOR2_X1 U22678 ( .A1(n19632), .A2(n19631), .ZN(n19908) );
  NAND2_X1 U22679 ( .A1(n19908), .A2(n20142), .ZN(n19637) );
  AOI21_X1 U22680 ( .B1(n19637), .B2(n20182), .A(n19704), .ZN(n19633) );
  NAND2_X1 U22681 ( .A1(n19639), .A2(n19633), .ZN(n19663) );
  INV_X1 U22682 ( .A(n19993), .ZN(n19708) );
  INV_X1 U22683 ( .A(n19992), .ZN(n19707) );
  OAI22_X1 U22684 ( .A1(n19663), .A2(n19708), .B1(n19707), .B2(n19662), .ZN(
        n19634) );
  INV_X1 U22685 ( .A(n19634), .ZN(n19643) );
  NOR2_X2 U22686 ( .A1(n19700), .A2(n19672), .ZN(n19694) );
  OAI21_X1 U22687 ( .B1(n19635), .B2(n19694), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19636) );
  NAND2_X1 U22688 ( .A1(n19637), .A2(n19636), .ZN(n19638) );
  AND3_X1 U22689 ( .A1(n19639), .A2(n19999), .A3(n19638), .ZN(n19640) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19967), .ZN(n19642) );
  OAI211_X1 U22691 ( .C1(n19920), .C2(n19668), .A(n19643), .B(n19642), .ZN(
        P2_U3080) );
  INV_X1 U22692 ( .A(n20006), .ZN(n19718) );
  INV_X1 U22693 ( .A(n20005), .ZN(n19717) );
  OAI22_X1 U22694 ( .A1(n19663), .A2(n19718), .B1(n19717), .B2(n19662), .ZN(
        n19644) );
  INV_X1 U22695 ( .A(n19644), .ZN(n19646) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19970), .ZN(n19645) );
  OAI211_X1 U22697 ( .C1(n19923), .C2(n19668), .A(n19646), .B(n19645), .ZN(
        P2_U3081) );
  INV_X1 U22698 ( .A(n20012), .ZN(n19723) );
  INV_X1 U22699 ( .A(n20011), .ZN(n19722) );
  OAI22_X1 U22700 ( .A1(n19663), .A2(n19723), .B1(n19722), .B2(n19662), .ZN(
        n19647) );
  INV_X1 U22701 ( .A(n19647), .ZN(n19649) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19973), .ZN(n19648) );
  OAI211_X1 U22703 ( .C1(n19926), .C2(n19668), .A(n19649), .B(n19648), .ZN(
        P2_U3082) );
  INV_X1 U22704 ( .A(n20018), .ZN(n19728) );
  INV_X1 U22705 ( .A(n20017), .ZN(n19727) );
  OAI22_X1 U22706 ( .A1(n19663), .A2(n19728), .B1(n19727), .B2(n19662), .ZN(
        n19650) );
  INV_X1 U22707 ( .A(n19650), .ZN(n19652) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19955), .ZN(n19651) );
  OAI211_X1 U22709 ( .C1(n19929), .C2(n19668), .A(n19652), .B(n19651), .ZN(
        P2_U3083) );
  INV_X1 U22710 ( .A(n20024), .ZN(n19733) );
  INV_X1 U22711 ( .A(n20023), .ZN(n19732) );
  OAI22_X1 U22712 ( .A1(n19663), .A2(n19733), .B1(n19732), .B2(n19662), .ZN(
        n19653) );
  INV_X1 U22713 ( .A(n19653), .ZN(n19655) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19976), .ZN(n19654) );
  OAI211_X1 U22715 ( .C1(n19932), .C2(n19668), .A(n19655), .B(n19654), .ZN(
        P2_U3084) );
  INV_X1 U22716 ( .A(n20030), .ZN(n19738) );
  INV_X1 U22717 ( .A(n20029), .ZN(n19737) );
  OAI22_X1 U22718 ( .A1(n19663), .A2(n19738), .B1(n19737), .B2(n19662), .ZN(
        n19656) );
  INV_X1 U22719 ( .A(n19656), .ZN(n19658) );
  AOI22_X1 U22720 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19979), .ZN(n19657) );
  OAI211_X1 U22721 ( .C1(n19935), .C2(n19668), .A(n19658), .B(n19657), .ZN(
        P2_U3085) );
  INV_X1 U22722 ( .A(n20036), .ZN(n19743) );
  INV_X1 U22723 ( .A(n20035), .ZN(n19742) );
  OAI22_X1 U22724 ( .A1(n19663), .A2(n19743), .B1(n19742), .B2(n19662), .ZN(
        n19659) );
  INV_X1 U22725 ( .A(n19659), .ZN(n19661) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19983), .ZN(n19660) );
  OAI211_X1 U22727 ( .C1(n19938), .C2(n19668), .A(n19661), .B(n19660), .ZN(
        P2_U3086) );
  INV_X1 U22728 ( .A(n20043), .ZN(n19749) );
  INV_X1 U22729 ( .A(n20041), .ZN(n19748) );
  OAI22_X1 U22730 ( .A1(n19663), .A2(n19749), .B1(n19748), .B2(n19662), .ZN(
        n19664) );
  INV_X1 U22731 ( .A(n19664), .ZN(n19667) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19665), .B1(
        n19694), .B2(n19941), .ZN(n19666) );
  OAI211_X1 U22733 ( .C1(n19946), .C2(n19668), .A(n19667), .B(n19666), .ZN(
        P2_U3087) );
  INV_X1 U22734 ( .A(n19672), .ZN(n19669) );
  AOI21_X1 U22735 ( .B1(n19762), .B2(n19669), .A(n20129), .ZN(n19673) );
  INV_X1 U22736 ( .A(n10555), .ZN(n19674) );
  NOR2_X1 U22737 ( .A1(n20166), .A2(n19676), .ZN(n19710) );
  AOI211_X1 U22738 ( .C1(n19674), .C2(n19670), .A(n19710), .B(n20152), .ZN(
        n19671) );
  AOI211_X2 U22739 ( .C1(n19673), .C2(n19676), .A(n19671), .B(n19913), .ZN(
        n19699) );
  INV_X1 U22740 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n20803) );
  NOR2_X2 U22741 ( .A1(n19757), .A2(n19672), .ZN(n19752) );
  AOI22_X1 U22742 ( .A1(n19967), .A2(n19752), .B1(n19992), .B2(n19710), .ZN(
        n19679) );
  INV_X1 U22743 ( .A(n19673), .ZN(n19677) );
  OAI21_X1 U22744 ( .B1(n19674), .B2(n19710), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19675) );
  OAI21_X1 U22745 ( .B1(n19677), .B2(n19676), .A(n19675), .ZN(n19695) );
  AOI22_X1 U22746 ( .A1(n19993), .A2(n19695), .B1(n19694), .B2(n20001), .ZN(
        n19678) );
  OAI211_X1 U22747 ( .C1(n19699), .C2(n20803), .A(n19679), .B(n19678), .ZN(
        P2_U3088) );
  AOI22_X1 U22748 ( .A1(n20007), .A2(n19694), .B1(n20005), .B2(n19710), .ZN(
        n19681) );
  AOI22_X1 U22749 ( .A1(n20006), .A2(n19695), .B1(n19752), .B2(n19970), .ZN(
        n19680) );
  OAI211_X1 U22750 ( .C1(n19699), .C2(n10414), .A(n19681), .B(n19680), .ZN(
        P2_U3089) );
  INV_X1 U22751 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19684) );
  AOI22_X1 U22752 ( .A1(n20013), .A2(n19694), .B1(n19710), .B2(n20011), .ZN(
        n19683) );
  AOI22_X1 U22753 ( .A1(n20012), .A2(n19695), .B1(n19752), .B2(n19973), .ZN(
        n19682) );
  OAI211_X1 U22754 ( .C1(n19699), .C2(n19684), .A(n19683), .B(n19682), .ZN(
        P2_U3090) );
  AOI22_X1 U22755 ( .A1(n19955), .A2(n19752), .B1(n20017), .B2(n19710), .ZN(
        n19686) );
  AOI22_X1 U22756 ( .A1(n20018), .A2(n19695), .B1(n19694), .B2(n20019), .ZN(
        n19685) );
  OAI211_X1 U22757 ( .C1(n19699), .C2(n10361), .A(n19686), .B(n19685), .ZN(
        P2_U3091) );
  INV_X1 U22758 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19689) );
  AOI22_X1 U22759 ( .A1(n20025), .A2(n19694), .B1(n20023), .B2(n19710), .ZN(
        n19688) );
  AOI22_X1 U22760 ( .A1(n20024), .A2(n19695), .B1(n19752), .B2(n19976), .ZN(
        n19687) );
  OAI211_X1 U22761 ( .C1(n19699), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P2_U3092) );
  AOI22_X1 U22762 ( .A1(n20031), .A2(n19694), .B1(n20029), .B2(n19710), .ZN(
        n19691) );
  AOI22_X1 U22763 ( .A1(n20030), .A2(n19695), .B1(n19752), .B2(n19979), .ZN(
        n19690) );
  OAI211_X1 U22764 ( .C1(n19699), .C2(n10556), .A(n19691), .B(n19690), .ZN(
        P2_U3093) );
  AOI22_X1 U22765 ( .A1(n20037), .A2(n19694), .B1(n19710), .B2(n20035), .ZN(
        n19693) );
  AOI22_X1 U22766 ( .A1(n20036), .A2(n19695), .B1(n19752), .B2(n19983), .ZN(
        n19692) );
  OAI211_X1 U22767 ( .C1(n19699), .C2(n10598), .A(n19693), .B(n19692), .ZN(
        P2_U3094) );
  INV_X1 U22768 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n19698) );
  AOI22_X1 U22769 ( .A1(n20045), .A2(n19694), .B1(n20041), .B2(n19710), .ZN(
        n19697) );
  AOI22_X1 U22770 ( .A1(n20043), .A2(n19695), .B1(n19752), .B2(n19941), .ZN(
        n19696) );
  OAI211_X1 U22771 ( .C1(n19699), .C2(n19698), .A(n19697), .B(n19696), .ZN(
        P2_U3095) );
  NOR2_X1 U22772 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19989), .ZN(
        n19766) );
  INV_X1 U22773 ( .A(n19766), .ZN(n19761) );
  NOR2_X1 U22774 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19761), .ZN(
        n19703) );
  INV_X1 U22775 ( .A(n19703), .ZN(n19747) );
  NAND2_X1 U22776 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19747), .ZN(n19701) );
  OR2_X1 U22777 ( .A1(n19702), .A2(n19701), .ZN(n19713) );
  NOR2_X1 U22778 ( .A1(n19710), .A2(n19703), .ZN(n19705) );
  AOI21_X1 U22779 ( .B1(n20182), .B2(n19705), .A(n19704), .ZN(n19706) );
  NAND2_X1 U22780 ( .A1(n19713), .A2(n19706), .ZN(n19750) );
  OAI22_X1 U22781 ( .A1(n19750), .A2(n19708), .B1(n19707), .B2(n19747), .ZN(
        n19709) );
  INV_X1 U22782 ( .A(n19709), .ZN(n19716) );
  INV_X1 U22783 ( .A(n19710), .ZN(n19712) );
  OAI21_X1 U22784 ( .B1(n19752), .B2(n19783), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19711) );
  OAI221_X1 U22785 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19712), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19711), .A(n19747), .ZN(n19714) );
  NAND3_X1 U22786 ( .A1(n19714), .A2(n19999), .A3(n19713), .ZN(n19753) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20001), .ZN(n19715) );
  OAI211_X1 U22788 ( .C1(n20004), .C2(n19756), .A(n19716), .B(n19715), .ZN(
        P2_U3096) );
  OAI22_X1 U22789 ( .A1(n19750), .A2(n19718), .B1(n19717), .B2(n19747), .ZN(
        n19719) );
  INV_X1 U22790 ( .A(n19719), .ZN(n19721) );
  AOI22_X1 U22791 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20007), .ZN(n19720) );
  OAI211_X1 U22792 ( .C1(n20010), .C2(n19756), .A(n19721), .B(n19720), .ZN(
        P2_U3097) );
  OAI22_X1 U22793 ( .A1(n19750), .A2(n19723), .B1(n19722), .B2(n19747), .ZN(
        n19724) );
  INV_X1 U22794 ( .A(n19724), .ZN(n19726) );
  AOI22_X1 U22795 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20013), .ZN(n19725) );
  OAI211_X1 U22796 ( .C1(n20016), .C2(n19756), .A(n19726), .B(n19725), .ZN(
        P2_U3098) );
  OAI22_X1 U22797 ( .A1(n19750), .A2(n19728), .B1(n19727), .B2(n19747), .ZN(
        n19729) );
  INV_X1 U22798 ( .A(n19729), .ZN(n19731) );
  AOI22_X1 U22799 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20019), .ZN(n19730) );
  OAI211_X1 U22800 ( .C1(n20022), .C2(n19756), .A(n19731), .B(n19730), .ZN(
        P2_U3099) );
  OAI22_X1 U22801 ( .A1(n19750), .A2(n19733), .B1(n19732), .B2(n19747), .ZN(
        n19734) );
  INV_X1 U22802 ( .A(n19734), .ZN(n19736) );
  AOI22_X1 U22803 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20025), .ZN(n19735) );
  OAI211_X1 U22804 ( .C1(n20028), .C2(n19756), .A(n19736), .B(n19735), .ZN(
        P2_U3100) );
  OAI22_X1 U22805 ( .A1(n19750), .A2(n19738), .B1(n19737), .B2(n19747), .ZN(
        n19739) );
  INV_X1 U22806 ( .A(n19739), .ZN(n19741) );
  AOI22_X1 U22807 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20031), .ZN(n19740) );
  OAI211_X1 U22808 ( .C1(n20034), .C2(n19756), .A(n19741), .B(n19740), .ZN(
        P2_U3101) );
  OAI22_X1 U22809 ( .A1(n19750), .A2(n19743), .B1(n19742), .B2(n19747), .ZN(
        n19744) );
  INV_X1 U22810 ( .A(n19744), .ZN(n19746) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20037), .ZN(n19745) );
  OAI211_X1 U22812 ( .C1(n20040), .C2(n19756), .A(n19746), .B(n19745), .ZN(
        P2_U3102) );
  OAI22_X1 U22813 ( .A1(n19750), .A2(n19749), .B1(n19748), .B2(n19747), .ZN(
        n19751) );
  INV_X1 U22814 ( .A(n19751), .ZN(n19755) );
  AOI22_X1 U22815 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19753), .B1(
        n19752), .B2(n20045), .ZN(n19754) );
  OAI211_X1 U22816 ( .C1(n20051), .C2(n19756), .A(n19755), .B(n19754), .ZN(
        P2_U3103) );
  INV_X1 U22817 ( .A(n19764), .ZN(n19759) );
  NOR2_X1 U22818 ( .A1(n20166), .A2(n19761), .ZN(n19792) );
  OAI21_X1 U22819 ( .B1(n19759), .B2(n19792), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19760) );
  OAI21_X1 U22820 ( .B1(n19761), .B2(n20129), .A(n19760), .ZN(n19782) );
  AOI22_X1 U22821 ( .A1(n19782), .A2(n19993), .B1(n19992), .B2(n19792), .ZN(
        n19769) );
  NAND2_X1 U22822 ( .A1(n19762), .A2(n19994), .ZN(n20130) );
  INV_X1 U22823 ( .A(n20130), .ZN(n19767) );
  INV_X1 U22824 ( .A(n19792), .ZN(n19763) );
  OAI211_X1 U22825 ( .C1(n19764), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19763), 
        .B(n20129), .ZN(n19765) );
  OAI211_X1 U22826 ( .C1(n19767), .C2(n19766), .A(n19999), .B(n19765), .ZN(
        n19784) );
  AOI22_X1 U22827 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20001), .ZN(n19768) );
  OAI211_X1 U22828 ( .C1(n20004), .C2(n19818), .A(n19769), .B(n19768), .ZN(
        P2_U3104) );
  AOI22_X1 U22829 ( .A1(n19782), .A2(n20006), .B1(n20005), .B2(n19792), .ZN(
        n19771) );
  AOI22_X1 U22830 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20007), .ZN(n19770) );
  OAI211_X1 U22831 ( .C1(n20010), .C2(n19818), .A(n19771), .B(n19770), .ZN(
        P2_U3105) );
  AOI22_X1 U22832 ( .A1(n19782), .A2(n20012), .B1(n20011), .B2(n19792), .ZN(
        n19773) );
  AOI22_X1 U22833 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20013), .ZN(n19772) );
  OAI211_X1 U22834 ( .C1(n20016), .C2(n19818), .A(n19773), .B(n19772), .ZN(
        P2_U3106) );
  AOI22_X1 U22835 ( .A1(n19782), .A2(n20018), .B1(n20017), .B2(n19792), .ZN(
        n19775) );
  AOI22_X1 U22836 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20019), .ZN(n19774) );
  OAI211_X1 U22837 ( .C1(n20022), .C2(n19818), .A(n19775), .B(n19774), .ZN(
        P2_U3107) );
  AOI22_X1 U22838 ( .A1(n19782), .A2(n20024), .B1(n20023), .B2(n19792), .ZN(
        n19777) );
  AOI22_X1 U22839 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20025), .ZN(n19776) );
  OAI211_X1 U22840 ( .C1(n20028), .C2(n19818), .A(n19777), .B(n19776), .ZN(
        P2_U3108) );
  AOI22_X1 U22841 ( .A1(n19782), .A2(n20030), .B1(n20029), .B2(n19792), .ZN(
        n19779) );
  AOI22_X1 U22842 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20031), .ZN(n19778) );
  OAI211_X1 U22843 ( .C1(n20034), .C2(n19818), .A(n19779), .B(n19778), .ZN(
        P2_U3109) );
  AOI22_X1 U22844 ( .A1(n19782), .A2(n20036), .B1(n20035), .B2(n19792), .ZN(
        n19781) );
  AOI22_X1 U22845 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20037), .ZN(n19780) );
  OAI211_X1 U22846 ( .C1(n20040), .C2(n19818), .A(n19781), .B(n19780), .ZN(
        P2_U3110) );
  AOI22_X1 U22847 ( .A1(n19782), .A2(n20043), .B1(n20041), .B2(n19792), .ZN(
        n19786) );
  AOI22_X1 U22848 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19784), .B1(
        n19783), .B2(n20045), .ZN(n19785) );
  OAI211_X1 U22849 ( .C1(n20051), .C2(n19818), .A(n19786), .B(n19785), .ZN(
        P2_U3111) );
  INV_X1 U22850 ( .A(n19851), .ZN(n19788) );
  INV_X1 U22851 ( .A(n19820), .ZN(n19787) );
  NAND2_X1 U22852 ( .A1(n20149), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19878) );
  NOR2_X1 U22853 ( .A1(n19878), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19823) );
  INV_X1 U22854 ( .A(n19823), .ZN(n19826) );
  NOR2_X1 U22855 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19826), .ZN(
        n19813) );
  AOI22_X1 U22856 ( .A1(n19967), .A2(n19838), .B1(n19992), .B2(n19813), .ZN(
        n19800) );
  INV_X1 U22857 ( .A(n10547), .ZN(n19789) );
  AOI21_X1 U22858 ( .B1(n19789), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19795) );
  INV_X1 U22859 ( .A(n19818), .ZN(n19790) );
  NOR2_X1 U22860 ( .A1(n19838), .A2(n19790), .ZN(n19791) );
  OAI21_X1 U22861 ( .B1(n19791), .B2(n13249), .A(n20152), .ZN(n19798) );
  INV_X1 U22862 ( .A(n19798), .ZN(n19793) );
  NOR2_X1 U22863 ( .A1(n19813), .A2(n19792), .ZN(n19796) );
  NAND2_X1 U22864 ( .A1(n19793), .A2(n19796), .ZN(n19794) );
  OAI211_X1 U22865 ( .C1(n19813), .C2(n19795), .A(n19794), .B(n19999), .ZN(
        n19815) );
  OAI21_X1 U22866 ( .B1(n10547), .B2(n19813), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19797) );
  AOI22_X1 U22867 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19815), .B1(
        n19993), .B2(n19814), .ZN(n19799) );
  OAI211_X1 U22868 ( .C1(n19920), .C2(n19818), .A(n19800), .B(n19799), .ZN(
        P2_U3112) );
  AOI22_X1 U22869 ( .A1(n19970), .A2(n19838), .B1(n20005), .B2(n19813), .ZN(
        n19802) );
  AOI22_X1 U22870 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19815), .B1(
        n20006), .B2(n19814), .ZN(n19801) );
  OAI211_X1 U22871 ( .C1(n19923), .C2(n19818), .A(n19802), .B(n19801), .ZN(
        P2_U3113) );
  AOI22_X1 U22872 ( .A1(n19973), .A2(n19838), .B1(n20011), .B2(n19813), .ZN(
        n19804) );
  AOI22_X1 U22873 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19815), .B1(
        n20012), .B2(n19814), .ZN(n19803) );
  OAI211_X1 U22874 ( .C1(n19926), .C2(n19818), .A(n19804), .B(n19803), .ZN(
        P2_U3114) );
  AOI22_X1 U22875 ( .A1(n19955), .A2(n19838), .B1(n20017), .B2(n19813), .ZN(
        n19806) );
  AOI22_X1 U22876 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19815), .B1(
        n20018), .B2(n19814), .ZN(n19805) );
  OAI211_X1 U22877 ( .C1(n19929), .C2(n19818), .A(n19806), .B(n19805), .ZN(
        P2_U3115) );
  AOI22_X1 U22878 ( .A1(n19976), .A2(n19838), .B1(n20023), .B2(n19813), .ZN(
        n19808) );
  AOI22_X1 U22879 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19815), .B1(
        n20024), .B2(n19814), .ZN(n19807) );
  OAI211_X1 U22880 ( .C1(n19932), .C2(n19818), .A(n19808), .B(n19807), .ZN(
        P2_U3116) );
  AOI22_X1 U22881 ( .A1(n19979), .A2(n19838), .B1(n20029), .B2(n19813), .ZN(
        n19810) );
  AOI22_X1 U22882 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19815), .B1(
        n20030), .B2(n19814), .ZN(n19809) );
  OAI211_X1 U22883 ( .C1(n19935), .C2(n19818), .A(n19810), .B(n19809), .ZN(
        P2_U3117) );
  AOI22_X1 U22884 ( .A1(n19983), .A2(n19838), .B1(n20035), .B2(n19813), .ZN(
        n19812) );
  AOI22_X1 U22885 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19815), .B1(
        n20036), .B2(n19814), .ZN(n19811) );
  OAI211_X1 U22886 ( .C1(n19938), .C2(n19818), .A(n19812), .B(n19811), .ZN(
        P2_U3118) );
  AOI22_X1 U22887 ( .A1(n19941), .A2(n19838), .B1(n20041), .B2(n19813), .ZN(
        n19817) );
  AOI22_X1 U22888 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19815), .B1(
        n20043), .B2(n19814), .ZN(n19816) );
  OAI211_X1 U22889 ( .C1(n19946), .C2(n19818), .A(n19817), .B(n19816), .ZN(
        P2_U3119) );
  NOR2_X1 U22890 ( .A1(n19819), .A2(n19878), .ZN(n19852) );
  AOI22_X1 U22891 ( .A1(n19967), .A2(n19853), .B1(n19992), .B2(n19852), .ZN(
        n19829) );
  OAI21_X1 U22892 ( .B1(n19882), .B2(n19820), .A(n20152), .ZN(n19827) );
  INV_X1 U22893 ( .A(n19852), .ZN(n19821) );
  OAI211_X1 U22894 ( .C1(n10554), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19821), 
        .B(n20129), .ZN(n19822) );
  OAI211_X1 U22895 ( .C1(n19827), .C2(n19823), .A(n19999), .B(n19822), .ZN(
        n19844) );
  OAI21_X1 U22896 ( .B1(n19824), .B2(n19852), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19825) );
  OAI21_X1 U22897 ( .B1(n19827), .B2(n19826), .A(n19825), .ZN(n19843) );
  AOI22_X1 U22898 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19844), .B1(
        n19993), .B2(n19843), .ZN(n19828) );
  OAI211_X1 U22899 ( .C1(n19920), .C2(n19847), .A(n19829), .B(n19828), .ZN(
        P2_U3120) );
  AOI22_X1 U22900 ( .A1(n19970), .A2(n19853), .B1(n20005), .B2(n19852), .ZN(
        n19831) );
  AOI22_X1 U22901 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19844), .B1(
        n20006), .B2(n19843), .ZN(n19830) );
  OAI211_X1 U22902 ( .C1(n19923), .C2(n19847), .A(n19831), .B(n19830), .ZN(
        P2_U3121) );
  AOI22_X1 U22903 ( .A1(n19973), .A2(n19853), .B1(n20011), .B2(n19852), .ZN(
        n19833) );
  AOI22_X1 U22904 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19844), .B1(
        n20012), .B2(n19843), .ZN(n19832) );
  OAI211_X1 U22905 ( .C1(n19926), .C2(n19847), .A(n19833), .B(n19832), .ZN(
        P2_U3122) );
  AOI22_X1 U22906 ( .A1(n20019), .A2(n19838), .B1(n20017), .B2(n19852), .ZN(
        n19835) );
  AOI22_X1 U22907 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19844), .B1(
        n20018), .B2(n19843), .ZN(n19834) );
  OAI211_X1 U22908 ( .C1(n20022), .C2(n19876), .A(n19835), .B(n19834), .ZN(
        P2_U3123) );
  AOI22_X1 U22909 ( .A1(n20025), .A2(n19838), .B1(n20023), .B2(n19852), .ZN(
        n19837) );
  AOI22_X1 U22910 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19844), .B1(
        n20024), .B2(n19843), .ZN(n19836) );
  OAI211_X1 U22911 ( .C1(n20028), .C2(n19876), .A(n19837), .B(n19836), .ZN(
        P2_U3124) );
  AOI22_X1 U22912 ( .A1(n20031), .A2(n19838), .B1(n20029), .B2(n19852), .ZN(
        n19840) );
  AOI22_X1 U22913 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19844), .B1(
        n20030), .B2(n19843), .ZN(n19839) );
  OAI211_X1 U22914 ( .C1(n20034), .C2(n19876), .A(n19840), .B(n19839), .ZN(
        P2_U3125) );
  AOI22_X1 U22915 ( .A1(n19983), .A2(n19853), .B1(n20035), .B2(n19852), .ZN(
        n19842) );
  AOI22_X1 U22916 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19844), .B1(
        n20036), .B2(n19843), .ZN(n19841) );
  OAI211_X1 U22917 ( .C1(n19938), .C2(n19847), .A(n19842), .B(n19841), .ZN(
        P2_U3126) );
  AOI22_X1 U22918 ( .A1(n19941), .A2(n19853), .B1(n20041), .B2(n19852), .ZN(
        n19846) );
  AOI22_X1 U22919 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19844), .B1(
        n20043), .B2(n19843), .ZN(n19845) );
  OAI211_X1 U22920 ( .C1(n19946), .C2(n19847), .A(n19846), .B(n19845), .ZN(
        P2_U3127) );
  NOR2_X1 U22921 ( .A1(n19848), .A2(n19878), .ZN(n19871) );
  OAI21_X1 U22922 ( .B1(n10549), .B2(n19871), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19849) );
  OAI21_X1 U22923 ( .B1(n19878), .B2(n19850), .A(n19849), .ZN(n19872) );
  AOI22_X1 U22924 ( .A1(n19872), .A2(n19993), .B1(n19992), .B2(n19871), .ZN(
        n19858) );
  INV_X1 U22925 ( .A(n10549), .ZN(n19855) );
  AOI221_X1 U22926 ( .B1(n19853), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19904), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19852), .ZN(n19854) );
  AOI211_X1 U22927 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19855), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19854), .ZN(n19856) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19967), .ZN(n19857) );
  OAI211_X1 U22929 ( .C1(n19920), .C2(n19876), .A(n19858), .B(n19857), .ZN(
        P2_U3128) );
  AOI22_X1 U22930 ( .A1(n19872), .A2(n20006), .B1(n20005), .B2(n19871), .ZN(
        n19860) );
  AOI22_X1 U22931 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19970), .ZN(n19859) );
  OAI211_X1 U22932 ( .C1(n19923), .C2(n19876), .A(n19860), .B(n19859), .ZN(
        P2_U3129) );
  AOI22_X1 U22933 ( .A1(n19872), .A2(n20012), .B1(n20011), .B2(n19871), .ZN(
        n19862) );
  AOI22_X1 U22934 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19973), .ZN(n19861) );
  OAI211_X1 U22935 ( .C1(n19926), .C2(n19876), .A(n19862), .B(n19861), .ZN(
        P2_U3130) );
  AOI22_X1 U22936 ( .A1(n19872), .A2(n20018), .B1(n20017), .B2(n19871), .ZN(
        n19864) );
  AOI22_X1 U22937 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19955), .ZN(n19863) );
  OAI211_X1 U22938 ( .C1(n19929), .C2(n19876), .A(n19864), .B(n19863), .ZN(
        P2_U3131) );
  AOI22_X1 U22939 ( .A1(n19872), .A2(n20024), .B1(n20023), .B2(n19871), .ZN(
        n19866) );
  AOI22_X1 U22940 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19976), .ZN(n19865) );
  OAI211_X1 U22941 ( .C1(n19932), .C2(n19876), .A(n19866), .B(n19865), .ZN(
        P2_U3132) );
  AOI22_X1 U22942 ( .A1(n19872), .A2(n20030), .B1(n20029), .B2(n19871), .ZN(
        n19868) );
  AOI22_X1 U22943 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19979), .ZN(n19867) );
  OAI211_X1 U22944 ( .C1(n19935), .C2(n19876), .A(n19868), .B(n19867), .ZN(
        P2_U3133) );
  AOI22_X1 U22945 ( .A1(n19872), .A2(n20036), .B1(n20035), .B2(n19871), .ZN(
        n19870) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19983), .ZN(n19869) );
  OAI211_X1 U22947 ( .C1(n19938), .C2(n19876), .A(n19870), .B(n19869), .ZN(
        P2_U3134) );
  AOI22_X1 U22948 ( .A1(n19872), .A2(n20043), .B1(n20041), .B2(n19871), .ZN(
        n19875) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19873), .B1(
        n19904), .B2(n19941), .ZN(n19874) );
  OAI211_X1 U22950 ( .C1(n19946), .C2(n19876), .A(n19875), .B(n19874), .ZN(
        P2_U3135) );
  OR2_X1 U22951 ( .A1(n20159), .A2(n19878), .ZN(n19885) );
  OR2_X1 U22952 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19885), .ZN(n19881) );
  NOR2_X1 U22953 ( .A1(n19879), .A2(n19878), .ZN(n19902) );
  NOR3_X1 U22954 ( .A1(n19880), .A2(n19902), .A3(n20182), .ZN(n19884) );
  AOI21_X1 U22955 ( .B1(n20182), .B2(n19881), .A(n19884), .ZN(n19903) );
  AOI22_X1 U22956 ( .A1(n19903), .A2(n19993), .B1(n19992), .B2(n19902), .ZN(
        n19889) );
  INV_X1 U22957 ( .A(n19882), .ZN(n19995) );
  INV_X1 U22958 ( .A(n20132), .ZN(n19883) );
  NAND2_X1 U22959 ( .A1(n19995), .A2(n19883), .ZN(n19886) );
  AOI21_X1 U22960 ( .B1(n19886), .B2(n19885), .A(n19884), .ZN(n19887) );
  OAI211_X1 U22961 ( .C1(n19902), .C2(n19670), .A(n19887), .B(n19999), .ZN(
        n19905) );
  AOI22_X1 U22962 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20001), .ZN(n19888) );
  OAI211_X1 U22963 ( .C1(n20004), .C2(n19945), .A(n19889), .B(n19888), .ZN(
        P2_U3136) );
  AOI22_X1 U22964 ( .A1(n19903), .A2(n20006), .B1(n20005), .B2(n19902), .ZN(
        n19891) );
  AOI22_X1 U22965 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20007), .ZN(n19890) );
  OAI211_X1 U22966 ( .C1(n20010), .C2(n19945), .A(n19891), .B(n19890), .ZN(
        P2_U3137) );
  AOI22_X1 U22967 ( .A1(n19903), .A2(n20012), .B1(n20011), .B2(n19902), .ZN(
        n19893) );
  AOI22_X1 U22968 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20013), .ZN(n19892) );
  OAI211_X1 U22969 ( .C1(n20016), .C2(n19945), .A(n19893), .B(n19892), .ZN(
        P2_U3138) );
  AOI22_X1 U22970 ( .A1(n19903), .A2(n20018), .B1(n20017), .B2(n19902), .ZN(
        n19895) );
  AOI22_X1 U22971 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20019), .ZN(n19894) );
  OAI211_X1 U22972 ( .C1(n20022), .C2(n19945), .A(n19895), .B(n19894), .ZN(
        P2_U3139) );
  AOI22_X1 U22973 ( .A1(n19903), .A2(n20024), .B1(n20023), .B2(n19902), .ZN(
        n19897) );
  AOI22_X1 U22974 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20025), .ZN(n19896) );
  OAI211_X1 U22975 ( .C1(n20028), .C2(n19945), .A(n19897), .B(n19896), .ZN(
        P2_U3140) );
  AOI22_X1 U22976 ( .A1(n19903), .A2(n20030), .B1(n20029), .B2(n19902), .ZN(
        n19899) );
  AOI22_X1 U22977 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20031), .ZN(n19898) );
  OAI211_X1 U22978 ( .C1(n20034), .C2(n19945), .A(n19899), .B(n19898), .ZN(
        P2_U3141) );
  AOI22_X1 U22979 ( .A1(n19903), .A2(n20036), .B1(n20035), .B2(n19902), .ZN(
        n19901) );
  AOI22_X1 U22980 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20037), .ZN(n19900) );
  OAI211_X1 U22981 ( .C1(n20040), .C2(n19945), .A(n19901), .B(n19900), .ZN(
        P2_U3142) );
  AOI22_X1 U22982 ( .A1(n19903), .A2(n20043), .B1(n20041), .B2(n19902), .ZN(
        n19907) );
  AOI22_X1 U22983 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19905), .B1(
        n19904), .B2(n20045), .ZN(n19906) );
  OAI211_X1 U22984 ( .C1(n20051), .C2(n19945), .A(n19907), .B(n19906), .ZN(
        P2_U3143) );
  NAND2_X1 U22985 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19908), .ZN(
        n19915) );
  OR2_X1 U22986 ( .A1(n19915), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19911) );
  NOR2_X1 U22987 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19909), .ZN(
        n19939) );
  NOR3_X1 U22988 ( .A1(n19910), .A2(n19939), .A3(n20182), .ZN(n19914) );
  AOI21_X1 U22989 ( .B1(n20182), .B2(n19911), .A(n19914), .ZN(n19940) );
  AOI22_X1 U22990 ( .A1(n19940), .A2(n19993), .B1(n19992), .B2(n19939), .ZN(
        n19919) );
  OAI21_X1 U22991 ( .B1(n19912), .B2(n19963), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19916) );
  AOI211_X1 U22992 ( .C1(n19916), .C2(n19915), .A(n19914), .B(n19913), .ZN(
        n19917) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19967), .ZN(n19918) );
  OAI211_X1 U22994 ( .C1(n19920), .C2(n19945), .A(n19919), .B(n19918), .ZN(
        P2_U3144) );
  AOI22_X1 U22995 ( .A1(n19940), .A2(n20006), .B1(n20005), .B2(n19939), .ZN(
        n19922) );
  AOI22_X1 U22996 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19970), .ZN(n19921) );
  OAI211_X1 U22997 ( .C1(n19923), .C2(n19945), .A(n19922), .B(n19921), .ZN(
        P2_U3145) );
  AOI22_X1 U22998 ( .A1(n19940), .A2(n20012), .B1(n20011), .B2(n19939), .ZN(
        n19925) );
  AOI22_X1 U22999 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19973), .ZN(n19924) );
  OAI211_X1 U23000 ( .C1(n19926), .C2(n19945), .A(n19925), .B(n19924), .ZN(
        P2_U3146) );
  AOI22_X1 U23001 ( .A1(n19940), .A2(n20018), .B1(n20017), .B2(n19939), .ZN(
        n19928) );
  AOI22_X1 U23002 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19955), .ZN(n19927) );
  OAI211_X1 U23003 ( .C1(n19929), .C2(n19945), .A(n19928), .B(n19927), .ZN(
        P2_U3147) );
  AOI22_X1 U23004 ( .A1(n19940), .A2(n20024), .B1(n20023), .B2(n19939), .ZN(
        n19931) );
  AOI22_X1 U23005 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19976), .ZN(n19930) );
  OAI211_X1 U23006 ( .C1(n19932), .C2(n19945), .A(n19931), .B(n19930), .ZN(
        P2_U3148) );
  AOI22_X1 U23007 ( .A1(n19940), .A2(n20030), .B1(n20029), .B2(n19939), .ZN(
        n19934) );
  AOI22_X1 U23008 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19979), .ZN(n19933) );
  OAI211_X1 U23009 ( .C1(n19935), .C2(n19945), .A(n19934), .B(n19933), .ZN(
        P2_U3149) );
  AOI22_X1 U23010 ( .A1(n19940), .A2(n20036), .B1(n20035), .B2(n19939), .ZN(
        n19937) );
  AOI22_X1 U23011 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19983), .ZN(n19936) );
  OAI211_X1 U23012 ( .C1(n19938), .C2(n19945), .A(n19937), .B(n19936), .ZN(
        P2_U3150) );
  AOI22_X1 U23013 ( .A1(n19940), .A2(n20043), .B1(n20041), .B2(n19939), .ZN(
        n19944) );
  AOI22_X1 U23014 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19942), .B1(
        n19963), .B2(n19941), .ZN(n19943) );
  OAI211_X1 U23015 ( .C1(n19946), .C2(n19945), .A(n19944), .B(n19943), .ZN(
        P2_U3151) );
  INV_X1 U23016 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19949) );
  AOI22_X1 U23017 ( .A1(n19962), .A2(n19993), .B1(n19961), .B2(n19992), .ZN(
        n19948) );
  AOI22_X1 U23018 ( .A1(n19963), .A2(n20001), .B1(n19984), .B2(n19967), .ZN(
        n19947) );
  OAI211_X1 U23019 ( .C1(n19966), .C2(n19949), .A(n19948), .B(n19947), .ZN(
        P2_U3152) );
  AOI22_X1 U23020 ( .A1(n19962), .A2(n20006), .B1(n19961), .B2(n20005), .ZN(
        n19951) );
  AOI22_X1 U23021 ( .A1(n19963), .A2(n20007), .B1(n19984), .B2(n19970), .ZN(
        n19950) );
  OAI211_X1 U23022 ( .C1(n19966), .C2(n20925), .A(n19951), .B(n19950), .ZN(
        P2_U3153) );
  INV_X1 U23023 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n19954) );
  AOI22_X1 U23024 ( .A1(n19962), .A2(n20012), .B1(n19961), .B2(n20011), .ZN(
        n19953) );
  AOI22_X1 U23025 ( .A1(n19963), .A2(n20013), .B1(n19984), .B2(n19973), .ZN(
        n19952) );
  OAI211_X1 U23026 ( .C1(n19966), .C2(n19954), .A(n19953), .B(n19952), .ZN(
        P2_U3154) );
  AOI22_X1 U23027 ( .A1(n19962), .A2(n20018), .B1(n19961), .B2(n20017), .ZN(
        n19957) );
  AOI22_X1 U23028 ( .A1(n19963), .A2(n20019), .B1(n19984), .B2(n19955), .ZN(
        n19956) );
  OAI211_X1 U23029 ( .C1(n19966), .C2(n10375), .A(n19957), .B(n19956), .ZN(
        P2_U3155) );
  INV_X1 U23030 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n19960) );
  AOI22_X1 U23031 ( .A1(n19962), .A2(n20024), .B1(n19961), .B2(n20023), .ZN(
        n19959) );
  AOI22_X1 U23032 ( .A1(n19963), .A2(n20025), .B1(n19984), .B2(n19976), .ZN(
        n19958) );
  OAI211_X1 U23033 ( .C1(n19966), .C2(n19960), .A(n19959), .B(n19958), .ZN(
        P2_U3156) );
  AOI22_X1 U23034 ( .A1(n19962), .A2(n20036), .B1(n19961), .B2(n20035), .ZN(
        n19965) );
  AOI22_X1 U23035 ( .A1(n19963), .A2(n20037), .B1(n19984), .B2(n19983), .ZN(
        n19964) );
  OAI211_X1 U23036 ( .C1(n19966), .C2(n10599), .A(n19965), .B(n19964), .ZN(
        P2_U3158) );
  AOI22_X1 U23037 ( .A1(n20001), .A2(n19984), .B1(n19982), .B2(n19992), .ZN(
        n19969) );
  AOI22_X1 U23038 ( .A1(n19993), .A2(n19985), .B1(n20046), .B2(n19967), .ZN(
        n19968) );
  OAI211_X1 U23039 ( .C1(n19988), .C2(n20807), .A(n19969), .B(n19968), .ZN(
        P2_U3160) );
  AOI22_X1 U23040 ( .A1(n20007), .A2(n19984), .B1(n19982), .B2(n20005), .ZN(
        n19972) );
  AOI22_X1 U23041 ( .A1(n20006), .A2(n19985), .B1(n20046), .B2(n19970), .ZN(
        n19971) );
  OAI211_X1 U23042 ( .C1(n19988), .C2(n14528), .A(n19972), .B(n19971), .ZN(
        P2_U3161) );
  AOI22_X1 U23043 ( .A1(n19973), .A2(n20046), .B1(n19982), .B2(n20011), .ZN(
        n19975) );
  AOI22_X1 U23044 ( .A1(n20012), .A2(n19985), .B1(n19984), .B2(n20013), .ZN(
        n19974) );
  OAI211_X1 U23045 ( .C1(n19988), .C2(n14559), .A(n19975), .B(n19974), .ZN(
        P2_U3162) );
  AOI22_X1 U23046 ( .A1(n20025), .A2(n19984), .B1(n19982), .B2(n20023), .ZN(
        n19978) );
  AOI22_X1 U23047 ( .A1(n20024), .A2(n19985), .B1(n20046), .B2(n19976), .ZN(
        n19977) );
  OAI211_X1 U23048 ( .C1(n19988), .C2(n14612), .A(n19978), .B(n19977), .ZN(
        P2_U3164) );
  AOI22_X1 U23049 ( .A1(n19979), .A2(n20046), .B1(n20029), .B2(n19982), .ZN(
        n19981) );
  AOI22_X1 U23050 ( .A1(n20030), .A2(n19985), .B1(n19984), .B2(n20031), .ZN(
        n19980) );
  OAI211_X1 U23051 ( .C1(n19988), .C2(n14638), .A(n19981), .B(n19980), .ZN(
        P2_U3165) );
  AOI22_X1 U23052 ( .A1(n19983), .A2(n20046), .B1(n19982), .B2(n20035), .ZN(
        n19987) );
  AOI22_X1 U23053 ( .A1(n20036), .A2(n19985), .B1(n19984), .B2(n20037), .ZN(
        n19986) );
  OAI211_X1 U23054 ( .C1(n19988), .C2(n14657), .A(n19987), .B(n19986), .ZN(
        P2_U3166) );
  OR2_X1 U23055 ( .A1(n20142), .A2(n19989), .ZN(n19997) );
  OR2_X1 U23056 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19997), .ZN(n19991) );
  NOR3_X1 U23057 ( .A1(n19990), .A2(n20042), .A3(n20182), .ZN(n19996) );
  AOI21_X1 U23058 ( .B1(n20182), .B2(n19991), .A(n19996), .ZN(n20044) );
  AOI22_X1 U23059 ( .A1(n20044), .A2(n19993), .B1(n20042), .B2(n19992), .ZN(
        n20003) );
  NAND2_X1 U23060 ( .A1(n19995), .A2(n19994), .ZN(n19998) );
  AOI21_X1 U23061 ( .B1(n19998), .B2(n19997), .A(n19996), .ZN(n20000) );
  OAI211_X1 U23062 ( .C1(n20042), .C2(n19670), .A(n20000), .B(n19999), .ZN(
        n20047) );
  AOI22_X1 U23063 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20001), .ZN(n20002) );
  OAI211_X1 U23064 ( .C1(n20004), .C2(n20050), .A(n20003), .B(n20002), .ZN(
        P2_U3168) );
  AOI22_X1 U23065 ( .A1(n20044), .A2(n20006), .B1(n20042), .B2(n20005), .ZN(
        n20009) );
  AOI22_X1 U23066 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20007), .ZN(n20008) );
  OAI211_X1 U23067 ( .C1(n20010), .C2(n20050), .A(n20009), .B(n20008), .ZN(
        P2_U3169) );
  AOI22_X1 U23068 ( .A1(n20044), .A2(n20012), .B1(n20042), .B2(n20011), .ZN(
        n20015) );
  AOI22_X1 U23069 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20013), .ZN(n20014) );
  OAI211_X1 U23070 ( .C1(n20016), .C2(n20050), .A(n20015), .B(n20014), .ZN(
        P2_U3170) );
  AOI22_X1 U23071 ( .A1(n20044), .A2(n20018), .B1(n20042), .B2(n20017), .ZN(
        n20021) );
  AOI22_X1 U23072 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20019), .ZN(n20020) );
  OAI211_X1 U23073 ( .C1(n20022), .C2(n20050), .A(n20021), .B(n20020), .ZN(
        P2_U3171) );
  AOI22_X1 U23074 ( .A1(n20044), .A2(n20024), .B1(n20042), .B2(n20023), .ZN(
        n20027) );
  AOI22_X1 U23075 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20025), .ZN(n20026) );
  OAI211_X1 U23076 ( .C1(n20028), .C2(n20050), .A(n20027), .B(n20026), .ZN(
        P2_U3172) );
  AOI22_X1 U23077 ( .A1(n20044), .A2(n20030), .B1(n20042), .B2(n20029), .ZN(
        n20033) );
  AOI22_X1 U23078 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20031), .ZN(n20032) );
  OAI211_X1 U23079 ( .C1(n20034), .C2(n20050), .A(n20033), .B(n20032), .ZN(
        P2_U3173) );
  AOI22_X1 U23080 ( .A1(n20044), .A2(n20036), .B1(n20042), .B2(n20035), .ZN(
        n20039) );
  AOI22_X1 U23081 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20037), .ZN(n20038) );
  OAI211_X1 U23082 ( .C1(n20040), .C2(n20050), .A(n20039), .B(n20038), .ZN(
        P2_U3174) );
  AOI22_X1 U23083 ( .A1(n20044), .A2(n20043), .B1(n20042), .B2(n20041), .ZN(
        n20049) );
  AOI22_X1 U23084 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20047), .B1(
        n20046), .B2(n20045), .ZN(n20048) );
  OAI211_X1 U23085 ( .C1(n20051), .C2(n20050), .A(n20049), .B(n20048), .ZN(
        P2_U3175) );
  INV_X1 U23086 ( .A(n20055), .ZN(n20053) );
  OAI211_X1 U23087 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n20190), .A(n20053), 
        .B(n20052), .ZN(n20058) );
  OAI211_X1 U23088 ( .C1(n20055), .C2(n20054), .A(n20183), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n20057) );
  OAI211_X1 U23089 ( .C1(n20059), .C2(n20058), .A(n20057), .B(n20056), .ZN(
        P2_U3177) );
  INV_X1 U23090 ( .A(n20128), .ZN(n20060) );
  AND2_X1 U23091 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20060), .ZN(
        P2_U3179) );
  AND2_X1 U23092 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20060), .ZN(
        P2_U3180) );
  AND2_X1 U23093 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20060), .ZN(
        P2_U3181) );
  AND2_X1 U23094 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20060), .ZN(
        P2_U3182) );
  AND2_X1 U23095 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20060), .ZN(
        P2_U3183) );
  AND2_X1 U23096 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20060), .ZN(
        P2_U3184) );
  AND2_X1 U23097 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20060), .ZN(
        P2_U3185) );
  AND2_X1 U23098 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20060), .ZN(
        P2_U3186) );
  AND2_X1 U23099 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20060), .ZN(
        P2_U3187) );
  AND2_X1 U23100 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20060), .ZN(
        P2_U3188) );
  AND2_X1 U23101 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20060), .ZN(
        P2_U3189) );
  AND2_X1 U23102 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20060), .ZN(
        P2_U3190) );
  AND2_X1 U23103 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20060), .ZN(
        P2_U3191) );
  AND2_X1 U23104 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20060), .ZN(
        P2_U3192) );
  AND2_X1 U23105 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20060), .ZN(
        P2_U3193) );
  AND2_X1 U23106 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20060), .ZN(
        P2_U3194) );
  INV_X1 U23107 ( .A(P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20712) );
  NOR2_X1 U23108 ( .A1(n20712), .A2(n20128), .ZN(P2_U3195) );
  AND2_X1 U23109 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20060), .ZN(
        P2_U3196) );
  AND2_X1 U23110 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20060), .ZN(
        P2_U3197) );
  AND2_X1 U23111 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20060), .ZN(
        P2_U3198) );
  NOR2_X1 U23112 ( .A1(n20741), .A2(n20128), .ZN(P2_U3199) );
  AND2_X1 U23113 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20060), .ZN(
        P2_U3200) );
  AND2_X1 U23114 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20060), .ZN(P2_U3201) );
  NOR2_X1 U23115 ( .A1(n20731), .A2(n20128), .ZN(P2_U3202) );
  AND2_X1 U23116 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20060), .ZN(P2_U3203) );
  AND2_X1 U23117 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20060), .ZN(P2_U3204) );
  AND2_X1 U23118 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20060), .ZN(P2_U3205) );
  AND2_X1 U23119 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20060), .ZN(P2_U3206) );
  INV_X1 U23120 ( .A(P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20756) );
  NOR2_X1 U23121 ( .A1(n20756), .A2(n20128), .ZN(P2_U3207) );
  AND2_X1 U23122 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20060), .ZN(P2_U3208) );
  INV_X1 U23123 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20066) );
  NOR2_X1 U23124 ( .A1(n20061), .A2(n20066), .ZN(n20065) );
  NAND2_X1 U23125 ( .A1(n20183), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n20073) );
  AOI21_X1 U23126 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(n20624), .A(n20062), .ZN(n20063) );
  INV_X1 U23127 ( .A(NA), .ZN(n20629) );
  NOR3_X1 U23128 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n20629), .ZN(n20078) );
  AOI21_X1 U23129 ( .B1(n20063), .B2(n20194), .A(n20078), .ZN(n20064) );
  OAI221_X1 U23130 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n20065), .C1(
        P2_STATE_REG_2__SCAN_IN), .C2(n20073), .A(n20064), .ZN(P2_U3209) );
  AOI21_X1 U23131 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20624), .A(n20079), 
        .ZN(n20071) );
  NOR3_X1 U23132 ( .A1(n20071), .A2(n20066), .A3(n20061), .ZN(n20067) );
  INV_X1 U23133 ( .A(n20073), .ZN(n20072) );
  NOR2_X1 U23134 ( .A1(n20067), .A2(n20072), .ZN(n20069) );
  OAI211_X1 U23135 ( .C1(n20624), .C2(n20070), .A(n20069), .B(n20068), .ZN(
        P2_U3210) );
  AOI21_X1 U23136 ( .B1(n20072), .B2(P2_STATE_REG_2__SCAN_IN), .A(n20071), 
        .ZN(n20077) );
  OAI22_X1 U23137 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n20074), .B1(NA), 
        .B2(n20073), .ZN(n20075) );
  OAI211_X1 U23138 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n20075), .ZN(n20076) );
  OAI21_X1 U23139 ( .B1(n20078), .B2(n20077), .A(n20076), .ZN(P2_U3211) );
  INV_X1 U23140 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20082) );
  NAND2_X1 U23141 ( .A1(n20193), .A2(n20079), .ZN(n20121) );
  CLKBUF_X1 U23142 ( .A(n20121), .Z(n20118) );
  OAI222_X1 U23143 ( .A1(n20119), .A2(n10986), .B1(n20080), .B2(n20193), .C1(
        n20082), .C2(n20118), .ZN(P2_U3212) );
  OAI222_X1 U23144 ( .A1(n20119), .A2(n20082), .B1(n20081), .B2(n20193), .C1(
        n11004), .C2(n20118), .ZN(P2_U3213) );
  OAI222_X1 U23145 ( .A1(n20119), .A2(n11004), .B1(n20083), .B2(n20193), .C1(
        n10868), .C2(n20118), .ZN(P2_U3214) );
  OAI222_X1 U23146 ( .A1(n20118), .A2(n13523), .B1(n20084), .B2(n20193), .C1(
        n10868), .C2(n20115), .ZN(P2_U3215) );
  OAI222_X1 U23147 ( .A1(n20121), .A2(n14014), .B1(n20085), .B2(n20193), .C1(
        n13523), .C2(n20115), .ZN(P2_U3216) );
  OAI222_X1 U23148 ( .A1(n20121), .A2(n10858), .B1(n20086), .B2(n20193), .C1(
        n14014), .C2(n20115), .ZN(P2_U3217) );
  OAI222_X1 U23149 ( .A1(n20121), .A2(n11037), .B1(n20087), .B2(n20193), .C1(
        n10858), .C2(n20115), .ZN(P2_U3218) );
  OAI222_X1 U23150 ( .A1(n20121), .A2(n11054), .B1(n20088), .B2(n20193), .C1(
        n11037), .C2(n20115), .ZN(P2_U3219) );
  OAI222_X1 U23151 ( .A1(n20121), .A2(n11067), .B1(n20089), .B2(n20193), .C1(
        n11054), .C2(n20115), .ZN(P2_U3220) );
  OAI222_X1 U23152 ( .A1(n20118), .A2(n11083), .B1(n20090), .B2(n20193), .C1(
        n11067), .C2(n20115), .ZN(P2_U3221) );
  OAI222_X1 U23153 ( .A1(n20118), .A2(n11097), .B1(n20091), .B2(n20193), .C1(
        n11083), .C2(n20115), .ZN(P2_U3222) );
  OAI222_X1 U23154 ( .A1(n20118), .A2(n10891), .B1(n20092), .B2(n20193), .C1(
        n11097), .C2(n20115), .ZN(P2_U3223) );
  OAI222_X1 U23155 ( .A1(n20118), .A2(n11129), .B1(n20093), .B2(n20193), .C1(
        n10891), .C2(n20115), .ZN(P2_U3224) );
  OAI222_X1 U23156 ( .A1(n20118), .A2(n20910), .B1(n20094), .B2(n20193), .C1(
        n11129), .C2(n20115), .ZN(P2_U3225) );
  OAI222_X1 U23157 ( .A1(n20118), .A2(n20808), .B1(n20095), .B2(n20193), .C1(
        n20910), .C2(n20119), .ZN(P2_U3226) );
  OAI222_X1 U23158 ( .A1(n20121), .A2(n20097), .B1(n20096), .B2(n20193), .C1(
        n20808), .C2(n20119), .ZN(P2_U3227) );
  OAI222_X1 U23159 ( .A1(n20121), .A2(n20099), .B1(n20098), .B2(n20193), .C1(
        n20097), .C2(n20119), .ZN(P2_U3228) );
  INV_X1 U23160 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20101) );
  OAI222_X1 U23161 ( .A1(n20121), .A2(n20101), .B1(n20100), .B2(n20193), .C1(
        n20099), .C2(n20115), .ZN(P2_U3229) );
  OAI222_X1 U23162 ( .A1(n20121), .A2(n20103), .B1(n20102), .B2(n20193), .C1(
        n20101), .C2(n20115), .ZN(P2_U3230) );
  OAI222_X1 U23163 ( .A1(n20121), .A2(n15663), .B1(n20104), .B2(n20193), .C1(
        n20103), .C2(n20115), .ZN(P2_U3231) );
  INV_X1 U23164 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n20106) );
  OAI222_X1 U23165 ( .A1(n20121), .A2(n20106), .B1(n20105), .B2(n20193), .C1(
        n15663), .C2(n20115), .ZN(P2_U3232) );
  OAI222_X1 U23166 ( .A1(n20118), .A2(n11157), .B1(n20107), .B2(n20193), .C1(
        n20106), .C2(n20115), .ZN(P2_U3233) );
  OAI222_X1 U23167 ( .A1(n20118), .A2(n20109), .B1(n20108), .B2(n20193), .C1(
        n11157), .C2(n20115), .ZN(P2_U3234) );
  OAI222_X1 U23168 ( .A1(n20118), .A2(n10925), .B1(n20842), .B2(n20193), .C1(
        n20109), .C2(n20115), .ZN(P2_U3235) );
  OAI222_X1 U23169 ( .A1(n20118), .A2(n20111), .B1(n20110), .B2(n20193), .C1(
        n10925), .C2(n20115), .ZN(P2_U3236) );
  OAI222_X1 U23170 ( .A1(n20118), .A2(n15608), .B1(n20112), .B2(n20193), .C1(
        n20111), .C2(n20115), .ZN(P2_U3237) );
  OAI222_X1 U23171 ( .A1(n20119), .A2(n15608), .B1(n20901), .B2(n20193), .C1(
        n20113), .C2(n20118), .ZN(P2_U3238) );
  OAI222_X1 U23172 ( .A1(n20118), .A2(n20116), .B1(n20114), .B2(n20193), .C1(
        n20113), .C2(n20115), .ZN(P2_U3239) );
  OAI222_X1 U23173 ( .A1(n20118), .A2(n20743), .B1(n20117), .B2(n20193), .C1(
        n20116), .C2(n20115), .ZN(P2_U3240) );
  OAI222_X1 U23174 ( .A1(n20121), .A2(n16414), .B1(n20120), .B2(n20193), .C1(
        n20743), .C2(n20119), .ZN(P2_U3241) );
  OAI22_X1 U23175 ( .A1(n20194), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20193), .ZN(n20122) );
  INV_X1 U23176 ( .A(n20122), .ZN(P2_U3585) );
  MUX2_X1 U23177 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20194), .Z(P2_U3586) );
  OAI22_X1 U23178 ( .A1(n20194), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20193), .ZN(n20123) );
  INV_X1 U23179 ( .A(n20123), .ZN(P2_U3587) );
  OAI22_X1 U23180 ( .A1(n20194), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20193), .ZN(n20124) );
  INV_X1 U23181 ( .A(n20124), .ZN(P2_U3588) );
  OAI21_X1 U23182 ( .B1(n20128), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20126), 
        .ZN(n20125) );
  INV_X1 U23183 ( .A(n20125), .ZN(P2_U3591) );
  OAI21_X1 U23184 ( .B1(n20128), .B2(n20127), .A(n20126), .ZN(P2_U3592) );
  OR2_X1 U23185 ( .A1(n20130), .A2(n20129), .ZN(n20140) );
  NAND2_X1 U23186 ( .A1(n20152), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20131) );
  OR2_X1 U23187 ( .A1(n20132), .A2(n20131), .ZN(n20143) );
  NAND2_X1 U23188 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n20133), .ZN(n20134) );
  OAI21_X1 U23189 ( .B1(n20153), .B2(n20134), .A(n20150), .ZN(n20144) );
  NAND2_X1 U23190 ( .A1(n20143), .A2(n20144), .ZN(n20138) );
  NOR2_X1 U23191 ( .A1(n20135), .A2(n19670), .ZN(n20136) );
  AOI21_X1 U23192 ( .B1(n20138), .B2(n20137), .A(n20136), .ZN(n20139) );
  AND2_X1 U23193 ( .A1(n20140), .A2(n20139), .ZN(n20141) );
  AOI22_X1 U23194 ( .A1(n20167), .A2(n20142), .B1(n20141), .B2(n20164), .ZN(
        P2_U3602) );
  OAI21_X1 U23195 ( .B1(n20145), .B2(n20144), .A(n20143), .ZN(n20146) );
  AOI21_X1 U23196 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20147), .A(n20146), 
        .ZN(n20148) );
  AOI22_X1 U23197 ( .A1(n20167), .A2(n20149), .B1(n20148), .B2(n20164), .ZN(
        P2_U3603) );
  INV_X1 U23198 ( .A(n20150), .ZN(n20160) );
  AND2_X1 U23199 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20151) );
  OR3_X1 U23200 ( .A1(n20153), .A2(n20160), .A3(n20151), .ZN(n20155) );
  NAND3_X1 U23201 ( .A1(n20153), .A2(n20152), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n20154) );
  NAND2_X1 U23202 ( .A1(n20155), .A2(n20154), .ZN(n20156) );
  AOI21_X1 U23203 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20157), .A(n20156), 
        .ZN(n20158) );
  AOI22_X1 U23204 ( .A1(n20167), .A2(n20159), .B1(n20158), .B2(n20164), .ZN(
        P2_U3604) );
  OAI22_X1 U23205 ( .A1(n20161), .A2(n20160), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19670), .ZN(n20162) );
  AOI21_X1 U23206 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20163), .A(n20162), 
        .ZN(n20165) );
  AOI22_X1 U23207 ( .A1(n20167), .A2(n20166), .B1(n20165), .B2(n20164), .ZN(
        P2_U3605) );
  INV_X1 U23208 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20168) );
  AOI22_X1 U23209 ( .A1(n20193), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20168), 
        .B2(n20194), .ZN(P2_U3608) );
  INV_X1 U23210 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n20177) );
  AOI22_X1 U23211 ( .A1(n20172), .A2(n20171), .B1(n20170), .B2(n20169), .ZN(
        n20175) );
  NOR2_X1 U23212 ( .A1(n20173), .A2(n20176), .ZN(n20174) );
  AOI22_X1 U23213 ( .A1(n20177), .A2(n20176), .B1(n20175), .B2(n20174), .ZN(
        P2_U3609) );
  OAI21_X1 U23214 ( .B1(n20179), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n20178), 
        .ZN(n20180) );
  NAND3_X1 U23215 ( .A1(n20181), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n20180), 
        .ZN(n20186) );
  OAI22_X1 U23216 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20184), .B1(n20183), 
        .B2(n20182), .ZN(n20185) );
  NAND2_X1 U23217 ( .A1(n20186), .A2(n20185), .ZN(n20192) );
  AOI21_X1 U23218 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20187), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20189) );
  AOI211_X1 U23219 ( .C1(n19454), .C2(n20190), .A(n20189), .B(n20188), .ZN(
        n20191) );
  MUX2_X1 U23220 ( .A(n20192), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n20191), 
        .Z(P2_U3610) );
  OAI22_X1 U23221 ( .A1(n20194), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20193), .ZN(n20195) );
  INV_X1 U23222 ( .A(n20195), .ZN(P2_U3611) );
  AOI21_X1 U23223 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20632), .A(n12770), 
        .ZN(n20625) );
  INV_X1 U23224 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n20196) );
  AOI21_X1 U23225 ( .B1(n20625), .B2(n20196), .A(n20693), .ZN(P1_U2802) );
  OAI21_X1 U23226 ( .B1(n20198), .B2(n20197), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n20199) );
  OAI21_X1 U23227 ( .B1(n20200), .B2(n10118), .A(n20199), .ZN(P1_U2803) );
  NOR2_X1 U23228 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20202) );
  OAI21_X1 U23229 ( .B1(n20202), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20691), .ZN(
        n20201) );
  OAI21_X1 U23230 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20691), .A(n20201), 
        .ZN(P1_U2804) );
  NOR2_X1 U23231 ( .A1(n20625), .A2(n20693), .ZN(n20683) );
  OAI21_X1 U23232 ( .B1(BS16), .B2(n20202), .A(n20683), .ZN(n20681) );
  OAI21_X1 U23233 ( .B1(n20683), .B2(n20818), .A(n20681), .ZN(P1_U2805) );
  OAI21_X1 U23234 ( .B1(n20205), .B2(n20204), .A(n20203), .ZN(P1_U2806) );
  NOR2_X1 U23235 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20975) );
  AOI211_X1 U23236 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_4__SCAN_IN), .B(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20206) );
  INV_X1 U23237 ( .A(P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20619) );
  INV_X1 U23238 ( .A(P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n20863) );
  NAND4_X1 U23239 ( .A1(n20975), .A2(n20206), .A3(n20619), .A4(n20863), .ZN(
        n20214) );
  OR4_X1 U23240 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20213) );
  OR4_X1 U23241 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n20212) );
  NOR4_X1 U23242 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20210) );
  NOR4_X1 U23243 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20209) );
  NOR4_X1 U23244 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n20208) );
  NOR4_X1 U23245 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20207) );
  NAND4_X1 U23246 ( .A1(n20210), .A2(n20209), .A3(n20208), .A4(n20207), .ZN(
        n20211) );
  INV_X1 U23247 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20216) );
  NOR3_X1 U23248 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20217) );
  OAI21_X1 U23249 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20217), .A(n20687), .ZN(
        n20215) );
  OAI21_X1 U23250 ( .B1(n20687), .B2(n20216), .A(n20215), .ZN(P1_U2807) );
  INV_X1 U23251 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20682) );
  AOI21_X1 U23252 ( .B1(n13275), .B2(n20682), .A(n20217), .ZN(n20219) );
  INV_X1 U23253 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20218) );
  INV_X1 U23254 ( .A(n20687), .ZN(n20689) );
  AOI22_X1 U23255 ( .A1(n20687), .A2(n20219), .B1(n20218), .B2(n20689), .ZN(
        P1_U2808) );
  AOI22_X1 U23256 ( .A1(n20263), .A2(P1_EBX_REG_9__SCAN_IN), .B1(n20221), .B2(
        n20220), .ZN(n20222) );
  OAI211_X1 U23257 ( .C1(n20257), .C2(n20969), .A(n20222), .B(n20254), .ZN(
        n20223) );
  AOI21_X1 U23258 ( .B1(n20253), .B2(n20278), .A(n20223), .ZN(n20226) );
  AOI22_X1 U23259 ( .A1(n20279), .A2(n20233), .B1(n14061), .B2(n20224), .ZN(
        n20225) );
  OAI211_X1 U23260 ( .C1(n20227), .C2(n14061), .A(n20226), .B(n20225), .ZN(
        P1_U2831) );
  AOI22_X1 U23261 ( .A1(n20263), .A2(P1_EBX_REG_7__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n20269), .ZN(n20228) );
  OAI211_X1 U23262 ( .C1(n20267), .C2(n20229), .A(n20228), .B(n20254), .ZN(
        n20230) );
  AOI221_X1 U23263 ( .B1(n20239), .B2(P1_REIP_REG_7__SCAN_IN), .C1(n20232), 
        .C2(n20231), .A(n20230), .ZN(n20236) );
  NAND2_X1 U23264 ( .A1(n20234), .A2(n20233), .ZN(n20235) );
  OAI211_X1 U23265 ( .C1(n20277), .C2(n20237), .A(n20236), .B(n20235), .ZN(
        P1_U2833) );
  INV_X1 U23266 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20238) );
  NOR4_X1 U23267 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20249), .A3(n20271), .A4(
        n20238), .ZN(n20245) );
  AOI21_X1 U23268 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20239), .A(n20349), .ZN(
        n20241) );
  AOI22_X1 U23269 ( .A1(n20263), .A2(P1_EBX_REG_6__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20269), .ZN(n20240) );
  OAI211_X1 U23270 ( .C1(n20243), .C2(n20242), .A(n20241), .B(n20240), .ZN(
        n20244) );
  AOI211_X1 U23271 ( .C1(n20246), .C2(n20253), .A(n20245), .B(n20244), .ZN(
        n20247) );
  OAI21_X1 U23272 ( .B1(n20248), .B2(n20277), .A(n20247), .ZN(P1_U2834) );
  NOR3_X1 U23273 ( .A1(n20271), .A2(n20249), .A3(P1_REIP_REG_5__SCAN_IN), .ZN(
        n20250) );
  AOI21_X1 U23274 ( .B1(n20263), .B2(P1_EBX_REG_5__SCAN_IN), .A(n20250), .ZN(
        n20260) );
  NOR2_X1 U23275 ( .A1(n20252), .A2(n20251), .ZN(n20274) );
  AOI22_X1 U23276 ( .A1(n20253), .A2(n20283), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n20274), .ZN(n20255) );
  OAI211_X1 U23277 ( .C1(n20257), .C2(n20256), .A(n20255), .B(n20254), .ZN(
        n20258) );
  AOI21_X1 U23278 ( .B1(n20284), .B2(n20272), .A(n20258), .ZN(n20259) );
  OAI211_X1 U23279 ( .C1(n20261), .C2(n20277), .A(n20260), .B(n20259), .ZN(
        P1_U2835) );
  INV_X1 U23280 ( .A(n20262), .ZN(n20264) );
  AOI22_X1 U23281 ( .A1(n20265), .A2(n20264), .B1(n20263), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n20266) );
  OAI21_X1 U23282 ( .B1(n20267), .B2(n20367), .A(n20266), .ZN(n20268) );
  AOI211_X1 U23283 ( .C1(n20269), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20349), .B(n20268), .ZN(n20276) );
  NAND3_X1 U23284 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n20270) );
  INV_X1 U23285 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20366) );
  OAI21_X1 U23286 ( .B1(n20271), .B2(n20270), .A(n20366), .ZN(n20273) );
  AOI22_X1 U23287 ( .A1(n20274), .A2(n20273), .B1(n20355), .B2(n20272), .ZN(
        n20275) );
  OAI211_X1 U23288 ( .C1(n20360), .C2(n20277), .A(n20276), .B(n20275), .ZN(
        P1_U2836) );
  AOI22_X1 U23289 ( .A1(n20279), .A2(n20708), .B1(n20706), .B2(n20278), .ZN(
        n20280) );
  OAI21_X1 U23290 ( .B1(n20282), .B2(n20281), .A(n20280), .ZN(P1_U2863) );
  AOI22_X1 U23291 ( .A1(n20284), .A2(n20708), .B1(n20706), .B2(n20283), .ZN(
        n20285) );
  OAI21_X1 U23292 ( .B1(n20282), .B2(n20286), .A(n20285), .ZN(P1_U2867) );
  INV_X1 U23293 ( .A(P1_UWORD_REG_2__SCAN_IN), .ZN(n20894) );
  INV_X1 U23294 ( .A(n20287), .ZN(n20288) );
  AOI22_X1 U23295 ( .A1(n20288), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n20318), .ZN(n20289) );
  OAI21_X1 U23296 ( .B1(n20894), .B2(n20698), .A(n20289), .ZN(P1_U2918) );
  AOI22_X1 U23297 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20297), .B1(n20318), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20290) );
  OAI21_X1 U23298 ( .B1(n20291), .B2(n20698), .A(n20290), .ZN(P1_U2921) );
  INV_X1 U23299 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20293) );
  AOI22_X1 U23300 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20292) );
  OAI21_X1 U23301 ( .B1(n20293), .B2(n20321), .A(n20292), .ZN(P1_U2922) );
  AOI22_X1 U23302 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(n20297), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20296), .ZN(n20294) );
  OAI21_X1 U23303 ( .B1(n20791), .B2(n20310), .A(n20294), .ZN(P1_U2923) );
  AOI22_X1 U23304 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20295) );
  OAI21_X1 U23305 ( .B1(n14291), .B2(n20321), .A(n20295), .ZN(P1_U2924) );
  AOI22_X1 U23306 ( .A1(P1_EAX_REG_11__SCAN_IN), .A2(n20297), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20296), .ZN(n20298) );
  OAI21_X1 U23307 ( .B1(n20733), .B2(n20310), .A(n20298), .ZN(P1_U2925) );
  INV_X1 U23308 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n20300) );
  AOI22_X1 U23309 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20299) );
  OAI21_X1 U23310 ( .B1(n20300), .B2(n20321), .A(n20299), .ZN(P1_U2926) );
  INV_X1 U23311 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20302) );
  AOI22_X1 U23312 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20301) );
  OAI21_X1 U23313 ( .B1(n20302), .B2(n20321), .A(n20301), .ZN(P1_U2927) );
  AOI22_X1 U23314 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20303) );
  OAI21_X1 U23315 ( .B1(n20304), .B2(n20321), .A(n20303), .ZN(P1_U2928) );
  INV_X1 U23316 ( .A(P1_LWORD_REG_7__SCAN_IN), .ZN(n20305) );
  INV_X1 U23317 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n20879) );
  OAI222_X1 U23318 ( .A1(n20698), .A2(n20305), .B1(n20321), .B2(n11833), .C1(
        n20879), .C2(n20310), .ZN(P1_U2929) );
  AOI22_X1 U23319 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20306) );
  OAI21_X1 U23320 ( .B1(n20307), .B2(n20321), .A(n20306), .ZN(P1_U2930) );
  AOI22_X1 U23321 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20308) );
  OAI21_X1 U23322 ( .B1(n13356), .B2(n20321), .A(n20308), .ZN(P1_U2931) );
  INV_X1 U23323 ( .A(P1_LWORD_REG_4__SCAN_IN), .ZN(n20815) );
  OAI222_X1 U23324 ( .A1(n20698), .A2(n20815), .B1(n20321), .B2(n20311), .C1(
        n20310), .C2(n20309), .ZN(P1_U2932) );
  AOI22_X1 U23325 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20312) );
  OAI21_X1 U23326 ( .B1(n20313), .B2(n20321), .A(n20312), .ZN(P1_U2933) );
  AOI22_X1 U23327 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20314) );
  OAI21_X1 U23328 ( .B1(n20315), .B2(n20321), .A(n20314), .ZN(P1_U2934) );
  AOI22_X1 U23329 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20316) );
  OAI21_X1 U23330 ( .B1(n20317), .B2(n20321), .A(n20316), .ZN(P1_U2935) );
  AOI22_X1 U23331 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20319), .B1(n20318), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20320) );
  OAI21_X1 U23332 ( .B1(n20322), .B2(n20321), .A(n20320), .ZN(P1_U2936) );
  AOI22_X1 U23333 ( .A1(n20323), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20345), .ZN(n20325) );
  NAND2_X1 U23334 ( .A1(n20333), .A2(n20324), .ZN(n20335) );
  NAND2_X1 U23335 ( .A1(n20325), .A2(n20335), .ZN(P1_U2946) );
  AOI22_X1 U23336 ( .A1(n20346), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20327) );
  NAND2_X1 U23337 ( .A1(n20333), .A2(n20326), .ZN(n20337) );
  NAND2_X1 U23338 ( .A1(n20327), .A2(n20337), .ZN(P1_U2947) );
  AOI22_X1 U23339 ( .A1(n20346), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20329) );
  NAND2_X1 U23340 ( .A1(n20333), .A2(n20328), .ZN(n20339) );
  NAND2_X1 U23341 ( .A1(n20329), .A2(n20339), .ZN(P1_U2948) );
  AOI22_X1 U23342 ( .A1(n20346), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20331) );
  NAND2_X1 U23343 ( .A1(n20333), .A2(n20330), .ZN(n20343) );
  NAND2_X1 U23344 ( .A1(n20331), .A2(n20343), .ZN(P1_U2950) );
  AOI22_X1 U23345 ( .A1(n20346), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20345), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20334) );
  NAND2_X1 U23346 ( .A1(n20333), .A2(n20332), .ZN(n20347) );
  NAND2_X1 U23347 ( .A1(n20334), .A2(n20347), .ZN(P1_U2951) );
  AOI22_X1 U23348 ( .A1(n20346), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20345), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20336) );
  NAND2_X1 U23349 ( .A1(n20336), .A2(n20335), .ZN(P1_U2961) );
  AOI22_X1 U23350 ( .A1(n20346), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20345), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20338) );
  NAND2_X1 U23351 ( .A1(n20338), .A2(n20337), .ZN(P1_U2962) );
  AOI22_X1 U23352 ( .A1(n20346), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20345), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20340) );
  NAND2_X1 U23353 ( .A1(n20340), .A2(n20339), .ZN(P1_U2963) );
  AOI22_X1 U23354 ( .A1(n20346), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20345), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20342) );
  NAND2_X1 U23355 ( .A1(n20342), .A2(n20341), .ZN(P1_U2964) );
  AOI22_X1 U23356 ( .A1(n20346), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20345), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20344) );
  NAND2_X1 U23357 ( .A1(n20344), .A2(n20343), .ZN(P1_U2965) );
  AOI22_X1 U23358 ( .A1(n20346), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20345), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20348) );
  NAND2_X1 U23359 ( .A1(n20348), .A2(n20347), .ZN(P1_U2966) );
  AOI22_X1 U23360 ( .A1(n20350), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20349), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20359) );
  OR2_X1 U23361 ( .A1(n20352), .A2(n20351), .ZN(n20353) );
  NAND2_X1 U23362 ( .A1(n20354), .A2(n20353), .ZN(n20365) );
  INV_X1 U23363 ( .A(n20365), .ZN(n20357) );
  AOI22_X1 U23364 ( .A1(n20357), .A2(n20356), .B1(n14067), .B2(n20355), .ZN(
        n20358) );
  OAI211_X1 U23365 ( .C1(n20361), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        P1_U2995) );
  NOR2_X1 U23366 ( .A1(n20363), .A2(n20362), .ZN(n20395) );
  NOR3_X1 U23367 ( .A1(n20384), .A2(n20395), .A3(n20383), .ZN(n20381) );
  AOI211_X1 U23368 ( .C1(n20963), .C2(n20380), .A(n20364), .B(n20375), .ZN(
        n20370) );
  NOR2_X1 U23369 ( .A1(n20365), .A2(n20385), .ZN(n20369) );
  OAI22_X1 U23370 ( .A1(n20392), .A2(n20367), .B1(n20366), .B2(n20254), .ZN(
        n20368) );
  NOR3_X1 U23371 ( .A1(n20370), .A2(n20369), .A3(n20368), .ZN(n20371) );
  OAI21_X1 U23372 ( .B1(n20381), .B2(n20963), .A(n20371), .ZN(P1_U3027) );
  AOI21_X1 U23373 ( .B1(n20374), .B2(n20373), .A(n20372), .ZN(n20379) );
  OAI22_X1 U23374 ( .A1(n20376), .A2(n20385), .B1(n20375), .B2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20377) );
  INV_X1 U23375 ( .A(n20377), .ZN(n20378) );
  OAI211_X1 U23376 ( .C1(n20381), .C2(n20380), .A(n20379), .B(n20378), .ZN(
        P1_U3028) );
  NAND2_X1 U23377 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20382), .ZN(
        n20399) );
  NOR2_X1 U23378 ( .A1(n20384), .A2(n20383), .ZN(n20398) );
  NOR3_X1 U23379 ( .A1(n20387), .A2(n20386), .A3(n20385), .ZN(n20396) );
  AND3_X1 U23380 ( .A1(n20389), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n20388), .ZN(n20394) );
  OAI21_X1 U23381 ( .B1(n20392), .B2(n20391), .A(n20390), .ZN(n20393) );
  NOR4_X1 U23382 ( .A1(n20396), .A2(n20395), .A3(n20394), .A4(n20393), .ZN(
        n20397) );
  OAI221_X1 U23383 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20399), .C1(
        n20962), .C2(n20398), .A(n20397), .ZN(P1_U3029) );
  AND2_X1 U23384 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20400), .ZN(
        P1_U3032) );
  AOI22_X1 U23385 ( .A1(n9857), .A2(n20415), .B1(n20414), .B2(n20461), .ZN(
        n20403) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20417), .B1(
        n20567), .B2(n20416), .ZN(n20402) );
  OAI211_X1 U23387 ( .C1(n20464), .C2(n20447), .A(n20403), .B(n20402), .ZN(
        P1_U3034) );
  AOI22_X1 U23388 ( .A1(n20574), .A2(n20415), .B1(n20414), .B2(n20465), .ZN(
        n20405) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20417), .B1(
        n20573), .B2(n20416), .ZN(n20404) );
  OAI211_X1 U23390 ( .C1(n20468), .C2(n20447), .A(n20405), .B(n20404), .ZN(
        P1_U3035) );
  AOI22_X1 U23391 ( .A1(n20580), .A2(n20415), .B1(n20414), .B2(n20469), .ZN(
        n20407) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20417), .B1(
        n20579), .B2(n20416), .ZN(n20406) );
  OAI211_X1 U23393 ( .C1(n20472), .C2(n20447), .A(n20407), .B(n20406), .ZN(
        P1_U3036) );
  AOI22_X1 U23394 ( .A1(n20586), .A2(n20415), .B1(n20414), .B2(n20473), .ZN(
        n20409) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20417), .B1(
        n20585), .B2(n20416), .ZN(n20408) );
  OAI211_X1 U23396 ( .C1(n20476), .C2(n20447), .A(n20409), .B(n20408), .ZN(
        P1_U3037) );
  AOI22_X1 U23397 ( .A1(n20592), .A2(n20415), .B1(n20414), .B2(n20477), .ZN(
        n20411) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20417), .B1(
        n20591), .B2(n20416), .ZN(n20410) );
  OAI211_X1 U23399 ( .C1(n20480), .C2(n20447), .A(n20411), .B(n20410), .ZN(
        P1_U3038) );
  AOI22_X1 U23400 ( .A1(n20598), .A2(n20415), .B1(n20414), .B2(n20481), .ZN(
        n20413) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20417), .B1(
        n20597), .B2(n20416), .ZN(n20412) );
  OAI211_X1 U23402 ( .C1(n20484), .C2(n20447), .A(n20413), .B(n20412), .ZN(
        P1_U3039) );
  AOI22_X1 U23403 ( .A1(n20606), .A2(n20415), .B1(n20414), .B2(n20487), .ZN(
        n20419) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20417), .B1(
        n20604), .B2(n20416), .ZN(n20418) );
  OAI211_X1 U23405 ( .C1(n20492), .C2(n20447), .A(n20419), .B(n20418), .ZN(
        P1_U3040) );
  NOR2_X1 U23406 ( .A1(n20549), .A2(n20422), .ZN(n20442) );
  INV_X1 U23407 ( .A(n20420), .ZN(n20550) );
  AOI21_X1 U23408 ( .B1(n20421), .B2(n20550), .A(n20442), .ZN(n20423) );
  OAI22_X1 U23409 ( .A1(n20423), .A2(n20559), .B1(n20422), .B2(n20616), .ZN(
        n20441) );
  AOI22_X1 U23410 ( .A1(n20554), .A2(n20442), .B1(n20441), .B2(n20553), .ZN(
        n20428) );
  OAI21_X1 U23411 ( .B1(n20424), .B2(n20524), .A(n20423), .ZN(n20425) );
  OAI221_X1 U23412 ( .B1(n20561), .B2(n20426), .C1(n20559), .C2(n20425), .A(
        n20557), .ZN(n20444) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20563), .ZN(n20427) );
  OAI211_X1 U23414 ( .C1(n20566), .C2(n20447), .A(n20428), .B(n20427), .ZN(
        P1_U3041) );
  AOI22_X1 U23415 ( .A1(n9857), .A2(n20442), .B1(n20441), .B2(n20567), .ZN(
        n20430) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20569), .ZN(n20429) );
  OAI211_X1 U23417 ( .C1(n20572), .C2(n20447), .A(n20430), .B(n20429), .ZN(
        P1_U3042) );
  AOI22_X1 U23418 ( .A1(n20574), .A2(n20442), .B1(n20441), .B2(n20573), .ZN(
        n20432) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20575), .ZN(n20431) );
  OAI211_X1 U23420 ( .C1(n20578), .C2(n20447), .A(n20432), .B(n20431), .ZN(
        P1_U3043) );
  AOI22_X1 U23421 ( .A1(n20580), .A2(n20442), .B1(n20441), .B2(n20579), .ZN(
        n20434) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20581), .ZN(n20433) );
  OAI211_X1 U23423 ( .C1(n20584), .C2(n20447), .A(n20434), .B(n20433), .ZN(
        P1_U3044) );
  AOI22_X1 U23424 ( .A1(n20586), .A2(n20442), .B1(n20441), .B2(n20585), .ZN(
        n20436) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20587), .ZN(n20435) );
  OAI211_X1 U23426 ( .C1(n20590), .C2(n20447), .A(n20436), .B(n20435), .ZN(
        P1_U3045) );
  AOI22_X1 U23427 ( .A1(n20592), .A2(n20442), .B1(n20441), .B2(n20591), .ZN(
        n20438) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20593), .ZN(n20437) );
  OAI211_X1 U23429 ( .C1(n20596), .C2(n20447), .A(n20438), .B(n20437), .ZN(
        P1_U3046) );
  AOI22_X1 U23430 ( .A1(n20598), .A2(n20442), .B1(n20597), .B2(n20441), .ZN(
        n20440) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20599), .ZN(n20439) );
  OAI211_X1 U23432 ( .C1(n20602), .C2(n20447), .A(n20440), .B(n20439), .ZN(
        P1_U3047) );
  AOI22_X1 U23433 ( .A1(n20606), .A2(n20442), .B1(n20441), .B2(n20604), .ZN(
        n20446) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20444), .B1(
        n20443), .B2(n20607), .ZN(n20445) );
  OAI211_X1 U23435 ( .C1(n20613), .C2(n20447), .A(n20446), .B(n20445), .ZN(
        P1_U3048) );
  NOR3_X1 U23436 ( .A1(n20788), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20498) );
  INV_X1 U23437 ( .A(n20498), .ZN(n20494) );
  NOR2_X1 U23438 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20494), .ZN(
        n20486) );
  NAND3_X1 U23439 ( .A1(n20493), .A2(n20561), .A3(n12613), .ZN(n20449) );
  OAI21_X1 U23440 ( .B1(n20451), .B2(n20450), .A(n20449), .ZN(n20485) );
  AOI22_X1 U23441 ( .A1(n20554), .A2(n20486), .B1(n20553), .B2(n20485), .ZN(
        n20459) );
  AOI21_X1 U23442 ( .B1(n20456), .B2(n20519), .A(n20818), .ZN(n20452) );
  AOI21_X1 U23443 ( .B1(n20493), .B2(n12613), .A(n20452), .ZN(n20453) );
  NOR2_X1 U23444 ( .A1(n20453), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20455) );
  AOI22_X1 U23445 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n20488), .B2(n20457), .ZN(n20458) );
  OAI211_X1 U23446 ( .C1(n20460), .C2(n20519), .A(n20459), .B(n20458), .ZN(
        P1_U3065) );
  AOI22_X1 U23447 ( .A1(n9857), .A2(n20486), .B1(n20567), .B2(n20485), .ZN(
        n20463) );
  AOI22_X1 U23448 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n20488), .B2(n20461), .ZN(n20462) );
  OAI211_X1 U23449 ( .C1(n20464), .C2(n20519), .A(n20463), .B(n20462), .ZN(
        P1_U3066) );
  AOI22_X1 U23450 ( .A1(n20574), .A2(n20486), .B1(n20573), .B2(n20485), .ZN(
        n20467) );
  AOI22_X1 U23451 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n20488), .B2(n20465), .ZN(n20466) );
  OAI211_X1 U23452 ( .C1(n20468), .C2(n20519), .A(n20467), .B(n20466), .ZN(
        P1_U3067) );
  AOI22_X1 U23453 ( .A1(n20580), .A2(n20486), .B1(n20579), .B2(n20485), .ZN(
        n20471) );
  AOI22_X1 U23454 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n20488), .B2(n20469), .ZN(n20470) );
  OAI211_X1 U23455 ( .C1(n20472), .C2(n20519), .A(n20471), .B(n20470), .ZN(
        P1_U3068) );
  AOI22_X1 U23456 ( .A1(n20586), .A2(n20486), .B1(n20585), .B2(n20485), .ZN(
        n20475) );
  AOI22_X1 U23457 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n20488), .B2(n20473), .ZN(n20474) );
  OAI211_X1 U23458 ( .C1(n20476), .C2(n20519), .A(n20475), .B(n20474), .ZN(
        P1_U3069) );
  AOI22_X1 U23459 ( .A1(n20592), .A2(n20486), .B1(n20591), .B2(n20485), .ZN(
        n20479) );
  AOI22_X1 U23460 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n20488), .B2(n20477), .ZN(n20478) );
  OAI211_X1 U23461 ( .C1(n20480), .C2(n20519), .A(n20479), .B(n20478), .ZN(
        P1_U3070) );
  AOI22_X1 U23462 ( .A1(n20598), .A2(n20486), .B1(n20597), .B2(n20485), .ZN(
        n20483) );
  AOI22_X1 U23463 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n20488), .B2(n20481), .ZN(n20482) );
  OAI211_X1 U23464 ( .C1(n20484), .C2(n20519), .A(n20483), .B(n20482), .ZN(
        P1_U3071) );
  AOI22_X1 U23465 ( .A1(n20606), .A2(n20486), .B1(n20604), .B2(n20485), .ZN(
        n20491) );
  AOI22_X1 U23466 ( .A1(n20489), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n20488), .B2(n20487), .ZN(n20490) );
  OAI211_X1 U23467 ( .C1(n20492), .C2(n20519), .A(n20491), .B(n20490), .ZN(
        P1_U3072) );
  NOR2_X1 U23468 ( .A1(n20549), .A2(n20494), .ZN(n20514) );
  AOI21_X1 U23469 ( .B1(n20493), .B2(n20550), .A(n20514), .ZN(n20495) );
  OAI22_X1 U23470 ( .A1(n20495), .A2(n20559), .B1(n20494), .B2(n20616), .ZN(
        n20513) );
  AOI22_X1 U23471 ( .A1(n20554), .A2(n20514), .B1(n20553), .B2(n20513), .ZN(
        n20500) );
  OAI21_X1 U23472 ( .B1(n20496), .B2(n20524), .A(n20495), .ZN(n20497) );
  OAI221_X1 U23473 ( .B1(n20561), .B2(n20498), .C1(n20559), .C2(n20497), .A(
        n20557), .ZN(n20516) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20563), .ZN(n20499) );
  OAI211_X1 U23475 ( .C1(n20566), .C2(n20519), .A(n20500), .B(n20499), .ZN(
        P1_U3073) );
  AOI22_X1 U23476 ( .A1(n9857), .A2(n20514), .B1(n20567), .B2(n20513), .ZN(
        n20502) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20569), .ZN(n20501) );
  OAI211_X1 U23478 ( .C1(n20572), .C2(n20519), .A(n20502), .B(n20501), .ZN(
        P1_U3074) );
  AOI22_X1 U23479 ( .A1(n20574), .A2(n20514), .B1(n20573), .B2(n20513), .ZN(
        n20504) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20575), .ZN(n20503) );
  OAI211_X1 U23481 ( .C1(n20578), .C2(n20519), .A(n20504), .B(n20503), .ZN(
        P1_U3075) );
  AOI22_X1 U23482 ( .A1(n20580), .A2(n20514), .B1(n20579), .B2(n20513), .ZN(
        n20506) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20581), .ZN(n20505) );
  OAI211_X1 U23484 ( .C1(n20584), .C2(n20519), .A(n20506), .B(n20505), .ZN(
        P1_U3076) );
  AOI22_X1 U23485 ( .A1(n20586), .A2(n20514), .B1(n20585), .B2(n20513), .ZN(
        n20508) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20587), .ZN(n20507) );
  OAI211_X1 U23487 ( .C1(n20590), .C2(n20519), .A(n20508), .B(n20507), .ZN(
        P1_U3077) );
  AOI22_X1 U23488 ( .A1(n20592), .A2(n20514), .B1(n20591), .B2(n20513), .ZN(
        n20510) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20593), .ZN(n20509) );
  OAI211_X1 U23490 ( .C1(n20596), .C2(n20519), .A(n20510), .B(n20509), .ZN(
        P1_U3078) );
  AOI22_X1 U23491 ( .A1(n20598), .A2(n20514), .B1(n20597), .B2(n20513), .ZN(
        n20512) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20599), .ZN(n20511) );
  OAI211_X1 U23493 ( .C1(n20602), .C2(n20519), .A(n20512), .B(n20511), .ZN(
        P1_U3079) );
  AOI22_X1 U23494 ( .A1(n20606), .A2(n20514), .B1(n20604), .B2(n20513), .ZN(
        n20518) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20516), .B1(
        n20515), .B2(n20607), .ZN(n20517) );
  OAI211_X1 U23496 ( .C1(n20613), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P1_U3080) );
  NOR2_X1 U23497 ( .A1(n20549), .A2(n20522), .ZN(n20543) );
  INV_X1 U23498 ( .A(n20520), .ZN(n20521) );
  AOI21_X1 U23499 ( .B1(n20521), .B2(n20550), .A(n20543), .ZN(n20523) );
  OAI22_X1 U23500 ( .A1(n20523), .A2(n20559), .B1(n20522), .B2(n20616), .ZN(
        n20542) );
  AOI22_X1 U23501 ( .A1(n20554), .A2(n20543), .B1(n20542), .B2(n20553), .ZN(
        n20529) );
  OAI21_X1 U23502 ( .B1(n20525), .B2(n20524), .A(n20523), .ZN(n20526) );
  OAI221_X1 U23503 ( .B1(n20561), .B2(n20527), .C1(n20559), .C2(n20526), .A(
        n20557), .ZN(n20545) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20563), .ZN(n20528) );
  OAI211_X1 U23505 ( .C1(n20566), .C2(n20548), .A(n20529), .B(n20528), .ZN(
        P1_U3105) );
  AOI22_X1 U23506 ( .A1(n9857), .A2(n20543), .B1(n20542), .B2(n20567), .ZN(
        n20531) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20569), .ZN(n20530) );
  OAI211_X1 U23508 ( .C1(n20572), .C2(n20548), .A(n20531), .B(n20530), .ZN(
        P1_U3106) );
  AOI22_X1 U23509 ( .A1(n20574), .A2(n20543), .B1(n20542), .B2(n20573), .ZN(
        n20533) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20575), .ZN(n20532) );
  OAI211_X1 U23511 ( .C1(n20578), .C2(n20548), .A(n20533), .B(n20532), .ZN(
        P1_U3107) );
  AOI22_X1 U23512 ( .A1(n20580), .A2(n20543), .B1(n20542), .B2(n20579), .ZN(
        n20535) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20581), .ZN(n20534) );
  OAI211_X1 U23514 ( .C1(n20584), .C2(n20548), .A(n20535), .B(n20534), .ZN(
        P1_U3108) );
  AOI22_X1 U23515 ( .A1(n20586), .A2(n20543), .B1(n20542), .B2(n20585), .ZN(
        n20537) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20587), .ZN(n20536) );
  OAI211_X1 U23517 ( .C1(n20590), .C2(n20548), .A(n20537), .B(n20536), .ZN(
        P1_U3109) );
  AOI22_X1 U23518 ( .A1(n20592), .A2(n20543), .B1(n20542), .B2(n20591), .ZN(
        n20539) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20593), .ZN(n20538) );
  OAI211_X1 U23520 ( .C1(n20596), .C2(n20548), .A(n20539), .B(n20538), .ZN(
        P1_U3110) );
  AOI22_X1 U23521 ( .A1(n20598), .A2(n20543), .B1(n20597), .B2(n20542), .ZN(
        n20541) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20599), .ZN(n20540) );
  OAI211_X1 U23523 ( .C1(n20602), .C2(n20548), .A(n20541), .B(n20540), .ZN(
        P1_U3111) );
  AOI22_X1 U23524 ( .A1(n20606), .A2(n20543), .B1(n20542), .B2(n20604), .ZN(
        n20547) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20545), .B1(
        n20544), .B2(n20607), .ZN(n20546) );
  OAI211_X1 U23526 ( .C1(n20613), .C2(n20548), .A(n20547), .B(n20546), .ZN(
        P1_U3112) );
  INV_X1 U23527 ( .A(n20560), .ZN(n20552) );
  NOR2_X1 U23528 ( .A1(n20549), .A2(n20552), .ZN(n20605) );
  AOI21_X1 U23529 ( .B1(n20551), .B2(n20550), .A(n20605), .ZN(n20555) );
  OAI22_X1 U23530 ( .A1(n20555), .A2(n20559), .B1(n20552), .B2(n20616), .ZN(
        n20603) );
  AOI22_X1 U23531 ( .A1(n20554), .A2(n20605), .B1(n20553), .B2(n20603), .ZN(
        n20565) );
  NAND2_X1 U23532 ( .A1(n20556), .A2(n20555), .ZN(n20558) );
  OAI221_X1 U23533 ( .B1(n20561), .B2(n20560), .C1(n20559), .C2(n20558), .A(
        n20557), .ZN(n20609) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20563), .ZN(n20564) );
  OAI211_X1 U23535 ( .C1(n20566), .C2(n20612), .A(n20565), .B(n20564), .ZN(
        P1_U3137) );
  AOI22_X1 U23536 ( .A1(n9857), .A2(n20605), .B1(n20567), .B2(n20603), .ZN(
        n20571) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20569), .ZN(n20570) );
  OAI211_X1 U23538 ( .C1(n20572), .C2(n20612), .A(n20571), .B(n20570), .ZN(
        P1_U3138) );
  AOI22_X1 U23539 ( .A1(n20574), .A2(n20605), .B1(n20573), .B2(n20603), .ZN(
        n20577) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20575), .ZN(n20576) );
  OAI211_X1 U23541 ( .C1(n20578), .C2(n20612), .A(n20577), .B(n20576), .ZN(
        P1_U3139) );
  AOI22_X1 U23542 ( .A1(n20580), .A2(n20605), .B1(n20579), .B2(n20603), .ZN(
        n20583) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20581), .ZN(n20582) );
  OAI211_X1 U23544 ( .C1(n20584), .C2(n20612), .A(n20583), .B(n20582), .ZN(
        P1_U3140) );
  AOI22_X1 U23545 ( .A1(n20586), .A2(n20605), .B1(n20585), .B2(n20603), .ZN(
        n20589) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20587), .ZN(n20588) );
  OAI211_X1 U23547 ( .C1(n20590), .C2(n20612), .A(n20589), .B(n20588), .ZN(
        P1_U3141) );
  AOI22_X1 U23548 ( .A1(n20592), .A2(n20605), .B1(n20591), .B2(n20603), .ZN(
        n20595) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20593), .ZN(n20594) );
  OAI211_X1 U23550 ( .C1(n20596), .C2(n20612), .A(n20595), .B(n20594), .ZN(
        P1_U3142) );
  AOI22_X1 U23551 ( .A1(n20598), .A2(n20605), .B1(n20597), .B2(n20603), .ZN(
        n20601) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20599), .ZN(n20600) );
  OAI211_X1 U23553 ( .C1(n20602), .C2(n20612), .A(n20601), .B(n20600), .ZN(
        P1_U3143) );
  AOI22_X1 U23554 ( .A1(n20606), .A2(n20605), .B1(n20604), .B2(n20603), .ZN(
        n20611) );
  AOI22_X1 U23555 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20609), .B1(
        n20608), .B2(n20607), .ZN(n20610) );
  OAI211_X1 U23556 ( .C1(n20613), .C2(n20612), .A(n20611), .B(n20610), .ZN(
        P1_U3144) );
  NOR2_X1 U23557 ( .A1(n10118), .A2(n20614), .ZN(n20617) );
  OAI21_X1 U23558 ( .B1(n20617), .B2(n20616), .A(n20615), .ZN(P1_U3163) );
  INV_X1 U23559 ( .A(n20683), .ZN(n20618) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20618), .ZN(
        P1_U3164) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20618), .ZN(
        P1_U3165) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20618), .ZN(
        P1_U3166) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20618), .ZN(
        P1_U3167) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20618), .ZN(
        P1_U3168) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20618), .ZN(
        P1_U3169) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20618), .ZN(
        P1_U3170) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20618), .ZN(
        P1_U3171) );
  AND2_X1 U23568 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20618), .ZN(
        P1_U3172) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20618), .ZN(
        P1_U3173) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20618), .ZN(
        P1_U3174) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20618), .ZN(
        P1_U3175) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20618), .ZN(
        P1_U3176) );
  NOR2_X1 U23573 ( .A1(n20683), .A2(n20863), .ZN(P1_U3177) );
  AND2_X1 U23574 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20618), .ZN(
        P1_U3178) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20618), .ZN(
        P1_U3179) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20618), .ZN(
        P1_U3180) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20618), .ZN(
        P1_U3181) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20618), .ZN(
        P1_U3182) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20618), .ZN(
        P1_U3183) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20618), .ZN(
        P1_U3184) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20618), .ZN(
        P1_U3185) );
  INV_X1 U23582 ( .A(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20945) );
  NOR2_X1 U23583 ( .A1(n20683), .A2(n20945), .ZN(P1_U3186) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20618), .ZN(P1_U3187) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20618), .ZN(P1_U3188) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20618), .ZN(P1_U3189) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20618), .ZN(P1_U3190) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20618), .ZN(P1_U3191) );
  NOR2_X1 U23589 ( .A1(n20683), .A2(n20619), .ZN(P1_U3192) );
  INV_X1 U23590 ( .A(P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n20775) );
  NOR2_X1 U23591 ( .A1(n20683), .A2(n20775), .ZN(P1_U3193) );
  NAND2_X1 U23592 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20623), .ZN(n20628) );
  INV_X1 U23593 ( .A(n20628), .ZN(n20622) );
  INV_X1 U23594 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20971) );
  AOI21_X1 U23595 ( .B1(n20632), .B2(n20971), .A(n20624), .ZN(n20620) );
  INV_X1 U23596 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20704) );
  AOI211_X1 U23597 ( .C1(NA), .C2(n12770), .A(n20620), .B(n20704), .ZN(n20621)
         );
  OAI22_X1 U23598 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20622), .B1(n20693), 
        .B2(n20621), .ZN(P1_U3194) );
  NOR3_X1 U23599 ( .A1(NA), .A2(n12770), .A3(n20623), .ZN(n20627) );
  AOI21_X1 U23600 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n20632), .A(n20624), .ZN(n20626) );
  AOI222_X1 U23601 ( .A1(n20627), .A2(n20626), .B1(n20627), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(n20626), .C2(n20625), .ZN(n20631)
         );
  OAI211_X1 U23602 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20629), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20628), .ZN(n20630) );
  NAND2_X1 U23603 ( .A1(n20631), .A2(n20630), .ZN(P1_U3196) );
  INV_X1 U23604 ( .A(n9720), .ZN(n20671) );
  NAND2_X1 U23605 ( .A1(n20632), .A2(n20693), .ZN(n20675) );
  INV_X1 U23606 ( .A(n20675), .ZN(n20669) );
  AOI22_X1 U23607 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20669), .ZN(n20633) );
  OAI21_X1 U23608 ( .B1(n13275), .B2(n20671), .A(n20633), .ZN(P1_U3197) );
  INV_X1 U23609 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20635) );
  AOI22_X1 U23610 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20669), .ZN(n20634) );
  OAI21_X1 U23611 ( .B1(n20635), .B2(n20671), .A(n20634), .ZN(P1_U3198) );
  INV_X1 U23612 ( .A(n20636), .ZN(P1_U3199) );
  AOI222_X1 U23613 ( .A1(n20669), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n9720), .ZN(n20637) );
  INV_X1 U23614 ( .A(n20637), .ZN(P1_U3200) );
  INV_X1 U23615 ( .A(n20638), .ZN(P1_U3201) );
  AOI222_X1 U23616 ( .A1(n20669), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n9720), .ZN(n20639) );
  INV_X1 U23617 ( .A(n20639), .ZN(P1_U3202) );
  INV_X1 U23618 ( .A(n20640), .ZN(P1_U3203) );
  AOI222_X1 U23619 ( .A1(n9720), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20669), .ZN(n20641) );
  INV_X1 U23620 ( .A(n20641), .ZN(P1_U3204) );
  AOI222_X1 U23621 ( .A1(n9720), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20669), .ZN(n20642) );
  INV_X1 U23622 ( .A(n20642), .ZN(P1_U3205) );
  AOI22_X1 U23623 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20669), .ZN(n20643) );
  OAI21_X1 U23624 ( .B1(n20644), .B2(n20671), .A(n20643), .ZN(P1_U3206) );
  INV_X1 U23625 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20646) );
  AOI22_X1 U23626 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20669), .ZN(n20645) );
  OAI21_X1 U23627 ( .B1(n20646), .B2(n20671), .A(n20645), .ZN(P1_U3207) );
  AOI22_X1 U23628 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n9720), .ZN(n20647) );
  OAI21_X1 U23629 ( .B1(n20649), .B2(n20675), .A(n20647), .ZN(P1_U3208) );
  AOI22_X1 U23630 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20669), .ZN(n20648) );
  OAI21_X1 U23631 ( .B1(n20649), .B2(n20671), .A(n20648), .ZN(P1_U3209) );
  AOI22_X1 U23632 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n9720), .ZN(n20650) );
  OAI21_X1 U23633 ( .B1(n15114), .B2(n20675), .A(n20650), .ZN(P1_U3210) );
  AOI222_X1 U23634 ( .A1(n9720), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20669), .ZN(n20651) );
  INV_X1 U23635 ( .A(n20651), .ZN(P1_U3211) );
  AOI22_X1 U23636 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20669), .ZN(n20652) );
  OAI21_X1 U23637 ( .B1(n15284), .B2(n20671), .A(n20652), .ZN(P1_U3212) );
  AOI22_X1 U23638 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n9720), .ZN(n20653) );
  OAI21_X1 U23639 ( .B1(n20654), .B2(n20675), .A(n20653), .ZN(P1_U3213) );
  AOI222_X1 U23640 ( .A1(n9720), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20669), .ZN(n20655) );
  INV_X1 U23641 ( .A(n20655), .ZN(P1_U3214) );
  AOI22_X1 U23642 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20669), .ZN(n20656) );
  OAI21_X1 U23643 ( .B1(n20657), .B2(n20671), .A(n20656), .ZN(P1_U3215) );
  AOI22_X1 U23644 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n9720), .ZN(n20658) );
  OAI21_X1 U23645 ( .B1(n15066), .B2(n20675), .A(n20658), .ZN(P1_U3216) );
  AOI222_X1 U23646 ( .A1(n20669), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n9720), .ZN(n20659) );
  INV_X1 U23647 ( .A(n20659), .ZN(P1_U3217) );
  AOI22_X1 U23648 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20669), .ZN(n20660) );
  OAI21_X1 U23649 ( .B1(n20661), .B2(n20671), .A(n20660), .ZN(P1_U3218) );
  AOI22_X1 U23650 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20691), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n9720), .ZN(n20662) );
  OAI21_X1 U23651 ( .B1(n20663), .B2(n20675), .A(n20662), .ZN(P1_U3219) );
  AOI222_X1 U23652 ( .A1(n9720), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20669), .ZN(n20664) );
  INV_X1 U23653 ( .A(n20664), .ZN(P1_U3220) );
  AOI222_X1 U23654 ( .A1(n9720), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20669), .ZN(n20665) );
  INV_X1 U23655 ( .A(n20665), .ZN(P1_U3221) );
  AOI222_X1 U23656 ( .A1(n9720), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20669), .ZN(n20666) );
  INV_X1 U23657 ( .A(n20666), .ZN(P1_U3222) );
  AOI222_X1 U23658 ( .A1(n9720), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20669), .ZN(n20667) );
  INV_X1 U23659 ( .A(n20667), .ZN(P1_U3223) );
  AOI222_X1 U23660 ( .A1(n9720), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20691), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20669), .ZN(n20668) );
  INV_X1 U23661 ( .A(n20668), .ZN(P1_U3224) );
  AOI22_X1 U23662 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20669), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20691), .ZN(n20670) );
  OAI21_X1 U23663 ( .B1(n20672), .B2(n20671), .A(n20670), .ZN(P1_U3225) );
  AOI22_X1 U23664 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n9720), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20691), .ZN(n20674) );
  OAI21_X1 U23665 ( .B1(n20986), .B2(n20675), .A(n20674), .ZN(P1_U3226) );
  OAI22_X1 U23666 ( .A1(n20691), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20693), .ZN(n20676) );
  INV_X1 U23667 ( .A(n20676), .ZN(P1_U3458) );
  OAI22_X1 U23668 ( .A1(n20691), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20693), .ZN(n20677) );
  INV_X1 U23669 ( .A(n20677), .ZN(P1_U3459) );
  OAI22_X1 U23670 ( .A1(n20691), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20693), .ZN(n20678) );
  INV_X1 U23671 ( .A(n20678), .ZN(P1_U3460) );
  OAI22_X1 U23672 ( .A1(n20691), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20693), .ZN(n20679) );
  INV_X1 U23673 ( .A(n20679), .ZN(P1_U3461) );
  OAI21_X1 U23674 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20683), .A(n20681), 
        .ZN(n20680) );
  INV_X1 U23675 ( .A(n20680), .ZN(P1_U3464) );
  OAI21_X1 U23676 ( .B1(n20683), .B2(n20682), .A(n20681), .ZN(P1_U3465) );
  AOI21_X1 U23677 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20684) );
  AOI22_X1 U23678 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20684), .B2(n13275), .ZN(n20686) );
  INV_X1 U23679 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20685) );
  AOI22_X1 U23680 ( .A1(n20687), .A2(n20686), .B1(n20685), .B2(n20689), .ZN(
        P1_U3481) );
  INV_X1 U23681 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20690) );
  NOR2_X1 U23682 ( .A1(n20689), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20688) );
  AOI22_X1 U23683 ( .A1(n20690), .A2(n20689), .B1(n13049), .B2(n20688), .ZN(
        P1_U3482) );
  AOI22_X1 U23684 ( .A1(n20693), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20692), 
        .B2(n20691), .ZN(P1_U3483) );
  INV_X1 U23685 ( .A(n20694), .ZN(n20695) );
  OAI211_X1 U23686 ( .C1(n20698), .C2(n20697), .A(n20696), .B(n20695), .ZN(
        n20705) );
  OAI211_X1 U23687 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20700), .A(n20699), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20701) );
  NAND3_X1 U23688 ( .A1(n20705), .A2(n20702), .A3(n20701), .ZN(n20703) );
  OAI21_X1 U23689 ( .B1(n20705), .B2(n20704), .A(n20703), .ZN(P1_U3485) );
  MUX2_X1 U23690 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20691), .Z(P1_U3486) );
  AOI222_X1 U23691 ( .A1(n20709), .A2(n20708), .B1(n20707), .B2(
        P1_EBX_REG_12__SCAN_IN), .C1(n20706), .C2(n9820), .ZN(n20959) );
  INV_X1 U23692 ( .A(READY22_REG_SCAN_IN), .ZN(n20711) );
  AOI22_X1 U23693 ( .A1(n20712), .A2(keyinput77), .B1(keyinput98), .B2(n20711), 
        .ZN(n20710) );
  OAI221_X1 U23694 ( .B1(n20712), .B2(keyinput77), .C1(n20711), .C2(keyinput98), .A(n20710), .ZN(n20723) );
  INV_X1 U23695 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n20978) );
  AOI22_X1 U23696 ( .A1(n20978), .A2(keyinput21), .B1(keyinput97), .B2(n20964), 
        .ZN(n20713) );
  OAI221_X1 U23697 ( .B1(n20978), .B2(keyinput21), .C1(n20964), .C2(keyinput97), .A(n20713), .ZN(n20722) );
  INV_X1 U23698 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20715) );
  AOI22_X1 U23699 ( .A1(n20716), .A2(keyinput96), .B1(n20715), .B2(keyinput35), 
        .ZN(n20714) );
  OAI221_X1 U23700 ( .B1(n20716), .B2(keyinput96), .C1(n20715), .C2(keyinput35), .A(n20714), .ZN(n20721) );
  AOI22_X1 U23701 ( .A1(n20719), .A2(keyinput84), .B1(keyinput99), .B2(n20718), 
        .ZN(n20717) );
  OAI221_X1 U23702 ( .B1(n20719), .B2(keyinput84), .C1(n20718), .C2(keyinput99), .A(n20717), .ZN(n20720) );
  NOR4_X1 U23703 ( .A1(n20723), .A2(n20722), .A3(n20721), .A4(n20720), .ZN(
        n20767) );
  AOI22_X1 U23704 ( .A1(n20725), .A2(keyinput111), .B1(n14603), .B2(keyinput28), .ZN(n20724) );
  OAI221_X1 U23705 ( .B1(n20725), .B2(keyinput111), .C1(n14603), .C2(
        keyinput28), .A(n20724), .ZN(n20729) );
  XOR2_X1 U23706 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B(keyinput107), .Z(
        n20728) );
  XNOR2_X1 U23707 ( .A(n20726), .B(keyinput83), .ZN(n20727) );
  OR3_X1 U23708 ( .A1(n20729), .A2(n20728), .A3(n20727), .ZN(n20736) );
  AOI22_X1 U23709 ( .A1(n20970), .A2(keyinput19), .B1(keyinput73), .B2(n20731), 
        .ZN(n20730) );
  OAI221_X1 U23710 ( .B1(n20970), .B2(keyinput19), .C1(n20731), .C2(keyinput73), .A(n20730), .ZN(n20735) );
  AOI22_X1 U23711 ( .A1(n13868), .A2(keyinput54), .B1(n20733), .B2(keyinput37), 
        .ZN(n20732) );
  OAI221_X1 U23712 ( .B1(n13868), .B2(keyinput54), .C1(n20733), .C2(keyinput37), .A(n20732), .ZN(n20734) );
  NOR3_X1 U23713 ( .A1(n20736), .A2(n20735), .A3(n20734), .ZN(n20766) );
  AOI22_X1 U23714 ( .A1(n20738), .A2(keyinput126), .B1(n20999), .B2(keyinput56), .ZN(n20737) );
  OAI221_X1 U23715 ( .B1(n20738), .B2(keyinput126), .C1(n20999), .C2(
        keyinput56), .A(n20737), .ZN(n20749) );
  INV_X1 U23716 ( .A(DATAI_23_), .ZN(n20740) );
  AOI22_X1 U23717 ( .A1(n20741), .A2(keyinput41), .B1(n20740), .B2(keyinput61), 
        .ZN(n20739) );
  OAI221_X1 U23718 ( .B1(n20741), .B2(keyinput41), .C1(n20740), .C2(keyinput61), .A(n20739), .ZN(n20748) );
  AOI22_X1 U23719 ( .A1(n20971), .A2(keyinput9), .B1(n20743), .B2(keyinput122), 
        .ZN(n20742) );
  OAI221_X1 U23720 ( .B1(n20971), .B2(keyinput9), .C1(n20743), .C2(keyinput122), .A(n20742), .ZN(n20747) );
  XOR2_X1 U23721 ( .A(n14484), .B(keyinput68), .Z(n20745) );
  XNOR2_X1 U23722 ( .A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B(keyinput32), .ZN(
        n20744) );
  NAND2_X1 U23723 ( .A1(n20745), .A2(n20744), .ZN(n20746) );
  NOR4_X1 U23724 ( .A1(n20749), .A2(n20748), .A3(n20747), .A4(n20746), .ZN(
        n20765) );
  AOI22_X1 U23725 ( .A1(n20751), .A2(keyinput10), .B1(n14094), .B2(keyinput85), 
        .ZN(n20750) );
  OAI221_X1 U23726 ( .B1(n20751), .B2(keyinput10), .C1(n14094), .C2(keyinput85), .A(n20750), .ZN(n20763) );
  AOI22_X1 U23727 ( .A1(n20754), .A2(keyinput120), .B1(n20753), .B2(keyinput31), .ZN(n20752) );
  OAI221_X1 U23728 ( .B1(n20754), .B2(keyinput120), .C1(n20753), .C2(
        keyinput31), .A(n20752), .ZN(n20762) );
  INV_X1 U23729 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20965) );
  AOI22_X1 U23730 ( .A1(n20756), .A2(keyinput58), .B1(n20965), .B2(keyinput87), 
        .ZN(n20755) );
  OAI221_X1 U23731 ( .B1(n20756), .B2(keyinput58), .C1(n20965), .C2(keyinput87), .A(n20755), .ZN(n20761) );
  AOI22_X1 U23732 ( .A1(n20759), .A2(keyinput70), .B1(keyinput115), .B2(n20758), .ZN(n20757) );
  OAI221_X1 U23733 ( .B1(n20759), .B2(keyinput70), .C1(n20758), .C2(
        keyinput115), .A(n20757), .ZN(n20760) );
  NOR4_X1 U23734 ( .A1(n20763), .A2(n20762), .A3(n20761), .A4(n20760), .ZN(
        n20764) );
  NAND4_X1 U23735 ( .A1(n20767), .A2(n20766), .A3(n20765), .A4(n20764), .ZN(
        n20957) );
  INV_X1 U23736 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n20993) );
  AOI22_X1 U23737 ( .A1(n20993), .A2(keyinput15), .B1(keyinput0), .B2(n20769), 
        .ZN(n20768) );
  OAI221_X1 U23738 ( .B1(n20993), .B2(keyinput15), .C1(n20769), .C2(keyinput0), 
        .A(n20768), .ZN(n20781) );
  AOI22_X1 U23739 ( .A1(n20772), .A2(keyinput25), .B1(keyinput89), .B2(n20771), 
        .ZN(n20770) );
  OAI221_X1 U23740 ( .B1(n20772), .B2(keyinput25), .C1(n20771), .C2(keyinput89), .A(n20770), .ZN(n20780) );
  AOI22_X1 U23741 ( .A1(n20775), .A2(keyinput124), .B1(n20774), .B2(keyinput94), .ZN(n20773) );
  OAI221_X1 U23742 ( .B1(n20775), .B2(keyinput124), .C1(n20774), .C2(
        keyinput94), .A(n20773), .ZN(n20779) );
  AOI22_X1 U23743 ( .A1(n10008), .A2(keyinput100), .B1(keyinput24), .B2(n20777), .ZN(n20776) );
  OAI221_X1 U23744 ( .B1(n10008), .B2(keyinput100), .C1(n20777), .C2(
        keyinput24), .A(n20776), .ZN(n20778) );
  NOR4_X1 U23745 ( .A1(n20781), .A2(n20780), .A3(n20779), .A4(n20778), .ZN(
        n20832) );
  AOI22_X1 U23746 ( .A1(n20987), .A2(keyinput27), .B1(keyinput2), .B2(n20783), 
        .ZN(n20782) );
  OAI221_X1 U23747 ( .B1(n20987), .B2(keyinput27), .C1(n20783), .C2(keyinput2), 
        .A(n20782), .ZN(n20795) );
  INV_X1 U23748 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n20786) );
  INV_X1 U23749 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U23750 ( .A1(n20786), .A2(keyinput43), .B1(n20785), .B2(keyinput65), 
        .ZN(n20784) );
  OAI221_X1 U23751 ( .B1(n20786), .B2(keyinput43), .C1(n20785), .C2(keyinput65), .A(n20784), .ZN(n20794) );
  AOI22_X1 U23752 ( .A1(n20789), .A2(keyinput104), .B1(n20788), .B2(keyinput64), .ZN(n20787) );
  OAI221_X1 U23753 ( .B1(n20789), .B2(keyinput104), .C1(n20788), .C2(
        keyinput64), .A(n20787), .ZN(n20793) );
  AOI22_X1 U23754 ( .A1(n20963), .A2(keyinput4), .B1(keyinput67), .B2(n20791), 
        .ZN(n20790) );
  OAI221_X1 U23755 ( .B1(n20963), .B2(keyinput4), .C1(n20791), .C2(keyinput67), 
        .A(n20790), .ZN(n20792) );
  NOR4_X1 U23756 ( .A1(n20795), .A2(n20794), .A3(n20793), .A4(n20792), .ZN(
        n20831) );
  INV_X1 U23757 ( .A(P3_LWORD_REG_2__SCAN_IN), .ZN(n20798) );
  AOI22_X1 U23758 ( .A1(n20798), .A2(keyinput51), .B1(n20797), .B2(keyinput6), 
        .ZN(n20796) );
  OAI221_X1 U23759 ( .B1(n20798), .B2(keyinput51), .C1(n20797), .C2(keyinput6), 
        .A(n20796), .ZN(n20801) );
  INV_X1 U23760 ( .A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20799) );
  XNOR2_X1 U23761 ( .A(n20799), .B(keyinput74), .ZN(n20800) );
  NOR2_X1 U23762 ( .A1(n20801), .A2(n20800), .ZN(n20813) );
  AOI22_X1 U23763 ( .A1(n20804), .A2(keyinput80), .B1(n20803), .B2(keyinput76), 
        .ZN(n20802) );
  OAI221_X1 U23764 ( .B1(n20804), .B2(keyinput80), .C1(n20803), .C2(keyinput76), .A(n20802), .ZN(n20805) );
  INV_X1 U23765 ( .A(n20805), .ZN(n20812) );
  AOI22_X1 U23766 ( .A1(n20808), .A2(keyinput86), .B1(n20807), .B2(keyinput49), 
        .ZN(n20806) );
  OAI221_X1 U23767 ( .B1(n20808), .B2(keyinput86), .C1(n20807), .C2(keyinput49), .A(n20806), .ZN(n20809) );
  INV_X1 U23768 ( .A(n20809), .ZN(n20811) );
  XNOR2_X1 U23769 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B(keyinput20), .ZN(
        n20810) );
  AND4_X1 U23770 ( .A1(n20813), .A2(n20812), .A3(n20811), .A4(n20810), .ZN(
        n20830) );
  AOI22_X1 U23771 ( .A1(n20816), .A2(keyinput48), .B1(keyinput102), .B2(n20815), .ZN(n20814) );
  OAI221_X1 U23772 ( .B1(n20816), .B2(keyinput48), .C1(n20815), .C2(
        keyinput102), .A(n20814), .ZN(n20828) );
  AOI22_X1 U23773 ( .A1(n20979), .A2(keyinput101), .B1(keyinput1), .B2(n20818), 
        .ZN(n20817) );
  OAI221_X1 U23774 ( .B1(n20979), .B2(keyinput101), .C1(n20818), .C2(keyinput1), .A(n20817), .ZN(n20827) );
  AOI22_X1 U23775 ( .A1(n20821), .A2(keyinput7), .B1(n20820), .B2(keyinput116), 
        .ZN(n20819) );
  OAI221_X1 U23776 ( .B1(n20821), .B2(keyinput7), .C1(n20820), .C2(keyinput116), .A(n20819), .ZN(n20826) );
  INV_X1 U23777 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20824) );
  INV_X1 U23778 ( .A(READY2), .ZN(n20823) );
  AOI22_X1 U23779 ( .A1(n20824), .A2(keyinput30), .B1(keyinput108), .B2(n20823), .ZN(n20822) );
  OAI221_X1 U23780 ( .B1(n20824), .B2(keyinput30), .C1(n20823), .C2(
        keyinput108), .A(n20822), .ZN(n20825) );
  NOR4_X1 U23781 ( .A1(n20828), .A2(n20827), .A3(n20826), .A4(n20825), .ZN(
        n20829) );
  NAND4_X1 U23782 ( .A1(n20832), .A2(n20831), .A3(n20830), .A4(n20829), .ZN(
        n20956) );
  AOI22_X1 U23783 ( .A1(n20835), .A2(keyinput62), .B1(n20834), .B2(keyinput91), 
        .ZN(n20833) );
  OAI221_X1 U23784 ( .B1(n20835), .B2(keyinput62), .C1(n20834), .C2(keyinput91), .A(n20833), .ZN(n20839) );
  XNOR2_X1 U23785 ( .A(n20836), .B(keyinput3), .ZN(n20838) );
  XOR2_X1 U23786 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B(keyinput117), .Z(
        n20837) );
  OR3_X1 U23787 ( .A1(n20839), .A2(n20838), .A3(n20837), .ZN(n20848) );
  AOI22_X1 U23788 ( .A1(n20842), .A2(keyinput71), .B1(keyinput5), .B2(n20841), 
        .ZN(n20840) );
  OAI221_X1 U23789 ( .B1(n20842), .B2(keyinput71), .C1(n20841), .C2(keyinput5), 
        .A(n20840), .ZN(n20847) );
  AOI22_X1 U23790 ( .A1(n20845), .A2(keyinput42), .B1(n20844), .B2(keyinput44), 
        .ZN(n20843) );
  OAI221_X1 U23791 ( .B1(n20845), .B2(keyinput42), .C1(n20844), .C2(keyinput44), .A(n20843), .ZN(n20846) );
  NOR3_X1 U23792 ( .A1(n20848), .A2(n20847), .A3(n20846), .ZN(n20892) );
  AOI22_X1 U23793 ( .A1(n20851), .A2(keyinput63), .B1(keyinput93), .B2(n20850), 
        .ZN(n20849) );
  OAI221_X1 U23794 ( .B1(n20851), .B2(keyinput63), .C1(n20850), .C2(keyinput93), .A(n20849), .ZN(n20860) );
  INV_X1 U23795 ( .A(P3_LWORD_REG_13__SCAN_IN), .ZN(n20853) );
  AOI22_X1 U23796 ( .A1(n20854), .A2(keyinput78), .B1(keyinput18), .B2(n20853), 
        .ZN(n20852) );
  OAI221_X1 U23797 ( .B1(n20854), .B2(keyinput78), .C1(n20853), .C2(keyinput18), .A(n20852), .ZN(n20859) );
  AOI22_X1 U23798 ( .A1(n20984), .A2(keyinput17), .B1(n20960), .B2(keyinput106), .ZN(n20855) );
  OAI221_X1 U23799 ( .B1(n20984), .B2(keyinput17), .C1(n20960), .C2(
        keyinput106), .A(n20855), .ZN(n20858) );
  AOI22_X1 U23800 ( .A1(n20986), .A2(keyinput46), .B1(n10522), .B2(keyinput29), 
        .ZN(n20856) );
  OAI221_X1 U23801 ( .B1(n20986), .B2(keyinput46), .C1(n10522), .C2(keyinput29), .A(n20856), .ZN(n20857) );
  NOR4_X1 U23802 ( .A1(n20860), .A2(n20859), .A3(n20858), .A4(n20857), .ZN(
        n20891) );
  AOI22_X1 U23803 ( .A1(n20863), .A2(keyinput112), .B1(n20862), .B2(keyinput8), 
        .ZN(n20861) );
  OAI221_X1 U23804 ( .B1(n20863), .B2(keyinput112), .C1(n20862), .C2(keyinput8), .A(n20861), .ZN(n20875) );
  AOI22_X1 U23805 ( .A1(n14095), .A2(keyinput110), .B1(n20865), .B2(keyinput38), .ZN(n20864) );
  OAI221_X1 U23806 ( .B1(n14095), .B2(keyinput110), .C1(n20865), .C2(
        keyinput38), .A(n20864), .ZN(n20874) );
  INV_X1 U23807 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20867) );
  AOI22_X1 U23808 ( .A1(n20868), .A2(keyinput81), .B1(keyinput59), .B2(n20867), 
        .ZN(n20866) );
  OAI221_X1 U23809 ( .B1(n20868), .B2(keyinput81), .C1(n20867), .C2(keyinput59), .A(n20866), .ZN(n20873) );
  AOI22_X1 U23810 ( .A1(n20871), .A2(keyinput47), .B1(keyinput52), .B2(n20870), 
        .ZN(n20869) );
  OAI221_X1 U23811 ( .B1(n20871), .B2(keyinput47), .C1(n20870), .C2(keyinput52), .A(n20869), .ZN(n20872) );
  NOR4_X1 U23812 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20890) );
  AOI22_X1 U23813 ( .A1(n10891), .A2(keyinput11), .B1(keyinput105), .B2(n20962), .ZN(n20876) );
  OAI221_X1 U23814 ( .B1(n10891), .B2(keyinput11), .C1(n20962), .C2(
        keyinput105), .A(n20876), .ZN(n20888) );
  INV_X1 U23815 ( .A(DATAI_18_), .ZN(n20878) );
  AOI22_X1 U23816 ( .A1(n20879), .A2(keyinput118), .B1(n20878), .B2(keyinput57), .ZN(n20877) );
  OAI221_X1 U23817 ( .B1(n20879), .B2(keyinput118), .C1(n20878), .C2(
        keyinput57), .A(n20877), .ZN(n20887) );
  AOI22_X1 U23818 ( .A1(n20881), .A2(keyinput16), .B1(keyinput72), .B2(n20983), 
        .ZN(n20880) );
  OAI221_X1 U23819 ( .B1(n20881), .B2(keyinput16), .C1(n20983), .C2(keyinput72), .A(n20880), .ZN(n20886) );
  AOI22_X1 U23820 ( .A1(n20884), .A2(keyinput109), .B1(n20883), .B2(keyinput22), .ZN(n20882) );
  OAI221_X1 U23821 ( .B1(n20884), .B2(keyinput109), .C1(n20883), .C2(
        keyinput22), .A(n20882), .ZN(n20885) );
  NOR4_X1 U23822 ( .A1(n20888), .A2(n20887), .A3(n20886), .A4(n20885), .ZN(
        n20889) );
  NAND4_X1 U23823 ( .A1(n20892), .A2(n20891), .A3(n20890), .A4(n20889), .ZN(
        n20955) );
  AOI22_X1 U23824 ( .A1(n20895), .A2(keyinput34), .B1(keyinput127), .B2(n20894), .ZN(n20893) );
  OAI221_X1 U23825 ( .B1(n20895), .B2(keyinput34), .C1(n20894), .C2(
        keyinput127), .A(n20893), .ZN(n20908) );
  AOI22_X1 U23826 ( .A1(n20898), .A2(keyinput50), .B1(n20897), .B2(keyinput13), 
        .ZN(n20896) );
  OAI221_X1 U23827 ( .B1(n20898), .B2(keyinput50), .C1(n20897), .C2(keyinput13), .A(n20896), .ZN(n20907) );
  INV_X1 U23828 ( .A(DATAI_1_), .ZN(n20900) );
  AOI22_X1 U23829 ( .A1(n20901), .A2(keyinput75), .B1(keyinput125), .B2(n20900), .ZN(n20899) );
  OAI221_X1 U23830 ( .B1(n20901), .B2(keyinput75), .C1(n20900), .C2(
        keyinput125), .A(n20899), .ZN(n20906) );
  INV_X1 U23831 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n20902) );
  XOR2_X1 U23832 ( .A(n20902), .B(keyinput33), .Z(n20904) );
  XNOR2_X1 U23833 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B(keyinput69), .ZN(
        n20903) );
  NAND2_X1 U23834 ( .A1(n20904), .A2(n20903), .ZN(n20905) );
  NOR4_X1 U23835 ( .A1(n20908), .A2(n20907), .A3(n20906), .A4(n20905), .ZN(
        n20953) );
  INV_X1 U23836 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n20911) );
  AOI22_X1 U23837 ( .A1(n20911), .A2(keyinput53), .B1(n20910), .B2(keyinput119), .ZN(n20909) );
  OAI221_X1 U23838 ( .B1(n20911), .B2(keyinput53), .C1(n20910), .C2(
        keyinput119), .A(n20909), .ZN(n20915) );
  XNOR2_X1 U23839 ( .A(n20912), .B(keyinput14), .ZN(n20914) );
  XOR2_X1 U23840 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B(keyinput121), .Z(
        n20913) );
  OR3_X1 U23841 ( .A1(n20915), .A2(n20914), .A3(n20913), .ZN(n20921) );
  AOI22_X1 U23842 ( .A1(n20961), .A2(keyinput92), .B1(n10012), .B2(keyinput123), .ZN(n20916) );
  OAI221_X1 U23843 ( .B1(n20961), .B2(keyinput92), .C1(n10012), .C2(
        keyinput123), .A(n20916), .ZN(n20920) );
  AOI22_X1 U23844 ( .A1(n20918), .A2(keyinput79), .B1(n20998), .B2(keyinput82), 
        .ZN(n20917) );
  OAI221_X1 U23845 ( .B1(n20918), .B2(keyinput79), .C1(n20998), .C2(keyinput82), .A(n20917), .ZN(n20919) );
  NOR3_X1 U23846 ( .A1(n20921), .A2(n20920), .A3(n20919), .ZN(n20952) );
  AOI22_X1 U23847 ( .A1(n20923), .A2(keyinput39), .B1(n20969), .B2(keyinput26), 
        .ZN(n20922) );
  OAI221_X1 U23848 ( .B1(n20923), .B2(keyinput39), .C1(n20969), .C2(keyinput26), .A(n20922), .ZN(n20934) );
  AOI22_X1 U23849 ( .A1(n20925), .A2(keyinput66), .B1(keyinput90), .B2(n12626), 
        .ZN(n20924) );
  OAI221_X1 U23850 ( .B1(n20925), .B2(keyinput66), .C1(n12626), .C2(keyinput90), .A(n20924), .ZN(n20933) );
  XOR2_X1 U23851 ( .A(n20926), .B(keyinput95), .Z(n20929) );
  XNOR2_X1 U23852 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B(keyinput12), .ZN(
        n20928) );
  XNOR2_X1 U23853 ( .A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B(keyinput40), .ZN(
        n20927) );
  NAND3_X1 U23854 ( .A1(n20929), .A2(n20928), .A3(n20927), .ZN(n20932) );
  XNOR2_X1 U23855 ( .A(n20930), .B(keyinput103), .ZN(n20931) );
  NOR4_X1 U23856 ( .A1(n20934), .A2(n20933), .A3(n20932), .A4(n20931), .ZN(
        n20951) );
  AOI22_X1 U23857 ( .A1(n20937), .A2(keyinput55), .B1(keyinput60), .B2(n20936), 
        .ZN(n20935) );
  OAI221_X1 U23858 ( .B1(n20937), .B2(keyinput55), .C1(n20936), .C2(keyinput60), .A(n20935), .ZN(n20949) );
  AOI22_X1 U23859 ( .A1(n20940), .A2(keyinput88), .B1(n20939), .B2(keyinput114), .ZN(n20938) );
  OAI221_X1 U23860 ( .B1(n20940), .B2(keyinput88), .C1(n20939), .C2(
        keyinput114), .A(n20938), .ZN(n20948) );
  AOI22_X1 U23861 ( .A1(n20943), .A2(keyinput36), .B1(keyinput45), .B2(n20942), 
        .ZN(n20941) );
  OAI221_X1 U23862 ( .B1(n20943), .B2(keyinput36), .C1(n20942), .C2(keyinput45), .A(n20941), .ZN(n20947) );
  AOI22_X1 U23863 ( .A1(n20945), .A2(keyinput23), .B1(keyinput113), .B2(n9992), 
        .ZN(n20944) );
  OAI221_X1 U23864 ( .B1(n20945), .B2(keyinput23), .C1(n9992), .C2(keyinput113), .A(n20944), .ZN(n20946) );
  NOR4_X1 U23865 ( .A1(n20949), .A2(n20948), .A3(n20947), .A4(n20946), .ZN(
        n20950) );
  NAND4_X1 U23866 ( .A1(n20953), .A2(n20952), .A3(n20951), .A4(n20950), .ZN(
        n20954) );
  NOR4_X1 U23867 ( .A1(n20957), .A2(n20956), .A3(n20955), .A4(n20954), .ZN(
        n20958) );
  XNOR2_X1 U23868 ( .A(n20959), .B(n20958), .ZN(n21025) );
  NOR4_X1 U23869 ( .A1(n20961), .A2(n20960), .A3(
        P1_INSTQUEUE_REG_11__2__SCAN_IN), .A4(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20968) );
  NAND4_X1 U23870 ( .A1(P1_EBX_REG_1__SCAN_IN), .A2(n20964), .A3(n20963), .A4(
        n20962), .ZN(n20966) );
  NOR3_X1 U23871 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20966), .A3(
        P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n20967) );
  NAND4_X1 U23872 ( .A1(n20968), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .A4(n20967), .ZN(n20973) );
  NAND4_X1 U23873 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n20971), .A3(
        n20970), .A4(n20969), .ZN(n20972) );
  NOR2_X1 U23874 ( .A1(n20973), .A2(n20972), .ZN(n21023) );
  NAND4_X1 U23875 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n20975), .A4(n20974), .ZN(
        n20982) );
  NOR3_X1 U23876 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_3__7__SCAN_IN), .A3(n20976), .ZN(n20977) );
  NAND3_X1 U23877 ( .A1(n20977), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A3(
        P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20981) );
  NAND4_X1 U23878 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12626), .A3(
        n20979), .A4(n20978), .ZN(n20980) );
  NOR3_X1 U23879 ( .A1(n20982), .A2(n20981), .A3(n20980), .ZN(n21022) );
  NOR4_X1 U23880 ( .A1(P1_EAX_REG_16__SCAN_IN), .A2(DATAI_18_), .A3(n20984), 
        .A4(n20983), .ZN(n20985) );
  NAND3_X1 U23881 ( .A1(BUF1_REG_30__SCAN_IN), .A2(BUF1_REG_26__SCAN_IN), .A3(
        n20985), .ZN(n20997) );
  NAND4_X1 U23882 ( .A1(READY2), .A2(P3_ADDRESS_REG_13__SCAN_IN), .A3(n20987), 
        .A4(n20986), .ZN(n20988) );
  NOR3_X1 U23883 ( .A1(DATAI_23_), .A2(BUF1_REG_20__SCAN_IN), .A3(n20988), 
        .ZN(n20995) );
  NAND4_X1 U23884 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_15__6__SCAN_IN), .A3(P3_REIP_REG_11__SCAN_IN), .A4(
        P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n20992) );
  NAND4_X1 U23885 ( .A1(P3_DATAO_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_UWORD_REG_4__SCAN_IN), .A4(
        P3_UWORD_REG_2__SCAN_IN), .ZN(n20991) );
  NAND4_X1 U23886 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_5__0__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n20990) );
  NAND4_X1 U23887 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A3(P3_REIP_REG_0__SCAN_IN), .A4(
        P3_EBX_REG_15__SCAN_IN), .ZN(n20989) );
  NOR4_X1 U23888 ( .A1(n20992), .A2(n20991), .A3(n20990), .A4(n20989), .ZN(
        n20994) );
  NAND4_X1 U23889 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20995), .A3(n20994), 
        .A4(n20993), .ZN(n20996) );
  NOR4_X1 U23890 ( .A1(n20999), .A2(n20998), .A3(n20997), .A4(n20996), .ZN(
        n21021) );
  NOR4_X1 U23891 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_DATAO_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        DATAI_1_), .ZN(n21003) );
  NOR4_X1 U23892 ( .A1(P3_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_11__SCAN_IN), .A3(READY22_REG_SCAN_IN), .A4(
        P3_W_R_N_REG_SCAN_IN), .ZN(n21002) );
  NOR4_X1 U23893 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_EAX_REG_26__SCAN_IN), .A3(P2_EAX_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_8__SCAN_IN), .ZN(n21001) );
  NOR4_X1 U23894 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(P1_EBX_REG_15__SCAN_IN), 
        .A3(P1_UWORD_REG_12__SCAN_IN), .A4(P2_UWORD_REG_5__SCAN_IN), .ZN(
        n21000) );
  NAND4_X1 U23895 ( .A1(n21003), .A2(n21002), .A3(n21001), .A4(n21000), .ZN(
        n21019) );
  NAND4_X1 U23896 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P1_UWORD_REG_2__SCAN_IN), 
        .A3(P1_LWORD_REG_4__SCAN_IN), .A4(P2_UWORD_REG_7__SCAN_IN), .ZN(n21007) );
  NAND4_X1 U23897 ( .A1(P3_ADDRESS_REG_25__SCAN_IN), .A2(
        P3_UWORD_REG_13__SCAN_IN), .A3(P3_LWORD_REG_5__SCAN_IN), .A4(
        P2_DATAO_REG_0__SCAN_IN), .ZN(n21006) );
  NAND4_X1 U23898 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_3__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_READREQUEST_REG_SCAN_IN), .ZN(n21005) );
  NAND4_X1 U23899 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(P2_REIP_REG_15__SCAN_IN), 
        .A3(P2_REIP_REG_16__SCAN_IN), .A4(P2_EAX_REG_13__SCAN_IN), .ZN(n21004)
         );
  OR4_X1 U23900 ( .A1(n21007), .A2(n21006), .A3(n21005), .A4(n21004), .ZN(
        n21018) );
  NOR4_X1 U23901 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .A3(BUF2_REG_17__SCAN_IN), .A4(
        BUF2_REG_20__SCAN_IN), .ZN(n21011) );
  NOR4_X1 U23902 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_DATAO_REG_22__SCAN_IN), .A3(P1_DATAO_REG_28__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n21010) );
  NOR4_X1 U23903 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(
        P2_EBX_REG_22__SCAN_IN), .A3(P2_REIP_REG_30__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21009) );
  NOR4_X1 U23904 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_8__6__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21008) );
  NAND4_X1 U23905 ( .A1(n21011), .A2(n21010), .A3(n21009), .A4(n21008), .ZN(
        n21017) );
  NOR4_X1 U23906 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_11__0__SCAN_IN), .A3(P3_INSTQUEUE_REG_10__2__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n21015) );
  NOR4_X1 U23907 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_LWORD_REG_2__SCAN_IN), .A3(P3_LWORD_REG_13__SCAN_IN), .A4(
        P3_DATAO_REG_13__SCAN_IN), .ZN(n21014) );
  NOR4_X1 U23908 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A3(P2_DATAO_REG_13__SCAN_IN), .A4(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n21013) );
  NOR4_X1 U23909 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_6__5__SCAN_IN), .A3(P3_INSTQUEUE_REG_12__6__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n21012) );
  NAND4_X1 U23910 ( .A1(n21015), .A2(n21014), .A3(n21013), .A4(n21012), .ZN(
        n21016) );
  NOR4_X1 U23911 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21020) );
  NAND4_X1 U23912 ( .A1(n21023), .A2(n21022), .A3(n21021), .A4(n21020), .ZN(
        n21024) );
  XNOR2_X1 U23913 ( .A(n21025), .B(n21024), .ZN(P1_U2860) );
  NAND2_X1 U12610 ( .A1(n10034), .A2(n10032), .ZN(n10766) );
  BUF_X1 U11180 ( .A(n12265), .Z(n9723) );
  BUF_X2 U11168 ( .A(n10369), .Z(n9750) );
  CLKBUF_X1 U11208 ( .A(n12049), .Z(n12032) );
  CLKBUF_X1 U11216 ( .A(n12470), .Z(n9737) );
  CLKBUF_X1 U11230 ( .A(n13438), .Z(n14335) );
  CLKBUF_X1 U11254 ( .A(n9741), .Z(n11210) );
  CLKBUF_X1 U11272 ( .A(n12191), .Z(n17414) );
  AND2_X1 U11509 ( .A1(n13872), .A2(n9963), .ZN(n14230) );
  CLKBUF_X1 U11619 ( .A(n15347), .Z(n16408) );
  CLKBUF_X1 U12191 ( .A(n16683), .Z(n9740) );
  CLKBUF_X1 U12431 ( .A(n15667), .Z(n16482) );
  CLKBUF_X1 U12443 ( .A(n14740), .Z(n14741) );
  CLKBUF_X1 U12593 ( .A(n12740), .Z(n12762) );
endmodule

