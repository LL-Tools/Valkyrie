

module b17_C_gen_AntiSAT_k_256_7 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, 
        keyinput_f65, keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, 
        keyinput_f70, keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, 
        keyinput_f75, keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, 
        keyinput_f80, keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, 
        keyinput_f85, keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, 
        keyinput_f90, keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, 
        keyinput_f95, keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, 
        keyinput_f100, keyinput_f101, keyinput_f102, keyinput_f103, 
        keyinput_f104, keyinput_f105, keyinput_f106, keyinput_f107, 
        keyinput_f108, keyinput_f109, keyinput_f110, keyinput_f111, 
        keyinput_f112, keyinput_f113, keyinput_f114, keyinput_f115, 
        keyinput_f116, keyinput_f117, keyinput_f118, keyinput_f119, 
        keyinput_f120, keyinput_f121, keyinput_f122, keyinput_f123, 
        keyinput_f124, keyinput_f125, keyinput_f126, keyinput_f127, 
        keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, 
        keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, 
        keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, 
        keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, 
        keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, 
        keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, 
        keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, 
        keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, 
        keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, 
        keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, 
        keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, 
        keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, 
        keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63, keyinput_g64, 
        keyinput_g65, keyinput_g66, keyinput_g67, keyinput_g68, keyinput_g69, 
        keyinput_g70, keyinput_g71, keyinput_g72, keyinput_g73, keyinput_g74, 
        keyinput_g75, keyinput_g76, keyinput_g77, keyinput_g78, keyinput_g79, 
        keyinput_g80, keyinput_g81, keyinput_g82, keyinput_g83, keyinput_g84, 
        keyinput_g85, keyinput_g86, keyinput_g87, keyinput_g88, keyinput_g89, 
        keyinput_g90, keyinput_g91, keyinput_g92, keyinput_g93, keyinput_g94, 
        keyinput_g95, keyinput_g96, keyinput_g97, keyinput_g98, keyinput_g99, 
        keyinput_g100, keyinput_g101, keyinput_g102, keyinput_g103, 
        keyinput_g104, keyinput_g105, keyinput_g106, keyinput_g107, 
        keyinput_g108, keyinput_g109, keyinput_g110, keyinput_g111, 
        keyinput_g112, keyinput_g113, keyinput_g114, keyinput_g115, 
        keyinput_g116, keyinput_g117, keyinput_g118, keyinput_g119, 
        keyinput_g120, keyinput_g121, keyinput_g122, keyinput_g123, 
        keyinput_g124, keyinput_g125, keyinput_g126, keyinput_g127, U355, U356, 
        U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, 
        U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, 
        U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, 
        U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, 
        U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, 
        U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, 
        U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, 
        U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, 
        P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, 
        P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, 
        P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, 
        P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, 
        P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, 
        P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, 
        P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, 
        P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, 
        P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, 
        P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, 
        P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, 
        P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, 
        P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, 
        P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, 
        P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, 
        P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, 
        P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, 
        P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, 
        P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, 
        P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, 
        P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, 
        P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, 
        P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, 
        P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, 
        P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, 
        P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, 
        P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, 
        P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, 
        P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, 
        P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, 
        P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, 
        P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, 
        P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, 
        P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, 
        P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, 
        P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, 
        P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, 
        P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, 
        P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, 
        P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, 
        P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, 
        P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, 
        P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, 
        P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, 
        P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, 
        P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, 
        P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, 
        P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, 
        P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, 
        P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, 
        P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, 
        P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, 
        P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, 
        P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, 
        P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, 
        P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, 
        P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, 
        P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, 
        P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, 
        P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, 
        P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, 
        P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, 
        P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, 
        P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, 
        P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, 
        P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, 
        P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, 
        P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, 
        P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, 
        P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, 
        P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, 
        P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, 
        P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, 
        P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, 
        P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, 
        P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, 
        P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, 
        P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, 
        P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, 
        P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, 
        P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, 
        P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, 
        P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, 
        P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, 
        P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, 
        P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, 
        P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, 
        P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, 
        P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, 
        P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, 
        P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, 
        P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, 
        P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, 
        P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, 
        P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, 
        P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, 
        P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, 
        P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, 
        P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, 
        P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, 
        P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, 
        P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, 
        P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, 
        P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, 
        P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, 
        P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, 
        P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, 
        P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, 
        P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, 
        P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, 
        P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, 
        P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, 
        P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, 
        P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, 
        P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, 
        P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, 
        P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, 
        P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, 
        P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, 
        P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, 
        P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, 
        P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, 
        P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, 
        P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, 
        P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, 
        P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, 
        P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, 
        P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, 
        P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, 
        P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, 
        P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, 
        P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, 
        P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, 
        P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, 
        P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, 
        P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, 
        P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, 
        P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, 
        P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, 
        P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, 
        P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, 
        P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, 
        P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, 
        P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, 
        P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, 
        P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, 
        P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, 
        P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, 
        P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, 
        P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, 
        P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, 
        P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, 
        P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, 
        P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, 
        P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, 
        P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, 
        P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, 
        P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, 
        P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, 
        P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, 
        P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, 
        P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, 
        P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, 
        P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, 
        P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, 
        P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, 
        P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, 
        P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, 
        P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, 
        P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, 
        P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, 
        P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, 
        P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, 
        P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, 
        P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, 
        P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, 
        P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, 
        P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, 
        P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, 
        P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9811, n9812, n9814, n9815, n9816, n9817, n9819, n9820, n9821, n9822,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
         n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148,
         n17149, n17150, n17151, n17152, n17153, n17154, n17155, n17156,
         n17157, n17158, n17159, n17160, n17161, n17162, n17163, n17164,
         n17165, n17166, n17167, n17168, n17169, n17170, n17171, n17172,
         n17173, n17174, n17175, n17176, n17177, n17178, n17179, n17180,
         n17181, n17182, n17183, n17184, n17185, n17186, n17187, n17188,
         n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
         n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204,
         n17205, n17206, n17207, n17208, n17209, n17210, n17211, n17212,
         n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220,
         n17221, n17222, n17223, n17224, n17225, n17226, n17227, n17228,
         n17229, n17230, n17231, n17232, n17233, n17234, n17235, n17236,
         n17237, n17238, n17239, n17240, n17241, n17242, n17243, n17244,
         n17245, n17246, n17247, n17248, n17249, n17250, n17251, n17252,
         n17253, n17254, n17255, n17256, n17257, n17258, n17259, n17260,
         n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268,
         n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
         n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284,
         n17285, n17286, n17287, n17288, n17289, n17290, n17291, n17292,
         n17293, n17294, n17295, n17296, n17297, n17298, n17299, n17300,
         n17301, n17302, n17303, n17304, n17305, n17306, n17307, n17308,
         n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
         n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324,
         n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332,
         n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340,
         n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
         n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356,
         n17357, n17358, n17359, n17360, n17361, n17362, n17363, n17364,
         n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
         n17373, n17374, n17375, n17376, n17377, n17378, n17379, n17380,
         n17381, n17382, n17383, n17384, n17385, n17386, n17387, n17388,
         n17389, n17390, n17391, n17392, n17393, n17394, n17395, n17396,
         n17397, n17398, n17399, n17400, n17401, n17402, n17403, n17404,
         n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412,
         n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420,
         n17421, n17422, n17423, n17424, n17425, n17426, n17427, n17428,
         n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
         n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444,
         n17445, n17446, n17447, n17448, n17449, n17450, n17451, n17452,
         n17453, n17454, n17455, n17456, n17457, n17458, n17459, n17460,
         n17461, n17462, n17463, n17464, n17465, n17466, n17467, n17468,
         n17469, n17470, n17471, n17472, n17473, n17474, n17475, n17476,
         n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484,
         n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492,
         n17493, n17494, n17495, n17496, n17497, n17498, n17499, n17500,
         n17501, n17502, n17503, n17504, n17505, n17506, n17507, n17508,
         n17509, n17510, n17511, n17512, n17513, n17514, n17515, n17516,
         n17517, n17518, n17519, n17520, n17521, n17522, n17523, n17524,
         n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
         n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540,
         n17541, n17542, n17543, n17544, n17545, n17546, n17547, n17548,
         n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556,
         n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564,
         n17565, n17566, n17567, n17568, n17569, n17570, n17571, n17572,
         n17573, n17574, n17575, n17576, n17577, n17578, n17579, n17580,
         n17581, n17582, n17583, n17584, n17585, n17586, n17587, n17588,
         n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596,
         n17597, n17598, n17599, n17600, n17601, n17602, n17603, n17604,
         n17605, n17606, n17607, n17608, n17609, n17610, n17611, n17612,
         n17613, n17614, n17615, n17616, n17617, n17618, n17619, n17620,
         n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628,
         n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636,
         n17637, n17638, n17639, n17640, n17641, n17642, n17643, n17644,
         n17645, n17646, n17647, n17648, n17649, n17650, n17651, n17652,
         n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
         n17661, n17662, n17663, n17664, n17665, n17666, n17667, n17668,
         n17669, n17670, n17671, n17672, n17673, n17674, n17675, n17676,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17714, n17715, n17716,
         n17717, n17718, n17719, n17720, n17721, n17722, n17723, n17724,
         n17725, n17726, n17727, n17728, n17729, n17730, n17731, n17732,
         n17733, n17734, n17735, n17736, n17737, n17738, n17739, n17740,
         n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
         n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756,
         n17757, n17758, n17759, n17760, n17761, n17762, n17763, n17764,
         n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772,
         n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780,
         n17781, n17782, n17783, n17784, n17785, n17786, n17787, n17788,
         n17789, n17790, n17791, n17792, n17793, n17794, n17795, n17796,
         n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804,
         n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
         n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820,
         n17821, n17822, n17823, n17824, n17825, n17826, n17827, n17828,
         n17829, n17830, n17831, n17832, n17833, n17834, n17835, n17836,
         n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844,
         n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
         n17853, n17854, n17855, n17856, n17857, n17858, n17859, n17860,
         n17861, n17862, n17863, n17864, n17865, n17866, n17867, n17868,
         n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
         n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884,
         n17885, n17886, n17887, n17888, n17889, n17890, n17891, n17892,
         n17893, n17894, n17895, n17896, n17897, n17898, n17899, n17900,
         n17901, n17902, n17903, n17904, n17905, n17906, n17907, n17908,
         n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916,
         n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924,
         n17925, n17926, n17927, n17928, n17929, n17930, n17931, n17932,
         n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
         n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948,
         n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
         n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964,
         n17965, n17966, n17967, n17968, n17969, n17970, n17971, n17972,
         n17973, n17974, n17975, n17976, n17977, n17978, n17979, n17980,
         n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988,
         n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996,
         n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
         n18005, n18006, n18007, n18008, n18009, n18010, n18011, n18012,
         n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020,
         n18021, n18022, n18023, n18024, n18025, n18026, n18027, n18028,
         n18029, n18030, n18031, n18032, n18033, n18034, n18035, n18036,
         n18037, n18038, n18039, n18040, n18041, n18042, n18043, n18044,
         n18045, n18046, n18047, n18048, n18049, n18050, n18051, n18052,
         n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060,
         n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068,
         n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18076,
         n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
         n18085, n18086, n18087, n18088, n18089, n18090, n18091, n18092,
         n18093, n18094, n18095, n18096, n18097, n18098, n18099, n18100,
         n18101, n18102, n18103, n18104, n18105, n18106, n18107, n18108,
         n18109, n18110, n18111, n18112, n18113, n18114, n18115, n18116,
         n18117, n18118, n18119, n18120, n18121, n18122, n18123, n18124,
         n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132,
         n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
         n18141, n18142, n18143, n18144, n18145, n18146, n18147, n18148,
         n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
         n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164,
         n18165, n18166, n18167, n18168, n18169, n18170, n18171, n18172,
         n18173, n18174, n18175, n18176, n18177, n18178, n18179, n18180,
         n18181, n18182, n18183, n18184, n18185, n18186, n18187, n18188,
         n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
         n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204,
         n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212,
         n18213, n18214, n18215, n18216, n18217, n18218, n18219, n18220,
         n18221, n18222, n18223, n18224, n18225, n18226, n18227, n18228,
         n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236,
         n18237, n18238, n18239, n18240, n18241, n18242, n18243, n18244,
         n18245, n18246, n18247, n18248, n18249, n18250, n18251, n18252,
         n18253, n18254, n18255, n18256, n18257, n18258, n18259, n18260,
         n18261, n18262, n18263, n18264, n18265, n18266, n18267, n18268,
         n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
         n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284,
         n18285, n18286, n18287, n18288, n18289, n18290, n18291, n18292,
         n18293, n18294, n18295, n18296, n18297, n18298, n18299, n18300,
         n18301, n18302, n18303, n18304, n18305, n18306, n18307, n18308,
         n18309, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18317, n18318, n18319, n18320, n18321, n18322, n18323, n18324,
         n18325, n18326, n18327, n18328, n18329, n18330, n18331, n18332,
         n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340,
         n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348,
         n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356,
         n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
         n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372,
         n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380,
         n18381, n18382, n18383, n18384, n18385, n18386, n18387, n18388,
         n18389, n18390, n18391, n18392, n18393, n18394, n18395, n18396,
         n18397, n18398, n18399, n18400, n18401, n18402, n18403, n18404,
         n18405, n18406, n18407, n18408, n18409, n18410, n18411, n18412,
         n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420,
         n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428,
         n18429, n18430, n18431, n18432, n18433, n18434, n18435, n18436,
         n18437, n18438, n18439, n18440, n18441, n18442, n18443, n18444,
         n18445, n18446, n18447, n18448, n18449, n18450, n18451, n18452,
         n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460,
         n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468,
         n18469, n18470, n18471, n18472, n18473, n18474, n18475, n18476,
         n18477, n18478, n18479, n18480, n18481, n18482, n18483, n18484,
         n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492,
         n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500,
         n18501, n18502, n18503, n18504, n18505, n18506, n18507, n18508,
         n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
         n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524,
         n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532,
         n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540,
         n18541, n18542, n18543, n18544, n18545, n18546, n18547, n18548,
         n18549, n18550, n18551, n18552, n18553, n18554, n18555, n18556,
         n18557, n18558, n18559, n18560, n18561, n18562, n18563, n18564,
         n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
         n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580,
         n18581, n18582, n18583, n18584, n18585, n18586, n18587, n18588,
         n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
         n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604,
         n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612,
         n18613, n18614, n18615, n18616, n18617, n18618, n18619, n18620,
         n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
         n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636,
         n18637, n18638, n18639, n18640, n18641, n18642, n18643, n18644,
         n18645, n18646, n18647, n18648, n18649, n18650, n18651, n18652,
         n18653, n18654, n18655, n18656, n18657, n18658, n18659, n18660,
         n18661, n18662, n18663, n18664, n18665, n18666, n18667, n18668,
         n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676,
         n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684,
         n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692,
         n18693, n18694, n18695, n18696, n18697, n18698, n18699, n18700,
         n18701, n18702, n18703, n18704, n18705, n18706, n18707, n18708,
         n18709, n18710, n18711, n18712, n18713, n18714, n18715, n18716,
         n18717, n18718, n18719, n18720, n18721, n18722, n18723, n18724,
         n18725, n18726, n18727, n18728, n18729, n18730, n18731, n18732,
         n18733, n18734, n18735, n18736, n18737, n18738, n18739, n18740,
         n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748,
         n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756,
         n18757, n18758, n18759, n18760, n18761, n18762, n18763, n18764,
         n18765, n18766, n18767, n18768, n18769, n18770, n18771, n18772,
         n18773, n18774, n18775, n18776, n18777, n18778, n18779, n18780,
         n18781, n18782, n18783, n18784, n18785, n18786, n18787, n18788,
         n18789, n18790, n18791, n18792, n18793, n18794, n18795, n18796,
         n18797, n18798, n18799, n18800, n18801, n18802, n18803, n18804,
         n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
         n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820,
         n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828,
         n18829, n18830, n18831, n18832, n18833, n18834, n18835, n18836,
         n18837, n18838, n18839, n18840, n18841, n18842, n18843, n18844,
         n18845, n18846, n18847, n18848, n18849, n18850, n18851, n18852,
         n18853, n18854, n18855, n18856, n18857, n18858, n18859, n18860,
         n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
         n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876,
         n18877, n18878, n18879, n18880, n18881, n18882, n18883, n18884,
         n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892,
         n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900,
         n18901, n18902, n18903, n18904, n18905, n18906, n18907, n18908,
         n18909, n18910, n18911, n18912, n18913, n18914, n18915, n18916,
         n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
         n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932,
         n18933, n18934, n18935, n18936, n18937, n18938, n18939, n18940,
         n18941, n18942, n18943, n18944, n18945, n18946, n18947, n18948,
         n18949, n18950, n18951, n18952, n18953, n18954, n18955, n18956,
         n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964,
         n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972,
         n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
         n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988,
         n18989, n18990, n18991, n18992, n18993, n18994, n18995, n18996,
         n18997, n18998, n18999, n19000, n19001, n19002, n19003, n19004,
         n19005, n19006, n19007, n19008, n19009, n19010, n19011, n19012,
         n19013, n19014, n19015, n19016, n19017, n19018, n19019, n19020,
         n19021, n19022, n19023, n19024, n19025, n19026, n19027, n19028,
         n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
         n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044,
         n19045, n19046, n19047, n19048, n19049, n19050, n19051, n19052,
         n19053, n19054, n19055, n19056, n19057, n19058, n19059, n19060,
         n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
         n19069, n19070, n19071, n19072, n19073, n19074, n19075, n19076,
         n19077, n19078, n19079, n19080, n19081, n19082, n19083, n19084,
         n19085, n19086, n19087, n19088, n19089, n19090, n19091, n19092,
         n19093, n19094, n19095, n19096, n19097, n19098, n19099, n19100,
         n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108,
         n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116,
         n19117, n19118, n19119, n19120, n19121, n19122, n19123, n19124,
         n19125, n19126, n19127, n19128, n19129, n19130, n19131, n19132,
         n19133, n19134, n19135, n19136, n19137, n19138, n19139, n19140,
         n19141, n19142, n19143, n19144, n19145, n19146, n19147, n19148,
         n19149, n19150, n19151, n19152, n19153, n19154, n19155, n19156,
         n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
         n19165, n19166, n19167, n19168, n19169, n19170, n19171, n19172,
         n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180,
         n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188,
         n19189, n19190, n19191, n19192, n19193, n19194, n19195, n19196,
         n19197, n19198, n19199, n19200, n19201, n19202, n19203, n19204,
         n19205, n19206, n19207, n19208, n19209, n19210, n19211, n19212,
         n19213, n19214, n19215, n19216, n19217, n19218, n19219, n19220,
         n19221, n19222, n19223, n19224, n19225, n19226, n19227, n19228,
         n19229, n19230, n19231, n19232, n19233, n19234, n19235, n19236,
         n19237, n19238, n19239, n19240, n19241, n19242, n19243, n19244,
         n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260,
         n19261, n19262, n19263, n19264, n19265, n19266, n19267, n19268,
         n19269, n19270, n19271, n19272, n19273, n19274, n19275, n19276,
         n19277, n19278, n19279, n19280, n19281, n19282, n19283, n19284,
         n19285, n19286, n19287, n19288, n19289, n19290, n19291, n19292,
         n19293, n19294, n19295, n19296, n19297, n19298, n19299, n19300,
         n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308,
         n19309, n19310, n19311, n19312, n19313, n19314, n19315, n19316,
         n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324,
         n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19339, n19340,
         n19341, n19342, n19343, n19344, n19345, n19346, n19347, n19348,
         n19349, n19350, n19351, n19352, n19353, n19354, n19355, n19356,
         n19357, n19358, n19359, n19360, n19361, n19362, n19363, n19364,
         n19365, n19366, n19367, n19368, n19369, n19370, n19371, n19372,
         n19373, n19374, n19375, n19376, n19377, n19378, n19379, n19380,
         n19381, n19382, n19383, n19384, n19385, n19386, n19387, n19388,
         n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396,
         n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19419, n19420,
         n19421, n19422, n19423, n19424, n19425, n19426, n19427, n19428,
         n19429, n19430, n19431, n19432, n19433, n19434, n19435, n19436,
         n19437, n19438, n19439, n19440, n19441, n19442, n19443, n19444,
         n19445, n19446, n19447, n19448, n19449, n19450, n19451, n19452,
         n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19460,
         n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468,
         n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476,
         n19477, n19478, n19479, n19480, n19481, n19482, n19483, n19484,
         n19485, n19486, n19487, n19488, n19489, n19490, n19491, n19492,
         n19493, n19494, n19495, n19496, n19497, n19498, n19499, n19500,
         n19501, n19502, n19503, n19504, n19505, n19506, n19507, n19508,
         n19509, n19510, n19511, n19512, n19513, n19514, n19515, n19516,
         n19517, n19518, n19519, n19520, n19521, n19522, n19523, n19524,
         n19525, n19526, n19527, n19528, n19529, n19530, n19531, n19532,
         n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540,
         n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
         n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556,
         n19557, n19558, n19559, n19560, n19561, n19562, n19563, n19564,
         n19565, n19566, n19567, n19568, n19569, n19570, n19571, n19572,
         n19573, n19574, n19575, n19576, n19577, n19578, n19579, n19580,
         n19581, n19582, n19583, n19584, n19585, n19586, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19604,
         n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612,
         n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
         n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628,
         n19629, n19630, n19631, n19632, n19633, n19634, n19635, n19636,
         n19637, n19638, n19639, n19640, n19641, n19642, n19643, n19644,
         n19645, n19646, n19647, n19648, n19649, n19650, n19651, n19652,
         n19653, n19654, n19655, n19656, n19657, n19658, n19659, n19660,
         n19661, n19662, n19663, n19664, n19665, n19666, n19667, n19668,
         n19669, n19670, n19671, n19672, n19673, n19674, n19675, n19676,
         n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684,
         n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
         n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700,
         n19701, n19702, n19703, n19704, n19705, n19706, n19707, n19708,
         n19709, n19710, n19711, n19712, n19713, n19714, n19715, n19716,
         n19717, n19718, n19719, n19720, n19721, n19722, n19723, n19724,
         n19725, n19726, n19727, n19728, n19729, n19730, n19731, n19732,
         n19733, n19734, n19735, n19736, n19737, n19738, n19739, n19740,
         n19741, n19742, n19743, n19744, n19745, n19746, n19747, n19748,
         n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756,
         n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
         n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772,
         n19773, n19774, n19775, n19776, n19777, n19778, n19779, n19780,
         n19781, n19782, n19783, n19784, n19785, n19786, n19787, n19788,
         n19789, n19790, n19791, n19792, n19793, n19794, n19795, n19796,
         n19797, n19798, n19799, n19800, n19801, n19802, n19803, n19804,
         n19805, n19806, n19807, n19808, n19809, n19810, n19811, n19812,
         n19813, n19814, n19815, n19816, n19817, n19818, n19819, n19820,
         n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828,
         n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
         n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844,
         n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852,
         n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860,
         n19861, n19862, n19863, n19864, n19865, n19866, n19867, n19868,
         n19869, n19870, n19871, n19872, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19890, n19891, n19892,
         n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900,
         n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
         n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916,
         n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924,
         n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932,
         n19933, n19934, n19935, n19936, n19937, n19938, n19939, n19940,
         n19941, n19942, n19943, n19944, n19945, n19946, n19947, n19948,
         n19949, n19950, n19951, n19952, n19953, n19954, n19955, n19956,
         n19957, n19958, n19959, n19960, n19961, n19962, n19963, n19964,
         n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972,
         n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
         n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988,
         n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996,
         n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004,
         n20005, n20006, n20007, n20008, n20009, n20010, n20011, n20012,
         n20013, n20014, n20015, n20016, n20017, n20018, n20019, n20020,
         n20021, n20022, n20023, n20024, n20025, n20026, n20027, n20028,
         n20029, n20030, n20031, n20032, n20033, n20034, n20035, n20036,
         n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044,
         n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
         n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060,
         n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068,
         n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076,
         n20077, n20078, n20079, n20080, n20081, n20082, n20083, n20084,
         n20085, n20086, n20087, n20088, n20089, n20090, n20091, n20092,
         n20093, n20094, n20095, n20096, n20097, n20098, n20099, n20100,
         n20101, n20102, n20103, n20104, n20105, n20106, n20107, n20108,
         n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116,
         n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
         n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132,
         n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140,
         n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148,
         n20149, n20150, n20151, n20152, n20153, n20154, n20155, n20156,
         n20157, n20158, n20159, n20160, n20161, n20162, n20163, n20164,
         n20165, n20166, n20167, n20168, n20169, n20170, n20171, n20172,
         n20173, n20174, n20175, n20176, n20177, n20178, n20179, n20180,
         n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188,
         n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
         n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204,
         n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212,
         n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220,
         n20221, n20222, n20223, n20224, n20225, n20226, n20227, n20228,
         n20229, n20230, n20231, n20232, n20233, n20234, n20235, n20236,
         n20237, n20238, n20239, n20240, n20241, n20242, n20243, n20244,
         n20245, n20246, n20247, n20248, n20249, n20250, n20251, n20252,
         n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260,
         n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
         n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276,
         n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284,
         n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292,
         n20293, n20294, n20295, n20296, n20297, n20298, n20299, n20300,
         n20301, n20302, n20303, n20304, n20305, n20306, n20307, n20308,
         n20309, n20310, n20311, n20312, n20313, n20314, n20315, n20316,
         n20317, n20318, n20319, n20320, n20321, n20322, n20323, n20324,
         n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332,
         n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
         n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348,
         n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356,
         n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364,
         n20365, n20366, n20367, n20368, n20369, n20370, n20371, n20372,
         n20373, n20374, n20375, n20376, n20377, n20378, n20379, n20380,
         n20381, n20382, n20383, n20384, n20385, n20386, n20387, n20388,
         n20389, n20390, n20391, n20392, n20393, n20394, n20395, n20396,
         n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404,
         n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
         n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420,
         n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428,
         n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436,
         n20437, n20438, n20439, n20440, n20441, n20442, n20443, n20444,
         n20445, n20446, n20447, n20448, n20449, n20450, n20451, n20452,
         n20453, n20454, n20455, n20456, n20457, n20458, n20459, n20460,
         n20461, n20462, n20463, n20464, n20465, n20466, n20467, n20468,
         n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476,
         n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
         n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492,
         n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500,
         n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508,
         n20509, n20510, n20511, n20512, n20513, n20514, n20515, n20516,
         n20517, n20518, n20519, n20520, n20521, n20522, n20523, n20524,
         n20525, n20526, n20527, n20528, n20529, n20530, n20531, n20532,
         n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
         n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548,
         n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556,
         n20557, n20558, n20559, n20560, n20561, n20562, n20563, n20564,
         n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572,
         n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580,
         n20581, n20582, n20583, n20584, n20585, n20586, n20587, n20588,
         n20589, n20590, n20591, n20592, n20593, n20594, n20595, n20596,
         n20597, n20598, n20599, n20600, n20601, n20602, n20603, n20604,
         n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
         n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620,
         n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628,
         n20629, n20630, n20631, n20632, n20633, n20634, n20635, n20636,
         n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644,
         n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652,
         n20653, n20654, n20655, n20656, n20657, n20658, n20659, n20660,
         n20661, n20662, n20663, n20664, n20665, n20666, n20667, n20668,
         n20669, n20670, n20671, n20672, n20673, n20674, n20675, n20676,
         n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
         n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692,
         n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700,
         n20701, n20702, n20703, n20704, n20705, n20706, n20707, n20708,
         n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716,
         n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724,
         n20725, n20726, n20727, n20728, n20729, n20730, n20731, n20732,
         n20733, n20734, n20735, n20736, n20737, n20738, n20739, n20740,
         n20741, n20742, n20743, n20744, n20745, n20746, n20747, n20748,
         n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
         n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764,
         n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772,
         n20773, n20774, n20775, n20776, n20777, n20778, n20779, n20780,
         n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788,
         n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796,
         n20797, n20798, n20799, n20800, n20801, n20802, n20803, n20804,
         n20805, n20806, n20807, n20808, n20809, n20810, n20811, n20812,
         n20813, n20814, n20815, n20816, n20817, n20818, n20819, n20820,
         n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
         n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836,
         n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844,
         n20845, n20846, n20847, n20848, n20849, n20850, n20851, n20852,
         n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860,
         n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868,
         n20869, n20870, n20871, n20872, n20873, n20874, n20875, n20876,
         n20877, n20878, n20879, n20880, n20881, n20882, n20883, n20884,
         n20885, n20886, n20887, n20888, n20889, n20890, n20891, n20892,
         n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
         n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908,
         n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916,
         n20917, n20918, n20919, n20920, n20921, n20922, n20923, n20924,
         n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932,
         n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940,
         n20941, n20942, n20943, n20944, n20945, n20946, n20947, n20948,
         n20949, n20950, n20951, n20952, n20953, n20954, n20955, n20956,
         n20957, n20958, n20959, n20960, n20961, n20962, n20963, n20964,
         n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
         n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980,
         n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988,
         n20989, n20990, n20991, n20992, n20993, n20994, n20995, n20996,
         n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004,
         n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012,
         n21013, n21014, n21015, n21016, n21017, n21018, n21019, n21020,
         n21021, n21022, n21023, n21024, n21025, n21026, n21027, n21028,
         n21029, n21030, n21031, n21032, n21033, n21034, n21035, n21036,
         n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
         n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052,
         n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060,
         n21061, n21062, n21063, n21064, n21065, n21066, n21067, n21068,
         n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076,
         n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084,
         n21085, n21086, n21087, n21088, n21089, n21090, n21091, n21092,
         n21093, n21094, n21095, n21096, n21097, n21098, n21099, n21100,
         n21101, n21102, n21103, n21104, n21105, n21106, n21107, n21108,
         n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
         n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124,
         n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132,
         n21133, n21134, n21135, n21136, n21137, n21138, n21139, n21140,
         n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148,
         n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156,
         n21157, n21158, n21159, n21160, n21161, n21162, n21163, n21164,
         n21165, n21166, n21167, n21168, n21169, n21170, n21171, n21172,
         n21173, n21174, n21175, n21176, n21177, n21178, n21179, n21180,
         n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
         n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196,
         n21197, n21198, n21199, n21200;

  OR2_X1 U11255 ( .A1(n17514), .A2(n17702), .ZN(n9942) );
  OAI21_X1 U11256 ( .B1(n11494), .B2(n11493), .A(n11498), .ZN(n18606) );
  NOR2_X1 U11257 ( .A1(n11399), .A2(n11398), .ZN(n16989) );
  CLKBUF_X2 U11258 ( .A(n11379), .Z(n17116) );
  INV_X1 U11259 ( .A(n12584), .ZN(n19976) );
  CLKBUF_X2 U11260 ( .A(n12581), .Z(n12584) );
  CLKBUF_X2 U11261 ( .A(n11876), .Z(n9816) );
  AND2_X1 U11262 ( .A1(n14262), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11862) );
  AND2_X1 U11263 ( .A1(n14265), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11881) );
  INV_X1 U11264 ( .A(n9858), .ZN(n14079) );
  CLKBUF_X2 U11265 ( .A(n9830), .Z(n17130) );
  CLKBUF_X2 U11266 ( .A(n11876), .Z(n9815) );
  CLKBUF_X2 U11267 ( .A(n12001), .Z(n14258) );
  BUF_X1 U11268 ( .A(n9812), .Z(n17077) );
  INV_X1 U11269 ( .A(n17147), .ZN(n15453) );
  CLKBUF_X2 U11270 ( .A(n10318), .Z(n10855) );
  NOR2_X2 U11271 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11190), .ZN(
        n17129) );
  BUF_X1 U11272 ( .A(n10441), .Z(n13596) );
  NAND2_X1 U11273 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18601) );
  INV_X2 U11274 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11412) );
  BUF_X1 U11275 ( .A(n13047), .Z(n9817) );
  INV_X2 U11276 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18764) );
  CLKBUF_X1 U11277 ( .A(n11065), .Z(n11030) );
  CLKBUF_X2 U11278 ( .A(n10443), .Z(n11051) );
  CLKBUF_X2 U11279 ( .A(n10315), .Z(n10983) );
  CLKBUF_X2 U11280 ( .A(n11066), .Z(n10906) );
  CLKBUF_X2 U11281 ( .A(n11075), .Z(n10935) );
  BUF_X1 U11282 ( .A(n10342), .Z(n11745) );
  AND4_X1 U11283 ( .A1(n10265), .A2(n10264), .A3(n10263), .A4(n10262), .ZN(
        n10266) );
  AND2_X1 U11284 ( .A1(n10254), .A2(n10260), .ZN(n11075) );
  OAI221_X2 U11285 ( .B1(n11446), .B2(n18587), .C1(n11446), .C2(n11445), .A(
        n18642), .ZN(n18127) );
  NOR3_X2 U11286 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18652), .A3(n18812), 
        .ZN(n18642) );
  CLKBUF_X1 U11287 ( .A(n18062), .Z(n9811) );
  NOR3_X1 U11288 ( .A1(n17319), .A2(n18588), .A3(n18127), .ZN(n18062) );
  AND4_X1 U11289 ( .A1(n10287), .A2(n10286), .A3(n10285), .A4(n10284), .ZN(
        n10288) );
  CLKBUF_X2 U11290 ( .A(n10343), .Z(n11076) );
  AND2_X2 U11291 ( .A1(n10242), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10260) );
  INV_X1 U11292 ( .A(n13489), .ZN(n12017) );
  AND3_X1 U11294 ( .A1(n10308), .A2(n10307), .A3(n10306), .ZN(n9840) );
  NAND2_X1 U11295 ( .A1(n12033), .A2(n15344), .ZN(n12582) );
  BUF_X1 U11296 ( .A(n12094), .Z(n12481) );
  BUF_X1 U11297 ( .A(n12481), .Z(n13970) );
  NAND2_X1 U11298 ( .A1(n12131), .A2(n16283), .ZN(n19564) );
  CLKBUF_X3 U11299 ( .A(n11245), .Z(n17152) );
  AND2_X1 U11300 ( .A1(n20149), .A2(n13447), .ZN(n13442) );
  OR2_X1 U11301 ( .A1(n9824), .A2(n11519), .ZN(n10240) );
  XNOR2_X1 U11302 ( .A(n12364), .B(n12362), .ZN(n14917) );
  INV_X1 U11304 ( .A(n17064), .ZN(n11326) );
  INV_X2 U11305 ( .A(n11326), .ZN(n17082) );
  INV_X1 U11306 ( .A(n17737), .ZN(n17528) );
  AND3_X1 U11307 ( .A1(n9942), .A2(n10229), .A3(n10163), .ZN(n11314) );
  INV_X1 U11308 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13577) );
  INV_X1 U11309 ( .A(n11227), .ZN(n11237) );
  AND2_X2 U11310 ( .A1(n13377), .A2(n11550), .ZN(n10173) );
  NOR2_X2 U11311 ( .A1(n17342), .A2(n17395), .ZN(n17312) );
  NAND2_X2 U11312 ( .A1(n12093), .A2(n12092), .ZN(n12109) );
  OAI21_X2 U11313 ( .B1(n14859), .B2(n10092), .A(n10094), .ZN(n14142) );
  AND2_X1 U11314 ( .A1(n14858), .A2(n14857), .ZN(n14859) );
  NAND2_X2 U11315 ( .A1(n10603), .A2(n10582), .ZN(n13589) );
  NOR2_X2 U11316 ( .A1(n16489), .A2(n17413), .ZN(n11498) );
  NAND2_X1 U11317 ( .A1(n10500), .A2(n11586), .ZN(n10513) );
  NOR2_X2 U11318 ( .A1(n11817), .A2(n12240), .ZN(n12241) );
  OAI21_X2 U11319 ( .B1(n11535), .B2(n20156), .A(n11534), .ZN(n11536) );
  OAI21_X2 U11320 ( .B1(n13513), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n10491), 
        .ZN(n11535) );
  NOR2_X2 U11322 ( .A1(n9817), .A2(n12045), .ZN(n12029) );
  NAND2_X2 U11323 ( .A1(n12071), .A2(n12070), .ZN(n9945) );
  NAND2_X2 U11324 ( .A1(n11829), .A2(n11828), .ZN(n12026) );
  CLKBUF_X3 U11325 ( .A(n11269), .Z(n9812) );
  NOR2_X1 U11326 ( .A1(n18601), .A2(n11192), .ZN(n11269) );
  INV_X8 U11327 ( .A(n15405), .ZN(n17142) );
  NOR2_X2 U11328 ( .A1(n13951), .A2(n14901), .ZN(n13865) );
  INV_X1 U11329 ( .A(n12148), .ZN(n15317) );
  AND2_X1 U11331 ( .A1(n14256), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11876) );
  NAND2_X2 U11332 ( .A1(n12226), .A2(n19004), .ZN(n12253) );
  NAND2_X1 U11335 ( .A1(n11582), .A2(n11581), .ZN(n13734) );
  NAND2_X1 U11336 ( .A1(n10131), .A2(n12221), .ZN(n12795) );
  INV_X8 U11337 ( .A(n14587), .ZN(n9820) );
  NAND2_X1 U11338 ( .A1(n10581), .A2(n10550), .ZN(n14716) );
  NAND2_X1 U11339 ( .A1(n11539), .A2(n11538), .ZN(n11541) );
  NOR2_X1 U11340 ( .A1(n15816), .A2(n15821), .ZN(n13622) );
  NAND2_X1 U11341 ( .A1(n9956), .A2(n9955), .ZN(n10106) );
  NAND2_X1 U11342 ( .A1(n10461), .A2(n10496), .ZN(n10500) );
  NAND2_X1 U11343 ( .A1(n13019), .A2(n13018), .ZN(n13025) );
  NOR2_X2 U11344 ( .A1(n17982), .A2(n18615), .ZN(n18053) );
  NAND2_X1 U11345 ( .A1(n10411), .A2(n10410), .ZN(n10481) );
  AND3_X1 U11346 ( .A1(n10397), .A2(n10396), .A3(n10395), .ZN(n10419) );
  OR2_X1 U11347 ( .A1(n17808), .A2(n17809), .ZN(n10193) );
  XNOR2_X1 U11348 ( .A(n11283), .B(n11449), .ZN(n11284) );
  NOR2_X1 U11349 ( .A1(n17829), .A2(n17820), .ZN(n17819) );
  OR2_X1 U11350 ( .A1(n10240), .A2(n11641), .ZN(n10395) );
  CLKBUF_X1 U11351 ( .A(n10388), .Z(n11641) );
  NAND2_X1 U11352 ( .A1(n10391), .A2(n10388), .ZN(n10342) );
  OR2_X1 U11353 ( .A1(n9934), .A2(n11242), .ZN(n11449) );
  INV_X2 U11354 ( .A(n19283), .ZN(n12023) );
  CLKBUF_X2 U11355 ( .A(n12022), .Z(n13016) );
  INV_X2 U11356 ( .A(n13443), .ZN(n20149) );
  INV_X2 U11357 ( .A(n13447), .ZN(n20156) );
  AND4_X1 U11358 ( .A1(n10355), .A2(n10354), .A3(n10353), .A4(n10352), .ZN(
        n10361) );
  OR2_X2 U11359 ( .A1(n10279), .A2(n10278), .ZN(n10325) );
  BUF_X2 U11360 ( .A(n9831), .Z(n17150) );
  AOI21_X1 U11361 ( .B1(n10315), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n10316), .ZN(n10322) );
  AND2_X2 U11362 ( .A1(n14258), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12726) );
  CLKBUF_X2 U11363 ( .A(n10370), .Z(n13325) );
  INV_X4 U11364 ( .A(n11237), .ZN(n17132) );
  BUF_X2 U11365 ( .A(n10434), .Z(n11068) );
  BUF_X2 U11366 ( .A(n11007), .Z(n11029) );
  BUF_X2 U11367 ( .A(n10448), .Z(n11070) );
  CLKBUF_X2 U11368 ( .A(n10369), .Z(n10894) );
  BUF_X2 U11369 ( .A(n10375), .Z(n11067) );
  OR2_X1 U11370 ( .A1(n16856), .A2(n11191), .ZN(n17108) );
  INV_X4 U11371 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11987) );
  NOR2_X2 U11372 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10261) );
  AND2_X1 U11373 ( .A1(n12812), .A2(n12811), .ZN(n12813) );
  AND2_X1 U11374 ( .A1(n12830), .A2(n12829), .ZN(n12831) );
  AOI211_X1 U11375 ( .C1(n13997), .C2(n19242), .A(n13976), .B(n13975), .ZN(
        n13977) );
  AOI211_X1 U11376 ( .C1(n13997), .C2(n19262), .A(n13996), .B(n13995), .ZN(
        n13998) );
  OR2_X1 U11377 ( .A1(n12821), .A2(n16172), .ZN(n12830) );
  AOI21_X1 U11378 ( .B1(n13852), .B2(n13851), .A(n13850), .ZN(n13853) );
  AND2_X1 U11379 ( .A1(n10226), .A2(n11791), .ZN(n11792) );
  AND2_X1 U11380 ( .A1(n15208), .A2(n15207), .ZN(n15231) );
  NAND2_X1 U11381 ( .A1(n10145), .A2(n13849), .ZN(n13847) );
  AND2_X1 U11382 ( .A1(n9958), .A2(n15018), .ZN(n15003) );
  OR2_X1 U11383 ( .A1(n14304), .A2(n20131), .ZN(n10226) );
  NAND2_X1 U11384 ( .A1(n10143), .A2(n9976), .ZN(n13848) );
  OR2_X1 U11385 ( .A1(n15203), .A2(n10224), .ZN(n15208) );
  NAND2_X1 U11386 ( .A1(n11783), .A2(n11785), .ZN(n14304) );
  OR2_X1 U11387 ( .A1(n10233), .A2(n11784), .ZN(n11785) );
  NAND2_X1 U11388 ( .A1(n11601), .A2(n11600), .ZN(n11604) );
  AND2_X1 U11389 ( .A1(n10214), .A2(n12804), .ZN(n10217) );
  NAND2_X1 U11390 ( .A1(n14175), .A2(n10102), .ZN(n14751) );
  AOI21_X1 U11391 ( .B1(n9939), .B2(n17739), .A(n9938), .ZN(n16335) );
  NOR2_X1 U11392 ( .A1(n14768), .A2(n14770), .ZN(n14769) );
  NAND2_X1 U11393 ( .A1(n14773), .A2(n14146), .ZN(n14172) );
  XNOR2_X1 U11394 ( .A(n13973), .B(n13972), .ZN(n16060) );
  NAND2_X1 U11395 ( .A1(n14145), .A2(n14144), .ZN(n14146) );
  OR2_X1 U11396 ( .A1(n11321), .A2(n17734), .ZN(n15555) );
  XNOR2_X1 U11397 ( .A(n12253), .B(n15272), .ZN(n13727) );
  CLKBUF_X1 U11398 ( .A(n13743), .Z(n13819) );
  NAND2_X1 U11399 ( .A1(n15296), .A2(n15297), .ZN(n15295) );
  NOR2_X1 U11400 ( .A1(n17702), .A2(n17482), .ZN(n16362) );
  AND2_X1 U11401 ( .A1(n12786), .A2(n19234), .ZN(n15296) );
  NOR2_X1 U11402 ( .A1(n13758), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10196) );
  NAND3_X1 U11403 ( .A1(n10172), .A2(n10174), .A3(n10171), .ZN(n13534) );
  NAND2_X1 U11404 ( .A1(n9820), .A2(n11591), .ZN(n13758) );
  BUF_X1 U11405 ( .A(n12787), .Z(n12789) );
  OR2_X1 U11406 ( .A1(n14797), .A2(n10099), .ZN(n14091) );
  NAND3_X1 U11407 ( .A1(n12180), .A2(n12781), .A3(n12234), .ZN(n12228) );
  NOR2_X1 U11408 ( .A1(n14791), .A2(n14792), .ZN(n14793) );
  AND2_X1 U11409 ( .A1(n12201), .A2(n12200), .ZN(n12227) );
  NAND2_X1 U11410 ( .A1(n9990), .A2(n9847), .ZN(n11567) );
  OR2_X1 U11411 ( .A1(n12198), .A2(n12197), .ZN(n12201) );
  CLKBUF_X1 U11412 ( .A(n11180), .Z(n14496) );
  XNOR2_X1 U11413 ( .A(n11541), .B(n11540), .ZN(n13304) );
  NAND2_X1 U11414 ( .A1(n19027), .A2(n13222), .ZN(n10097) );
  OAI21_X1 U11415 ( .B1(n13097), .B2(n13098), .A(n13220), .ZN(n19925) );
  AND2_X1 U11416 ( .A1(n13394), .A2(n13395), .ZN(n13916) );
  NAND2_X2 U11417 ( .A1(n14502), .A2(n13280), .ZN(n14499) );
  NAND2_X1 U11418 ( .A1(n12117), .A2(n12116), .ZN(n19734) );
  AND2_X1 U11419 ( .A1(n10207), .A2(n13910), .ZN(n19423) );
  AND2_X1 U11420 ( .A1(n10207), .A2(n12112), .ZN(n15354) );
  NAND2_X1 U11421 ( .A1(n20078), .A2(n13608), .ZN(n14439) );
  OR2_X1 U11422 ( .A1(n12142), .A2(n12141), .ZN(n12181) );
  OR2_X1 U11423 ( .A1(n12130), .A2(n16283), .ZN(n12185) );
  INV_X1 U11424 ( .A(n17703), .ZN(n9944) );
  OR2_X1 U11425 ( .A1(n12142), .A2(n12136), .ZN(n19660) );
  OR2_X1 U11426 ( .A1(n12132), .A2(n19251), .ZN(n19620) );
  OR2_X2 U11427 ( .A1(n12113), .A2(n12112), .ZN(n15332) );
  OR2_X1 U11428 ( .A1(n12115), .A2(n12141), .ZN(n19595) );
  AND2_X1 U11429 ( .A1(n19029), .A2(n13096), .ZN(n13098) );
  OR2_X1 U11430 ( .A1(n12132), .A2(n16283), .ZN(n19765) );
  AND2_X1 U11431 ( .A1(n9872), .A2(n10184), .ZN(n17703) );
  OR2_X1 U11432 ( .A1(n13221), .A2(n13095), .ZN(n13096) );
  OR2_X1 U11433 ( .A1(n13099), .A2(n12138), .ZN(n12140) );
  NAND2_X2 U11434 ( .A1(n10106), .A2(n12488), .ZN(n13099) );
  OAI211_X1 U11435 ( .C1(n10106), .C2(n10105), .A(n13094), .B(n10104), .ZN(
        n13221) );
  NOR2_X2 U11436 ( .A1(n18808), .A2(n16474), .ZN(n17822) );
  INV_X2 U11437 ( .A(n17283), .ZN(n17337) );
  XNOR2_X1 U11438 ( .A(n13025), .B(n13039), .ZN(n13038) );
  NOR2_X1 U11439 ( .A1(n17641), .A2(n11300), .ZN(n11301) );
  NOR2_X1 U11440 ( .A1(n13683), .A2(n15340), .ZN(n19126) );
  NOR2_X1 U11441 ( .A1(n13683), .A2(n15338), .ZN(n19127) );
  OR2_X1 U11442 ( .A1(n12313), .A2(n12311), .ZN(n12308) );
  OR2_X1 U11443 ( .A1(n10527), .A2(n10528), .ZN(n10525) );
  NAND2_X1 U11444 ( .A1(n12274), .A2(n12279), .ZN(n12313) );
  XNOR2_X1 U11445 ( .A(n11299), .B(n11300), .ZN(n17749) );
  AND2_X1 U11446 ( .A1(n12487), .A2(n12107), .ZN(n12108) );
  AND2_X2 U11447 ( .A1(n12111), .A2(n12086), .ZN(n19076) );
  XNOR2_X1 U11448 ( .A(n10481), .B(n10479), .ZN(n10502) );
  NAND2_X1 U11449 ( .A1(n12277), .A2(n12350), .ZN(n12274) );
  CLKBUF_X2 U11450 ( .A(n12081), .Z(n12111) );
  OR2_X1 U11451 ( .A1(n11294), .A2(n11297), .ZN(n10178) );
  NOR2_X2 U11452 ( .A1(n13837), .A2(n18606), .ZN(n18617) );
  OR2_X1 U11453 ( .A1(n12069), .A2(n12068), .ZN(n12070) );
  NOR2_X1 U11454 ( .A1(n12266), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10072) );
  NAND2_X1 U11455 ( .A1(n12257), .A2(n12256), .ZN(n12266) );
  NAND3_X1 U11456 ( .A1(n10486), .A2(n10408), .A3(n10407), .ZN(n10519) );
  NOR2_X1 U11457 ( .A1(n10428), .A2(n10427), .ZN(n10479) );
  AOI21_X1 U11458 ( .B1(n12102), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12079), .ZN(n12090) );
  NAND2_X1 U11459 ( .A1(n12100), .A2(n12099), .ZN(n12106) );
  AND3_X1 U11460 ( .A1(n11895), .A2(n9844), .A3(n10075), .ZN(n12257) );
  CLKBUF_X1 U11461 ( .A(n12078), .Z(n12102) );
  NAND2_X1 U11462 ( .A1(n10424), .A2(n10475), .ZN(n10407) );
  NOR2_X1 U11463 ( .A1(n17416), .A2(n11491), .ZN(n16473) );
  NAND2_X2 U11464 ( .A1(n17416), .A2(n17415), .ZN(n17443) );
  OR2_X1 U11465 ( .A1(n12095), .A2(n13507), .ZN(n12097) );
  NAND2_X1 U11466 ( .A1(n12578), .A2(n12039), .ZN(n12058) );
  AND2_X1 U11467 ( .A1(n12019), .A2(n12018), .ZN(n12020) );
  CLKBUF_X1 U11468 ( .A(n12578), .Z(n16266) );
  NAND2_X1 U11469 ( .A1(n11115), .A2(n10154), .ZN(n10153) );
  NOR2_X1 U11470 ( .A1(n12072), .A2(n12061), .ZN(n12062) );
  BUF_X2 U11471 ( .A(n12072), .Z(n13873) );
  AND2_X1 U11472 ( .A1(n10364), .A2(n20156), .ZN(n10169) );
  AND2_X1 U11473 ( .A1(n12862), .A2(n12402), .ZN(n12578) );
  NOR2_X1 U11474 ( .A1(n17332), .A2(n11457), .ZN(n11268) );
  CLKBUF_X1 U11475 ( .A(n12028), .Z(n13048) );
  INV_X1 U11476 ( .A(n12028), .ZN(n12468) );
  AND2_X1 U11477 ( .A1(n10086), .A2(n10083), .ZN(n12010) );
  NAND2_X2 U11478 ( .A1(n9873), .A2(n12583), .ZN(n12759) );
  NAND2_X1 U11479 ( .A1(n17203), .A2(n18180), .ZN(n15584) );
  NAND2_X1 U11480 ( .A1(n11659), .A2(n10421), .ZN(n13106) );
  NOR2_X1 U11481 ( .A1(n12015), .A2(n12582), .ZN(n12016) );
  AND2_X1 U11482 ( .A1(n12032), .A2(n19984), .ZN(n12407) );
  INV_X1 U11483 ( .A(n18157), .ZN(n15442) );
  INV_X1 U11484 ( .A(n10240), .ZN(n15538) );
  INV_X1 U11485 ( .A(n18808), .ZN(n18164) );
  AND2_X1 U11486 ( .A1(n13328), .A2(n20149), .ZN(n10417) );
  OR2_X1 U11487 ( .A1(n11850), .A2(n11849), .ZN(n12603) );
  NAND3_X1 U11488 ( .A1(n11378), .A2(n11377), .A3(n11376), .ZN(n18157) );
  INV_X1 U11489 ( .A(n11411), .ZN(n18180) );
  NOR2_X1 U11490 ( .A1(n11367), .A2(n11366), .ZN(n11411) );
  CLKBUF_X1 U11491 ( .A(n10391), .Z(n11531) );
  NAND2_X1 U11492 ( .A1(n9935), .A2(n9936), .ZN(n9934) );
  NAND3_X1 U11493 ( .A1(n11281), .A2(n11280), .A3(n11279), .ZN(n15585) );
  NAND4_X2 U11494 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n13443) );
  OR2_X2 U11495 ( .A1(n16423), .A2(n16374), .ZN(n16426) );
  INV_X1 U11496 ( .A(n12033), .ZN(n10206) );
  NAND2_X1 U11497 ( .A1(n11988), .A2(n11987), .ZN(n10084) );
  NAND2_X1 U11498 ( .A1(n11993), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10085) );
  AND4_X1 U11499 ( .A1(n10379), .A2(n10378), .A3(n10377), .A4(n10376), .ZN(
        n10385) );
  NAND2_X1 U11500 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  NAND2_X2 U11501 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19892), .ZN(n19899) );
  CLKBUF_X3 U11502 ( .A(n17129), .Z(n17148) );
  AND4_X1 U11503 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10362) );
  AND4_X1 U11504 ( .A1(n10374), .A2(n10373), .A3(n10372), .A4(n10371), .ZN(
        n10386) );
  AND4_X1 U11505 ( .A1(n10248), .A2(n10247), .A3(n10246), .A4(n10245), .ZN(
        n10269) );
  AND4_X1 U11506 ( .A1(n10347), .A2(n10346), .A3(n10345), .A4(n10344), .ZN(
        n10363) );
  AND4_X1 U11507 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10384) );
  AND4_X1 U11508 ( .A1(n10253), .A2(n10252), .A3(n10251), .A4(n10250), .ZN(
        n10268) );
  AND4_X1 U11509 ( .A1(n10258), .A2(n10257), .A3(n10256), .A4(n10255), .ZN(
        n10267) );
  AND4_X1 U11510 ( .A1(n11992), .A2(n11991), .A3(n11990), .A4(n11989), .ZN(
        n11993) );
  AND4_X1 U11511 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n11988) );
  AND4_X1 U11512 ( .A1(n10368), .A2(n10367), .A3(n10366), .A4(n10365), .ZN(
        n10387) );
  AND4_X1 U11513 ( .A1(n10359), .A2(n10358), .A3(n10357), .A4(n10356), .ZN(
        n10360) );
  AND4_X1 U11514 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n10299) );
  AND4_X1 U11515 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10298) );
  INV_X2 U11516 ( .A(n18036), .ZN(n9821) );
  INV_X2 U11517 ( .A(n20759), .ZN(n9822) );
  CLKBUF_X2 U11518 ( .A(n11379), .Z(n17151) );
  INV_X2 U11519 ( .A(n16454), .ZN(U215) );
  BUF_X2 U11520 ( .A(n15367), .Z(n9830) );
  BUF_X2 U11521 ( .A(n9812), .Z(n17131) );
  INV_X4 U11522 ( .A(n17108), .ZN(n17050) );
  CLKBUF_X3 U11523 ( .A(n11223), .Z(n17149) );
  CLKBUF_X3 U11524 ( .A(n17024), .Z(n17144) );
  BUF_X2 U11525 ( .A(n15448), .Z(n9831) );
  CLKBUF_X3 U11526 ( .A(n11271), .Z(n17143) );
  CLKBUF_X2 U11527 ( .A(n11249), .Z(n17024) );
  INV_X2 U11528 ( .A(n18799), .ZN(n18733) );
  INV_X2 U11529 ( .A(n19990), .ZN(n19892) );
  INV_X2 U11530 ( .A(n16464), .ZN(n16466) );
  NAND2_X1 U11531 ( .A1(n11412), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11191) );
  OR2_X1 U11532 ( .A1(n18782), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11193) );
  CLKBUF_X1 U11533 ( .A(n10847), .Z(n13432) );
  AND2_X1 U11534 ( .A1(n11798), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13690) );
  AND2_X1 U11535 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15309) );
  NOR2_X1 U11536 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11793) );
  OR2_X2 U11537 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n16856) );
  INV_X2 U11538 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18782) );
  INV_X2 U11539 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18789) );
  NAND4_X1 U11540 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n9824) );
  AND2_X1 U11541 ( .A1(n10167), .A2(n11640), .ZN(n10170) );
  AND2_X2 U11542 ( .A1(n13342), .A2(n13330), .ZN(n10315) );
  NOR2_X2 U11543 ( .A1(n15031), .A2(n15030), .ZN(n14804) );
  INV_X2 U11544 ( .A(n12962), .ZN(n10166) );
  AND2_X4 U11545 ( .A1(n12031), .A2(n19971), .ZN(n12594) );
  NOR2_X2 U11546 ( .A1(n15477), .A2(n16342), .ZN(n15476) );
  NAND2_X1 U11547 ( .A1(n19273), .A2(n12455), .ZN(n13047) );
  INV_X1 U11548 ( .A(n12455), .ZN(n19278) );
  MUX2_X1 U11549 ( .A(n10310), .B(n11638), .S(n10394), .Z(n10341) );
  AND2_X4 U11550 ( .A1(n10249), .A2(n13330), .ZN(n10369) );
  NAND2_X1 U11551 ( .A1(n13424), .A2(n13861), .ZN(n9966) );
  INV_X4 U11552 ( .A(n10325), .ZN(n10416) );
  AND2_X1 U11553 ( .A1(n10261), .A2(n13311), .ZN(n9825) );
  NAND4_X1 U11554 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n9826) );
  NAND4_X1 U11555 ( .A1(n10363), .A2(n10362), .A3(n10361), .A4(n10360), .ZN(
        n9827) );
  XNOR2_X1 U11556 ( .A(n12234), .B(n12233), .ZN(n13424) );
  XNOR2_X2 U11557 ( .A(n12111), .B(n12125), .ZN(n12112) );
  NAND3_X2 U11558 ( .A1(n10389), .A2(n11530), .A3(n11129), .ZN(n12962) );
  INV_X2 U11559 ( .A(n10402), .ZN(n11530) );
  AND2_X4 U11560 ( .A1(n10261), .A2(n13311), .ZN(n10328) );
  INV_X2 U11561 ( .A(n12026), .ZN(n13045) );
  AND2_X1 U11562 ( .A1(n13330), .A2(n13311), .ZN(n9828) );
  AND2_X1 U11563 ( .A1(n13330), .A2(n13311), .ZN(n10343) );
  AND2_X1 U11564 ( .A1(n10260), .A2(n13342), .ZN(n9829) );
  NOR2_X1 U11565 ( .A1(n18764), .A2(n11190), .ZN(n15367) );
  NOR2_X1 U11566 ( .A1(n11193), .A2(n11191), .ZN(n15448) );
  INV_X2 U11567 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11872) );
  NAND2_X2 U11568 ( .A1(n11547), .A2(n11546), .ZN(n13377) );
  OR2_X2 U11569 ( .A1(n13589), .A2(n11585), .ZN(n11547) );
  NAND2_X2 U11570 ( .A1(n10500), .A2(n10499), .ZN(n11527) );
  XNOR2_X2 U11571 ( .A(n13103), .B(n11536), .ZN(n13228) );
  AND2_X1 U11572 ( .A1(n10254), .A2(n10260), .ZN(n9832) );
  NOR2_X2 U11573 ( .A1(n13666), .A2(n13665), .ZN(n13677) );
  NAND2_X2 U11574 ( .A1(n10097), .A2(n10095), .ZN(n13666) );
  XNOR2_X2 U11575 ( .A(n11548), .B(n13384), .ZN(n13376) );
  XNOR2_X2 U11576 ( .A(n12080), .B(n9945), .ZN(n13029) );
  OAI21_X2 U11577 ( .B1(n13088), .B2(n13087), .A(n13086), .ZN(n13097) );
  OR2_X1 U11578 ( .A1(n14421), .A2(n14371), .ZN(n14356) );
  NAND2_X1 U11579 ( .A1(n14530), .A2(n11616), .ZN(n9980) );
  CLKBUF_X1 U11580 ( .A(n10328), .Z(n10981) );
  BUF_X1 U11581 ( .A(n11069), .Z(n10982) );
  OR2_X1 U11582 ( .A1(n10474), .A2(n10473), .ZN(n11529) );
  OR2_X1 U11583 ( .A1(n13596), .A2(n20718), .ZN(n10566) );
  OR2_X1 U11584 ( .A1(n9827), .A2(n20718), .ZN(n10565) );
  NAND3_X1 U11585 ( .A1(n13596), .A2(n9827), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11143) );
  AND2_X1 U11586 ( .A1(n10144), .A2(n14926), .ZN(n9976) );
  AND2_X1 U11587 ( .A1(n11854), .A2(n11853), .ZN(n11871) );
  OR2_X1 U11588 ( .A1(n12437), .A2(n12372), .ZN(n11854) );
  NAND2_X1 U11589 ( .A1(n10033), .A2(n14340), .ZN(n10032) );
  INV_X1 U11590 ( .A(n14327), .ZN(n10033) );
  INV_X1 U11591 ( .A(n13776), .ZN(n10025) );
  NAND2_X1 U11592 ( .A1(n13635), .A2(n13744), .ZN(n13743) );
  INV_X1 U11593 ( .A(n10847), .ZN(n11093) );
  NAND2_X1 U11594 ( .A1(n13217), .A2(n11669), .ZN(n11732) );
  OR2_X1 U11595 ( .A1(n10440), .A2(n10439), .ZN(n11588) );
  INV_X1 U11596 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10242) );
  INV_X1 U11597 ( .A(n14142), .ZN(n14145) );
  OAI211_X1 U11598 ( .C1(n9952), .C2(n15272), .A(n9951), .B(n12794), .ZN(
        n12800) );
  CLKBUF_X1 U11599 ( .A(n12768), .Z(n12792) );
  NAND2_X1 U11600 ( .A1(n12789), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15298) );
  NAND2_X1 U11601 ( .A1(n11518), .A2(n9824), .ZN(n10421) );
  NOR2_X1 U11602 ( .A1(n11783), .A2(n14292), .ZN(n14291) );
  NAND2_X1 U11603 ( .A1(n10951), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10994) );
  INV_X1 U11604 ( .A(n13217), .ZN(n13129) );
  NAND2_X1 U11605 ( .A1(n10065), .A2(n10063), .ZN(n10062) );
  NOR2_X1 U11606 ( .A1(n10067), .A2(n10066), .ZN(n10065) );
  INV_X1 U11607 ( .A(n14311), .ZN(n10066) );
  NAND2_X1 U11608 ( .A1(n11567), .A2(n11587), .ZN(n11593) );
  AND2_X1 U11609 ( .A1(n11637), .A2(n13153), .ZN(n11761) );
  NAND2_X1 U11610 ( .A1(n12366), .A2(n12367), .ZN(n13855) );
  AND2_X1 U11611 ( .A1(n14012), .A2(n13678), .ZN(n10098) );
  AOI21_X1 U11612 ( .B1(n13420), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n9965), .ZN(n9964) );
  NOR2_X1 U11613 ( .A1(n13420), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9963) );
  INV_X1 U11614 ( .A(n13503), .ZN(n9965) );
  NOR2_X1 U11615 ( .A1(n14901), .A2(n13952), .ZN(n13953) );
  NOR2_X1 U11616 ( .A1(n14963), .A2(n10137), .ZN(n10132) );
  NAND2_X1 U11617 ( .A1(n12328), .A2(n12327), .ZN(n12341) );
  AOI21_X1 U11618 ( .B1(n15235), .B2(n15232), .A(n14956), .ZN(n16113) );
  AND2_X1 U11619 ( .A1(n17734), .A2(n17960), .ZN(n11305) );
  INV_X1 U11620 ( .A(n13128), .ZN(n13153) );
  NAND2_X1 U11621 ( .A1(n13172), .A2(n12971), .ZN(n20798) );
  NAND2_X1 U11622 ( .A1(n14681), .A2(n20127), .ZN(n14557) );
  INV_X1 U11623 ( .A(n12228), .ZN(n12202) );
  NAND2_X1 U11624 ( .A1(n9990), .A2(n9991), .ZN(n10652) );
  NOR2_X1 U11625 ( .A1(n9898), .A2(n10602), .ZN(n9991) );
  OR2_X1 U11626 ( .A1(n10599), .A2(n10598), .ZN(n11551) );
  INV_X1 U11627 ( .A(n10565), .ZN(n10475) );
  INV_X1 U11628 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n10155) );
  XNOR2_X1 U11629 ( .A(n10487), .B(n10486), .ZN(n20252) );
  INV_X1 U11630 ( .A(n14092), .ZN(n10093) );
  XNOR2_X1 U11631 ( .A(n12228), .B(n12227), .ZN(n12787) );
  AND4_X1 U11632 ( .A1(n11922), .A2(n11921), .A3(n11920), .A4(n11919), .ZN(
        n11938) );
  OR2_X1 U11633 ( .A1(n11869), .A2(n11868), .ZN(n12612) );
  NAND4_X1 U11634 ( .A1(n10212), .A2(n12168), .A3(n10211), .A4(n10210), .ZN(
        n10209) );
  NOR2_X1 U11635 ( .A1(n12177), .A2(n12174), .ZN(n10212) );
  NOR2_X1 U11636 ( .A1(n12176), .A2(n12173), .ZN(n10211) );
  AND2_X1 U11637 ( .A1(n11840), .A2(n19971), .ZN(n10129) );
  NAND2_X1 U11638 ( .A1(n13099), .A2(n12127), .ZN(n12132) );
  NAND2_X1 U11639 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19958), .ZN(
        n12372) );
  AND2_X1 U11640 ( .A1(n11496), .A2(n11487), .ZN(n11490) );
  NOR2_X1 U11641 ( .A1(n16989), .A2(n18157), .ZN(n11431) );
  OR2_X1 U11642 ( .A1(n17325), .A2(n11291), .ZN(n11295) );
  NOR2_X1 U11643 ( .A1(n15697), .A2(n15685), .ZN(n10070) );
  NOR2_X1 U11644 ( .A1(n14315), .A2(n10032), .ZN(n10031) );
  XNOR2_X1 U11645 ( .A(n11567), .B(n10655), .ZN(n11574) );
  INV_X1 U11646 ( .A(n13569), .ZN(n10020) );
  INV_X1 U11647 ( .A(n13362), .ZN(n10613) );
  INV_X1 U11648 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13323) );
  AND2_X1 U11649 ( .A1(n9892), .A2(n10069), .ZN(n10068) );
  INV_X1 U11650 ( .A(n14396), .ZN(n10069) );
  INV_X1 U11651 ( .A(n11549), .ZN(n10175) );
  AND2_X1 U11652 ( .A1(n11692), .A2(n13217), .ZN(n11717) );
  INV_X1 U11653 ( .A(n11732), .ZN(n11735) );
  NAND2_X1 U11654 ( .A1(n10515), .A2(n10514), .ZN(n10548) );
  AND2_X1 U11655 ( .A1(n9849), .A2(n14778), .ZN(n10079) );
  NAND2_X1 U11656 ( .A1(n12350), .A2(n12296), .ZN(n12300) );
  OR2_X1 U11657 ( .A1(n12317), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12296) );
  NAND2_X1 U11658 ( .A1(n9945), .A2(n12088), .ZN(n12093) );
  INV_X1 U11659 ( .A(n12106), .ZN(n12103) );
  NAND2_X1 U11660 ( .A1(n10103), .A2(n9875), .ZN(n14175) );
  INV_X1 U11661 ( .A(n14769), .ZN(n10103) );
  AND2_X1 U11662 ( .A1(n13024), .A2(n19976), .ZN(n14198) );
  AND2_X1 U11663 ( .A1(n12023), .A2(n12033), .ZN(n9962) );
  INV_X1 U11664 ( .A(n15287), .ZN(n10120) );
  NOR2_X1 U11665 ( .A1(n11918), .A2(n11917), .ZN(n12626) );
  AND2_X1 U11666 ( .A1(n10018), .A2(n9922), .ZN(n10017) );
  NOR2_X1 U11667 ( .A1(n14969), .A2(n10019), .ZN(n10018) );
  INV_X1 U11668 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10019) );
  AND2_X1 U11669 ( .A1(n10109), .A2(n10108), .ZN(n10107) );
  INV_X1 U11670 ( .A(n14799), .ZN(n10108) );
  NOR2_X1 U11671 ( .A1(n10110), .A2(n15007), .ZN(n10109) );
  NOR2_X1 U11672 ( .A1(n10013), .A2(n15045), .ZN(n10012) );
  INV_X1 U11673 ( .A(n10015), .ZN(n10013) );
  NAND2_X1 U11674 ( .A1(n12796), .A2(n13959), .ZN(n12802) );
  INV_X1 U11675 ( .A(n12795), .ZN(n12796) );
  NAND2_X1 U11676 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10002) );
  NAND2_X1 U11677 ( .A1(n9947), .A2(n12780), .ZN(n12782) );
  NAND2_X1 U11678 ( .A1(n13424), .A2(n13423), .ZN(n9947) );
  XNOR2_X1 U11679 ( .A(n9946), .B(n12781), .ZN(n12783) );
  NAND2_X1 U11680 ( .A1(n12180), .A2(n12234), .ZN(n9946) );
  NAND2_X1 U11681 ( .A1(n12350), .A2(n12358), .ZN(n13955) );
  AND2_X1 U11682 ( .A1(n10144), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10142) );
  OR2_X1 U11683 ( .A1(n15999), .A2(n13861), .ZN(n13849) );
  NOR2_X1 U11684 ( .A1(n16044), .A2(n13861), .ZN(n12354) );
  NAND2_X1 U11685 ( .A1(n12622), .A2(n13502), .ZN(n10121) );
  AND2_X1 U11686 ( .A1(n12241), .A2(n12237), .ZN(n12236) );
  MUX2_X1 U11687 ( .A(n19283), .B(n12033), .S(n12022), .Z(n12009) );
  AND3_X1 U11688 ( .A1(n15344), .A2(n13045), .A3(n19273), .ZN(n10083) );
  OAI21_X1 U11689 ( .B1(n12037), .B2(n13016), .A(n12455), .ZN(n12034) );
  NOR2_X1 U11690 ( .A1(n13099), .A2(n12136), .ZN(n10207) );
  NAND2_X1 U11691 ( .A1(n13099), .A2(n12137), .ZN(n12130) );
  OR2_X1 U11692 ( .A1(n13029), .A2(n19076), .ZN(n12141) );
  AND2_X1 U11693 ( .A1(n12386), .A2(n11893), .ZN(n12416) );
  AND2_X1 U11694 ( .A1(n12584), .A2(n16274), .ZN(n16312) );
  NOR2_X1 U11695 ( .A1(n16473), .A2(n18810), .ZN(n16489) );
  NOR2_X1 U11696 ( .A1(n10049), .A2(n10053), .ZN(n10048) );
  INV_X1 U11697 ( .A(n10050), .ZN(n10049) );
  INV_X1 U11698 ( .A(n10048), .ZN(n10046) );
  NAND3_X1 U11699 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(n18782), .ZN(n11190) );
  NAND2_X1 U11700 ( .A1(n18764), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11192) );
  NOR3_X1 U11701 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18601), .ZN(n11249) );
  NOR2_X1 U11702 ( .A1(n15463), .A2(n16856), .ZN(n11272) );
  NOR2_X1 U11703 ( .A1(n17776), .A2(n10042), .ZN(n10041) );
  INV_X1 U11704 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10042) );
  INV_X1 U11705 ( .A(n11431), .ZN(n11494) );
  NAND2_X1 U11706 ( .A1(n10164), .A2(n17515), .ZN(n10159) );
  INV_X1 U11707 ( .A(n17535), .ZN(n10162) );
  AND2_X1 U11708 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11289), .ZN(
        n11290) );
  INV_X1 U11709 ( .A(n15584), .ZN(n18616) );
  OAI21_X1 U11710 ( .B1(n11437), .B2(n11444), .A(n11436), .ZN(n16471) );
  NAND2_X1 U11711 ( .A1(n14353), .A2(n14340), .ZN(n14339) );
  INV_X1 U11712 ( .A(n10032), .ZN(n10030) );
  AND2_X1 U11713 ( .A1(n14559), .A2(n13432), .ZN(n10972) );
  INV_X1 U11714 ( .A(n14369), .ZN(n10956) );
  NOR2_X1 U11715 ( .A1(n9845), .A2(n9925), .ZN(n10023) );
  AND2_X1 U11716 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10584), .ZN(
        n10605) );
  NOR2_X1 U11717 ( .A1(n9820), .A2(n11614), .ZN(n11615) );
  INV_X1 U11718 ( .A(n10063), .ZN(n10061) );
  NOR2_X1 U11719 ( .A1(n14357), .A2(n14342), .ZN(n14341) );
  BUF_X1 U11720 ( .A(n11610), .Z(n14572) );
  INV_X1 U11721 ( .A(n10186), .ZN(n10185) );
  OAI21_X1 U11722 ( .B1(n10187), .B2(n15734), .A(n9820), .ZN(n10186) );
  NAND2_X1 U11723 ( .A1(n14593), .A2(n10188), .ZN(n10187) );
  OR2_X1 U11724 ( .A1(n15676), .A2(n11700), .ZN(n15668) );
  AND2_X1 U11725 ( .A1(n9870), .A2(n11594), .ZN(n10198) );
  AND2_X1 U11726 ( .A1(n11691), .A2(n11690), .ZN(n15673) );
  NAND2_X1 U11727 ( .A1(n10176), .A2(n11549), .ZN(n11554) );
  INV_X1 U11728 ( .A(n10455), .ZN(n10497) );
  OR2_X1 U11729 ( .A1(n14716), .A2(n10580), .ZN(n20368) );
  INV_X1 U11730 ( .A(n20500), .ZN(n20494) );
  NOR2_X1 U11731 ( .A1(n20458), .A2(n20289), .ZN(n20606) );
  OR2_X2 U11732 ( .A1(n10324), .A2(n10323), .ZN(n13608) );
  NAND2_X1 U11733 ( .A1(n12390), .A2(n12389), .ZN(n12442) );
  OR2_X1 U11734 ( .A1(n12388), .A2(n12387), .ZN(n12390) );
  AND2_X1 U11735 ( .A1(n16303), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12387) );
  NAND2_X1 U11736 ( .A1(n11853), .A2(n11852), .ZN(n12437) );
  AND2_X1 U11737 ( .A1(n13955), .A2(n12360), .ZN(n12366) );
  NAND2_X1 U11738 ( .A1(n10010), .A2(n10009), .ZN(n10008) );
  INV_X1 U11739 ( .A(n16027), .ZN(n10009) );
  OR2_X1 U11740 ( .A1(n10004), .A2(n16092), .ZN(n10010) );
  AND2_X1 U11741 ( .A1(n12555), .A2(n12554), .ZN(n14792) );
  NOR2_X1 U11742 ( .A1(n12247), .A2(n12246), .ZN(n12248) );
  OR2_X1 U11743 ( .A1(n16267), .A2(n13007), .ZN(n12863) );
  OR2_X1 U11744 ( .A1(n13392), .A2(n13391), .ZN(n13540) );
  OR2_X1 U11745 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  AND2_X1 U11746 ( .A1(n14936), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14928) );
  NOR2_X1 U11747 ( .A1(n15962), .A2(n16028), .ZN(n14936) );
  OR2_X1 U11748 ( .A1(n14913), .A2(n9931), .ZN(n14909) );
  NOR3_X1 U11749 ( .A1(n13857), .A2(n13861), .A3(n14910), .ZN(n14901) );
  INV_X1 U11750 ( .A(n12371), .ZN(n9973) );
  NOR2_X1 U11751 ( .A1(n9973), .A2(n15081), .ZN(n9972) );
  INV_X1 U11752 ( .A(n12363), .ZN(n12362) );
  AND2_X1 U11753 ( .A1(n15100), .A2(n12480), .ZN(n15079) );
  NAND2_X1 U11754 ( .A1(n15026), .A2(n14959), .ZN(n9958) );
  NAND2_X1 U11755 ( .A1(n10150), .A2(n9897), .ZN(n9977) );
  AND2_X1 U11756 ( .A1(n12263), .A2(n10149), .ZN(n10148) );
  INV_X1 U11757 ( .A(n13929), .ZN(n10149) );
  XNOR2_X1 U11758 ( .A(n12800), .B(n12798), .ZN(n15055) );
  AOI21_X1 U11759 ( .B1(n9950), .B2(n9949), .A(n9876), .ZN(n9952) );
  INV_X1 U11760 ( .A(n12792), .ZN(n9949) );
  OAI21_X1 U11761 ( .B1(n15283), .B2(n15284), .A(n12252), .ZN(n13728) );
  NOR2_X1 U11762 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19972) );
  AND2_X1 U11763 ( .A1(n12449), .A2(n19829), .ZN(n12810) );
  XNOR2_X1 U11764 ( .A(n13054), .B(n12596), .ZN(n13288) );
  NAND2_X1 U11765 ( .A1(n13038), .A2(n13037), .ZN(n13042) );
  INV_X1 U11766 ( .A(n15306), .ZN(n16282) );
  OR2_X1 U11767 ( .A1(n12825), .A2(n12824), .ZN(n19776) );
  NOR2_X1 U11768 ( .A1(n19916), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12825) );
  NOR2_X1 U11769 ( .A1(n18808), .A2(n11492), .ZN(n17413) );
  NAND2_X1 U11770 ( .A1(n17666), .A2(n10043), .ZN(n17624) );
  AND2_X1 U11771 ( .A1(n17664), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10043) );
  INV_X1 U11772 ( .A(n16362), .ZN(n10204) );
  NOR2_X1 U11773 ( .A1(n18588), .A2(n17319), .ZN(n10203) );
  AND2_X1 U11774 ( .A1(n10200), .A2(n10199), .ZN(n17469) );
  INV_X1 U11775 ( .A(n17470), .ZN(n10199) );
  NOR2_X1 U11776 ( .A1(n11476), .A2(n17505), .ZN(n17842) );
  NAND2_X1 U11777 ( .A1(n11313), .A2(n17702), .ZN(n17513) );
  AOI21_X1 U11778 ( .B1(n17638), .B2(n11304), .A(n17734), .ZN(n17620) );
  NAND2_X1 U11779 ( .A1(n11445), .A2(n11432), .ZN(n18588) );
  NAND2_X1 U11780 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15463) );
  NAND2_X1 U11781 ( .A1(n13434), .A2(n13433), .ZN(n15629) );
  INV_X1 U11782 ( .A(n14536), .ZN(n14454) );
  AND2_X1 U11783 ( .A1(n14502), .A2(n13281), .ZN(n14495) );
  NAND2_X1 U11784 ( .A1(n11167), .A2(n11166), .ZN(n14502) );
  NAND2_X1 U11785 ( .A1(n13149), .A2(n13153), .ZN(n11167) );
  XNOR2_X1 U11786 ( .A(n14291), .B(n11096), .ZN(n14282) );
  OR2_X1 U11787 ( .A1(n20127), .A2(n11788), .ZN(n15790) );
  NOR2_X2 U11788 ( .A1(n15530), .A2(n13128), .ZN(n20127) );
  MUX2_X1 U11789 ( .A(n14296), .B(n11681), .S(n9886), .Z(n11743) );
  NAND2_X1 U11790 ( .A1(n14507), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11619) );
  NAND2_X1 U11791 ( .A1(n14551), .A2(n14550), .ZN(n14553) );
  NAND2_X1 U11792 ( .A1(n14549), .A2(n9820), .ZN(n14551) );
  AND2_X1 U11793 ( .A1(n11761), .A2(n11644), .ZN(n15933) );
  AND2_X1 U11794 ( .A1(n11761), .A2(n11645), .ZN(n15932) );
  CLKBUF_X1 U11795 ( .A(n13513), .Z(n13514) );
  INV_X1 U11796 ( .A(n9985), .ZN(n13412) );
  INV_X1 U11797 ( .A(n20602), .ZN(n20638) );
  XNOR2_X1 U11798 ( .A(n15203), .B(n12530), .ZN(n10091) );
  OR2_X1 U11799 ( .A1(n12869), .A2(n12584), .ZN(n16173) );
  NAND2_X1 U11800 ( .A1(n10114), .A2(n10112), .ZN(n15067) );
  OR2_X1 U11801 ( .A1(n15989), .A2(n16253), .ZN(n10114) );
  AOI21_X1 U11802 ( .B1(n15063), .B2(n19257), .A(n10113), .ZN(n10112) );
  INV_X1 U11803 ( .A(n15062), .ZN(n10113) );
  AND2_X1 U11804 ( .A1(n12810), .A2(n19963), .ZN(n19263) );
  NOR2_X1 U11805 ( .A1(n19683), .A2(n19560), .ZN(n19602) );
  NOR2_X2 U11806 ( .A1(n17319), .A2(n17833), .ZN(n17739) );
  INV_X1 U11807 ( .A(n17822), .ZN(n17833) );
  XNOR2_X1 U11808 ( .A(n15557), .B(n16336), .ZN(n9939) );
  AND2_X1 U11809 ( .A1(n11138), .A2(n11157), .ZN(n11123) );
  CLKBUF_X1 U11810 ( .A(n10402), .Z(n10403) );
  NOR2_X1 U11811 ( .A1(n9819), .A2(n9961), .ZN(n9960) );
  OR2_X1 U11812 ( .A1(n11423), .A2(n11422), .ZN(n11414) );
  NAND2_X1 U11813 ( .A1(n15721), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11612) );
  INV_X1 U11814 ( .A(n10603), .ZN(n9990) );
  OR2_X1 U11815 ( .A1(n10644), .A2(n10643), .ZN(n11576) );
  AND2_X1 U11816 ( .A1(n10601), .A2(n10600), .ZN(n10602) );
  NAND2_X1 U11817 ( .A1(n10424), .A2(n13439), .ZN(n10425) );
  NOR2_X1 U11818 ( .A1(n10543), .A2(n10542), .ZN(n11517) );
  INV_X1 U11819 ( .A(n11517), .ZN(n10154) );
  NAND2_X1 U11820 ( .A1(n10441), .A2(n13608), .ZN(n10339) );
  AOI21_X1 U11821 ( .B1(n11104), .B2(n11103), .A(n11102), .ZN(n11147) );
  AND2_X1 U11822 ( .A1(n12030), .A2(n12581), .ZN(n12052) );
  AND2_X1 U11823 ( .A1(n12862), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12019) );
  INV_X1 U11824 ( .A(n12022), .ZN(n12014) );
  AND2_X1 U11825 ( .A1(n10146), .A2(n14934), .ZN(n10144) );
  INV_X1 U11826 ( .A(n14958), .ZN(n10140) );
  NAND2_X1 U11827 ( .A1(n10215), .A2(n16158), .ZN(n10214) );
  INV_X1 U11828 ( .A(n12801), .ZN(n10215) );
  AOI22_X1 U11829 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19356), .B1(
        n12114), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12124) );
  AND2_X1 U11830 ( .A1(n12264), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U11831 ( .A1(n13045), .A2(n12033), .ZN(n12037) );
  INV_X1 U11832 ( .A(n9819), .ZN(n12458) );
  NAND2_X1 U11833 ( .A1(n9954), .A2(n19251), .ZN(n12129) );
  INV_X1 U11834 ( .A(n12139), .ZN(n9954) );
  NAND2_X1 U11835 ( .A1(n11874), .A2(n11873), .ZN(n11888) );
  NOR2_X1 U11836 ( .A1(n18789), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11435) );
  AND2_X1 U11837 ( .A1(n11147), .A2(n11145), .ZN(n11158) );
  AND3_X1 U11838 ( .A1(n11668), .A2(n11710), .A3(n11667), .ZN(n13702) );
  AND2_X1 U11839 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n10950), .ZN(
        n10951) );
  INV_X1 U11840 ( .A(n10949), .ZN(n10950) );
  AND2_X1 U11841 ( .A1(n10027), .A2(n10028), .ZN(n10026) );
  INV_X1 U11842 ( .A(n14418), .ZN(n10027) );
  AND2_X1 U11843 ( .A1(n14472), .A2(n14424), .ZN(n10028) );
  INV_X1 U11844 ( .A(n11058), .ZN(n11090) );
  NOR2_X1 U11845 ( .A1(n10401), .A2(n20718), .ZN(n11058) );
  INV_X1 U11846 ( .A(n13824), .ZN(n10024) );
  NOR2_X1 U11847 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n10847) );
  NOR2_X1 U11848 ( .A1(n10064), .A2(n14342), .ZN(n10063) );
  INV_X1 U11849 ( .A(n14329), .ZN(n10064) );
  INV_X1 U11850 ( .A(n15805), .ZN(n10188) );
  NAND2_X1 U11851 ( .A1(n10055), .A2(n14384), .ZN(n10054) );
  INV_X1 U11852 ( .A(n11708), .ZN(n10055) );
  INV_X1 U11853 ( .A(n14434), .ZN(n10056) );
  OR2_X1 U11854 ( .A1(n9820), .A2(n15844), .ZN(n14599) );
  OR2_X1 U11855 ( .A1(n15928), .A2(n13702), .ZN(n13700) );
  INV_X1 U11856 ( .A(n13462), .ZN(n10060) );
  NAND2_X1 U11857 ( .A1(n11647), .A2(n11646), .ZN(n11649) );
  MUX2_X1 U11858 ( .A(n11732), .B(n11681), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11647) );
  OR2_X1 U11859 ( .A1(n10454), .A2(n10453), .ZN(n11528) );
  AND3_X1 U11860 ( .A1(n10478), .A2(n10477), .A3(n10476), .ZN(n10511) );
  OR2_X1 U11861 ( .A1(n10576), .A2(n10575), .ZN(n11545) );
  AND2_X2 U11862 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13330) );
  OR2_X1 U11863 ( .A1(n10486), .A2(n10518), .ZN(n10530) );
  AND2_X1 U11864 ( .A1(n10562), .A2(n20707), .ZN(n20401) );
  NAND2_X1 U11865 ( .A1(n10490), .A2(n10489), .ZN(n20193) );
  AOI22_X1 U11866 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10680), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U11867 ( .A1(n11143), .A2(n11585), .ZN(n11151) );
  NAND2_X1 U11868 ( .A1(n10566), .A2(n10565), .ZN(n11148) );
  NAND2_X1 U11869 ( .A1(n10205), .A2(n11987), .ZN(n10130) );
  NAND2_X1 U11870 ( .A1(n11839), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11840) );
  NAND2_X1 U11871 ( .A1(n19949), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11853) );
  OR2_X1 U11872 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n11946), .ZN(n12358) );
  INV_X1 U11873 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10080) );
  NOR2_X1 U11874 ( .A1(n10074), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10073) );
  INV_X1 U11875 ( .A(n11941), .ZN(n10074) );
  NAND2_X1 U11876 ( .A1(n10072), .A2(n10071), .ZN(n12277) );
  AND2_X1 U11877 ( .A1(n13399), .A2(n12509), .ZN(n10071) );
  NOR2_X1 U11878 ( .A1(n10078), .A2(n12224), .ZN(n10077) );
  INV_X1 U11879 ( .A(n12229), .ZN(n10078) );
  OR2_X1 U11880 ( .A1(n11906), .A2(n11905), .ZN(n12199) );
  NAND2_X1 U11881 ( .A1(n12025), .A2(n12024), .ZN(n12053) );
  NAND2_X1 U11882 ( .A1(n13048), .A2(n12455), .ZN(n12024) );
  NAND2_X1 U11883 ( .A1(n12046), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12048) );
  CLKBUF_X3 U11884 ( .A(n12000), .Z(n14257) );
  NAND2_X1 U11885 ( .A1(n9890), .A2(n14780), .ZN(n10094) );
  NAND2_X1 U11886 ( .A1(n10093), .A2(n9890), .ZN(n10092) );
  OR2_X1 U11887 ( .A1(n10100), .A2(n16065), .ZN(n10099) );
  NOR2_X1 U11888 ( .A1(n15186), .A2(n10122), .ZN(n12751) );
  NAND2_X1 U11889 ( .A1(n10101), .A2(n14790), .ZN(n10100) );
  INV_X1 U11890 ( .A(n16069), .ZN(n10101) );
  NOR2_X1 U11891 ( .A1(n16230), .A2(n10124), .ZN(n10123) );
  INV_X1 U11892 ( .A(n15273), .ZN(n10124) );
  NOR2_X1 U11893 ( .A1(n14776), .A2(n14765), .ZN(n10116) );
  NOR2_X1 U11894 ( .A1(n18930), .A2(n10016), .ZN(n10015) );
  INV_X1 U11895 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10016) );
  INV_X1 U11896 ( .A(n15492), .ZN(n10014) );
  INV_X1 U11897 ( .A(n13855), .ZN(n13859) );
  INV_X1 U11898 ( .A(n13849), .ZN(n13851) );
  NOR2_X1 U11899 ( .A1(n12348), .A2(n9895), .ZN(n9974) );
  AND2_X1 U11900 ( .A1(n14962), .A2(n10136), .ZN(n10135) );
  AND2_X1 U11901 ( .A1(n14959), .A2(n10138), .ZN(n10136) );
  NOR2_X1 U11902 ( .A1(n10140), .A2(n10139), .ZN(n10138) );
  INV_X1 U11903 ( .A(n15232), .ZN(n10139) );
  NOR2_X1 U11904 ( .A1(n14976), .A2(n12326), .ZN(n12327) );
  INV_X1 U11905 ( .A(n14964), .ZN(n12328) );
  AND2_X1 U11906 ( .A1(n15017), .A2(n15019), .ZN(n14959) );
  AND2_X1 U11907 ( .A1(n15238), .A2(n16197), .ZN(n10128) );
  AND2_X1 U11908 ( .A1(n10128), .A2(n16181), .ZN(n10127) );
  INV_X1 U11909 ( .A(n13873), .ZN(n13965) );
  NAND2_X1 U11910 ( .A1(n12220), .A2(n12219), .ZN(n12790) );
  OR2_X1 U11911 ( .A1(n12218), .A2(n12217), .ZN(n12220) );
  AND4_X1 U11912 ( .A1(n11930), .A2(n11929), .A3(n11928), .A4(n11927), .ZN(
        n11936) );
  AND4_X1 U11913 ( .A1(n11926), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11937) );
  OAI21_X1 U11914 ( .B1(n10209), .B2(n10208), .A(n19976), .ZN(n12179) );
  AND3_X1 U11915 ( .A1(n12412), .A2(n12409), .A3(n12456), .ZN(n12452) );
  OAI21_X1 U11916 ( .B1(n12584), .B2(n12056), .A(n19971), .ZN(n12587) );
  NOR2_X1 U11917 ( .A1(n11804), .A2(n11803), .ZN(n12769) );
  OR2_X1 U11918 ( .A1(n14166), .A2(n19272), .ZN(n13039) );
  CLKBUF_X1 U11919 ( .A(n12424), .Z(n15314) );
  INV_X1 U11920 ( .A(n11243), .ZN(n9936) );
  AOI21_X1 U11921 ( .B1(n17152), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A(n9933), .ZN(n9935) );
  INV_X1 U11922 ( .A(n11244), .ZN(n9933) );
  NOR4_X2 U11923 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A4(n18789), .ZN(n11245) );
  NOR2_X1 U11924 ( .A1(n18601), .A2(n11191), .ZN(n11271) );
  NOR2_X1 U11925 ( .A1(n11192), .A2(n16856), .ZN(n11223) );
  NOR2_X1 U11926 ( .A1(n17825), .A2(n10051), .ZN(n10050) );
  INV_X1 U11927 ( .A(n17621), .ZN(n11311) );
  OR2_X1 U11928 ( .A1(n17748), .A2(n11301), .ZN(n9941) );
  INV_X1 U11929 ( .A(n9941), .ZN(n11302) );
  OAI21_X1 U11930 ( .B1(n9857), .B2(n10178), .A(n10177), .ZN(n11299) );
  NAND2_X1 U11931 ( .A1(n17766), .A2(n10179), .ZN(n10177) );
  AND3_X1 U11932 ( .A1(n11488), .A2(n11426), .A3(n11410), .ZN(n11432) );
  NOR2_X1 U11933 ( .A1(n11389), .A2(n11388), .ZN(n15439) );
  INV_X1 U11934 ( .A(n20046), .ZN(n15688) );
  AND2_X1 U11935 ( .A1(n11688), .A2(n11687), .ZN(n14396) );
  NAND2_X1 U11936 ( .A1(n13747), .A2(n9892), .ZN(n15686) );
  AND2_X1 U11937 ( .A1(n11676), .A2(n11675), .ZN(n13746) );
  OAI21_X1 U11938 ( .B1(n11097), .B2(n15543), .A(n11163), .ZN(n13149) );
  AND2_X1 U11939 ( .A1(n20721), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n11094) );
  AND2_X1 U11940 ( .A1(n11061), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13435) );
  AND2_X1 U11941 ( .A1(n10031), .A2(n11784), .ZN(n10029) );
  AND2_X1 U11942 ( .A1(n11022), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11023) );
  NAND2_X1 U11943 ( .A1(n11023), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11062) );
  NOR2_X1 U11944 ( .A1(n10887), .A2(n10886), .ZN(n10888) );
  NOR2_X1 U11945 ( .A1(n10852), .A2(n10851), .ZN(n10853) );
  NAND2_X1 U11946 ( .A1(n10853), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10887) );
  NOR2_X1 U11947 ( .A1(n10829), .A2(n14607), .ZN(n10830) );
  NOR2_X1 U11948 ( .A1(n10783), .A2(n10708), .ZN(n10784) );
  NAND2_X1 U11949 ( .A1(n10784), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10829) );
  NAND2_X1 U11950 ( .A1(n10723), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10783) );
  NOR2_X1 U11951 ( .A1(n10778), .A2(n14398), .ZN(n10723) );
  OR2_X1 U11952 ( .A1(n10763), .A2(n15689), .ZN(n10778) );
  AND2_X1 U11953 ( .A1(n10707), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10739) );
  NOR2_X1 U11954 ( .A1(n10691), .A2(n10690), .ZN(n10707) );
  NAND2_X1 U11955 ( .A1(n10675), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10691) );
  INV_X1 U11956 ( .A(n13584), .ZN(n10021) );
  AND2_X1 U11957 ( .A1(n10647), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10656) );
  NOR2_X1 U11958 ( .A1(n10628), .A2(n20033), .ZN(n10647) );
  AOI21_X1 U11959 ( .B1(n10634), .B2(n10775), .A(n10633), .ZN(n13569) );
  INV_X1 U11960 ( .A(n10632), .ZN(n10633) );
  NAND2_X1 U11961 ( .A1(n10613), .A2(n10612), .ZN(n13568) );
  AND2_X1 U11962 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U11963 ( .A1(n10583), .A2(n10775), .ZN(n10588) );
  NAND2_X1 U11964 ( .A1(n13270), .A2(n10558), .ZN(n13364) );
  OAI21_X1 U11965 ( .B1(n14716), .B2(n10627), .A(n10554), .ZN(n10555) );
  NAND2_X1 U11966 ( .A1(n10557), .A2(n10556), .ZN(n13270) );
  INV_X1 U11967 ( .A(n13267), .ZN(n10557) );
  INV_X1 U11968 ( .A(n13268), .ZN(n10556) );
  NOR2_X1 U11969 ( .A1(n9903), .A2(n11615), .ZN(n9979) );
  AND2_X1 U11970 ( .A1(n14331), .A2(n14316), .ZN(n14318) );
  OR2_X1 U11971 ( .A1(n14356), .A2(n11729), .ZN(n14357) );
  NOR2_X1 U11972 ( .A1(n9820), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10151) );
  NAND2_X1 U11973 ( .A1(n9989), .A2(n9929), .ZN(n9988) );
  INV_X1 U11974 ( .A(n15569), .ZN(n9989) );
  NOR2_X1 U11975 ( .A1(n9836), .A2(n15612), .ZN(n15611) );
  NOR3_X1 U11976 ( .A1(n15668), .A2(n10056), .A3(n11708), .ZN(n14436) );
  OR2_X1 U11977 ( .A1(n9820), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14586) );
  NOR2_X1 U11978 ( .A1(n15668), .A2(n11708), .ZN(n15648) );
  OR2_X1 U11979 ( .A1(n9820), .A2(n11603), .ZN(n14615) );
  NAND2_X1 U11980 ( .A1(n13747), .A2(n9900), .ZN(n15676) );
  AND2_X1 U11981 ( .A1(n13747), .A2(n10068), .ZN(n15674) );
  NAND2_X1 U11982 ( .A1(n13747), .A2(n13746), .ZN(n15696) );
  NOR2_X1 U11983 ( .A1(n11770), .A2(n13618), .ZN(n15888) );
  NOR2_X1 U11984 ( .A1(n15886), .A2(n13620), .ZN(n15825) );
  CLKBUF_X1 U11985 ( .A(n14636), .Z(n15765) );
  NOR2_X1 U11986 ( .A1(n13700), .A2(n13586), .ZN(n13641) );
  AND2_X1 U11987 ( .A1(n13641), .A2(n13640), .ZN(n13747) );
  NAND2_X1 U11988 ( .A1(n10195), .A2(n13734), .ZN(n9987) );
  NOR2_X1 U11989 ( .A1(n10197), .A2(n10196), .ZN(n10195) );
  INV_X1 U11990 ( .A(n11584), .ZN(n10197) );
  AND2_X1 U11991 ( .A1(n11666), .A2(n11665), .ZN(n15929) );
  NAND2_X1 U11992 ( .A1(n10059), .A2(n10058), .ZN(n15928) );
  AND3_X1 U11993 ( .A1(n13579), .A2(n9839), .A3(n15929), .ZN(n10058) );
  NOR2_X1 U11994 ( .A1(n13365), .A2(n10057), .ZN(n15930) );
  NAND2_X1 U11995 ( .A1(n13579), .A2(n9839), .ZN(n10057) );
  AND2_X1 U11996 ( .A1(n15942), .A2(n20718), .ZN(n11787) );
  NAND2_X1 U11997 ( .A1(n10175), .A2(n11550), .ZN(n10174) );
  NOR2_X1 U11998 ( .A1(n11540), .A2(n20146), .ZN(n13380) );
  NAND2_X1 U11999 ( .A1(n10059), .A2(n9926), .ZN(n13463) );
  AND2_X1 U12000 ( .A1(n11652), .A2(n11651), .ZN(n13271) );
  NAND2_X1 U12001 ( .A1(n11761), .A2(n13314), .ZN(n15886) );
  AND2_X1 U12002 ( .A1(n13447), .A2(n9827), .ZN(n13217) );
  AND3_X1 U12003 ( .A1(n10416), .A2(n10388), .A3(n13608), .ZN(n10389) );
  NAND2_X1 U12004 ( .A1(n10456), .A2(n10497), .ZN(n10461) );
  AND2_X1 U12005 ( .A1(n13589), .A2(n14716), .ZN(n20250) );
  INV_X1 U12006 ( .A(n20250), .ZN(n20262) );
  INV_X1 U12007 ( .A(n20453), .ZN(n20596) );
  NAND3_X1 U12008 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20718), .A3(n13595), 
        .ZN(n20179) );
  OR2_X1 U12009 ( .A1(n14716), .A2(n13408), .ZN(n20649) );
  INV_X1 U12010 ( .A(n20257), .ZN(n20657) );
  NAND2_X2 U12011 ( .A1(n15786), .A2(n13594), .ZN(n20186) );
  AND2_X1 U12012 ( .A1(n15536), .A2(n15535), .ZN(n15549) );
  INV_X1 U12013 ( .A(n16312), .ZN(n12459) );
  OR2_X1 U12014 ( .A1(n12423), .A2(n12459), .ZN(n12809) );
  OR2_X1 U12015 ( .A1(n19965), .A2(n12809), .ZN(n12817) );
  XNOR2_X1 U12016 ( .A(n13855), .B(n13858), .ZN(n15986) );
  AND2_X1 U12017 ( .A1(n12285), .A2(n9849), .ZN(n12353) );
  NAND2_X1 U12018 ( .A1(n12343), .A2(n12350), .ZN(n12285) );
  NOR2_X1 U12019 ( .A1(n12345), .A2(n10082), .ZN(n10081) );
  NOR2_X1 U12020 ( .A1(n16041), .A2(n16042), .ZN(n16040) );
  NOR2_X1 U12021 ( .A1(n15497), .A2(n15498), .ZN(n15964) );
  INV_X1 U12022 ( .A(n18849), .ZN(n9996) );
  OR2_X1 U12023 ( .A1(n18856), .A2(n10004), .ZN(n9997) );
  NAND2_X1 U12024 ( .A1(n12299), .A2(n11941), .ZN(n12322) );
  NOR2_X1 U12025 ( .A1(n15492), .A2(n10011), .ZN(n15022) );
  NAND2_X1 U12026 ( .A1(n10012), .A2(n9902), .ZN(n10011) );
  AND2_X1 U12027 ( .A1(n12264), .A2(n11939), .ZN(n11940) );
  INV_X1 U12028 ( .A(n10072), .ZN(n12267) );
  INV_X1 U12029 ( .A(n12108), .ZN(n9956) );
  INV_X1 U12030 ( .A(n12109), .ZN(n9955) );
  NAND2_X1 U12031 ( .A1(n12108), .A2(n12109), .ZN(n12488) );
  NOR2_X1 U12032 ( .A1(n14762), .A2(n12573), .ZN(n14744) );
  OR2_X1 U12033 ( .A1(n13662), .A2(n13661), .ZN(n19085) );
  AND2_X1 U12034 ( .A1(n12488), .A2(n12487), .ZN(n19025) );
  CLKBUF_X2 U12035 ( .A(n12609), .Z(n13988) );
  NOR2_X1 U12036 ( .A1(n14814), .A2(n13882), .ZN(n13991) );
  INV_X1 U12037 ( .A(n14751), .ZN(n14222) );
  NOR2_X1 U12038 ( .A1(n9835), .A2(n12762), .ZN(n14812) );
  NOR3_X1 U12039 ( .A1(n14864), .A2(n10126), .A3(n14851), .ZN(n14833) );
  XNOR2_X1 U12040 ( .A(n14142), .B(n14144), .ZN(n14775) );
  NOR2_X1 U12041 ( .A1(n14864), .A2(n14851), .ZN(n14850) );
  INV_X1 U12042 ( .A(n12751), .ZN(n15145) );
  NOR3_X1 U12043 ( .A1(n15186), .A2(n14881), .A3(n15157), .ZN(n10237) );
  NOR2_X1 U12044 ( .A1(n14797), .A2(n16069), .ZN(n16068) );
  INV_X1 U12045 ( .A(n12582), .ZN(n12583) );
  OR2_X1 U12046 ( .A1(n13676), .A2(n13675), .ZN(n13678) );
  NOR2_X1 U12047 ( .A1(n16211), .A2(n12672), .ZN(n15261) );
  NAND2_X1 U12048 ( .A1(n15274), .A2(n15273), .ZN(n16229) );
  INV_X1 U12049 ( .A(n10117), .ZN(n13720) );
  NOR2_X1 U12050 ( .A1(n10121), .A2(n10120), .ZN(n10119) );
  AND2_X2 U12051 ( .A1(n12026), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12977) );
  AND2_X1 U12052 ( .A1(n12976), .A2(n19977), .ZN(n19197) );
  NOR2_X1 U12053 ( .A1(n12862), .A2(n12863), .ZN(n13480) );
  INV_X1 U12054 ( .A(n12860), .ZN(n15340) );
  NAND2_X1 U12055 ( .A1(n14928), .A2(n9848), .ZN(n14905) );
  AND2_X1 U12056 ( .A1(n14928), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14919) );
  NAND2_X1 U12057 ( .A1(n10116), .A2(n10115), .ZN(n14762) );
  INV_X1 U12058 ( .A(n14760), .ZN(n10115) );
  INV_X1 U12059 ( .A(n10116), .ZN(n14767) );
  NAND2_X1 U12060 ( .A1(n14985), .A2(n9919), .ZN(n15962) );
  AND2_X1 U12061 ( .A1(n14985), .A2(n10017), .ZN(n15963) );
  AND2_X1 U12062 ( .A1(n15147), .A2(n14793), .ZN(n15148) );
  NAND2_X1 U12063 ( .A1(n14985), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14986) );
  NAND2_X1 U12064 ( .A1(n15022), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15012) );
  AND2_X1 U12065 ( .A1(n12545), .A2(n12544), .ZN(n14799) );
  AND2_X1 U12066 ( .A1(n14804), .A2(n10107), .ZN(n14983) );
  AND2_X1 U12067 ( .A1(n12540), .A2(n12539), .ZN(n15007) );
  NAND2_X1 U12068 ( .A1(n14804), .A2(n10109), .ZN(n15008) );
  AND2_X1 U12069 ( .A1(n13916), .A2(n9866), .ZN(n16102) );
  NAND2_X1 U12070 ( .A1(n10014), .A2(n10015), .ZN(n15493) );
  AND2_X1 U12071 ( .A1(n13916), .A2(n9864), .ZN(n16103) );
  AND2_X1 U12072 ( .A1(n13916), .A2(n13915), .ZN(n13918) );
  NAND2_X1 U12073 ( .A1(n15483), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15492) );
  NAND2_X1 U12074 ( .A1(n13943), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15491) );
  NAND2_X1 U12075 ( .A1(n10001), .A2(n9999), .ZN(n15490) );
  NOR2_X1 U12076 ( .A1(n10002), .A2(n10000), .ZN(n9999) );
  NAND2_X1 U12077 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10000) );
  AND2_X1 U12078 ( .A1(n13260), .A2(n13275), .ZN(n16150) );
  OR2_X1 U12079 ( .A1(n10002), .A2(n18994), .ZN(n9998) );
  OR2_X1 U12080 ( .A1(n15486), .A2(n10002), .ZN(n15488) );
  NOR2_X1 U12081 ( .A1(n15486), .A2(n16178), .ZN(n15489) );
  NAND2_X1 U12082 ( .A1(n12782), .A2(n12783), .ZN(n19233) );
  INV_X1 U12083 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13504) );
  NOR2_X1 U12084 ( .A1(n13472), .A2(n13504), .ZN(n15487) );
  NAND2_X1 U12085 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13472) );
  OR2_X1 U12086 ( .A1(n14742), .A2(n13876), .ZN(n13973) );
  NAND2_X1 U12087 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n10222), .ZN(
        n10221) );
  NOR2_X1 U12088 ( .A1(n14910), .A2(n12472), .ZN(n10222) );
  XNOR2_X1 U12089 ( .A(n12355), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14926) );
  NAND2_X1 U12090 ( .A1(n12807), .A2(n9953), .ZN(n14939) );
  AND2_X1 U12091 ( .A1(n9854), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9953) );
  OR3_X1 U12092 ( .A1(n16029), .A2(n13861), .A3(n15102), .ZN(n14933) );
  NOR2_X1 U12093 ( .A1(n14949), .A2(n14784), .ZN(n14785) );
  NAND2_X1 U12094 ( .A1(n12807), .A2(n12806), .ZN(n14980) );
  OAI21_X1 U12095 ( .B1(n15003), .B2(n14961), .A(n9957), .ZN(n14977) );
  AND2_X1 U12096 ( .A1(n15002), .A2(n14993), .ZN(n9957) );
  AOI21_X1 U12097 ( .B1(n15042), .B2(n14958), .A(n14957), .ZN(n15028) );
  NAND2_X1 U12098 ( .A1(n15028), .A2(n15027), .ZN(n15026) );
  NAND2_X1 U12099 ( .A1(n13916), .A2(n9871), .ZN(n15031) );
  AND2_X1 U12100 ( .A1(n12529), .A2(n12528), .ZN(n15030) );
  NAND2_X1 U12101 ( .A1(n13911), .A2(n9841), .ZN(n10133) );
  OR2_X1 U12102 ( .A1(n12282), .A2(n12275), .ZN(n10134) );
  NAND2_X1 U12103 ( .A1(n13914), .A2(n13923), .ZN(n15250) );
  AND2_X1 U12104 ( .A1(n9868), .A2(n16141), .ZN(n10111) );
  NOR2_X1 U12105 ( .A1(n13223), .A2(n13224), .ZN(n13261) );
  AOI21_X1 U12106 ( .B1(n19230), .B2(n19231), .A(n12250), .ZN(n15284) );
  NOR2_X1 U12107 ( .A1(n10118), .A2(n10121), .ZN(n19031) );
  INV_X1 U12108 ( .A(n13501), .ZN(n10118) );
  OR2_X1 U12109 ( .A1(n12608), .A2(n12611), .ZN(n13073) );
  AOI21_X1 U12110 ( .B1(n12112), .B2(n13089), .A(n13027), .ZN(n13037) );
  INV_X1 U12111 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11798) );
  NOR2_X2 U12112 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16280) );
  OR2_X1 U12113 ( .A1(n12466), .A2(n12465), .ZN(n15306) );
  INV_X1 U12114 ( .A(n13001), .ZN(n16272) );
  CLKBUF_X1 U12115 ( .A(n12402), .Z(n13011) );
  AND2_X1 U12116 ( .A1(n15325), .A2(n19923), .ZN(n15329) );
  NAND2_X1 U12117 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19776), .ZN(n19287) );
  INV_X1 U12118 ( .A(n19287), .ZN(n19291) );
  INV_X1 U12119 ( .A(n19776), .ZN(n19503) );
  NOR2_X2 U12120 ( .A1(n15340), .A2(n15339), .ZN(n19294) );
  NOR2_X2 U12121 ( .A1(n15338), .A2(n15339), .ZN(n19295) );
  INV_X1 U12122 ( .A(n19926), .ZN(n19771) );
  NAND2_X1 U12123 ( .A1(n12442), .A2(n12419), .ZN(n16267) );
  OR2_X1 U12124 ( .A1(n12418), .A2(n12417), .ZN(n12419) );
  NOR3_X1 U12125 ( .A1(n16489), .A2(n17413), .A3(n18604), .ZN(n18585) );
  NOR2_X1 U12126 ( .A1(n16525), .A2(n16524), .ZN(n16523) );
  NOR2_X1 U12127 ( .A1(n17486), .A2(n16545), .ZN(n16544) );
  NOR2_X1 U12128 ( .A1(n17538), .A2(n16588), .ZN(n16587) );
  NOR2_X1 U12129 ( .A1(n16609), .A2(n16608), .ZN(n16607) );
  OR2_X1 U12130 ( .A1(n16339), .A2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10047) );
  NAND2_X1 U12131 ( .A1(n16339), .A2(n10045), .ZN(n10044) );
  NOR2_X1 U12132 ( .A1(n10046), .A2(n10052), .ZN(n10045) );
  NOR2_X2 U12133 ( .A1(n11337), .A2(n11336), .ZN(n17203) );
  AND2_X1 U12134 ( .A1(n11272), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11221) );
  NOR2_X1 U12135 ( .A1(n17414), .A2(n17350), .ZN(n17381) );
  NAND2_X1 U12136 ( .A1(n17611), .A2(n9846), .ZN(n17559) );
  NOR2_X1 U12137 ( .A1(n17591), .A2(n10037), .ZN(n10036) );
  INV_X1 U12138 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U12139 ( .A1(n17611), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17589) );
  NOR2_X1 U12140 ( .A1(n17624), .A2(n17623), .ZN(n17611) );
  AND3_X1 U12141 ( .A1(n10040), .A2(n10039), .A3(n10041), .ZN(n17666) );
  INV_X1 U12142 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17719) );
  NOR2_X1 U12143 ( .A1(n17777), .A2(n17776), .ZN(n17768) );
  AND2_X1 U12144 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17792) );
  NAND2_X1 U12145 ( .A1(n17791), .A2(n17830), .ZN(n17707) );
  AND2_X1 U12146 ( .A1(n17512), .A2(n17841), .ZN(n17843) );
  NAND2_X1 U12147 ( .A1(n10160), .A2(n10159), .ZN(n10157) );
  NOR2_X1 U12148 ( .A1(n10165), .A2(n17878), .ZN(n10161) );
  NAND2_X1 U12149 ( .A1(n11312), .A2(n10159), .ZN(n10156) );
  NOR2_X1 U12150 ( .A1(n10158), .A2(n11312), .ZN(n17514) );
  AND2_X1 U12151 ( .A1(n17576), .A2(n11310), .ZN(n17525) );
  OR3_X1 U12152 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17555), .ZN(n11309) );
  NOR2_X1 U12153 ( .A1(n17734), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17604) );
  NOR2_X1 U12154 ( .A1(n18021), .A2(n16353), .ZN(n17891) );
  INV_X1 U12155 ( .A(n18021), .ZN(n17997) );
  OAI21_X1 U12156 ( .B1(n18593), .B2(n18606), .A(n18592), .ZN(n18615) );
  NAND2_X1 U12157 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17639), .ZN(
        n18021) );
  NOR2_X1 U12158 ( .A1(n11347), .A2(n11346), .ZN(n11487) );
  INV_X1 U12159 ( .A(n16471), .ZN(n18586) );
  INV_X1 U12160 ( .A(n11286), .ZN(n10194) );
  INV_X1 U12161 ( .A(n18613), .ZN(n17936) );
  NAND2_X1 U12162 ( .A1(n15585), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17829) );
  NOR2_X1 U12163 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18156), .ZN(n18452) );
  NOR2_X1 U12164 ( .A1(n11409), .A2(n11408), .ZN(n18171) );
  INV_X1 U12165 ( .A(n15439), .ZN(n18176) );
  OAI22_X1 U12166 ( .A1(n18582), .A2(n18017), .B1(n12833), .B2(n18588), .ZN(
        n18638) );
  OR2_X1 U12167 ( .A1(n12946), .A2(n13128), .ZN(n12971) );
  OR2_X1 U12168 ( .A1(n13451), .A2(n13450), .ZN(n15630) );
  INV_X1 U12169 ( .A(n20067), .ZN(n20049) );
  AND2_X1 U12170 ( .A1(n15629), .A2(n13441), .ZN(n20053) );
  AND2_X1 U12171 ( .A1(n15629), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20024) );
  INV_X1 U12172 ( .A(n20053), .ZN(n20063) );
  AND3_X1 U12173 ( .A1(n13449), .A2(n13444), .A3(n13445), .ZN(n20067) );
  NAND2_X2 U12174 ( .A1(n13132), .A2(n13131), .ZN(n20078) );
  OR2_X1 U12175 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  OR2_X1 U12176 ( .A1(n13145), .A2(n13128), .ZN(n13132) );
  INV_X1 U12177 ( .A(n14493), .ZN(n14488) );
  OR2_X1 U12178 ( .A1(n14495), .A2(n13283), .ZN(n13772) );
  INV_X1 U12179 ( .A(n13772), .ZN(n14504) );
  AND2_X1 U12180 ( .A1(n13156), .A2(n15537), .ZN(n20082) );
  INV_X1 U12181 ( .A(n20080), .ZN(n20801) );
  AND2_X1 U12182 ( .A1(n13255), .A2(n20156), .ZN(n20121) );
  INV_X1 U12183 ( .A(n20121), .ZN(n13257) );
  AND2_X1 U12184 ( .A1(n9860), .A2(n14328), .ZN(n14536) );
  AND2_X1 U12185 ( .A1(n14381), .A2(n14433), .ZN(n15638) );
  INV_X1 U12186 ( .A(n15664), .ZN(n15738) );
  CLKBUF_X1 U12187 ( .A(n13304), .Z(n13305) );
  INV_X1 U12188 ( .A(n20127), .ZN(n19996) );
  INV_X1 U12189 ( .A(n15790), .ZN(n20125) );
  INV_X1 U12190 ( .A(n11615), .ZN(n9978) );
  INV_X1 U12191 ( .A(n15906), .ZN(n15927) );
  INV_X1 U12192 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20570) );
  CLKBUF_X1 U12193 ( .A(n10502), .Z(n10503) );
  INV_X1 U12194 ( .A(n9982), .ZN(n20789) );
  INV_X1 U12195 ( .A(n13337), .ZN(n9983) );
  INV_X1 U12196 ( .A(n15551), .ZN(n20786) );
  INV_X1 U12197 ( .A(n20244), .ZN(n20239) );
  OAI21_X1 U12198 ( .B1(n20306), .B2(n20290), .A(n20606), .ZN(n20308) );
  NOR2_X2 U12199 ( .A1(n20262), .A2(n20499), .ZN(n20307) );
  OR2_X1 U12200 ( .A1(n20368), .A2(n20596), .ZN(n20360) );
  INV_X1 U12201 ( .A(n20360), .ZN(n20396) );
  OAI211_X1 U12202 ( .C1(n20424), .C2(n20537), .A(n20460), .B(n20408), .ZN(
        n20426) );
  INV_X1 U12203 ( .A(n20464), .ZN(n20485) );
  NOR2_X2 U12204 ( .A1(n20500), .A2(n20569), .ZN(n20484) );
  OAI211_X1 U12205 ( .C1(n20557), .C2(n20537), .A(n20606), .B(n20536), .ZN(
        n20565) );
  INV_X1 U12206 ( .A(n20561), .ZN(n20592) );
  INV_X1 U12207 ( .A(n20682), .ZN(n20624) );
  INV_X1 U12208 ( .A(n20683), .ZN(n20625) );
  OAI211_X1 U12209 ( .C1(n20636), .C2(n20607), .A(n20606), .B(n20605), .ZN(
        n20639) );
  INV_X1 U12210 ( .A(n20708), .ZN(n20637) );
  INV_X1 U12211 ( .A(n20540), .ZN(n20647) );
  INV_X1 U12212 ( .A(n20543), .ZN(n20664) );
  INV_X1 U12213 ( .A(n20549), .ZN(n20676) );
  INV_X1 U12214 ( .A(n20555), .ZN(n20689) );
  INV_X1 U12215 ( .A(n20560), .ZN(n20698) );
  OR2_X1 U12216 ( .A1(n20649), .A2(n20499), .ZN(n20715) );
  NOR2_X1 U12217 ( .A1(n13155), .A2(n20537), .ZN(n15551) );
  INV_X1 U12218 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20717) );
  INV_X1 U12219 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20537) );
  INV_X1 U12220 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20718) );
  NAND2_X1 U12221 ( .A1(n12031), .A2(n13045), .ZN(n19984) );
  OR2_X1 U12222 ( .A1(n15985), .A2(n15968), .ZN(n15973) );
  NOR2_X1 U12223 ( .A1(n15973), .A2(n15972), .ZN(n15974) );
  NOR2_X1 U12224 ( .A1(n15983), .A2(n19046), .ZN(n9994) );
  NAND2_X1 U12225 ( .A1(n12370), .A2(n13855), .ZN(n15999) );
  OAI21_X1 U12226 ( .B1(n10006), .B2(n10004), .A(n10003), .ZN(n16016) );
  NAND2_X1 U12227 ( .A1(n10008), .A2(n10005), .ZN(n10003) );
  NOR2_X1 U12229 ( .A1(n16040), .A2(n10004), .ZN(n16026) );
  INV_X1 U12230 ( .A(n9997), .ZN(n18848) );
  AND2_X1 U12231 ( .A1(n14794), .A2(n15149), .ZN(n18847) );
  AOI21_X1 U12232 ( .B1(n18881), .B2(n18882), .A(n10004), .ZN(n18868) );
  AND2_X1 U12233 ( .A1(n13486), .A2(n16311), .ZN(n19069) );
  OR2_X1 U12234 ( .A1(n19053), .A2(n19971), .ZN(n19049) );
  INV_X1 U12235 ( .A(n19049), .ZN(n19081) );
  INV_X1 U12236 ( .A(n19046), .ZN(n19075) );
  OAI21_X1 U12237 ( .B1(n14744), .B2(n14743), .A(n14742), .ZN(n15989) );
  OR2_X1 U12238 ( .A1(n13541), .A2(n13540), .ZN(n13542) );
  OR2_X1 U12239 ( .A1(n12640), .A2(n12639), .ZN(n19108) );
  NOR2_X1 U12240 ( .A1(n10096), .A2(n9850), .ZN(n10095) );
  INV_X1 U12241 ( .A(n19943), .ZN(n19361) );
  INV_X1 U12242 ( .A(n19117), .ZN(n19107) );
  AND2_X2 U12243 ( .A1(n13015), .A2(n19829), .ZN(n19121) );
  NOR2_X1 U12244 ( .A1(n14859), .A2(n14092), .ZN(n14781) );
  OR2_X1 U12245 ( .A1(n13051), .A2(n13050), .ZN(n13052) );
  NOR2_X1 U12246 ( .A1(n19176), .A2(n19187), .ZN(n19172) );
  INV_X1 U12247 ( .A(n19191), .ZN(n19176) );
  AND2_X1 U12248 ( .A1(n19162), .A2(n13064), .ZN(n19187) );
  INV_X1 U12249 ( .A(n19162), .ZN(n19186) );
  INV_X1 U12250 ( .A(n19164), .ZN(n19195) );
  NOR2_X1 U12251 ( .A1(n19197), .A2(n13117), .ZN(n19196) );
  BUF_X1 U12252 ( .A(n19196), .Z(n19227) );
  XNOR2_X1 U12253 ( .A(n13469), .B(n13468), .ZN(n13964) );
  NAND2_X1 U12254 ( .A1(n16159), .A2(n16158), .ZN(n16157) );
  NAND2_X1 U12255 ( .A1(n15269), .A2(n12801), .ZN(n16159) );
  INV_X1 U12256 ( .A(n16170), .ZN(n19247) );
  NAND2_X1 U12257 ( .A1(n12869), .A2(n12822), .ZN(n16179) );
  AND2_X1 U12258 ( .A1(n16179), .A2(n12954), .ZN(n16170) );
  INV_X1 U12259 ( .A(n16179), .ZN(n19239) );
  AOI21_X1 U12260 ( .B1(n15969), .B2(n19257), .A(n13992), .ZN(n13993) );
  XNOR2_X1 U12261 ( .A(n13963), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n13997) );
  NOR2_X1 U12262 ( .A1(n10221), .A2(n13984), .ZN(n10220) );
  XNOR2_X1 U12263 ( .A(n13961), .B(n10238), .ZN(n13999) );
  XNOR2_X1 U12264 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n13960), .ZN(
        n10238) );
  NAND2_X1 U12265 ( .A1(n13954), .A2(n13953), .ZN(n13961) );
  NAND2_X1 U12266 ( .A1(n14917), .A2(n9972), .ZN(n9967) );
  NAND2_X1 U12267 ( .A1(n14917), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14916) );
  NOR2_X1 U12268 ( .A1(n14942), .A2(n12348), .ZN(n15111) );
  NOR2_X1 U12269 ( .A1(n13935), .A2(n12477), .ZN(n15174) );
  OR2_X1 U12270 ( .A1(n15253), .A2(n12275), .ZN(n10141) );
  AND2_X1 U12271 ( .A1(n10147), .A2(n10148), .ZN(n16136) );
  NAND2_X1 U12272 ( .A1(n13914), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16144) );
  NOR2_X1 U12273 ( .A1(n12475), .A2(n15288), .ZN(n16224) );
  NAND2_X1 U12274 ( .A1(n13718), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13717) );
  NAND2_X1 U12275 ( .A1(n9952), .A2(n12791), .ZN(n13718) );
  INV_X1 U12276 ( .A(n19257), .ZN(n16215) );
  INV_X1 U12277 ( .A(n16253), .ZN(n19255) );
  NAND2_X1 U12278 ( .A1(n9966), .A2(n13503), .ZN(n13422) );
  NAND2_X1 U12279 ( .A1(n15202), .A2(n15204), .ZN(n16257) );
  AND2_X1 U12280 ( .A1(n12810), .A2(n12580), .ZN(n19257) );
  INV_X1 U12281 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19958) );
  OR2_X1 U12282 ( .A1(n13025), .A2(n13021), .ZN(n19952) );
  INV_X1 U12283 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19949) );
  INV_X1 U12284 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16303) );
  XNOR2_X1 U12285 ( .A(n13038), .B(n13037), .ZN(n19943) );
  NAND2_X1 U12286 ( .A1(n16272), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19916) );
  INV_X1 U12287 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13013) );
  INV_X1 U12288 ( .A(n19416), .ZN(n19406) );
  INV_X1 U12289 ( .A(n19443), .ZN(n19446) );
  INV_X1 U12290 ( .A(n19464), .ZN(n19474) );
  NOR2_X1 U12291 ( .A1(n19499), .A2(n19684), .ZN(n19490) );
  INV_X1 U12292 ( .A(n19523), .ZN(n19513) );
  AND2_X1 U12293 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13090), .ZN(
        n19534) );
  OAI21_X1 U12294 ( .B1(n19597), .B2(n19613), .A(n19776), .ZN(n19615) );
  INV_X1 U12295 ( .A(n19787), .ZN(n19741) );
  INV_X1 U12296 ( .A(n19756), .ZN(n19758) );
  OAI21_X1 U12297 ( .B1(n19738), .B2(n19737), .A(n19736), .ZN(n19760) );
  INV_X1 U12298 ( .A(n19697), .ZN(n19778) );
  AND2_X1 U12299 ( .A1(n16274), .A2(n19291), .ZN(n19769) );
  AND2_X1 U12300 ( .A1(n19976), .A2(n19291), .ZN(n19782) );
  INV_X1 U12301 ( .A(n19707), .ZN(n19796) );
  INV_X1 U12302 ( .A(n19711), .ZN(n19802) );
  INV_X1 U12303 ( .A(n19715), .ZN(n19808) );
  INV_X1 U12304 ( .A(n19719), .ZN(n19814) );
  INV_X1 U12305 ( .A(n19764), .ZN(n19822) );
  AND2_X1 U12306 ( .A1(n16317), .A2(n16316), .ZN(n19836) );
  INV_X1 U12307 ( .A(n19836), .ZN(n16325) );
  NAND2_X1 U12308 ( .A1(n18824), .A2(n18157), .ZN(n18822) );
  INV_X1 U12309 ( .A(n18810), .ZN(n18820) );
  NAND2_X1 U12310 ( .A1(n18642), .A2(n18586), .ZN(n17414) );
  NOR2_X1 U12311 ( .A1(n18585), .A2(n17414), .ZN(n18824) );
  NAND2_X1 U12312 ( .A1(n18642), .A2(n18638), .ZN(n16474) );
  NOR2_X1 U12313 ( .A1(n16568), .A2(n16567), .ZN(n16566) );
  NOR2_X1 U12314 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16614), .ZN(n16597) );
  INV_X1 U12315 ( .A(n16828), .ZN(n16864) );
  NOR2_X1 U12316 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16759), .ZN(n16738) );
  NOR2_X1 U12317 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16803), .ZN(n16787) );
  NOR2_X2 U12318 ( .A1(n18822), .A2(n18644), .ZN(n16828) );
  INV_X1 U12319 ( .A(n16877), .ZN(n16868) );
  OAI211_X1 U12320 ( .C1(n18652), .C2(n18645), .A(n16823), .B(n18819), .ZN(
        n16877) );
  NOR2_X1 U12321 ( .A1(n16593), .A2(n16940), .ZN(n16946) );
  NOR2_X1 U12322 ( .A1(n17017), .A2(n17006), .ZN(n17002) );
  NOR2_X1 U12323 ( .A1(n16762), .A2(n17162), .ZN(n17140) );
  NOR2_X1 U12324 ( .A1(n16821), .A2(n17177), .ZN(n17181) );
  NOR3_X1 U12325 ( .A1(n17367), .A2(n17278), .A3(n17251), .ZN(n17243) );
  NOR3_X1 U12326 ( .A1(n18188), .A2(n17278), .A3(n17419), .ZN(n17270) );
  NAND2_X1 U12327 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17282), .ZN(n17278) );
  AND2_X1 U12328 ( .A1(n18188), .A2(n15587), .ZN(n17283) );
  AND2_X1 U12329 ( .A1(n17313), .A2(n17345), .ZN(n17321) );
  NOR2_X1 U12330 ( .A1(n11199), .A2(n11198), .ZN(n17761) );
  NOR2_X1 U12331 ( .A1(n11209), .A2(n11208), .ZN(n17325) );
  AOI21_X1 U12332 ( .B1(n18642), .B2(n15583), .A(n15582), .ZN(n17342) );
  INV_X1 U12333 ( .A(n17316), .ZN(n17348) );
  NOR2_X1 U12334 ( .A1(n17342), .A2(n15584), .ZN(n17316) );
  CLKBUF_X1 U12335 ( .A(n17377), .Z(n17409) );
  NOR2_X1 U12336 ( .A1(n17476), .A2(n17477), .ZN(n16339) );
  NOR2_X1 U12337 ( .A1(n17508), .A2(n17509), .ZN(n17496) );
  AND2_X1 U12338 ( .A1(n17611), .A2(n10034), .ZN(n17549) );
  AND2_X1 U12339 ( .A1(n9846), .A2(n10035), .ZN(n10034) );
  INV_X1 U12340 ( .A(n17560), .ZN(n10035) );
  NAND2_X1 U12341 ( .A1(n17319), .A2(n17822), .ZN(n17737) );
  INV_X1 U12342 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17670) );
  INV_X1 U12343 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17681) );
  INV_X1 U12344 ( .A(n17739), .ZN(n17717) );
  INV_X1 U12345 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17776) );
  INV_X1 U12346 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17800) );
  INV_X1 U12347 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17816) );
  OAI21_X1 U12348 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18803), .A(n16474), 
        .ZN(n17830) );
  INV_X1 U12349 ( .A(n17818), .ZN(n17834) );
  INV_X1 U12350 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18813) );
  NAND2_X1 U12351 ( .A1(n10204), .A2(n10203), .ZN(n10202) );
  INV_X1 U12352 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18812) );
  AND2_X1 U12353 ( .A1(n11307), .A2(n11306), .ZN(n17610) );
  NAND2_X1 U12354 ( .A1(n10181), .A2(n10180), .ZN(n18065) );
  NOR2_X1 U12355 ( .A1(n9857), .A2(n11294), .ZN(n17767) );
  INV_X1 U12356 ( .A(n17986), .ZN(n18129) );
  INV_X1 U12357 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18628) );
  INV_X1 U12358 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18632) );
  INV_X1 U12359 ( .A(n18787), .ZN(n18790) );
  INV_X1 U12360 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18758) );
  NAND2_X1 U12362 ( .A1(n14282), .A2(n11168), .ZN(n11185) );
  NAND2_X1 U12363 ( .A1(n14557), .A2(n14556), .ZN(n14558) );
  AND2_X1 U12364 ( .A1(n11778), .A2(n11777), .ZN(n11779) );
  AOI211_X1 U12365 ( .C1(n15932), .C2(n14408), .A(n13978), .B(n11769), .ZN(
        n11778) );
  OAI21_X1 U12366 ( .B1(n9995), .B2(n15974), .A(n9993), .ZN(P2_U2825) );
  INV_X1 U12367 ( .A(n15982), .ZN(n9995) );
  NOR2_X1 U12368 ( .A1(n9994), .A2(n15981), .ZN(n9993) );
  AOI21_X1 U12369 ( .B1(n15973), .B2(n15972), .A(n19834), .ZN(n15982) );
  AOI21_X1 U12370 ( .B1(n18896), .B2(n19250), .A(n15025), .ZN(n10089) );
  NAND2_X1 U12371 ( .A1(n10091), .A2(n19242), .ZN(n10090) );
  OR2_X1 U12372 ( .A1(n15218), .A2(n16173), .ZN(n10088) );
  AOI211_X1 U12373 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15068), .A(
        n15067), .B(n15066), .ZN(n15071) );
  OR2_X1 U12374 ( .A1(n16334), .A2(n16333), .ZN(n9938) );
  AOI21_X1 U12375 ( .B1(n9939), .B2(n9811), .A(n9937), .ZN(n15560) );
  OR2_X1 U12376 ( .A1(n15559), .A2(n16329), .ZN(n9937) );
  OR2_X1 U12377 ( .A1(n13743), .A2(n9845), .ZN(n9833) );
  INV_X1 U12378 ( .A(n11895), .ZN(n12246) );
  INV_X2 U12379 ( .A(n15967), .ZN(n10004) );
  AND2_X1 U12380 ( .A1(n9853), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9834) );
  INV_X1 U12381 ( .A(n11234), .ZN(n17147) );
  OR3_X1 U12382 ( .A1(n14864), .A2(n10125), .A3(n14825), .ZN(n9835) );
  OR3_X1 U12383 ( .A1(n15668), .A2(n10054), .A3(n9901), .ZN(n9836) );
  AND2_X1 U12384 ( .A1(n14382), .A2(n9911), .ZN(n9837) );
  AND2_X1 U12385 ( .A1(n12807), .A2(n9834), .ZN(n9838) );
  INV_X1 U12386 ( .A(n12033), .ZN(n12011) );
  NAND2_X1 U12387 ( .A1(n14492), .A2(n10850), .ZN(n14381) );
  INV_X1 U12388 ( .A(n12031), .ZN(n12581) );
  AND2_X1 U12389 ( .A1(n9926), .A2(n10060), .ZN(n9839) );
  NAND2_X1 U12390 ( .A1(n14382), .A2(n10028), .ZN(n14416) );
  INV_X2 U12391 ( .A(n11593), .ZN(n14587) );
  NAND2_X1 U12392 ( .A1(n13912), .A2(n12276), .ZN(n9841) );
  AND2_X1 U12393 ( .A1(n11549), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9842) );
  AND2_X1 U12394 ( .A1(n12254), .A2(n9899), .ZN(n9843) );
  AND2_X1 U12395 ( .A1(n10076), .A2(n10077), .ZN(n9844) );
  NAND2_X1 U12396 ( .A1(n13677), .A2(n13678), .ZN(n14000) );
  OR2_X1 U12397 ( .A1(n9889), .A2(n10024), .ZN(n9845) );
  AND2_X1 U12398 ( .A1(n10036), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9846) );
  AND2_X1 U12399 ( .A1(n9991), .A2(n10653), .ZN(n9847) );
  AND2_X1 U12400 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n9848) );
  INV_X1 U12401 ( .A(n13365), .ZN(n10059) );
  INV_X1 U12402 ( .A(n13310), .ZN(n9981) );
  AND2_X1 U12403 ( .A1(n10081), .A2(n10080), .ZN(n9849) );
  NAND2_X1 U12404 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n9850) );
  AND2_X1 U12405 ( .A1(n9848), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9851) );
  INV_X1 U12406 ( .A(n10168), .ZN(n11629) );
  AND2_X1 U12407 ( .A1(n12301), .A2(n14795), .ZN(n9852) );
  AND2_X1 U12408 ( .A1(n12806), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9853) );
  AND2_X1 U12409 ( .A1(n9834), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9854) );
  AND2_X1 U12410 ( .A1(n13923), .A2(n16196), .ZN(n9855) );
  AND2_X2 U12411 ( .A1(n14265), .A2(n11987), .ZN(n11912) );
  NAND2_X1 U12412 ( .A1(n14636), .A2(n11594), .ZN(n14597) );
  AND2_X1 U12413 ( .A1(n10143), .A2(n10146), .ZN(n9856) );
  NOR2_X1 U12414 ( .A1(n17772), .A2(n18084), .ZN(n9857) );
  NAND2_X1 U12415 ( .A1(n14063), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9858) );
  AND2_X1 U12416 ( .A1(n12285), .A2(n12342), .ZN(n9859) );
  NOR2_X1 U12417 ( .A1(n14381), .A2(n14383), .ZN(n14382) );
  NAND2_X1 U12418 ( .A1(n14353), .A2(n10030), .ZN(n9860) );
  INV_X1 U12419 ( .A(n13439), .ZN(n12958) );
  OR2_X1 U12420 ( .A1(n10603), .A2(n10602), .ZN(n9861) );
  OR2_X1 U12421 ( .A1(n9820), .A2(n15907), .ZN(n9862) );
  INV_X1 U12422 ( .A(n9975), .ZN(n14942) );
  AND2_X1 U12423 ( .A1(n12807), .A2(n9853), .ZN(n14967) );
  AND2_X1 U12424 ( .A1(n14382), .A2(n14424), .ZN(n14422) );
  NOR2_X1 U12425 ( .A1(n11233), .A2(n11232), .ZN(n17349) );
  INV_X1 U12426 ( .A(n17349), .ZN(n11283) );
  AND4_X1 U12427 ( .A1(n10305), .A2(n10304), .A3(n10303), .A4(n10302), .ZN(
        n9863) );
  INV_X1 U12428 ( .A(n13029), .ZN(n16283) );
  NAND2_X1 U12430 ( .A1(n10147), .A2(n12263), .ZN(n13930) );
  AND2_X1 U12431 ( .A1(n13403), .A2(n13915), .ZN(n9864) );
  AND2_X1 U12432 ( .A1(n16149), .A2(n13275), .ZN(n9865) );
  AND2_X1 U12433 ( .A1(n9864), .A2(n16104), .ZN(n9866) );
  NAND2_X1 U12434 ( .A1(n14578), .A2(n14593), .ZN(n14577) );
  INV_X1 U12435 ( .A(n12129), .ZN(n12192) );
  AND4_X1 U12436 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n9867) );
  AND2_X1 U12437 ( .A1(n9865), .A2(n13359), .ZN(n9868) );
  NAND2_X1 U12438 ( .A1(n12807), .A2(n9854), .ZN(n9869) );
  AND2_X1 U12439 ( .A1(n15744), .A2(n11598), .ZN(n9870) );
  INV_X1 U12440 ( .A(n16158), .ZN(n10218) );
  XNOR2_X1 U12441 ( .A(n12802), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16158) );
  NAND2_X1 U12442 ( .A1(n12977), .A2(n12031), .ZN(n12045) );
  AND2_X1 U12443 ( .A1(n9866), .A2(n13546), .ZN(n9871) );
  OR2_X1 U12444 ( .A1(n11302), .A2(n17642), .ZN(n9872) );
  AND2_X1 U12445 ( .A1(n10129), .A2(n10130), .ZN(n9873) );
  AND2_X1 U12446 ( .A1(n11592), .A2(n9862), .ZN(n9874) );
  NAND2_X1 U12447 ( .A1(n17609), .A2(n17702), .ZN(n17576) );
  NAND2_X1 U12448 ( .A1(n12808), .A2(n12479), .ZN(n14913) );
  OR2_X1 U12449 ( .A1(n14174), .A2(n14173), .ZN(n9875) );
  NOR2_X1 U12450 ( .A1(n11284), .A2(n18112), .ZN(n11285) );
  AND2_X1 U12451 ( .A1(n14382), .A2(n10026), .ZN(n14368) );
  AND2_X1 U12452 ( .A1(n15294), .A2(n12790), .ZN(n9876) );
  AND2_X1 U12453 ( .A1(n13914), .A2(n9855), .ZN(n9877) );
  OR2_X1 U12454 ( .A1(n12371), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9878) );
  AND2_X1 U12455 ( .A1(n10141), .A2(n12276), .ZN(n9879) );
  AND2_X1 U12456 ( .A1(n9980), .A2(n9978), .ZN(n9880) );
  INV_X1 U12457 ( .A(n12112), .ZN(n13910) );
  AND2_X1 U12458 ( .A1(n10218), .A2(n12804), .ZN(n9881) );
  AND2_X1 U12459 ( .A1(n10216), .A2(n12805), .ZN(n9882) );
  INV_X1 U12460 ( .A(n12759), .ZN(n13989) );
  NOR2_X1 U12461 ( .A1(n10237), .A2(n15158), .ZN(n9883) );
  AND2_X1 U12462 ( .A1(n10014), .A2(n10012), .ZN(n9884) );
  AND2_X1 U12463 ( .A1(n14985), .A2(n10018), .ZN(n9885) );
  OR2_X1 U12464 ( .A1(n14357), .A2(n10062), .ZN(n9886) );
  NOR3_X1 U12465 ( .A1(n13581), .A2(n13630), .A3(n10021), .ZN(n13582) );
  NOR2_X1 U12466 ( .A1(n15222), .A2(n13680), .ZN(n13679) );
  OR2_X1 U12467 ( .A1(n14797), .A2(n10100), .ZN(n14789) );
  NOR2_X1 U12468 ( .A1(n13743), .A2(n10782), .ZN(n13775) );
  AND2_X1 U12469 ( .A1(n15237), .A2(n10128), .ZN(n16180) );
  NAND2_X1 U12470 ( .A1(n13364), .A2(n13363), .ZN(n13362) );
  NOR2_X1 U12471 ( .A1(n15012), .A2(n14996), .ZN(n14985) );
  NOR2_X1 U12472 ( .A1(n15490), .A2(n18972), .ZN(n13943) );
  NOR2_X1 U12473 ( .A1(n15491), .A2(n18955), .ZN(n15483) );
  NOR2_X1 U12474 ( .A1(n15486), .A2(n9998), .ZN(n15056) );
  NOR2_X1 U12475 ( .A1(n15492), .A2(n18930), .ZN(n15482) );
  AND2_X1 U12476 ( .A1(n14804), .A2(n14803), .ZN(n9887) );
  NAND2_X1 U12477 ( .A1(n15237), .A2(n10127), .ZN(n9888) );
  OR2_X1 U12478 ( .A1(n10782), .A2(n10025), .ZN(n9889) );
  INV_X1 U12479 ( .A(n10165), .ZN(n10164) );
  NAND2_X1 U12480 ( .A1(n14118), .A2(n14117), .ZN(n9890) );
  NOR2_X1 U12481 ( .A1(n13743), .A2(n9889), .ZN(n13774) );
  AND2_X1 U12482 ( .A1(n13582), .A2(n13636), .ZN(n13635) );
  OR2_X1 U12483 ( .A1(n15186), .A2(n14881), .ZN(n9891) );
  AND2_X1 U12484 ( .A1(n13746), .A2(n10070), .ZN(n9892) );
  NAND2_X1 U12485 ( .A1(n13734), .A2(n11584), .ZN(n13757) );
  INV_X1 U12486 ( .A(n12260), .ZN(n10076) );
  NAND2_X1 U12487 ( .A1(n9987), .A2(n11592), .ZN(n13782) );
  NAND2_X1 U12488 ( .A1(n13447), .A2(n11531), .ZN(n11585) );
  AND3_X1 U12489 ( .A1(n10020), .A2(n10613), .A3(n10612), .ZN(n13567) );
  NAND2_X1 U12491 ( .A1(n14775), .A2(n14774), .ZN(n14773) );
  NAND2_X1 U12492 ( .A1(n10406), .A2(n10364), .ZN(n10168) );
  NAND2_X1 U12493 ( .A1(n12023), .A2(n12410), .ZN(n12409) );
  NOR2_X1 U12494 ( .A1(n14781), .A2(n14780), .ZN(n9893) );
  OR3_X1 U12495 ( .A1(n15668), .A2(n10054), .A3(n10056), .ZN(n9894) );
  AND2_X1 U12496 ( .A1(n12354), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9895) );
  NAND2_X1 U12497 ( .A1(n12236), .A2(n12235), .ZN(n12247) );
  OR2_X1 U12498 ( .A1(n14864), .A2(n10125), .ZN(n9896) );
  AND2_X1 U12499 ( .A1(n10148), .A2(n16138), .ZN(n9897) );
  AND2_X1 U12500 ( .A1(n10625), .A2(n10624), .ZN(n9898) );
  AND2_X1 U12501 ( .A1(n10578), .A2(n10577), .ZN(n13408) );
  INV_X1 U12502 ( .A(n13408), .ZN(n10580) );
  AND2_X1 U12503 ( .A1(n16151), .A2(n16153), .ZN(n9899) );
  AND2_X1 U12504 ( .A1(n10068), .A2(n15673), .ZN(n9900) );
  INV_X1 U12505 ( .A(n10653), .ZN(n9992) );
  OR2_X1 U12506 ( .A1(n10056), .A2(n14425), .ZN(n9901) );
  AND2_X1 U12507 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9902) );
  OR2_X1 U12508 ( .A1(n9820), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9903) );
  OR2_X1 U12509 ( .A1(n11887), .A2(n11886), .ZN(n12781) );
  INV_X1 U12510 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18994) );
  INV_X1 U12511 ( .A(n17702), .ZN(n17734) );
  NAND2_X1 U12512 ( .A1(n11298), .A2(n16354), .ZN(n17702) );
  AND2_X1 U12513 ( .A1(n10123), .A2(n13934), .ZN(n9904) );
  NOR2_X1 U12514 ( .A1(n12597), .A2(n12626), .ZN(n9905) );
  AND2_X1 U12515 ( .A1(n10127), .A2(n15220), .ZN(n9906) );
  AND2_X1 U12516 ( .A1(n10073), .A2(n9852), .ZN(n9907) );
  NOR2_X1 U12517 ( .A1(n13457), .A2(n9984), .ZN(n9908) );
  AND2_X1 U12518 ( .A1(n10107), .A2(n14982), .ZN(n9909) );
  AND2_X1 U12519 ( .A1(n9997), .A2(n9996), .ZN(n9910) );
  AND2_X1 U12520 ( .A1(n10956), .A2(n10026), .ZN(n9911) );
  AND2_X1 U12521 ( .A1(n10073), .A2(n12301), .ZN(n9912) );
  INV_X1 U12522 ( .A(n12977), .ZN(n12376) );
  OAI22_X1 U12523 ( .A1(n13964), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n13470), 
        .B2(n13969), .ZN(n15967) );
  INV_X1 U12524 ( .A(n10004), .ZN(n10005) );
  OR2_X1 U12525 ( .A1(n13608), .A2(n20721), .ZN(n9913) );
  NOR2_X1 U12526 ( .A1(n14919), .A2(n14918), .ZN(n9914) );
  NAND2_X1 U12527 ( .A1(n10097), .A2(n19028), .ZN(n13258) );
  NAND2_X1 U12528 ( .A1(n10166), .A2(n13447), .ZN(n11097) );
  NAND2_X1 U12529 ( .A1(n12629), .A2(n12628), .ZN(n15274) );
  AND2_X1 U12530 ( .A1(n12820), .A2(n12584), .ZN(n19242) );
  AND2_X1 U12531 ( .A1(n15274), .A2(n10123), .ZN(n13933) );
  AND2_X1 U12532 ( .A1(n13260), .A2(n10111), .ZN(n13394) );
  AND2_X1 U12533 ( .A1(n13260), .A2(n9868), .ZN(n13357) );
  AND2_X1 U12534 ( .A1(n13260), .A2(n9865), .ZN(n13356) );
  AND2_X1 U12535 ( .A1(n10059), .A2(n9839), .ZN(n9915) );
  AND2_X1 U12536 ( .A1(n16339), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9916) );
  INV_X1 U12537 ( .A(n16353), .ZN(n9943) );
  INV_X1 U12538 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n9961) );
  INV_X1 U12539 ( .A(n14200), .ZN(n10102) );
  INV_X1 U12540 ( .A(n20283), .ZN(n9986) );
  AND2_X1 U12541 ( .A1(n13261), .A2(n13262), .ZN(n13260) );
  INV_X1 U12542 ( .A(n12342), .ZN(n10082) );
  AND2_X1 U12543 ( .A1(n13677), .A2(n10098), .ZN(n9917) );
  AND2_X1 U12544 ( .A1(n15237), .A2(n15238), .ZN(n15239) );
  AND2_X1 U12545 ( .A1(n13220), .A2(n13219), .ZN(n19027) );
  NAND2_X1 U12546 ( .A1(n15965), .A2(n10004), .ZN(n9918) );
  AND2_X1 U12547 ( .A1(n10017), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9919) );
  NOR2_X1 U12548 ( .A1(n17767), .A2(n17766), .ZN(n9920) );
  NAND2_X1 U12549 ( .A1(n10560), .A2(n10533), .ZN(n13310) );
  AND2_X1 U12550 ( .A1(n9851), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9921) );
  AND2_X1 U12551 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n9922) );
  AND2_X1 U12552 ( .A1(n14928), .A2(n9851), .ZN(n9923) );
  AND2_X1 U12553 ( .A1(n16339), .A2(n10050), .ZN(n9924) );
  INV_X1 U12554 ( .A(n17777), .ZN(n10040) );
  INV_X1 U12555 ( .A(n14803), .ZN(n10110) );
  INV_X1 U12556 ( .A(n19028), .ZN(n10096) );
  NAND2_X1 U12557 ( .A1(n10832), .A2(n10831), .ZN(n9925) );
  NAND2_X1 U12558 ( .A1(n11656), .A2(n11655), .ZN(n9926) );
  AND2_X1 U12559 ( .A1(n10190), .A2(n10189), .ZN(n9927) );
  INV_X1 U12560 ( .A(n14316), .ZN(n10067) );
  INV_X1 U12561 ( .A(n16232), .ZN(n19016) );
  INV_X1 U12562 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10051) );
  AND2_X1 U12563 ( .A1(n17611), .A2(n10036), .ZN(n9928) );
  AND2_X1 U12564 ( .A1(n14581), .A2(n15835), .ZN(n9929) );
  AND2_X1 U12565 ( .A1(n13470), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13089) );
  INV_X1 U12566 ( .A(n13089), .ZN(n10105) );
  AND2_X1 U12567 ( .A1(n9855), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9930) );
  INV_X1 U12568 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10052) );
  INV_X1 U12569 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10053) );
  OR2_X1 U12570 ( .A1(n15081), .A2(n12472), .ZN(n9931) );
  NAND2_X1 U12571 ( .A1(n15257), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10087) );
  NAND2_X2 U12572 ( .A1(n18821), .A2(n18652), .ZN(n18036) );
  INV_X1 U12573 ( .A(n16798), .ZN(n16818) );
  NOR2_X1 U12574 ( .A1(n16798), .A2(n16505), .ZN(n16620) );
  OAI22_X2 U12575 ( .A1(n20152), .A2(n20184), .B1(n21135), .B2(n20186), .ZN(
        n20660) );
  OAI22_X2 U12576 ( .A1(n21118), .A2(n20186), .B1(n13685), .B2(n20184), .ZN(
        n20666) );
  NAND2_X2 U12577 ( .A1(n15786), .A2(n13593), .ZN(n20184) );
  OAI22_X2 U12578 ( .A1(n20163), .A2(n20184), .B1(n21033), .B2(n20186), .ZN(
        n20672) );
  OAI22_X2 U12579 ( .A1(n20170), .A2(n20186), .B1(n14887), .B2(n20184), .ZN(
        n20678) );
  NOR3_X2 U12580 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18523), .A3(
        n18328), .ZN(n18345) );
  NOR3_X2 U12581 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18523), .A3(
        n18424), .ZN(n18392) );
  NOR3_X2 U12582 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18523), .A3(
        n18284), .ZN(n18302) );
  OAI22_X2 U12583 ( .A1(n14876), .A2(n20184), .B1(n21024), .B2(n20186), .ZN(
        n20691) );
  NOR3_X2 U12584 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18523), .A3(
        n18196), .ZN(n18212) );
  OAI22_X2 U12585 ( .A1(n20957), .A2(n20186), .B1(n16375), .B2(n20184), .ZN(
        n20710) );
  NOR4_X4 U12586 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .A4(n18813), .ZN(n18653) );
  OR2_X1 U12587 ( .A1(n19925), .A2(n19527), .ZN(n19725) );
  OR2_X1 U12588 ( .A1(n19925), .A2(n19952), .ZN(n19683) );
  NAND2_X1 U12589 ( .A1(n19925), .A2(n19952), .ZN(n19422) );
  AND3_X2 U12590 ( .A1(n10190), .A2(n10189), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17796) );
  NOR2_X1 U12591 ( .A1(n17796), .A2(n9932), .ZN(n18099) );
  NOR2_X1 U12592 ( .A1(n9927), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n9932) );
  XNOR2_X1 U12593 ( .A(n11293), .B(n11292), .ZN(n17772) );
  NOR2_X1 U12594 ( .A1(n17788), .A2(n11290), .ZN(n11293) );
  NOR2_X1 U12595 ( .A1(n9941), .A2(n9940), .ZN(n11304) );
  NAND4_X1 U12596 ( .A1(n18009), .A2(n17642), .A3(n17987), .A4(n11303), .ZN(
        n9940) );
  NOR2_X2 U12597 ( .A1(n17749), .A2(n18071), .ZN(n17748) );
  NAND4_X1 U12598 ( .A1(n17513), .A2(n10157), .A3(n17851), .A4(n10156), .ZN(
        n10163) );
  NAND2_X2 U12599 ( .A1(n9944), .A2(n9943), .ZN(n17621) );
  NAND2_X2 U12600 ( .A1(n11969), .A2(n11970), .ZN(n12455) );
  INV_X1 U12601 ( .A(n15295), .ZN(n9950) );
  INV_X1 U12602 ( .A(n12791), .ZN(n9948) );
  NAND2_X1 U12603 ( .A1(n9948), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9951) );
  INV_X1 U12604 ( .A(n14939), .ZN(n15112) );
  OR2_X2 U12605 ( .A1(n12126), .A2(n13099), .ZN(n12139) );
  AND2_X4 U12606 ( .A1(n12029), .A2(n12468), .ZN(n13966) );
  NAND3_X1 U12607 ( .A1(n12468), .A2(n9960), .A3(n9959), .ZN(n12064) );
  INV_X1 U12608 ( .A(n12045), .ZN(n9959) );
  NAND3_X1 U12609 ( .A1(n9962), .A2(n13064), .A3(n13016), .ZN(n12028) );
  AOI21_X2 U12610 ( .B1(n9966), .B2(n9964), .A(n9963), .ZN(n19230) );
  OAI21_X2 U12611 ( .B1(n15253), .B2(n10134), .A(n10133), .ZN(n15235) );
  NAND2_X2 U12612 ( .A1(n9977), .A2(n12272), .ZN(n15253) );
  NAND2_X1 U12613 ( .A1(n12365), .A2(n9878), .ZN(n9969) );
  NAND3_X1 U12614 ( .A1(n9970), .A2(n9968), .A3(n9967), .ZN(n12819) );
  OAI21_X1 U12615 ( .B1(n12365), .B2(n12371), .A(n9969), .ZN(n9968) );
  NAND3_X1 U12616 ( .A1(n9971), .A2(n12365), .A3(n9973), .ZN(n9970) );
  INV_X1 U12617 ( .A(n14917), .ZN(n9971) );
  NAND2_X2 U12618 ( .A1(n9975), .A2(n9974), .ZN(n10143) );
  OR2_X2 U12619 ( .A1(n14944), .A2(n14943), .ZN(n9975) );
  NAND2_X2 U12620 ( .A1(n12011), .A2(n12014), .ZN(n12030) );
  NAND3_X1 U12621 ( .A1(n12409), .A2(n15344), .A3(n12403), .ZN(n12454) );
  NAND2_X1 U12622 ( .A1(n12030), .A2(n19283), .ZN(n12403) );
  XNOR2_X1 U12623 ( .A(n12033), .B(n12022), .ZN(n12410) );
  NAND2_X1 U12624 ( .A1(n9980), .A2(n9979), .ZN(n14508) );
  XNOR2_X1 U12625 ( .A(n10560), .B(n20283), .ZN(n9985) );
  NAND2_X1 U12626 ( .A1(n9985), .A2(n20718), .ZN(n10578) );
  NAND2_X1 U12627 ( .A1(n13412), .A2(n13310), .ZN(n20254) );
  NOR2_X1 U12628 ( .A1(n13412), .A2(n9981), .ZN(n20492) );
  OAI21_X1 U12629 ( .B1(n13412), .B2(n14721), .A(n9983), .ZN(n9982) );
  AND2_X1 U12630 ( .A1(n20065), .A2(n9985), .ZN(n9984) );
  NAND2_X2 U12631 ( .A1(n9987), .A2(n9874), .ZN(n14636) );
  OAI21_X2 U12632 ( .B1(n14578), .B2(n9988), .A(n14587), .ZN(n15720) );
  NAND2_X2 U12633 ( .A1(n11604), .A2(n15734), .ZN(n14578) );
  AOI21_X1 U12634 ( .B1(n18856), .B2(n9996), .A(n10004), .ZN(n15497) );
  NAND2_X1 U12635 ( .A1(n14928), .A2(n9921), .ZN(n13469) );
  INV_X1 U12636 ( .A(n15486), .ZN(n10001) );
  AOI21_X1 U12637 ( .B1(n16041), .B2(n10005), .A(n10008), .ZN(n10007) );
  INV_X1 U12638 ( .A(n16041), .ZN(n10006) );
  NAND4_X1 U12639 ( .A1(n10020), .A2(n13632), .A3(n10613), .A4(n10612), .ZN(
        n13581) );
  AOI21_X1 U12640 ( .B1(n11574), .B2(n10775), .A(n10660), .ZN(n13630) );
  INV_X1 U12641 ( .A(n13743), .ZN(n10022) );
  NAND2_X1 U12642 ( .A1(n10022), .A2(n10023), .ZN(n14431) );
  NAND2_X2 U12643 ( .A1(n10547), .A2(n10546), .ZN(n10581) );
  AND2_X1 U12644 ( .A1(n14353), .A2(n10031), .ZN(n10233) );
  NAND2_X1 U12645 ( .A1(n14353), .A2(n10029), .ZN(n11783) );
  INV_X1 U12646 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10038) );
  INV_X1 U12647 ( .A(n16690), .ZN(n10039) );
  NAND2_X1 U12648 ( .A1(n10040), .A2(n10041), .ZN(n17691) );
  OAI211_X2 U12649 ( .C1(n10048), .C2(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n10047), .B(n10044), .ZN(n16798) );
  NOR2_X1 U12650 ( .A1(n14357), .A2(n10061), .ZN(n14331) );
  AND2_X1 U12651 ( .A1(n12300), .A2(n9912), .ZN(n12286) );
  AND2_X1 U12652 ( .A1(n12300), .A2(n12301), .ZN(n12299) );
  NAND2_X1 U12653 ( .A1(n12300), .A2(n9907), .ZN(n12343) );
  INV_X1 U12654 ( .A(n12247), .ZN(n10075) );
  NAND3_X1 U12655 ( .A1(n10075), .A2(n11895), .A3(n10077), .ZN(n12261) );
  NAND3_X1 U12656 ( .A1(n11895), .A2(n10075), .A3(n12229), .ZN(n12231) );
  NAND2_X1 U12657 ( .A1(n12285), .A2(n10079), .ZN(n11946) );
  NAND2_X1 U12658 ( .A1(n12285), .A2(n10081), .ZN(n12349) );
  NAND2_X1 U12659 ( .A1(n12030), .A2(n19278), .ZN(n10086) );
  NAND2_X2 U12660 ( .A1(n11958), .A2(n11957), .ZN(n12022) );
  NAND2_X2 U12661 ( .A1(n11816), .A2(n11815), .ZN(n12033) );
  NAND2_X4 U12662 ( .A1(n10085), .A2(n10084), .ZN(n19273) );
  NAND2_X1 U12663 ( .A1(n13914), .A2(n9930), .ZN(n15035) );
  NAND3_X1 U12664 ( .A1(n10090), .A2(n10089), .A3(n10088), .ZN(P2_U2997) );
  NAND3_X1 U12665 ( .A1(n12109), .A2(n13089), .A3(n12108), .ZN(n10104) );
  NAND2_X1 U12666 ( .A1(n14804), .A2(n9909), .ZN(n14791) );
  NAND2_X2 U12667 ( .A1(n10130), .A2(n11840), .ZN(n12031) );
  AOI21_X1 U12668 ( .B1(n13501), .B2(n10119), .A(n9905), .ZN(n10117) );
  NAND2_X1 U12669 ( .A1(n13501), .A2(n13502), .ZN(n13500) );
  NAND3_X1 U12670 ( .A1(n12745), .A2(n12747), .A3(n14872), .ZN(n10122) );
  NAND2_X1 U12671 ( .A1(n15274), .A2(n9904), .ZN(n16211) );
  NAND3_X1 U12672 ( .A1(n14840), .A2(n14834), .A3(n12756), .ZN(n10125) );
  INV_X1 U12673 ( .A(n14840), .ZN(n10126) );
  NAND2_X1 U12674 ( .A1(n15237), .A2(n9906), .ZN(n15222) );
  NAND2_X1 U12675 ( .A1(n12768), .A2(n13861), .ZN(n12226) );
  AND2_X2 U12676 ( .A1(n12795), .A2(n12223), .ZN(n12768) );
  INV_X1 U12677 ( .A(n12222), .ZN(n10131) );
  OAI21_X2 U12678 ( .B1(n12341), .B2(n15235), .A(n10132), .ZN(n15137) );
  NAND2_X1 U12679 ( .A1(n14960), .A2(n10135), .ZN(n10137) );
  NAND3_X1 U12680 ( .A1(n10143), .A2(n14926), .A3(n10142), .ZN(n10145) );
  INV_X1 U12681 ( .A(n15109), .ZN(n10146) );
  NAND2_X1 U12682 ( .A1(n12255), .A2(n9843), .ZN(n10150) );
  CLKBUF_X1 U12683 ( .A(n10150), .Z(n10147) );
  NAND2_X1 U12684 ( .A1(n12255), .A2(n12254), .ZN(n15051) );
  NAND2_X1 U12685 ( .A1(n11608), .A2(n10151), .ZN(n14550) );
  AND2_X2 U12686 ( .A1(n14562), .A2(n11606), .ZN(n11608) );
  NAND2_X1 U12687 ( .A1(n10152), .A2(n10153), .ZN(n10545) );
  NAND3_X1 U12688 ( .A1(n10560), .A2(n10533), .A3(n10155), .ZN(n10152) );
  NAND3_X1 U12689 ( .A1(n10157), .A2(n17513), .A3(n10156), .ZN(n17495) );
  NAND2_X1 U12690 ( .A1(n10162), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10158) );
  NAND2_X1 U12691 ( .A1(n10162), .A2(n10161), .ZN(n10160) );
  INV_X1 U12692 ( .A(n10163), .ZN(n17494) );
  NOR2_X1 U12693 ( .A1(n17702), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10165) );
  NAND2_X1 U12694 ( .A1(n10166), .A2(n11623), .ZN(n10167) );
  NAND2_X1 U12695 ( .A1(n10392), .A2(n10417), .ZN(n11640) );
  NAND3_X1 U12696 ( .A1(n11097), .A2(n10170), .A3(n11154), .ZN(n10393) );
  NAND2_X2 U12697 ( .A1(n10406), .A2(n10169), .ZN(n11154) );
  AND3_X2 U12698 ( .A1(n10340), .A2(n10341), .A3(n10231), .ZN(n10406) );
  NAND2_X1 U12699 ( .A1(n10176), .A2(n9842), .ZN(n10172) );
  NAND2_X1 U12700 ( .A1(n13376), .A2(n13377), .ZN(n10176) );
  NAND2_X1 U12701 ( .A1(n13534), .A2(n13535), .ZN(n11556) );
  NAND2_X1 U12702 ( .A1(n10173), .A2(n13376), .ZN(n10171) );
  INV_X1 U12703 ( .A(n11297), .ZN(n10179) );
  NAND3_X1 U12704 ( .A1(n10181), .A2(n10180), .A3(n17702), .ZN(n10184) );
  OAI21_X1 U12705 ( .B1(n17748), .B2(n11301), .A(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10180) );
  NAND2_X1 U12706 ( .A1(n10183), .A2(n10182), .ZN(n10181) );
  NOR2_X1 U12707 ( .A1(n11301), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10182) );
  INV_X1 U12708 ( .A(n17748), .ZN(n10183) );
  INV_X1 U12709 ( .A(n10184), .ZN(n17733) );
  OAI21_X2 U12710 ( .B1(n11604), .B2(n10187), .A(n10185), .ZN(n15721) );
  NAND3_X1 U12711 ( .A1(n10193), .A2(n10192), .A3(n11286), .ZN(n10189) );
  NAND2_X1 U12712 ( .A1(n10191), .A2(n10194), .ZN(n10190) );
  INV_X1 U12713 ( .A(n10193), .ZN(n17807) );
  NAND2_X1 U12714 ( .A1(n10193), .A2(n10192), .ZN(n10191) );
  INV_X1 U12715 ( .A(n11285), .ZN(n10192) );
  NOR2_X1 U12716 ( .A1(n17807), .A2(n11285), .ZN(n11287) );
  NAND2_X1 U12717 ( .A1(n14636), .A2(n10198), .ZN(n15735) );
  NAND3_X1 U12718 ( .A1(n11307), .A2(n17950), .A3(n11306), .ZN(n17609) );
  INV_X1 U12719 ( .A(n10200), .ZN(n17471) );
  NOR2_X1 U12720 ( .A1(n10202), .A2(n17469), .ZN(n16363) );
  NAND2_X1 U12721 ( .A1(n17483), .A2(n10201), .ZN(n10200) );
  NAND2_X1 U12722 ( .A1(n17482), .A2(n17734), .ZN(n10201) );
  NAND3_X1 U12723 ( .A1(n10581), .A2(n10550), .A3(n11627), .ZN(n11523) );
  NAND2_X1 U12724 ( .A1(n9867), .A2(n11834), .ZN(n10205) );
  NAND3_X1 U12725 ( .A1(n12044), .A2(n13053), .A3(n10206), .ZN(n12423) );
  NAND3_X1 U12726 ( .A1(n12017), .A2(n12423), .A3(n19273), .ZN(n12018) );
  NAND3_X1 U12727 ( .A1(n12167), .A2(n12169), .A3(n12166), .ZN(n10208) );
  NAND2_X1 U12728 ( .A1(n12114), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10210) );
  NAND2_X1 U12729 ( .A1(n9882), .A2(n10213), .ZN(n14979) );
  NAND2_X1 U12730 ( .A1(n10217), .A2(n15269), .ZN(n10213) );
  NAND2_X1 U12731 ( .A1(n10214), .A2(n9881), .ZN(n10216) );
  OAI21_X2 U12732 ( .B1(n15269), .B2(n10218), .A(n10217), .ZN(n13914) );
  INV_X1 U12733 ( .A(n14913), .ZN(n10219) );
  NOR2_X1 U12734 ( .A1(n14913), .A2(n10221), .ZN(n13962) );
  NAND2_X1 U12735 ( .A1(n10219), .A2(n10220), .ZN(n13963) );
  NOR2_X1 U12736 ( .A1(n14913), .A2(n15081), .ZN(n14914) );
  OR2_X1 U12737 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  NAND2_X1 U12738 ( .A1(n13033), .A2(n13032), .ZN(n13035) );
  XNOR2_X1 U12739 ( .A(n14091), .B(n14118), .ZN(n14858) );
  NAND2_X1 U12740 ( .A1(n13036), .A2(n13086), .ZN(n13088) );
  NAND2_X1 U12741 ( .A1(n13035), .A2(n13034), .ZN(n13086) );
  NAND2_X1 U12742 ( .A1(n12834), .A2(n9811), .ZN(n11515) );
  CLKBUF_X1 U12743 ( .A(n12058), .Z(n15313) );
  NAND2_X1 U12744 ( .A1(n15148), .A2(n14946), .ZN(n14949) );
  NOR3_X1 U12745 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n11193), .ZN(n11379) );
  NAND2_X1 U12746 ( .A1(n17621), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11307) );
  NAND2_X1 U12747 ( .A1(n11608), .A2(n11607), .ZN(n11609) );
  NAND2_X1 U12748 ( .A1(n17576), .A2(n17564), .ZN(n17565) );
  INV_X1 U12749 ( .A(n14979), .ZN(n12807) );
  NOR2_X1 U12750 ( .A1(n12062), .A2(n10230), .ZN(n12063) );
  NAND2_X1 U12751 ( .A1(n15556), .A2(n11317), .ZN(n11325) );
  AND2_X1 U12752 ( .A1(n14262), .A2(n11987), .ZN(n12154) );
  INV_X1 U12753 ( .A(n15344), .ZN(n13064) );
  AND2_X2 U12754 ( .A1(n12022), .A2(n15344), .ZN(n13053) );
  OR2_X2 U12755 ( .A1(n12413), .A2(n12045), .ZN(n12072) );
  AND2_X4 U12756 ( .A1(n10260), .A2(n13342), .ZN(n10680) );
  NAND2_X1 U12758 ( .A1(n10519), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10411) );
  AND2_X2 U12759 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13311) );
  NOR2_X1 U12762 ( .A1(n14745), .A2(n14250), .ZN(n14274) );
  NAND2_X1 U12763 ( .A1(n13142), .A2(n11518), .ZN(n10402) );
  NAND2_X1 U12764 ( .A1(n12044), .A2(n12016), .ZN(n12862) );
  INV_X1 U12765 ( .A(n14939), .ZN(n12808) );
  INV_X1 U12766 ( .A(n13966), .ZN(n13870) );
  NAND2_X1 U12767 ( .A1(n13029), .A2(n16252), .ZN(n12136) );
  NAND2_X1 U12768 ( .A1(n13099), .A2(n13910), .ZN(n12142) );
  NAND2_X1 U12769 ( .A1(n13099), .A2(n12112), .ZN(n12115) );
  NOR2_X1 U12770 ( .A1(n12582), .A2(n13016), .ZN(n12043) );
  NAND2_X2 U12771 ( .A1(n11543), .A2(n11542), .ZN(n11548) );
  AND2_X4 U12772 ( .A1(n10249), .A2(n10260), .ZN(n11065) );
  INV_X1 U12773 ( .A(n11272), .ZN(n15405) );
  NOR2_X1 U12774 ( .A1(n20456), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10223) );
  AND2_X1 U12775 ( .A1(n16264), .A2(n15202), .ZN(n10224) );
  AND2_X1 U12776 ( .A1(n12083), .A2(n12084), .ZN(n10225) );
  OR2_X1 U12777 ( .A1(n15984), .A2(n15985), .ZN(n10227) );
  CLKBUF_X3 U12778 ( .A(n11327), .Z(n17109) );
  NOR2_X1 U12779 ( .A1(n11193), .A2(n11192), .ZN(n11327) );
  AND2_X1 U12780 ( .A1(n12122), .A2(n12121), .ZN(n10228) );
  NAND2_X1 U12781 ( .A1(n17734), .A2(n11476), .ZN(n10229) );
  AND2_X1 U12782 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U12783 ( .A1(n10339), .A2(n10390), .ZN(n10231) );
  INV_X1 U12784 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10559) );
  NOR2_X1 U12785 ( .A1(n13666), .A2(n13542), .ZN(n10232) );
  NAND2_X1 U12786 ( .A1(n17507), .A2(n17830), .ZN(n17608) );
  INV_X1 U12787 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n13030) );
  OR2_X1 U12788 ( .A1(n17414), .A2(n18643), .ZN(n17463) );
  NAND2_X1 U12789 ( .A1(n19972), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10234) );
  INV_X1 U12790 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20148) );
  INV_X1 U12791 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11606) );
  INV_X1 U12792 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15689) );
  INV_X1 U12793 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11851) );
  INV_X1 U12794 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n13470) );
  OR2_X1 U12795 ( .A1(n18868), .A2(n15496), .ZN(n10235) );
  NAND2_X1 U12796 ( .A1(n15495), .A2(n10004), .ZN(n10236) );
  NAND2_X1 U12797 ( .A1(n13098), .A2(n13097), .ZN(n13220) );
  NAND3_X2 U12798 ( .A1(n19728), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19776), 
        .ZN(n15339) );
  INV_X1 U12799 ( .A(n13861), .ZN(n13959) );
  INV_X1 U12800 ( .A(n10370), .ZN(n10429) );
  AND2_X1 U12801 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10239) );
  INV_X1 U12802 ( .A(n10421), .ZN(n11692) );
  INV_X1 U12803 ( .A(n11692), .ZN(n11669) );
  INV_X1 U12804 ( .A(n11148), .ZN(n11130) );
  NOR2_X1 U12805 ( .A1(n11130), .A2(n11156), .ZN(n11132) );
  OR2_X1 U12806 ( .A1(n11120), .A2(n20156), .ZN(n11138) );
  INV_X1 U12807 ( .A(n10422), .ZN(n10326) );
  NAND2_X1 U12808 ( .A1(n11999), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11830) );
  NAND2_X1 U12809 ( .A1(n11871), .A2(n11870), .ZN(n11874) );
  INV_X1 U12810 ( .A(n11105), .ZN(n11118) );
  INV_X1 U12811 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10244) );
  INV_X1 U12812 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10516) );
  NAND2_X1 U12813 ( .A1(n10521), .A2(n10520), .ZN(n10527) );
  OR2_X1 U12814 ( .A1(n10513), .A2(n10512), .ZN(n10514) );
  INV_X1 U12815 ( .A(n11888), .ZN(n11892) );
  INV_X1 U12816 ( .A(n14143), .ZN(n14144) );
  AOI22_X1 U12817 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19454), .B1(
        n19529), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12143) );
  OAI21_X1 U12818 ( .B1(n11412), .B2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n11414), .ZN(n11415) );
  NAND2_X1 U12819 ( .A1(n11101), .A2(n11100), .ZN(n11104) );
  NAND2_X1 U12820 ( .A1(n10426), .A2(n10425), .ZN(n10427) );
  OR2_X1 U12821 ( .A1(n13800), .A2(n13765), .ZN(n10782) );
  OR2_X1 U12822 ( .A1(n13103), .A2(n11537), .ZN(n11538) );
  OR2_X1 U12823 ( .A1(n10623), .A2(n10622), .ZN(n11560) );
  XNOR2_X1 U12824 ( .A(n10545), .B(n10544), .ZN(n10549) );
  AOI21_X1 U12825 ( .B1(n11892), .B2(n11891), .A(n11890), .ZN(n12386) );
  NAND2_X1 U12826 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11834) );
  AND4_X1 U12827 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11935) );
  INV_X1 U12828 ( .A(n12790), .ZN(n12221) );
  NAND2_X1 U12829 ( .A1(n12584), .A2(n12612), .ZN(n12178) );
  AND2_X1 U12830 ( .A1(n14198), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n13034) );
  AOI22_X1 U12831 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U12832 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11997) );
  NOR2_X1 U12833 ( .A1(n15463), .A2(n11193), .ZN(n11234) );
  AND2_X1 U12834 ( .A1(n11434), .A2(n11435), .ZN(n11413) );
  NOR2_X1 U12835 ( .A1(n10994), .A2(n14554), .ZN(n10995) );
  INV_X1 U12836 ( .A(n14432), .ZN(n10850) );
  INV_X1 U12837 ( .A(n10388), .ZN(n10441) );
  INV_X1 U12838 ( .A(n14173), .ZN(n14169) );
  INV_X1 U12839 ( .A(n19273), .ZN(n12396) );
  OR2_X1 U12840 ( .A1(n13025), .A2(n13040), .ZN(n13041) );
  INV_X1 U12841 ( .A(n12115), .ZN(n12117) );
  NOR2_X1 U12842 ( .A1(n11296), .A2(n17760), .ZN(n11297) );
  AOI21_X1 U12843 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18623), .A(
        n11413), .ZN(n11423) );
  AND2_X1 U12844 ( .A1(n11114), .A2(n9826), .ZN(n11129) );
  AND3_X1 U12845 ( .A1(n13448), .A2(n13450), .A3(n13449), .ZN(n20046) );
  NAND2_X1 U12846 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n10344) );
  NAND2_X1 U12847 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10368) );
  NAND2_X1 U12848 ( .A1(n10995), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11021) );
  INV_X1 U12849 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10690) );
  AND2_X1 U12850 ( .A1(n14599), .A2(n14615), .ZN(n15734) );
  AND2_X1 U12851 ( .A1(n11753), .A2(n11748), .ZN(n13314) );
  NAND2_X1 U12852 ( .A1(n10564), .A2(n10563), .ZN(n20283) );
  INV_X1 U12853 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n15515) );
  INV_X1 U12854 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20531) );
  NOR2_X1 U12855 ( .A1(n19273), .A2(n19283), .ZN(n12012) );
  NAND2_X1 U12856 ( .A1(n12257), .A2(n10206), .ZN(n12350) );
  INV_X1 U12857 ( .A(n13970), .ZN(n13875) );
  OR2_X1 U12858 ( .A1(n13543), .A2(n13542), .ZN(n13663) );
  AND2_X1 U12859 ( .A1(n16064), .A2(n14118), .ZN(n14092) );
  AND2_X1 U12860 ( .A1(n12347), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12348) );
  NAND2_X1 U12861 ( .A1(n13042), .A2(n13041), .ZN(n13087) );
  AND2_X1 U12862 ( .A1(n12398), .A2(n12395), .ZN(n13001) );
  OR2_X1 U12863 ( .A1(n18594), .A2(n11495), .ZN(n13842) );
  NOR2_X1 U12864 ( .A1(n18616), .A2(n18176), .ZN(n11489) );
  INV_X1 U12865 ( .A(n15556), .ZN(n11320) );
  OAI21_X1 U12866 ( .B1(n17621), .B2(n17526), .A(n11309), .ZN(n11310) );
  NAND2_X1 U12867 ( .A1(n17565), .A2(n17884), .ZN(n17535) );
  NOR2_X1 U12868 ( .A1(n17761), .A2(n11295), .ZN(n11298) );
  XOR2_X1 U12869 ( .A(n11295), .B(n17759), .Z(n11296) );
  NAND2_X1 U12870 ( .A1(n18617), .A2(n17936), .ZN(n17982) );
  INV_X1 U12871 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14398) );
  NAND2_X1 U12872 ( .A1(n10605), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10628) );
  INV_X1 U12873 ( .A(n11717), .ZN(n11742) );
  INV_X1 U12874 ( .A(n10627), .ZN(n10775) );
  OAI211_X1 U12875 ( .C1(n9913), .C2(n10651), .A(n10650), .B(n10649), .ZN(
        n13632) );
  OR2_X1 U12876 ( .A1(n13155), .A2(n11782), .ZN(n15530) );
  OR3_X1 U12877 ( .A1(n15795), .A2(n15796), .A3(n14516), .ZN(n14664) );
  NAND2_X1 U12878 ( .A1(n15864), .A2(n11772), .ZN(n15804) );
  AND2_X1 U12879 ( .A1(n11680), .A2(n11679), .ZN(n15697) );
  OAI21_X1 U12880 ( .B1(n20804), .B2(n15949), .A(n20786), .ZN(n13595) );
  OR2_X1 U12881 ( .A1(n20368), .A2(n20569), .ZN(n20336) );
  INV_X1 U12882 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20489) );
  OR2_X1 U12883 ( .A1(n13589), .A2(n13407), .ZN(n20500) );
  OR2_X1 U12884 ( .A1(n20649), .A2(n20526), .ZN(n20561) );
  OR2_X1 U12885 ( .A1(n13155), .A2(n15563), .ZN(n15543) );
  AOI21_X1 U12886 ( .B1(n15979), .B2(n19069), .A(n15978), .ZN(n15980) );
  INV_X1 U12887 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18972) );
  NAND2_X1 U12888 ( .A1(n9917), .A2(n14798), .ZN(n14797) );
  AND2_X1 U12889 ( .A1(n15205), .A2(n16187), .ZN(n15206) );
  OR3_X1 U12890 ( .A1(n18941), .A2(n13861), .A3(n12512), .ZN(n13911) );
  NAND2_X1 U12891 ( .A1(n12810), .A2(n12453), .ZN(n15202) );
  INV_X1 U12892 ( .A(n16257), .ZN(n15285) );
  AND3_X1 U12893 ( .A1(n13004), .A2(n13003), .A3(n13002), .ZN(n16293) );
  OR3_X1 U12894 ( .A1(n19310), .A2(n19500), .A3(n19305), .ZN(n19350) );
  OR2_X1 U12895 ( .A1(n19940), .A2(n19943), .ZN(n19560) );
  NOR2_X2 U12896 ( .A1(n13842), .A2(n18820), .ZN(n18613) );
  NOR2_X1 U12897 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16682), .ZN(n16667) );
  NOR2_X1 U12898 ( .A1(n18582), .A2(n13842), .ZN(n15441) );
  AOI211_X1 U12899 ( .C1(n17131), .C2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n11278), .B(n11277), .ZN(n11281) );
  NAND2_X1 U12900 ( .A1(n12840), .A2(n17818), .ZN(n12841) );
  NOR2_X1 U12901 ( .A1(n17526), .A2(n17970), .ZN(n17527) );
  NOR2_X1 U12902 ( .A1(n17681), .A2(n17670), .ZN(n17664) );
  INV_X1 U12903 ( .A(n11510), .ZN(n11511) );
  INV_X1 U12904 ( .A(n18615), .ZN(n18605) );
  NOR2_X1 U12905 ( .A1(n17325), .A2(n11453), .ZN(n17758) );
  AOI211_X1 U12906 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n11375), .B(n11374), .ZN(n11376) );
  NAND2_X1 U12907 ( .A1(n18808), .A2(n18053), .ZN(n18017) );
  AND2_X1 U12908 ( .A1(n11153), .A2(n11152), .ZN(n13155) );
  OR2_X1 U12909 ( .A1(n15548), .A2(n20718), .ZN(n13128) );
  NAND2_X1 U12910 ( .A1(n10830), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10852) );
  AND2_X1 U12911 ( .A1(n15629), .A2(n13438), .ZN(n20025) );
  INV_X1 U12912 ( .A(n15630), .ZN(n15644) );
  INV_X1 U12913 ( .A(n15688), .ZN(n20061) );
  INV_X1 U12914 ( .A(n14439), .ZN(n20074) );
  INV_X1 U12915 ( .A(n15712), .ZN(n20073) );
  AND2_X1 U12916 ( .A1(n10885), .A2(n10884), .ZN(n14424) );
  INV_X1 U12917 ( .A(n14502), .ZN(n14487) );
  OR2_X1 U12918 ( .A1(n13130), .A2(n12958), .ZN(n11166) );
  INV_X1 U12919 ( .A(n13256), .ZN(n13251) );
  AOI21_X1 U12920 ( .B1(n15783), .B2(n14307), .A(n11790), .ZN(n11791) );
  NAND2_X1 U12921 ( .A1(n10888), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10949) );
  AOI21_X1 U12922 ( .B1(n9925), .B2(n9833), .A(n14492), .ZN(n15708) );
  NAND2_X1 U12923 ( .A1(n10739), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10763) );
  AND2_X1 U12924 ( .A1(n10656), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10675) );
  AND2_X1 U12925 ( .A1(n15790), .A2(n20124), .ZN(n15783) );
  NOR2_X1 U12926 ( .A1(n15804), .A2(n15570), .ZN(n15808) );
  OR2_X1 U12927 ( .A1(n13229), .A2(n15816), .ZN(n15827) );
  AND2_X1 U12928 ( .A1(n15927), .A2(n11771), .ZN(n15864) );
  INV_X1 U12929 ( .A(n15822), .ZN(n15821) );
  AND2_X1 U12930 ( .A1(n11787), .A2(n20721), .ZN(n15935) );
  AND2_X1 U12931 ( .A1(n11761), .A2(n15506), .ZN(n15816) );
  NAND2_X1 U12932 ( .A1(n20718), .A2(n13595), .ZN(n20289) );
  NOR2_X1 U12933 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15942) );
  AND2_X1 U12934 ( .A1(n20250), .A2(n20400), .ZN(n20216) );
  OAI21_X1 U12935 ( .B1(n20225), .B2(n20224), .A(n20223), .ZN(n20246) );
  NOR2_X2 U12936 ( .A1(n20262), .A2(n20596), .ZN(n20278) );
  OR2_X1 U12937 ( .A1(n20220), .A2(n13590), .ZN(n20526) );
  INV_X1 U12938 ( .A(n20336), .ZN(n20363) );
  INV_X1 U12939 ( .A(n20393), .ZN(n20389) );
  INV_X1 U12940 ( .A(n20404), .ZN(n20425) );
  INV_X1 U12941 ( .A(n20526), .ZN(n20400) );
  INV_X1 U12942 ( .A(n20524), .ZN(n20479) );
  AND2_X1 U12943 ( .A1(n20220), .A2(n11527), .ZN(n20453) );
  NOR2_X2 U12944 ( .A1(n20500), .A2(n20499), .ZN(n20564) );
  INV_X1 U12945 ( .A(n20289), .ZN(n20196) );
  OR2_X1 U12946 ( .A1(n20220), .A2(n11527), .ZN(n20569) );
  INV_X1 U12947 ( .A(n20706), .ZN(n20635) );
  INV_X1 U12948 ( .A(n20546), .ZN(n20670) );
  INV_X1 U12949 ( .A(n20715), .ZN(n20692) );
  NAND2_X1 U12950 ( .A1(n20220), .A2(n13590), .ZN(n20499) );
  INV_X1 U12951 ( .A(n15980), .ZN(n15981) );
  OR2_X1 U12952 ( .A1(n12736), .A2(n12735), .ZN(n13545) );
  OR2_X1 U12953 ( .A1(n12655), .A2(n12654), .ZN(n13355) );
  INV_X1 U12954 ( .A(n19952), .ZN(n19527) );
  INV_X1 U12955 ( .A(n12910), .ZN(n12930) );
  AND2_X1 U12956 ( .A1(n13480), .A2(n12584), .ZN(n13486) );
  INV_X1 U12957 ( .A(n16173), .ZN(n19240) );
  OR2_X1 U12958 ( .A1(n14917), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15073) );
  NOR2_X1 U12959 ( .A1(n16189), .A2(n15206), .ZN(n15207) );
  INV_X1 U12960 ( .A(n16264), .ZN(n19262) );
  XNOR2_X1 U12961 ( .A(n13088), .B(n13043), .ZN(n19940) );
  OAI21_X1 U12962 ( .B1(n15329), .B2(n15330), .A(n15327), .ZN(n19296) );
  NOR2_X2 U12963 ( .A1(n19560), .A2(n19422), .ZN(n19352) );
  NOR2_X1 U12964 ( .A1(n19560), .A2(n19499), .ZN(n19370) );
  OR2_X1 U12965 ( .A1(n19940), .A2(n19361), .ZN(n19630) );
  NAND2_X1 U12966 ( .A1(n19940), .A2(n19361), .ZN(n19684) );
  OR2_X1 U12967 ( .A1(n15356), .A2(n15355), .ZN(n19495) );
  NAND2_X1 U12968 ( .A1(n19940), .A2(n19943), .ZN(n19926) );
  NOR2_X1 U12969 ( .A1(n19725), .A2(n19560), .ZN(n19575) );
  NOR2_X1 U12970 ( .A1(n19683), .A2(n19630), .ZN(n19656) );
  INV_X1 U12971 ( .A(n19827), .ZN(n19753) );
  AND2_X1 U12972 ( .A1(n19283), .A2(n19291), .ZN(n19800) );
  AND2_X1 U12973 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n12448), .ZN(n19829) );
  XNOR2_X1 U12974 ( .A(n18808), .B(n15442), .ZN(n18810) );
  INV_X1 U12975 ( .A(n16872), .ZN(n16863) );
  NOR2_X1 U12976 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16637), .ZN(n16621) );
  NOR2_X1 U12977 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16654), .ZN(n16643) );
  NOR2_X1 U12978 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16711), .ZN(n16693) );
  NOR2_X1 U12979 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16732), .ZN(n16715) );
  NOR2_X1 U12980 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16784), .ZN(n16763) );
  INV_X1 U12981 ( .A(n16857), .ZN(n16851) );
  NOR2_X1 U12982 ( .A1(n16988), .A2(n17003), .ZN(n16972) );
  OAI21_X1 U12983 ( .B1(n15441), .B2(n15440), .A(n18642), .ZN(n15581) );
  NOR2_X1 U12984 ( .A1(n17357), .A2(n17227), .ZN(n17221) );
  NAND2_X1 U12985 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17237), .ZN(n17236) );
  NOR2_X1 U12986 ( .A1(n17373), .A2(n17266), .ZN(n17261) );
  NOR2_X1 U12987 ( .A1(n17464), .A2(n17288), .ZN(n17282) );
  NOR2_X1 U12988 ( .A1(n17700), .A2(n16353), .ZN(n17616) );
  NAND2_X1 U12989 ( .A1(n9943), .A2(n18018), .ZN(n17970) );
  NAND2_X1 U12990 ( .A1(n11475), .A2(n17735), .ZN(n18018) );
  INV_X1 U12991 ( .A(n18498), .ZN(n18529) );
  NOR2_X2 U12992 ( .A1(n18813), .A2(n17707), .ZN(n17685) );
  INV_X1 U12993 ( .A(n16343), .ZN(n16367) );
  INV_X1 U12994 ( .A(n18036), .ZN(n18042) );
  NOR2_X1 U12995 ( .A1(n17874), .A2(n17524), .ZN(n17512) );
  INV_X1 U12996 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18009) );
  INV_X1 U12997 ( .A(n18127), .ZN(n18137) );
  NOR2_X1 U12998 ( .A1(n18588), .A2(n18127), .ZN(n18136) );
  INV_X1 U12999 ( .A(n18446), .ZN(n18517) );
  INV_X1 U13000 ( .A(n16989), .ZN(n18188) );
  OR2_X1 U13001 ( .A1(n13155), .A2(n12943), .ZN(n13172) );
  INV_X1 U13002 ( .A(n20024), .ZN(n20064) );
  INV_X1 U13003 ( .A(n20025), .ZN(n15623) );
  INV_X1 U13004 ( .A(n20041), .ZN(n20071) );
  NAND2_X1 U13005 ( .A1(n20078), .A2(n13133), .ZN(n15712) );
  INV_X1 U13006 ( .A(n20082), .ZN(n20108) );
  NOR2_X1 U13007 ( .A1(n13172), .A2(n13171), .ZN(n13255) );
  INV_X1 U13008 ( .A(n15783), .ZN(n15782) );
  INV_X1 U13009 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20033) );
  INV_X1 U13010 ( .A(n15932), .ZN(n20137) );
  INV_X1 U13011 ( .A(n15935), .ZN(n20135) );
  NOR2_X1 U13012 ( .A1(n15825), .A2(n15888), .ZN(n15906) );
  INV_X1 U13013 ( .A(n15933), .ZN(n20138) );
  INV_X1 U13014 ( .A(n13603), .ZN(n20191) );
  NAND2_X1 U13015 ( .A1(n20250), .A2(n20192), .ZN(n20244) );
  AOI22_X1 U13016 ( .A1(n20222), .A2(n20224), .B1(n20458), .B2(n10223), .ZN(
        n20249) );
  AOI22_X1 U13017 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20256), .B1(n20255), 
        .B2(n20260), .ZN(n20282) );
  OR2_X1 U13018 ( .A1(n20368), .A2(n20526), .ZN(n20335) );
  AOI22_X1 U13019 ( .A1(n20342), .A2(n20339), .B1(n10223), .B2(n20530), .ZN(
        n20367) );
  OR2_X1 U13020 ( .A1(n20368), .A2(n20499), .ZN(n20404) );
  NAND2_X1 U13021 ( .A1(n20494), .A2(n20400), .ZN(n20452) );
  AOI22_X1 U13022 ( .A1(n20463), .A2(n20459), .B1(n20458), .B2(n20457), .ZN(
        n20488) );
  NAND2_X1 U13023 ( .A1(n20494), .A2(n20453), .ZN(n20524) );
  AOI22_X1 U13024 ( .A1(n20535), .A2(n20532), .B1(n20530), .B2(n20529), .ZN(
        n20568) );
  OR2_X1 U13025 ( .A1(n20649), .A2(n20569), .ZN(n20602) );
  OR2_X1 U13026 ( .A1(n20649), .A2(n20596), .ZN(n20695) );
  INV_X1 U13027 ( .A(n20784), .ZN(n20780) );
  INV_X1 U13028 ( .A(n20758), .ZN(n20771) );
  NAND2_X1 U13029 ( .A1(n12818), .A2(n19829), .ZN(n12869) );
  INV_X1 U13030 ( .A(n19069), .ZN(n19055) );
  AND2_X1 U13031 ( .A1(n13052), .A2(n19829), .ZN(n19162) );
  NAND2_X1 U13032 ( .A1(n13062), .A2(n19162), .ZN(n19191) );
  INV_X1 U13033 ( .A(n19197), .ZN(n19229) );
  INV_X1 U13034 ( .A(n13486), .ZN(n12975) );
  INV_X1 U13035 ( .A(n19242), .ZN(n16172) );
  INV_X1 U13036 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18955) );
  INV_X1 U13037 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16178) );
  INV_X1 U13038 ( .A(n19263), .ZN(n16246) );
  NAND2_X1 U13039 ( .A1(n12810), .A2(n19964), .ZN(n16264) );
  AND2_X1 U13040 ( .A1(n15337), .A2(n15336), .ZN(n19300) );
  INV_X1 U13041 ( .A(n19370), .ZN(n19386) );
  OR2_X1 U13042 ( .A1(n19422), .A2(n19630), .ZN(n19416) );
  OR2_X1 U13043 ( .A1(n19499), .A2(n19630), .ZN(n19443) );
  OR2_X1 U13044 ( .A1(n19422), .A2(n19684), .ZN(n19464) );
  INV_X1 U13045 ( .A(n19490), .ZN(n19498) );
  OR2_X1 U13046 ( .A1(n19499), .A2(n19926), .ZN(n19557) );
  INV_X1 U13047 ( .A(n19575), .ZN(n19588) );
  INV_X1 U13048 ( .A(n19602), .ZN(n19618) );
  INV_X1 U13049 ( .A(n19656), .ZN(n19682) );
  NAND2_X1 U13050 ( .A1(n19685), .A2(n19689), .ZN(n19756) );
  NAND2_X1 U13051 ( .A1(n19726), .A2(n19771), .ZN(n19827) );
  INV_X1 U13052 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19979) );
  INV_X1 U13053 ( .A(n19911), .ZN(n19837) );
  INV_X1 U13054 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18652) );
  NAND2_X1 U13055 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n16877), .ZN(n16857) );
  INV_X1 U13056 ( .A(n16873), .ZN(n16860) );
  NOR2_X1 U13057 ( .A1(n16882), .A2(n16930), .ZN(n16935) );
  NOR2_X1 U13058 ( .A1(n16733), .A2(n17103), .ZN(n17105) );
  AND2_X1 U13059 ( .A1(n17200), .A2(n18188), .ZN(n17197) );
  INV_X2 U13060 ( .A(n17197), .ZN(n17191) );
  INV_X1 U13061 ( .A(n16354), .ZN(n17319) );
  NOR2_X1 U13062 ( .A1(n11219), .A2(n11218), .ZN(n17332) );
  NOR2_X1 U13063 ( .A1(n18805), .A2(n17381), .ZN(n17377) );
  INV_X1 U13064 ( .A(n17381), .ZN(n17411) );
  INV_X1 U13065 ( .A(n17461), .ZN(n17451) );
  INV_X1 U13066 ( .A(n17685), .ZN(n17669) );
  INV_X1 U13067 ( .A(n17616), .ZN(n17633) );
  AOI22_X1 U13068 ( .A1(n17528), .A2(n17997), .B1(n17818), .B2(n18018), .ZN(
        n17700) );
  NOR2_X1 U13069 ( .A1(n17685), .A2(n17539), .ZN(n17813) );
  INV_X1 U13070 ( .A(n9811), .ZN(n18039) );
  INV_X1 U13071 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18623) );
  INV_X1 U13072 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18677) );
  NAND2_X1 U13073 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18677), .ZN(n18799) );
  NAND2_X1 U13074 ( .A1(n11185), .A2(n11184), .ZN(P1_U2873) );
  OAI21_X1 U13075 ( .B1(n14659), .B2(n19996), .A(n11792), .ZN(P1_U2970) );
  INV_X1 U13076 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10241) );
  AND2_X2 U13077 ( .A1(n10241), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10249) );
  NAND2_X1 U13078 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10248) );
  NAND2_X1 U13079 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10247) );
  INV_X1 U13080 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10243) );
  AND2_X2 U13081 ( .A1(n10243), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10259) );
  AND2_X2 U13082 ( .A1(n10249), .A2(n10259), .ZN(n10448) );
  NAND2_X1 U13083 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10246) );
  AND2_X2 U13084 ( .A1(n10244), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10254) );
  AND2_X2 U13085 ( .A1(n10254), .A2(n13330), .ZN(n10375) );
  NAND2_X1 U13086 ( .A1(n10375), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10245) );
  AND2_X2 U13087 ( .A1(n10249), .A2(n10261), .ZN(n10443) );
  NAND2_X1 U13088 ( .A1(n10443), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10253) );
  AND2_X2 U13089 ( .A1(n10254), .A2(n10259), .ZN(n11066) );
  NAND2_X1 U13090 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10252) );
  NAND2_X1 U13091 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10251) );
  AND2_X2 U13092 ( .A1(n10260), .A2(n13311), .ZN(n10370) );
  NAND2_X1 U13093 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10250) );
  AND2_X2 U13094 ( .A1(n10254), .A2(n10261), .ZN(n11007) );
  NAND2_X1 U13095 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10258) );
  NOR2_X4 U13096 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13342) );
  AND2_X2 U13097 ( .A1(n10259), .A2(n13342), .ZN(n10434) );
  NAND2_X1 U13098 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10257) );
  NAND2_X1 U13099 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n10256) );
  NAND2_X1 U13100 ( .A1(n10328), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10255) );
  AND2_X2 U13101 ( .A1(n10259), .A2(n13311), .ZN(n10318) );
  NAND2_X1 U13102 ( .A1(n10318), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10265) );
  NAND2_X1 U13103 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10264) );
  AND2_X2 U13104 ( .A1(n10261), .A2(n13342), .ZN(n10317) );
  NAND2_X1 U13105 ( .A1(n10317), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10263) );
  NAND2_X1 U13106 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10262) );
  NAND4_X4 U13107 ( .A1(n10269), .A2(n10268), .A3(n10267), .A4(n10266), .ZN(
        n10391) );
  AOI22_X1 U13108 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9832), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13109 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10443), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10272) );
  AOI22_X1 U13110 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13111 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10315), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10270) );
  NAND4_X1 U13112 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10279) );
  AOI22_X1 U13113 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10375), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13114 ( .A1(n10318), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10276) );
  AOI22_X1 U13115 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9828), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10275) );
  AOI22_X1 U13116 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10317), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10274) );
  NAND4_X1 U13117 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n10278) );
  NAND2_X1 U13118 ( .A1(n10391), .A2(n10325), .ZN(n10310) );
  NAND2_X1 U13119 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10282) );
  NAND2_X1 U13120 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n10281) );
  NAND2_X1 U13121 ( .A1(n10443), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10280) );
  NAND3_X1 U13122 ( .A1(n10282), .A2(n10281), .A3(n10280), .ZN(n10283) );
  NOR2_X1 U13123 ( .A1(n10283), .A2(n10239), .ZN(n10289) );
  NAND2_X1 U13124 ( .A1(n10318), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U13125 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10286) );
  NAND2_X1 U13126 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10285) );
  NAND2_X1 U13127 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n10284) );
  NAND2_X1 U13128 ( .A1(n10289), .A2(n10288), .ZN(n10301) );
  NAND2_X1 U13129 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10293) );
  NAND2_X1 U13130 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10292) );
  NAND2_X1 U13131 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n10291) );
  NAND2_X1 U13132 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U13133 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10297) );
  NAND2_X1 U13134 ( .A1(n10375), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10296) );
  NAND2_X1 U13135 ( .A1(n10328), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10295) );
  NAND2_X1 U13136 ( .A1(n10317), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n10294) );
  NOR2_X2 U13137 ( .A1(n10301), .A2(n10300), .ZN(n10388) );
  INV_X1 U13138 ( .A(n10342), .ZN(n11638) );
  AOI22_X1 U13139 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10305) );
  AOI22_X1 U13140 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10375), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10304) );
  AOI22_X1 U13141 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U13142 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10315), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10302) );
  AOI22_X1 U13143 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10343), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U13144 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10307) );
  AOI22_X1 U13145 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10443), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10306) );
  CLKBUF_X3 U13146 ( .A(n10317), .Z(n11069) );
  AOI22_X1 U13147 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10309) );
  NAND3_X2 U13148 ( .A1(n9863), .A2(n9840), .A3(n10309), .ZN(n10394) );
  AOI22_X1 U13149 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11075), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10314) );
  AOI22_X1 U13150 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10313) );
  AOI22_X1 U13151 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10370), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13152 ( .A1(n10443), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10343), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10311) );
  NAND4_X1 U13153 ( .A1(n10314), .A2(n10313), .A3(n10312), .A4(n10311), .ZN(
        n10324) );
  AND2_X1 U13154 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10316) );
  AOI22_X1 U13155 ( .A1(n10375), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10317), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10321) );
  AOI22_X1 U13156 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10320) );
  AOI22_X1 U13157 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10319) );
  NAND4_X1 U13158 ( .A1(n10322), .A2(n10321), .A3(n10320), .A4(n10319), .ZN(
        n10323) );
  INV_X1 U13159 ( .A(n10339), .ZN(n10327) );
  NAND2_X1 U13160 ( .A1(n10416), .A2(n10391), .ZN(n10422) );
  NAND2_X1 U13161 ( .A1(n10327), .A2(n10326), .ZN(n10400) );
  AOI22_X1 U13162 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10370), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10331) );
  AOI22_X1 U13163 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10443), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13164 ( .A1(n10317), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13165 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n10338) );
  AOI22_X1 U13166 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11075), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13167 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10375), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U13168 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10343), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13169 ( .A1(n10318), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10315), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U13170 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10337) );
  NAND2_X1 U13171 ( .A1(n10400), .A2(n11518), .ZN(n10340) );
  NAND2_X1 U13172 ( .A1(n10325), .A2(n13608), .ZN(n10390) );
  NAND2_X1 U13173 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n10347) );
  NAND2_X1 U13174 ( .A1(n11075), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10346) );
  NAND2_X1 U13175 ( .A1(n10443), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10345) );
  NAND2_X1 U13176 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10351) );
  NAND2_X1 U13177 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10350) );
  NAND2_X1 U13178 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10349) );
  NAND2_X1 U13179 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10348) );
  NAND2_X1 U13180 ( .A1(n10318), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n10355) );
  NAND2_X1 U13181 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10354) );
  NAND2_X1 U13182 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10353) );
  NAND2_X1 U13183 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10352) );
  NAND2_X1 U13184 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10359) );
  NAND2_X1 U13185 ( .A1(n10375), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10358) );
  NAND2_X1 U13186 ( .A1(n10328), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10357) );
  NAND2_X1 U13187 ( .A1(n10317), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10356) );
  NOR2_X1 U13188 ( .A1(n11745), .A2(n9827), .ZN(n10364) );
  NAND2_X1 U13189 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10367) );
  NAND2_X1 U13190 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10366) );
  NAND2_X1 U13191 ( .A1(n10343), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10365) );
  NAND2_X1 U13192 ( .A1(n10443), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10374) );
  NAND2_X1 U13193 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10373) );
  NAND2_X1 U13194 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10372) );
  NAND2_X1 U13195 ( .A1(n10370), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10371) );
  NAND2_X1 U13196 ( .A1(n10375), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10379) );
  NAND2_X1 U13197 ( .A1(n10434), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10378) );
  NAND2_X1 U13198 ( .A1(n10318), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n10377) );
  NAND2_X1 U13199 ( .A1(n10317), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10376) );
  NAND2_X1 U13200 ( .A1(n10448), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10383) );
  NAND2_X1 U13201 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13202 ( .A1(n10328), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10381) );
  NAND2_X1 U13203 ( .A1(n10315), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10380) );
  NAND4_X4 U13204 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n13447) );
  INV_X2 U13205 ( .A(n10394), .ZN(n13142) );
  INV_X2 U13206 ( .A(n10391), .ZN(n11114) );
  INV_X1 U13207 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20728) );
  XNOR2_X1 U13208 ( .A(n20728), .B(P1_STATE_REG_2__SCAN_IN), .ZN(n11623) );
  NOR3_X1 U13209 ( .A1(n10390), .A2(n11531), .A3(n13447), .ZN(n10392) );
  NOR2_X2 U13210 ( .A1(n11518), .A2(n10394), .ZN(n13328) );
  NAND2_X1 U13211 ( .A1(n10393), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10486) );
  INV_X1 U13212 ( .A(n13442), .ZN(n11107) );
  NAND2_X1 U13213 ( .A1(n10394), .A2(n13443), .ZN(n11752) );
  AND2_X1 U13214 ( .A1(n11107), .A2(n11752), .ZN(n10397) );
  NOR2_X1 U13215 ( .A1(n11745), .A2(n10421), .ZN(n13135) );
  INV_X1 U13216 ( .A(n13135), .ZN(n10396) );
  INV_X1 U13217 ( .A(n13443), .ZN(n11519) );
  NAND2_X1 U13218 ( .A1(n11114), .A2(n10325), .ZN(n10398) );
  AND2_X1 U13219 ( .A1(n10398), .A2(n13608), .ZN(n10413) );
  OR2_X2 U13220 ( .A1(n11745), .A2(n10325), .ZN(n10399) );
  AND2_X2 U13221 ( .A1(n10413), .A2(n10399), .ZN(n11749) );
  NAND2_X1 U13222 ( .A1(n11749), .A2(n11641), .ZN(n10412) );
  BUF_X1 U13223 ( .A(n10400), .Z(n10401) );
  NAND2_X1 U13224 ( .A1(n10412), .A2(n10401), .ZN(n10404) );
  INV_X1 U13225 ( .A(n10417), .ZN(n11750) );
  INV_X1 U13226 ( .A(n11518), .ZN(n20167) );
  NAND2_X1 U13227 ( .A1(n20167), .A2(n13443), .ZN(n11659) );
  NAND2_X1 U13228 ( .A1(n13106), .A2(n10403), .ZN(n11747) );
  NAND4_X1 U13229 ( .A1(n10419), .A2(n10404), .A3(n11750), .A4(n11747), .ZN(
        n10405) );
  NAND2_X1 U13230 ( .A1(n10405), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10408) );
  INV_X1 U13231 ( .A(n10406), .ZN(n10424) );
  NAND2_X1 U13232 ( .A1(n20717), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15548) );
  INV_X1 U13233 ( .A(n15548), .ZN(n10409) );
  INV_X1 U13234 ( .A(n11787), .ZN(n10482) );
  MUX2_X1 U13235 ( .A(n10409), .B(n10482), .S(n20570), .Z(n10410) );
  NAND3_X1 U13236 ( .A1(n10412), .A2(n13447), .A3(n10401), .ZN(n10420) );
  INV_X1 U13237 ( .A(n10413), .ZN(n10415) );
  NAND2_X1 U13238 ( .A1(n15942), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10414) );
  AOI21_X1 U13239 ( .B1(n10415), .B2(n15538), .A(n10414), .ZN(n10418) );
  NAND2_X1 U13240 ( .A1(n10417), .A2(n10416), .ZN(n11758) );
  NAND4_X1 U13241 ( .A1(n10420), .A2(n10419), .A3(n10418), .A4(n11758), .ZN(
        n10428) );
  AOI21_X1 U13242 ( .B1(n10422), .B2(n11518), .A(n11692), .ZN(n10423) );
  NOR2_X1 U13243 ( .A1(n13447), .A2(n13443), .ZN(n13439) );
  NAND2_X1 U13244 ( .A1(n10423), .A2(n12958), .ZN(n10426) );
  NAND2_X1 U13245 ( .A1(n10502), .A2(n20718), .ZN(n10456) );
  AOI22_X1 U13246 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10433) );
  AOI22_X1 U13247 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13248 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10370), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U13249 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10430) );
  NAND4_X1 U13250 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10440) );
  AOI22_X1 U13251 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U13252 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13253 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10436) );
  AOI22_X1 U13254 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10435) );
  NAND4_X1 U13255 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10439) );
  INV_X1 U13256 ( .A(n11588), .ZN(n10442) );
  NOR2_X1 U13257 ( .A1(n10442), .A2(n10566), .ZN(n10462) );
  NOR2_X1 U13258 ( .A1(n10566), .A2(n11588), .ZN(n10463) );
  AOI22_X1 U13259 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10447) );
  AOI22_X1 U13260 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10446) );
  AOI22_X1 U13261 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10445) );
  AOI22_X1 U13262 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10444) );
  NAND4_X1 U13263 ( .A1(n10447), .A2(n10446), .A3(n10445), .A4(n10444), .ZN(
        n10454) );
  AOI22_X1 U13264 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10452) );
  AOI22_X1 U13265 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10370), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10451) );
  AOI22_X1 U13266 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10450) );
  AOI22_X1 U13267 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10449) );
  NAND4_X1 U13268 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10453) );
  MUX2_X1 U13269 ( .A(n10462), .B(n10463), .S(n11528), .Z(n10455) );
  INV_X1 U13270 ( .A(n11528), .ZN(n10458) );
  NAND2_X1 U13271 ( .A1(n13596), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10457) );
  MUX2_X1 U13272 ( .A(n10458), .B(n10457), .S(n9827), .Z(n10460) );
  AOI21_X1 U13273 ( .B1(n11641), .B2(n11588), .A(n20718), .ZN(n10459) );
  NAND2_X1 U13274 ( .A1(n10460), .A2(n10459), .ZN(n10496) );
  INV_X1 U13275 ( .A(n10462), .ZN(n11586) );
  INV_X1 U13276 ( .A(n10463), .ZN(n10478) );
  INV_X1 U13277 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10464) );
  OR2_X1 U13278 ( .A1(n11143), .A2(n10464), .ZN(n10477) );
  AOI22_X1 U13279 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10468) );
  AOI22_X1 U13280 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10467) );
  AOI22_X1 U13281 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10466) );
  AOI22_X1 U13282 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10465) );
  NAND4_X1 U13283 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10474) );
  AOI22_X1 U13284 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10472) );
  AOI22_X1 U13285 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10471) );
  AOI22_X1 U13286 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13287 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10469) );
  NAND4_X1 U13288 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n10473) );
  NAND2_X1 U13289 ( .A1(n10475), .A2(n11529), .ZN(n10476) );
  XNOR2_X2 U13290 ( .A(n10513), .B(n10511), .ZN(n10510) );
  INV_X1 U13291 ( .A(n10479), .ZN(n10480) );
  NAND2_X1 U13292 ( .A1(n10481), .A2(n10480), .ZN(n10489) );
  INV_X1 U13293 ( .A(n10489), .ZN(n10488) );
  NAND2_X1 U13294 ( .A1(n10519), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10485) );
  NAND2_X1 U13295 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n10523) );
  OAI21_X1 U13296 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n10523), .ZN(n20456) );
  NAND2_X1 U13297 ( .A1(n15548), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10517) );
  OAI21_X1 U13298 ( .B1(n10482), .B2(n20456), .A(n10517), .ZN(n10483) );
  INV_X1 U13299 ( .A(n10483), .ZN(n10484) );
  NAND2_X1 U13300 ( .A1(n10485), .A2(n10484), .ZN(n10487) );
  NAND2_X1 U13301 ( .A1(n10488), .A2(n20252), .ZN(n10532) );
  INV_X1 U13302 ( .A(n20252), .ZN(n10490) );
  NAND2_X1 U13303 ( .A1(n10532), .A2(n20193), .ZN(n13513) );
  INV_X1 U13304 ( .A(n10566), .ZN(n11115) );
  NAND2_X1 U13305 ( .A1(n11115), .A2(n11529), .ZN(n10491) );
  INV_X1 U13306 ( .A(n11535), .ZN(n10509) );
  XNOR2_X2 U13307 ( .A(n10510), .B(n10509), .ZN(n20220) );
  NAND2_X1 U13308 ( .A1(n10416), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10627) );
  NAND2_X1 U13309 ( .A1(n20220), .A2(n10775), .ZN(n10495) );
  INV_X2 U13310 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20721) );
  INV_X2 U13311 ( .A(n9913), .ZN(n11095) );
  AOI22_X1 U13312 ( .A1(n11095), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20721), .ZN(n10493) );
  INV_X1 U13313 ( .A(n10390), .ZN(n13282) );
  NAND2_X1 U13314 ( .A1(n13282), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n10589) );
  INV_X1 U13315 ( .A(n10589), .ZN(n10606) );
  NAND2_X1 U13316 ( .A1(n10606), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10492) );
  AND2_X1 U13317 ( .A1(n10493), .A2(n10492), .ZN(n10494) );
  NAND2_X1 U13318 ( .A1(n10495), .A2(n10494), .ZN(n13215) );
  INV_X1 U13319 ( .A(n10496), .ZN(n10498) );
  NAND2_X1 U13320 ( .A1(n10498), .A2(n10497), .ZN(n10499) );
  NAND2_X1 U13321 ( .A1(n11527), .A2(n10416), .ZN(n10501) );
  NAND2_X1 U13322 ( .A1(n10501), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13125) );
  AOI22_X1 U13323 ( .A1(n11095), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20721), .ZN(n10505) );
  NAND2_X1 U13324 ( .A1(n10606), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13325 ( .A1(n10505), .A2(n10504), .ZN(n10506) );
  AOI21_X1 U13326 ( .B1(n10503), .B2(n10775), .A(n10506), .ZN(n13124) );
  OR2_X1 U13327 ( .A1(n13125), .A2(n13124), .ZN(n13127) );
  INV_X1 U13328 ( .A(n13124), .ZN(n10507) );
  OR2_X1 U13329 ( .A1(n10507), .A2(n11093), .ZN(n10508) );
  NAND2_X1 U13330 ( .A1(n13127), .A2(n10508), .ZN(n13214) );
  NAND2_X1 U13331 ( .A1(n13215), .A2(n13214), .ZN(n13267) );
  NAND2_X1 U13332 ( .A1(n10510), .A2(n10509), .ZN(n10515) );
  INV_X1 U13333 ( .A(n10511), .ZN(n10512) );
  INV_X1 U13334 ( .A(n10548), .ZN(n10547) );
  AND2_X1 U13335 ( .A1(n10517), .A2(n10516), .ZN(n10518) );
  NAND2_X1 U13336 ( .A1(n10532), .A2(n10530), .ZN(n10526) );
  NAND2_X1 U13337 ( .A1(n10561), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10521) );
  NAND2_X1 U13338 ( .A1(n15548), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10520) );
  INV_X1 U13339 ( .A(n10523), .ZN(n10522) );
  NAND2_X1 U13340 ( .A1(n10522), .A2(n15515), .ZN(n20490) );
  NAND2_X1 U13341 ( .A1(n10523), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10524) );
  NAND2_X1 U13342 ( .A1(n20490), .A2(n10524), .ZN(n13598) );
  AND2_X1 U13343 ( .A1(n11787), .A2(n13598), .ZN(n10528) );
  NAND2_X1 U13344 ( .A1(n10526), .A2(n10525), .ZN(n10560) );
  INV_X1 U13345 ( .A(n10527), .ZN(n10531) );
  INV_X1 U13346 ( .A(n10528), .ZN(n10529) );
  NAND4_X1 U13347 ( .A1(n10532), .A2(n10531), .A3(n10530), .A4(n10529), .ZN(
        n10533) );
  AOI22_X1 U13348 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10537) );
  AOI22_X1 U13349 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13350 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13351 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13352 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10543) );
  AOI22_X1 U13353 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13354 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13355 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10539) );
  AOI22_X1 U13356 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10538) );
  NAND4_X1 U13357 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10542) );
  INV_X1 U13358 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20166) );
  OAI22_X1 U13359 ( .A1(n11143), .A2(n20166), .B1(n11517), .B2(n10565), .ZN(
        n10544) );
  INV_X1 U13360 ( .A(n10549), .ZN(n10546) );
  NAND2_X1 U13361 ( .A1(n10549), .A2(n10548), .ZN(n10550) );
  XNOR2_X1 U13362 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13530) );
  AOI21_X1 U13363 ( .B1(n13432), .B2(n13530), .A(n11094), .ZN(n10552) );
  NAND2_X1 U13364 ( .A1(n11095), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n10551) );
  OAI211_X1 U13365 ( .C1(n10589), .C2(n13323), .A(n10552), .B(n10551), .ZN(
        n10553) );
  INV_X1 U13366 ( .A(n10553), .ZN(n10554) );
  NAND2_X1 U13367 ( .A1(n11094), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13368 ( .A1(n10555), .A2(n10558), .ZN(n13268) );
  NAND2_X1 U13369 ( .A1(n10561), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10564) );
  NOR3_X1 U13370 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15515), .A3(
        n20531), .ZN(n20375) );
  NAND2_X1 U13371 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20375), .ZN(
        n20394) );
  NAND2_X1 U13372 ( .A1(n20489), .A2(n20394), .ZN(n10562) );
  NAND3_X1 U13373 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20597) );
  INV_X1 U13374 ( .A(n20597), .ZN(n20659) );
  NAND2_X1 U13375 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20659), .ZN(
        n20707) );
  AOI22_X1 U13376 ( .A1(n11787), .A2(n20401), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15548), .ZN(n10563) );
  INV_X1 U13377 ( .A(n11143), .ZN(n11131) );
  AOI22_X1 U13378 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13379 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13380 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10568) );
  INV_X1 U13381 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20173) );
  AOI22_X1 U13382 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10567) );
  NAND4_X1 U13383 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n10576) );
  AOI22_X1 U13384 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13385 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10573) );
  AOI22_X1 U13386 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10572) );
  AOI22_X1 U13387 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10571) );
  NAND4_X1 U13388 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10575) );
  AOI22_X1 U13389 ( .A1(n11131), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11148), .B2(n11545), .ZN(n10577) );
  INV_X1 U13390 ( .A(n10581), .ZN(n10579) );
  NAND2_X2 U13391 ( .A1(n10580), .A2(n10579), .ZN(n10603) );
  NAND2_X1 U13392 ( .A1(n10581), .A2(n13408), .ZN(n10582) );
  INV_X1 U13393 ( .A(n13589), .ZN(n10583) );
  NOR2_X1 U13394 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n10584), .ZN(
        n10585) );
  NOR2_X1 U13395 ( .A1(n10605), .A2(n10585), .ZN(n13564) );
  INV_X1 U13396 ( .A(n11094), .ZN(n10811) );
  INV_X1 U13397 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13560) );
  OAI22_X1 U13398 ( .A1(n13564), .A2(n11093), .B1(n10811), .B2(n13560), .ZN(
        n10586) );
  AOI21_X1 U13399 ( .B1(n11095), .B2(P1_EAX_REG_3__SCAN_IN), .A(n10586), .ZN(
        n10587) );
  OAI211_X1 U13400 ( .C1(n10589), .C2(n10559), .A(n10588), .B(n10587), .ZN(
        n13363) );
  INV_X1 U13401 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13604) );
  OR2_X1 U13402 ( .A1(n11143), .A2(n13604), .ZN(n10601) );
  AOI22_X1 U13403 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U13404 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10680), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10592) );
  AOI22_X1 U13405 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11067), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U13406 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11070), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10590) );
  NAND4_X1 U13407 ( .A1(n10593), .A2(n10592), .A3(n10591), .A4(n10590), .ZN(
        n10599) );
  AOI22_X1 U13408 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n10894), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10597) );
  AOI22_X1 U13409 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10596) );
  AOI22_X1 U13410 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10595) );
  AOI22_X1 U13411 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n11068), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10594) );
  NAND4_X1 U13412 ( .A1(n10597), .A2(n10596), .A3(n10595), .A4(n10594), .ZN(
        n10598) );
  NAND2_X1 U13413 ( .A1(n11148), .A2(n11551), .ZN(n10600) );
  NAND2_X1 U13414 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  NAND2_X1 U13415 ( .A1(n9861), .A2(n10604), .ZN(n11553) );
  INV_X1 U13416 ( .A(n11553), .ZN(n10611) );
  OAI21_X1 U13417 ( .B1(n10605), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n10628), .ZN(n20043) );
  AOI22_X1 U13418 ( .A1(n11095), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20721), .ZN(n10608) );
  NAND2_X1 U13419 ( .A1(n10606), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10607) );
  NAND2_X1 U13420 ( .A1(n10608), .A2(n10607), .ZN(n10609) );
  MUX2_X1 U13421 ( .A(n20043), .B(n10609), .S(n11093), .Z(n10610) );
  AOI21_X1 U13422 ( .B1(n10611), .B2(n10775), .A(n10610), .ZN(n13460) );
  INV_X1 U13423 ( .A(n13460), .ZN(n10612) );
  AOI22_X1 U13424 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10617) );
  AOI22_X1 U13425 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10616) );
  AOI22_X1 U13426 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10615) );
  INV_X1 U13427 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20178) );
  AOI22_X1 U13428 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10614) );
  NAND4_X1 U13429 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10623) );
  AOI22_X1 U13430 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10318), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10621) );
  AOI22_X1 U13431 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10620) );
  AOI22_X1 U13432 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10619) );
  AOI22_X1 U13433 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13434 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10622) );
  NAND2_X1 U13435 ( .A1(n11148), .A2(n11560), .ZN(n10625) );
  OR2_X1 U13436 ( .A1(n11143), .A2(n20178), .ZN(n10624) );
  NAND2_X1 U13437 ( .A1(n9861), .A2(n9898), .ZN(n10626) );
  NAND2_X1 U13438 ( .A1(n10652), .A2(n10626), .ZN(n11557) );
  INV_X1 U13439 ( .A(n11557), .ZN(n10634) );
  AND2_X1 U13440 ( .A1(n10628), .A2(n20033), .ZN(n10629) );
  OR2_X1 U13441 ( .A1(n10629), .A2(n10647), .ZN(n20039) );
  NAND2_X1 U13442 ( .A1(n20039), .A2(n13432), .ZN(n10630) );
  OAI21_X1 U13443 ( .B1(n20033), .B2(n10811), .A(n10630), .ZN(n10631) );
  AOI21_X1 U13444 ( .B1(n11095), .B2(P1_EAX_REG_5__SCAN_IN), .A(n10631), .ZN(
        n10632) );
  INV_X1 U13445 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n10651) );
  AOI22_X1 U13446 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13447 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10637) );
  AOI22_X1 U13448 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U13449 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10635) );
  NAND4_X1 U13450 ( .A1(n10638), .A2(n10637), .A3(n10636), .A4(n10635), .ZN(
        n10644) );
  AOI22_X1 U13451 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10642) );
  AOI22_X1 U13452 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10680), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10641) );
  AOI22_X1 U13453 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10640) );
  AOI22_X1 U13454 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10639) );
  NAND4_X1 U13455 ( .A1(n10642), .A2(n10641), .A3(n10640), .A4(n10639), .ZN(
        n10643) );
  NAND2_X1 U13456 ( .A1(n11148), .A2(n11576), .ZN(n10646) );
  INV_X1 U13457 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20190) );
  OR2_X1 U13458 ( .A1(n11143), .A2(n20190), .ZN(n10645) );
  NAND2_X1 U13459 ( .A1(n10646), .A2(n10645), .ZN(n10653) );
  NAND2_X1 U13460 ( .A1(n10652), .A2(n9992), .ZN(n11568) );
  NAND2_X1 U13461 ( .A1(n11568), .A2(n10775), .ZN(n10650) );
  NOR2_X1 U13462 ( .A1(n10647), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10648) );
  OR2_X1 U13463 ( .A1(n10656), .A2(n10648), .ZN(n20029) );
  AOI22_X1 U13464 ( .A1(n20029), .A2(n10847), .B1(n11094), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10649) );
  INV_X1 U13465 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13611) );
  NAND2_X1 U13466 ( .A1(n11148), .A2(n11588), .ZN(n10654) );
  OAI21_X1 U13467 ( .B1(n13611), .B2(n11143), .A(n10654), .ZN(n10655) );
  INV_X1 U13468 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n10659) );
  NOR2_X1 U13469 ( .A1(n10656), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10657) );
  OR2_X1 U13470 ( .A1(n10675), .A2(n10657), .ZN(n20020) );
  AOI22_X1 U13471 ( .A1(n20020), .A2(n10847), .B1(n11094), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10658) );
  OAI21_X1 U13472 ( .B1(n9913), .B2(n10659), .A(n10658), .ZN(n10660) );
  AOI22_X1 U13473 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13474 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10663) );
  AOI22_X1 U13475 ( .A1(n10982), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10662) );
  AOI22_X1 U13476 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10661) );
  NAND4_X1 U13477 ( .A1(n10664), .A2(n10663), .A3(n10662), .A4(n10661), .ZN(
        n10670) );
  AOI22_X1 U13478 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10668) );
  AOI22_X1 U13479 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10667) );
  AOI22_X1 U13480 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13481 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10665) );
  NAND4_X1 U13482 ( .A1(n10668), .A2(n10667), .A3(n10666), .A4(n10665), .ZN(
        n10669) );
  OAI21_X1 U13483 ( .B1(n10670), .B2(n10669), .A(n10775), .ZN(n10674) );
  NAND2_X1 U13484 ( .A1(n11095), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n10673) );
  XNOR2_X1 U13485 ( .A(n10675), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13760) );
  NAND2_X1 U13486 ( .A1(n13760), .A2(n10847), .ZN(n10672) );
  NAND2_X1 U13487 ( .A1(n11094), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10671) );
  NAND4_X1 U13488 ( .A1(n10674), .A2(n10673), .A3(n10672), .A4(n10671), .ZN(
        n13584) );
  XNOR2_X1 U13489 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n10691), .ZN(
        n13787) );
  AOI22_X1 U13490 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10679) );
  AOI22_X1 U13491 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13492 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10677) );
  AOI22_X1 U13493 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10676) );
  NAND4_X1 U13494 ( .A1(n10679), .A2(n10678), .A3(n10677), .A4(n10676), .ZN(
        n10686) );
  AOI22_X1 U13496 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10684) );
  AOI22_X1 U13497 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10683) );
  AOI22_X1 U13498 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10682) );
  AOI22_X1 U13499 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10681) );
  NAND4_X1 U13500 ( .A1(n10684), .A2(n10683), .A3(n10682), .A4(n10681), .ZN(
        n10685) );
  OR2_X1 U13501 ( .A1(n10686), .A2(n10685), .ZN(n10687) );
  AOI22_X1 U13502 ( .A1(n10775), .A2(n10687), .B1(n11094), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10689) );
  NAND2_X1 U13503 ( .A1(n11095), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n10688) );
  OAI211_X1 U13504 ( .C1(n13787), .C2(n11093), .A(n10689), .B(n10688), .ZN(
        n13636) );
  XNOR2_X1 U13505 ( .A(n10707), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14635) );
  NAND2_X1 U13506 ( .A1(n14635), .A2(n10847), .ZN(n10706) );
  INV_X1 U13507 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14640) );
  AOI22_X1 U13508 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10695) );
  AOI22_X1 U13509 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13510 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13511 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10692) );
  NAND4_X1 U13512 ( .A1(n10695), .A2(n10694), .A3(n10693), .A4(n10692), .ZN(
        n10701) );
  AOI22_X1 U13513 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U13514 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13515 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13516 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10696) );
  NAND4_X1 U13517 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10700) );
  OAI21_X1 U13518 ( .B1(n10701), .B2(n10700), .A(n10775), .ZN(n10703) );
  NAND2_X1 U13519 ( .A1(n11095), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n10702) );
  OAI211_X1 U13520 ( .C1(n10811), .C2(n14640), .A(n10703), .B(n10702), .ZN(
        n10704) );
  INV_X1 U13521 ( .A(n10704), .ZN(n10705) );
  NAND2_X1 U13522 ( .A1(n10706), .A2(n10705), .ZN(n13744) );
  INV_X1 U13523 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10708) );
  XNOR2_X1 U13524 ( .A(n10783), .B(n10708), .ZN(n14619) );
  AOI22_X1 U13525 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10712) );
  AOI22_X1 U13526 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13527 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10710) );
  AOI22_X1 U13528 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10709) );
  NAND4_X1 U13529 ( .A1(n10712), .A2(n10711), .A3(n10710), .A4(n10709), .ZN(
        n10718) );
  AOI22_X1 U13530 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10369), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10716) );
  AOI22_X1 U13531 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10715) );
  AOI22_X1 U13532 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10714) );
  AOI22_X1 U13533 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10713) );
  NAND4_X1 U13534 ( .A1(n10716), .A2(n10715), .A3(n10714), .A4(n10713), .ZN(
        n10717) );
  OAI21_X1 U13535 ( .B1(n10718), .B2(n10717), .A(n10775), .ZN(n10721) );
  NAND2_X1 U13536 ( .A1(n11095), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n10720) );
  NAND2_X1 U13537 ( .A1(n11094), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10719) );
  NAND3_X1 U13538 ( .A1(n10721), .A2(n10720), .A3(n10719), .ZN(n10722) );
  AOI21_X1 U13539 ( .B1(n14619), .B2(n10847), .A(n10722), .ZN(n13800) );
  XOR2_X1 U13540 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n10723), .Z(
        n15748) );
  INV_X1 U13541 ( .A(n15748), .ZN(n10738) );
  AOI22_X1 U13542 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10727) );
  AOI22_X1 U13543 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10726) );
  AOI22_X1 U13544 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10725) );
  AOI22_X1 U13545 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10724) );
  NAND4_X1 U13546 ( .A1(n10727), .A2(n10726), .A3(n10725), .A4(n10724), .ZN(
        n10733) );
  AOI22_X1 U13547 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11029), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10731) );
  AOI22_X1 U13548 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U13549 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10729) );
  AOI22_X1 U13550 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10728) );
  NAND4_X1 U13551 ( .A1(n10731), .A2(n10730), .A3(n10729), .A4(n10728), .ZN(
        n10732) );
  OAI21_X1 U13552 ( .B1(n10733), .B2(n10732), .A(n10775), .ZN(n10736) );
  NAND2_X1 U13553 ( .A1(n11095), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U13554 ( .A1(n11094), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10734) );
  NAND3_X1 U13555 ( .A1(n10736), .A2(n10735), .A3(n10734), .ZN(n10737) );
  AOI21_X1 U13556 ( .B1(n10738), .B2(n13432), .A(n10737), .ZN(n13767) );
  NAND2_X1 U13557 ( .A1(n11095), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n10741) );
  OAI21_X1 U13558 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n10739), .A(
        n10763), .ZN(n15772) );
  AOI22_X1 U13559 ( .A1(n10847), .A2(n15772), .B1(n11094), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10740) );
  NAND2_X1 U13560 ( .A1(n10741), .A2(n10740), .ZN(n13817) );
  AOI22_X1 U13561 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10745) );
  AOI22_X1 U13562 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10744) );
  AOI22_X1 U13563 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U13564 ( .A1(n10680), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10742) );
  NAND4_X1 U13565 ( .A1(n10745), .A2(n10744), .A3(n10743), .A4(n10742), .ZN(
        n10751) );
  AOI22_X1 U13566 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10749) );
  AOI22_X1 U13567 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10748) );
  AOI22_X1 U13568 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10747) );
  AOI22_X1 U13569 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10746) );
  NAND4_X1 U13570 ( .A1(n10749), .A2(n10748), .A3(n10747), .A4(n10746), .ZN(
        n10750) );
  OR2_X1 U13571 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  AND2_X1 U13572 ( .A1(n10775), .A2(n10752), .ZN(n13770) );
  INV_X1 U13573 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U13574 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n11067), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10756) );
  AOI22_X1 U13575 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9829), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10755) );
  AOI22_X1 U13576 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10754) );
  AOI22_X1 U13577 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10328), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10753) );
  NAND4_X1 U13578 ( .A1(n10756), .A2(n10755), .A3(n10754), .A4(n10753), .ZN(
        n10762) );
  AOI22_X1 U13579 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10760) );
  AOI22_X1 U13580 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10759) );
  AOI22_X1 U13581 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10758) );
  AOI22_X1 U13582 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10855), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10757) );
  NAND4_X1 U13583 ( .A1(n10760), .A2(n10759), .A3(n10758), .A4(n10757), .ZN(
        n10761) );
  OAI21_X1 U13584 ( .B1(n10762), .B2(n10761), .A(n10775), .ZN(n10766) );
  XNOR2_X1 U13585 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n10763), .ZN(
        n15759) );
  OAI22_X1 U13586 ( .A1(n15759), .A2(n11093), .B1(n10811), .B2(n15689), .ZN(
        n10764) );
  INV_X1 U13587 ( .A(n10764), .ZN(n10765) );
  OAI211_X1 U13588 ( .C1(n9913), .C2(n13823), .A(n10766), .B(n10765), .ZN(
        n13821) );
  INV_X1 U13589 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14503) );
  AOI22_X1 U13590 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10770) );
  AOI22_X1 U13591 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10769) );
  AOI22_X1 U13592 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9825), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10768) );
  AOI22_X1 U13593 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10767) );
  NAND4_X1 U13594 ( .A1(n10770), .A2(n10769), .A3(n10768), .A4(n10767), .ZN(
        n10777) );
  AOI22_X1 U13595 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10774) );
  AOI22_X1 U13596 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10773) );
  AOI22_X1 U13597 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10772) );
  AOI22_X1 U13598 ( .A1(n9829), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10771) );
  NAND4_X1 U13599 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n10771), .ZN(
        n10776) );
  OAI21_X1 U13600 ( .B1(n10777), .B2(n10776), .A(n10775), .ZN(n10781) );
  INV_X1 U13601 ( .A(n10778), .ZN(n10779) );
  XNOR2_X1 U13602 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n10779), .ZN(
        n14631) );
  AOI22_X1 U13603 ( .A1(n10847), .A2(n14631), .B1(n11094), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10780) );
  OAI211_X1 U13604 ( .C1(n9913), .C2(n14503), .A(n10781), .B(n10780), .ZN(
        n14391) );
  OAI211_X1 U13605 ( .C1(n13817), .C2(n13770), .A(n13821), .B(n14391), .ZN(
        n13766) );
  OR2_X1 U13606 ( .A1(n13767), .A2(n13766), .ZN(n13765) );
  OR2_X1 U13607 ( .A1(n10784), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10785) );
  NAND2_X1 U13608 ( .A1(n10785), .A2(n10829), .ZN(n15741) );
  INV_X1 U13609 ( .A(n15741), .ZN(n15663) );
  AOI22_X1 U13610 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10789) );
  AOI22_X1 U13611 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10788) );
  AOI22_X1 U13612 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10787) );
  AOI22_X1 U13613 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10786) );
  NAND4_X1 U13614 ( .A1(n10789), .A2(n10788), .A3(n10787), .A4(n10786), .ZN(
        n10795) );
  AOI22_X1 U13615 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10793) );
  AOI22_X1 U13616 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10792) );
  AOI22_X1 U13617 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10791) );
  AOI22_X1 U13618 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10790) );
  NAND4_X1 U13619 ( .A1(n10793), .A2(n10792), .A3(n10791), .A4(n10790), .ZN(
        n10794) );
  OR2_X1 U13620 ( .A1(n10795), .A2(n10794), .ZN(n10798) );
  INV_X1 U13621 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13778) );
  NAND2_X1 U13622 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10796) );
  OAI211_X1 U13623 ( .C1(n9913), .C2(n13778), .A(n11093), .B(n10796), .ZN(
        n10797) );
  AOI21_X1 U13624 ( .B1(n11058), .B2(n10798), .A(n10797), .ZN(n10799) );
  AOI21_X1 U13625 ( .B1(n15663), .B2(n10847), .A(n10799), .ZN(n13776) );
  AOI22_X1 U13626 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10803) );
  AOI22_X1 U13627 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10802) );
  AOI22_X1 U13628 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10801) );
  AOI22_X1 U13629 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10800) );
  NAND4_X1 U13630 ( .A1(n10803), .A2(n10802), .A3(n10801), .A4(n10800), .ZN(
        n10809) );
  AOI22_X1 U13631 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10807) );
  AOI22_X1 U13632 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10806) );
  AOI22_X1 U13633 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10805) );
  AOI22_X1 U13634 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10804) );
  NAND4_X1 U13635 ( .A1(n10807), .A2(n10806), .A3(n10805), .A4(n10804), .ZN(
        n10808) );
  OR2_X1 U13636 ( .A1(n10809), .A2(n10808), .ZN(n10810) );
  NAND2_X1 U13637 ( .A1(n11058), .A2(n10810), .ZN(n10814) );
  XNOR2_X1 U13638 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n10829), .ZN(
        n14609) );
  INV_X1 U13639 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14607) );
  OAI22_X1 U13640 ( .A1(n11093), .A2(n14609), .B1(n10811), .B2(n14607), .ZN(
        n10812) );
  AOI21_X1 U13641 ( .B1(n11095), .B2(P1_EAX_REG_17__SCAN_IN), .A(n10812), .ZN(
        n10813) );
  NAND2_X1 U13642 ( .A1(n10814), .A2(n10813), .ZN(n13824) );
  AOI22_X1 U13643 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13644 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10817) );
  AOI22_X1 U13645 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10816) );
  AOI22_X1 U13646 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10815) );
  NAND4_X1 U13647 ( .A1(n10818), .A2(n10817), .A3(n10816), .A4(n10815), .ZN(
        n10824) );
  AOI22_X1 U13648 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10822) );
  AOI22_X1 U13649 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10821) );
  AOI22_X1 U13650 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10820) );
  AOI22_X1 U13651 ( .A1(n10982), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10819) );
  NAND4_X1 U13652 ( .A1(n10822), .A2(n10821), .A3(n10820), .A4(n10819), .ZN(
        n10823) );
  NOR2_X1 U13653 ( .A1(n10824), .A2(n10823), .ZN(n10828) );
  NAND2_X1 U13654 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10825) );
  NAND2_X1 U13655 ( .A1(n11093), .A2(n10825), .ZN(n10826) );
  AOI21_X1 U13656 ( .B1(n11095), .B2(P1_EAX_REG_18__SCAN_IN), .A(n10826), .ZN(
        n10827) );
  OAI21_X1 U13657 ( .B1(n11090), .B2(n10828), .A(n10827), .ZN(n10832) );
  OAI21_X1 U13658 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10830), .A(
        n10852), .ZN(n15656) );
  OR2_X1 U13659 ( .A1(n11093), .A2(n15656), .ZN(n10831) );
  AOI22_X1 U13660 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10836) );
  AOI22_X1 U13661 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13662 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10834) );
  AOI22_X1 U13663 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10833) );
  NAND4_X1 U13664 ( .A1(n10836), .A2(n10835), .A3(n10834), .A4(n10833), .ZN(
        n10842) );
  AOI22_X1 U13665 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10840) );
  AOI22_X1 U13666 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10839) );
  AOI22_X1 U13667 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10838) );
  AOI22_X1 U13668 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10837) );
  NAND4_X1 U13669 ( .A1(n10840), .A2(n10839), .A3(n10838), .A4(n10837), .ZN(
        n10841) );
  NOR2_X1 U13670 ( .A1(n10842), .A2(n10841), .ZN(n10846) );
  NAND2_X1 U13671 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10843) );
  NAND2_X1 U13672 ( .A1(n11093), .A2(n10843), .ZN(n10844) );
  AOI21_X1 U13673 ( .B1(n11095), .B2(P1_EAX_REG_19__SCAN_IN), .A(n10844), .ZN(
        n10845) );
  OAI21_X1 U13674 ( .B1(n11090), .B2(n10846), .A(n10845), .ZN(n10849) );
  XNOR2_X1 U13675 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n10852), .ZN(
        n15632) );
  NAND2_X1 U13676 ( .A1(n15632), .A2(n10847), .ZN(n10848) );
  NAND2_X1 U13677 ( .A1(n10849), .A2(n10848), .ZN(n14432) );
  INV_X1 U13678 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10851) );
  OR2_X1 U13679 ( .A1(n10853), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10854) );
  NAND2_X1 U13680 ( .A1(n10854), .A2(n10887), .ZN(n15727) );
  AOI22_X1 U13681 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n11051), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10859) );
  AOI22_X1 U13682 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10894), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13683 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n10855), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10857) );
  AOI22_X1 U13684 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11070), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10856) );
  NAND4_X1 U13685 ( .A1(n10859), .A2(n10858), .A3(n10857), .A4(n10856), .ZN(
        n10865) );
  AOI22_X1 U13686 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U13687 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10862) );
  AOI22_X1 U13688 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10861) );
  AOI22_X1 U13689 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10860) );
  NAND4_X1 U13690 ( .A1(n10863), .A2(n10862), .A3(n10861), .A4(n10860), .ZN(
        n10864) );
  NOR2_X1 U13691 ( .A1(n10865), .A2(n10864), .ZN(n10866) );
  NOR2_X1 U13692 ( .A1(n11090), .A2(n10866), .ZN(n10869) );
  INV_X1 U13693 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14481) );
  NAND2_X1 U13694 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10867) );
  OAI211_X1 U13695 ( .C1(n9913), .C2(n14481), .A(n11093), .B(n10867), .ZN(
        n10868) );
  OAI22_X1 U13696 ( .A1(n15727), .A2(n11093), .B1(n10869), .B2(n10868), .ZN(
        n14383) );
  AOI22_X1 U13697 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10873) );
  AOI22_X1 U13698 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10872) );
  AOI22_X1 U13699 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10871) );
  AOI22_X1 U13700 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10870) );
  NAND4_X1 U13701 ( .A1(n10873), .A2(n10872), .A3(n10871), .A4(n10870), .ZN(
        n10879) );
  AOI22_X1 U13702 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10877) );
  AOI22_X1 U13703 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10876) );
  AOI22_X1 U13704 ( .A1(n13325), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10875) );
  AOI22_X1 U13705 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10874) );
  NAND4_X1 U13706 ( .A1(n10877), .A2(n10876), .A3(n10875), .A4(n10874), .ZN(
        n10878) );
  NOR2_X1 U13707 ( .A1(n10879), .A2(n10878), .ZN(n10883) );
  NAND2_X1 U13708 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10880) );
  NAND2_X1 U13709 ( .A1(n11093), .A2(n10880), .ZN(n10881) );
  AOI21_X1 U13710 ( .B1(n11095), .B2(P1_EAX_REG_21__SCAN_IN), .A(n10881), .ZN(
        n10882) );
  OAI21_X1 U13711 ( .B1(n11090), .B2(n10883), .A(n10882), .ZN(n10885) );
  XNOR2_X1 U13712 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n10887), .ZN(
        n15626) );
  NAND2_X1 U13713 ( .A1(n15626), .A2(n13432), .ZN(n10884) );
  INV_X1 U13714 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10886) );
  OR2_X1 U13715 ( .A1(n10888), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10889) );
  NAND2_X1 U13716 ( .A1(n10889), .A2(n10949), .ZN(n15726) );
  INV_X1 U13717 ( .A(n15726), .ZN(n10905) );
  AOI22_X1 U13718 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13719 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10892) );
  AOI22_X1 U13720 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10891) );
  AOI22_X1 U13721 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10890) );
  NAND4_X1 U13722 ( .A1(n10893), .A2(n10892), .A3(n10891), .A4(n10890), .ZN(
        n10900) );
  AOI22_X1 U13723 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10898) );
  AOI22_X1 U13724 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U13725 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10896) );
  AOI22_X1 U13726 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10895) );
  NAND4_X1 U13727 ( .A1(n10898), .A2(n10897), .A3(n10896), .A4(n10895), .ZN(
        n10899) );
  OR2_X1 U13728 ( .A1(n10900), .A2(n10899), .ZN(n10903) );
  INV_X1 U13729 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14474) );
  NAND2_X1 U13730 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10901) );
  OAI211_X1 U13731 ( .C1(n9913), .C2(n14474), .A(n11093), .B(n10901), .ZN(
        n10902) );
  AOI21_X1 U13732 ( .B1(n11058), .B2(n10903), .A(n10902), .ZN(n10904) );
  AOI21_X1 U13733 ( .B1(n10905), .B2(n13432), .A(n10904), .ZN(n14472) );
  AOI22_X1 U13734 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11029), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10910) );
  AOI22_X1 U13735 ( .A1(n11030), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10369), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10909) );
  AOI22_X1 U13736 ( .A1(n10906), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10908) );
  AOI22_X1 U13737 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10907) );
  NAND4_X1 U13738 ( .A1(n10910), .A2(n10909), .A3(n10908), .A4(n10907), .ZN(
        n10916) );
  AOI22_X1 U13739 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13740 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10913) );
  AOI22_X1 U13741 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10912) );
  AOI22_X1 U13742 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10911) );
  NAND4_X1 U13743 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(
        n10915) );
  NOR2_X1 U13744 ( .A1(n10916), .A2(n10915), .ZN(n10933) );
  AOI22_X1 U13745 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13746 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10919) );
  AOI22_X1 U13747 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10918) );
  AOI22_X1 U13748 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10917) );
  NAND4_X1 U13749 ( .A1(n10920), .A2(n10919), .A3(n10918), .A4(n10917), .ZN(
        n10926) );
  AOI22_X1 U13750 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11029), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13751 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13752 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10922) );
  AOI22_X1 U13753 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10921) );
  NAND4_X1 U13754 ( .A1(n10924), .A2(n10923), .A3(n10922), .A4(n10921), .ZN(
        n10925) );
  NOR2_X1 U13755 ( .A1(n10926), .A2(n10925), .ZN(n10934) );
  XOR2_X1 U13756 ( .A(n10933), .B(n10934), .Z(n10927) );
  NAND2_X1 U13757 ( .A1(n10927), .A2(n11058), .ZN(n10930) );
  INV_X1 U13758 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15609) );
  OAI21_X1 U13759 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15609), .A(n11093), 
        .ZN(n10928) );
  AOI21_X1 U13760 ( .B1(n11095), .B2(P1_EAX_REG_23__SCAN_IN), .A(n10928), .ZN(
        n10929) );
  NAND2_X1 U13761 ( .A1(n10930), .A2(n10929), .ZN(n10932) );
  XNOR2_X1 U13762 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n10949), .ZN(
        n15606) );
  NAND2_X1 U13763 ( .A1(n15606), .A2(n13432), .ZN(n10931) );
  NAND2_X1 U13764 ( .A1(n10932), .A2(n10931), .ZN(n14418) );
  NOR2_X1 U13765 ( .A1(n10934), .A2(n10933), .ZN(n10958) );
  AOI22_X1 U13766 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U13767 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13768 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13769 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10936) );
  NAND4_X1 U13770 ( .A1(n10939), .A2(n10938), .A3(n10937), .A4(n10936), .ZN(
        n10945) );
  AOI22_X1 U13771 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13772 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U13773 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10941) );
  AOI22_X1 U13774 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10940) );
  NAND4_X1 U13775 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(
        n10944) );
  OR2_X1 U13776 ( .A1(n10945), .A2(n10944), .ZN(n10957) );
  XNOR2_X1 U13777 ( .A(n10958), .B(n10957), .ZN(n10948) );
  INV_X1 U13778 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14377) );
  AOI21_X1 U13779 ( .B1(n14377), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n10946) );
  AOI21_X1 U13780 ( .B1(n11095), .B2(P1_EAX_REG_24__SCAN_IN), .A(n10946), .ZN(
        n10947) );
  OAI21_X1 U13781 ( .B1(n10948), .B2(n11090), .A(n10947), .ZN(n10955) );
  INV_X1 U13782 ( .A(n10951), .ZN(n10952) );
  NAND2_X1 U13783 ( .A1(n10952), .A2(n14377), .ZN(n10953) );
  AND2_X1 U13784 ( .A1(n10994), .A2(n10953), .ZN(n14372) );
  NAND2_X1 U13785 ( .A1(n14372), .A2(n13432), .ZN(n10954) );
  NAND2_X1 U13786 ( .A1(n10955), .A2(n10954), .ZN(n14369) );
  NAND2_X1 U13787 ( .A1(n10958), .A2(n10957), .ZN(n10975) );
  AOI22_X1 U13788 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10962) );
  AOI22_X1 U13789 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U13790 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U13791 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10959) );
  NAND4_X1 U13792 ( .A1(n10962), .A2(n10961), .A3(n10960), .A4(n10959), .ZN(
        n10968) );
  AOI22_X1 U13793 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11029), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10966) );
  AOI22_X1 U13794 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U13795 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U13796 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10963) );
  NAND4_X1 U13797 ( .A1(n10966), .A2(n10965), .A3(n10964), .A4(n10963), .ZN(
        n10967) );
  NOR2_X1 U13798 ( .A1(n10968), .A2(n10967), .ZN(n10976) );
  XOR2_X1 U13799 ( .A(n10975), .B(n10976), .Z(n10969) );
  NAND2_X1 U13800 ( .A1(n10969), .A2(n11058), .ZN(n10974) );
  NAND2_X1 U13801 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10970) );
  NAND2_X1 U13802 ( .A1(n11093), .A2(n10970), .ZN(n10971) );
  AOI21_X1 U13803 ( .B1(n11095), .B2(P1_EAX_REG_25__SCAN_IN), .A(n10971), .ZN(
        n10973) );
  XNOR2_X1 U13804 ( .A(n10994), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14559) );
  AOI21_X1 U13805 ( .B1(n10974), .B2(n10973), .A(n10972), .ZN(n14355) );
  AND2_X2 U13806 ( .A1(n9837), .A2(n14355), .ZN(n14353) );
  NOR2_X1 U13807 ( .A1(n10976), .A2(n10975), .ZN(n11002) );
  AOI22_X1 U13808 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U13809 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10979) );
  AOI22_X1 U13810 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U13811 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10977) );
  NAND4_X1 U13812 ( .A1(n10980), .A2(n10979), .A3(n10978), .A4(n10977), .ZN(
        n10989) );
  AOI22_X1 U13813 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U13814 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U13815 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U13816 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10984) );
  NAND4_X1 U13817 ( .A1(n10987), .A2(n10986), .A3(n10985), .A4(n10984), .ZN(
        n10988) );
  OR2_X1 U13818 ( .A1(n10989), .A2(n10988), .ZN(n11001) );
  INV_X1 U13819 ( .A(n11001), .ZN(n10990) );
  XNOR2_X1 U13820 ( .A(n11002), .B(n10990), .ZN(n10991) );
  NAND2_X1 U13821 ( .A1(n10991), .A2(n11058), .ZN(n11000) );
  NAND2_X1 U13822 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10992) );
  NAND2_X1 U13823 ( .A1(n11093), .A2(n10992), .ZN(n10993) );
  AOI21_X1 U13824 ( .B1(n11095), .B2(P1_EAX_REG_26__SCAN_IN), .A(n10993), .ZN(
        n10999) );
  INV_X1 U13825 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14554) );
  INV_X1 U13826 ( .A(n10995), .ZN(n10996) );
  INV_X1 U13827 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U13828 ( .A1(n10996), .A2(n14343), .ZN(n10997) );
  NAND2_X1 U13829 ( .A1(n11021), .A2(n10997), .ZN(n14543) );
  NOR2_X1 U13830 ( .A1(n14543), .A2(n11093), .ZN(n10998) );
  AOI21_X1 U13831 ( .B1(n11000), .B2(n10999), .A(n10998), .ZN(n14340) );
  NAND2_X1 U13832 ( .A1(n11002), .A2(n11001), .ZN(n11027) );
  AOI22_X1 U13833 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n11070), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U13834 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n11067), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U13835 ( .A1(n10369), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U13836 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11003) );
  NAND4_X1 U13837 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(
        n11013) );
  AOI22_X1 U13838 ( .A1(n11007), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11051), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11011) );
  AOI22_X1 U13839 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U13840 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11009) );
  AOI22_X1 U13841 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11008) );
  NAND4_X1 U13842 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11012) );
  NOR2_X1 U13843 ( .A1(n11013), .A2(n11012), .ZN(n11028) );
  XOR2_X1 U13844 ( .A(n11027), .B(n11028), .Z(n11014) );
  NAND2_X1 U13845 ( .A1(n11014), .A2(n11058), .ZN(n11018) );
  NAND2_X1 U13846 ( .A1(n20721), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U13847 ( .A1(n11093), .A2(n11015), .ZN(n11016) );
  AOI21_X1 U13848 ( .B1(n11095), .B2(P1_EAX_REG_27__SCAN_IN), .A(n11016), .ZN(
        n11017) );
  NAND2_X1 U13849 ( .A1(n11018), .A2(n11017), .ZN(n11020) );
  XNOR2_X1 U13850 ( .A(n11021), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14532) );
  NAND2_X1 U13851 ( .A1(n14532), .A2(n13432), .ZN(n11019) );
  NAND2_X1 U13852 ( .A1(n11020), .A2(n11019), .ZN(n14327) );
  INV_X1 U13853 ( .A(n11021), .ZN(n11022) );
  INV_X1 U13854 ( .A(n11023), .ZN(n11025) );
  INV_X1 U13855 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U13856 ( .A1(n11025), .A2(n11024), .ZN(n11026) );
  NAND2_X1 U13857 ( .A1(n11062), .A2(n11026), .ZN(n14525) );
  NOR2_X1 U13858 ( .A1(n11028), .A2(n11027), .ZN(n11046) );
  AOI22_X1 U13859 ( .A1(n11029), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10935), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U13860 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11030), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U13861 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11032) );
  AOI22_X1 U13862 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11031) );
  NAND4_X1 U13863 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11040) );
  AOI22_X1 U13864 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10855), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11038) );
  AOI22_X1 U13865 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11037) );
  AOI22_X1 U13866 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11036) );
  AOI22_X1 U13867 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11035) );
  NAND4_X1 U13868 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(
        n11039) );
  OR2_X1 U13869 ( .A1(n11040), .A2(n11039), .ZN(n11045) );
  XNOR2_X1 U13870 ( .A(n11046), .B(n11045), .ZN(n11043) );
  AOI21_X1 U13871 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n20721), .A(
        n13432), .ZN(n11042) );
  NAND2_X1 U13872 ( .A1(n11095), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n11041) );
  OAI211_X1 U13873 ( .C1(n11043), .C2(n11090), .A(n11042), .B(n11041), .ZN(
        n11044) );
  OAI21_X1 U13874 ( .B1(n11093), .B2(n14525), .A(n11044), .ZN(n14315) );
  NAND2_X1 U13875 ( .A1(n11046), .A2(n11045), .ZN(n11084) );
  AOI22_X1 U13876 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11029), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U13877 ( .A1(n11065), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11049) );
  AOI22_X1 U13878 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11048) );
  AOI22_X1 U13879 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11047) );
  NAND4_X1 U13880 ( .A1(n11050), .A2(n11049), .A3(n11048), .A4(n11047), .ZN(
        n11057) );
  AOI22_X1 U13881 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11068), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U13882 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11077), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U13883 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11053) );
  AOI22_X1 U13884 ( .A1(n11067), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U13885 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n11056) );
  NOR2_X1 U13886 ( .A1(n11057), .A2(n11056), .ZN(n11085) );
  XOR2_X1 U13887 ( .A(n11084), .B(n11085), .Z(n11059) );
  NAND2_X1 U13888 ( .A1(n11059), .A2(n11058), .ZN(n11064) );
  INV_X1 U13889 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14310) );
  AOI21_X1 U13890 ( .B1(n14310), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n11060) );
  AOI21_X1 U13891 ( .B1(n11095), .B2(P1_EAX_REG_29__SCAN_IN), .A(n11060), .ZN(
        n11063) );
  INV_X1 U13892 ( .A(n11062), .ZN(n11061) );
  AOI21_X1 U13893 ( .B1(n11062), .B2(n14310), .A(n13435), .ZN(n14307) );
  AOI22_X1 U13894 ( .A1(n11064), .A2(n11063), .B1(n13432), .B2(n14307), .ZN(
        n11784) );
  XNOR2_X1 U13895 ( .A(n13435), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14512) );
  AOI22_X1 U13896 ( .A1(n11066), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11065), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U13897 ( .A1(n11068), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11067), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U13898 ( .A1(n10894), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U13899 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11069), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U13900 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n11083) );
  AOI22_X1 U13901 ( .A1(n10935), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11029), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U13902 ( .A1(n10855), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13325), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U13903 ( .A1(n11051), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11076), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U13904 ( .A1(n11077), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11078) );
  NAND4_X1 U13905 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11082) );
  NOR2_X1 U13906 ( .A1(n11083), .A2(n11082), .ZN(n11087) );
  NOR2_X1 U13907 ( .A1(n11085), .A2(n11084), .ZN(n11086) );
  XOR2_X1 U13908 ( .A(n11087), .B(n11086), .Z(n11091) );
  AOI21_X1 U13909 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20721), .A(
        n13432), .ZN(n11089) );
  NAND2_X1 U13910 ( .A1(n11095), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n11088) );
  OAI211_X1 U13911 ( .C1(n11091), .C2(n11090), .A(n11089), .B(n11088), .ZN(
        n11092) );
  OAI21_X1 U13912 ( .B1(n11093), .B2(n14512), .A(n11092), .ZN(n14292) );
  AOI22_X1 U13913 ( .A1(n11095), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n11094), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11096) );
  XNOR2_X1 U13914 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11119) );
  NAND2_X1 U13915 ( .A1(n20570), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11105) );
  NAND2_X1 U13916 ( .A1(n11119), .A2(n11118), .ZN(n11099) );
  NAND2_X1 U13917 ( .A1(n20531), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11098) );
  NAND2_X1 U13918 ( .A1(n11099), .A2(n11098), .ZN(n11128) );
  MUX2_X1 U13919 ( .A(n15515), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11127) );
  NAND2_X1 U13920 ( .A1(n11128), .A2(n11127), .ZN(n11101) );
  NAND2_X1 U13921 ( .A1(n15515), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11100) );
  MUX2_X1 U13922 ( .A(n20489), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11103) );
  NOR2_X1 U13923 ( .A1(n10559), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11102) );
  NOR2_X1 U13924 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20148), .ZN(
        n11145) );
  XNOR2_X1 U13925 ( .A(n11104), .B(n11103), .ZN(n11155) );
  NAND2_X1 U13926 ( .A1(n11143), .A2(n11155), .ZN(n11141) );
  OAI21_X1 U13927 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20570), .A(
        n11105), .ZN(n11109) );
  INV_X1 U13928 ( .A(n11151), .ZN(n11106) );
  OAI21_X1 U13929 ( .B1(n11130), .B2(n11109), .A(n11106), .ZN(n11113) );
  INV_X1 U13930 ( .A(n11129), .ZN(n11108) );
  OAI211_X1 U13931 ( .C1(n11115), .C2(n20156), .A(n11108), .B(n11107), .ZN(
        n11111) );
  INV_X1 U13932 ( .A(n11109), .ZN(n11110) );
  NAND2_X1 U13933 ( .A1(n11111), .A2(n11110), .ZN(n11112) );
  NAND2_X1 U13934 ( .A1(n11113), .A2(n11112), .ZN(n11122) );
  INV_X1 U13935 ( .A(n11122), .ZN(n11126) );
  OAI21_X1 U13936 ( .B1(n13442), .B2(n11114), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11117) );
  NAND2_X1 U13937 ( .A1(n11115), .A2(n13447), .ZN(n11116) );
  NAND2_X1 U13938 ( .A1(n11117), .A2(n11116), .ZN(n11120) );
  XNOR2_X1 U13939 ( .A(n11119), .B(n11118), .ZN(n11157) );
  INV_X1 U13940 ( .A(n11123), .ZN(n11125) );
  AOI21_X1 U13941 ( .B1(n11131), .B2(n11157), .A(n11120), .ZN(n11121) );
  AOI21_X1 U13942 ( .B1(n11123), .B2(n11122), .A(n11121), .ZN(n11124) );
  AOI21_X1 U13943 ( .B1(n11126), .B2(n11125), .A(n11124), .ZN(n11137) );
  XNOR2_X1 U13944 ( .A(n11128), .B(n11127), .ZN(n11156) );
  NOR2_X1 U13945 ( .A1(n11129), .A2(n13447), .ZN(n11133) );
  AOI211_X1 U13946 ( .C1(n11131), .C2(n11156), .A(n11133), .B(n11132), .ZN(
        n11136) );
  INV_X1 U13947 ( .A(n11132), .ZN(n11135) );
  INV_X1 U13948 ( .A(n11133), .ZN(n11134) );
  OAI22_X1 U13949 ( .A1(n11137), .A2(n11136), .B1(n11135), .B2(n11134), .ZN(
        n11140) );
  INV_X1 U13950 ( .A(n11138), .ZN(n11139) );
  AOI222_X1 U13951 ( .A1(n11141), .A2(n11140), .B1(n11139), .B2(n11158), .C1(
        n11155), .C2(n11151), .ZN(n11142) );
  AOI21_X1 U13952 ( .B1(n11158), .B2(n11143), .A(n11142), .ZN(n11144) );
  AOI21_X1 U13953 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20718), .A(
        n11144), .ZN(n11150) );
  NAND2_X1 U13954 ( .A1(n20148), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11146) );
  AOI21_X1 U13955 ( .B1(n11147), .B2(n11146), .A(n11145), .ZN(n11160) );
  NAND2_X1 U13956 ( .A1(n11160), .A2(n11148), .ZN(n11149) );
  NAND2_X1 U13957 ( .A1(n11150), .A2(n11149), .ZN(n11153) );
  NAND2_X1 U13958 ( .A1(n11151), .A2(n11160), .ZN(n11152) );
  NAND2_X1 U13959 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20800) );
  INV_X1 U13960 ( .A(n20800), .ZN(n15563) );
  AOI21_X1 U13961 ( .B1(n10401), .B2(n20149), .A(n10403), .ZN(n11639) );
  NAND2_X1 U13962 ( .A1(n11639), .A2(n13439), .ZN(n13313) );
  NOR4_X1 U13963 ( .A1(n11158), .A2(n11157), .A3(n11156), .A4(n11155), .ZN(
        n11159) );
  OR2_X1 U13964 ( .A1(n11160), .A2(n11159), .ZN(n12964) );
  OR2_X1 U13965 ( .A1(n12964), .A2(n15563), .ZN(n11161) );
  OAI22_X1 U13966 ( .A1(n13155), .A2(n13313), .B1(n11154), .B2(n11161), .ZN(
        n11162) );
  INV_X1 U13967 ( .A(n11162), .ZN(n11163) );
  NOR2_X1 U13968 ( .A1(n13596), .A2(n13128), .ZN(n11165) );
  NOR2_X1 U13969 ( .A1(n13608), .A2(n11531), .ZN(n11164) );
  NAND4_X1 U13970 ( .A1(n13328), .A2(n11165), .A3(n11164), .A4(n10325), .ZN(
        n13130) );
  INV_X1 U13971 ( .A(n13608), .ZN(n13133) );
  AND2_X1 U13972 ( .A1(n14502), .A2(n13133), .ZN(n11168) );
  NOR4_X1 U13973 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n11172) );
  NOR4_X1 U13974 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n11171) );
  NOR4_X1 U13975 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n11170) );
  NOR4_X1 U13976 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n11169) );
  AND4_X1 U13977 ( .A1(n11172), .A2(n11171), .A3(n11170), .A4(n11169), .ZN(
        n11177) );
  NOR4_X1 U13978 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n11175) );
  NOR4_X1 U13979 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n11174) );
  NOR4_X1 U13980 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n11173) );
  INV_X1 U13981 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20738) );
  AND4_X1 U13982 ( .A1(n11175), .A2(n11174), .A3(n11173), .A4(n20738), .ZN(
        n11176) );
  NAND2_X1 U13983 ( .A1(n11177), .A2(n11176), .ZN(n11178) );
  AND2_X2 U13984 ( .A1(n11178), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n13593)
         );
  INV_X1 U13985 ( .A(n13593), .ZN(n13594) );
  NOR2_X1 U13986 ( .A1(n10390), .A2(n13594), .ZN(n11179) );
  NAND2_X1 U13987 ( .A1(n14502), .A2(n11179), .ZN(n14493) );
  INV_X1 U13988 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16375) );
  NOR2_X1 U13989 ( .A1(n14493), .A2(n16375), .ZN(n11183) );
  NOR3_X1 U13990 ( .A1(n14487), .A2(n13593), .A3(n10390), .ZN(n11180) );
  AOI22_X1 U13991 ( .A1(n14496), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14487), .ZN(n11181) );
  INV_X1 U13992 ( .A(n11181), .ZN(n11182) );
  NOR2_X1 U13993 ( .A1(n11183), .A2(n11182), .ZN(n11184) );
  AOI22_X1 U13994 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11189) );
  AOI22_X1 U13995 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11188) );
  AOI22_X1 U13996 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11187) );
  AOI22_X1 U13997 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11186) );
  NAND4_X1 U13998 ( .A1(n11189), .A2(n11188), .A3(n11187), .A4(n11186), .ZN(
        n11199) );
  AOI22_X1 U13999 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11197) );
  NOR2_X2 U14000 ( .A1(n18601), .A2(n15463), .ZN(n17064) );
  AOI22_X1 U14001 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11196) );
  OR3_X2 U14002 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n16856), .ZN(n11369) );
  INV_X4 U14003 ( .A(n11369), .ZN(n17141) );
  AOI22_X1 U14004 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11195) );
  NOR4_X2 U14005 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(n18789), .A4(n18764), .ZN(
        n11227) );
  AOI22_X1 U14006 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11194) );
  NAND4_X1 U14007 ( .A1(n11197), .A2(n11196), .A3(n11195), .A4(n11194), .ZN(
        n11198) );
  AOI22_X1 U14008 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14009 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14010 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14011 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11200) );
  NAND4_X1 U14012 ( .A1(n11203), .A2(n11202), .A3(n11201), .A4(n11200), .ZN(
        n11209) );
  AOI22_X1 U14013 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11207) );
  AOI22_X1 U14014 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11206) );
  AOI22_X1 U14015 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11205) );
  AOI22_X1 U14016 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11204) );
  NAND4_X1 U14017 ( .A1(n11207), .A2(n11206), .A3(n11205), .A4(n11204), .ZN(
        n11208) );
  AOI22_X1 U14018 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11213) );
  AOI22_X1 U14019 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14020 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14021 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11327), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11210) );
  NAND4_X1 U14022 ( .A1(n11213), .A2(n11212), .A3(n11211), .A4(n11210), .ZN(
        n11219) );
  AOI22_X1 U14023 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11217) );
  AOI22_X1 U14024 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14025 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14026 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11214) );
  NAND4_X1 U14027 ( .A1(n11217), .A2(n11216), .A3(n11215), .A4(n11214), .ZN(
        n11218) );
  AOI22_X1 U14028 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11226) );
  INV_X1 U14029 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17192) );
  AOI22_X1 U14030 ( .A1(n11249), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11327), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11220) );
  OAI21_X1 U14031 ( .B1(n11326), .B2(n17192), .A(n11220), .ZN(n11222) );
  NOR2_X1 U14032 ( .A1(n11222), .A2(n11221), .ZN(n11225) );
  AOI22_X1 U14033 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11223), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11224) );
  NAND3_X1 U14034 ( .A1(n11226), .A2(n11225), .A3(n11224), .ZN(n11233) );
  AOI22_X1 U14035 ( .A1(n17141), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11231) );
  AOI22_X1 U14036 ( .A1(n11227), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11245), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14037 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11271), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14038 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11228) );
  NAND4_X1 U14039 ( .A1(n11231), .A2(n11230), .A3(n11229), .A4(n11228), .ZN(
        n11232) );
  INV_X1 U14040 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17107) );
  AOI22_X1 U14041 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14042 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11234), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11235) );
  OAI211_X1 U14043 ( .C1(n11237), .C2(n17107), .A(n11236), .B(n11235), .ZN(
        n11243) );
  AOI22_X1 U14044 ( .A1(n11272), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11271), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14045 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11327), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14046 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14047 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11238) );
  NAND4_X1 U14048 ( .A1(n11241), .A2(n11240), .A3(n11239), .A4(n11238), .ZN(
        n11242) );
  AOI22_X1 U14049 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11244) );
  NAND2_X1 U14050 ( .A1(n11283), .A2(n11449), .ZN(n11457) );
  AOI22_X1 U14051 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11257) );
  INV_X1 U14052 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14053 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11247) );
  AOI22_X1 U14054 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11246) );
  OAI211_X1 U14055 ( .C1(n11237), .C2(n11248), .A(n11247), .B(n11246), .ZN(
        n11255) );
  AOI22_X1 U14056 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11253) );
  AOI22_X1 U14057 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11252) );
  AOI22_X1 U14058 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11251) );
  AOI22_X1 U14059 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11250) );
  NAND4_X1 U14060 ( .A1(n11253), .A2(n11252), .A3(n11251), .A4(n11250), .ZN(
        n11254) );
  AOI211_X1 U14061 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n11255), .B(n11254), .ZN(n11256) );
  NAND2_X1 U14062 ( .A1(n11257), .A2(n11256), .ZN(n11451) );
  NAND2_X1 U14063 ( .A1(n11268), .A2(n11451), .ZN(n11291) );
  AOI22_X1 U14064 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11267) );
  AOI22_X1 U14065 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11266) );
  INV_X1 U14066 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17168) );
  INV_X2 U14067 ( .A(n17147), .ZN(n17124) );
  AOI22_X1 U14068 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11258) );
  OAI21_X1 U14069 ( .B1(n11326), .B2(n17168), .A(n11258), .ZN(n11264) );
  AOI22_X1 U14070 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11262) );
  AOI22_X1 U14071 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11261) );
  AOI22_X1 U14072 ( .A1(n17141), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11260) );
  AOI22_X1 U14073 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11259) );
  NAND4_X1 U14074 ( .A1(n11262), .A2(n11261), .A3(n11260), .A4(n11259), .ZN(
        n11263) );
  AOI211_X1 U14075 ( .C1(n17142), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n11264), .B(n11263), .ZN(n11265) );
  NAND3_X1 U14076 ( .A1(n11267), .A2(n11266), .A3(n11265), .ZN(n16354) );
  INV_X1 U14077 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17515) );
  INV_X1 U14078 ( .A(n11451), .ZN(n17329) );
  XNOR2_X1 U14079 ( .A(n11268), .B(n17329), .ZN(n11289) );
  INV_X1 U14080 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18102) );
  INV_X1 U14081 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18767) );
  NOR2_X1 U14082 ( .A1(n11283), .A2(n18767), .ZN(n11282) );
  INV_X1 U14083 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U14084 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11270) );
  OAI21_X1 U14085 ( .B1(n11326), .B2(n17146), .A(n11270), .ZN(n11278) );
  AOI22_X1 U14086 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11276) );
  AOI22_X1 U14087 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11327), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11275) );
  AOI22_X1 U14088 ( .A1(n11272), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11271), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11274) );
  AOI22_X1 U14089 ( .A1(n11227), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11245), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11273) );
  NAND4_X1 U14090 ( .A1(n11276), .A2(n11275), .A3(n11274), .A4(n11273), .ZN(
        n11277) );
  AOI22_X1 U14091 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14092 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11279) );
  XNOR2_X1 U14093 ( .A(n17349), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17820) );
  NOR2_X1 U14094 ( .A1(n11282), .A2(n17819), .ZN(n17809) );
  INV_X1 U14095 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18112) );
  XNOR2_X1 U14096 ( .A(n18112), .B(n11284), .ZN(n17808) );
  XNOR2_X1 U14097 ( .A(n11457), .B(n17332), .ZN(n11286) );
  NOR2_X1 U14098 ( .A1(n11287), .A2(n11286), .ZN(n11288) );
  NOR2_X2 U14099 ( .A1(n17796), .A2(n11288), .ZN(n17790) );
  XNOR2_X1 U14100 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11289), .ZN(
        n17789) );
  NOR2_X1 U14101 ( .A1(n17790), .A2(n17789), .ZN(n17788) );
  XNOR2_X1 U14102 ( .A(n11291), .B(n17325), .ZN(n11292) );
  INV_X1 U14103 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18084) );
  NOR2_X1 U14104 ( .A1(n11293), .A2(n11292), .ZN(n11294) );
  INV_X1 U14105 ( .A(n17761), .ZN(n17759) );
  INV_X1 U14106 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n17760) );
  XNOR2_X1 U14107 ( .A(n11296), .B(n17760), .ZN(n17766) );
  OAI21_X1 U14108 ( .B1(n11298), .B2(n16354), .A(n17702), .ZN(n11300) );
  INV_X1 U14109 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18071) );
  INV_X1 U14110 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17642) );
  INV_X1 U14111 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18041) );
  INV_X1 U14112 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17701) );
  NOR2_X1 U14113 ( .A1(n18041), .A2(n17701), .ZN(n18024) );
  NAND2_X1 U14114 ( .A1(n18024), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18010) );
  NOR2_X1 U14115 ( .A1(n18010), .A2(n18009), .ZN(n18006) );
  NAND2_X1 U14116 ( .A1(n18006), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17985) );
  INV_X1 U14117 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17987) );
  NOR2_X1 U14118 ( .A1(n17985), .A2(n17987), .ZN(n17968) );
  NAND2_X1 U14119 ( .A1(n17968), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16353) );
  NAND2_X1 U14120 ( .A1(n18041), .A2(n17701), .ZN(n17713) );
  NOR3_X1 U14121 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n17713), .ZN(n17638) );
  INV_X1 U14122 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11303) );
  INV_X1 U14123 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17960) );
  NOR2_X1 U14124 ( .A1(n17620), .A2(n11305), .ZN(n11306) );
  INV_X1 U14125 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17950) );
  NOR2_X1 U14126 ( .A1(n17960), .A2(n17950), .ZN(n17940) );
  INV_X1 U14127 ( .A(n17940), .ZN(n16352) );
  NAND2_X1 U14128 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17898) );
  INV_X1 U14129 ( .A(n17898), .ZN(n17916) );
  NAND3_X1 U14130 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17916), .ZN(n17900) );
  NOR2_X1 U14131 ( .A1(n16352), .A2(n17900), .ZN(n17895) );
  NAND3_X1 U14132 ( .A1(n17895), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17526) );
  INV_X1 U14133 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17929) );
  NAND2_X1 U14134 ( .A1(n17604), .A2(n17929), .ZN(n11308) );
  NOR2_X1 U14135 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11308), .ZN(
        n17566) );
  INV_X1 U14136 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17897) );
  NAND2_X1 U14137 ( .A1(n17566), .A2(n17897), .ZN(n17555) );
  INV_X1 U14138 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17524) );
  NAND2_X1 U14139 ( .A1(n17525), .A2(n17524), .ZN(n11313) );
  INV_X1 U14140 ( .A(n11313), .ZN(n11312) );
  NAND2_X1 U14141 ( .A1(n17940), .A2(n11311), .ZN(n17564) );
  INV_X1 U14142 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17543) );
  NOR2_X1 U14143 ( .A1(n17900), .A2(n17543), .ZN(n17884) );
  INV_X1 U14144 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17878) );
  INV_X1 U14145 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17851) );
  NOR2_X1 U14146 ( .A1(n17515), .A2(n17851), .ZN(n17841) );
  INV_X1 U14147 ( .A(n17841), .ZN(n11476) );
  NAND2_X1 U14148 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11314), .ZN(
        n17482) );
  OR2_X2 U14149 ( .A1(n11314), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17483) );
  NOR2_X2 U14150 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17483), .ZN(
        n11315) );
  OAI22_X1 U14151 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17702), .B1(
        n16362), .B2(n11315), .ZN(n15477) );
  INV_X1 U14152 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16342) );
  NAND2_X1 U14153 ( .A1(n15476), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15556) );
  NAND2_X1 U14154 ( .A1(n16342), .A2(n11315), .ZN(n11321) );
  INV_X1 U14155 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16336) );
  NOR2_X1 U14156 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16336), .ZN(
        n11316) );
  AOI21_X1 U14157 ( .B1(n11321), .B2(n17702), .A(n11316), .ZN(n11317) );
  INV_X1 U14158 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18768) );
  AOI21_X1 U14159 ( .B1(n17734), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n18768), .ZN(n11319) );
  AND2_X1 U14160 ( .A1(n17734), .A2(n18768), .ZN(n11318) );
  NOR2_X1 U14161 ( .A1(n11319), .A2(n11318), .ZN(n11324) );
  NAND2_X1 U14162 ( .A1(n11320), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11323) );
  NAND2_X1 U14163 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16336), .ZN(
        n11507) );
  OAI22_X1 U14164 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17702), .B1(
        n11507), .B2(n15555), .ZN(n11322) );
  AOI22_X1 U14166 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14167 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14168 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14169 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11328) );
  NAND4_X1 U14170 ( .A1(n11331), .A2(n11330), .A3(n11329), .A4(n11328), .ZN(
        n11337) );
  AOI22_X1 U14171 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11335) );
  AOI22_X1 U14172 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14173 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14174 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11332) );
  NAND4_X1 U14175 ( .A1(n11335), .A2(n11334), .A3(n11333), .A4(n11332), .ZN(
        n11336) );
  AOI22_X1 U14176 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14177 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14178 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11339) );
  AOI22_X1 U14179 ( .A1(n17077), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11338) );
  NAND4_X1 U14180 ( .A1(n11341), .A2(n11340), .A3(n11339), .A4(n11338), .ZN(
        n11347) );
  AOI22_X1 U14181 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11345) );
  AOI22_X1 U14182 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11344) );
  AOI22_X1 U14183 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11343) );
  AOI22_X1 U14184 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11342) );
  NAND4_X1 U14185 ( .A1(n11345), .A2(n11344), .A3(n11343), .A4(n11342), .ZN(
        n11346) );
  AOI22_X1 U14186 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14187 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11350) );
  AOI22_X1 U14188 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11349) );
  AOI22_X1 U14189 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11348) );
  NAND4_X1 U14190 ( .A1(n11351), .A2(n11350), .A3(n11349), .A4(n11348), .ZN(
        n11357) );
  AOI22_X1 U14191 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14192 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14193 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14194 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11352) );
  NAND4_X1 U14195 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n11356) );
  NOR2_X4 U14196 ( .A1(n11357), .A2(n11356), .ZN(n18808) );
  NAND2_X1 U14197 ( .A1(n11487), .A2(n18164), .ZN(n11438) );
  NOR2_X1 U14198 ( .A1(n17203), .A2(n11438), .ZN(n11445) );
  AOI22_X1 U14199 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11361) );
  AOI22_X1 U14200 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14201 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14202 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11358) );
  NAND4_X1 U14203 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n11367) );
  AOI22_X1 U14204 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11365) );
  AOI22_X1 U14205 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11364) );
  AOI22_X1 U14206 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11363) );
  AOI22_X1 U14207 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11362) );
  NAND4_X1 U14208 ( .A1(n11365), .A2(n11364), .A3(n11363), .A4(n11362), .ZN(
        n11366) );
  INV_X1 U14209 ( .A(n17203), .ZN(n18184) );
  NAND2_X1 U14210 ( .A1(n11411), .A2(n18184), .ZN(n11488) );
  AOI22_X1 U14211 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14212 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14213 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11368) );
  OAI21_X1 U14214 ( .B1(n11369), .B2(n17146), .A(n11368), .ZN(n11375) );
  AOI22_X1 U14215 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14216 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11372) );
  AOI22_X1 U14217 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11371) );
  AOI22_X1 U14218 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11370) );
  NAND4_X1 U14219 ( .A1(n11373), .A2(n11372), .A3(n11371), .A4(n11370), .ZN(
        n11374) );
  NAND2_X1 U14220 ( .A1(n15442), .A2(n18164), .ZN(n11426) );
  AOI22_X1 U14221 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14222 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14223 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17116), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14224 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11380) );
  NAND4_X1 U14225 ( .A1(n11383), .A2(n11382), .A3(n11381), .A4(n11380), .ZN(
        n11389) );
  AOI22_X1 U14226 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14227 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11386) );
  AOI22_X1 U14228 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11385) );
  AOI22_X1 U14229 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11384) );
  NAND4_X1 U14230 ( .A1(n11387), .A2(n11386), .A3(n11385), .A4(n11384), .ZN(
        n11388) );
  AOI22_X1 U14231 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17124), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17109), .ZN(n11393) );
  AOI22_X1 U14232 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14233 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17149), .ZN(n11391) );
  AOI22_X1 U14234 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17150), .ZN(n11390) );
  NAND4_X1 U14235 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11399) );
  AOI22_X1 U14236 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11397) );
  AOI22_X1 U14237 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17141), .B1(
        P3_INSTQUEUE_REG_8__7__SCAN_IN), .B2(n17050), .ZN(n11396) );
  AOI22_X1 U14238 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17024), .ZN(n11395) );
  AOI22_X1 U14239 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17132), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11394) );
  NAND4_X1 U14240 ( .A1(n11397), .A2(n11396), .A3(n11395), .A4(n11394), .ZN(
        n11398) );
  AOI22_X1 U14241 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11403) );
  AOI22_X1 U14242 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14243 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14244 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11400) );
  NAND4_X1 U14245 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n11409) );
  AOI22_X1 U14246 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14247 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14248 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14249 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11404) );
  NAND4_X1 U14250 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11408) );
  NOR2_X1 U14251 ( .A1(n16989), .A2(n18171), .ZN(n11496) );
  OAI21_X1 U14252 ( .B1(n15439), .B2(n18616), .A(n11490), .ZN(n11495) );
  INV_X1 U14253 ( .A(n11495), .ZN(n11410) );
  NOR2_X1 U14254 ( .A1(n17203), .A2(n11411), .ZN(n11430) );
  AOI21_X1 U14255 ( .B1(n11487), .B2(n11430), .A(n18176), .ZN(n11441) );
  INV_X1 U14256 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18639) );
  OAI22_X1 U14257 ( .A1(n18782), .A2(n18623), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14258 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18628), .B2(n11412), .ZN(
        n11422) );
  OAI22_X1 U14259 ( .A1(n18632), .A2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(
        n11415), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11420) );
  NAND2_X1 U14260 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11415), .ZN(
        n11418) );
  AND2_X1 U14261 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11418), .ZN(
        n11416) );
  OAI22_X1 U14262 ( .A1(n18639), .A2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(
        n11420), .B2(n11416), .ZN(n11417) );
  INV_X1 U14263 ( .A(n11417), .ZN(n11436) );
  NOR2_X1 U14264 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18632), .ZN(
        n11419) );
  AOI22_X1 U14265 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11420), .B1(
        n11419), .B2(n11418), .ZN(n11424) );
  NAND2_X1 U14266 ( .A1(n11423), .A2(n11422), .ZN(n11421) );
  OAI211_X1 U14267 ( .C1(n11423), .C2(n11422), .A(n11424), .B(n11421), .ZN(
        n11444) );
  AOI21_X1 U14268 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n18789), .A(
        n11435), .ZN(n11442) );
  NAND3_X1 U14269 ( .A1(n11434), .A2(n11424), .A3(n11442), .ZN(n11425) );
  NAND3_X1 U14270 ( .A1(n11436), .A2(n11444), .A3(n11425), .ZN(n18582) );
  AOI211_X1 U14271 ( .C1(n18188), .C2(n15584), .A(n15442), .B(n18164), .ZN(
        n11481) );
  AOI21_X1 U14272 ( .B1(n11487), .B2(n11426), .A(n11430), .ZN(n11429) );
  NAND2_X1 U14273 ( .A1(n17203), .A2(n18176), .ZN(n18594) );
  AOI21_X1 U14274 ( .B1(n18594), .B2(n18180), .A(n16989), .ZN(n11427) );
  NAND3_X1 U14275 ( .A1(n11487), .A2(n18594), .A3(n11488), .ZN(n11483) );
  OAI22_X1 U14276 ( .A1(n11489), .A2(n11427), .B1(n18157), .B2(n11483), .ZN(
        n11428) );
  AOI211_X1 U14277 ( .C1(n18171), .C2(n11494), .A(n11429), .B(n11428), .ZN(
        n11484) );
  NAND4_X1 U14278 ( .A1(n15439), .A2(n18171), .A3(n11431), .A4(n11430), .ZN(
        n11486) );
  NOR2_X1 U14279 ( .A1(n11487), .A2(n11486), .ZN(n11491) );
  AOI21_X1 U14280 ( .B1(n11432), .B2(n11484), .A(n11491), .ZN(n11433) );
  NOR2_X1 U14281 ( .A1(n11481), .A2(n11433), .ZN(n13844) );
  XNOR2_X1 U14282 ( .A(n11435), .B(n11434), .ZN(n11437) );
  INV_X1 U14283 ( .A(n11487), .ZN(n18167) );
  NAND2_X2 U14284 ( .A1(n18733), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18743) );
  INV_X1 U14285 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18671) );
  INV_X1 U14286 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18679) );
  NAND2_X1 U14287 ( .A1(n18671), .A2(n18679), .ZN(n18661) );
  NAND3_X1 U14288 ( .A1(n18677), .A2(n18743), .A3(n18661), .ZN(n18806) );
  INV_X1 U14289 ( .A(n18806), .ZN(n13840) );
  AOI21_X1 U14290 ( .B1(n18808), .B2(n18167), .A(n13840), .ZN(n11439) );
  NAND2_X1 U14291 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18809) );
  INV_X1 U14292 ( .A(n18809), .ZN(n18669) );
  AOI21_X1 U14293 ( .B1(n11439), .B2(n11438), .A(n18669), .ZN(n16472) );
  NAND2_X1 U14294 ( .A1(n11487), .A2(n18180), .ZN(n11482) );
  NAND3_X1 U14295 ( .A1(n18586), .A2(n16472), .A3(n11482), .ZN(n11440) );
  OAI211_X1 U14296 ( .C1(n11441), .C2(n18582), .A(n13844), .B(n11440), .ZN(
        n11446) );
  INV_X1 U14297 ( .A(n11442), .ZN(n11443) );
  OAI21_X1 U14298 ( .B1(n11444), .B2(n11443), .A(n18586), .ZN(n12833) );
  INV_X1 U14299 ( .A(n12833), .ZN(n18587) );
  NAND2_X1 U14300 ( .A1(n11302), .A2(n17702), .ZN(n17639) );
  INV_X1 U14301 ( .A(n17526), .ZN(n11447) );
  NAND2_X1 U14302 ( .A1(n17891), .A2(n11447), .ZN(n17874) );
  NAND2_X1 U14303 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11500) );
  INV_X1 U14304 ( .A(n11500), .ZN(n11477) );
  NAND2_X1 U14305 ( .A1(n17843), .A2(n11477), .ZN(n16343) );
  NOR3_X1 U14306 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16342), .A3(
        n16336), .ZN(n11509) );
  NAND2_X1 U14307 ( .A1(n11477), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16328) );
  INV_X1 U14308 ( .A(n16328), .ZN(n11478) );
  NAND2_X1 U14309 ( .A1(n17843), .A2(n11478), .ZN(n16327) );
  OR2_X1 U14310 ( .A1(n16336), .A2(n16327), .ZN(n11448) );
  AOI22_X1 U14311 ( .A1(n16367), .A2(n11509), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n11448), .ZN(n12835) );
  NAND2_X1 U14312 ( .A1(n17319), .A2(n18136), .ZN(n18064) );
  OR2_X1 U14313 ( .A1(n12835), .A2(n18064), .ZN(n11513) );
  NAND2_X1 U14314 ( .A1(n11283), .A2(n15585), .ZN(n11458) );
  INV_X1 U14315 ( .A(n11449), .ZN(n17338) );
  NAND2_X1 U14316 ( .A1(n11458), .A2(n17338), .ZN(n11455) );
  INV_X1 U14317 ( .A(n11455), .ZN(n11450) );
  NOR2_X1 U14318 ( .A1(n17332), .A2(n11450), .ZN(n11454) );
  NAND2_X1 U14319 ( .A1(n11454), .A2(n11451), .ZN(n11453) );
  NAND2_X1 U14320 ( .A1(n17758), .A2(n17759), .ZN(n11452) );
  NOR2_X1 U14321 ( .A1(n17319), .A2(n11452), .ZN(n11474) );
  XOR2_X1 U14322 ( .A(n17319), .B(n11452), .Z(n11470) );
  XOR2_X1 U14323 ( .A(n17325), .B(n11453), .Z(n11466) );
  AND2_X1 U14324 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11466), .ZN(
        n11467) );
  XNOR2_X1 U14325 ( .A(n17329), .B(n11454), .ZN(n11464) );
  AND2_X1 U14326 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11464), .ZN(
        n11465) );
  XNOR2_X1 U14327 ( .A(n17332), .B(n11455), .ZN(n11462) );
  AND2_X1 U14328 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11462), .ZN(
        n11463) );
  INV_X1 U14329 ( .A(n15585), .ZN(n11456) );
  OAI21_X1 U14330 ( .B1(n11457), .B2(n11456), .A(n11455), .ZN(n11459) );
  AND2_X1 U14331 ( .A1(n11459), .A2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11461) );
  NOR2_X1 U14332 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15585), .ZN(
        n17827) );
  NAND2_X1 U14333 ( .A1(n17827), .A2(n17820), .ZN(n17817) );
  OAI211_X1 U14334 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n11283), .A(
        n11458), .B(n17817), .ZN(n17811) );
  XNOR2_X1 U14335 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11459), .ZN(
        n17810) );
  NOR2_X1 U14336 ( .A1(n17811), .A2(n17810), .ZN(n11460) );
  NOR2_X1 U14337 ( .A1(n11461), .A2(n11460), .ZN(n17799) );
  XNOR2_X1 U14338 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11462), .ZN(
        n17798) );
  NOR2_X1 U14339 ( .A1(n17799), .A2(n17798), .ZN(n17797) );
  NOR2_X1 U14340 ( .A1(n11463), .A2(n17797), .ZN(n17785) );
  XNOR2_X1 U14341 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11464), .ZN(
        n17784) );
  NOR2_X1 U14342 ( .A1(n17785), .A2(n17784), .ZN(n17783) );
  NOR2_X1 U14343 ( .A1(n11465), .A2(n17783), .ZN(n17775) );
  XNOR2_X1 U14344 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11466), .ZN(
        n17774) );
  NOR2_X1 U14345 ( .A1(n17775), .A2(n17774), .ZN(n17773) );
  NOR2_X1 U14346 ( .A1(n11467), .A2(n17773), .ZN(n17757) );
  XOR2_X1 U14347 ( .A(n17761), .B(n17758), .Z(n11468) );
  AOI222_X1 U14348 ( .A1(n17757), .A2(n17760), .B1(n17757), .B2(n11468), .C1(
        n17760), .C2(n11468), .ZN(n11471) );
  NOR2_X1 U14349 ( .A1(n11470), .A2(n11471), .ZN(n17750) );
  NOR2_X1 U14350 ( .A1(n17750), .A2(n18071), .ZN(n11469) );
  NAND2_X1 U14351 ( .A1(n11474), .A2(n11469), .ZN(n11475) );
  INV_X1 U14352 ( .A(n11469), .ZN(n11473) );
  AND2_X1 U14353 ( .A1(n11471), .A2(n11470), .ZN(n17751) );
  AOI21_X1 U14354 ( .B1(n11474), .B2(n11473), .A(n17751), .ZN(n11472) );
  OAI21_X1 U14355 ( .B1(n11474), .B2(n11473), .A(n11472), .ZN(n17736) );
  NAND2_X1 U14356 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17736), .ZN(
        n17735) );
  NAND2_X1 U14357 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17527), .ZN(
        n17505) );
  NAND2_X1 U14358 ( .A1(n11477), .A2(n17842), .ZN(n16364) );
  INV_X1 U14359 ( .A(n11509), .ZN(n11480) );
  NAND2_X1 U14360 ( .A1(n11478), .A2(n17842), .ZN(n16326) );
  OAI21_X1 U14361 ( .B1(n16336), .B2(n16326), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11479) );
  OAI21_X1 U14362 ( .B1(n16364), .B2(n11480), .A(n11479), .ZN(n12840) );
  AOI21_X1 U14363 ( .B1(n11483), .B2(n11482), .A(n11481), .ZN(n11485) );
  OAI21_X1 U14364 ( .B1(n18171), .B2(n11485), .A(n11484), .ZN(n11497) );
  NOR2_X2 U14365 ( .A1(n11486), .A2(n11497), .ZN(n13837) );
  NAND2_X1 U14366 ( .A1(n18171), .A2(n11487), .ZN(n18593) );
  NOR2_X1 U14367 ( .A1(n11488), .A2(n18593), .ZN(n15438) );
  NAND2_X1 U14368 ( .A1(n18808), .A2(n15438), .ZN(n11493) );
  NAND4_X1 U14369 ( .A1(n18157), .A2(n17203), .A3(n11490), .A4(n11489), .ZN(
        n11492) );
  INV_X1 U14370 ( .A(n11492), .ZN(n17416) );
  NOR2_X1 U14371 ( .A1(n18808), .A2(n11496), .ZN(n11499) );
  AOI21_X1 U14372 ( .B1(n11499), .B2(n11498), .A(n11497), .ZN(n18592) );
  NOR2_X1 U14373 ( .A1(n18017), .A2(n18127), .ZN(n18126) );
  AOI21_X1 U14374 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18050) );
  NAND2_X1 U14375 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18077) );
  NOR3_X1 U14376 ( .A1(n17760), .A2(n18102), .A3(n18077), .ZN(n18068) );
  NAND3_X1 U14377 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18068), .ZN(n16355) );
  OR2_X1 U14378 ( .A1(n18050), .A2(n16355), .ZN(n17957) );
  NOR3_X1 U14379 ( .A1(n16353), .A2(n16352), .A3(n17957), .ZN(n17892) );
  AND2_X1 U14380 ( .A1(n18613), .A2(n17892), .ZN(n16356) );
  INV_X1 U14381 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18786) );
  OAI21_X1 U14382 ( .B1(n18605), .B2(n18786), .A(n18617), .ZN(n18113) );
  NOR2_X1 U14383 ( .A1(n18112), .A2(n18767), .ZN(n18114) );
  INV_X1 U14384 ( .A(n16355), .ZN(n17937) );
  NAND2_X1 U14385 ( .A1(n18114), .A2(n17937), .ZN(n17956) );
  NOR2_X1 U14386 ( .A1(n16353), .A2(n17956), .ZN(n17939) );
  NAND2_X1 U14387 ( .A1(n17895), .A2(n17939), .ZN(n17840) );
  NOR2_X1 U14388 ( .A1(n17543), .A2(n17840), .ZN(n11501) );
  AOI22_X1 U14389 ( .A1(n17884), .A2(n16356), .B1(n18113), .B2(n11501), .ZN(
        n17858) );
  NOR2_X1 U14390 ( .A1(n17878), .A2(n17524), .ZN(n17860) );
  NAND2_X1 U14391 ( .A1(n17841), .A2(n17860), .ZN(n11503) );
  NOR4_X1 U14392 ( .A1(n17858), .A2(n18127), .A3(n11500), .A4(n11503), .ZN(
        n15472) );
  INV_X1 U14393 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18740) );
  NAND2_X1 U14394 ( .A1(n18813), .A2(n18758), .ZN(n18771) );
  NOR2_X1 U14395 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18771), .ZN(n18821) );
  NOR2_X1 U14396 ( .A1(n18740), .A2(n18036), .ZN(n12839) );
  NOR2_X1 U14397 ( .A1(n18053), .A2(n18127), .ZN(n18130) );
  NAND2_X1 U14398 ( .A1(n18036), .A2(n18127), .ZN(n17986) );
  NAND2_X1 U14399 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n11501), .ZN(
        n17838) );
  INV_X1 U14400 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17836) );
  OR2_X1 U14401 ( .A1(n17836), .A2(n11503), .ZN(n16359) );
  OAI21_X1 U14402 ( .B1(n17838), .B2(n16359), .A(n18615), .ZN(n11506) );
  INV_X1 U14403 ( .A(n11501), .ZN(n11502) );
  INV_X1 U14404 ( .A(n18617), .ZN(n18131) );
  OAI21_X1 U14405 ( .B1(n11502), .B2(n11503), .A(n18131), .ZN(n11505) );
  NAND2_X1 U14406 ( .A1(n17884), .A2(n17892), .ZN(n17837) );
  OAI21_X1 U14407 ( .B1(n11503), .B2(n17837), .A(n18613), .ZN(n11504) );
  NAND4_X1 U14408 ( .A1(n17986), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n15473) );
  AOI22_X1 U14409 ( .A1(n18130), .A2(n16328), .B1(n18036), .B2(n15473), .ZN(
        n15562) );
  INV_X1 U14410 ( .A(n18130), .ZN(n18078) );
  OAI22_X1 U14411 ( .A1(n15562), .A2(n18768), .B1(n11507), .B2(n18078), .ZN(
        n11508) );
  AOI211_X1 U14412 ( .C1(n11509), .C2(n15472), .A(n12839), .B(n11508), .ZN(
        n11510) );
  AOI21_X1 U14413 ( .B1(n12840), .B2(n18126), .A(n11511), .ZN(n11512) );
  AND2_X1 U14414 ( .A1(n11513), .A2(n11512), .ZN(n11514) );
  NAND2_X1 U14415 ( .A1(n11515), .A2(n11514), .ZN(P3_U2831) );
  NAND2_X1 U14416 ( .A1(n11529), .A2(n11528), .ZN(n11516) );
  NAND2_X1 U14417 ( .A1(n11516), .A2(n11517), .ZN(n11544) );
  OAI21_X1 U14418 ( .B1(n11517), .B2(n11516), .A(n11544), .ZN(n11521) );
  NAND2_X1 U14419 ( .A1(n20149), .A2(n11518), .ZN(n11524) );
  INV_X1 U14420 ( .A(n11524), .ZN(n11520) );
  AOI21_X1 U14421 ( .B1(n11521), .B2(n15538), .A(n11520), .ZN(n11522) );
  NAND2_X1 U14422 ( .A1(n11523), .A2(n11522), .ZN(n13303) );
  OAI21_X1 U14423 ( .B1(n10240), .B2(n11528), .A(n11524), .ZN(n11525) );
  INV_X1 U14424 ( .A(n11525), .ZN(n11526) );
  OAI21_X2 U14425 ( .B1(n11527), .B2(n11585), .A(n11526), .ZN(n13102) );
  NAND2_X2 U14426 ( .A1(n13102), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13103) );
  XNOR2_X1 U14427 ( .A(n11529), .B(n11528), .ZN(n11532) );
  OAI211_X1 U14428 ( .C1(n11532), .C2(n10240), .A(n11530), .B(n11531), .ZN(
        n11533) );
  INV_X1 U14429 ( .A(n11533), .ZN(n11534) );
  NAND2_X1 U14430 ( .A1(n13228), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11539) );
  INV_X1 U14431 ( .A(n11536), .ZN(n11537) );
  INV_X1 U14432 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11540) );
  NAND2_X1 U14433 ( .A1(n13303), .A2(n13304), .ZN(n11543) );
  NAND2_X1 U14434 ( .A1(n11541), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11542) );
  INV_X1 U14435 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13384) );
  NAND2_X1 U14436 ( .A1(n11544), .A2(n11545), .ZN(n11559) );
  OAI211_X1 U14437 ( .C1(n11545), .C2(n11544), .A(n11559), .B(n15538), .ZN(
        n11546) );
  NAND2_X1 U14438 ( .A1(n11548), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11549) );
  INV_X1 U14439 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11550) );
  INV_X1 U14440 ( .A(n11551), .ZN(n11558) );
  XNOR2_X1 U14441 ( .A(n11559), .B(n11558), .ZN(n11552) );
  OAI22_X1 U14442 ( .A1(n11553), .A2(n11585), .B1(n11552), .B2(n10240), .ZN(
        n13535) );
  NAND2_X1 U14443 ( .A1(n11554), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11555) );
  NAND2_X1 U14444 ( .A1(n11556), .A2(n11555), .ZN(n13616) );
  OR2_X1 U14445 ( .A1(n11557), .A2(n11585), .ZN(n11563) );
  NOR2_X1 U14446 ( .A1(n11559), .A2(n11558), .ZN(n11561) );
  NAND2_X1 U14447 ( .A1(n11561), .A2(n11560), .ZN(n11575) );
  OAI211_X1 U14448 ( .C1(n11561), .C2(n11560), .A(n11575), .B(n15538), .ZN(
        n11562) );
  NAND2_X1 U14449 ( .A1(n11563), .A2(n11562), .ZN(n11564) );
  INV_X1 U14450 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11770) );
  XNOR2_X1 U14451 ( .A(n11564), .B(n11770), .ZN(n13617) );
  NAND2_X1 U14452 ( .A1(n13616), .A2(n13617), .ZN(n11566) );
  NAND2_X1 U14453 ( .A1(n11564), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11565) );
  NAND2_X1 U14454 ( .A1(n11566), .A2(n11565), .ZN(n15776) );
  INV_X1 U14455 ( .A(n11585), .ZN(n11627) );
  NAND3_X1 U14456 ( .A1(n11567), .A2(n11568), .A3(n11627), .ZN(n11571) );
  XNOR2_X1 U14457 ( .A(n11575), .B(n11576), .ZN(n11569) );
  NAND2_X1 U14458 ( .A1(n11569), .A2(n15538), .ZN(n11570) );
  NAND2_X1 U14459 ( .A1(n11571), .A2(n11570), .ZN(n11572) );
  OR2_X1 U14460 ( .A1(n11572), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15778) );
  NAND2_X1 U14461 ( .A1(n15776), .A2(n15778), .ZN(n11573) );
  NAND2_X1 U14462 ( .A1(n11572), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15777) );
  NAND2_X1 U14463 ( .A1(n11573), .A2(n15777), .ZN(n13731) );
  INV_X1 U14464 ( .A(n13731), .ZN(n11582) );
  NAND2_X1 U14465 ( .A1(n11574), .A2(n11627), .ZN(n11580) );
  INV_X1 U14466 ( .A(n11575), .ZN(n11577) );
  NAND2_X1 U14467 ( .A1(n11577), .A2(n11576), .ZN(n11590) );
  XNOR2_X1 U14468 ( .A(n11590), .B(n11588), .ZN(n11578) );
  NAND2_X1 U14469 ( .A1(n11578), .A2(n15538), .ZN(n11579) );
  NAND2_X1 U14470 ( .A1(n11580), .A2(n11579), .ZN(n11583) );
  XNOR2_X1 U14471 ( .A(n11583), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13732) );
  INV_X1 U14472 ( .A(n13732), .ZN(n11581) );
  OR2_X1 U14473 ( .A1(n11583), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11584) );
  NOR2_X1 U14474 ( .A1(n11586), .A2(n11585), .ZN(n11587) );
  NAND2_X1 U14475 ( .A1(n15538), .A2(n11588), .ZN(n11589) );
  OR2_X1 U14476 ( .A1(n11590), .A2(n11589), .ZN(n11591) );
  NAND2_X1 U14477 ( .A1(n13758), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11592) );
  INV_X1 U14478 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15907) );
  NAND2_X1 U14479 ( .A1(n9820), .A2(n15907), .ZN(n11594) );
  INV_X1 U14480 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15878) );
  OR2_X1 U14481 ( .A1(n9820), .A2(n15878), .ZN(n15742) );
  NAND2_X1 U14482 ( .A1(n9820), .A2(n15878), .ZN(n11595) );
  NAND2_X1 U14483 ( .A1(n15742), .A2(n11595), .ZN(n14628) );
  INV_X1 U14484 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n14627) );
  NAND2_X1 U14485 ( .A1(n9820), .A2(n14627), .ZN(n15754) );
  NAND2_X1 U14486 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11596) );
  NAND2_X1 U14487 ( .A1(n9820), .A2(n11596), .ZN(n14626) );
  NAND2_X1 U14488 ( .A1(n15754), .A2(n14626), .ZN(n11597) );
  NOR2_X1 U14489 ( .A1(n14628), .A2(n11597), .ZN(n15744) );
  INV_X1 U14490 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15863) );
  NAND2_X1 U14491 ( .A1(n9820), .A2(n15863), .ZN(n11598) );
  XNOR2_X1 U14492 ( .A(n9820), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15737) );
  INV_X1 U14493 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15844) );
  NAND2_X1 U14494 ( .A1(n9820), .A2(n15844), .ZN(n14613) );
  NAND2_X1 U14495 ( .A1(n15737), .A2(n14613), .ZN(n14601) );
  NOR2_X1 U14496 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11599) );
  OAI22_X1 U14497 ( .A1(n15735), .A2(n14601), .B1(n11599), .B2(n9820), .ZN(
        n11601) );
  INV_X1 U14498 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14605) );
  NAND2_X1 U14499 ( .A1(n9820), .A2(n14605), .ZN(n11600) );
  INV_X1 U14500 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U14501 ( .A1(n15768), .A2(n15763), .ZN(n14598) );
  NAND3_X1 U14502 ( .A1(n15863), .A2(n15878), .A3(n14627), .ZN(n11602) );
  NOR2_X1 U14503 ( .A1(n14598), .A2(n11602), .ZN(n11603) );
  NAND2_X1 U14504 ( .A1(n9820), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14505 ( .A1(n14586), .A2(n11605), .ZN(n14593) );
  AND2_X1 U14506 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11773) );
  NAND2_X1 U14507 ( .A1(n11773), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15805) );
  INV_X1 U14508 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14708) );
  INV_X1 U14509 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15572) );
  NAND2_X1 U14510 ( .A1(n14708), .A2(n15572), .ZN(n15569) );
  INV_X1 U14511 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14581) );
  INV_X1 U14512 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15835) );
  NAND2_X1 U14513 ( .A1(n11612), .A2(n15720), .ZN(n11610) );
  INV_X1 U14514 ( .A(n11610), .ZN(n14562) );
  INV_X1 U14515 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14552) );
  INV_X1 U14516 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14689) );
  NAND2_X1 U14517 ( .A1(n14552), .A2(n14689), .ZN(n14518) );
  INV_X1 U14518 ( .A(n14518), .ZN(n11607) );
  NAND2_X1 U14519 ( .A1(n11609), .A2(n14587), .ZN(n14539) );
  NAND2_X1 U14520 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14687) );
  INV_X1 U14521 ( .A(n14687), .ZN(n11611) );
  NAND2_X1 U14522 ( .A1(n11611), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15796) );
  NAND2_X1 U14523 ( .A1(n14572), .A2(n15796), .ZN(n11613) );
  NAND2_X1 U14524 ( .A1(n11612), .A2(n9820), .ZN(n14548) );
  NAND3_X1 U14525 ( .A1(n11613), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14548), .ZN(n14529) );
  NAND2_X1 U14526 ( .A1(n14539), .A2(n14529), .ZN(n14530) );
  NAND2_X1 U14527 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14666) );
  NAND2_X1 U14528 ( .A1(n9820), .A2(n14666), .ZN(n11616) );
  INV_X1 U14529 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14675) );
  INV_X1 U14530 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14660) );
  NAND2_X1 U14531 ( .A1(n14675), .A2(n14660), .ZN(n14665) );
  INV_X1 U14532 ( .A(n14665), .ZN(n11614) );
  INV_X1 U14533 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11780) );
  INV_X1 U14534 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11617) );
  NAND2_X1 U14535 ( .A1(n14508), .A2(n11617), .ZN(n11620) );
  NOR2_X1 U14536 ( .A1(n14666), .A2(n11780), .ZN(n11775) );
  AND2_X1 U14537 ( .A1(n9820), .A2(n11775), .ZN(n11618) );
  NAND2_X1 U14538 ( .A1(n14530), .A2(n11618), .ZN(n14507) );
  NAND2_X1 U14539 ( .A1(n11620), .A2(n11619), .ZN(n11621) );
  XNOR2_X1 U14540 ( .A(n11621), .B(n14729), .ZN(n13983) );
  AND2_X1 U14541 ( .A1(n11114), .A2(n13608), .ZN(n13281) );
  NAND4_X1 U14542 ( .A1(n11530), .A2(n11641), .A3(n13281), .A4(n10416), .ZN(
        n13141) );
  OAI21_X1 U14543 ( .B1(n13141), .B2(n15563), .A(n13443), .ZN(n11625) );
  INV_X1 U14544 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n11622) );
  NAND2_X1 U14545 ( .A1(n11623), .A2(n11622), .ZN(n15564) );
  NAND2_X1 U14546 ( .A1(n15538), .A2(n15564), .ZN(n11624) );
  AOI21_X1 U14547 ( .B1(n11625), .B2(n11624), .A(n13282), .ZN(n11626) );
  OR2_X1 U14548 ( .A1(n11626), .A2(n10394), .ZN(n11636) );
  NOR2_X1 U14549 ( .A1(n10401), .A2(n20156), .ZN(n11748) );
  NAND2_X1 U14550 ( .A1(n13155), .A2(n11748), .ZN(n11635) );
  AOI21_X1 U14551 ( .B1(n11627), .B2(n10416), .A(n20149), .ZN(n11628) );
  NAND2_X1 U14552 ( .A1(n10412), .A2(n11628), .ZN(n11755) );
  NAND3_X1 U14553 ( .A1(n11755), .A2(n11749), .A3(n11639), .ZN(n11630) );
  NAND2_X1 U14554 ( .A1(n11630), .A2(n10168), .ZN(n13144) );
  NAND2_X1 U14555 ( .A1(n13447), .A2(n15564), .ZN(n11631) );
  NAND3_X1 U14556 ( .A1(n11631), .A2(n10394), .A3(n20800), .ZN(n11632) );
  OR2_X1 U14557 ( .A1(n12964), .A2(n11632), .ZN(n11633) );
  AND2_X1 U14558 ( .A1(n13144), .A2(n11633), .ZN(n11634) );
  OAI211_X1 U14559 ( .C1(n13155), .C2(n11636), .A(n11635), .B(n11634), .ZN(
        n11637) );
  NAND3_X1 U14560 ( .A1(n11639), .A2(n11638), .A3(n11749), .ZN(n11782) );
  NAND2_X1 U14561 ( .A1(n11782), .A2(n13313), .ZN(n12963) );
  OAI21_X1 U14562 ( .B1(n11640), .B2(n11641), .A(n11097), .ZN(n11642) );
  NOR2_X1 U14563 ( .A1(n12963), .A2(n11642), .ZN(n11643) );
  NAND2_X1 U14564 ( .A1(n11643), .A2(n11154), .ZN(n11644) );
  OAI22_X1 U14565 ( .A1(n11640), .A2(n13596), .B1(n12962), .B2(n13447), .ZN(
        n11645) );
  AOI22_X1 U14566 ( .A1(n13106), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13129), .ZN(n11744) );
  AOI22_X1 U14567 ( .A1(n13106), .A2(P1_EBX_REG_30__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n13129), .ZN(n14296) );
  INV_X1 U14568 ( .A(n11692), .ZN(n11681) );
  OR2_X1 U14569 ( .A1(n13106), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11646) );
  INV_X1 U14570 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11648) );
  OAI22_X1 U14571 ( .A1(n11737), .A2(n11648), .B1(n11681), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13107) );
  XNOR2_X1 U14572 ( .A(n11649), .B(n13107), .ZN(n13515) );
  AOI21_X1 U14573 ( .B1(n13515), .B2(n13217), .A(n11649), .ZN(n13272) );
  INV_X1 U14574 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n21030) );
  NAND2_X1 U14575 ( .A1(n11735), .A2(n21030), .ZN(n11652) );
  NAND2_X1 U14576 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11650) );
  OAI211_X1 U14577 ( .C1(n13129), .C2(P1_EBX_REG_2__SCAN_IN), .A(n11737), .B(
        n11650), .ZN(n11651) );
  NAND2_X1 U14578 ( .A1(n13272), .A2(n13271), .ZN(n13365) );
  INV_X1 U14579 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n21172) );
  NAND2_X1 U14580 ( .A1(n11717), .A2(n21172), .ZN(n11656) );
  NAND2_X1 U14581 ( .A1(n11737), .A2(n13384), .ZN(n11654) );
  NAND2_X1 U14582 ( .A1(n13217), .A2(n21172), .ZN(n11653) );
  NAND3_X1 U14583 ( .A1(n11654), .A2(n11681), .A3(n11653), .ZN(n11655) );
  NAND2_X1 U14584 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11657) );
  OAI211_X1 U14585 ( .C1(n13129), .C2(P1_EBX_REG_4__SCAN_IN), .A(n11737), .B(
        n11657), .ZN(n11658) );
  OAI21_X1 U14586 ( .B1(n11732), .B2(P1_EBX_REG_4__SCAN_IN), .A(n11658), .ZN(
        n13462) );
  MUX2_X1 U14587 ( .A(n11742), .B(n11737), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n11663) );
  INV_X1 U14588 ( .A(n11659), .ZN(n11660) );
  NAND2_X1 U14589 ( .A1(n11660), .A2(n13129), .ZN(n11710) );
  NAND2_X1 U14590 ( .A1(n13129), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11661) );
  AND2_X1 U14591 ( .A1(n11710), .A2(n11661), .ZN(n11662) );
  NAND2_X1 U14592 ( .A1(n11663), .A2(n11662), .ZN(n13579) );
  INV_X1 U14593 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20077) );
  NAND2_X1 U14594 ( .A1(n11735), .A2(n20077), .ZN(n11666) );
  NAND2_X1 U14595 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11664) );
  OAI211_X1 U14596 ( .C1(n13129), .C2(P1_EBX_REG_6__SCAN_IN), .A(n11737), .B(
        n11664), .ZN(n11665) );
  MUX2_X1 U14597 ( .A(n11742), .B(n11737), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n11668) );
  NAND2_X1 U14598 ( .A1(n13129), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11667) );
  NAND2_X1 U14599 ( .A1(n11669), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11670) );
  OAI211_X1 U14600 ( .C1(n13129), .C2(P1_EBX_REG_8__SCAN_IN), .A(n11737), .B(
        n11670), .ZN(n11671) );
  OAI21_X1 U14601 ( .B1(n11732), .B2(P1_EBX_REG_8__SCAN_IN), .A(n11671), .ZN(
        n13586) );
  MUX2_X1 U14602 ( .A(n11742), .B(n11737), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n11674) );
  NAND2_X1 U14603 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n13129), .ZN(
        n11672) );
  AND2_X1 U14604 ( .A1(n11710), .A2(n11672), .ZN(n11673) );
  NAND2_X1 U14605 ( .A1(n11674), .A2(n11673), .ZN(n13640) );
  MUX2_X1 U14606 ( .A(n11732), .B(n11681), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11676) );
  OR2_X1 U14607 ( .A1(n13106), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11675) );
  INV_X1 U14608 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15719) );
  NAND2_X1 U14609 ( .A1(n11717), .A2(n15719), .ZN(n11680) );
  NAND2_X1 U14610 ( .A1(n11737), .A2(n15768), .ZN(n11678) );
  NAND2_X1 U14611 ( .A1(n13217), .A2(n15719), .ZN(n11677) );
  NAND3_X1 U14612 ( .A1(n11678), .A2(n11681), .A3(n11677), .ZN(n11679) );
  NAND2_X1 U14613 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11682) );
  OAI211_X1 U14614 ( .C1(n13129), .C2(P1_EBX_REG_12__SCAN_IN), .A(n11737), .B(
        n11682), .ZN(n11683) );
  OAI21_X1 U14615 ( .B1(n11732), .B2(P1_EBX_REG_12__SCAN_IN), .A(n11683), .ZN(
        n15685) );
  INV_X1 U14616 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n11684) );
  NAND2_X1 U14617 ( .A1(n11717), .A2(n11684), .ZN(n11688) );
  NAND2_X1 U14618 ( .A1(n11737), .A2(n15878), .ZN(n11686) );
  NAND2_X1 U14619 ( .A1(n13217), .A2(n11684), .ZN(n11685) );
  NAND3_X1 U14620 ( .A1(n11686), .A2(n11681), .A3(n11685), .ZN(n11687) );
  MUX2_X1 U14621 ( .A(n11732), .B(n11681), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11691) );
  INV_X1 U14622 ( .A(n13106), .ZN(n11689) );
  NAND2_X1 U14623 ( .A1(n15863), .A2(n11689), .ZN(n11690) );
  INV_X1 U14624 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n21134) );
  NAND2_X1 U14625 ( .A1(n11735), .A2(n21134), .ZN(n11695) );
  NAND2_X1 U14626 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11693) );
  OAI211_X1 U14627 ( .C1(n13129), .C2(P1_EBX_REG_16__SCAN_IN), .A(n11737), .B(
        n11693), .ZN(n11694) );
  AND2_X1 U14628 ( .A1(n11695), .A2(n11694), .ZN(n15665) );
  INV_X1 U14629 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n21009) );
  NAND2_X1 U14630 ( .A1(n11717), .A2(n21009), .ZN(n11699) );
  NAND2_X1 U14631 ( .A1(n11737), .A2(n15844), .ZN(n11697) );
  NAND2_X1 U14632 ( .A1(n13217), .A2(n21009), .ZN(n11696) );
  NAND3_X1 U14633 ( .A1(n11697), .A2(n11681), .A3(n11696), .ZN(n11698) );
  NAND2_X1 U14634 ( .A1(n11699), .A2(n11698), .ZN(n13801) );
  NAND2_X1 U14635 ( .A1(n15665), .A2(n13801), .ZN(n11700) );
  MUX2_X1 U14636 ( .A(n11732), .B(n11669), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11702) );
  OR2_X1 U14637 ( .A1(n13106), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11701) );
  NAND2_X1 U14638 ( .A1(n11702), .A2(n11701), .ZN(n15650) );
  INV_X1 U14639 ( .A(n15650), .ZN(n11707) );
  INV_X1 U14640 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n21156) );
  NAND2_X1 U14641 ( .A1(n11717), .A2(n21156), .ZN(n11706) );
  NAND2_X1 U14642 ( .A1(n11737), .A2(n14605), .ZN(n11704) );
  NAND2_X1 U14643 ( .A1(n13217), .A2(n21156), .ZN(n11703) );
  NAND3_X1 U14644 ( .A1(n11704), .A2(n11681), .A3(n11703), .ZN(n11705) );
  NAND2_X1 U14645 ( .A1(n11706), .A2(n11705), .ZN(n15649) );
  NAND2_X1 U14646 ( .A1(n11707), .A2(n15649), .ZN(n11708) );
  MUX2_X1 U14647 ( .A(n11742), .B(n11737), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11712) );
  NAND2_X1 U14648 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n13129), .ZN(
        n11709) );
  AND2_X1 U14649 ( .A1(n11710), .A2(n11709), .ZN(n11711) );
  NAND2_X1 U14650 ( .A1(n11712), .A2(n11711), .ZN(n14434) );
  INV_X1 U14651 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n11713) );
  NAND2_X1 U14652 ( .A1(n11735), .A2(n11713), .ZN(n11716) );
  NAND2_X1 U14653 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11714) );
  OAI211_X1 U14654 ( .C1(n13129), .C2(P1_EBX_REG_20__SCAN_IN), .A(n11737), .B(
        n11714), .ZN(n11715) );
  AND2_X1 U14655 ( .A1(n11716), .A2(n11715), .ZN(n14384) );
  INV_X1 U14656 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n14427) );
  NAND2_X1 U14657 ( .A1(n11717), .A2(n14427), .ZN(n11721) );
  NAND2_X1 U14658 ( .A1(n11737), .A2(n14581), .ZN(n11719) );
  NAND2_X1 U14659 ( .A1(n13217), .A2(n14427), .ZN(n11718) );
  NAND3_X1 U14660 ( .A1(n11719), .A2(n11669), .A3(n11718), .ZN(n11720) );
  AND2_X1 U14661 ( .A1(n11721), .A2(n11720), .ZN(n14425) );
  NAND2_X1 U14662 ( .A1(n11681), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11722) );
  OAI211_X1 U14663 ( .C1(n13129), .C2(P1_EBX_REG_22__SCAN_IN), .A(n11737), .B(
        n11722), .ZN(n11723) );
  OAI21_X1 U14664 ( .B1(n11732), .B2(P1_EBX_REG_22__SCAN_IN), .A(n11723), .ZN(
        n15612) );
  MUX2_X1 U14665 ( .A(n11742), .B(n11737), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n11725) );
  NAND2_X1 U14666 ( .A1(n13129), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14667 ( .A1(n11725), .A2(n11724), .ZN(n14419) );
  NAND2_X1 U14668 ( .A1(n15611), .A2(n14419), .ZN(n14421) );
  MUX2_X1 U14669 ( .A(n11732), .B(n11669), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11726) );
  OAI21_X1 U14670 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n13106), .A(
        n11726), .ZN(n14371) );
  MUX2_X1 U14671 ( .A(n11742), .B(n11737), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n11728) );
  NAND2_X1 U14672 ( .A1(n13129), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14673 ( .A1(n11728), .A2(n11727), .ZN(n14358) );
  INV_X1 U14674 ( .A(n14358), .ZN(n11729) );
  NAND2_X1 U14675 ( .A1(n11669), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11730) );
  OAI211_X1 U14676 ( .C1(n13129), .C2(P1_EBX_REG_26__SCAN_IN), .A(n11737), .B(
        n11730), .ZN(n11731) );
  OAI21_X1 U14677 ( .B1(n11732), .B2(P1_EBX_REG_26__SCAN_IN), .A(n11731), .ZN(
        n14342) );
  NAND2_X1 U14678 ( .A1(n11737), .A2(n14675), .ZN(n11733) );
  OAI211_X1 U14679 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n13129), .A(n11733), .B(
        n11681), .ZN(n11734) );
  OAI21_X1 U14680 ( .B1(n11742), .B2(P1_EBX_REG_27__SCAN_IN), .A(n11734), .ZN(
        n14329) );
  INV_X1 U14681 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n20945) );
  NAND2_X1 U14682 ( .A1(n11735), .A2(n20945), .ZN(n11739) );
  NAND2_X1 U14683 ( .A1(n11669), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11736) );
  OAI211_X1 U14684 ( .C1(n13129), .C2(P1_EBX_REG_28__SCAN_IN), .A(n11737), .B(
        n11736), .ZN(n11738) );
  AND2_X1 U14685 ( .A1(n11739), .A2(n11738), .ZN(n14316) );
  OR2_X1 U14686 ( .A1(n13106), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11741) );
  INV_X1 U14687 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n20990) );
  NAND2_X1 U14688 ( .A1(n13217), .A2(n20990), .ZN(n11740) );
  NAND2_X1 U14689 ( .A1(n11741), .A2(n11740), .ZN(n14294) );
  OAI22_X1 U14690 ( .A1(n14294), .A2(n11692), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11742), .ZN(n14311) );
  XOR2_X1 U14691 ( .A(n11744), .B(n11743), .Z(n14408) );
  INV_X1 U14692 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20965) );
  NOR2_X1 U14693 ( .A1(n20135), .A2(n20965), .ZN(n13978) );
  NAND2_X1 U14694 ( .A1(n13442), .A2(n11745), .ZN(n11746) );
  AND2_X1 U14695 ( .A1(n11747), .A2(n11746), .ZN(n11753) );
  NAND2_X1 U14696 ( .A1(n11750), .A2(n11749), .ZN(n11751) );
  NAND2_X1 U14697 ( .A1(n11751), .A2(n13447), .ZN(n11754) );
  AND3_X1 U14698 ( .A1(n11754), .A2(n11753), .A3(n11752), .ZN(n11756) );
  OAI211_X1 U14699 ( .C1(n10406), .C2(n12958), .A(n11756), .B(n11755), .ZN(
        n13137) );
  NAND2_X1 U14700 ( .A1(n13135), .A2(n20149), .ZN(n11757) );
  NAND2_X1 U14701 ( .A1(n11758), .A2(n11757), .ZN(n11759) );
  OR2_X1 U14702 ( .A1(n13137), .A2(n11759), .ZN(n11760) );
  NAND2_X1 U14703 ( .A1(n11761), .A2(n11760), .ZN(n15822) );
  NAND2_X1 U14704 ( .A1(n15886), .A2(n15822), .ZN(n13229) );
  NOR2_X1 U14705 ( .A1(n10168), .A2(n20156), .ZN(n15506) );
  INV_X1 U14706 ( .A(n15827), .ZN(n15846) );
  INV_X1 U14707 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15823) );
  INV_X2 U14708 ( .A(n20135), .ZN(n15899) );
  NOR2_X1 U14709 ( .A1(n15899), .A2(n11761), .ZN(n15819) );
  AOI21_X1 U14710 ( .B1(n15821), .B2(n15823), .A(n15819), .ZN(n11768) );
  INV_X1 U14711 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14729) );
  INV_X1 U14712 ( .A(n14666), .ZN(n11767) );
  NAND2_X1 U14713 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15807) );
  INV_X1 U14714 ( .A(n15886), .ZN(n20143) );
  NOR2_X1 U14715 ( .A1(n11550), .A2(n13384), .ZN(n13553) );
  INV_X1 U14716 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14730) );
  OAI21_X1 U14717 ( .B1(n15823), .B2(n14730), .A(n11540), .ZN(n20133) );
  NAND2_X1 U14718 ( .A1(n13553), .A2(n20133), .ZN(n13623) );
  NOR2_X1 U14719 ( .A1(n11770), .A2(n13623), .ZN(n15817) );
  INV_X1 U14720 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15768) );
  INV_X1 U14721 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15923) );
  INV_X1 U14722 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15922) );
  INV_X1 U14723 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13736) );
  NOR3_X1 U14724 ( .A1(n15923), .A2(n15922), .A3(n13736), .ZN(n13794) );
  NAND3_X1 U14725 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n13794), .ZN(n15883) );
  NOR2_X1 U14726 ( .A1(n15768), .A2(n15883), .ZN(n15887) );
  NAND2_X1 U14727 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15887), .ZN(
        n15813) );
  NOR2_X1 U14728 ( .A1(n15878), .A2(n15813), .ZN(n11771) );
  NAND4_X1 U14729 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15829) );
  NOR2_X1 U14730 ( .A1(n15835), .A2(n15829), .ZN(n11772) );
  NAND3_X1 U14731 ( .A1(n15817), .A2(n11771), .A3(n11772), .ZN(n11763) );
  AND3_X1 U14732 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n13553), .ZN(n13621) );
  NAND2_X1 U14733 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13621), .ZN(
        n15882) );
  NOR2_X1 U14734 ( .A1(n15813), .A2(n15882), .ZN(n15812) );
  INV_X1 U14735 ( .A(n15812), .ZN(n15873) );
  NOR2_X1 U14736 ( .A1(n15878), .A2(n15873), .ZN(n15814) );
  AOI21_X1 U14737 ( .B1(n11772), .B2(n15814), .A(n13622), .ZN(n11762) );
  INV_X1 U14738 ( .A(n11768), .ZN(n13619) );
  AOI211_X1 U14739 ( .C1(n20143), .C2(n11763), .A(n11762), .B(n13619), .ZN(
        n15573) );
  NOR2_X1 U14740 ( .A1(n15827), .A2(n13619), .ZN(n13790) );
  AOI21_X1 U14741 ( .B1(n11773), .B2(n15573), .A(n13790), .ZN(n15809) );
  AOI21_X1 U14742 ( .B1(n15807), .B2(n15827), .A(n15809), .ZN(n14695) );
  NAND2_X1 U14743 ( .A1(n15827), .A2(n14687), .ZN(n11764) );
  NAND2_X1 U14744 ( .A1(n14695), .A2(n11764), .ZN(n15793) );
  NAND2_X1 U14745 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11765) );
  AND2_X1 U14746 ( .A1(n15827), .A2(n11765), .ZN(n11766) );
  NOR2_X1 U14747 ( .A1(n15793), .A2(n11766), .ZN(n14670) );
  OAI21_X1 U14748 ( .B1(n11767), .B2(n15846), .A(n14670), .ZN(n14657) );
  AOI211_X1 U14749 ( .C1(n11780), .C2(n15827), .A(n11617), .B(n14657), .ZN(
        n14647) );
  AOI211_X1 U14750 ( .C1(n15846), .C2(n11768), .A(n14729), .B(n14647), .ZN(
        n11769) );
  INV_X1 U14751 ( .A(n15817), .ZN(n13620) );
  NOR2_X1 U14752 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15816), .ZN(
        n13231) );
  NOR2_X1 U14753 ( .A1(n13231), .A2(n13622), .ZN(n14688) );
  NAND2_X1 U14754 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14688), .ZN(
        n20146) );
  NAND2_X1 U14755 ( .A1(n13553), .A2(n13380), .ZN(n13618) );
  INV_X1 U14756 ( .A(n11773), .ZN(n15570) );
  AND2_X1 U14757 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11774) );
  NAND2_X1 U14758 ( .A1(n15808), .A2(n11774), .ZN(n15795) );
  INV_X1 U14759 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14516) );
  INV_X1 U14760 ( .A(n11775), .ZN(n11776) );
  NOR2_X1 U14761 ( .A1(n14664), .A2(n11776), .ZN(n14649) );
  NAND3_X1 U14762 ( .A1(n14649), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n14729), .ZN(n11777) );
  OAI21_X1 U14763 ( .B1(n13983), .B2(n20138), .A(n11779), .ZN(P1_U3000) );
  XNOR2_X1 U14764 ( .A(n9820), .B(n11780), .ZN(n11781) );
  XNOR2_X1 U14765 ( .A(n9880), .B(n11781), .ZN(n14659) );
  NAND3_X1 U14766 ( .A1(n20718), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15947) );
  INV_X1 U14767 ( .A(n15947), .ZN(n11786) );
  NOR2_X2 U14768 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20658) );
  AND2_X2 U14769 ( .A1(n11786), .A2(n20658), .ZN(n15786) );
  INV_X1 U14770 ( .A(n15786), .ZN(n20131) );
  OR2_X1 U14771 ( .A1(n11787), .A2(n20658), .ZN(n20799) );
  AND2_X1 U14772 ( .A1(n20799), .A2(n20718), .ZN(n11788) );
  NAND2_X1 U14773 ( .A1(n20718), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15540) );
  INV_X1 U14774 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21127) );
  NAND2_X1 U14775 ( .A1(n21127), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n11789) );
  NAND2_X1 U14776 ( .A1(n15540), .A2(n11789), .ZN(n20124) );
  NAND2_X1 U14777 ( .A1(n15935), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14653) );
  OAI21_X1 U14778 ( .B1(n15790), .B2(n14310), .A(n14653), .ZN(n11790) );
  AND2_X2 U14779 ( .A1(n11851), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13691) );
  AND2_X4 U14780 ( .A1(n13691), .A2(n11872), .ZN(n12000) );
  AND2_X2 U14781 ( .A1(n14257), .A2(n11987), .ZN(n12149) );
  AND2_X4 U14782 ( .A1(n13691), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11999) );
  CLKBUF_X3 U14783 ( .A(n11999), .Z(n14256) );
  AOI22_X1 U14784 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12149), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11797) );
  AND2_X2 U14785 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12424) );
  AND2_X4 U14786 ( .A1(n12424), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14063) );
  AND2_X1 U14787 ( .A1(n14063), .A2(n11987), .ZN(n12148) );
  INV_X1 U14788 ( .A(n15317), .ZN(n14001) );
  AND2_X4 U14789 ( .A1(n15309), .A2(n11872), .ZN(n14262) );
  AOI22_X1 U14790 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12148), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11796) );
  AND2_X4 U14791 ( .A1(n11793), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14264) );
  AND2_X1 U14792 ( .A1(n14264), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11863) );
  AOI22_X1 U14793 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n11863), .ZN(n11795) );
  AND2_X1 U14794 ( .A1(n14264), .A2(n11987), .ZN(n12147) );
  AND2_X4 U14795 ( .A1(n16280), .A2(n13577), .ZN(n14265) );
  AOI22_X1 U14796 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12147), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11794) );
  NAND4_X1 U14797 ( .A1(n11797), .A2(n11796), .A3(n11795), .A4(n11794), .ZN(
        n11804) );
  AND2_X4 U14798 ( .A1(n13690), .A2(n11872), .ZN(n14263) );
  AND2_X2 U14799 ( .A1(n14263), .A2(n11987), .ZN(n12155) );
  AOI22_X1 U14800 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11802) );
  AND2_X4 U14801 ( .A1(n12424), .A2(n13577), .ZN(n12001) );
  AOI22_X1 U14802 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n12726), .B1(
        n11912), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11801) );
  AND2_X2 U14803 ( .A1(n14256), .A2(n11987), .ZN(n11896) );
  AOI22_X1 U14804 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14079), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11800) );
  AND2_X2 U14805 ( .A1(n14263), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14027) );
  NAND2_X1 U14806 ( .A1(n14258), .A2(n11987), .ZN(n14035) );
  INV_X2 U14807 ( .A(n14035), .ZN(n14078) );
  AOI22_X1 U14808 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11799) );
  NAND4_X1 U14809 ( .A1(n11802), .A2(n11801), .A3(n11800), .A4(n11799), .ZN(
        n11803) );
  AOI22_X1 U14810 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11805) );
  AND2_X1 U14811 ( .A1(n11805), .A2(n11987), .ZN(n11809) );
  AOI22_X1 U14812 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11808) );
  AOI22_X1 U14813 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11807) );
  AOI22_X1 U14814 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11806) );
  NAND4_X1 U14815 ( .A1(n11809), .A2(n11808), .A3(n11807), .A4(n11806), .ZN(
        n11816) );
  AOI22_X1 U14816 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11810) );
  AND2_X1 U14817 ( .A1(n11810), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11814) );
  AOI22_X1 U14818 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11813) );
  AOI22_X1 U14819 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14820 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11811) );
  NAND4_X1 U14821 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11815) );
  MUX2_X1 U14823 ( .A(n12769), .B(P2_EBX_REG_1__SCAN_IN), .S(n12264), .Z(
        n11817) );
  INV_X1 U14824 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13485) );
  AOI22_X1 U14825 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11821) );
  AOI22_X1 U14826 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11820) );
  AOI22_X1 U14827 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11819) );
  AOI22_X1 U14828 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11818) );
  NAND4_X1 U14829 ( .A1(n11821), .A2(n11820), .A3(n11819), .A4(n11818), .ZN(
        n11822) );
  NAND2_X1 U14830 ( .A1(n11822), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11829) );
  AOI22_X1 U14831 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U14832 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11825) );
  AOI22_X1 U14833 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U14834 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11823) );
  NAND4_X1 U14835 ( .A1(n11826), .A2(n11825), .A3(n11824), .A4(n11823), .ZN(
        n11827) );
  NAND2_X1 U14836 ( .A1(n11827), .A2(n11987), .ZN(n11828) );
  AOI22_X1 U14837 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14838 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14839 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14840 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14841 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14842 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14843 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U14844 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11839) );
  NAND2_X2 U14845 ( .A1(n12026), .A2(n12031), .ZN(n13489) );
  AOI22_X1 U14846 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n11896), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14847 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12149), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11843) );
  AOI22_X1 U14848 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n12148), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14849 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11841) );
  NAND4_X1 U14850 ( .A1(n11844), .A2(n11843), .A3(n11842), .A4(n11841), .ZN(
        n11850) );
  AOI22_X1 U14851 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14852 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14853 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12147), .B1(
        n11912), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U14854 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11863), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U14855 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11849) );
  NAND2_X1 U14856 ( .A1(n12017), .A2(n12603), .ZN(n11857) );
  MUX2_X1 U14857 ( .A(n13030), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n11856) );
  INV_X1 U14858 ( .A(n11856), .ZN(n11855) );
  NAND2_X1 U14859 ( .A1(n11851), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11852) );
  MUX2_X1 U14860 ( .A(n11856), .B(n11855), .S(n11871), .Z(n12415) );
  INV_X1 U14861 ( .A(n12415), .ZN(n12374) );
  NAND2_X1 U14862 ( .A1(n13489), .A2(n12374), .ZN(n12378) );
  NAND2_X1 U14863 ( .A1(n11857), .A2(n12378), .ZN(n12439) );
  MUX2_X1 U14864 ( .A(n13485), .B(n12439), .S(n10206), .Z(n12237) );
  AOI22_X1 U14865 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14866 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n9814), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14867 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n14078), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14868 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n14079), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11858) );
  NAND4_X1 U14869 ( .A1(n11861), .A2(n11860), .A3(n11859), .A4(n11858), .ZN(
        n11869) );
  AOI22_X1 U14870 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14871 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14872 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11912), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11865) );
  AOI22_X1 U14873 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12147), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11864) );
  NAND4_X1 U14874 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11868) );
  NAND2_X1 U14875 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13030), .ZN(
        n11870) );
  NAND2_X1 U14876 ( .A1(n11872), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11873) );
  XNOR2_X1 U14877 ( .A(n11987), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11889) );
  XNOR2_X1 U14878 ( .A(n11888), .B(n11889), .ZN(n12414) );
  INV_X1 U14879 ( .A(n12414), .ZN(n11875) );
  MUX2_X1 U14880 ( .A(n12612), .B(n11875), .S(n13489), .Z(n12382) );
  INV_X1 U14881 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13507) );
  MUX2_X1 U14882 ( .A(n12382), .B(n13507), .S(n12264), .Z(n12235) );
  AOI22_X1 U14883 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11880) );
  AOI22_X1 U14884 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n9814), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11879) );
  AOI22_X1 U14885 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n14079), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14886 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14078), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11877) );
  NAND4_X1 U14887 ( .A1(n11880), .A2(n11879), .A3(n11878), .A4(n11877), .ZN(
        n11887) );
  AOI22_X1 U14888 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14889 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14890 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12147), .B1(
        n11912), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14891 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n11863), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11882) );
  NAND4_X1 U14892 ( .A1(n11885), .A2(n11884), .A3(n11883), .A4(n11882), .ZN(
        n11886) );
  INV_X1 U14893 ( .A(n11889), .ZN(n11891) );
  NOR2_X1 U14894 ( .A1(n11987), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11890) );
  NOR2_X1 U14895 ( .A1(n16303), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11893) );
  INV_X1 U14896 ( .A(n12416), .ZN(n11894) );
  MUX2_X1 U14897 ( .A(n12781), .B(n11894), .S(n13489), .Z(n12383) );
  INV_X1 U14898 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19120) );
  MUX2_X1 U14899 ( .A(n12383), .B(n19120), .S(n12264), .Z(n11895) );
  AOI22_X1 U14900 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12149), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14901 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14902 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U14903 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11897) );
  NAND4_X1 U14904 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11906) );
  AOI22_X1 U14905 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14906 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14907 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14908 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11901) );
  NAND4_X1 U14909 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11905) );
  INV_X1 U14910 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n11907) );
  MUX2_X1 U14911 ( .A(n12199), .B(n11907), .S(n12264), .Z(n12229) );
  AOI22_X1 U14912 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11911) );
  AOI22_X1 U14913 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n9814), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11910) );
  AOI22_X1 U14914 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12148), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11909) );
  AOI22_X1 U14915 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11908) );
  NAND4_X1 U14916 ( .A1(n11911), .A2(n11910), .A3(n11909), .A4(n11908), .ZN(
        n11918) );
  AOI22_X1 U14917 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U14918 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11863), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U14919 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U14920 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U14921 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11917) );
  MUX2_X1 U14922 ( .A(n12626), .B(P2_EBX_REG_6__SCAN_IN), .S(n12264), .Z(
        n12224) );
  NAND2_X1 U14923 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U14924 ( .A1(n12149), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11921) );
  NAND2_X1 U14925 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11920) );
  NAND2_X1 U14926 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11919) );
  NAND2_X1 U14927 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U14928 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11925) );
  NAND2_X1 U14929 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11924) );
  NAND2_X1 U14930 ( .A1(n11862), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U14931 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11930) );
  NAND2_X1 U14932 ( .A1(n11863), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11929) );
  NAND2_X1 U14933 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11928) );
  NAND2_X1 U14934 ( .A1(n12147), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11927) );
  NAND2_X1 U14935 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11934) );
  NAND2_X1 U14936 ( .A1(n12726), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11933) );
  NAND2_X1 U14937 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11932) );
  NAND2_X1 U14938 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11931) );
  AND4_X2 U14939 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n13861) );
  MUX2_X1 U14940 ( .A(n13861), .B(P2_EBX_REG_7__SCAN_IN), .S(n12264), .Z(
        n12260) );
  INV_X1 U14941 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13399) );
  NAND2_X1 U14942 ( .A1(n12264), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12256) );
  NAND2_X1 U14943 ( .A1(n12264), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n12279) );
  AND2_X1 U14944 ( .A1(n12264), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12311) );
  INV_X1 U14945 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n12524) );
  INV_X1 U14946 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U14947 ( .A1(n12524), .A2(n12521), .ZN(n11939) );
  OR2_X2 U14948 ( .A1(n12308), .A2(n11940), .ZN(n12317) );
  NAND2_X1 U14949 ( .A1(n12264), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12301) );
  OAI21_X1 U14950 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(P2_EBX_REG_18__SCAN_IN), 
        .A(n12264), .ZN(n11941) );
  INV_X1 U14951 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14795) );
  NAND2_X1 U14952 ( .A1(n12264), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12342) );
  AND2_X1 U14953 ( .A1(n12264), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12345) );
  INV_X1 U14954 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14778) );
  AND3_X1 U14955 ( .A1(n12264), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n11946), .ZN(
        n11942) );
  NOR2_X1 U14956 ( .A1(n13955), .A2(n11942), .ZN(n16018) );
  NAND2_X1 U14957 ( .A1(n16018), .A2(n13959), .ZN(n12355) );
  NOR2_X1 U14958 ( .A1(n12353), .A2(n14778), .ZN(n11943) );
  NAND2_X1 U14959 ( .A1(n12264), .A2(n11943), .ZN(n11944) );
  AND2_X1 U14960 ( .A1(n12350), .A2(n11944), .ZN(n11945) );
  NAND2_X1 U14961 ( .A1(n11946), .A2(n11945), .ZN(n16029) );
  INV_X1 U14962 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15102) );
  OAI21_X1 U14963 ( .B1(n16029), .B2(n13861), .A(n15102), .ZN(n14934) );
  AOI22_X1 U14964 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U14965 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U14966 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U14967 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U14968 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NAND2_X1 U14969 ( .A1(n11951), .A2(n11987), .ZN(n11958) );
  AOI22_X1 U14970 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11955) );
  AOI22_X1 U14971 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U14972 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U14973 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11952) );
  NAND4_X1 U14974 ( .A1(n11955), .A2(n11954), .A3(n11953), .A4(n11952), .ZN(
        n11956) );
  NAND2_X1 U14975 ( .A1(n11956), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11957) );
  AOI22_X1 U14976 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11959) );
  AND2_X1 U14977 ( .A1(n11959), .A2(n11987), .ZN(n11963) );
  AOI22_X1 U14978 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U14979 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U14980 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11960) );
  NAND4_X1 U14981 ( .A1(n11963), .A2(n11962), .A3(n11961), .A4(n11960), .ZN(
        n11970) );
  AOI22_X1 U14982 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11964) );
  AND2_X1 U14983 ( .A1(n11964), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11968) );
  AOI22_X1 U14984 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11967) );
  AOI22_X1 U14985 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U14986 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11965) );
  NAND4_X1 U14987 ( .A1(n11968), .A2(n11967), .A3(n11966), .A4(n11965), .ZN(
        n11969) );
  AOI22_X1 U14988 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11974) );
  AOI22_X1 U14989 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11973) );
  AOI22_X1 U14990 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11972) );
  AOI22_X1 U14991 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11971) );
  NAND4_X1 U14992 ( .A1(n11974), .A2(n11973), .A3(n11972), .A4(n11971), .ZN(
        n11975) );
  NAND2_X1 U14993 ( .A1(n11975), .A2(n11987), .ZN(n11982) );
  AOI22_X1 U14994 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U14995 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11978) );
  AOI22_X1 U14996 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U14997 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11976) );
  NAND4_X1 U14998 ( .A1(n11979), .A2(n11978), .A3(n11977), .A4(n11976), .ZN(
        n11980) );
  NAND2_X1 U14999 ( .A1(n11980), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11981) );
  NAND2_X4 U15000 ( .A1(n11982), .A2(n11981), .ZN(n15344) );
  AOI22_X1 U15001 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15002 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15003 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15004 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11983) );
  AOI22_X1 U15005 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11999), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15006 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15007 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U15008 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15009 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15010 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15011 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11994) );
  NAND4_X1 U15012 ( .A1(n11997), .A2(n11996), .A3(n11995), .A4(n11994), .ZN(
        n11998) );
  NAND2_X1 U15013 ( .A1(n11998), .A2(n11987), .ZN(n12008) );
  AOI22_X1 U15014 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15015 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12003) );
  AOI22_X1 U15016 ( .A1(n14063), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12001), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12002) );
  NAND4_X1 U15017 ( .A1(n12005), .A2(n12004), .A3(n12003), .A4(n12002), .ZN(
        n12006) );
  NAND2_X1 U15018 ( .A1(n12006), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12007) );
  NAND2_X2 U15019 ( .A1(n12008), .A2(n12007), .ZN(n19283) );
  NAND2_X1 U15020 ( .A1(n12010), .A2(n12009), .ZN(n12450) );
  NOR2_X1 U15021 ( .A1(n12026), .A2(n19278), .ZN(n12013) );
  NAND4_X1 U15022 ( .A1(n12013), .A2(n12012), .A3(n12011), .A4(n13053), .ZN(
        n12402) );
  NAND2_X1 U15023 ( .A1(n12450), .A2(n12402), .ZN(n12457) );
  NAND2_X1 U15024 ( .A1(n12457), .A2(n12052), .ZN(n12021) );
  AND3_X2 U15025 ( .A1(n19273), .A2(n12023), .A3(n19278), .ZN(n12044) );
  NAND2_X1 U15026 ( .A1(n12014), .A2(n12026), .ZN(n12015) );
  NAND2_X1 U15027 ( .A1(n12021), .A2(n12020), .ZN(n12042) );
  NAND2_X1 U15028 ( .A1(n12454), .A2(n19278), .ZN(n12025) );
  NAND2_X1 U15029 ( .A1(n12053), .A2(n9959), .ZN(n12027) );
  NAND2_X1 U15030 ( .A1(n12042), .A2(n12027), .ZN(n12078) );
  OAI22_X1 U15031 ( .A1(n12078), .A2(n12029), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n13966), .ZN(n12083) );
  INV_X1 U15032 ( .A(n12030), .ZN(n13062) );
  AND2_X1 U15033 ( .A1(n15344), .A2(n19283), .ZN(n12032) );
  OAI211_X1 U15034 ( .C1(n13062), .C2(n12455), .A(n12407), .B(n12034), .ZN(
        n12576) );
  INV_X1 U15035 ( .A(n12576), .ZN(n12035) );
  NAND2_X1 U15036 ( .A1(n12035), .A2(n12458), .ZN(n12041) );
  INV_X1 U15037 ( .A(n12041), .ZN(n12036) );
  NAND2_X1 U15038 ( .A1(n12036), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12084) );
  NAND3_X1 U15039 ( .A1(n12083), .A2(n10234), .A3(n12084), .ZN(n12057) );
  INV_X1 U15040 ( .A(n12037), .ZN(n12038) );
  NAND4_X1 U15041 ( .A1(n12458), .A2(n12038), .A3(n12581), .A4(n13053), .ZN(
        n12039) );
  NAND2_X1 U15042 ( .A1(n12058), .A2(n12581), .ZN(n12040) );
  NAND2_X2 U15043 ( .A1(n12041), .A2(n12040), .ZN(n12575) );
  NAND2_X1 U15044 ( .A1(n12575), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12094) );
  INV_X1 U15045 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n12056) );
  INV_X1 U15046 ( .A(n12042), .ZN(n12051) );
  NAND2_X1 U15047 ( .A1(n13966), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n12049) );
  INV_X1 U15048 ( .A(n19972), .ZN(n16313) );
  NAND2_X1 U15049 ( .A1(n12044), .A2(n12043), .ZN(n12413) );
  INV_X1 U15050 ( .A(n12072), .ZN(n12046) );
  NAND2_X1 U15051 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15052 ( .A1(n12049), .A2(n16313), .A3(n12048), .A4(n12047), .ZN(
        n12050) );
  NOR2_X1 U15053 ( .A1(n12051), .A2(n12050), .ZN(n12055) );
  INV_X1 U15054 ( .A(n12052), .ZN(n12462) );
  NAND3_X1 U15055 ( .A1(n12053), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12462), 
        .ZN(n12054) );
  OAI211_X2 U15056 ( .C1(n12094), .C2(n12056), .A(n12055), .B(n12054), .ZN(
        n12082) );
  NAND2_X1 U15057 ( .A1(n12057), .A2(n12082), .ZN(n12081) );
  NAND2_X1 U15058 ( .A1(n12078), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12060) );
  AOI22_X1 U15059 ( .A1(n12058), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n19972), .ZN(n12059) );
  NAND2_X1 U15060 ( .A1(n12060), .A2(n12059), .ZN(n12068) );
  AND2_X1 U15061 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12066) );
  INV_X1 U15062 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n12061) );
  NAND2_X1 U15063 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  AOI21_X2 U15064 ( .B1(n12575), .B2(n12066), .A(n12065), .ZN(n12067) );
  XNOR2_X1 U15065 ( .A(n12068), .B(n12067), .ZN(n12110) );
  NAND2_X1 U15066 ( .A1(n12081), .A2(n12110), .ZN(n12071) );
  INV_X1 U15067 ( .A(n12067), .ZN(n12069) );
  INV_X1 U15068 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12245) );
  INV_X1 U15069 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n12075) );
  NAND2_X1 U15070 ( .A1(n13966), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U15071 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12073) );
  OAI211_X1 U15072 ( .C1(n13873), .C2(n12075), .A(n12074), .B(n12073), .ZN(
        n12076) );
  INV_X1 U15073 ( .A(n12076), .ZN(n12077) );
  OAI21_X2 U15074 ( .B1(n12481), .B2(n12245), .A(n12077), .ZN(n12089) );
  INV_X1 U15075 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13474) );
  OAI21_X1 U15076 ( .B1(n13030), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n13474), 
        .ZN(n12079) );
  XNOR2_X1 U15077 ( .A(n12089), .B(n12090), .ZN(n12080) );
  INV_X1 U15078 ( .A(n12082), .ZN(n12085) );
  NAND2_X1 U15079 ( .A1(n12085), .A2(n10225), .ZN(n12086) );
  INV_X1 U15080 ( .A(n12090), .ZN(n12087) );
  NAND2_X1 U15081 ( .A1(n12089), .A2(n12087), .ZN(n12088) );
  INV_X1 U15082 ( .A(n12089), .ZN(n12091) );
  NAND2_X1 U15083 ( .A1(n12091), .A2(n12090), .ZN(n12092) );
  INV_X1 U15084 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13419) );
  OR2_X1 U15085 ( .A1(n12094), .A2(n13419), .ZN(n12100) );
  INV_X1 U15086 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13425) );
  INV_X1 U15087 ( .A(n13966), .ZN(n12095) );
  NAND2_X1 U15088 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12096) );
  OAI211_X1 U15089 ( .C1(n13873), .C2(n13425), .A(n12097), .B(n12096), .ZN(
        n12098) );
  INV_X1 U15090 ( .A(n12098), .ZN(n12099) );
  AND2_X1 U15091 ( .A1(n19972), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12101) );
  AOI21_X1 U15092 ( .B1(n12102), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12101), .ZN(n12104) );
  NAND2_X1 U15093 ( .A1(n12103), .A2(n12104), .ZN(n12487) );
  INV_X1 U15094 ( .A(n12104), .ZN(n12105) );
  NAND2_X1 U15095 ( .A1(n12106), .A2(n12105), .ZN(n12107) );
  OR2_X2 U15096 ( .A1(n12141), .A2(n13099), .ZN(n12113) );
  NOR2_X2 U15097 ( .A1(n12113), .A2(n13910), .ZN(n19356) );
  INV_X1 U15098 ( .A(n15332), .ZN(n12114) );
  INV_X1 U15099 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12118) );
  INV_X1 U15100 ( .A(n19076), .ZN(n16252) );
  INV_X1 U15101 ( .A(n12136), .ZN(n12116) );
  INV_X1 U15102 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14102) );
  OAI22_X1 U15103 ( .A1(n12118), .A2(n19595), .B1(n19734), .B2(n14102), .ZN(
        n12119) );
  INV_X1 U15104 ( .A(n12119), .ZN(n12123) );
  INV_X1 U15105 ( .A(n12125), .ZN(n12120) );
  AND2_X1 U15106 ( .A1(n19076), .A2(n12120), .ZN(n12137) );
  INV_X1 U15107 ( .A(n12185), .ZN(n19686) );
  AOI21_X1 U15108 ( .B1(n19686), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n12584), .ZN(n12122) );
  INV_X1 U15109 ( .A(n19660), .ZN(n19653) );
  NAND2_X1 U15110 ( .A1(n19653), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12121) );
  NAND3_X1 U15111 ( .A1(n12124), .A2(n12123), .A3(n10228), .ZN(n12165) );
  AND2_X1 U15112 ( .A1(n12125), .A2(n19076), .ZN(n12127) );
  INV_X1 U15113 ( .A(n12127), .ZN(n12126) );
  INV_X1 U15114 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14093) );
  INV_X1 U15115 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12128) );
  OAI22_X1 U15116 ( .A1(n12129), .A2(n14093), .B1(n19620), .B2(n12128), .ZN(
        n12135) );
  INV_X1 U15117 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12133) );
  INV_X1 U15118 ( .A(n12130), .ZN(n12131) );
  INV_X1 U15119 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14101) );
  OAI22_X1 U15120 ( .A1(n12133), .A2(n19564), .B1(n19765), .B2(n14101), .ZN(
        n12134) );
  NOR2_X1 U15121 ( .A1(n12135), .A2(n12134), .ZN(n12146) );
  AOI22_X1 U15122 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19423), .B1(
        n15354), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12145) );
  INV_X1 U15123 ( .A(n12137), .ZN(n12138) );
  NOR2_X2 U15124 ( .A1(n12140), .A2(n19251), .ZN(n19302) );
  NOR2_X2 U15125 ( .A1(n12139), .A2(n19251), .ZN(n19392) );
  AOI22_X1 U15126 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19302), .B1(
        n19392), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12144) );
  NOR2_X2 U15127 ( .A1(n12140), .A2(n16283), .ZN(n19454) );
  INV_X1 U15128 ( .A(n12181), .ZN(n19529) );
  NAND4_X1 U15129 ( .A1(n12146), .A2(n12145), .A3(n12144), .A4(n12143), .ZN(
        n12164) );
  AOI22_X1 U15130 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12153) );
  AOI22_X1 U15131 ( .A1(n12149), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U15132 ( .A1(n14078), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15133 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14079), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12150) );
  NAND4_X1 U15134 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12162) );
  AOI22_X1 U15135 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11912), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15136 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15137 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15138 ( .A1(n9814), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12157) );
  NAND4_X1 U15139 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12161) );
  NOR2_X1 U15140 ( .A1(n12162), .A2(n12161), .ZN(n12770) );
  OR2_X1 U15141 ( .A1(n12770), .A2(n19976), .ZN(n12953) );
  NOR2_X1 U15142 ( .A1(n12953), .A2(n12769), .ZN(n12774) );
  OR2_X1 U15143 ( .A1(n12774), .A2(n12603), .ZN(n12163) );
  OAI21_X2 U15144 ( .B1(n12165), .B2(n12164), .A(n12163), .ZN(n12233) );
  INV_X1 U15145 ( .A(n12233), .ZN(n12180) );
  AOI22_X1 U15146 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19356), .B1(
        n15354), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15147 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19392), .B1(
        n12192), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12166) );
  AOI22_X1 U15148 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19454), .B1(
        n19302), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12169) );
  NAND2_X1 U15149 ( .A1(n19423), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n12168) );
  INV_X1 U15150 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12171) );
  INV_X1 U15151 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12170) );
  OAI22_X1 U15152 ( .A1(n12171), .A2(n12185), .B1(n19564), .B2(n12170), .ZN(
        n12174) );
  INV_X1 U15153 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12172) );
  INV_X1 U15154 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14155) );
  OAI22_X1 U15155 ( .A1(n12172), .A2(n19620), .B1(n19765), .B2(n14155), .ZN(
        n12173) );
  INV_X1 U15156 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14157) );
  INV_X1 U15157 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14156) );
  OAI22_X1 U15158 ( .A1(n14157), .A2(n12181), .B1(n19734), .B2(n14156), .ZN(
        n12177) );
  INV_X1 U15159 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12175) );
  INV_X1 U15160 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14158) );
  OAI22_X1 U15161 ( .A1(n12175), .A2(n19595), .B1(n19660), .B2(n14158), .ZN(
        n12176) );
  NAND2_X2 U15162 ( .A1(n12179), .A2(n12178), .ZN(n12234) );
  INV_X1 U15163 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14204) );
  INV_X1 U15164 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14213) );
  INV_X1 U15165 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14212) );
  OAI22_X1 U15166 ( .A1(n14213), .A2(n12181), .B1(n19734), .B2(n14212), .ZN(
        n12184) );
  INV_X1 U15167 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12182) );
  INV_X1 U15168 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14214) );
  OAI22_X1 U15169 ( .A1(n12182), .A2(n19595), .B1(n19660), .B2(n14214), .ZN(
        n12183) );
  NOR2_X1 U15170 ( .A1(n12184), .A2(n12183), .ZN(n12191) );
  INV_X1 U15171 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12186) );
  INV_X1 U15172 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14034) );
  OAI22_X1 U15173 ( .A1(n12186), .A2(n12185), .B1(n19564), .B2(n14034), .ZN(
        n12189) );
  INV_X1 U15174 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12187) );
  INV_X1 U15175 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14211) );
  OAI22_X1 U15176 ( .A1(n12187), .A2(n19620), .B1(n19765), .B2(n14211), .ZN(
        n12188) );
  NOR2_X1 U15177 ( .A1(n12189), .A2(n12188), .ZN(n12190) );
  OAI211_X1 U15178 ( .C1(n14204), .C2(n15332), .A(n12191), .B(n12190), .ZN(
        n12198) );
  AOI22_X1 U15179 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19356), .B1(
        n15354), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15180 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19392), .B1(
        n12192), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15181 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19454), .B1(
        n19302), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12194) );
  NAND2_X1 U15182 ( .A1(n19423), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n12193) );
  NAND4_X1 U15183 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12197) );
  INV_X1 U15184 ( .A(n12199), .ZN(n12623) );
  NAND2_X1 U15185 ( .A1(n12623), .A2(n12584), .ZN(n12200) );
  NAND2_X1 U15186 ( .A1(n12202), .A2(n12227), .ZN(n12222) );
  INV_X1 U15187 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19299) );
  INV_X1 U15188 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14238) );
  INV_X1 U15189 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14234) );
  OAI22_X1 U15190 ( .A1(n14238), .A2(n19660), .B1(n19734), .B2(n14234), .ZN(
        n12205) );
  INV_X1 U15191 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12203) );
  INV_X1 U15192 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14236) );
  OAI22_X1 U15193 ( .A1(n12203), .A2(n19595), .B1(n12181), .B2(n14236), .ZN(
        n12204) );
  NOR2_X1 U15194 ( .A1(n12205), .A2(n12204), .ZN(n12212) );
  INV_X1 U15195 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12207) );
  INV_X1 U15196 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12206) );
  OAI22_X1 U15197 ( .A1(n12207), .A2(n19564), .B1(n19620), .B2(n12206), .ZN(
        n12210) );
  INV_X1 U15198 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12208) );
  INV_X1 U15199 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14232) );
  OAI22_X1 U15200 ( .A1(n12208), .A2(n12185), .B1(n19765), .B2(n14232), .ZN(
        n12209) );
  NOR2_X1 U15201 ( .A1(n12210), .A2(n12209), .ZN(n12211) );
  OAI211_X1 U15202 ( .C1(n19299), .C2(n15332), .A(n12212), .B(n12211), .ZN(
        n12218) );
  AOI22_X1 U15203 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19356), .B1(
        n15354), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12216) );
  AOI22_X1 U15204 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19302), .B1(
        n19392), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12215) );
  AOI22_X1 U15205 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19454), .B1(
        n12192), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12214) );
  NAND2_X1 U15206 ( .A1(n19423), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n12213) );
  NAND4_X1 U15207 ( .A1(n12216), .A2(n12215), .A3(n12214), .A4(n12213), .ZN(
        n12217) );
  NAND2_X1 U15208 ( .A1(n12626), .A2(n12584), .ZN(n12219) );
  NAND2_X1 U15209 ( .A1(n12222), .A2(n12790), .ZN(n12223) );
  NAND2_X1 U15210 ( .A1(n12231), .A2(n12224), .ZN(n12225) );
  NAND2_X1 U15211 ( .A1(n12261), .A2(n12225), .ZN(n19004) );
  INV_X1 U15212 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15272) );
  NAND2_X1 U15213 ( .A1(n12787), .A2(n13861), .ZN(n12232) );
  OR2_X1 U15214 ( .A1(n12248), .A2(n12229), .ZN(n12230) );
  NAND2_X1 U15215 ( .A1(n12231), .A2(n12230), .ZN(n19014) );
  NAND2_X2 U15216 ( .A1(n12232), .A2(n19014), .ZN(n12251) );
  XNOR2_X2 U15217 ( .A(n12251), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15283) );
  OAI21_X1 U15218 ( .B1(n12236), .B2(n12235), .A(n12247), .ZN(n13503) );
  INV_X1 U15219 ( .A(n12236), .ZN(n12239) );
  OR2_X1 U15220 ( .A1(n12241), .A2(n12237), .ZN(n12238) );
  NAND2_X1 U15221 ( .A1(n12239), .A2(n12238), .ZN(n13490) );
  OAI21_X1 U15222 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19958), .A(
        n12372), .ZN(n12375) );
  MUX2_X1 U15223 ( .A(n12770), .B(n12375), .S(n13489), .Z(n12438) );
  INV_X1 U15224 ( .A(n12240), .ZN(n12243) );
  OAI21_X1 U15225 ( .B1(n12438), .B2(n12264), .A(n12243), .ZN(n19063) );
  NAND2_X1 U15226 ( .A1(n19063), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13890) );
  INV_X1 U15227 ( .A(n12241), .ZN(n12242) );
  OAI21_X1 U15228 ( .B1(n9961), .B2(n12243), .A(n12242), .ZN(n19050) );
  NOR2_X1 U15229 ( .A1(n13890), .A2(n19050), .ZN(n12244) );
  NAND2_X1 U15230 ( .A1(n13890), .A2(n19050), .ZN(n13889) );
  OAI21_X1 U15231 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12244), .A(
        n13889), .ZN(n13069) );
  XNOR2_X1 U15232 ( .A(n13490), .B(n12245), .ZN(n13068) );
  OR2_X1 U15233 ( .A1(n13069), .A2(n13068), .ZN(n13071) );
  OAI21_X1 U15234 ( .B1(n13490), .B2(n12245), .A(n13071), .ZN(n13420) );
  AND2_X1 U15235 ( .A1(n12247), .A2(n12246), .ZN(n12249) );
  OR2_X1 U15236 ( .A1(n12249), .A2(n12248), .ZN(n19037) );
  XNOR2_X1 U15237 ( .A(n19037), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19231) );
  INV_X1 U15238 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19259) );
  NOR2_X1 U15239 ( .A1(n19037), .A2(n19259), .ZN(n12250) );
  NAND2_X1 U15240 ( .A1(n12251), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12252) );
  NAND2_X1 U15241 ( .A1(n13727), .A2(n13728), .ZN(n12255) );
  NAND2_X1 U15242 ( .A1(n12253), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12254) );
  OR2_X1 U15243 ( .A1(n12257), .A2(n12256), .ZN(n12258) );
  NAND2_X1 U15244 ( .A1(n12266), .A2(n12258), .ZN(n18983) );
  INV_X1 U15245 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16227) );
  OR2_X1 U15246 ( .A1(n13861), .A2(n16227), .ZN(n12259) );
  OR2_X1 U15247 ( .A1(n18983), .A2(n12259), .ZN(n16151) );
  XNOR2_X1 U15248 ( .A(n12261), .B(n10076), .ZN(n18992) );
  NAND2_X1 U15249 ( .A1(n18992), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16153) );
  OR2_X1 U15250 ( .A1(n18983), .A2(n13861), .ZN(n12262) );
  NAND2_X1 U15251 ( .A1(n12262), .A2(n16227), .ZN(n16152) );
  OR2_X1 U15252 ( .A1(n18992), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15052) );
  AND2_X1 U15253 ( .A1(n16152), .A2(n15052), .ZN(n12263) );
  NAND2_X1 U15254 ( .A1(n12264), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12265) );
  XNOR2_X1 U15255 ( .A(n12266), .B(n12265), .ZN(n18970) );
  NAND2_X1 U15256 ( .A1(n18970), .A2(n13959), .ZN(n12271) );
  INV_X1 U15257 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n13936) );
  AND2_X1 U15258 ( .A1(n12271), .A2(n13936), .ZN(n13929) );
  OR2_X1 U15259 ( .A1(n12267), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12269) );
  NAND3_X1 U15260 ( .A1(n12267), .A2(n12264), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n12268) );
  NAND3_X1 U15261 ( .A1(n12269), .A2(n12268), .A3(n12350), .ZN(n18962) );
  INV_X1 U15262 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12506) );
  OAI21_X1 U15263 ( .B1(n18962), .B2(n13861), .A(n12506), .ZN(n16138) );
  OR2_X1 U15264 ( .A1(n13861), .A2(n12506), .ZN(n12270) );
  OR2_X1 U15265 ( .A1(n18962), .A2(n12270), .ZN(n16137) );
  OR2_X1 U15266 ( .A1(n12271), .A2(n13936), .ZN(n13928) );
  AND2_X1 U15267 ( .A1(n16137), .A2(n13928), .ZN(n12272) );
  AND3_X1 U15268 ( .A1(n12264), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n12269), .ZN(
        n12273) );
  NOR2_X1 U15269 ( .A1(n12274), .A2(n12273), .ZN(n18953) );
  NAND2_X1 U15270 ( .A1(n18953), .A2(n13959), .ZN(n15251) );
  INV_X1 U15271 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15258) );
  NOR2_X1 U15272 ( .A1(n15251), .A2(n15258), .ZN(n12275) );
  NAND2_X1 U15273 ( .A1(n15251), .A2(n15258), .ZN(n12276) );
  INV_X1 U15274 ( .A(n12277), .ZN(n12278) );
  OR2_X1 U15275 ( .A1(n12279), .A2(n12278), .ZN(n12280) );
  NAND2_X1 U15276 ( .A1(n12313), .A2(n12280), .ZN(n18941) );
  OR2_X1 U15277 ( .A1(n18941), .A2(n13861), .ZN(n12281) );
  INV_X1 U15278 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12512) );
  NAND2_X1 U15279 ( .A1(n12281), .A2(n12512), .ZN(n13912) );
  INV_X1 U15280 ( .A(n13911), .ZN(n12282) );
  NAND2_X1 U15281 ( .A1(n12264), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12283) );
  NOR2_X1 U15282 ( .A1(n12286), .A2(n12283), .ZN(n12284) );
  OR2_X1 U15283 ( .A1(n12285), .A2(n12284), .ZN(n18851) );
  NOR2_X1 U15284 ( .A1(n18851), .A2(n13861), .ZN(n12339) );
  NOR2_X1 U15285 ( .A1(n12339), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14964) );
  INV_X1 U15286 ( .A(n12286), .ZN(n12289) );
  NAND2_X1 U15287 ( .A1(n12264), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12287) );
  MUX2_X1 U15288 ( .A(n12264), .B(n12287), .S(n12322), .Z(n12288) );
  NAND2_X1 U15289 ( .A1(n12289), .A2(n12288), .ZN(n18861) );
  INV_X1 U15290 ( .A(n18861), .ZN(n12290) );
  AOI21_X1 U15291 ( .B1(n12290), .B2(n13959), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14976) );
  NAND2_X1 U15292 ( .A1(n12264), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12291) );
  MUX2_X1 U15293 ( .A(n12291), .B(n12264), .S(n12299), .Z(n12293) );
  INV_X1 U15294 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n12292) );
  NAND2_X1 U15295 ( .A1(n12299), .A2(n12292), .ZN(n12321) );
  NAND2_X1 U15296 ( .A1(n12293), .A2(n12321), .ZN(n18879) );
  INV_X1 U15297 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15196) );
  OAI21_X1 U15298 ( .B1(n18879), .B2(n13861), .A(n15196), .ZN(n15002) );
  AND2_X1 U15299 ( .A1(n12264), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12295) );
  INV_X1 U15300 ( .A(n12350), .ZN(n12294) );
  AOI21_X1 U15301 ( .B1(n12317), .B2(n12295), .A(n12294), .ZN(n12297) );
  NAND2_X1 U15302 ( .A1(n12297), .A2(n12296), .ZN(n18901) );
  NOR2_X1 U15303 ( .A1(n18901), .A2(n13861), .ZN(n12298) );
  INV_X1 U15304 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15230) );
  XNOR2_X1 U15305 ( .A(n12298), .B(n15230), .ZN(n15027) );
  INV_X1 U15306 ( .A(n12299), .ZN(n12305) );
  INV_X1 U15307 ( .A(n12300), .ZN(n12303) );
  INV_X1 U15308 ( .A(n12301), .ZN(n12302) );
  NAND2_X1 U15309 ( .A1(n12303), .A2(n12302), .ZN(n12304) );
  NAND2_X1 U15310 ( .A1(n12305), .A2(n12304), .ZN(n18893) );
  OR2_X1 U15311 ( .A1(n18893), .A2(n13861), .ZN(n12306) );
  INV_X1 U15312 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12530) );
  NAND2_X1 U15313 ( .A1(n12306), .A2(n12530), .ZN(n15018) );
  NAND2_X1 U15314 ( .A1(n12264), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12307) );
  MUX2_X1 U15315 ( .A(n12264), .B(n12307), .S(n12308), .Z(n12309) );
  OR2_X1 U15316 ( .A1(n12308), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12316) );
  NAND2_X1 U15317 ( .A1(n12309), .A2(n12316), .ZN(n18920) );
  OR2_X1 U15318 ( .A1(n18920), .A2(n13861), .ZN(n12310) );
  INV_X1 U15319 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16210) );
  NAND2_X1 U15320 ( .A1(n12310), .A2(n16210), .ZN(n16111) );
  INV_X1 U15321 ( .A(n12311), .ZN(n12312) );
  XNOR2_X1 U15322 ( .A(n12313), .B(n12312), .ZN(n18933) );
  NAND2_X1 U15323 ( .A1(n18933), .A2(n13959), .ZN(n12314) );
  INV_X1 U15324 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15242) );
  NAND2_X1 U15325 ( .A1(n12314), .A2(n15242), .ZN(n15233) );
  AND2_X1 U15326 ( .A1(n12264), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12315) );
  NAND2_X1 U15327 ( .A1(n12316), .A2(n12315), .ZN(n12318) );
  NAND2_X1 U15328 ( .A1(n12318), .A2(n12317), .ZN(n18910) );
  OR2_X1 U15329 ( .A1(n18910), .A2(n13861), .ZN(n12319) );
  INV_X1 U15330 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16187) );
  NAND2_X1 U15331 ( .A1(n12319), .A2(n16187), .ZN(n15041) );
  AND4_X1 U15332 ( .A1(n15018), .A2(n16111), .A3(n15233), .A4(n15041), .ZN(
        n12325) );
  AND2_X1 U15333 ( .A1(n12264), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U15334 ( .A1(n12321), .A2(n12320), .ZN(n12323) );
  NAND2_X1 U15335 ( .A1(n12323), .A2(n12322), .ZN(n18872) );
  OR2_X1 U15336 ( .A1(n18872), .A2(n13861), .ZN(n12324) );
  INV_X1 U15337 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15177) );
  NAND2_X1 U15338 ( .A1(n12324), .A2(n15177), .ZN(n14993) );
  NAND4_X1 U15339 ( .A1(n15002), .A2(n15027), .A3(n12325), .A4(n14993), .ZN(
        n12326) );
  INV_X1 U15340 ( .A(n18879), .ZN(n12330) );
  NOR2_X1 U15341 ( .A1(n13861), .A2(n15196), .ZN(n12329) );
  NAND2_X1 U15342 ( .A1(n12330), .A2(n12329), .ZN(n15001) );
  OR2_X1 U15343 ( .A1(n13861), .A2(n15177), .ZN(n12331) );
  OR2_X1 U15344 ( .A1(n18872), .A2(n12331), .ZN(n14992) );
  AND2_X1 U15345 ( .A1(n15001), .A2(n14992), .ZN(n14960) );
  OR2_X1 U15346 ( .A1(n13861), .A2(n12530), .ZN(n12332) );
  OR2_X1 U15347 ( .A1(n18893), .A2(n12332), .ZN(n15017) );
  INV_X1 U15348 ( .A(n18901), .ZN(n12334) );
  NOR2_X1 U15349 ( .A1(n13861), .A2(n15230), .ZN(n12333) );
  NAND2_X1 U15350 ( .A1(n12334), .A2(n12333), .ZN(n15019) );
  OR2_X1 U15351 ( .A1(n13861), .A2(n16210), .ZN(n12335) );
  OR2_X1 U15352 ( .A1(n18920), .A2(n12335), .ZN(n16110) );
  OR2_X1 U15353 ( .A1(n13861), .A2(n16187), .ZN(n12336) );
  OR2_X1 U15354 ( .A1(n18910), .A2(n12336), .ZN(n15040) );
  AND2_X1 U15355 ( .A1(n16110), .A2(n15040), .ZN(n14958) );
  NOR2_X1 U15356 ( .A1(n13861), .A2(n15242), .ZN(n12337) );
  NAND2_X1 U15357 ( .A1(n18933), .A2(n12337), .ZN(n15232) );
  INV_X1 U15358 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15164) );
  OR2_X1 U15359 ( .A1(n13861), .A2(n15164), .ZN(n12338) );
  NOR2_X1 U15360 ( .A1(n18861), .A2(n12338), .ZN(n14975) );
  INV_X1 U15361 ( .A(n14975), .ZN(n14962) );
  INV_X1 U15362 ( .A(n12339), .ZN(n12340) );
  INV_X1 U15363 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15588) );
  NOR2_X1 U15364 ( .A1(n12340), .A2(n15588), .ZN(n14963) );
  AOI21_X1 U15365 ( .B1(n10082), .B2(n12343), .A(n9859), .ZN(n15480) );
  NAND2_X1 U15366 ( .A1(n15480), .A2(n13959), .ZN(n12344) );
  INV_X1 U15367 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15141) );
  NAND2_X1 U15368 ( .A1(n12344), .A2(n15141), .ZN(n15133) );
  NOR2_X1 U15369 ( .A1(n12344), .A2(n15141), .ZN(n15135) );
  AOI21_X1 U15370 ( .B1(n15137), .B2(n15133), .A(n15135), .ZN(n14944) );
  XNOR2_X1 U15371 ( .A(n9859), .B(n12345), .ZN(n16052) );
  NAND2_X1 U15372 ( .A1(n16052), .A2(n13959), .ZN(n12346) );
  XOR2_X1 U15373 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n12346), .Z(
        n14943) );
  INV_X1 U15374 ( .A(n12346), .ZN(n12347) );
  NAND3_X1 U15375 ( .A1(n12349), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n12264), 
        .ZN(n12351) );
  NAND2_X1 U15376 ( .A1(n12351), .A2(n12350), .ZN(n12352) );
  OR2_X1 U15377 ( .A1(n12353), .A2(n12352), .ZN(n16044) );
  NOR2_X1 U15378 ( .A1(n12354), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15109) );
  INV_X1 U15379 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15091) );
  OR2_X1 U15380 ( .A1(n12355), .A2(n15091), .ZN(n12356) );
  NAND2_X1 U15381 ( .A1(n14933), .A2(n12356), .ZN(n13850) );
  INV_X1 U15382 ( .A(n13850), .ZN(n12357) );
  AND2_X2 U15383 ( .A1(n13848), .A2(n12357), .ZN(n12364) );
  NAND2_X1 U15384 ( .A1(n12264), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12360) );
  INV_X1 U15385 ( .A(n12358), .ZN(n12359) );
  NOR2_X1 U15386 ( .A1(n12360), .A2(n12359), .ZN(n12361) );
  NOR2_X1 U15387 ( .A1(n12366), .A2(n12361), .ZN(n16005) );
  NAND2_X1 U15388 ( .A1(n16005), .A2(n13959), .ZN(n12363) );
  OR2_X1 U15389 ( .A1(n12364), .A2(n12363), .ZN(n12365) );
  NAND2_X1 U15390 ( .A1(n12264), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12367) );
  INV_X1 U15391 ( .A(n12366), .ZN(n12369) );
  INV_X1 U15392 ( .A(n12367), .ZN(n12368) );
  NAND2_X1 U15393 ( .A1(n12369), .A2(n12368), .ZN(n12370) );
  XOR2_X1 U15394 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n13849), .Z(
        n12371) );
  INV_X1 U15395 ( .A(n12375), .ZN(n12427) );
  XNOR2_X1 U15396 ( .A(n12437), .B(n12372), .ZN(n12418) );
  OAI21_X1 U15397 ( .B1(n19976), .B2(n12415), .A(n12418), .ZN(n12373) );
  OAI211_X1 U15398 ( .C1(n12374), .C2(n12427), .A(n12373), .B(n13045), .ZN(
        n12381) );
  OAI21_X1 U15399 ( .B1(n12375), .B2(n12437), .A(n12017), .ZN(n12380) );
  NAND2_X1 U15400 ( .A1(n12376), .A2(n19976), .ZN(n12377) );
  NAND2_X1 U15401 ( .A1(n12377), .A2(n12415), .ZN(n12379) );
  AOI22_X1 U15402 ( .A1(n12381), .A2(n12380), .B1(n12379), .B2(n12378), .ZN(
        n12385) );
  NAND2_X1 U15403 ( .A1(n12383), .A2(n12382), .ZN(n12444) );
  NAND2_X1 U15404 ( .A1(n12444), .A2(n13489), .ZN(n12384) );
  OAI21_X1 U15405 ( .B1(n12414), .B2(n12385), .A(n12384), .ZN(n12392) );
  INV_X1 U15406 ( .A(n12386), .ZN(n12388) );
  NAND2_X1 U15407 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13013), .ZN(
        n12389) );
  NAND2_X1 U15408 ( .A1(n12017), .A2(n12416), .ZN(n12391) );
  NAND3_X1 U15409 ( .A1(n12392), .A2(n12442), .A3(n12391), .ZN(n12393) );
  MUX2_X1 U15410 ( .A(n12393), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n13470), .Z(n12398) );
  INV_X1 U15411 ( .A(n12442), .ZN(n12394) );
  NAND2_X1 U15412 ( .A1(n12394), .A2(n12977), .ZN(n12395) );
  NOR2_X1 U15413 ( .A1(n13001), .A2(n12584), .ZN(n12397) );
  NOR2_X1 U15414 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19847) );
  AOI211_X1 U15415 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19847), .ZN(n19977) );
  NAND2_X1 U15416 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19838) );
  NAND2_X1 U15417 ( .A1(n19977), .A2(n19838), .ZN(n13482) );
  INV_X1 U15418 ( .A(n13482), .ZN(n12994) );
  NAND3_X1 U15419 ( .A1(n12397), .A2(n12994), .A3(n12396), .ZN(n12447) );
  INV_X1 U15420 ( .A(n12397), .ZN(n12400) );
  AOI21_X1 U15421 ( .B1(n12398), .B2(n13045), .A(n12023), .ZN(n12399) );
  NAND2_X1 U15422 ( .A1(n12400), .A2(n12399), .ZN(n12446) );
  INV_X1 U15423 ( .A(n13045), .ZN(n16274) );
  NAND2_X1 U15424 ( .A1(n16274), .A2(n15344), .ZN(n12401) );
  NAND2_X1 U15425 ( .A1(n12401), .A2(n19273), .ZN(n12406) );
  NAND2_X1 U15426 ( .A1(n12403), .A2(n19273), .ZN(n12404) );
  NAND2_X1 U15427 ( .A1(n13011), .A2(n12404), .ZN(n12405) );
  OAI211_X1 U15428 ( .C1(n12407), .C2(n12406), .A(n12405), .B(n9819), .ZN(
        n12408) );
  INV_X1 U15429 ( .A(n12408), .ZN(n12412) );
  OR2_X1 U15430 ( .A1(n12410), .A2(n13064), .ZN(n12411) );
  NAND2_X1 U15431 ( .A1(n12411), .A2(n16312), .ZN(n12456) );
  INV_X1 U15432 ( .A(n12413), .ZN(n12421) );
  NOR3_X1 U15433 ( .A1(n12416), .A2(n12415), .A3(n12414), .ZN(n12426) );
  INV_X1 U15434 ( .A(n12426), .ZN(n12417) );
  INV_X1 U15435 ( .A(n16267), .ZN(n12420) );
  NAND3_X1 U15436 ( .A1(n12421), .A2(n12420), .A3(n12994), .ZN(n12422) );
  NAND2_X1 U15437 ( .A1(n12452), .A2(n12422), .ZN(n12996) );
  MUX2_X1 U15438 ( .A(n12413), .B(n19273), .S(n12584), .Z(n12435) );
  INV_X1 U15439 ( .A(n19838), .ZN(n19980) );
  OR2_X1 U15440 ( .A1(n16267), .A2(n19980), .ZN(n12434) );
  NAND2_X1 U15441 ( .A1(n15314), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12425) );
  NAND2_X1 U15442 ( .A1(n12425), .A2(n13013), .ZN(n13009) );
  INV_X1 U15443 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n13006) );
  OAI211_X1 U15444 ( .C1(n9815), .C2(n13009), .A(P2_STATE2_REG_1__SCAN_IN), 
        .B(n13006), .ZN(n19954) );
  AOI21_X1 U15445 ( .B1(n12427), .B2(n12426), .A(n16267), .ZN(n12428) );
  INV_X1 U15446 ( .A(n12428), .ZN(n12429) );
  NAND2_X1 U15447 ( .A1(n13474), .A2(n12429), .ZN(n12430) );
  NAND2_X1 U15448 ( .A1(n19954), .A2(n12430), .ZN(n19962) );
  INV_X1 U15449 ( .A(n19962), .ZN(n12431) );
  NAND2_X1 U15450 ( .A1(n12431), .A2(n19976), .ZN(n12432) );
  NOR2_X1 U15451 ( .A1(n12423), .A2(n12432), .ZN(n12815) );
  INV_X1 U15452 ( .A(n12815), .ZN(n12433) );
  OAI21_X1 U15453 ( .B1(n12435), .B2(n12434), .A(n12433), .ZN(n12436) );
  NOR2_X1 U15454 ( .A1(n12996), .A2(n12436), .ZN(n12445) );
  INV_X1 U15455 ( .A(n12437), .ZN(n12441) );
  INV_X1 U15456 ( .A(n12438), .ZN(n12440) );
  AOI21_X1 U15457 ( .B1(n12441), .B2(n12440), .A(n12439), .ZN(n12443) );
  OAI21_X1 U15458 ( .B1(n12444), .B2(n12443), .A(n12442), .ZN(n19965) );
  NAND4_X1 U15459 ( .A1(n12447), .A2(n12446), .A3(n12445), .A4(n12817), .ZN(
        n12449) );
  NAND2_X1 U15460 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13474), .ZN(n13475) );
  INV_X1 U15461 ( .A(n13475), .ZN(n12448) );
  NOR2_X1 U15462 ( .A1(n12423), .A2(n13489), .ZN(n19963) );
  NAND2_X1 U15463 ( .A1(n12819), .A2(n19263), .ZN(n12814) );
  AND2_X1 U15464 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12806) );
  NAND2_X1 U15465 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16223) );
  INV_X1 U15466 ( .A(n16223), .ZN(n12470) );
  INV_X1 U15467 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15289) );
  NOR3_X1 U15468 ( .A1(n13419), .A2(n15289), .A3(n19259), .ZN(n13724) );
  NAND2_X1 U15469 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13724), .ZN(
        n12475) );
  INV_X1 U15470 ( .A(n12450), .ZN(n12451) );
  NAND2_X1 U15471 ( .A1(n12452), .A2(n12451), .ZN(n16271) );
  INV_X1 U15472 ( .A(n16271), .ZN(n12453) );
  INV_X1 U15473 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13894) );
  NOR2_X1 U15474 ( .A1(n12056), .A2(n13894), .ZN(n13888) );
  NAND2_X1 U15475 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13888), .ZN(
        n13078) );
  NOR2_X1 U15476 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13888), .ZN(
        n13067) );
  AOI21_X1 U15477 ( .B1(n15202), .B2(n13078), .A(n13067), .ZN(n16241) );
  NAND2_X1 U15478 ( .A1(n12454), .A2(n19976), .ZN(n13571) );
  AOI21_X1 U15479 ( .B1(n13571), .B2(n12456), .A(n12455), .ZN(n12466) );
  AND2_X1 U15480 ( .A1(n19273), .A2(n16274), .ZN(n12464) );
  AND2_X1 U15481 ( .A1(n13048), .A2(n12458), .ZN(n12461) );
  NAND2_X1 U15482 ( .A1(n12459), .A2(n19984), .ZN(n12867) );
  NAND2_X1 U15483 ( .A1(n9817), .A2(n12023), .ZN(n12460) );
  AOI22_X1 U15484 ( .A1(n12462), .A2(n12461), .B1(n12867), .B2(n12460), .ZN(
        n12463) );
  OAI21_X1 U15485 ( .B1(n12457), .B2(n12464), .A(n12463), .ZN(n12465) );
  NOR2_X1 U15486 ( .A1(n9819), .A2(n13489), .ZN(n12467) );
  NAND2_X1 U15487 ( .A1(n12468), .A2(n12467), .ZN(n15307) );
  NAND2_X1 U15488 ( .A1(n16282), .A2(n15307), .ZN(n12469) );
  NAND2_X1 U15489 ( .A1(n12810), .A2(n12469), .ZN(n15204) );
  NAND2_X1 U15490 ( .A1(n16241), .A2(n16257), .ZN(n15288) );
  NAND2_X1 U15491 ( .A1(n12470), .A2(n16224), .ZN(n13935) );
  AND2_X1 U15492 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16196) );
  AND2_X1 U15493 ( .A1(n16196), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15191) );
  AND2_X1 U15494 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15257) );
  AND2_X1 U15495 ( .A1(n15257), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13923) );
  AND2_X1 U15496 ( .A1(n15191), .A2(n13923), .ZN(n15183) );
  AND2_X1 U15497 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15005) );
  NAND2_X1 U15498 ( .A1(n15005), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15192) );
  NOR2_X1 U15499 ( .A1(n15192), .A2(n15196), .ZN(n12471) );
  AND2_X1 U15500 ( .A1(n15183), .A2(n12471), .ZN(n12805) );
  INV_X1 U15501 ( .A(n12805), .ZN(n12477) );
  NAND2_X1 U15502 ( .A1(n12806), .A2(n15174), .ZN(n15589) );
  NOR2_X1 U15503 ( .A1(n15588), .A2(n15589), .ZN(n15138) );
  INV_X1 U15504 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15127) );
  NOR2_X1 U15505 ( .A1(n15127), .A2(n15141), .ZN(n15123) );
  NAND2_X1 U15506 ( .A1(n15138), .A2(n15123), .ZN(n15114) );
  INV_X1 U15507 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15115) );
  NOR2_X1 U15508 ( .A1(n15114), .A2(n15115), .ZN(n15103) );
  NAND2_X1 U15509 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15086) );
  INV_X1 U15510 ( .A(n15086), .ZN(n12479) );
  NAND2_X1 U15511 ( .A1(n15103), .A2(n12479), .ZN(n15074) );
  INV_X1 U15512 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12472) );
  INV_X1 U15513 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15081) );
  NOR2_X1 U15514 ( .A1(n12472), .A2(n15081), .ZN(n15064) );
  OR2_X1 U15515 ( .A1(n15204), .A2(n13888), .ZN(n12474) );
  INV_X1 U15516 ( .A(n12810), .ZN(n12473) );
  NOR2_X2 U15517 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19728) );
  AND2_X1 U15518 ( .A1(n19972), .A2(n19728), .ZN(n12763) );
  INV_X1 U15519 ( .A(n12763), .ZN(n16232) );
  NAND2_X1 U15520 ( .A1(n12473), .A2(n16232), .ZN(n16254) );
  NAND2_X1 U15521 ( .A1(n12474), .A2(n16254), .ZN(n13080) );
  NOR2_X1 U15522 ( .A1(n13080), .A2(n16257), .ZN(n15255) );
  INV_X1 U15523 ( .A(n15255), .ZN(n15185) );
  NOR3_X1 U15524 ( .A1(n13067), .A2(n12475), .A3(n16223), .ZN(n12476) );
  NOR2_X1 U15525 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15204), .ZN(
        n13083) );
  NOR2_X1 U15526 ( .A1(n13083), .A2(n13080), .ZN(n13721) );
  OAI21_X1 U15527 ( .B1(n15285), .B2(n12476), .A(n13721), .ZN(n15182) );
  OAI21_X1 U15528 ( .B1(n15182), .B2(n12477), .A(n15185), .ZN(n15176) );
  OAI211_X1 U15529 ( .C1(n12806), .C2(n15255), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n15176), .ZN(n15593) );
  NAND2_X1 U15530 ( .A1(n15185), .A2(n15593), .ZN(n15140) );
  OAI211_X1 U15531 ( .C1(n15123), .C2(n15285), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15140), .ZN(n12478) );
  INV_X1 U15532 ( .A(n12478), .ZN(n15113) );
  OR2_X1 U15533 ( .A1(n15255), .A2(n15113), .ZN(n15100) );
  OR2_X1 U15534 ( .A1(n15255), .A2(n12479), .ZN(n12480) );
  OAI21_X1 U15535 ( .B1(n15074), .B2(n15064), .A(n15079), .ZN(n15068) );
  OR2_X1 U15536 ( .A1(n13970), .A2(n15141), .ZN(n12486) );
  INV_X1 U15537 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12750) );
  NAND2_X1 U15538 ( .A1(n13966), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15539 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12482) );
  OAI211_X1 U15540 ( .C1(n13873), .C2(n12750), .A(n12483), .B(n12482), .ZN(
        n12484) );
  INV_X1 U15541 ( .A(n12484), .ZN(n12485) );
  NAND2_X1 U15542 ( .A1(n12486), .A2(n12485), .ZN(n15147) );
  OR2_X1 U15543 ( .A1(n13970), .A2(n19259), .ZN(n12490) );
  AOI22_X1 U15544 ( .A1(n13965), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12489) );
  OAI211_X1 U15545 ( .C1(n13870), .C2(n19120), .A(n12490), .B(n12489), .ZN(
        n19024) );
  NAND2_X1 U15546 ( .A1(n19025), .A2(n19024), .ZN(n13223) );
  INV_X1 U15547 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n15291) );
  OAI22_X1 U15548 ( .A1(n13873), .A2(n15291), .B1(n13474), .B2(n16178), .ZN(
        n12492) );
  NOR2_X1 U15549 ( .A1(n13970), .A2(n15289), .ZN(n12491) );
  AOI211_X1 U15550 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n13966), .A(n12492), .B(
        n12491), .ZN(n13224) );
  OR2_X1 U15551 ( .A1(n13970), .A2(n15272), .ZN(n12498) );
  INV_X1 U15552 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12495) );
  NAND2_X1 U15553 ( .A1(n13966), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U15554 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12493) );
  OAI211_X1 U15555 ( .C1(n13873), .C2(n12495), .A(n12494), .B(n12493), .ZN(
        n12496) );
  INV_X1 U15556 ( .A(n12496), .ZN(n12497) );
  NAND2_X1 U15557 ( .A1(n12498), .A2(n12497), .ZN(n13262) );
  INV_X1 U15558 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13277) );
  INV_X1 U15559 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16225) );
  OR2_X1 U15560 ( .A1(n13970), .A2(n16225), .ZN(n12500) );
  AOI22_X1 U15561 ( .A1(n13965), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12499) );
  OAI211_X1 U15562 ( .C1(n13277), .C2(n13870), .A(n12500), .B(n12499), .ZN(
        n13275) );
  INV_X1 U15563 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n19110) );
  OR2_X1 U15564 ( .A1(n13970), .A2(n16227), .ZN(n12502) );
  AOI22_X1 U15565 ( .A1(n13965), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12501) );
  OAI211_X1 U15566 ( .C1(n19110), .C2(n13870), .A(n12502), .B(n12501), .ZN(
        n16149) );
  INV_X1 U15567 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n12505) );
  OR2_X1 U15568 ( .A1(n13970), .A2(n13936), .ZN(n12504) );
  AOI22_X1 U15569 ( .A1(n13965), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12503) );
  OAI211_X1 U15570 ( .C1(n12505), .C2(n13870), .A(n12504), .B(n12503), .ZN(
        n13359) );
  INV_X1 U15571 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n12509) );
  OR2_X1 U15572 ( .A1(n13970), .A2(n12506), .ZN(n12508) );
  AOI22_X1 U15573 ( .A1(n13965), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12507) );
  OAI211_X1 U15574 ( .C1(n12509), .C2(n13870), .A(n12508), .B(n12507), .ZN(
        n16141) );
  OR2_X1 U15575 ( .A1(n13970), .A2(n15258), .ZN(n12511) );
  AOI22_X1 U15576 ( .A1(n13965), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n12510) );
  OAI211_X1 U15577 ( .C1(n13399), .C2(n13870), .A(n12511), .B(n12510), .ZN(
        n13395) );
  INV_X1 U15578 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n12515) );
  OR2_X1 U15579 ( .A1(n13970), .A2(n12512), .ZN(n12514) );
  AOI22_X1 U15580 ( .A1(n13965), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12513) );
  OAI211_X1 U15581 ( .C1(n12515), .C2(n13870), .A(n12514), .B(n12513), .ZN(
        n13915) );
  INV_X1 U15582 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n12518) );
  OR2_X1 U15583 ( .A1(n13970), .A2(n15242), .ZN(n12517) );
  AOI22_X1 U15584 ( .A1(n13965), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n12516) );
  OAI211_X1 U15585 ( .C1(n12518), .C2(n13870), .A(n12517), .B(n12516), .ZN(
        n13403) );
  OR2_X1 U15586 ( .A1(n13970), .A2(n16210), .ZN(n12520) );
  AOI22_X1 U15587 ( .A1(n13965), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n12519) );
  OAI211_X1 U15588 ( .C1(n12521), .C2(n13870), .A(n12520), .B(n12519), .ZN(
        n16104) );
  OR2_X1 U15589 ( .A1(n13970), .A2(n16187), .ZN(n12523) );
  AOI22_X1 U15590 ( .A1(n13965), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n12522) );
  OAI211_X1 U15591 ( .C1(n12524), .C2(n13870), .A(n12523), .B(n12522), .ZN(
        n13546) );
  OR2_X1 U15592 ( .A1(n13970), .A2(n15230), .ZN(n12529) );
  INV_X1 U15593 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19873) );
  NAND2_X1 U15594 ( .A1(n13966), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12526) );
  NAND2_X1 U15595 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12525) );
  OAI211_X1 U15596 ( .C1(n13873), .C2(n19873), .A(n12526), .B(n12525), .ZN(
        n12527) );
  INV_X1 U15597 ( .A(n12527), .ZN(n12528) );
  OR2_X1 U15598 ( .A1(n13970), .A2(n12530), .ZN(n12535) );
  INV_X1 U15599 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19875) );
  NAND2_X1 U15600 ( .A1(n13966), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n12532) );
  NAND2_X1 U15601 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12531) );
  OAI211_X1 U15602 ( .C1(n13873), .C2(n19875), .A(n12532), .B(n12531), .ZN(
        n12533) );
  INV_X1 U15603 ( .A(n12533), .ZN(n12534) );
  NAND2_X1 U15604 ( .A1(n12535), .A2(n12534), .ZN(n14803) );
  OR2_X1 U15605 ( .A1(n13970), .A2(n15196), .ZN(n12540) );
  INV_X1 U15606 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15010) );
  NAND2_X1 U15607 ( .A1(n13966), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12537) );
  NAND2_X1 U15608 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12536) );
  OAI211_X1 U15609 ( .C1(n13873), .C2(n15010), .A(n12537), .B(n12536), .ZN(
        n12538) );
  INV_X1 U15610 ( .A(n12538), .ZN(n12539) );
  OR2_X1 U15611 ( .A1(n13970), .A2(n15177), .ZN(n12545) );
  INV_X1 U15612 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19878) );
  NAND2_X1 U15613 ( .A1(n13966), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12542) );
  NAND2_X1 U15614 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12541) );
  OAI211_X1 U15615 ( .C1(n13873), .C2(n19878), .A(n12542), .B(n12541), .ZN(
        n12543) );
  INV_X1 U15616 ( .A(n12543), .ZN(n12544) );
  OR2_X1 U15617 ( .A1(n13970), .A2(n15164), .ZN(n12550) );
  INV_X1 U15618 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19880) );
  NAND2_X1 U15619 ( .A1(n13966), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12547) );
  NAND2_X1 U15620 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n12546) );
  OAI211_X1 U15621 ( .C1(n13873), .C2(n19880), .A(n12547), .B(n12546), .ZN(
        n12548) );
  INV_X1 U15622 ( .A(n12548), .ZN(n12549) );
  NAND2_X1 U15623 ( .A1(n12550), .A2(n12549), .ZN(n14982) );
  OR2_X1 U15624 ( .A1(n13970), .A2(n15588), .ZN(n12555) );
  NAND2_X1 U15625 ( .A1(n13966), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12552) );
  NAND2_X1 U15626 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12551) );
  OAI211_X1 U15627 ( .C1(n13873), .C2(n19882), .A(n12552), .B(n12551), .ZN(
        n12553) );
  INV_X1 U15628 ( .A(n12553), .ZN(n12554) );
  INV_X1 U15629 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n12558) );
  OR2_X1 U15630 ( .A1(n13970), .A2(n15127), .ZN(n12557) );
  AOI22_X1 U15631 ( .A1(n13965), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n12556) );
  OAI211_X1 U15632 ( .C1(n13870), .C2(n12558), .A(n12557), .B(n12556), .ZN(
        n14946) );
  INV_X1 U15633 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U15634 ( .A1(n13966), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U15635 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12559) );
  OAI211_X1 U15636 ( .C1(n13873), .C2(n12755), .A(n12560), .B(n12559), .ZN(
        n12561) );
  AOI21_X1 U15637 ( .B1(n13875), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n12561), .ZN(n14784) );
  OR2_X1 U15638 ( .A1(n13970), .A2(n15102), .ZN(n12563) );
  AOI22_X1 U15639 ( .A1(n13965), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n12562) );
  OAI211_X1 U15640 ( .C1(n13870), .C2(n14778), .A(n12563), .B(n12562), .ZN(
        n14777) );
  NAND2_X1 U15641 ( .A1(n14785), .A2(n14777), .ZN(n14776) );
  INV_X1 U15642 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19890) );
  NAND2_X1 U15643 ( .A1(n13966), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12565) );
  NAND2_X1 U15644 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12564) );
  OAI211_X1 U15645 ( .C1(n13873), .C2(n19890), .A(n12565), .B(n12564), .ZN(
        n12566) );
  AOI21_X1 U15646 ( .B1(n13875), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n12566), .ZN(n14765) );
  INV_X1 U15647 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19894) );
  NAND2_X1 U15648 ( .A1(n13966), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12568) );
  NAND2_X1 U15649 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12567) );
  OAI211_X1 U15650 ( .C1(n13873), .C2(n19894), .A(n12568), .B(n12567), .ZN(
        n12569) );
  AOI21_X1 U15651 ( .B1(n13875), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n12569), .ZN(n14760) );
  INV_X1 U15652 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U15653 ( .A1(n13966), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12571) );
  NAND2_X1 U15654 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12570) );
  OAI211_X1 U15655 ( .C1(n13873), .C2(n12764), .A(n12571), .B(n12570), .ZN(
        n12572) );
  AOI21_X1 U15656 ( .B1(n13875), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12572), .ZN(n12573) );
  AND2_X1 U15657 ( .A1(n14762), .A2(n12573), .ZN(n12574) );
  OR2_X1 U15658 ( .A1(n12574), .A2(n14744), .ZN(n16004) );
  NAND2_X1 U15659 ( .A1(n12810), .A2(n12575), .ZN(n16253) );
  NAND2_X1 U15660 ( .A1(n19273), .A2(n19976), .ZN(n12577) );
  NOR2_X1 U15661 ( .A1(n12576), .A2(n12577), .ZN(n16269) );
  NOR2_X1 U15662 ( .A1(n16266), .A2(n12584), .ZN(n12579) );
  OR2_X1 U15663 ( .A1(n16269), .A2(n12579), .ZN(n12580) );
  INV_X2 U15664 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19971) );
  NOR2_X1 U15665 ( .A1(n15344), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15666 ( .A1(n13988), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12585) );
  OAI21_X1 U15667 ( .B1(n12759), .B2(n12764), .A(n12585), .ZN(n12586) );
  INV_X1 U15668 ( .A(n12586), .ZN(n12762) );
  INV_X1 U15669 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19066) );
  INV_X1 U15670 ( .A(n12587), .ZN(n12589) );
  NAND2_X1 U15671 ( .A1(n13064), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12588) );
  OAI211_X1 U15672 ( .C1(n12759), .C2(n19066), .A(n12589), .B(n12588), .ZN(
        n13056) );
  NAND2_X1 U15673 ( .A1(n12594), .A2(n13062), .ZN(n12604) );
  OAI22_X1 U15674 ( .A1(n15344), .A2(P2_STATE2_REG_3__SCAN_IN), .B1(n19958), 
        .B2(n19971), .ZN(n12590) );
  INV_X1 U15675 ( .A(n12590), .ZN(n12591) );
  AND2_X1 U15676 ( .A1(n12604), .A2(n12591), .ZN(n12593) );
  NAND2_X1 U15677 ( .A1(n10206), .A2(n9873), .ZN(n12597) );
  OR2_X1 U15678 ( .A1(n12770), .A2(n12597), .ZN(n12592) );
  NAND2_X1 U15679 ( .A1(n12593), .A2(n12592), .ZN(n13055) );
  AND2_X2 U15680 ( .A1(n13056), .A2(n13055), .ZN(n13054) );
  AOI22_X1 U15681 ( .A1(n12609), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12595) );
  OAI21_X1 U15682 ( .B1(n12759), .B2(n12061), .A(n12595), .ZN(n12602) );
  INV_X1 U15683 ( .A(n12602), .ZN(n12596) );
  OR2_X1 U15684 ( .A1(n12769), .A2(n12597), .ZN(n12601) );
  NAND2_X1 U15685 ( .A1(n15344), .A2(n19971), .ZN(n12598) );
  OAI22_X1 U15686 ( .A1(n13062), .A2(n12598), .B1(n19971), .B2(n19949), .ZN(
        n12599) );
  INV_X1 U15687 ( .A(n12599), .ZN(n12600) );
  AND2_X1 U15688 ( .A1(n12601), .A2(n12600), .ZN(n13287) );
  NAND2_X1 U15689 ( .A1(n13288), .A2(n13287), .ZN(n13286) );
  OR2_X1 U15690 ( .A1(n13054), .A2(n12602), .ZN(n12607) );
  INV_X1 U15691 ( .A(n12603), .ZN(n12775) );
  OR2_X1 U15692 ( .A1(n12597), .A2(n12775), .ZN(n12605) );
  OAI211_X1 U15693 ( .C1(n19971), .C2(n13030), .A(n12605), .B(n12604), .ZN(
        n12606) );
  AND3_X1 U15694 ( .A1(n13286), .A2(n12607), .A3(n12606), .ZN(n12608) );
  AOI21_X2 U15695 ( .B1(n13286), .B2(n12607), .A(n12606), .ZN(n12611) );
  AOI22_X1 U15696 ( .A1(n13988), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12610) );
  OAI21_X1 U15697 ( .B1(n12759), .B2(n12075), .A(n12610), .ZN(n13072) );
  NOR2_X1 U15698 ( .A1(n13073), .A2(n13072), .ZN(n13074) );
  NOR2_X2 U15699 ( .A1(n13074), .A2(n12611), .ZN(n13501) );
  NAND2_X1 U15700 ( .A1(n13989), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12617) );
  AOI22_X1 U15701 ( .A1(n12594), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12616) );
  INV_X1 U15702 ( .A(n12612), .ZN(n12613) );
  OR2_X1 U15703 ( .A1(n12597), .A2(n12613), .ZN(n12615) );
  NAND2_X1 U15704 ( .A1(n13988), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12614) );
  NAND4_X1 U15705 ( .A1(n12617), .A2(n12616), .A3(n12615), .A4(n12614), .ZN(
        n13502) );
  INV_X1 U15706 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15707 ( .A1(n13988), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12620) );
  INV_X1 U15708 ( .A(n12781), .ZN(n12618) );
  OR2_X1 U15709 ( .A1(n12597), .A2(n12618), .ZN(n12619) );
  OAI211_X1 U15710 ( .C1(n12759), .C2(n12621), .A(n12620), .B(n12619), .ZN(
        n12622) );
  INV_X1 U15711 ( .A(n12622), .ZN(n19032) );
  AOI22_X1 U15712 ( .A1(n13988), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12625) );
  OR2_X1 U15713 ( .A1(n12597), .A2(n12623), .ZN(n12624) );
  OAI211_X1 U15714 ( .C1(n12759), .C2(n15291), .A(n12625), .B(n12624), .ZN(
        n15287) );
  AOI22_X1 U15715 ( .A1(n13988), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12627) );
  OAI21_X1 U15716 ( .B1(n12759), .B2(n12495), .A(n12627), .ZN(n13719) );
  NAND2_X1 U15717 ( .A1(n13720), .A2(n13719), .ZN(n12629) );
  OR2_X1 U15718 ( .A1(n12597), .A2(n13861), .ZN(n12628) );
  INV_X1 U15719 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19862) );
  AOI22_X1 U15720 ( .A1(n13988), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n12630) );
  OAI21_X1 U15721 ( .B1(n12759), .B2(n19862), .A(n12630), .ZN(n15273) );
  INV_X1 U15722 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12644) );
  AOI22_X1 U15723 ( .A1(n13988), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12643) );
  AOI22_X1 U15724 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15725 ( .A1(n12149), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12633) );
  AOI22_X1 U15726 ( .A1(n14001), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12632) );
  AOI22_X1 U15727 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12631) );
  NAND4_X1 U15728 ( .A1(n12634), .A2(n12633), .A3(n12632), .A4(n12631), .ZN(
        n12640) );
  AOI22_X1 U15729 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12638) );
  AOI22_X1 U15730 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12637) );
  AOI22_X1 U15731 ( .A1(n11863), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11912), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12636) );
  AOI22_X1 U15732 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12635) );
  NAND4_X1 U15733 ( .A1(n12638), .A2(n12637), .A3(n12636), .A4(n12635), .ZN(
        n12639) );
  INV_X1 U15734 ( .A(n19108), .ZN(n12641) );
  OR2_X1 U15735 ( .A1(n12597), .A2(n12641), .ZN(n12642) );
  OAI211_X1 U15736 ( .C1(n12759), .C2(n12644), .A(n12643), .B(n12642), .ZN(
        n12645) );
  INV_X1 U15737 ( .A(n12645), .ZN(n16230) );
  AOI22_X1 U15738 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12649) );
  AOI22_X1 U15739 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9814), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15740 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12726), .B1(
        n14001), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15741 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12646) );
  NAND4_X1 U15742 ( .A1(n12649), .A2(n12648), .A3(n12647), .A4(n12646), .ZN(
        n12655) );
  AOI22_X1 U15743 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15744 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12652) );
  AOI22_X1 U15745 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12651) );
  AOI22_X1 U15746 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12650) );
  NAND4_X1 U15747 ( .A1(n12653), .A2(n12652), .A3(n12651), .A4(n12650), .ZN(
        n12654) );
  INV_X1 U15748 ( .A(n13355), .ZN(n12658) );
  NAND2_X1 U15749 ( .A1(n13989), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12657) );
  AOI22_X1 U15750 ( .A1(n13988), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12594), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12656) );
  OAI211_X1 U15751 ( .C1(n12658), .C2(n12597), .A(n12657), .B(n12656), .ZN(
        n13934) );
  INV_X1 U15752 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12671) );
  AOI22_X1 U15753 ( .A1(n13988), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12670) );
  AOI22_X1 U15754 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11896), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15755 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12149), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15756 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12726), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15757 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n14079), .B1(
        n14001), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12659) );
  NAND4_X1 U15758 ( .A1(n12662), .A2(n12661), .A3(n12660), .A4(n12659), .ZN(
        n12668) );
  AOI22_X1 U15759 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12666) );
  AOI22_X1 U15760 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15761 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15762 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12663) );
  NAND4_X1 U15763 ( .A1(n12666), .A2(n12665), .A3(n12664), .A4(n12663), .ZN(
        n12667) );
  OR2_X1 U15764 ( .A1(n12668), .A2(n12667), .ZN(n19102) );
  INV_X1 U15765 ( .A(n19102), .ZN(n13387) );
  OR2_X1 U15766 ( .A1(n12597), .A2(n13387), .ZN(n12669) );
  OAI211_X1 U15767 ( .C1(n12759), .C2(n12671), .A(n12670), .B(n12669), .ZN(
        n16213) );
  INV_X1 U15768 ( .A(n16213), .ZN(n12672) );
  INV_X1 U15769 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15770 ( .A1(n13988), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15771 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12676) );
  AOI22_X1 U15772 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n9814), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U15773 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12726), .B1(
        n14001), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15774 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12673) );
  NAND4_X1 U15775 ( .A1(n12676), .A2(n12675), .A3(n12674), .A4(n12673), .ZN(
        n12682) );
  AOI22_X1 U15776 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12680) );
  AOI22_X1 U15777 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12679) );
  AOI22_X1 U15778 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12678) );
  AOI22_X1 U15779 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12677) );
  NAND4_X1 U15780 ( .A1(n12680), .A2(n12679), .A3(n12678), .A4(n12677), .ZN(
        n12681) );
  OR2_X1 U15781 ( .A1(n12682), .A2(n12681), .ZN(n13388) );
  INV_X1 U15782 ( .A(n13388), .ZN(n13386) );
  OR2_X1 U15783 ( .A1(n12597), .A2(n13386), .ZN(n12683) );
  OAI211_X1 U15784 ( .C1(n12759), .C2(n12685), .A(n12684), .B(n12683), .ZN(
        n15262) );
  NAND2_X1 U15785 ( .A1(n15261), .A2(n15262), .ZN(n13919) );
  INV_X1 U15786 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U15787 ( .A1(n13988), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12697) );
  AOI22_X1 U15788 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12149), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12689) );
  AOI22_X1 U15789 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11896), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U15790 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12726), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12687) );
  AOI22_X1 U15791 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n14079), .B1(
        n14001), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12686) );
  NAND4_X1 U15792 ( .A1(n12689), .A2(n12688), .A3(n12687), .A4(n12686), .ZN(
        n12695) );
  AOI22_X1 U15793 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U15794 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15795 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11912), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12691) );
  AOI22_X1 U15796 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12147), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12690) );
  NAND4_X1 U15797 ( .A1(n12693), .A2(n12692), .A3(n12691), .A4(n12690), .ZN(
        n12694) );
  NOR2_X1 U15798 ( .A1(n12695), .A2(n12694), .ZN(n19098) );
  OR2_X1 U15799 ( .A1(n12597), .A2(n19098), .ZN(n12696) );
  OAI211_X1 U15800 ( .C1(n12759), .C2(n12698), .A(n12697), .B(n12696), .ZN(
        n12699) );
  INV_X1 U15801 ( .A(n12699), .ZN(n13920) );
  NOR2_X2 U15802 ( .A1(n13919), .A2(n13920), .ZN(n15237) );
  INV_X1 U15803 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15804 ( .A1(n13988), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15805 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12149), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12703) );
  AOI22_X1 U15806 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12702) );
  AOI22_X1 U15807 ( .A1(n14001), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12701) );
  AOI22_X1 U15808 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12700) );
  NAND4_X1 U15809 ( .A1(n12703), .A2(n12702), .A3(n12701), .A4(n12700), .ZN(
        n12709) );
  AOI22_X1 U15810 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12155), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12707) );
  AOI22_X1 U15811 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12706) );
  AOI22_X1 U15812 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15813 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12704) );
  NAND4_X1 U15814 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n12704), .ZN(
        n12708) );
  OR2_X1 U15815 ( .A1(n12709), .A2(n12708), .ZN(n13401) );
  INV_X1 U15816 ( .A(n13401), .ZN(n13400) );
  OR2_X1 U15817 ( .A1(n12597), .A2(n13400), .ZN(n12710) );
  OAI211_X1 U15818 ( .C1(n12759), .C2(n12712), .A(n12711), .B(n12710), .ZN(
        n15238) );
  INV_X1 U15819 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12725) );
  AOI22_X1 U15820 ( .A1(n13988), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15821 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11896), .B1(
        n9814), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15822 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12149), .B1(
        n9815), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12715) );
  AOI22_X1 U15823 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12726), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U15824 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n14079), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12713) );
  NAND4_X1 U15825 ( .A1(n12716), .A2(n12715), .A3(n12714), .A4(n12713), .ZN(
        n12722) );
  AOI22_X1 U15826 ( .A1(n12155), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12154), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12720) );
  AOI22_X1 U15827 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12719) );
  AOI22_X1 U15828 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n11912), .B1(
        n11881), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15829 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12147), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12717) );
  NAND4_X1 U15830 ( .A1(n12720), .A2(n12719), .A3(n12718), .A4(n12717), .ZN(
        n12721) );
  NOR2_X1 U15831 ( .A1(n12722), .A2(n12721), .ZN(n19093) );
  OR2_X1 U15832 ( .A1(n12597), .A2(n19093), .ZN(n12723) );
  OAI211_X1 U15833 ( .C1(n12759), .C2(n12725), .A(n12724), .B(n12723), .ZN(
        n16197) );
  INV_X1 U15834 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U15835 ( .A1(n13988), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12738) );
  AOI22_X1 U15836 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15837 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n9814), .B1(
        n9816), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15838 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15839 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U15840 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12736) );
  AOI22_X1 U15841 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12734) );
  AOI22_X1 U15842 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15843 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U15844 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12731) );
  NAND4_X1 U15845 ( .A1(n12734), .A2(n12733), .A3(n12732), .A4(n12731), .ZN(
        n12735) );
  INV_X1 U15846 ( .A(n13545), .ZN(n13543) );
  OR2_X1 U15847 ( .A1(n12597), .A2(n13543), .ZN(n12737) );
  OAI211_X1 U15848 ( .C1(n12759), .C2(n12739), .A(n12738), .B(n12737), .ZN(
        n16181) );
  AOI22_X1 U15849 ( .A1(n13988), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12740) );
  OAI21_X1 U15850 ( .B1(n12759), .B2(n19873), .A(n12740), .ZN(n15220) );
  AOI22_X1 U15851 ( .A1(n13988), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12741) );
  OAI21_X1 U15852 ( .B1(n12759), .B2(n19875), .A(n12741), .ZN(n12742) );
  INV_X1 U15853 ( .A(n12742), .ZN(n13680) );
  AOI22_X1 U15854 ( .A1(n13988), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12743) );
  OAI21_X1 U15855 ( .B1(n12759), .B2(n15010), .A(n12743), .ZN(n15187) );
  NAND2_X1 U15856 ( .A1(n13679), .A2(n15187), .ZN(n15186) );
  AOI22_X1 U15857 ( .A1(n13988), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12744) );
  OAI21_X1 U15858 ( .B1(n12759), .B2(n19878), .A(n12744), .ZN(n12745) );
  INV_X1 U15859 ( .A(n12745), .ZN(n14881) );
  AOI22_X1 U15860 ( .A1(n13988), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12746) );
  OAI21_X1 U15861 ( .B1(n12759), .B2(n19880), .A(n12746), .ZN(n12747) );
  INV_X1 U15862 ( .A(n12747), .ZN(n15157) );
  INV_X1 U15863 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19882) );
  AOI22_X1 U15864 ( .A1(n13988), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12748) );
  OAI21_X1 U15865 ( .B1(n12759), .B2(n19882), .A(n12748), .ZN(n14872) );
  AOI22_X1 U15866 ( .A1(n13988), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12749) );
  OAI21_X1 U15867 ( .B1(n12759), .B2(n12750), .A(n12749), .ZN(n15143) );
  NAND2_X1 U15868 ( .A1(n12751), .A2(n15143), .ZN(n14861) );
  INV_X1 U15869 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19885) );
  AOI22_X1 U15870 ( .A1(n13988), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12752) );
  OAI21_X1 U15871 ( .B1(n12759), .B2(n19885), .A(n12752), .ZN(n12753) );
  INV_X1 U15872 ( .A(n12753), .ZN(n14862) );
  OR2_X2 U15873 ( .A1(n14861), .A2(n14862), .ZN(n14864) );
  AOI22_X1 U15874 ( .A1(n13988), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12754) );
  OAI21_X1 U15875 ( .B1(n12759), .B2(n12755), .A(n12754), .ZN(n12756) );
  INV_X1 U15876 ( .A(n12756), .ZN(n14851) );
  INV_X1 U15877 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19888) );
  AOI22_X1 U15878 ( .A1(n13988), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12757) );
  OAI21_X1 U15879 ( .B1(n12759), .B2(n19888), .A(n12757), .ZN(n14840) );
  AOI22_X1 U15880 ( .A1(n13988), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12758) );
  OAI21_X1 U15881 ( .B1(n12759), .B2(n19890), .A(n12758), .ZN(n14834) );
  AOI22_X1 U15882 ( .A1(n13988), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12760) );
  OAI21_X1 U15883 ( .B1(n12759), .B2(n19894), .A(n12760), .ZN(n12761) );
  INV_X1 U15884 ( .A(n12761), .ZN(n14825) );
  AOI21_X1 U15885 ( .B1(n12762), .B2(n9835), .A(n14812), .ZN(n16002) );
  NOR2_X1 U15886 ( .A1(n16232), .A2(n12764), .ZN(n12826) );
  AOI21_X1 U15887 ( .B1(n19257), .B2(n16002), .A(n12826), .ZN(n12765) );
  OAI21_X1 U15888 ( .B1(n16004), .B2(n16253), .A(n12765), .ZN(n12767) );
  NOR3_X1 U15889 ( .A1(n15074), .A2(n15064), .A3(n15081), .ZN(n12766) );
  AOI211_X1 U15890 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15068), .A(
        n12767), .B(n12766), .ZN(n12812) );
  NAND2_X1 U15891 ( .A1(n12953), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12952) );
  INV_X1 U15892 ( .A(n12952), .ZN(n12771) );
  XOR2_X1 U15893 ( .A(n12770), .B(n12769), .Z(n12772) );
  NAND2_X1 U15894 ( .A1(n12771), .A2(n12772), .ZN(n12773) );
  XNOR2_X1 U15895 ( .A(n12772), .B(n12952), .ZN(n13896) );
  NAND2_X1 U15896 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13896), .ZN(
        n13895) );
  NAND2_X1 U15897 ( .A1(n12773), .A2(n13895), .ZN(n12776) );
  XOR2_X1 U15898 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12776), .Z(
        n13082) );
  XOR2_X1 U15899 ( .A(n12775), .B(n12774), .Z(n13081) );
  NAND2_X1 U15900 ( .A1(n13082), .A2(n13081), .ZN(n12778) );
  NAND2_X1 U15901 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12776), .ZN(
        n12777) );
  NAND2_X1 U15902 ( .A1(n12778), .A2(n12777), .ZN(n12779) );
  XNOR2_X1 U15903 ( .A(n12779), .B(n13419), .ZN(n13423) );
  NAND2_X1 U15904 ( .A1(n12779), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12780) );
  NAND2_X1 U15905 ( .A1(n19233), .A2(n19259), .ZN(n12786) );
  INV_X1 U15906 ( .A(n12782), .ZN(n12785) );
  INV_X1 U15907 ( .A(n12783), .ZN(n12784) );
  NAND2_X1 U15908 ( .A1(n12785), .A2(n12784), .ZN(n19234) );
  INV_X1 U15909 ( .A(n12789), .ZN(n12788) );
  NAND2_X1 U15910 ( .A1(n12788), .A2(n15289), .ZN(n15297) );
  NAND3_X1 U15911 ( .A1(n15295), .A2(n15298), .A3(n12792), .ZN(n12791) );
  INV_X1 U15912 ( .A(n15298), .ZN(n15294) );
  NAND2_X1 U15913 ( .A1(n15295), .A2(n15298), .ZN(n12793) );
  NAND2_X1 U15914 ( .A1(n12793), .A2(n12792), .ZN(n12794) );
  NAND2_X1 U15915 ( .A1(n12795), .A2(n13861), .ZN(n12797) );
  NAND2_X1 U15916 ( .A1(n12802), .A2(n12797), .ZN(n12798) );
  NAND2_X1 U15917 ( .A1(n15055), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15269) );
  INV_X1 U15918 ( .A(n12798), .ZN(n12799) );
  NAND2_X1 U15919 ( .A1(n12800), .A2(n12799), .ZN(n12801) );
  INV_X1 U15920 ( .A(n12802), .ZN(n12803) );
  NAND2_X1 U15921 ( .A1(n12803), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12804) );
  INV_X1 U15922 ( .A(n12806), .ZN(n15161) );
  OAI21_X1 U15923 ( .B1(n14914), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14909), .ZN(n12821) );
  INV_X1 U15924 ( .A(n12809), .ZN(n19964) );
  OR2_X1 U15925 ( .A1(n12821), .A2(n16264), .ZN(n12811) );
  NAND2_X1 U15926 ( .A1(n12814), .A2(n12813), .ZN(P2_U3018) );
  NAND2_X1 U15927 ( .A1(n12815), .A2(n16274), .ZN(n12816) );
  NAND2_X1 U15928 ( .A1(n12817), .A2(n12816), .ZN(n12818) );
  NAND2_X1 U15929 ( .A1(n12819), .A2(n19240), .ZN(n12832) );
  INV_X1 U15930 ( .A(n12869), .ZN(n12820) );
  NAND2_X1 U15931 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n15487), .ZN(
        n15486) );
  INV_X1 U15932 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18930) );
  INV_X1 U15933 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15045) );
  INV_X1 U15934 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14996) );
  INV_X1 U15935 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14969) );
  INV_X1 U15936 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16028) );
  OAI21_X1 U15937 ( .B1(n14919), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14905), .ZN(n15965) );
  INV_X1 U15938 ( .A(n15965), .ZN(n15996) );
  NOR2_X1 U15939 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19831) );
  OR2_X1 U15940 ( .A1(n19728), .A2(n19831), .ZN(n19950) );
  NAND2_X1 U15941 ( .A1(n19950), .A2(n13470), .ZN(n12822) );
  INV_X1 U15942 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19920) );
  NAND2_X1 U15943 ( .A1(n19920), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12823) );
  NAND2_X1 U15944 ( .A1(n10105), .A2(n12823), .ZN(n12954) );
  AOI21_X1 U15945 ( .B1(n19979), .B2(n13474), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19982) );
  NAND2_X1 U15946 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13005) );
  AND2_X1 U15947 ( .A1(n19982), .A2(n13005), .ZN(n12824) );
  INV_X1 U15948 ( .A(n15339), .ZN(n19250) );
  AOI21_X1 U15949 ( .B1(n19239), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12826), .ZN(n12827) );
  OAI21_X1 U15950 ( .B1(n16004), .B2(n15339), .A(n12827), .ZN(n12828) );
  AOI21_X1 U15951 ( .B1(n15996), .B2(n16170), .A(n12828), .ZN(n12829) );
  NAND2_X1 U15952 ( .A1(n12832), .A2(n12831), .ZN(P2_U2986) );
  NAND2_X1 U15953 ( .A1(n12834), .A2(n17739), .ZN(n12846) );
  OR2_X1 U15954 ( .A1(n12835), .A2(n17737), .ZN(n12844) );
  NAND2_X1 U15955 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17791) );
  OAI21_X1 U15956 ( .B1(n18813), .B2(n18812), .A(n18758), .ZN(n18803) );
  NAND2_X1 U15957 ( .A1(n17792), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17777) );
  NAND2_X1 U15958 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17740) );
  NOR2_X1 U15959 ( .A1(n17740), .A2(n17719), .ZN(n17692) );
  NAND3_X1 U15960 ( .A1(n17692), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16690) );
  NAND2_X1 U15961 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17623) );
  NAND2_X1 U15962 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17591) );
  NAND2_X1 U15963 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17560) );
  NAND2_X1 U15964 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17549), .ZN(
        n17508) );
  NAND2_X1 U15965 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17509) );
  NAND2_X1 U15966 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17496), .ZN(
        n17476) );
  NAND2_X1 U15967 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17477) );
  INV_X1 U15968 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17825) );
  NOR2_X1 U15969 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18812), .ZN(n17507) );
  NOR2_X1 U15970 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18758), .ZN(
        n18783) );
  AOI22_X1 U15971 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .B1(n18812), .B2(n18813), .ZN(n18656) );
  NOR2_X1 U15972 ( .A1(n18783), .A2(n18656), .ZN(n18156) );
  INV_X1 U15973 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18807) );
  NOR3_X1 U15974 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .A3(n18807), .ZN(n18448) );
  NAND2_X1 U15975 ( .A1(n18452), .A2(n18448), .ZN(n18498) );
  OAI21_X1 U15976 ( .B1(n17608), .B2(n17825), .A(n18498), .ZN(n17663) );
  NAND2_X1 U15977 ( .A1(n9916), .A2(n17663), .ZN(n16332) );
  XOR2_X1 U15978 ( .A(n10052), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(
        n12837) );
  NOR2_X1 U15979 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17608), .ZN(
        n16347) );
  INV_X1 U15980 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17489) );
  INV_X1 U15981 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16564) );
  NOR2_X1 U15982 ( .A1(n17825), .A2(n17508), .ZN(n16500) );
  NAND3_X1 U15983 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A3(n16500), .ZN(n17467) );
  NOR2_X1 U15984 ( .A1(n16564), .A2(n17467), .ZN(n16497) );
  INV_X1 U15985 ( .A(n16497), .ZN(n16496) );
  NOR2_X1 U15986 ( .A1(n17489), .A2(n16496), .ZN(n16495) );
  NAND2_X1 U15987 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16495), .ZN(
        n16493) );
  INV_X1 U15988 ( .A(n17830), .ZN(n17801) );
  NOR2_X1 U15989 ( .A1(n18498), .A2(n9916), .ZN(n16338) );
  AOI211_X1 U15990 ( .C1(n16493), .C2(n17507), .A(n17801), .B(n16338), .ZN(
        n12836) );
  INV_X1 U15991 ( .A(n12836), .ZN(n16337) );
  NOR2_X1 U15992 ( .A1(n16347), .A2(n16337), .ZN(n16331) );
  OAI22_X1 U15993 ( .A1(n16332), .A2(n12837), .B1(n16331), .B2(n10052), .ZN(
        n12838) );
  AOI211_X1 U15994 ( .C1(n17685), .C2(n16818), .A(n12839), .B(n12838), .ZN(
        n12842) );
  NOR2_X2 U15995 ( .A1(n18164), .A2(n16474), .ZN(n17818) );
  AND2_X1 U15996 ( .A1(n12842), .A2(n12841), .ZN(n12843) );
  AND2_X1 U15997 ( .A1(n12844), .A2(n12843), .ZN(n12845) );
  NAND2_X1 U15998 ( .A1(n12846), .A2(n12845), .ZN(P3_U2799) );
  NOR2_X1 U15999 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12848) );
  NOR4_X1 U16000 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12847) );
  NAND4_X1 U16001 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12848), .A4(n12847), .ZN(n12861) );
  NOR2_X1 U16002 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12861), .ZN(n16460)
         );
  INV_X1 U16003 ( .A(P1_M_IO_N_REG_SCAN_IN), .ZN(n20947) );
  INV_X1 U16004 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20968) );
  NOR4_X1 U16005 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        n20947), .A4(n20968), .ZN(n12850) );
  NOR4_X1 U16006 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n12849)
         );
  NAND3_X1 U16007 ( .A1(n13593), .A2(n12850), .A3(n12849), .ZN(U214) );
  NOR4_X1 U16008 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12854) );
  NOR4_X1 U16009 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12853) );
  NOR4_X1 U16010 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12852) );
  NOR4_X1 U16011 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12851) );
  NAND4_X1 U16012 ( .A1(n12854), .A2(n12853), .A3(n12852), .A4(n12851), .ZN(
        n12859) );
  NOR4_X1 U16013 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12857) );
  NOR4_X1 U16014 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n12856) );
  NOR4_X1 U16015 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12855) );
  INV_X1 U16016 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19858) );
  NAND4_X1 U16017 ( .A1(n12857), .A2(n12856), .A3(n12855), .A4(n19858), .ZN(
        n12858) );
  OAI21_X1 U16018 ( .B1(n12859), .B2(n12858), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12860) );
  INV_X2 U16019 ( .A(n15340), .ZN(n15338) );
  NOR2_X1 U16020 ( .A1(n15338), .A2(n12861), .ZN(n16374) );
  NAND2_X1 U16021 ( .A1(n16374), .A2(U214), .ZN(U212) );
  INV_X1 U16022 ( .A(n19829), .ZN(n13007) );
  NOR2_X1 U16023 ( .A1(n12863), .A2(n13011), .ZN(n19077) );
  INV_X1 U16024 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12865) );
  INV_X1 U16025 ( .A(n13480), .ZN(n12870) );
  AND2_X1 U16026 ( .A1(n19728), .A2(n13474), .ZN(n18826) );
  INV_X1 U16027 ( .A(n18826), .ZN(n12864) );
  OAI211_X1 U16028 ( .C1(n19077), .C2(n12865), .A(n12870), .B(n12864), .ZN(
        P2_U2814) );
  NOR2_X1 U16029 ( .A1(n16266), .A2(n16267), .ZN(n12999) );
  NAND2_X1 U16030 ( .A1(n12999), .A2(n19829), .ZN(n19974) );
  OAI21_X1 U16031 ( .B1(P2_READREQUEST_REG_SCAN_IN), .B2(n18826), .A(n19974), 
        .ZN(n12866) );
  OAI21_X1 U16032 ( .B1(n19974), .B2(n12867), .A(n12866), .ZN(P2_U3612) );
  INV_X1 U16033 ( .A(n12999), .ZN(n12868) );
  NOR2_X1 U16034 ( .A1(n12867), .A2(n19980), .ZN(n12998) );
  NOR3_X1 U16035 ( .A1(n12868), .A2(n12998), .A3(n12994), .ZN(n16306) );
  NOR2_X1 U16036 ( .A1(n16306), .A2(n13007), .ZN(n19961) );
  OAI21_X1 U16037 ( .B1(n19961), .B2(n13006), .A(n12869), .ZN(P2_U2819) );
  INV_X1 U16038 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12872) );
  INV_X1 U16039 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12871) );
  AOI21_X1 U16040 ( .B1(n19976), .B2(n19980), .A(n12870), .ZN(n12876) );
  NAND3_X1 U16041 ( .A1(n13480), .A2(n19976), .A3(n19838), .ZN(n12910) );
  AOI22_X1 U16042 ( .A1(n15340), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15338), .ZN(n19136) );
  OAI222_X1 U16043 ( .A1(n12975), .A2(n12872), .B1(n12871), .B2(n12876), .C1(
        n12910), .C2(n19136), .ZN(P2_U2982) );
  INV_X1 U16044 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12874) );
  INV_X1 U16045 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12873) );
  INV_X1 U16046 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16427) );
  INV_X1 U16047 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18158) );
  AOI22_X1 U16048 ( .A1(n15340), .A2(n16427), .B1(n18158), .B2(n15338), .ZN(
        n19124) );
  INV_X1 U16049 ( .A(n19124), .ZN(n15328) );
  OAI222_X1 U16050 ( .A1(n12975), .A2(n12874), .B1(n12873), .B2(n12876), .C1(
        n12910), .C2(n15328), .ZN(P2_U2967) );
  INV_X1 U16051 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13121) );
  INV_X1 U16052 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n12875) );
  OAI222_X1 U16053 ( .A1(n12910), .A2(n15328), .B1(n12975), .B2(n13121), .C1(
        n12875), .C2(n12876), .ZN(P2_U2952) );
  INV_X1 U16054 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13119) );
  INV_X2 U16055 ( .A(n12876), .ZN(n12940) );
  NAND2_X1 U16056 ( .A1(n12940), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12879) );
  NAND2_X1 U16057 ( .A1(n15338), .A2(BUF2_REG_10__SCAN_IN), .ZN(n12878) );
  INV_X1 U16058 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16405) );
  OR2_X1 U16059 ( .A1(n15338), .A2(n16405), .ZN(n12877) );
  NAND2_X1 U16060 ( .A1(n12878), .A2(n12877), .ZN(n19150) );
  NAND2_X1 U16061 ( .A1(n12930), .A2(n19150), .ZN(n12886) );
  OAI211_X1 U16062 ( .C1(n13119), .C2(n12975), .A(n12879), .B(n12886), .ZN(
        P2_U2962) );
  INV_X1 U16063 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19200) );
  NAND2_X1 U16064 ( .A1(n12940), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n12882) );
  NAND2_X1 U16065 ( .A1(n15338), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12881) );
  INV_X1 U16066 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16397) );
  OR2_X1 U16067 ( .A1(n15338), .A2(n16397), .ZN(n12880) );
  NAND2_X1 U16068 ( .A1(n12881), .A2(n12880), .ZN(n19139) );
  NAND2_X1 U16069 ( .A1(n12930), .A2(n19139), .ZN(n12890) );
  OAI211_X1 U16070 ( .C1(n19200), .C2(n12975), .A(n12882), .B(n12890), .ZN(
        P2_U2981) );
  INV_X1 U16071 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12989) );
  NAND2_X1 U16072 ( .A1(n12940), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12885) );
  NAND2_X1 U16073 ( .A1(n15338), .A2(BUF2_REG_12__SCAN_IN), .ZN(n12884) );
  INV_X1 U16074 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16401) );
  OR2_X1 U16075 ( .A1(n15338), .A2(n16401), .ZN(n12883) );
  NAND2_X1 U16076 ( .A1(n12884), .A2(n12883), .ZN(n19145) );
  NAND2_X1 U16077 ( .A1(n12930), .A2(n19145), .ZN(n12888) );
  OAI211_X1 U16078 ( .C1(n12989), .C2(n12975), .A(n12885), .B(n12888), .ZN(
        P2_U2964) );
  INV_X1 U16079 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19208) );
  NAND2_X1 U16080 ( .A1(n12940), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12887) );
  OAI211_X1 U16081 ( .C1(n19208), .C2(n12975), .A(n12887), .B(n12886), .ZN(
        P2_U2977) );
  INV_X1 U16082 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19204) );
  NAND2_X1 U16083 ( .A1(n12940), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12889) );
  OAI211_X1 U16084 ( .C1(n19204), .C2(n12975), .A(n12889), .B(n12888), .ZN(
        P2_U2979) );
  INV_X1 U16085 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13115) );
  NAND2_X1 U16086 ( .A1(n12940), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12891) );
  OAI211_X1 U16087 ( .C1(n13115), .C2(n12975), .A(n12891), .B(n12890), .ZN(
        P2_U2966) );
  INV_X1 U16088 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19212) );
  NAND2_X1 U16089 ( .A1(n12940), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12894) );
  NAND2_X1 U16090 ( .A1(n15338), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12893) );
  INV_X1 U16091 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16408) );
  OR2_X1 U16092 ( .A1(n15338), .A2(n16408), .ZN(n12892) );
  NAND2_X1 U16093 ( .A1(n12893), .A2(n12892), .ZN(n19156) );
  NAND2_X1 U16094 ( .A1(n12930), .A2(n19156), .ZN(n12895) );
  OAI211_X1 U16095 ( .C1(n19212), .C2(n12975), .A(n12894), .B(n12895), .ZN(
        P2_U2975) );
  INV_X1 U16096 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12986) );
  NAND2_X1 U16097 ( .A1(n12940), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12896) );
  OAI211_X1 U16098 ( .C1(n12986), .C2(n12975), .A(n12896), .B(n12895), .ZN(
        P2_U2960) );
  AOI22_X1 U16099 ( .A1(n12940), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(n13486), .ZN(n12901) );
  INV_X1 U16100 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12897) );
  OR2_X1 U16101 ( .A1(n15338), .A2(n12897), .ZN(n12899) );
  NAND2_X1 U16102 ( .A1(n15338), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12898) );
  AND2_X1 U16103 ( .A1(n12899), .A2(n12898), .ZN(n19153) );
  INV_X1 U16104 ( .A(n19153), .ZN(n12900) );
  NAND2_X1 U16105 ( .A1(n12930), .A2(n12900), .ZN(n12932) );
  NAND2_X1 U16106 ( .A1(n12901), .A2(n12932), .ZN(P2_U2961) );
  AOI22_X1 U16107 ( .A1(n12940), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16108 ( .A1(n15340), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15338), .ZN(n19279) );
  INV_X1 U16109 ( .A(n19279), .ZN(n12902) );
  NAND2_X1 U16110 ( .A1(n12930), .A2(n12902), .ZN(n12914) );
  NAND2_X1 U16111 ( .A1(n12903), .A2(n12914), .ZN(P2_U2955) );
  AOI22_X1 U16112 ( .A1(n12940), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(
        P2_EAX_REG_17__SCAN_IN), .B2(n13486), .ZN(n12905) );
  AOI22_X1 U16113 ( .A1(n15340), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15338), .ZN(n19269) );
  INV_X1 U16114 ( .A(n19269), .ZN(n12904) );
  NAND2_X1 U16115 ( .A1(n12930), .A2(n12904), .ZN(n12912) );
  NAND2_X1 U16116 ( .A1(n12905), .A2(n12912), .ZN(P2_U2953) );
  AOI22_X1 U16117 ( .A1(n12940), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(
        P2_EAX_REG_5__SCAN_IN), .B2(n13486), .ZN(n12906) );
  AOI22_X1 U16118 ( .A1(n15340), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15338), .ZN(n19288) );
  INV_X1 U16119 ( .A(n19288), .ZN(n19165) );
  NAND2_X1 U16120 ( .A1(n12930), .A2(n19165), .ZN(n12936) );
  NAND2_X1 U16121 ( .A1(n12906), .A2(n12936), .ZN(P2_U2972) );
  AOI22_X1 U16122 ( .A1(n12940), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(
        P2_EAX_REG_22__SCAN_IN), .B2(n13486), .ZN(n12907) );
  INV_X1 U16123 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16412) );
  INV_X1 U16124 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18185) );
  AOI22_X1 U16125 ( .A1(n15340), .A2(n16412), .B1(n18185), .B2(n15338), .ZN(
        n19161) );
  NAND2_X1 U16126 ( .A1(n12930), .A2(n19161), .ZN(n12908) );
  NAND2_X1 U16127 ( .A1(n12907), .A2(n12908), .ZN(P2_U2958) );
  AOI22_X1 U16128 ( .A1(n12940), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12909) );
  NAND2_X1 U16129 ( .A1(n12909), .A2(n12908), .ZN(P2_U2973) );
  AOI22_X1 U16130 ( .A1(n12940), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12911) );
  INV_X1 U16131 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16420) );
  INV_X1 U16132 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U16133 ( .A1(n15340), .A2(n16420), .B1(n18168), .B2(n15338), .ZN(
        n16082) );
  INV_X1 U16134 ( .A(n16082), .ZN(n19274) );
  OR2_X1 U16135 ( .A1(n12910), .A2(n19274), .ZN(n12941) );
  NAND2_X1 U16136 ( .A1(n12911), .A2(n12941), .ZN(P2_U2969) );
  AOI22_X1 U16137 ( .A1(n12940), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_1__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U16138 ( .A1(n12913), .A2(n12912), .ZN(P2_U2968) );
  AOI22_X1 U16139 ( .A1(n12940), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(
        P2_EAX_REG_3__SCAN_IN), .B2(n13486), .ZN(n12915) );
  NAND2_X1 U16140 ( .A1(n12915), .A2(n12914), .ZN(P2_U2970) );
  AOI22_X1 U16141 ( .A1(n12940), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16142 ( .A1(n15340), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15338), .ZN(n19159) );
  INV_X1 U16143 ( .A(n19159), .ZN(n12916) );
  NAND2_X1 U16144 ( .A1(n12930), .A2(n12916), .ZN(n12934) );
  NAND2_X1 U16145 ( .A1(n12917), .A2(n12934), .ZN(P2_U2974) );
  AOI22_X1 U16146 ( .A1(n12940), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_29__SCAN_IN), .B2(n13486), .ZN(n12921) );
  INV_X1 U16147 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16399) );
  OR2_X1 U16148 ( .A1(n15338), .A2(n16399), .ZN(n12919) );
  NAND2_X1 U16149 ( .A1(n15338), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12918) );
  AND2_X1 U16150 ( .A1(n12919), .A2(n12918), .ZN(n19142) );
  INV_X1 U16151 ( .A(n19142), .ZN(n12920) );
  NAND2_X1 U16152 ( .A1(n12930), .A2(n12920), .ZN(n12922) );
  NAND2_X1 U16153 ( .A1(n12921), .A2(n12922), .ZN(P2_U2965) );
  AOI22_X1 U16154 ( .A1(n12940), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(
        P2_EAX_REG_13__SCAN_IN), .B2(n13486), .ZN(n12923) );
  NAND2_X1 U16155 ( .A1(n12923), .A2(n12922), .ZN(P2_U2980) );
  AOI22_X1 U16156 ( .A1(n12940), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_27__SCAN_IN), .B2(n13486), .ZN(n12927) );
  INV_X1 U16157 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16403) );
  OR2_X1 U16158 ( .A1(n15338), .A2(n16403), .ZN(n12925) );
  NAND2_X1 U16159 ( .A1(n15338), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12924) );
  AND2_X1 U16160 ( .A1(n12925), .A2(n12924), .ZN(n19148) );
  INV_X1 U16161 ( .A(n19148), .ZN(n12926) );
  NAND2_X1 U16162 ( .A1(n12930), .A2(n12926), .ZN(n12928) );
  NAND2_X1 U16163 ( .A1(n12927), .A2(n12928), .ZN(P2_U2963) );
  AOI22_X1 U16164 ( .A1(n12940), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(
        P2_EAX_REG_11__SCAN_IN), .B2(n13486), .ZN(n12929) );
  NAND2_X1 U16165 ( .A1(n12929), .A2(n12928), .ZN(P2_U2978) );
  AOI22_X1 U16166 ( .A1(n12940), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_4__SCAN_IN), .B2(n13486), .ZN(n12931) );
  INV_X1 U16167 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16416) );
  INV_X1 U16168 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U16169 ( .A1(n15340), .A2(n16416), .B1(n18177), .B2(n15338), .ZN(
        n19173) );
  NAND2_X1 U16170 ( .A1(n12930), .A2(n19173), .ZN(n12938) );
  NAND2_X1 U16171 ( .A1(n12931), .A2(n12938), .ZN(P2_U2971) );
  AOI22_X1 U16172 ( .A1(n12940), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(
        P2_EAX_REG_9__SCAN_IN), .B2(n13486), .ZN(n12933) );
  NAND2_X1 U16173 ( .A1(n12933), .A2(n12932), .ZN(P2_U2976) );
  AOI22_X1 U16174 ( .A1(n12940), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16175 ( .A1(n12935), .A2(n12934), .ZN(P2_U2959) );
  AOI22_X1 U16176 ( .A1(n12940), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n13486), 
        .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12937) );
  NAND2_X1 U16177 ( .A1(n12937), .A2(n12936), .ZN(P2_U2957) );
  AOI22_X1 U16178 ( .A1(n12940), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(
        P2_EAX_REG_20__SCAN_IN), .B2(n13486), .ZN(n12939) );
  NAND2_X1 U16179 ( .A1(n12939), .A2(n12938), .ZN(P2_U2956) );
  AOI22_X1 U16180 ( .A1(n12940), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(
        P2_EAX_REG_18__SCAN_IN), .B2(n13486), .ZN(n12942) );
  NAND2_X1 U16181 ( .A1(n12942), .A2(n12941), .ZN(P2_U2954) );
  OR2_X1 U16182 ( .A1(n12962), .A2(n13128), .ZN(n12943) );
  INV_X1 U16183 ( .A(n12964), .ZN(n12944) );
  NAND2_X1 U16184 ( .A1(n11629), .A2(n12944), .ZN(n12946) );
  INV_X1 U16185 ( .A(n20658), .ZN(n20651) );
  NOR2_X1 U16186 ( .A1(n20651), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12970) );
  AOI21_X1 U16187 ( .B1(n12971), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n12970), 
        .ZN(n12945) );
  NAND2_X1 U16188 ( .A1(n13172), .A2(n12945), .ZN(P1_U2801) );
  AND2_X1 U16189 ( .A1(n12946), .A2(n12962), .ZN(n12947) );
  AOI21_X1 U16190 ( .B1(n13155), .B2(n12958), .A(n12947), .ZN(n12960) );
  AND2_X1 U16191 ( .A1(n12960), .A2(n13153), .ZN(n12950) );
  INV_X1 U16192 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n12949) );
  NAND3_X1 U16193 ( .A1(n15942), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n20721), 
        .ZN(n12948) );
  OAI21_X1 U16194 ( .B1(n12950), .B2(n12949), .A(n12948), .ZN(P1_U2803) );
  OR2_X1 U16195 ( .A1(n19063), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12951) );
  AND2_X1 U16196 ( .A1(n13890), .A2(n12951), .ZN(n16256) );
  OAI21_X1 U16197 ( .B1(n12953), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12952), .ZN(n16263) );
  OAI21_X1 U16198 ( .B1(n19239), .B2(n12954), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12955) );
  NAND2_X1 U16199 ( .A1(n12763), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n16261) );
  OAI211_X1 U16200 ( .C1(n16172), .C2(n16263), .A(n12955), .B(n16261), .ZN(
        n12956) );
  AOI21_X1 U16201 ( .B1(n19240), .B2(n16256), .A(n12956), .ZN(n12957) );
  OAI21_X1 U16202 ( .B1(n16252), .B2(n15339), .A(n12957), .ZN(P2_U3014) );
  NAND3_X1 U16203 ( .A1(n12958), .A2(n15564), .A3(n13129), .ZN(n12959) );
  NAND2_X1 U16204 ( .A1(n12959), .A2(n20800), .ZN(n20803) );
  AND2_X1 U16205 ( .A1(n12960), .A2(n20803), .ZN(n15528) );
  NOR2_X1 U16206 ( .A1(n15528), .A2(n13128), .ZN(n19997) );
  INV_X1 U16207 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15526) );
  INV_X1 U16208 ( .A(n13314), .ZN(n12961) );
  OR2_X1 U16209 ( .A1(n13155), .A2(n12961), .ZN(n12968) );
  NAND2_X1 U16210 ( .A1(n13155), .A2(n10166), .ZN(n12967) );
  NAND2_X1 U16211 ( .A1(n13155), .A2(n12963), .ZN(n12966) );
  NAND2_X1 U16212 ( .A1(n11629), .A2(n12964), .ZN(n12965) );
  NAND4_X1 U16213 ( .A1(n12968), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        n15525) );
  NAND2_X1 U16214 ( .A1(n19997), .A2(n15525), .ZN(n12969) );
  OAI21_X1 U16215 ( .B1(n19997), .B2(n15526), .A(n12969), .ZN(P1_U3484) );
  NOR2_X1 U16216 ( .A1(n12970), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12973)
         );
  OAI21_X1 U16217 ( .B1(n11692), .B2(n13439), .A(n20798), .ZN(n12972) );
  OAI21_X1 U16218 ( .B1(n12973), .B2(n20798), .A(n12972), .ZN(P1_U3487) );
  INV_X1 U16219 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n12979) );
  NOR2_X1 U16220 ( .A1(n13011), .A2(n12584), .ZN(n12974) );
  NAND2_X1 U16221 ( .A1(n16272), .A2(n12974), .ZN(n12993) );
  OAI21_X1 U16222 ( .B1(n12993), .B2(n13007), .A(n12975), .ZN(n12976) );
  NAND2_X1 U16223 ( .A1(n19197), .A2(n12977), .ZN(n13123) );
  OR2_X1 U16224 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13005), .ZN(n19975) );
  INV_X2 U16225 ( .A(n19975), .ZN(n13117) );
  AOI22_X1 U16226 ( .A1(n13117), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12978) );
  OAI21_X1 U16227 ( .B1(n12979), .B2(n13123), .A(n12978), .ZN(P2_U2929) );
  INV_X1 U16228 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U16229 ( .A1(n13117), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12980) );
  OAI21_X1 U16230 ( .B1(n14874), .B2(n13123), .A(n12980), .ZN(P2_U2930) );
  INV_X1 U16231 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14842) );
  AOI22_X1 U16232 ( .A1(n13117), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12981) );
  OAI21_X1 U16233 ( .B1(n14842), .B2(n13123), .A(n12981), .ZN(P2_U2926) );
  INV_X1 U16234 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14883) );
  AOI22_X1 U16235 ( .A1(n13117), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12982) );
  OAI21_X1 U16236 ( .B1(n14883), .B2(n13123), .A(n12982), .ZN(P2_U2932) );
  INV_X1 U16237 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16238 ( .A1(n13117), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12983) );
  OAI21_X1 U16239 ( .B1(n12984), .B2(n13123), .A(n12983), .ZN(P2_U2931) );
  AOI22_X1 U16240 ( .A1(n13117), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12985) );
  OAI21_X1 U16241 ( .B1(n12986), .B2(n13123), .A(n12985), .ZN(P2_U2927) );
  INV_X1 U16242 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n14865) );
  AOI22_X1 U16243 ( .A1(n13117), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12987) );
  OAI21_X1 U16244 ( .B1(n14865), .B2(n13123), .A(n12987), .ZN(P2_U2928) );
  AOI22_X1 U16245 ( .A1(n13117), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12988) );
  OAI21_X1 U16246 ( .B1(n12989), .B2(n13123), .A(n12988), .ZN(P2_U2923) );
  INV_X1 U16247 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14827) );
  AOI22_X1 U16248 ( .A1(n13117), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12990) );
  OAI21_X1 U16249 ( .B1(n14827), .B2(n13123), .A(n12990), .ZN(P2_U2924) );
  INV_X1 U16250 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16251 ( .A1(n13117), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19196), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12991) );
  OAI21_X1 U16252 ( .B1(n12992), .B2(n13123), .A(n12991), .ZN(P2_U2933) );
  INV_X1 U16253 ( .A(n12993), .ZN(n12995) );
  NAND2_X1 U16254 ( .A1(n12995), .A2(n12994), .ZN(n13004) );
  NAND2_X1 U16255 ( .A1(n13001), .A2(n16269), .ZN(n13014) );
  INV_X1 U16256 ( .A(n12996), .ZN(n12997) );
  AND2_X1 U16257 ( .A1(n13014), .A2(n12997), .ZN(n13003) );
  NAND2_X1 U16258 ( .A1(n12999), .A2(n12998), .ZN(n13000) );
  OAI21_X1 U16259 ( .B1(n13001), .B2(n16271), .A(n13000), .ZN(n13051) );
  INV_X1 U16260 ( .A(n13051), .ZN(n13002) );
  INV_X1 U16261 ( .A(n13005), .ZN(n19955) );
  NAND2_X1 U16262 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19955), .ZN(n16324) );
  OAI22_X1 U16263 ( .A1(n16293), .A2(n13007), .B1(n13006), .B2(n16324), .ZN(
        n13008) );
  AOI21_X1 U16264 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13470), .A(n13008), 
        .ZN(n19918) );
  INV_X1 U16265 ( .A(n19918), .ZN(n13578) );
  INV_X1 U16266 ( .A(n13009), .ZN(n13010) );
  NOR3_X1 U16267 ( .A1(n13011), .A2(n13010), .A3(n19976), .ZN(n16273) );
  NAND3_X1 U16268 ( .A1(n13578), .A2(n19831), .A3(n16273), .ZN(n13012) );
  OAI21_X1 U16269 ( .B1(n13578), .B2(n13013), .A(n13012), .ZN(P2_U3595) );
  NAND2_X1 U16270 ( .A1(n13014), .A2(n15307), .ZN(n13015) );
  INV_X1 U16271 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n19064) );
  NAND2_X1 U16272 ( .A1(n19076), .A2(n13089), .ZN(n13019) );
  NAND2_X1 U16273 ( .A1(n13016), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13017) );
  NAND2_X1 U16274 ( .A1(n13017), .A2(n19971), .ZN(n13093) );
  AOI22_X1 U16275 ( .A1(n13093), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19728), .B2(n19958), .ZN(n13018) );
  NOR2_X1 U16276 ( .A1(n13016), .A2(n13470), .ZN(n13024) );
  AOI21_X1 U16277 ( .B1(n19976), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13020) );
  AND2_X1 U16278 ( .A1(n13024), .A2(n13020), .ZN(n13021) );
  NAND2_X1 U16279 ( .A1(n19121), .A2(n15344), .ZN(n19117) );
  NAND2_X1 U16280 ( .A1(n19527), .A2(n19107), .ZN(n13023) );
  NAND2_X1 U16281 ( .A1(n19076), .A2(n19121), .ZN(n13022) );
  OAI211_X1 U16282 ( .C1(n19121), .C2(n19064), .A(n13023), .B(n13022), .ZN(
        P2_U2887) );
  INV_X1 U16283 ( .A(n14198), .ZN(n14166) );
  INV_X1 U16284 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19272) );
  NAND2_X1 U16285 ( .A1(n13093), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13026) );
  XNOR2_X1 U16286 ( .A(n19958), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19417) );
  NAND2_X1 U16287 ( .A1(n19417), .A2(n19728), .ZN(n19592) );
  NAND2_X1 U16288 ( .A1(n13026), .A2(n19592), .ZN(n13027) );
  MUX2_X1 U16289 ( .A(n9961), .B(n13910), .S(n19121), .Z(n13028) );
  OAI21_X1 U16290 ( .B1(n19361), .B2(n19117), .A(n13028), .ZN(P2_U2886) );
  NAND2_X1 U16291 ( .A1(n13029), .A2(n13089), .ZN(n13033) );
  NAND2_X1 U16292 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19622) );
  NAND2_X1 U16293 ( .A1(n19622), .A2(n13030), .ZN(n13031) );
  NOR2_X1 U16294 ( .A1(n13030), .A2(n19949), .ZN(n19727) );
  NAND2_X1 U16295 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19727), .ZN(
        n15326) );
  AND2_X1 U16296 ( .A1(n13031), .A2(n15326), .ZN(n19418) );
  AOI22_X1 U16297 ( .A1(n13093), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n19728), .B2(n19418), .ZN(n13032) );
  INV_X1 U16298 ( .A(n13039), .ZN(n13040) );
  INV_X1 U16299 ( .A(n13087), .ZN(n13043) );
  INV_X1 U16300 ( .A(n19940), .ZN(n19917) );
  MUX2_X1 U16301 ( .A(n13485), .B(n16283), .S(n19121), .Z(n13044) );
  OAI21_X1 U16302 ( .B1(n19917), .B2(n19117), .A(n13044), .ZN(P2_U2885) );
  NAND2_X1 U16303 ( .A1(n12584), .A2(n13045), .ZN(n13046) );
  OR2_X1 U16304 ( .A1(n9819), .A2(n13046), .ZN(n13049) );
  NOR2_X1 U16305 ( .A1(n13049), .A2(n13048), .ZN(n13050) );
  NAND2_X1 U16306 ( .A1(n19162), .A2(n12583), .ZN(n14884) );
  NAND2_X1 U16307 ( .A1(n19162), .A2(n13053), .ZN(n13683) );
  NAND2_X1 U16308 ( .A1(n14884), .A2(n13683), .ZN(n19164) );
  INV_X1 U16309 ( .A(n13054), .ZN(n13060) );
  INV_X1 U16310 ( .A(n13055), .ZN(n13058) );
  INV_X1 U16311 ( .A(n13056), .ZN(n13057) );
  NAND2_X1 U16312 ( .A1(n13058), .A2(n13057), .ZN(n13059) );
  NAND2_X1 U16313 ( .A1(n13060), .A2(n13059), .ZN(n13061) );
  INV_X1 U16314 ( .A(n13061), .ZN(n19070) );
  NOR2_X1 U16315 ( .A1(n19952), .A2(n13061), .ZN(n19190) );
  INV_X1 U16316 ( .A(n19190), .ZN(n13063) );
  OAI211_X1 U16317 ( .C1(n19527), .C2(n19070), .A(n13063), .B(n19176), .ZN(
        n13066) );
  AOI22_X1 U16318 ( .A1(n19187), .A2(n19070), .B1(n19186), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13065) );
  OAI211_X1 U16319 ( .C1(n19195), .C2(n15328), .A(n13066), .B(n13065), .ZN(
        P2_U2919) );
  NOR2_X1 U16320 ( .A1(n16232), .A2(n12075), .ZN(n19244) );
  INV_X1 U16321 ( .A(n13067), .ZN(n13722) );
  NAND2_X1 U16322 ( .A1(n13069), .A2(n13068), .ZN(n13070) );
  AND2_X1 U16323 ( .A1(n13071), .A2(n13070), .ZN(n19241) );
  NAND2_X1 U16324 ( .A1(n13073), .A2(n13072), .ZN(n13076) );
  INV_X1 U16325 ( .A(n13074), .ZN(n13075) );
  AND2_X1 U16326 ( .A1(n13076), .A2(n13075), .ZN(n19935) );
  INV_X1 U16327 ( .A(n19935), .ZN(n13293) );
  AOI22_X1 U16328 ( .A1(n19241), .A2(n19263), .B1(n13293), .B2(n19257), .ZN(
        n13077) );
  OAI221_X1 U16329 ( .B1(n15202), .B2(n13722), .C1(n15202), .C2(n13078), .A(
        n13077), .ZN(n13079) );
  AOI211_X1 U16330 ( .C1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .C2(n13080), .A(
        n19244), .B(n13079), .ZN(n13085) );
  XOR2_X1 U16331 ( .A(n13082), .B(n13081), .Z(n19243) );
  AOI22_X1 U16332 ( .A1(n19262), .A2(n19243), .B1(n13888), .B2(n13083), .ZN(
        n13084) );
  OAI211_X1 U16333 ( .C1(n16283), .C2(n16253), .A(n13085), .B(n13084), .ZN(
        P2_U3044) );
  INV_X1 U16334 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19933) );
  NAND2_X1 U16335 ( .A1(n19727), .A2(n19933), .ZN(n19504) );
  INV_X1 U16336 ( .A(n19504), .ZN(n13090) );
  INV_X1 U16337 ( .A(n19534), .ZN(n19531) );
  NAND2_X1 U16338 ( .A1(n15326), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13091) );
  NAND2_X1 U16339 ( .A1(n19531), .A2(n13091), .ZN(n13092) );
  AND2_X1 U16340 ( .A1(n13092), .A2(n19728), .ZN(n19652) );
  AOI21_X1 U16341 ( .B1(n13093), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19652), .ZN(n13094) );
  AND2_X1 U16342 ( .A1(n14198), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13095) );
  NAND2_X1 U16343 ( .A1(n13221), .A2(n13095), .ZN(n19029) );
  INV_X2 U16344 ( .A(n19121), .ZN(n19116) );
  INV_X1 U16345 ( .A(n13099), .ZN(n16244) );
  NOR2_X1 U16346 ( .A1(n16244), .A2(n19116), .ZN(n13100) );
  AOI21_X1 U16347 ( .B1(P2_EBX_REG_3__SCAN_IN), .B2(n19116), .A(n13100), .ZN(
        n13101) );
  OAI21_X1 U16348 ( .B1(n19925), .B2(n19117), .A(n13101), .ZN(P2_U2884) );
  INV_X1 U16349 ( .A(n13102), .ZN(n13105) );
  INV_X1 U16350 ( .A(n13103), .ZN(n13104) );
  AOI21_X1 U16351 ( .B1(n13105), .B2(n15823), .A(n13104), .ZN(n20126) );
  INV_X1 U16352 ( .A(n20126), .ZN(n13113) );
  NOR2_X1 U16353 ( .A1(n13106), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13108) );
  OR2_X1 U16354 ( .A1(n13108), .A2(n13107), .ZN(n13134) );
  INV_X1 U16355 ( .A(n13134), .ZN(n20066) );
  AND2_X1 U16356 ( .A1(n15823), .A2(n13229), .ZN(n13110) );
  NAND2_X1 U16357 ( .A1(n15899), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20129) );
  INV_X1 U16358 ( .A(n20129), .ZN(n13109) );
  AOI211_X1 U16359 ( .C1(n15932), .C2(n20066), .A(n13110), .B(n13109), .ZN(
        n13112) );
  OAI21_X1 U16360 ( .B1(n15816), .B2(n15819), .A(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13111) );
  OAI211_X1 U16361 ( .C1(n20138), .C2(n13113), .A(n13112), .B(n13111), .ZN(
        P1_U3031) );
  AOI22_X1 U16362 ( .A1(n13117), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n19227), .ZN(n13114) );
  OAI21_X1 U16363 ( .B1(n13115), .B2(n13123), .A(n13114), .ZN(P2_U2921) );
  INV_X1 U16364 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14815) );
  AOI22_X1 U16365 ( .A1(n13117), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13116) );
  OAI21_X1 U16366 ( .B1(n14815), .B2(n13123), .A(n13116), .ZN(P2_U2922) );
  AOI22_X1 U16367 ( .A1(n13117), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13118) );
  OAI21_X1 U16368 ( .B1(n13119), .B2(n13123), .A(n13118), .ZN(P2_U2925) );
  AOI22_X1 U16369 ( .A1(n13117), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13120) );
  OAI21_X1 U16370 ( .B1(n13121), .B2(n13123), .A(n13120), .ZN(P2_U2935) );
  INV_X1 U16371 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13682) );
  AOI22_X1 U16372 ( .A1(n13117), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13122) );
  OAI21_X1 U16373 ( .B1(n13682), .B2(n13123), .A(n13122), .ZN(P2_U2934) );
  NAND2_X1 U16374 ( .A1(n13125), .A2(n13124), .ZN(n13126) );
  NAND2_X1 U16375 ( .A1(n13127), .A2(n13126), .ZN(n20132) );
  NAND2_X1 U16376 ( .A1(n13155), .A2(n13314), .ZN(n13145) );
  OAI222_X1 U16377 ( .A1(n20132), .A2(n14439), .B1(n20078), .B2(n11648), .C1(
        n13134), .C2(n15712), .ZN(P1_U2872) );
  INV_X1 U16378 ( .A(n11154), .ZN(n15941) );
  OR2_X1 U16379 ( .A1(n13135), .A2(n11114), .ZN(n13136) );
  OR3_X1 U16380 ( .A1(n13137), .A2(n15941), .A3(n13136), .ZN(n13338) );
  NAND2_X1 U16381 ( .A1(n10503), .A2(n13338), .ZN(n13139) );
  INV_X1 U16382 ( .A(n10401), .ZN(n14724) );
  NAND2_X1 U16383 ( .A1(n14724), .A2(n10241), .ZN(n13138) );
  NAND2_X1 U16384 ( .A1(n13139), .A2(n13138), .ZN(n15508) );
  OAI22_X1 U16385 ( .A1(n20717), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20786), .ZN(n13140) );
  AOI21_X1 U16386 ( .B1(n15508), .B2(n15942), .A(n13140), .ZN(n13152) );
  INV_X1 U16387 ( .A(n13141), .ZN(n15539) );
  INV_X1 U16388 ( .A(n15564), .ZN(n15537) );
  OAI21_X1 U16389 ( .B1(n15506), .B2(n15539), .A(n15537), .ZN(n13147) );
  NAND2_X1 U16390 ( .A1(n13442), .A2(n13142), .ZN(n13143) );
  AND2_X1 U16391 ( .A1(n13144), .A2(n13143), .ZN(n13146) );
  OAI211_X1 U16392 ( .C1(n15543), .C2(n13147), .A(n13146), .B(n13145), .ZN(
        n13148) );
  OR2_X1 U16393 ( .A1(n13149), .A2(n13148), .ZN(n15505) );
  NAND2_X1 U16394 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15954) );
  NOR2_X1 U16395 ( .A1(n20718), .A2(n15954), .ZN(n13349) );
  AOI22_X1 U16396 ( .A1(n15505), .A2(n13153), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n13349), .ZN(n15940) );
  OAI21_X1 U16397 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n20537), .A(n15940), 
        .ZN(n20790) );
  INV_X1 U16398 ( .A(n20790), .ZN(n13151) );
  AOI21_X1 U16399 ( .B1(n15506), .B2(n15942), .A(n13151), .ZN(n13150) );
  OAI22_X1 U16400 ( .A1(n13152), .A2(n13151), .B1(n13150), .B2(n10241), .ZN(
        P1_U3474) );
  NAND2_X1 U16401 ( .A1(n15506), .A2(n13153), .ZN(n13154) );
  OAI22_X1 U16402 ( .A1(n13172), .A2(n13447), .B1(n13155), .B2(n13154), .ZN(
        n13156) );
  NAND2_X1 U16403 ( .A1(n20082), .A2(n13443), .ZN(n13375) );
  NOR2_X1 U16404 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15954), .ZN(n20106) );
  INV_X1 U16405 ( .A(n20106), .ZN(n20080) );
  NOR2_X4 U16406 ( .A1(n20082), .A2(n20801), .ZN(n15566) );
  AOI22_X1 U16407 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13157) );
  OAI21_X1 U16408 ( .B1(n14474), .B2(n13375), .A(n13157), .ZN(P1_U2914) );
  INV_X1 U16409 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13242) );
  AOI22_X1 U16410 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13158) );
  OAI21_X1 U16411 ( .B1(n13242), .B2(n13375), .A(n13158), .ZN(P1_U2908) );
  INV_X1 U16412 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13160) );
  AOI22_X1 U16413 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13159) );
  OAI21_X1 U16414 ( .B1(n13160), .B2(n13375), .A(n13159), .ZN(P1_U2917) );
  INV_X1 U16415 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13239) );
  AOI22_X1 U16416 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13161) );
  OAI21_X1 U16417 ( .B1(n13239), .B2(n13375), .A(n13161), .ZN(P1_U2911) );
  INV_X1 U16418 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13163) );
  AOI22_X1 U16419 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13162) );
  OAI21_X1 U16420 ( .B1(n13163), .B2(n13375), .A(n13162), .ZN(P1_U2912) );
  INV_X1 U16421 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U16422 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13164) );
  OAI21_X1 U16423 ( .B1(n20890), .B2(n13375), .A(n13164), .ZN(P1_U2909) );
  AOI22_X1 U16424 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U16425 ( .B1(n14481), .B2(n13375), .A(n13165), .ZN(P1_U2916) );
  INV_X1 U16426 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n21036) );
  AOI22_X1 U16427 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13166) );
  OAI21_X1 U16428 ( .B1(n21036), .B2(n13375), .A(n13166), .ZN(P1_U2913) );
  INV_X1 U16429 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16430 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13167) );
  OAI21_X1 U16431 ( .B1(n13168), .B2(n13375), .A(n13167), .ZN(P1_U2915) );
  INV_X1 U16432 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13170) );
  AOI22_X1 U16433 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13169) );
  OAI21_X1 U16434 ( .B1(n13170), .B2(n13375), .A(n13169), .ZN(P1_U2918) );
  NOR2_X1 U16435 ( .A1(n15538), .A2(n20800), .ZN(n13171) );
  INV_X2 U16436 ( .A(n13255), .ZN(n20120) );
  AOI22_X1 U16437 ( .A1(n20121), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13175) );
  NAND2_X1 U16438 ( .A1(n13255), .A2(n13447), .ZN(n13256) );
  INV_X1 U16439 ( .A(DATAI_1_), .ZN(n13174) );
  NAND2_X1 U16440 ( .A1(n13593), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13173) );
  OAI21_X1 U16441 ( .B1(n13593), .B2(n13174), .A(n13173), .ZN(n20158) );
  NAND2_X1 U16442 ( .A1(n13251), .A2(n20158), .ZN(n13197) );
  NAND2_X1 U16443 ( .A1(n13175), .A2(n13197), .ZN(P1_U2938) );
  AOI22_X1 U16444 ( .A1(n20121), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13178) );
  INV_X1 U16445 ( .A(DATAI_0_), .ZN(n21108) );
  NAND2_X1 U16446 ( .A1(n13594), .A2(n21108), .ZN(n13177) );
  NAND2_X1 U16447 ( .A1(n13593), .A2(n16427), .ZN(n13176) );
  AND2_X1 U16448 ( .A1(n13177), .A2(n13176), .ZN(n20151) );
  NAND2_X1 U16449 ( .A1(n13251), .A2(n20151), .ZN(n13212) );
  NAND2_X1 U16450 ( .A1(n13178), .A2(n13212), .ZN(P1_U2952) );
  AOI22_X1 U16451 ( .A1(n20121), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13179) );
  MUX2_X1 U16452 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n13593), .Z(
        n14465) );
  NAND2_X1 U16453 ( .A1(n13251), .A2(n14465), .ZN(n13236) );
  NAND2_X1 U16454 ( .A1(n13179), .A2(n13236), .ZN(P1_U2945) );
  AOI22_X1 U16455 ( .A1(n20121), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13182) );
  INV_X1 U16456 ( .A(DATAI_3_), .ZN(n20984) );
  NAND2_X1 U16457 ( .A1(n13594), .A2(n20984), .ZN(n13181) );
  INV_X1 U16458 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16418) );
  NAND2_X1 U16459 ( .A1(n13593), .A2(n16418), .ZN(n13180) );
  AND2_X1 U16460 ( .A1(n13181), .A2(n13180), .ZN(n20169) );
  NAND2_X1 U16461 ( .A1(n13251), .A2(n20169), .ZN(n13186) );
  NAND2_X1 U16462 ( .A1(n13182), .A2(n13186), .ZN(P1_U2955) );
  AOI22_X1 U16463 ( .A1(n20121), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13185) );
  INV_X1 U16464 ( .A(DATAI_2_), .ZN(n21119) );
  NAND2_X1 U16465 ( .A1(n13594), .A2(n21119), .ZN(n13184) );
  NAND2_X1 U16466 ( .A1(n13593), .A2(n16420), .ZN(n13183) );
  AND2_X1 U16467 ( .A1(n13184), .A2(n13183), .ZN(n20162) );
  NAND2_X1 U16468 ( .A1(n13251), .A2(n20162), .ZN(n13199) );
  NAND2_X1 U16469 ( .A1(n13185), .A2(n13199), .ZN(P1_U2939) );
  AOI22_X1 U16470 ( .A1(n20121), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13187) );
  NAND2_X1 U16471 ( .A1(n13187), .A2(n13186), .ZN(P1_U2940) );
  AOI22_X1 U16472 ( .A1(n20121), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13190) );
  INV_X1 U16473 ( .A(DATAI_4_), .ZN(n20931) );
  NAND2_X1 U16474 ( .A1(n13594), .A2(n20931), .ZN(n13189) );
  NAND2_X1 U16475 ( .A1(n13593), .A2(n16416), .ZN(n13188) );
  AND2_X1 U16476 ( .A1(n13189), .A2(n13188), .ZN(n14483) );
  NAND2_X1 U16477 ( .A1(n13251), .A2(n14483), .ZN(n13204) );
  NAND2_X1 U16478 ( .A1(n13190), .A2(n13204), .ZN(P1_U2941) );
  AOI22_X1 U16479 ( .A1(n20121), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13193) );
  INV_X1 U16480 ( .A(DATAI_5_), .ZN(n20894) );
  NAND2_X1 U16481 ( .A1(n13594), .A2(n20894), .ZN(n13192) );
  INV_X1 U16482 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16414) );
  NAND2_X1 U16483 ( .A1(n13593), .A2(n16414), .ZN(n13191) );
  AND2_X1 U16484 ( .A1(n13192), .A2(n13191), .ZN(n20175) );
  NAND2_X1 U16485 ( .A1(n13251), .A2(n20175), .ZN(n13206) );
  NAND2_X1 U16486 ( .A1(n13193), .A2(n13206), .ZN(P1_U2942) );
  AOI22_X1 U16487 ( .A1(n20121), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13196) );
  INV_X1 U16488 ( .A(DATAI_6_), .ZN(n20983) );
  NAND2_X1 U16489 ( .A1(n13594), .A2(n20983), .ZN(n13195) );
  NAND2_X1 U16490 ( .A1(n13593), .A2(n16412), .ZN(n13194) );
  AND2_X1 U16491 ( .A1(n13195), .A2(n13194), .ZN(n20183) );
  NAND2_X1 U16492 ( .A1(n13251), .A2(n20183), .ZN(n13208) );
  NAND2_X1 U16493 ( .A1(n13196), .A2(n13208), .ZN(P1_U2943) );
  AOI22_X1 U16494 ( .A1(n20121), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13198) );
  NAND2_X1 U16495 ( .A1(n13198), .A2(n13197), .ZN(P1_U2953) );
  AOI22_X1 U16496 ( .A1(n20121), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13200) );
  NAND2_X1 U16497 ( .A1(n13200), .A2(n13199), .ZN(P1_U2954) );
  AOI22_X1 U16498 ( .A1(n20121), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13203) );
  INV_X1 U16499 ( .A(DATAI_7_), .ZN(n20956) );
  NAND2_X1 U16500 ( .A1(n13594), .A2(n20956), .ZN(n13202) );
  INV_X1 U16501 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16410) );
  NAND2_X1 U16502 ( .A1(n13593), .A2(n16410), .ZN(n13201) );
  AND2_X1 U16503 ( .A1(n13202), .A2(n13201), .ZN(n14469) );
  NAND2_X1 U16504 ( .A1(n13251), .A2(n14469), .ZN(n13210) );
  NAND2_X1 U16505 ( .A1(n13203), .A2(n13210), .ZN(P1_U2944) );
  AOI22_X1 U16506 ( .A1(n20121), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13205) );
  NAND2_X1 U16507 ( .A1(n13205), .A2(n13204), .ZN(P1_U2956) );
  AOI22_X1 U16508 ( .A1(n20121), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13207) );
  NAND2_X1 U16509 ( .A1(n13207), .A2(n13206), .ZN(P1_U2957) );
  AOI22_X1 U16510 ( .A1(n20121), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13209) );
  NAND2_X1 U16511 ( .A1(n13209), .A2(n13208), .ZN(P1_U2958) );
  AOI22_X1 U16512 ( .A1(n20121), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20120), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13211) );
  NAND2_X1 U16513 ( .A1(n13211), .A2(n13210), .ZN(P1_U2959) );
  AOI22_X1 U16514 ( .A1(n20121), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20120), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13213) );
  NAND2_X1 U16515 ( .A1(n13213), .A2(n13212), .ZN(P1_U2937) );
  OR2_X1 U16516 ( .A1(n13215), .A2(n13214), .ZN(n13216) );
  NAND2_X1 U16517 ( .A1(n13267), .A2(n13216), .ZN(n13523) );
  XNOR2_X1 U16518 ( .A(n13515), .B(n13217), .ZN(n13234) );
  INV_X1 U16519 ( .A(n20078), .ZN(n14437) );
  AOI22_X1 U16520 ( .A1(n20073), .A2(n13234), .B1(n14437), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13218) );
  OAI21_X1 U16521 ( .B1(n14439), .B2(n13523), .A(n13218), .ZN(P1_U2871) );
  NAND2_X1 U16522 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13016), .ZN(
        n13219) );
  NAND2_X1 U16523 ( .A1(n13221), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13222) );
  AND2_X1 U16524 ( .A1(n14198), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n19028) );
  XOR2_X1 U16525 ( .A(n13258), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13227)
         );
  AOI21_X1 U16526 ( .B1(n13224), .B2(n13223), .A(n13261), .ZN(n19020) );
  NOR2_X1 U16527 ( .A1(n19121), .A2(n11907), .ZN(n13225) );
  AOI21_X1 U16528 ( .B1(n19020), .B2(n19121), .A(n13225), .ZN(n13226) );
  OAI21_X1 U16529 ( .B1(n13227), .B2(n19117), .A(n13226), .ZN(P2_U2882) );
  XNOR2_X1 U16530 ( .A(n13228), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13302) );
  AOI21_X1 U16531 ( .B1(n15823), .B2(n13229), .A(n15819), .ZN(n13230) );
  NAND2_X1 U16532 ( .A1(n15935), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13297) );
  OAI21_X1 U16533 ( .B1(n14730), .B2(n13230), .A(n13297), .ZN(n13233) );
  NOR3_X1 U16534 ( .A1(n15846), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n13231), .ZN(n13232) );
  AOI211_X1 U16535 ( .C1(n15932), .C2(n13234), .A(n13233), .B(n13232), .ZN(
        n13235) );
  OAI21_X1 U16536 ( .B1(n13302), .B2(n20138), .A(n13235), .ZN(P1_U3030) );
  INV_X1 U16537 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20093) );
  NAND2_X1 U16538 ( .A1(n20120), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13237) );
  OAI211_X1 U16539 ( .C1(n13257), .C2(n20093), .A(n13237), .B(n13236), .ZN(
        P1_U2960) );
  MUX2_X1 U16540 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n13593), .Z(
        n14462) );
  NAND2_X1 U16541 ( .A1(n13251), .A2(n14462), .ZN(n20110) );
  NAND2_X1 U16542 ( .A1(n20120), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n13238) );
  OAI211_X1 U16543 ( .C1(n13257), .C2(n13239), .A(n20110), .B(n13238), .ZN(
        P1_U2946) );
  INV_X1 U16544 ( .A(DATAI_12_), .ZN(n21016) );
  MUX2_X1 U16545 ( .A(n21016), .B(n16401), .S(n13593), .Z(n14446) );
  INV_X1 U16546 ( .A(n14446), .ZN(n13240) );
  NAND2_X1 U16547 ( .A1(n13251), .A2(n13240), .ZN(n20116) );
  NAND2_X1 U16548 ( .A1(n20120), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13241) );
  OAI211_X1 U16549 ( .C1(n13257), .C2(n13242), .A(n20116), .B(n13241), .ZN(
        P1_U2949) );
  INV_X1 U16550 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13369) );
  INV_X1 U16551 ( .A(DATAI_13_), .ZN(n20993) );
  NAND2_X1 U16552 ( .A1(n13593), .A2(BUF1_REG_13__SCAN_IN), .ZN(n13243) );
  OAI21_X1 U16553 ( .B1(n13593), .B2(n20993), .A(n13243), .ZN(n14501) );
  NAND2_X1 U16554 ( .A1(n13251), .A2(n14501), .ZN(n20118) );
  NAND2_X1 U16555 ( .A1(n20120), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n13244) );
  OAI211_X1 U16556 ( .C1(n13257), .C2(n13369), .A(n20118), .B(n13244), .ZN(
        P1_U2950) );
  INV_X1 U16557 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21002) );
  INV_X1 U16558 ( .A(DATAI_10_), .ZN(n13245) );
  MUX2_X1 U16559 ( .A(n13245), .B(n16405), .S(n13593), .Z(n14456) );
  INV_X1 U16560 ( .A(n14456), .ZN(n13246) );
  NAND2_X1 U16561 ( .A1(n13251), .A2(n13246), .ZN(n20112) );
  NAND2_X1 U16562 ( .A1(n20120), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n13247) );
  OAI211_X1 U16563 ( .C1(n13257), .C2(n21002), .A(n20112), .B(n13247), .ZN(
        P1_U2947) );
  INV_X1 U16564 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20936) );
  INV_X1 U16565 ( .A(DATAI_14_), .ZN(n20896) );
  NAND2_X1 U16566 ( .A1(n13593), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13248) );
  OAI21_X1 U16567 ( .B1(n13593), .B2(n20896), .A(n13248), .ZN(n14440) );
  NAND2_X1 U16568 ( .A1(n13251), .A2(n14440), .ZN(n20122) );
  NAND2_X1 U16569 ( .A1(n20120), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13249) );
  OAI211_X1 U16570 ( .C1(n13257), .C2(n20936), .A(n20122), .B(n13249), .ZN(
        P1_U2951) );
  INV_X1 U16571 ( .A(DATAI_11_), .ZN(n20919) );
  NAND2_X1 U16572 ( .A1(n13593), .A2(BUF1_REG_11__SCAN_IN), .ZN(n13250) );
  OAI21_X1 U16573 ( .B1(n13593), .B2(n20919), .A(n13250), .ZN(n14451) );
  NAND2_X1 U16574 ( .A1(n13251), .A2(n14451), .ZN(n20114) );
  NAND2_X1 U16575 ( .A1(n20120), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13252) );
  OAI211_X1 U16576 ( .C1(n13257), .C2(n20890), .A(n20114), .B(n13252), .ZN(
        P1_U2948) );
  INV_X1 U16577 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13815) );
  INV_X1 U16578 ( .A(DATAI_15_), .ZN(n13253) );
  NOR2_X1 U16579 ( .A1(n13593), .A2(n13253), .ZN(n13254) );
  AOI21_X1 U16580 ( .B1(n13593), .B2(BUF1_REG_15__SCAN_IN), .A(n13254), .ZN(
        n13816) );
  INV_X1 U16581 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20081) );
  OAI222_X1 U16582 ( .A1(n13257), .A2(n13815), .B1(n13256), .B2(n13816), .C1(
        n13255), .C2(n20081), .ZN(P1_U2967) );
  INV_X1 U16583 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13266) );
  NOR2_X1 U16584 ( .A1(n13258), .A2(n14204), .ZN(n13259) );
  OAI211_X1 U16585 ( .C1(n13259), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n19107), .B(n13666), .ZN(n13265) );
  NOR2_X1 U16586 ( .A1(n13262), .A2(n13261), .ZN(n13263) );
  NOR2_X1 U16587 ( .A1(n13260), .A2(n13263), .ZN(n19009) );
  NAND2_X1 U16588 ( .A1(n19009), .A2(n19121), .ZN(n13264) );
  OAI211_X1 U16589 ( .C1(n19121), .C2(n13266), .A(n13265), .B(n13264), .ZN(
        P2_U2881) );
  NAND2_X1 U16590 ( .A1(n13268), .A2(n13267), .ZN(n13269) );
  NAND2_X1 U16591 ( .A1(n13270), .A2(n13269), .ZN(n13533) );
  OAI21_X1 U16592 ( .B1(n13272), .B2(n13271), .A(n13365), .ZN(n20136) );
  INV_X1 U16593 ( .A(n20136), .ZN(n13273) );
  AOI22_X1 U16594 ( .A1(n20073), .A2(n13273), .B1(n14437), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13274) );
  OAI21_X1 U16595 ( .B1(n13533), .B2(n14439), .A(n13274), .ZN(P1_U2870) );
  XOR2_X1 U16596 ( .A(n13666), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n13279)
         );
  NOR2_X1 U16597 ( .A1(n13260), .A2(n13275), .ZN(n13276) );
  NOR2_X1 U16598 ( .A1(n16150), .A2(n13276), .ZN(n18999) );
  INV_X1 U16599 ( .A(n18999), .ZN(n15057) );
  MUX2_X1 U16600 ( .A(n13277), .B(n15057), .S(n19121), .Z(n13278) );
  OAI21_X1 U16601 ( .B1(n13279), .B2(n19117), .A(n13278), .ZN(P2_U2880) );
  NOR2_X1 U16602 ( .A1(n13281), .A2(n13282), .ZN(n13280) );
  AND2_X1 U16603 ( .A1(n14502), .A2(n13282), .ZN(n13283) );
  INV_X1 U16604 ( .A(n20158), .ZN(n13284) );
  INV_X1 U16605 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20105) );
  OAI222_X1 U16606 ( .A1(n13523), .A2(n14499), .B1(n14504), .B2(n13284), .C1(
        n14502), .C2(n20105), .ZN(P1_U2903) );
  INV_X1 U16607 ( .A(n20162), .ZN(n13285) );
  INV_X1 U16608 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20103) );
  OAI222_X1 U16609 ( .A1(n13533), .A2(n14499), .B1(n13285), .B2(n14504), .C1(
        n14502), .C2(n20103), .ZN(P1_U2902) );
  XOR2_X1 U16610 ( .A(n19935), .B(n19940), .Z(n13292) );
  OAI21_X1 U16611 ( .B1(n13288), .B2(n13287), .A(n13286), .ZN(n19947) );
  INV_X1 U16612 ( .A(n19947), .ZN(n19056) );
  NAND2_X1 U16613 ( .A1(n19361), .A2(n19056), .ZN(n13289) );
  OAI21_X1 U16614 ( .B1(n19361), .B2(n19056), .A(n13289), .ZN(n19189) );
  NOR2_X1 U16615 ( .A1(n19189), .A2(n19190), .ZN(n19188) );
  INV_X1 U16616 ( .A(n13289), .ZN(n13290) );
  NOR2_X1 U16617 ( .A1(n19188), .A2(n13290), .ZN(n13291) );
  NOR2_X1 U16618 ( .A1(n13291), .A2(n13292), .ZN(n19166) );
  AOI21_X1 U16619 ( .B1(n13292), .B2(n13291), .A(n19166), .ZN(n13296) );
  AOI22_X1 U16620 ( .A1(n13293), .A2(n19187), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19186), .ZN(n13295) );
  NAND2_X1 U16621 ( .A1(n19164), .A2(n16082), .ZN(n13294) );
  OAI211_X1 U16622 ( .C1(n13296), .C2(n19191), .A(n13295), .B(n13294), .ZN(
        P2_U2917) );
  INV_X1 U16623 ( .A(n13523), .ZN(n13300) );
  NAND2_X1 U16624 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13298) );
  OAI211_X1 U16625 ( .C1(n15782), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13298), .B(n13297), .ZN(n13299) );
  AOI21_X1 U16626 ( .B1(n15786), .B2(n13300), .A(n13299), .ZN(n13301) );
  OAI21_X1 U16627 ( .B1(n13302), .B2(n19996), .A(n13301), .ZN(P1_U2998) );
  XNOR2_X1 U16628 ( .A(n13303), .B(n13305), .ZN(n20139) );
  INV_X1 U16629 ( .A(n13533), .ZN(n13308) );
  AOI22_X1 U16630 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13306) );
  OAI21_X1 U16631 ( .B1(n15782), .B2(n13530), .A(n13306), .ZN(n13307) );
  AOI21_X1 U16632 ( .B1(n15786), .B2(n13308), .A(n13307), .ZN(n13309) );
  OAI21_X1 U16633 ( .B1(n19996), .B2(n20139), .A(n13309), .ZN(P1_U2997) );
  INV_X1 U16634 ( .A(n13338), .ZN(n14721) );
  OR2_X1 U16635 ( .A1(n13310), .A2(n14721), .ZN(n13322) );
  INV_X1 U16636 ( .A(n13311), .ZN(n14723) );
  NAND2_X1 U16637 ( .A1(n14723), .A2(n13323), .ZN(n13331) );
  NAND2_X1 U16638 ( .A1(n13311), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13326) );
  NAND2_X1 U16639 ( .A1(n13331), .A2(n13326), .ZN(n13316) );
  INV_X1 U16640 ( .A(n13316), .ZN(n14738) );
  NAND2_X1 U16641 ( .A1(n13328), .A2(n14738), .ZN(n13319) );
  NAND2_X1 U16642 ( .A1(n15506), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13312) );
  NAND2_X1 U16643 ( .A1(n15506), .A2(n10516), .ZN(n14726) );
  MUX2_X1 U16644 ( .A(n13312), .B(n14726), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n13318) );
  INV_X1 U16645 ( .A(n13313), .ZN(n13315) );
  OR2_X1 U16646 ( .A1(n13315), .A2(n13314), .ZN(n13333) );
  NAND2_X1 U16647 ( .A1(n13333), .A2(n13316), .ZN(n13317) );
  OAI211_X1 U16648 ( .C1(n13338), .C2(n13319), .A(n13318), .B(n13317), .ZN(
        n13320) );
  INV_X1 U16649 ( .A(n13320), .ZN(n13321) );
  AND2_X1 U16650 ( .A1(n13322), .A2(n13321), .ZN(n14740) );
  MUX2_X1 U16651 ( .A(n13323), .B(n14740), .S(n15505), .Z(n15518) );
  NOR2_X1 U16652 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20717), .ZN(n13346) );
  INV_X1 U16653 ( .A(n13346), .ZN(n13324) );
  OAI22_X1 U16654 ( .A1(n15518), .A2(P1_STATE2_REG_1__SCAN_IN), .B1(n13324), 
        .B2(n13323), .ZN(n13341) );
  NAND2_X1 U16655 ( .A1(n13326), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13327) );
  NAND2_X1 U16656 ( .A1(n10429), .A2(n13327), .ZN(n20785) );
  NAND2_X1 U16657 ( .A1(n13328), .A2(n20785), .ZN(n13336) );
  NAND2_X1 U16658 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13329) );
  AOI22_X1 U16659 ( .A1(n13330), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n10559), .B2(n13329), .ZN(n13334) );
  XNOR2_X1 U16660 ( .A(n13331), .B(n10559), .ZN(n13332) );
  AOI22_X1 U16661 ( .A1(n15506), .A2(n13334), .B1(n13333), .B2(n13332), .ZN(
        n13335) );
  OAI21_X1 U16662 ( .B1(n13338), .B2(n13336), .A(n13335), .ZN(n13337) );
  NAND2_X1 U16663 ( .A1(n15505), .A2(n20789), .ZN(n13339) );
  OAI21_X1 U16664 ( .B1(n15505), .B2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13339), .ZN(n15523) );
  AOI22_X1 U16665 ( .A1(n15523), .A2(n13324), .B1(P1_STATE2_REG_1__SCAN_IN), 
        .B2(n10559), .ZN(n13340) );
  NAND2_X1 U16666 ( .A1(n13341), .A2(n13340), .ZN(n15534) );
  OR2_X1 U16667 ( .A1(n10560), .A2(n9986), .ZN(n13343) );
  XNOR2_X1 U16668 ( .A(n13343), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20045) );
  NAND2_X1 U16669 ( .A1(n20045), .A2(n15941), .ZN(n13344) );
  NAND2_X1 U16670 ( .A1(n15505), .A2(n13344), .ZN(n13345) );
  OAI211_X1 U16671 ( .C1(n15505), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13345), .B(n20717), .ZN(n13348) );
  NAND2_X1 U16672 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13346), .ZN(
        n13347) );
  AND2_X1 U16673 ( .A1(n13348), .A2(n13347), .ZN(n15532) );
  OAI21_X1 U16674 ( .B1(n15534), .B2(n13342), .A(n15532), .ZN(n13351) );
  OAI21_X1 U16675 ( .B1(n13351), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13349), .ZN(
        n13350) );
  NAND2_X1 U16676 ( .A1(n20721), .A2(n20717), .ZN(n15951) );
  INV_X1 U16677 ( .A(n15951), .ZN(n20804) );
  INV_X1 U16678 ( .A(n15954), .ZN(n15949) );
  NAND2_X1 U16679 ( .A1(n13350), .A2(n20289), .ZN(n20147) );
  NOR2_X1 U16680 ( .A1(n13351), .A2(n15954), .ZN(n15546) );
  INV_X1 U16681 ( .A(n10503), .ZN(n13352) );
  AND2_X1 U16682 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20537), .ZN(n14719) );
  OAI22_X1 U16683 ( .A1(n11527), .A2(n20651), .B1(n13352), .B2(n14719), .ZN(
        n13353) );
  OAI21_X1 U16684 ( .B1(n15546), .B2(n13353), .A(n20147), .ZN(n13354) );
  OAI21_X1 U16685 ( .B1(n20147), .B2(n20570), .A(n13354), .ZN(P1_U3478) );
  INV_X1 U16686 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13391) );
  NOR2_X1 U16687 ( .A1(n13666), .A2(n13391), .ZN(n19109) );
  AND2_X1 U16688 ( .A1(n19109), .A2(n19108), .ZN(n19111) );
  AND2_X1 U16689 ( .A1(n13355), .A2(n19108), .ZN(n13389) );
  NAND2_X1 U16690 ( .A1(n19109), .A2(n13389), .ZN(n19103) );
  OAI211_X1 U16691 ( .C1(n19111), .C2(n13355), .A(n19103), .B(n19107), .ZN(
        n13361) );
  INV_X1 U16692 ( .A(n13357), .ZN(n13358) );
  OAI21_X1 U16693 ( .B1(n13356), .B2(n13359), .A(n13358), .ZN(n18981) );
  INV_X1 U16694 ( .A(n18981), .ZN(n13939) );
  NAND2_X1 U16695 ( .A1(n13939), .A2(n19121), .ZN(n13360) );
  OAI211_X1 U16696 ( .C1(n19121), .C2(n12505), .A(n13361), .B(n13360), .ZN(
        P2_U2878) );
  OAI21_X1 U16697 ( .B1(n13364), .B2(n13363), .A(n13362), .ZN(n13561) );
  OAI21_X1 U16698 ( .B1(n10059), .B2(n9926), .A(n13463), .ZN(n13456) );
  INV_X1 U16699 ( .A(n13456), .ZN(n13366) );
  AOI22_X1 U16700 ( .A1(n20073), .A2(n13366), .B1(n14437), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13367) );
  OAI21_X1 U16701 ( .B1(n13561), .B2(n14439), .A(n13367), .ZN(P1_U2869) );
  AOI22_X1 U16702 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13368) );
  OAI21_X1 U16703 ( .B1(n13369), .B2(n13375), .A(n13368), .ZN(P1_U2907) );
  AOI22_X1 U16704 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U16705 ( .B1(n13778), .B2(n13375), .A(n13370), .ZN(P1_U2920) );
  AOI22_X1 U16706 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13371) );
  OAI21_X1 U16707 ( .B1(n21002), .B2(n13375), .A(n13371), .ZN(P1_U2910) );
  INV_X1 U16708 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13373) );
  AOI22_X1 U16709 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13372) );
  OAI21_X1 U16710 ( .B1(n13373), .B2(n13375), .A(n13372), .ZN(P1_U2919) );
  AOI22_X1 U16711 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20801), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n15566), .ZN(n13374) );
  OAI21_X1 U16712 ( .B1(n20936), .B2(n13375), .A(n13374), .ZN(P1_U2906) );
  XNOR2_X1 U16713 ( .A(n13376), .B(n13377), .ZN(n13566) );
  INV_X1 U16714 ( .A(n20133), .ZN(n13378) );
  NOR2_X1 U16715 ( .A1(n15886), .A2(n13378), .ZN(n13379) );
  OR2_X1 U16716 ( .A1(n13380), .A2(n13379), .ZN(n13552) );
  INV_X1 U16717 ( .A(n13622), .ZN(n15881) );
  NAND2_X1 U16718 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13381) );
  AOI21_X1 U16719 ( .B1(n15881), .B2(n13381), .A(n13619), .ZN(n20145) );
  OAI21_X1 U16720 ( .B1(n15886), .B2(n20133), .A(n20145), .ZN(n13549) );
  NAND2_X1 U16721 ( .A1(n13549), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13382) );
  NAND2_X1 U16722 ( .A1(n15935), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13559) );
  OAI211_X1 U16723 ( .C1(n20137), .C2(n13456), .A(n13382), .B(n13559), .ZN(
        n13383) );
  AOI21_X1 U16724 ( .B1(n13384), .B2(n13552), .A(n13383), .ZN(n13385) );
  OAI21_X1 U16725 ( .B1(n20138), .B2(n13566), .A(n13385), .ZN(P1_U3028) );
  OAI21_X1 U16726 ( .B1(n19103), .B2(n13387), .A(n13386), .ZN(n13393) );
  AND2_X1 U16727 ( .A1(n19102), .A2(n13388), .ZN(n13390) );
  NAND2_X1 U16728 ( .A1(n13390), .A2(n13389), .ZN(n13392) );
  OR2_X1 U16729 ( .A1(n13666), .A2(n13540), .ZN(n19097) );
  NAND3_X1 U16730 ( .A1(n13393), .A2(n19107), .A3(n19097), .ZN(n13398) );
  NOR2_X1 U16731 ( .A1(n13394), .A2(n13395), .ZN(n13396) );
  NOR2_X1 U16732 ( .A1(n13916), .A2(n13396), .ZN(n18947) );
  NAND2_X1 U16733 ( .A1(n18947), .A2(n19121), .ZN(n13397) );
  OAI211_X1 U16734 ( .C1(n19121), .C2(n13399), .A(n13398), .B(n13397), .ZN(
        P2_U2876) );
  NOR2_X1 U16735 ( .A1(n19097), .A2(n19098), .ZN(n13402) );
  OR2_X1 U16736 ( .A1(n13400), .A2(n19098), .ZN(n13539) );
  OR2_X1 U16737 ( .A1(n19097), .A2(n13539), .ZN(n19092) );
  OAI211_X1 U16738 ( .C1(n13402), .C2(n13401), .A(n19092), .B(n19107), .ZN(
        n13406) );
  NOR2_X1 U16739 ( .A1(n13918), .A2(n13403), .ZN(n13404) );
  NOR2_X1 U16740 ( .A1(n16103), .A2(n13404), .ZN(n18935) );
  NAND2_X1 U16741 ( .A1(n18935), .A2(n19121), .ZN(n13405) );
  OAI211_X1 U16742 ( .C1(n19121), .C2(n12518), .A(n13406), .B(n13405), .ZN(
        P2_U2874) );
  INV_X1 U16743 ( .A(n14716), .ZN(n13407) );
  NOR2_X1 U16744 ( .A1(n20500), .A2(n20651), .ZN(n13414) );
  AND2_X1 U16745 ( .A1(n20658), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13409) );
  NAND2_X1 U16746 ( .A1(n20220), .A2(n13409), .ZN(n14717) );
  NOR2_X1 U16747 ( .A1(n20368), .A2(n14717), .ZN(n20374) );
  INV_X1 U16748 ( .A(n13409), .ZN(n13410) );
  OR2_X1 U16749 ( .A1(n20220), .A2(n13410), .ZN(n13411) );
  NOR2_X1 U16750 ( .A1(n20649), .A2(n13411), .ZN(n20574) );
  NAND2_X1 U16751 ( .A1(n20658), .A2(n21127), .ZN(n20527) );
  OAI22_X1 U16752 ( .A1(n13589), .A2(n20527), .B1(n13412), .B2(n14719), .ZN(
        n13413) );
  OR4_X1 U16753 ( .A1(n13414), .A2(n20374), .A3(n20574), .A4(n13413), .ZN(
        n13415) );
  NAND2_X1 U16754 ( .A1(n20147), .A2(n13415), .ZN(n13416) );
  OAI21_X1 U16755 ( .B1(n20147), .B2(n20489), .A(n13416), .ZN(P1_U3475) );
  INV_X1 U16756 ( .A(n20169), .ZN(n13417) );
  INV_X1 U16757 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20101) );
  OAI222_X1 U16758 ( .A1(n13561), .A2(n14499), .B1(n13417), .B2(n14504), .C1(
        n14502), .C2(n20101), .ZN(P1_U2901) );
  INV_X1 U16759 ( .A(n20151), .ZN(n13418) );
  INV_X1 U16760 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20109) );
  OAI222_X1 U16761 ( .A1(n20132), .A2(n14499), .B1(n13418), .B2(n14504), .C1(
        n14502), .C2(n20109), .ZN(P1_U2904) );
  XNOR2_X1 U16762 ( .A(n13420), .B(n13419), .ZN(n13421) );
  XNOR2_X1 U16763 ( .A(n13422), .B(n13421), .ZN(n16247) );
  XNOR2_X1 U16764 ( .A(n13424), .B(n13423), .ZN(n16245) );
  AOI21_X1 U16765 ( .B1(n13504), .B2(n13472), .A(n15487), .ZN(n15485) );
  OAI22_X1 U16766 ( .A1(n16179), .A2(n13504), .B1(n13425), .B2(n16232), .ZN(
        n13426) );
  AOI21_X1 U16767 ( .B1(n16170), .B2(n15485), .A(n13426), .ZN(n13428) );
  NAND2_X1 U16768 ( .A1(n13099), .A2(n19250), .ZN(n13427) );
  OAI211_X1 U16769 ( .C1(n16245), .C2(n16172), .A(n13428), .B(n13427), .ZN(
        n13429) );
  INV_X1 U16770 ( .A(n13429), .ZN(n13430) );
  OAI21_X1 U16771 ( .B1(n16247), .B2(n16173), .A(n13430), .ZN(P2_U3011) );
  NOR2_X1 U16772 ( .A1(n20537), .A2(n15951), .ZN(n15545) );
  AOI211_X1 U16773 ( .C1(P1_STATE2_REG_0__SCAN_IN), .C2(n15545), .A(n15899), 
        .B(n20798), .ZN(n13434) );
  AND2_X1 U16774 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20718), .ZN(n13431) );
  NAND2_X1 U16775 ( .A1(n13432), .A2(n13431), .ZN(n13433) );
  NAND2_X1 U16776 ( .A1(n13435), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13437) );
  INV_X1 U16777 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13436) );
  XNOR2_X1 U16778 ( .A(n13437), .B(n13436), .ZN(n13980) );
  NOR2_X1 U16779 ( .A1(n13980), .A2(n20717), .ZN(n13438) );
  AND2_X1 U16780 ( .A1(n13439), .A2(n20798), .ZN(n13440) );
  OR2_X1 U16781 ( .A1(n20025), .A2(n13440), .ZN(n20041) );
  AND2_X1 U16782 ( .A1(n13980), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13441) );
  AND2_X1 U16783 ( .A1(n13442), .A2(n20798), .ZN(n20065) );
  AND2_X1 U16784 ( .A1(n9827), .A2(n20798), .ZN(n13449) );
  AND2_X1 U16785 ( .A1(n13447), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13444) );
  NAND2_X1 U16786 ( .A1(n20800), .A2(n21127), .ZN(n13445) );
  INV_X1 U16787 ( .A(n13444), .ZN(n13448) );
  INV_X1 U16788 ( .A(n13445), .ZN(n13446) );
  OAI21_X1 U16789 ( .B1(n13447), .B2(n15537), .A(n13446), .ZN(n13450) );
  INV_X1 U16790 ( .A(n13449), .ZN(n13451) );
  NAND3_X1 U16791 ( .A1(n15644), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .ZN(n13453) );
  NOR2_X1 U16792 ( .A1(n15630), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13525) );
  OAI21_X1 U16793 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n15630), .A(n15629), .ZN(
        n13524) );
  OAI21_X1 U16794 ( .B1(n13525), .B2(n13524), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n13452) );
  OAI21_X1 U16795 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(n13453), .A(n13452), .ZN(
        n13454) );
  AOI21_X1 U16796 ( .B1(n20046), .B2(P1_EBX_REG_3__SCAN_IN), .A(n13454), .ZN(
        n13455) );
  OAI21_X1 U16797 ( .B1(n13456), .B2(n20049), .A(n13455), .ZN(n13457) );
  OAI21_X1 U16798 ( .B1(n20064), .B2(n13560), .A(n9908), .ZN(n13458) );
  AOI21_X1 U16799 ( .B1(n13564), .B2(n20053), .A(n13458), .ZN(n13459) );
  OAI21_X1 U16800 ( .B1(n20071), .B2(n13561), .A(n13459), .ZN(P1_U2837) );
  NAND2_X1 U16801 ( .A1(n13362), .A2(n13460), .ZN(n13461) );
  AND2_X1 U16802 ( .A1(n13568), .A2(n13461), .ZN(n20042) );
  INV_X1 U16803 ( .A(n20042), .ZN(n13467) );
  AND2_X1 U16804 ( .A1(n13463), .A2(n13462), .ZN(n13464) );
  NOR2_X1 U16805 ( .A1(n9915), .A2(n13464), .ZN(n20044) );
  AOI22_X1 U16806 ( .A1(n20073), .A2(n20044), .B1(n14437), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13465) );
  OAI21_X1 U16807 ( .B1(n13467), .B2(n14439), .A(n13465), .ZN(P1_U2868) );
  INV_X1 U16808 ( .A(n14483), .ZN(n13466) );
  INV_X1 U16809 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20099) );
  OAI222_X1 U16810 ( .A1(n13467), .A2(n14499), .B1(n13466), .B2(n14504), .C1(
        n14502), .C2(n20099), .ZN(P1_U2900) );
  INV_X1 U16811 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14906) );
  INV_X1 U16812 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13468) );
  INV_X1 U16813 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13969) );
  INV_X1 U16814 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U16815 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12056), .B1(n13471), 
        .B2(n13470), .ZN(n19078) );
  AOI22_X1 U16816 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13894), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n13470), .ZN(n13695) );
  NOR2_X1 U16817 ( .A1(n19078), .A2(n13695), .ZN(n13694) );
  NOR2_X1 U16818 ( .A1(n10004), .A2(n13694), .ZN(n13473) );
  OAI21_X1 U16819 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13472), .ZN(n19248) );
  XNOR2_X1 U16820 ( .A(n13473), .B(n19248), .ZN(n13496) );
  NOR4_X4 U16821 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .A4(n13474), .ZN(n19058) );
  OR2_X1 U16822 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19980), .ZN(n13487) );
  OR3_X1 U16823 ( .A1(n19974), .A2(n13489), .A3(n13487), .ZN(n19046) );
  NAND2_X1 U16824 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19979), .ZN(n19303) );
  NOR2_X1 U16825 ( .A1(n13475), .A2(n19303), .ZN(n16265) );
  OR2_X1 U16826 ( .A1(n19016), .A2(n19058), .ZN(n13476) );
  NOR2_X1 U16827 ( .A1(n16265), .A2(n13476), .ZN(n13477) );
  AND2_X2 U16828 ( .A1(n19974), .A2(n13477), .ZN(n19053) );
  INV_X1 U16829 ( .A(n13487), .ZN(n13478) );
  NOR2_X1 U16830 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13478), .ZN(n13479) );
  AND2_X1 U16831 ( .A1(n13480), .A2(n13479), .ZN(n13481) );
  OR2_X1 U16832 ( .A1(n13486), .A2(n13481), .ZN(n13484) );
  NOR2_X1 U16833 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13482), .ZN(n16311) );
  INV_X1 U16834 ( .A(n16311), .ZN(n13483) );
  AND2_X2 U16835 ( .A1(n13484), .A2(n13483), .ZN(n19047) );
  INV_X1 U16836 ( .A(n19047), .ZN(n19065) );
  INV_X1 U16837 ( .A(n19053), .ZN(n19067) );
  OAI22_X1 U16838 ( .A1(n13485), .A2(n19065), .B1(n12075), .B2(n19067), .ZN(
        n13492) );
  NAND2_X1 U16839 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13487), .ZN(n13488) );
  OR3_X1 U16840 ( .A1(n19974), .A2(n13489), .A3(n13488), .ZN(n19072) );
  OAI22_X1 U16841 ( .A1(n19935), .A2(n19055), .B1(n13490), .B2(n19072), .ZN(
        n13491) );
  AOI211_X1 U16842 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19081), .A(
        n13492), .B(n13491), .ZN(n13494) );
  NAND2_X1 U16843 ( .A1(n19940), .A2(n19077), .ZN(n13493) );
  OAI211_X1 U16844 ( .C1(n16283), .C2(n19046), .A(n13494), .B(n13493), .ZN(
        n13495) );
  AOI21_X1 U16845 ( .B1(n13496), .B2(n19058), .A(n13495), .ZN(n13497) );
  INV_X1 U16846 ( .A(n13497), .ZN(P2_U2853) );
  INV_X1 U16847 ( .A(n19077), .ZN(n13512) );
  NAND2_X1 U16848 ( .A1(n13694), .A2(n19248), .ZN(n15484) );
  NAND2_X1 U16849 ( .A1(n10005), .A2(n15484), .ZN(n13498) );
  XNOR2_X1 U16850 ( .A(n15485), .B(n13498), .ZN(n13499) );
  NAND2_X1 U16851 ( .A1(n13499), .A2(n19058), .ZN(n13511) );
  OAI21_X1 U16852 ( .B1(n13502), .B2(n13501), .A(n13500), .ZN(n19167) );
  OAI22_X1 U16853 ( .A1(n13504), .A2(n19049), .B1(n13503), .B2(n19072), .ZN(
        n13505) );
  INV_X1 U16854 ( .A(n13505), .ZN(n13506) );
  OAI21_X1 U16855 ( .B1(n19055), .B2(n19167), .A(n13506), .ZN(n13509) );
  OAI22_X1 U16856 ( .A1(n13507), .A2(n19065), .B1(n13425), .B2(n19067), .ZN(
        n13508) );
  AOI211_X1 U16857 ( .C1(n19075), .C2(n13099), .A(n13509), .B(n13508), .ZN(
        n13510) );
  OAI211_X1 U16858 ( .C1(n13512), .C2(n19925), .A(n13511), .B(n13510), .ZN(
        P2_U2852) );
  INV_X1 U16859 ( .A(n15629), .ZN(n14332) );
  INV_X1 U16860 ( .A(n20065), .ZN(n13518) );
  INV_X1 U16861 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20904) );
  AOI22_X1 U16862 ( .A1(n15644), .A2(n20904), .B1(n20046), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13517) );
  NAND2_X1 U16863 ( .A1(n13515), .A2(n20067), .ZN(n13516) );
  OAI211_X1 U16864 ( .C1(n13514), .C2(n13518), .A(n13517), .B(n13516), .ZN(
        n13519) );
  AOI21_X1 U16865 ( .B1(n14332), .B2(P1_REIP_REG_1__SCAN_IN), .A(n13519), .ZN(
        n13520) );
  OAI21_X1 U16866 ( .B1(n20063), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13520), .ZN(n13521) );
  AOI21_X1 U16867 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20024), .A(
        n13521), .ZN(n13522) );
  OAI21_X1 U16868 ( .B1(n20071), .B2(n13523), .A(n13522), .ZN(P1_U2839) );
  AOI22_X1 U16869 ( .A1(n20061), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n13524), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n13527) );
  NAND2_X1 U16870 ( .A1(n13525), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13526) );
  OAI211_X1 U16871 ( .C1(n20136), .C2(n20049), .A(n13527), .B(n13526), .ZN(
        n13528) );
  AOI21_X1 U16872 ( .B1(n9981), .B2(n20065), .A(n13528), .ZN(n13529) );
  OAI21_X1 U16873 ( .B1(n20063), .B2(n13530), .A(n13529), .ZN(n13531) );
  AOI21_X1 U16874 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n20024), .A(
        n13531), .ZN(n13532) );
  OAI21_X1 U16875 ( .B1(n20071), .B2(n13533), .A(n13532), .ZN(P1_U2838) );
  XNOR2_X1 U16876 ( .A(n13534), .B(n13535), .ZN(n13558) );
  NAND2_X1 U16877 ( .A1(n15935), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n13551) );
  NAND2_X1 U16878 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13536) );
  OAI211_X1 U16879 ( .C1(n15782), .C2(n20043), .A(n13551), .B(n13536), .ZN(
        n13537) );
  AOI21_X1 U16880 ( .B1(n20042), .B2(n15786), .A(n13537), .ZN(n13538) );
  OAI21_X1 U16881 ( .B1(n13558), .B2(n19996), .A(n13538), .ZN(P1_U2995) );
  OR2_X1 U16882 ( .A1(n13539), .A2(n19093), .ZN(n13541) );
  NOR2_X1 U16883 ( .A1(n13666), .A2(n13663), .ZN(n19086) );
  INV_X1 U16884 ( .A(n19086), .ZN(n13544) );
  OAI211_X1 U16885 ( .C1(n10232), .C2(n13545), .A(n13544), .B(n19107), .ZN(
        n13548) );
  OAI21_X1 U16886 ( .B1(n16102), .B2(n13546), .A(n15031), .ZN(n15047) );
  INV_X1 U16887 ( .A(n15047), .ZN(n18916) );
  NAND2_X1 U16888 ( .A1(n18916), .A2(n19121), .ZN(n13547) );
  OAI211_X1 U16889 ( .C1(n19121), .C2(n12524), .A(n13548), .B(n13547), .ZN(
        P2_U2872) );
  NAND2_X1 U16890 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13549), .ZN(
        n13550) );
  NAND2_X1 U16891 ( .A1(n13551), .A2(n13550), .ZN(n13556) );
  INV_X1 U16892 ( .A(n13552), .ZN(n13554) );
  AOI211_X1 U16893 ( .C1(n11550), .C2(n13384), .A(n13554), .B(n13553), .ZN(
        n13555) );
  AOI211_X1 U16894 ( .C1(n15932), .C2(n20044), .A(n13556), .B(n13555), .ZN(
        n13557) );
  OAI21_X1 U16895 ( .B1(n20138), .B2(n13558), .A(n13557), .ZN(P1_U3027) );
  OAI21_X1 U16896 ( .B1(n15790), .B2(n13560), .A(n13559), .ZN(n13563) );
  NOR2_X1 U16897 ( .A1(n13561), .A2(n20131), .ZN(n13562) );
  AOI211_X1 U16898 ( .C1(n15783), .C2(n13564), .A(n13563), .B(n13562), .ZN(
        n13565) );
  OAI21_X1 U16899 ( .B1(n19996), .B2(n13566), .A(n13565), .ZN(P1_U2996) );
  AOI21_X1 U16900 ( .B1(n13569), .B2(n13568), .A(n13567), .ZN(n15785) );
  INV_X1 U16901 ( .A(n15785), .ZN(n20034) );
  INV_X1 U16902 ( .A(n20175), .ZN(n13570) );
  INV_X1 U16903 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n20097) );
  OAI222_X1 U16904 ( .A1(n20034), .A2(n14499), .B1(n13570), .B2(n14504), .C1(
        n14502), .C2(n20097), .ZN(P1_U2899) );
  NOR2_X1 U16905 ( .A1(n13025), .A2(n19916), .ZN(n13575) );
  NAND2_X1 U16906 ( .A1(n13571), .A2(n12576), .ZN(n13689) );
  MUX2_X1 U16907 ( .A(n13689), .B(n15313), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13572) );
  AOI21_X1 U16908 ( .B1(n19076), .B2(n15306), .A(n13572), .ZN(n16290) );
  INV_X1 U16909 ( .A(n19831), .ZN(n19922) );
  OAI22_X1 U16910 ( .A1(n15967), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19078), .B2(n10004), .ZN(n13696) );
  INV_X1 U16911 ( .A(n13696), .ZN(n13573) );
  OAI22_X1 U16912 ( .A1(n16290), .A2(n19922), .B1(n13474), .B2(n13573), .ZN(
        n13574) );
  OAI21_X1 U16913 ( .B1(n13575), .B2(n13574), .A(n13578), .ZN(n13576) );
  OAI21_X1 U16914 ( .B1(n13578), .B2(n13577), .A(n13576), .ZN(P2_U3601) );
  NOR2_X1 U16915 ( .A1(n9915), .A2(n13579), .ZN(n13580) );
  OR2_X1 U16916 ( .A1(n15930), .A2(n13580), .ZN(n20030) );
  INV_X1 U16917 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n21157) );
  OAI222_X1 U16918 ( .A1(n20030), .A2(n15712), .B1(n20078), .B2(n21157), .C1(
        n14439), .C2(n20034), .ZN(P1_U2867) );
  NOR2_X1 U16919 ( .A1(n13581), .A2(n13630), .ZN(n13629) );
  INV_X1 U16920 ( .A(n13582), .ZN(n13583) );
  OAI21_X1 U16921 ( .B1(n13629), .B2(n13584), .A(n13583), .ZN(n13764) );
  AOI22_X1 U16922 ( .A1(n13772), .A2(n14465), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14487), .ZN(n13585) );
  OAI21_X1 U16923 ( .B1(n13764), .B2(n14499), .A(n13585), .ZN(P1_U2896) );
  AND2_X1 U16924 ( .A1(n13700), .A2(n13586), .ZN(n13587) );
  OR2_X1 U16925 ( .A1(n13587), .A2(n13641), .ZN(n13706) );
  INV_X1 U16926 ( .A(n13706), .ZN(n15918) );
  AOI22_X1 U16927 ( .A1(n20073), .A2(n15918), .B1(n14437), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n13588) );
  OAI21_X1 U16928 ( .B1(n13764), .B2(n14439), .A(n13588), .ZN(P1_U2864) );
  INV_X1 U16929 ( .A(n11527), .ZN(n13590) );
  OAI21_X1 U16930 ( .B1(n20216), .B2(n20692), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n13591) );
  NAND2_X1 U16931 ( .A1(n13591), .A2(n20658), .ZN(n13602) );
  INV_X1 U16932 ( .A(n13514), .ZN(n20598) );
  OR2_X1 U16933 ( .A1(n20254), .A2(n20598), .ZN(n13597) );
  INV_X1 U16934 ( .A(n20401), .ZN(n13592) );
  NAND2_X1 U16935 ( .A1(n13592), .A2(n20456), .ZN(n20285) );
  NOR2_X1 U16936 ( .A1(n13598), .A2(n20721), .ZN(n20458) );
  INV_X1 U16937 ( .A(n20458), .ZN(n20402) );
  OAI22_X1 U16938 ( .A1(n13602), .A2(n13597), .B1(n20285), .B2(n20402), .ZN(
        n20187) );
  INV_X1 U16939 ( .A(n20187), .ZN(n13615) );
  NAND2_X1 U16940 ( .A1(n20196), .A2(n14483), .ZN(n20682) );
  INV_X1 U16941 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16389) );
  INV_X1 U16942 ( .A(DATAI_20_), .ZN(n21003) );
  OAI22_X1 U16943 ( .A1(n16389), .A2(n20184), .B1(n21003), .B2(n20186), .ZN(
        n20509) );
  INV_X1 U16944 ( .A(n20179), .ZN(n13609) );
  NAND2_X1 U16945 ( .A1(n13609), .A2(n13596), .ZN(n20683) );
  NAND3_X1 U16946 ( .A1(n20489), .A2(n15515), .A3(n20531), .ZN(n20195) );
  NOR2_X1 U16947 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20195), .ZN(
        n20182) );
  INV_X1 U16948 ( .A(n20182), .ZN(n13610) );
  INV_X1 U16949 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16379) );
  INV_X1 U16950 ( .A(DATAI_28_), .ZN(n21166) );
  OAI22_X2 U16951 ( .A1(n16379), .A2(n20184), .B1(n21166), .B2(n20186), .ZN(
        n20685) );
  INV_X1 U16952 ( .A(n20685), .ZN(n20512) );
  OAI22_X1 U16953 ( .A1(n20683), .A2(n13610), .B1(n20715), .B2(n20512), .ZN(
        n13606) );
  INV_X1 U16954 ( .A(n13597), .ZN(n13601) );
  NAND2_X1 U16955 ( .A1(n13598), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20600) );
  NAND2_X1 U16956 ( .A1(n20196), .A2(n20600), .ZN(n20403) );
  AOI21_X1 U16957 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n13610), .A(n20403), 
        .ZN(n13600) );
  NAND2_X1 U16958 ( .A1(n20285), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13599) );
  OAI211_X1 U16959 ( .C1(n13602), .C2(n13601), .A(n13600), .B(n13599), .ZN(
        n13603) );
  NOR2_X1 U16960 ( .A1(n20191), .A2(n13604), .ZN(n13605) );
  AOI211_X1 U16961 ( .C1(n20216), .C2(n20509), .A(n13606), .B(n13605), .ZN(
        n13607) );
  OAI21_X1 U16962 ( .B1(n13615), .B2(n20682), .A(n13607), .ZN(P1_U3037) );
  NAND2_X1 U16963 ( .A1(n20196), .A2(n14469), .ZN(n20706) );
  INV_X1 U16964 ( .A(DATAI_23_), .ZN(n21122) );
  INV_X1 U16965 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16385) );
  OAI22_X1 U16966 ( .A1(n21122), .A2(n20186), .B1(n16385), .B2(n20184), .ZN(
        n20520) );
  NAND2_X1 U16967 ( .A1(n13609), .A2(n13608), .ZN(n20708) );
  INV_X1 U16968 ( .A(DATAI_31_), .ZN(n20957) );
  INV_X1 U16969 ( .A(n20710), .ZN(n20525) );
  OAI22_X1 U16970 ( .A1(n20708), .A2(n13610), .B1(n20715), .B2(n20525), .ZN(
        n13613) );
  NOR2_X1 U16971 ( .A1(n20191), .A2(n13611), .ZN(n13612) );
  AOI211_X1 U16972 ( .C1(n20216), .C2(n20520), .A(n13613), .B(n13612), .ZN(
        n13614) );
  OAI21_X1 U16973 ( .B1(n13615), .B2(n20706), .A(n13614), .ZN(P1_U3040) );
  XOR2_X1 U16974 ( .A(n13616), .B(n13617), .Z(n15787) );
  INV_X1 U16975 ( .A(n15787), .ZN(n13628) );
  NOR2_X1 U16976 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13618), .ZN(
        n13737) );
  INV_X1 U16977 ( .A(n13737), .ZN(n13627) );
  AOI21_X1 U16978 ( .B1(n20143), .B2(n13620), .A(n13619), .ZN(n15885) );
  OAI21_X1 U16979 ( .B1(n13622), .B2(n13621), .A(n15885), .ZN(n13735) );
  NOR3_X1 U16980 ( .A1(n15886), .A2(n13623), .A3(n15817), .ZN(n13625) );
  NAND2_X1 U16981 ( .A1(n15935), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15788) );
  OAI21_X1 U16982 ( .B1(n20137), .B2(n20030), .A(n15788), .ZN(n13624) );
  AOI211_X1 U16983 ( .C1(n13735), .C2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13625), .B(n13624), .ZN(n13626) );
  OAI211_X1 U16984 ( .C1(n13628), .C2(n20138), .A(n13627), .B(n13626), .ZN(
        P1_U3026) );
  AOI21_X1 U16985 ( .B1(n13630), .B2(n13581), .A(n13629), .ZN(n20017) );
  INV_X1 U16986 ( .A(n20017), .ZN(n13703) );
  INV_X1 U16987 ( .A(n14469), .ZN(n13631) );
  OAI222_X1 U16988 ( .A1(n13703), .A2(n14499), .B1(n13631), .B2(n14504), .C1(
        n14502), .C2(n10659), .ZN(P1_U2897) );
  XOR2_X1 U16989 ( .A(n13567), .B(n13632), .Z(n20075) );
  INV_X1 U16990 ( .A(n20075), .ZN(n13634) );
  INV_X1 U16991 ( .A(n20183), .ZN(n13633) );
  OAI222_X1 U16992 ( .A1(n14499), .A2(n13634), .B1(n13633), .B2(n14504), .C1(
        n14502), .C2(n10651), .ZN(P1_U2898) );
  NOR2_X1 U16993 ( .A1(n13582), .A2(n13636), .ZN(n13637) );
  OR2_X1 U16994 ( .A1(n13635), .A2(n13637), .ZN(n13784) );
  AOI22_X1 U16995 ( .A1(n13772), .A2(n14462), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14487), .ZN(n13638) );
  OAI21_X1 U16996 ( .B1(n13784), .B2(n14499), .A(n13638), .ZN(P1_U2895) );
  NAND4_X1 U16997 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .A4(P1_REIP_REG_6__SCAN_IN), .ZN(n13805)
         );
  NAND3_X1 U16998 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n13639) );
  NOR2_X1 U16999 ( .A1(n15630), .A2(n13639), .ZN(n20040) );
  NAND2_X1 U17000 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20040), .ZN(n15677) );
  NOR2_X1 U17001 ( .A1(n13805), .A2(n15677), .ZN(n14399) );
  INV_X1 U17002 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n21029) );
  NAND2_X1 U17003 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13650) );
  NAND2_X1 U17004 ( .A1(n20053), .A2(n13787), .ZN(n13649) );
  NOR2_X1 U17005 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  OR2_X1 U17006 ( .A1(n13747), .A2(n13642), .ZN(n13793) );
  NAND4_X1 U17007 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n13831)
         );
  NOR3_X1 U17008 ( .A1(n14332), .A2(n13831), .A3(n13805), .ZN(n13745) );
  NAND2_X1 U17009 ( .A1(n15629), .A2(n15630), .ZN(n20062) );
  NAND2_X1 U17010 ( .A1(n20062), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n13643) );
  OR2_X1 U17011 ( .A1(n13745), .A2(n13643), .ZN(n13645) );
  NAND2_X1 U17012 ( .A1(n20046), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n13644) );
  AND2_X1 U17013 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  OAI21_X1 U17014 ( .B1(n20049), .B2(n13793), .A(n13646), .ZN(n13647) );
  INV_X1 U17015 ( .A(n13647), .ZN(n13648) );
  NAND4_X1 U17016 ( .A1(n13650), .A2(n13649), .A3(n20135), .A4(n13648), .ZN(
        n13651) );
  AOI21_X1 U17017 ( .B1(n14399), .B2(n21029), .A(n13651), .ZN(n13652) );
  OAI21_X1 U17018 ( .B1(n15623), .B2(n13784), .A(n13652), .ZN(P1_U2831) );
  AOI22_X1 U17019 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12149), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13656) );
  AOI22_X1 U17020 ( .A1(n9816), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13655) );
  AOI22_X1 U17021 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13654) );
  AOI22_X1 U17022 ( .A1(n14079), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13653) );
  NAND4_X1 U17023 ( .A1(n13656), .A2(n13655), .A3(n13654), .A4(n13653), .ZN(
        n13662) );
  AOI22_X1 U17024 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12155), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13660) );
  AOI22_X1 U17025 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13659) );
  AOI22_X1 U17026 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13658) );
  AOI22_X1 U17027 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13657) );
  NAND4_X1 U17028 ( .A1(n13660), .A2(n13659), .A3(n13658), .A4(n13657), .ZN(
        n13661) );
  INV_X1 U17029 ( .A(n19085), .ZN(n13664) );
  AOI22_X1 U17030 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13670) );
  AOI22_X1 U17031 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n9815), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13669) );
  AOI22_X1 U17032 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13668) );
  AOI22_X1 U17033 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13667) );
  NAND4_X1 U17034 ( .A1(n13670), .A2(n13669), .A3(n13668), .A4(n13667), .ZN(
        n13676) );
  AOI22_X1 U17035 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13674) );
  AOI22_X1 U17036 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13673) );
  AOI22_X1 U17037 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13672) );
  AOI22_X1 U17038 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13671) );
  NAND4_X1 U17039 ( .A1(n13674), .A2(n13673), .A3(n13672), .A4(n13671), .ZN(
        n13675) );
  OAI21_X1 U17040 ( .B1(n13677), .B2(n13678), .A(n14000), .ZN(n14808) );
  AND2_X1 U17041 ( .A1(n15222), .A2(n13680), .ZN(n13681) );
  NOR2_X1 U17042 ( .A1(n13679), .A2(n13681), .ZN(n18895) );
  OAI22_X1 U17043 ( .A1(n14884), .A2(n19269), .B1(n19162), .B2(n13682), .ZN(
        n13687) );
  INV_X1 U17044 ( .A(n19127), .ZN(n14888) );
  INV_X1 U17045 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n13685) );
  INV_X1 U17046 ( .A(n19126), .ZN(n14886) );
  INV_X1 U17047 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13684) );
  OAI22_X1 U17048 ( .A1(n14888), .A2(n13685), .B1(n14886), .B2(n13684), .ZN(
        n13686) );
  AOI211_X1 U17049 ( .C1(n19187), .C2(n18895), .A(n13687), .B(n13686), .ZN(
        n13688) );
  OAI21_X1 U17050 ( .B1(n14808), .B2(n19191), .A(n13688), .ZN(P2_U2902) );
  OAI21_X1 U17051 ( .B1(n13691), .B2(n13690), .A(n13689), .ZN(n13693) );
  NAND2_X1 U17052 ( .A1(n15313), .A2(n11851), .ZN(n13692) );
  OAI211_X1 U17053 ( .C1(n13910), .C2(n16282), .A(n13693), .B(n13692), .ZN(
        n16292) );
  AOI211_X1 U17054 ( .C1(n19078), .C2(n13695), .A(n10004), .B(n13694), .ZN(
        n19059) );
  AOI21_X1 U17055 ( .B1(n10004), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n19059), .ZN(n19914) );
  NOR2_X1 U17056 ( .A1(n13474), .A2(n13696), .ZN(n19912) );
  INV_X1 U17057 ( .A(n19916), .ZN(n13697) );
  AOI222_X1 U17058 ( .A1(n16292), .A2(n19831), .B1(n19914), .B2(n19912), .C1(
        n13697), .C2(n19943), .ZN(n13699) );
  NAND2_X1 U17059 ( .A1(n19918), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13698) );
  OAI21_X1 U17060 ( .B1(n19918), .B2(n13699), .A(n13698), .ZN(P2_U3600) );
  INV_X1 U17061 ( .A(n13700), .ZN(n13701) );
  AOI21_X1 U17062 ( .B1(n13702), .B2(n15928), .A(n13701), .ZN(n20012) );
  INV_X1 U17063 ( .A(n20012), .ZN(n13738) );
  INV_X1 U17064 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13704) );
  OAI222_X1 U17065 ( .A1(n13738), .A2(n15712), .B1(n20078), .B2(n13704), .C1(
        n14439), .C2(n13703), .ZN(P1_U2865) );
  INV_X1 U17066 ( .A(n13764), .ZN(n13715) );
  NAND2_X1 U17067 ( .A1(n20062), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n13711) );
  AOI21_X1 U17068 ( .B1(n20046), .B2(P1_EBX_REG_8__SCAN_IN), .A(n15899), .ZN(
        n13705) );
  OAI21_X1 U17069 ( .B1(n13706), .B2(n20049), .A(n13705), .ZN(n13707) );
  AOI21_X1 U17070 ( .B1(n20024), .B2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n13707), .ZN(n13710) );
  INV_X1 U17071 ( .A(n13760), .ZN(n13708) );
  NAND2_X1 U17072 ( .A1(n20053), .A2(n13708), .ZN(n13709) );
  OAI211_X1 U17073 ( .C1(n13745), .C2(n13711), .A(n13710), .B(n13709), .ZN(
        n13714) );
  NAND3_X1 U17074 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .ZN(n13712) );
  NOR3_X1 U17075 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13712), .A3(n15677), .ZN(
        n13713) );
  AOI211_X1 U17076 ( .C1(n13715), .C2(n20025), .A(n13714), .B(n13713), .ZN(
        n13716) );
  INV_X1 U17077 ( .A(n13716), .ZN(P1_U2832) );
  INV_X1 U17078 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n21000) );
  OAI222_X1 U17079 ( .A1(n13793), .A2(n15712), .B1(n20078), .B2(n21000), .C1(
        n14439), .C2(n13784), .ZN(P1_U2863) );
  OAI21_X1 U17080 ( .B1(n13718), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n13717), .ZN(n16163) );
  XNOR2_X1 U17081 ( .A(n13720), .B(n13719), .ZN(n19163) );
  OAI21_X1 U17082 ( .B1(n15202), .B2(n13722), .A(n13721), .ZN(n15286) );
  INV_X1 U17083 ( .A(n15286), .ZN(n16251) );
  OAI21_X1 U17084 ( .B1(n15285), .B2(n13724), .A(n16251), .ZN(n15271) );
  AOI22_X1 U17085 ( .A1(n19016), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15271), .ZN(n13723) );
  OAI21_X1 U17086 ( .B1(n16215), .B2(n19163), .A(n13723), .ZN(n13726) );
  AND4_X1 U17087 ( .A1(n16241), .A2(n13724), .A3(n15272), .A4(n16257), .ZN(
        n13725) );
  AOI211_X1 U17088 ( .C1(n19009), .C2(n19255), .A(n13726), .B(n13725), .ZN(
        n13730) );
  XNOR2_X1 U17089 ( .A(n13728), .B(n13727), .ZN(n16166) );
  OR2_X1 U17090 ( .A1(n16166), .A2(n16246), .ZN(n13729) );
  OAI211_X1 U17091 ( .C1(n16163), .C2(n16264), .A(n13730), .B(n13729), .ZN(
        P2_U3040) );
  NOR2_X1 U17092 ( .A1(n15906), .A2(n13736), .ZN(n15921) );
  INV_X1 U17093 ( .A(n15921), .ZN(n13742) );
  NAND2_X1 U17094 ( .A1(n13731), .A2(n13732), .ZN(n13733) );
  NAND2_X1 U17095 ( .A1(n13734), .A2(n13733), .ZN(n15773) );
  NAND2_X1 U17096 ( .A1(n15773), .A2(n15933), .ZN(n13741) );
  NOR3_X1 U17097 ( .A1(n13737), .A2(n13736), .A3(n13735), .ZN(n15939) );
  NOR2_X1 U17098 ( .A1(n13790), .A2(n15939), .ZN(n15919) );
  INV_X1 U17099 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n21008) );
  OAI22_X1 U17100 ( .A1(n20137), .A2(n13738), .B1(n21008), .B2(n20135), .ZN(
        n13739) );
  AOI21_X1 U17101 ( .B1(n15919), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13739), .ZN(n13740) );
  OAI211_X1 U17102 ( .C1(n13742), .C2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13741), .B(n13740), .ZN(P1_U3024) );
  OAI21_X1 U17103 ( .B1(n13635), .B2(n13744), .A(n13819), .ZN(n14644) );
  NOR2_X1 U17104 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n21029), .ZN(n13752) );
  NAND2_X1 U17105 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .ZN(n13804) );
  INV_X1 U17106 ( .A(n13804), .ZN(n14400) );
  INV_X1 U17107 ( .A(n20062), .ZN(n20016) );
  AOI21_X1 U17108 ( .B1(n14400), .B2(n13745), .A(n20016), .ZN(n15702) );
  OAI21_X1 U17109 ( .B1(n13747), .B2(n13746), .A(n15696), .ZN(n13756) );
  INV_X1 U17110 ( .A(n13756), .ZN(n15910) );
  AOI22_X1 U17111 ( .A1(n15910), .A2(n20067), .B1(n20046), .B2(
        P1_EBX_REG_10__SCAN_IN), .ZN(n13748) );
  OAI211_X1 U17112 ( .C1(n20064), .C2(n14640), .A(n13748), .B(n20135), .ZN(
        n13749) );
  AOI21_X1 U17113 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15702), .A(n13749), 
        .ZN(n13750) );
  OAI21_X1 U17114 ( .B1(n14635), .B2(n20063), .A(n13750), .ZN(n13751) );
  AOI21_X1 U17115 ( .B1(n14399), .B2(n13752), .A(n13751), .ZN(n13753) );
  OAI21_X1 U17116 ( .B1(n15623), .B2(n14644), .A(n13753), .ZN(P1_U2830) );
  INV_X1 U17117 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13754) );
  OAI222_X1 U17118 ( .A1(n14644), .A2(n14499), .B1(n14456), .B2(n14504), .C1(
        n13754), .C2(n14502), .ZN(P1_U2894) );
  INV_X1 U17119 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13755) );
  OAI222_X1 U17120 ( .A1(n13756), .A2(n15712), .B1(n13755), .B2(n20078), .C1(
        n14439), .C2(n14644), .ZN(P1_U2862) );
  XOR2_X1 U17121 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13758), .Z(
        n13759) );
  XNOR2_X1 U17122 ( .A(n13757), .B(n13759), .ZN(n15920) );
  NAND2_X1 U17123 ( .A1(n15920), .A2(n20127), .ZN(n13763) );
  AND2_X1 U17124 ( .A1(n15899), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15917) );
  NOR2_X1 U17125 ( .A1(n15782), .A2(n13760), .ZN(n13761) );
  AOI211_X1 U17126 ( .C1(n20125), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15917), .B(n13761), .ZN(n13762) );
  OAI211_X1 U17127 ( .C1(n20131), .C2(n13764), .A(n13763), .B(n13762), .ZN(
        P1_U2991) );
  OR2_X1 U17128 ( .A1(n13819), .A2(n13765), .ZN(n13799) );
  OR2_X1 U17129 ( .A1(n13819), .A2(n13766), .ZN(n14392) );
  NAND2_X1 U17130 ( .A1(n14392), .A2(n13767), .ZN(n13768) );
  NAND2_X1 U17131 ( .A1(n13799), .A2(n13768), .ZN(n15713) );
  AOI22_X1 U17132 ( .A1(n13772), .A2(n14440), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14487), .ZN(n13769) );
  OAI21_X1 U17133 ( .B1(n15713), .B2(n14499), .A(n13769), .ZN(P1_U2890) );
  XNOR2_X1 U17134 ( .A(n13819), .B(n13817), .ZN(n13771) );
  NAND2_X1 U17135 ( .A1(n13771), .A2(n13770), .ZN(n13818) );
  OAI21_X1 U17136 ( .B1(n13771), .B2(n13770), .A(n13818), .ZN(n15703) );
  AOI22_X1 U17137 ( .A1(n13772), .A2(n14451), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n14487), .ZN(n13773) );
  OAI21_X1 U17138 ( .B1(n15703), .B2(n14499), .A(n13773), .ZN(P1_U2893) );
  NOR2_X1 U17139 ( .A1(n13775), .A2(n13776), .ZN(n13777) );
  OR2_X1 U17140 ( .A1(n13774), .A2(n13777), .ZN(n15664) );
  INV_X1 U17141 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20152) );
  OAI22_X1 U17142 ( .A1(n14493), .A2(n20152), .B1(n13778), .B2(n14502), .ZN(
        n13779) );
  INV_X1 U17143 ( .A(n13779), .ZN(n13781) );
  AOI22_X1 U17144 ( .A1(n14496), .A2(DATAI_16_), .B1(n14495), .B2(n20151), 
        .ZN(n13780) );
  OAI211_X1 U17145 ( .C1(n15664), .C2(n14499), .A(n13781), .B(n13780), .ZN(
        P1_U2888) );
  XNOR2_X1 U17146 ( .A(n9820), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13783) );
  XNOR2_X1 U17147 ( .A(n13782), .B(n13783), .ZN(n13798) );
  NAND2_X1 U17148 ( .A1(n15935), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n13792) );
  OAI21_X1 U17149 ( .B1(n15790), .B2(n10690), .A(n13792), .ZN(n13786) );
  NOR2_X1 U17150 ( .A1(n13784), .A2(n20131), .ZN(n13785) );
  AOI211_X1 U17151 ( .C1(n15783), .C2(n13787), .A(n13786), .B(n13785), .ZN(
        n13788) );
  OAI21_X1 U17152 ( .B1(n13798), .B2(n19996), .A(n13788), .ZN(P1_U2990) );
  INV_X1 U17153 ( .A(n15885), .ZN(n13789) );
  AOI21_X1 U17154 ( .B1(n15881), .B2(n15882), .A(n13789), .ZN(n13791) );
  AOI21_X1 U17155 ( .B1(n13794), .B2(n13791), .A(n13790), .ZN(n15912) );
  OAI21_X1 U17156 ( .B1(n20137), .B2(n13793), .A(n13792), .ZN(n13796) );
  NAND2_X1 U17157 ( .A1(n13794), .A2(n15927), .ZN(n15916) );
  NOR2_X1 U17158 ( .A1(n15916), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13795) );
  AOI211_X1 U17159 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n15912), .A(
        n13796), .B(n13795), .ZN(n13797) );
  OAI21_X1 U17160 ( .B1(n13798), .B2(n20138), .A(n13797), .ZN(P1_U3022) );
  AOI21_X1 U17161 ( .B1(n13800), .B2(n13799), .A(n13775), .ZN(n13814) );
  INV_X1 U17162 ( .A(n13801), .ZN(n15667) );
  XNOR2_X1 U17163 ( .A(n15676), .B(n15667), .ZN(n15853) );
  OAI22_X1 U17164 ( .A1(n15853), .A2(n15712), .B1(n21009), .B2(n20078), .ZN(
        n13802) );
  AOI21_X1 U17165 ( .B1(n13814), .B2(n20074), .A(n13802), .ZN(n13803) );
  INV_X1 U17166 ( .A(n13803), .ZN(P1_U2857) );
  INV_X1 U17167 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21138) );
  NAND2_X1 U17168 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .ZN(n14401) );
  NOR4_X1 U17169 ( .A1(n21138), .A2(n13805), .A3(n13804), .A4(n14401), .ZN(
        n15679) );
  NAND2_X1 U17170 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n15679), .ZN(n13830) );
  NOR2_X1 U17171 ( .A1(n13830), .A2(n15677), .ZN(n15657) );
  INV_X1 U17172 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21124) );
  NAND2_X1 U17173 ( .A1(n15657), .A2(n21124), .ZN(n13811) );
  INV_X1 U17174 ( .A(n13830), .ZN(n13806) );
  AOI21_X1 U17175 ( .B1(n15644), .B2(n13831), .A(n14332), .ZN(n20060) );
  OAI21_X1 U17176 ( .B1(n13806), .B2(n20016), .A(n20060), .ZN(n15678) );
  INV_X1 U17177 ( .A(n14619), .ZN(n13807) );
  AOI22_X1 U17178 ( .A1(n20053), .A2(n13807), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n20061), .ZN(n13808) );
  OAI211_X1 U17179 ( .C1(n20064), .C2(n10708), .A(n13808), .B(n20135), .ZN(
        n13809) );
  AOI21_X1 U17180 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15678), .A(n13809), 
        .ZN(n13810) );
  OAI211_X1 U17181 ( .C1(n15853), .C2(n20049), .A(n13811), .B(n13810), .ZN(
        n13812) );
  AOI21_X1 U17182 ( .B1(n13814), .B2(n20025), .A(n13812), .ZN(n13813) );
  INV_X1 U17183 ( .A(n13813), .ZN(P1_U2825) );
  INV_X1 U17184 ( .A(n13814), .ZN(n14623) );
  OAI222_X1 U17185 ( .A1(n14623), .A2(n14499), .B1(n14504), .B2(n13816), .C1(
        n14502), .C2(n13815), .ZN(P1_U2889) );
  INV_X1 U17186 ( .A(n13817), .ZN(n13820) );
  OAI21_X1 U17187 ( .B1(n13820), .B2(n13819), .A(n13818), .ZN(n13822) );
  NAND2_X1 U17188 ( .A1(n13822), .A2(n13821), .ZN(n14395) );
  OAI21_X1 U17189 ( .B1(n13822), .B2(n13821), .A(n14395), .ZN(n15691) );
  OAI222_X1 U17190 ( .A1(n15691), .A2(n14499), .B1(n14446), .B2(n14504), .C1(
        n13823), .C2(n14502), .ZN(P1_U2892) );
  OAI21_X1 U17191 ( .B1(n13774), .B2(n13824), .A(n9833), .ZN(n14612) );
  XNOR2_X1 U17192 ( .A(n15668), .B(n15649), .ZN(n15837) );
  AOI22_X1 U17193 ( .A1(n15837), .A2(n20073), .B1(n14437), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n13825) );
  OAI21_X1 U17194 ( .B1(n14612), .B2(n14439), .A(n13825), .ZN(P1_U2855) );
  AOI21_X1 U17195 ( .B1(n20046), .B2(P1_EBX_REG_17__SCAN_IN), .A(n15935), .ZN(
        n13827) );
  NAND2_X1 U17196 ( .A1(n15837), .A2(n20067), .ZN(n13826) );
  OAI211_X1 U17197 ( .C1(n20064), .C2(n14607), .A(n13827), .B(n13826), .ZN(
        n13828) );
  AOI21_X1 U17198 ( .B1(n20053), .B2(n14609), .A(n13828), .ZN(n13834) );
  INV_X1 U17199 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20752) );
  NAND2_X1 U17200 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15657), .ZN(n15659) );
  INV_X1 U17201 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20754) );
  OAI21_X1 U17202 ( .B1(n20752), .B2(n15659), .A(n20754), .ZN(n13832) );
  NAND3_X1 U17203 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_17__SCAN_IN), 
        .A3(P1_REIP_REG_16__SCAN_IN), .ZN(n13829) );
  NOR3_X1 U17204 ( .A1(n13831), .A2(n13830), .A3(n13829), .ZN(n15643) );
  OAI21_X1 U17205 ( .B1(n15643), .B2(n15630), .A(n15629), .ZN(n15642) );
  NAND2_X1 U17206 ( .A1(n13832), .A2(n15642), .ZN(n13833) );
  OAI211_X1 U17207 ( .C1(n14612), .C2(n15623), .A(n13834), .B(n13833), .ZN(
        P1_U2823) );
  AOI22_X1 U17208 ( .A1(n14488), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14487), .ZN(n13836) );
  AOI22_X1 U17209 ( .A1(n14496), .A2(DATAI_17_), .B1(n14495), .B2(n20158), 
        .ZN(n13835) );
  OAI211_X1 U17210 ( .C1(n14612), .C2(n14499), .A(n13836), .B(n13835), .ZN(
        P1_U2887) );
  INV_X1 U17211 ( .A(n13837), .ZN(n13838) );
  NOR2_X2 U17212 ( .A1(n13838), .A2(n18606), .ZN(n18604) );
  OAI21_X1 U17213 ( .B1(n15463), .B2(n18782), .A(n18639), .ZN(n13839) );
  NAND2_X1 U17214 ( .A1(n18604), .A2(n13839), .ZN(n18591) );
  NOR2_X1 U17215 ( .A1(n18771), .A2(n18591), .ZN(n13846) );
  INV_X1 U17216 ( .A(n18642), .ZN(n18649) );
  NAND2_X1 U17217 ( .A1(n16489), .A2(n13840), .ZN(n17350) );
  NAND2_X1 U17218 ( .A1(n18586), .A2(n18809), .ZN(n13845) );
  NOR2_X1 U17219 ( .A1(n17413), .A2(n18604), .ZN(n13841) );
  NOR3_X2 U17220 ( .A1(n18669), .A2(n13841), .A3(n16471), .ZN(n15583) );
  NOR2_X1 U17221 ( .A1(n15583), .A2(n15441), .ZN(n13843) );
  OAI211_X1 U17222 ( .C1(n17350), .C2(n13845), .A(n13844), .B(n13843), .ZN(
        n18614) );
  INV_X1 U17223 ( .A(n18614), .ZN(n18626) );
  NAND2_X1 U17224 ( .A1(n18652), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18155) );
  INV_X1 U17225 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16475) );
  NAND3_X1 U17226 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18756)
         );
  OR2_X1 U17227 ( .A1(n16475), .A2(n18756), .ZN(n15465) );
  OAI211_X1 U17228 ( .C1(n18649), .C2(n18626), .A(n18155), .B(n15465), .ZN(
        n18787) );
  MUX2_X1 U17229 ( .A(n13846), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18790), .Z(P3_U3284) );
  NAND2_X1 U17230 ( .A1(n13847), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13854) );
  NAND2_X1 U17231 ( .A1(n13848), .A2(n15081), .ZN(n13852) );
  NAND2_X1 U17232 ( .A1(n13854), .A2(n13853), .ZN(n14902) );
  NAND2_X1 U17233 ( .A1(n12264), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13858) );
  AOI21_X1 U17234 ( .B1(n15986), .B2(n13959), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14900) );
  INV_X1 U17235 ( .A(n14900), .ZN(n13856) );
  AND2_X2 U17236 ( .A1(n14902), .A2(n13856), .ZN(n13951) );
  INV_X1 U17237 ( .A(n15986), .ZN(n13857) );
  INV_X1 U17238 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14910) );
  NAND2_X1 U17239 ( .A1(n13859), .A2(n13858), .ZN(n13956) );
  AND2_X1 U17240 ( .A1(n12264), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13860) );
  XNOR2_X1 U17241 ( .A(n13956), .B(n13860), .ZN(n15977) );
  INV_X1 U17242 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13984) );
  OR2_X1 U17243 ( .A1(n13861), .A2(n13984), .ZN(n13862) );
  NOR2_X1 U17244 ( .A1(n15977), .A2(n13862), .ZN(n13952) );
  INV_X1 U17245 ( .A(n13952), .ZN(n13863) );
  OAI21_X1 U17246 ( .B1(n15977), .B2(n13861), .A(n13984), .ZN(n13950) );
  NAND2_X1 U17247 ( .A1(n13863), .A2(n13950), .ZN(n13864) );
  XNOR2_X1 U17248 ( .A(n13865), .B(n13864), .ZN(n14899) );
  NAND2_X1 U17249 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15064), .ZN(
        n13985) );
  NAND2_X1 U17250 ( .A1(n16257), .A2(n13985), .ZN(n13866) );
  NAND2_X1 U17251 ( .A1(n15079), .A2(n13866), .ZN(n13987) );
  INV_X1 U17252 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n13869) );
  OR2_X1 U17253 ( .A1(n13970), .A2(n14910), .ZN(n13868) );
  AOI22_X1 U17254 ( .A1(n13965), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n13867) );
  OAI211_X1 U17255 ( .C1(n13870), .C2(n13869), .A(n13868), .B(n13867), .ZN(
        n14743) );
  NAND2_X1 U17256 ( .A1(n14744), .A2(n14743), .ZN(n14742) );
  INV_X1 U17257 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U17258 ( .A1(n13966), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13872) );
  NAND2_X1 U17259 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13871) );
  OAI211_X1 U17260 ( .C1(n13873), .C2(n13879), .A(n13872), .B(n13871), .ZN(
        n13874) );
  AOI21_X1 U17261 ( .B1(n13875), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n13874), .ZN(n13876) );
  NAND2_X1 U17262 ( .A1(n14742), .A2(n13876), .ZN(n13877) );
  NAND2_X1 U17263 ( .A1(n13973), .A2(n13877), .ZN(n15983) );
  NAND2_X1 U17264 ( .A1(n12763), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U17265 ( .A1(n13988), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n13878) );
  OAI21_X1 U17266 ( .B1(n12759), .B2(n13879), .A(n13878), .ZN(n13880) );
  INV_X1 U17267 ( .A(n13880), .ZN(n13882) );
  INV_X1 U17268 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19896) );
  AOI22_X1 U17269 ( .A1(n13988), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12594), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13881) );
  OAI21_X1 U17270 ( .B1(n12759), .B2(n19896), .A(n13881), .ZN(n14811) );
  NAND2_X1 U17271 ( .A1(n14812), .A2(n14811), .ZN(n14814) );
  AOI21_X1 U17272 ( .B1(n13882), .B2(n14814), .A(n13991), .ZN(n15979) );
  NAND2_X1 U17273 ( .A1(n15979), .A2(n19257), .ZN(n13883) );
  OAI211_X1 U17274 ( .C1(n15983), .C2(n16253), .A(n14894), .B(n13883), .ZN(
        n13885) );
  NOR3_X1 U17275 ( .A1(n15074), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n13985), .ZN(n13884) );
  AOI211_X1 U17276 ( .C1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n13987), .A(
        n13885), .B(n13884), .ZN(n13887) );
  XNOR2_X1 U17277 ( .A(n13962), .B(n13984), .ZN(n14897) );
  NAND2_X1 U17278 ( .A1(n14897), .A2(n19262), .ZN(n13886) );
  OAI211_X1 U17279 ( .C1(n14899), .C2(n16246), .A(n13887), .B(n13886), .ZN(
        P2_U3016) );
  AOI211_X1 U17280 ( .C1(n13894), .C2(n12056), .A(n13888), .B(n15285), .ZN(
        n13899) );
  OAI21_X1 U17281 ( .B1(n13890), .B2(n19050), .A(n13889), .ZN(n13891) );
  XNOR2_X1 U17282 ( .A(n13891), .B(n13894), .ZN(n13905) );
  INV_X1 U17283 ( .A(n13905), .ZN(n13892) );
  NAND2_X1 U17284 ( .A1(n13892), .A2(n19263), .ZN(n13893) );
  NAND2_X1 U17285 ( .A1(n12763), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n13903) );
  OAI211_X1 U17286 ( .C1(n16254), .C2(n13894), .A(n13893), .B(n13903), .ZN(
        n13898) );
  OAI21_X1 U17287 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13896), .A(
        n13895), .ZN(n13901) );
  OAI22_X1 U17288 ( .A1(n16215), .A2(n19056), .B1(n13901), .B2(n16264), .ZN(
        n13897) );
  NOR3_X1 U17289 ( .A1(n13899), .A2(n13898), .A3(n13897), .ZN(n13900) );
  OAI21_X1 U17290 ( .B1(n13910), .B2(n16253), .A(n13900), .ZN(P2_U3045) );
  INV_X1 U17291 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13908) );
  INV_X1 U17292 ( .A(n13901), .ZN(n13902) );
  NAND2_X1 U17293 ( .A1(n13902), .A2(n19242), .ZN(n13904) );
  OAI211_X1 U17294 ( .C1(n13908), .C2(n16179), .A(n13904), .B(n13903), .ZN(
        n13907) );
  NOR2_X1 U17295 ( .A1(n13905), .A2(n16173), .ZN(n13906) );
  AOI211_X1 U17296 ( .C1(n16170), .C2(n13908), .A(n13907), .B(n13906), .ZN(
        n13909) );
  OAI21_X1 U17297 ( .B1(n13910), .B2(n15339), .A(n13909), .ZN(P2_U3013) );
  NAND2_X1 U17298 ( .A1(n13912), .A2(n13911), .ZN(n13913) );
  XOR2_X1 U17299 ( .A(n13913), .B(n9879), .Z(n16125) );
  AND2_X1 U17300 ( .A1(n15250), .A2(n12512), .ZN(n16123) );
  NOR2_X1 U17301 ( .A1(n15250), .A2(n12512), .ZN(n16124) );
  OR3_X1 U17302 ( .A1(n16123), .A2(n16124), .A3(n16264), .ZN(n13927) );
  OAI21_X1 U17303 ( .B1(n15182), .B2(n10087), .A(n15185), .ZN(n16209) );
  INV_X1 U17304 ( .A(n16209), .ZN(n15247) );
  NOR2_X1 U17305 ( .A1(n13916), .A2(n13915), .ZN(n13917) );
  NOR2_X1 U17306 ( .A1(n13918), .A2(n13917), .ZN(n18943) );
  INV_X1 U17307 ( .A(n18943), .ZN(n19101) );
  NAND2_X1 U17308 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19016), .ZN(n13922) );
  AOI21_X1 U17309 ( .B1(n13920), .B2(n13919), .A(n15237), .ZN(n19144) );
  NAND2_X1 U17310 ( .A1(n19257), .A2(n19144), .ZN(n13921) );
  OAI211_X1 U17311 ( .C1(n19101), .C2(n16253), .A(n13922), .B(n13921), .ZN(
        n13925) );
  INV_X1 U17312 ( .A(n13935), .ZN(n15256) );
  NAND2_X1 U17313 ( .A1(n15256), .A2(n13923), .ZN(n16201) );
  NOR2_X1 U17314 ( .A1(n16201), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13924) );
  AOI211_X1 U17315 ( .C1(n15247), .C2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n13925), .B(n13924), .ZN(n13926) );
  OAI211_X1 U17316 ( .C1(n16125), .C2(n16246), .A(n13927), .B(n13926), .ZN(
        P2_U3034) );
  INV_X1 U17317 ( .A(n13928), .ZN(n16135) );
  NOR2_X1 U17318 ( .A1(n16135), .A2(n13929), .ZN(n13931) );
  XOR2_X1 U17319 ( .A(n13931), .B(n13930), .Z(n13949) );
  INV_X1 U17320 ( .A(n13914), .ZN(n13932) );
  NAND2_X1 U17321 ( .A1(n13932), .A2(n13936), .ZN(n13942) );
  NAND3_X1 U17322 ( .A1(n13942), .A2(n19262), .A3(n16144), .ZN(n13941) );
  XOR2_X1 U17323 ( .A(n13933), .B(n13934), .Z(n18978) );
  INV_X1 U17324 ( .A(n18978), .ZN(n19154) );
  NAND2_X1 U17325 ( .A1(n12763), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n13944) );
  OAI21_X1 U17326 ( .B1(n16215), .B2(n19154), .A(n13944), .ZN(n13938) );
  NOR2_X1 U17327 ( .A1(n13936), .A2(n15182), .ZN(n15254) );
  AOI21_X1 U17328 ( .B1(n13936), .B2(n13935), .A(n15254), .ZN(n13937) );
  AOI211_X1 U17329 ( .C1(n13939), .C2(n19255), .A(n13938), .B(n13937), .ZN(
        n13940) );
  OAI211_X1 U17330 ( .C1(n13949), .C2(n16246), .A(n13941), .B(n13940), .ZN(
        P2_U3037) );
  NAND3_X1 U17331 ( .A1(n13942), .A2(n19242), .A3(n16144), .ZN(n13948) );
  AOI21_X1 U17332 ( .B1(n18972), .B2(n15490), .A(n13943), .ZN(n18976) );
  AOI22_X1 U17333 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n16170), .B2(n18976), .ZN(n13945) );
  OAI211_X1 U17334 ( .C1(n15339), .C2(n18981), .A(n13945), .B(n13944), .ZN(
        n13946) );
  INV_X1 U17335 ( .A(n13946), .ZN(n13947) );
  OAI211_X1 U17336 ( .C1(n16173), .C2(n13949), .A(n13948), .B(n13947), .ZN(
        P2_U3005) );
  NAND2_X1 U17337 ( .A1(n13951), .A2(n13950), .ZN(n13954) );
  INV_X1 U17338 ( .A(n13955), .ZN(n13958) );
  NOR2_X1 U17339 ( .A1(n13956), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13957) );
  MUX2_X1 U17340 ( .A(n13958), .B(n13957), .S(n12264), .Z(n15956) );
  NAND2_X1 U17341 ( .A1(n15956), .A2(n13959), .ZN(n13960) );
  NOR2_X1 U17342 ( .A1(n13964), .A2(n19247), .ZN(n13976) );
  AOI22_X1 U17343 ( .A1(n13965), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n13968) );
  NAND2_X1 U17344 ( .A1(n13966), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13967) );
  OAI211_X1 U17345 ( .C1(n13970), .C2(n13969), .A(n13968), .B(n13967), .ZN(
        n13971) );
  INV_X1 U17346 ( .A(n13971), .ZN(n13972) );
  AND2_X1 U17347 ( .A1(n19016), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n13992) );
  AOI21_X1 U17348 ( .B1(n19239), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13992), .ZN(n13974) );
  OAI21_X1 U17349 ( .B1(n16060), .B2(n15339), .A(n13974), .ZN(n13975) );
  OAI21_X1 U17350 ( .B1(n13999), .B2(n16173), .A(n13977), .ZN(P2_U2983) );
  AOI21_X1 U17351 ( .B1(n20125), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n13978), .ZN(n13979) );
  OAI21_X1 U17352 ( .B1(n15782), .B2(n13980), .A(n13979), .ZN(n13981) );
  AOI21_X1 U17353 ( .B1(n14282), .B2(n15786), .A(n13981), .ZN(n13982) );
  OAI21_X1 U17354 ( .B1(n13983), .B2(n19996), .A(n13982), .ZN(P1_U2968) );
  NOR4_X1 U17355 ( .A1(n15074), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n13985), .A4(n13984), .ZN(n13996) );
  NOR2_X1 U17356 ( .A1(n15285), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13986) );
  OAI21_X1 U17357 ( .B1(n13987), .B2(n13986), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13994) );
  AOI222_X1 U17358 ( .A1(n13989), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n13988), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12594), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13990) );
  XNOR2_X1 U17359 ( .A(n13991), .B(n13990), .ZN(n15969) );
  OAI211_X1 U17360 ( .C1(n16060), .C2(n16253), .A(n13994), .B(n13993), .ZN(
        n13995) );
  OAI21_X1 U17361 ( .B1(n13999), .B2(n16246), .A(n13998), .ZN(P2_U3015) );
  AOI22_X1 U17362 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14005) );
  AOI22_X1 U17363 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n9816), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14004) );
  AOI22_X1 U17364 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14003) );
  AOI22_X1 U17365 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14002) );
  NAND4_X1 U17366 ( .A1(n14005), .A2(n14004), .A3(n14003), .A4(n14002), .ZN(
        n14011) );
  AOI22_X1 U17367 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14009) );
  AOI22_X1 U17368 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14008) );
  AOI22_X1 U17369 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14007) );
  AOI22_X1 U17370 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14006) );
  NAND4_X1 U17371 ( .A1(n14009), .A2(n14008), .A3(n14007), .A4(n14006), .ZN(
        n14010) );
  NOR2_X1 U17372 ( .A1(n14011), .A2(n14010), .ZN(n16071) );
  INV_X1 U17373 ( .A(n16071), .ZN(n14012) );
  AOI22_X1 U17374 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n14016) );
  AOI22_X1 U17375 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n9816), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14015) );
  AOI22_X1 U17376 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14014) );
  AOI22_X1 U17377 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14013) );
  NAND4_X1 U17378 ( .A1(n14016), .A2(n14015), .A3(n14014), .A4(n14013), .ZN(
        n14022) );
  AOI22_X1 U17379 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14020) );
  AOI22_X1 U17380 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14019) );
  AOI22_X1 U17381 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14018) );
  AOI22_X1 U17382 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14017) );
  NAND4_X1 U17383 ( .A1(n14020), .A2(n14019), .A3(n14018), .A4(n14017), .ZN(
        n14021) );
  OR2_X1 U17384 ( .A1(n14022), .A2(n14021), .ZN(n14798) );
  AOI22_X1 U17385 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14026) );
  AOI22_X1 U17386 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n9815), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14025) );
  AOI22_X1 U17387 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14024) );
  AOI22_X1 U17388 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14023) );
  NAND4_X1 U17389 ( .A1(n14026), .A2(n14025), .A3(n14024), .A4(n14023), .ZN(
        n14033) );
  AOI22_X1 U17390 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U17391 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17392 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14029) );
  AOI22_X1 U17393 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14028) );
  NAND4_X1 U17394 ( .A1(n14031), .A2(n14030), .A3(n14029), .A4(n14028), .ZN(
        n14032) );
  NOR2_X1 U17395 ( .A1(n14033), .A2(n14032), .ZN(n16069) );
  AOI22_X1 U17396 ( .A1(n11896), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12149), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U17397 ( .A1(n9815), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17398 ( .A1(n12148), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12726), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14039) );
  INV_X1 U17399 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14036) );
  OAI22_X1 U17400 ( .A1(n14036), .A2(n9858), .B1(n14035), .B2(n14034), .ZN(
        n14037) );
  INV_X1 U17401 ( .A(n14037), .ZN(n14038) );
  NAND4_X1 U17402 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14047) );
  AOI22_X1 U17403 ( .A1(n14027), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12155), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U17404 ( .A1(n11881), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U17405 ( .A1(n11912), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U17406 ( .A1(n12154), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14042) );
  NAND4_X1 U17407 ( .A1(n14045), .A2(n14044), .A3(n14043), .A4(n14042), .ZN(
        n14046) );
  OR2_X1 U17408 ( .A1(n14047), .A2(n14046), .ZN(n14790) );
  AOI22_X1 U17409 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17410 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n9815), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U17411 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U17412 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14048) );
  NAND4_X1 U17413 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14057) );
  AOI22_X1 U17414 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17415 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17416 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14053) );
  AOI22_X1 U17417 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14052) );
  NAND4_X1 U17418 ( .A1(n14055), .A2(n14054), .A3(n14053), .A4(n14052), .ZN(
        n14056) );
  NOR2_X1 U17419 ( .A1(n14057), .A2(n14056), .ZN(n16065) );
  INV_X1 U17420 ( .A(n14263), .ZN(n14235) );
  INV_X1 U17421 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15362) );
  INV_X1 U17422 ( .A(n14262), .ZN(n14233) );
  INV_X1 U17423 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14058) );
  OAI22_X1 U17424 ( .A1(n14235), .A2(n15362), .B1(n14233), .B2(n14058), .ZN(
        n14062) );
  INV_X1 U17425 ( .A(n14265), .ZN(n14239) );
  INV_X1 U17426 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14060) );
  INV_X1 U17427 ( .A(n14264), .ZN(n14237) );
  INV_X1 U17428 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14059) );
  OAI22_X1 U17429 ( .A1(n14239), .A2(n14060), .B1(n14237), .B2(n14059), .ZN(
        n14061) );
  NOR2_X1 U17430 ( .A1(n14062), .A2(n14061), .ZN(n14066) );
  AOI22_X1 U17431 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14065) );
  INV_X1 U17432 ( .A(n14063), .ZN(n16277) );
  INV_X1 U17433 ( .A(n16277), .ZN(n14259) );
  AOI22_X1 U17434 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14064) );
  XNOR2_X1 U17435 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14253) );
  NAND4_X1 U17436 ( .A1(n14066), .A2(n14065), .A3(n14064), .A4(n14253), .ZN(
        n14077) );
  INV_X1 U17437 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14068) );
  INV_X1 U17438 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14067) );
  OAI22_X1 U17439 ( .A1(n14235), .A2(n14068), .B1(n14233), .B2(n14067), .ZN(
        n14072) );
  INV_X1 U17440 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14070) );
  INV_X1 U17441 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n14069) );
  OAI22_X1 U17442 ( .A1(n14239), .A2(n14070), .B1(n14237), .B2(n14069), .ZN(
        n14071) );
  NOR2_X1 U17443 ( .A1(n14072), .A2(n14071), .ZN(n14075) );
  AOI22_X1 U17444 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14074) );
  INV_X1 U17445 ( .A(n14253), .ZN(n14267) );
  AOI22_X1 U17446 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14073) );
  NAND4_X1 U17447 ( .A1(n14075), .A2(n14074), .A3(n14267), .A4(n14073), .ZN(
        n14076) );
  AND2_X1 U17448 ( .A1(n14077), .A2(n14076), .ZN(n14112) );
  NAND2_X1 U17449 ( .A1(n19976), .A2(n14112), .ZN(n14090) );
  AOI22_X1 U17450 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12149), .B1(
        n11896), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17451 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n9816), .B1(n9814), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17452 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12726), .B1(
        n12148), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17453 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n14079), .B1(
        n14078), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14080) );
  NAND4_X1 U17454 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14089) );
  AOI22_X1 U17455 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n12155), .B1(
        n14027), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U17456 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n11881), .B1(
        n11863), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14086) );
  AOI22_X1 U17457 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n11912), .B1(
        n12147), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14085) );
  AOI22_X1 U17458 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12154), .B1(
        n11862), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14084) );
  NAND4_X1 U17459 ( .A1(n14087), .A2(n14086), .A3(n14085), .A4(n14084), .ZN(
        n14088) );
  OR2_X1 U17460 ( .A1(n14089), .A2(n14088), .ZN(n14113) );
  XNOR2_X1 U17461 ( .A(n14090), .B(n14113), .ZN(n14118) );
  INV_X1 U17462 ( .A(n14112), .ZN(n14116) );
  NOR2_X1 U17463 ( .A1(n19976), .A2(n14116), .ZN(n14857) );
  INV_X1 U17464 ( .A(n14091), .ZN(n16064) );
  INV_X1 U17465 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14094) );
  OAI22_X1 U17466 ( .A1(n14235), .A2(n14094), .B1(n14233), .B2(n14093), .ZN(
        n14097) );
  INV_X1 U17467 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14095) );
  OAI22_X1 U17468 ( .A1(n14239), .A2(n14095), .B1(n14237), .B2(n19272), .ZN(
        n14096) );
  NOR2_X1 U17469 ( .A1(n14097), .A2(n14096), .ZN(n14100) );
  AOI22_X1 U17470 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14099) );
  AOI22_X1 U17471 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n14098) );
  NAND4_X1 U17472 ( .A1(n14100), .A2(n14099), .A3(n14098), .A4(n14253), .ZN(
        n14111) );
  OAI22_X1 U17473 ( .A1(n14235), .A2(n14102), .B1(n14233), .B2(n14101), .ZN(
        n14106) );
  INV_X1 U17474 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14104) );
  INV_X1 U17475 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n14103) );
  OAI22_X1 U17476 ( .A1(n14239), .A2(n14104), .B1(n14237), .B2(n14103), .ZN(
        n14105) );
  NOR2_X1 U17477 ( .A1(n14106), .A2(n14105), .ZN(n14109) );
  AOI22_X1 U17478 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17479 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14107) );
  NAND4_X1 U17480 ( .A1(n14109), .A2(n14108), .A3(n14267), .A4(n14107), .ZN(
        n14110) );
  AND2_X1 U17481 ( .A1(n14111), .A2(n14110), .ZN(n14115) );
  AND2_X1 U17482 ( .A1(n14113), .A2(n14112), .ZN(n14114) );
  NAND2_X1 U17483 ( .A1(n14114), .A2(n14115), .ZN(n14119) );
  OAI211_X1 U17484 ( .C1(n14115), .C2(n14114), .A(n14198), .B(n14119), .ZN(
        n14780) );
  NAND2_X1 U17485 ( .A1(n12584), .A2(n14115), .ZN(n14783) );
  NOR2_X1 U17486 ( .A1(n14783), .A2(n14116), .ZN(n14117) );
  INV_X1 U17487 ( .A(n14119), .ZN(n14139) );
  INV_X1 U17488 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14121) );
  INV_X1 U17489 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14120) );
  OAI22_X1 U17490 ( .A1(n14235), .A2(n14121), .B1(n14233), .B2(n14120), .ZN(
        n14124) );
  INV_X1 U17491 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14122) );
  INV_X1 U17492 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19277) );
  OAI22_X1 U17493 ( .A1(n14239), .A2(n14122), .B1(n14237), .B2(n19277), .ZN(
        n14123) );
  NOR2_X1 U17494 ( .A1(n14124), .A2(n14123), .ZN(n14127) );
  AOI22_X1 U17495 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14126) );
  AOI22_X1 U17496 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14125) );
  NAND4_X1 U17497 ( .A1(n14127), .A2(n14126), .A3(n14125), .A4(n14253), .ZN(
        n14138) );
  INV_X1 U17498 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14129) );
  INV_X1 U17499 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14128) );
  OAI22_X1 U17500 ( .A1(n14235), .A2(n14129), .B1(n14233), .B2(n14128), .ZN(
        n14133) );
  INV_X1 U17501 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14131) );
  INV_X1 U17502 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n14130) );
  OAI22_X1 U17503 ( .A1(n14239), .A2(n14131), .B1(n14237), .B2(n14130), .ZN(
        n14132) );
  NOR2_X1 U17504 ( .A1(n14133), .A2(n14132), .ZN(n14136) );
  AOI22_X1 U17505 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14135) );
  AOI22_X1 U17506 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14134) );
  NAND4_X1 U17507 ( .A1(n14136), .A2(n14135), .A3(n14267), .A4(n14134), .ZN(
        n14137) );
  AND2_X1 U17508 ( .A1(n14138), .A2(n14137), .ZN(n14140) );
  NAND2_X1 U17509 ( .A1(n14139), .A2(n14140), .ZN(n14167) );
  OAI211_X1 U17510 ( .C1(n14139), .C2(n14140), .A(n14198), .B(n14167), .ZN(
        n14143) );
  INV_X1 U17511 ( .A(n14140), .ZN(n14141) );
  NOR2_X1 U17512 ( .A1(n19976), .A2(n14141), .ZN(n14774) );
  INV_X1 U17513 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14148) );
  INV_X1 U17514 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14147) );
  OAI22_X1 U17515 ( .A1(n14235), .A2(n14148), .B1(n14233), .B2(n14147), .ZN(
        n14151) );
  INV_X1 U17516 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14149) );
  INV_X1 U17517 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19282) );
  OAI22_X1 U17518 ( .A1(n14239), .A2(n14149), .B1(n14237), .B2(n19282), .ZN(
        n14150) );
  NOR2_X1 U17519 ( .A1(n14151), .A2(n14150), .ZN(n14154) );
  AOI22_X1 U17520 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14153) );
  AOI22_X1 U17521 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14152) );
  NAND4_X1 U17522 ( .A1(n14154), .A2(n14153), .A3(n14152), .A4(n14253), .ZN(
        n14165) );
  OAI22_X1 U17523 ( .A1(n14235), .A2(n14156), .B1(n14233), .B2(n14155), .ZN(
        n14160) );
  OAI22_X1 U17524 ( .A1(n14239), .A2(n14158), .B1(n14237), .B2(n14157), .ZN(
        n14159) );
  NOR2_X1 U17525 ( .A1(n14160), .A2(n14159), .ZN(n14163) );
  AOI22_X1 U17526 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U17527 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14161) );
  NAND4_X1 U17528 ( .A1(n14163), .A2(n14162), .A3(n14267), .A4(n14161), .ZN(
        n14164) );
  NAND2_X1 U17529 ( .A1(n14165), .A2(n14164), .ZN(n14170) );
  AOI21_X1 U17530 ( .B1(n14167), .B2(n14170), .A(n14166), .ZN(n14168) );
  OR2_X1 U17531 ( .A1(n14167), .A2(n14170), .ZN(n14197) );
  NAND2_X1 U17532 ( .A1(n14168), .A2(n14197), .ZN(n14173) );
  XNOR2_X1 U17533 ( .A(n14172), .B(n14169), .ZN(n14768) );
  INV_X1 U17534 ( .A(n14170), .ZN(n14171) );
  NAND2_X1 U17535 ( .A1(n12584), .A2(n14171), .ZN(n14770) );
  INV_X1 U17536 ( .A(n14172), .ZN(n14174) );
  INV_X1 U17537 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14177) );
  INV_X1 U17538 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14176) );
  OAI22_X1 U17539 ( .A1(n14235), .A2(n14177), .B1(n14233), .B2(n14176), .ZN(
        n14181) );
  INV_X1 U17540 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14179) );
  INV_X1 U17541 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14178) );
  OAI22_X1 U17542 ( .A1(n14239), .A2(n14179), .B1(n14237), .B2(n14178), .ZN(
        n14180) );
  NOR2_X1 U17543 ( .A1(n14181), .A2(n14180), .ZN(n14184) );
  AOI22_X1 U17544 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14183) );
  AOI22_X1 U17545 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14182) );
  NAND4_X1 U17546 ( .A1(n14184), .A2(n14183), .A3(n14182), .A4(n14253), .ZN(
        n14195) );
  INV_X1 U17547 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14186) );
  INV_X1 U17548 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14185) );
  OAI22_X1 U17549 ( .A1(n14235), .A2(n14186), .B1(n14233), .B2(n14185), .ZN(
        n14190) );
  INV_X1 U17550 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14188) );
  INV_X1 U17551 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n14187) );
  OAI22_X1 U17552 ( .A1(n14239), .A2(n14188), .B1(n14237), .B2(n14187), .ZN(
        n14189) );
  NOR2_X1 U17553 ( .A1(n14190), .A2(n14189), .ZN(n14193) );
  AOI22_X1 U17554 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14192) );
  AOI22_X1 U17555 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14191) );
  NAND4_X1 U17556 ( .A1(n14193), .A2(n14192), .A3(n14267), .A4(n14191), .ZN(
        n14194) );
  NAND2_X1 U17557 ( .A1(n14195), .A2(n14194), .ZN(n14196) );
  INV_X1 U17558 ( .A(n14196), .ZN(n14201) );
  INV_X1 U17559 ( .A(n14197), .ZN(n14199) );
  OR2_X1 U17560 ( .A1(n14197), .A2(n14196), .ZN(n14750) );
  OAI211_X1 U17561 ( .C1(n14201), .C2(n14199), .A(n14750), .B(n14198), .ZN(
        n14200) );
  OAI21_X1 U17562 ( .B1(n14175), .B2(n10102), .A(n14751), .ZN(n14758) );
  NAND2_X1 U17563 ( .A1(n12584), .A2(n14201), .ZN(n14757) );
  NOR2_X1 U17564 ( .A1(n14758), .A2(n14757), .ZN(n14756) );
  INV_X1 U17565 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14203) );
  INV_X1 U17566 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14202) );
  OAI22_X1 U17567 ( .A1(n14235), .A2(n14203), .B1(n14233), .B2(n14202), .ZN(
        n14207) );
  INV_X1 U17568 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14205) );
  OAI22_X1 U17569 ( .A1(n14239), .A2(n14205), .B1(n14237), .B2(n14204), .ZN(
        n14206) );
  NOR2_X1 U17570 ( .A1(n14207), .A2(n14206), .ZN(n14210) );
  AOI22_X1 U17571 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14209) );
  AOI22_X1 U17572 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14208) );
  NAND4_X1 U17573 ( .A1(n14210), .A2(n14209), .A3(n14208), .A4(n14253), .ZN(
        n14221) );
  OAI22_X1 U17574 ( .A1(n14235), .A2(n14212), .B1(n14233), .B2(n14211), .ZN(
        n14216) );
  OAI22_X1 U17575 ( .A1(n14239), .A2(n14214), .B1(n14237), .B2(n14213), .ZN(
        n14215) );
  NOR2_X1 U17576 ( .A1(n14216), .A2(n14215), .ZN(n14219) );
  AOI22_X1 U17577 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14218) );
  AOI22_X1 U17578 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14217) );
  NAND4_X1 U17579 ( .A1(n14219), .A2(n14218), .A3(n14267), .A4(n14217), .ZN(
        n14220) );
  AND2_X1 U17580 ( .A1(n14221), .A2(n14220), .ZN(n14752) );
  OAI21_X1 U17581 ( .B1(n14756), .B2(n14222), .A(n14752), .ZN(n14747) );
  NAND2_X1 U17582 ( .A1(n19976), .A2(n14752), .ZN(n14223) );
  NOR2_X1 U17583 ( .A1(n14750), .A2(n14223), .ZN(n14248) );
  INV_X1 U17584 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14225) );
  INV_X1 U17585 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14224) );
  OAI22_X1 U17586 ( .A1(n14235), .A2(n14225), .B1(n14233), .B2(n14224), .ZN(
        n14228) );
  INV_X1 U17587 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14226) );
  OAI22_X1 U17588 ( .A1(n14239), .A2(n14226), .B1(n14237), .B2(n19299), .ZN(
        n14227) );
  NOR2_X1 U17589 ( .A1(n14228), .A2(n14227), .ZN(n14231) );
  AOI22_X1 U17590 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14230) );
  AOI22_X1 U17591 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14229) );
  NAND4_X1 U17592 ( .A1(n14231), .A2(n14230), .A3(n14229), .A4(n14253), .ZN(
        n14246) );
  OAI22_X1 U17593 ( .A1(n14235), .A2(n14234), .B1(n14233), .B2(n14232), .ZN(
        n14241) );
  OAI22_X1 U17594 ( .A1(n14239), .A2(n14238), .B1(n14237), .B2(n14236), .ZN(
        n14240) );
  NOR2_X1 U17595 ( .A1(n14241), .A2(n14240), .ZN(n14244) );
  AOI22_X1 U17596 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14243) );
  AOI22_X1 U17597 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14242) );
  NAND4_X1 U17598 ( .A1(n14244), .A2(n14243), .A3(n14267), .A4(n14242), .ZN(
        n14245) );
  AND2_X1 U17599 ( .A1(n14246), .A2(n14245), .ZN(n14247) );
  NAND2_X1 U17600 ( .A1(n14248), .A2(n14247), .ZN(n14249) );
  OAI21_X1 U17601 ( .B1(n14248), .B2(n14247), .A(n14249), .ZN(n14746) );
  NOR2_X1 U17602 ( .A1(n14747), .A2(n14746), .ZN(n14745) );
  INV_X1 U17603 ( .A(n14249), .ZN(n14250) );
  AOI22_X1 U17604 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14252) );
  AOI22_X1 U17605 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n14251) );
  NAND2_X1 U17606 ( .A1(n14252), .A2(n14251), .ZN(n14272) );
  AOI22_X1 U17607 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U17608 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14254) );
  NAND3_X1 U17609 ( .A1(n14255), .A2(n14254), .A3(n14253), .ZN(n14271) );
  AOI22_X1 U17610 ( .A1(n14257), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14256), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14261) );
  AOI22_X1 U17611 ( .A1(n14259), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14258), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14260) );
  NAND2_X1 U17612 ( .A1(n14261), .A2(n14260), .ZN(n14270) );
  AOI22_X1 U17613 ( .A1(n14263), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14262), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14268) );
  AOI22_X1 U17614 ( .A1(n14265), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n14264), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14266) );
  NAND3_X1 U17615 ( .A1(n14268), .A2(n14267), .A3(n14266), .ZN(n14269) );
  OAI22_X1 U17616 ( .A1(n14272), .A2(n14271), .B1(n14270), .B2(n14269), .ZN(
        n14273) );
  XNOR2_X1 U17617 ( .A(n14274), .B(n14273), .ZN(n14281) );
  NOR2_X1 U17618 ( .A1(n15983), .A2(n19116), .ZN(n14275) );
  AOI21_X1 U17619 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19116), .A(n14275), .ZN(
        n14276) );
  OAI21_X1 U17620 ( .B1(n14281), .B2(n19117), .A(n14276), .ZN(P2_U2857) );
  INV_X1 U17621 ( .A(n19139), .ZN(n14277) );
  OAI22_X1 U17622 ( .A1(n14884), .A2(n14277), .B1(n19162), .B2(n13115), .ZN(
        n14278) );
  AOI21_X1 U17623 ( .B1(n15979), .B2(n19187), .A(n14278), .ZN(n14280) );
  AOI22_X1 U17624 ( .A1(n19127), .A2(BUF1_REG_30__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14279) );
  OAI211_X1 U17625 ( .C1(n14281), .C2(n19191), .A(n14280), .B(n14279), .ZN(
        P2_U2889) );
  INV_X1 U17626 ( .A(n14282), .ZN(n14290) );
  INV_X1 U17627 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21027) );
  INV_X1 U17628 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21140) );
  INV_X1 U17629 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20763) );
  AND4_X1 U17630 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .A4(n15643), .ZN(n15619) );
  AND2_X1 U17631 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15619), .ZN(n15613) );
  NAND2_X1 U17632 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15613), .ZN(n15600) );
  NOR2_X1 U17633 ( .A1(n20763), .A2(n15600), .ZN(n14374) );
  NAND2_X1 U17634 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n14374), .ZN(n14359) );
  NOR2_X1 U17635 ( .A1(n21140), .A2(n14359), .ZN(n14346) );
  NAND2_X1 U17636 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(n14346), .ZN(n14347) );
  NOR2_X1 U17637 ( .A1(n21027), .A2(n14347), .ZN(n14284) );
  AND3_X1 U17638 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n14284), .A3(n15629), 
        .ZN(n14305) );
  NAND3_X1 U17639 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .A3(n14305), .ZN(n14283) );
  NAND2_X1 U17640 ( .A1(n20062), .A2(n14283), .ZN(n14298) );
  AND2_X1 U17641 ( .A1(n15644), .A2(n14284), .ZN(n14320) );
  NAND3_X1 U17642 ( .A1(n14320), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14299) );
  INV_X1 U17643 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14510) );
  NOR3_X1 U17644 ( .A1(n14299), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14510), 
        .ZN(n14285) );
  AOI21_X1 U17645 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(n20061), .A(n14285), .ZN(
        n14287) );
  NAND2_X1 U17646 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14286) );
  OAI211_X1 U17647 ( .C1(n14298), .C2(n20965), .A(n14287), .B(n14286), .ZN(
        n14288) );
  AOI21_X1 U17648 ( .B1(n14408), .B2(n20067), .A(n14288), .ZN(n14289) );
  OAI21_X1 U17649 ( .B1(n14290), .B2(n15623), .A(n14289), .ZN(P1_U2809) );
  AOI21_X1 U17650 ( .B1(n14292), .B2(n11783), .A(n14291), .ZN(n14514) );
  INV_X1 U17651 ( .A(n14514), .ZN(n14443) );
  NAND2_X1 U17652 ( .A1(n9886), .A2(n11692), .ZN(n14295) );
  INV_X1 U17653 ( .A(n14318), .ZN(n14293) );
  AOI22_X1 U17654 ( .A1(n14295), .A2(n14294), .B1(n14293), .B2(n11669), .ZN(
        n14297) );
  XNOR2_X1 U17655 ( .A(n14297), .B(n14296), .ZN(n14646) );
  AOI21_X1 U17656 ( .B1(n14510), .B2(n14299), .A(n14298), .ZN(n14302) );
  AOI22_X1 U17657 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n20061), .ZN(n14300) );
  OAI21_X1 U17658 ( .B1(n20063), .B2(n14512), .A(n14300), .ZN(n14301) );
  AOI211_X1 U17659 ( .C1(n14646), .C2(n20067), .A(n14302), .B(n14301), .ZN(
        n14303) );
  OAI21_X1 U17660 ( .B1(n14443), .B2(n15623), .A(n14303), .ZN(P1_U2810) );
  NOR2_X1 U17661 ( .A1(n20016), .A2(n14305), .ZN(n14319) );
  INV_X1 U17662 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14523) );
  NOR2_X1 U17663 ( .A1(n14523), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14306) );
  AOI22_X1 U17664 ( .A1(n14320), .A2(n14306), .B1(n20046), .B2(
        P1_EBX_REG_29__SCAN_IN), .ZN(n14309) );
  NAND2_X1 U17665 ( .A1(n20053), .A2(n14307), .ZN(n14308) );
  OAI211_X1 U17666 ( .C1(n20064), .C2(n14310), .A(n14309), .B(n14308), .ZN(
        n14313) );
  XNOR2_X1 U17667 ( .A(n14318), .B(n14311), .ZN(n14654) );
  NOR2_X1 U17668 ( .A1(n14654), .A2(n20049), .ZN(n14312) );
  AOI211_X1 U17669 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(n14319), .A(n14313), 
        .B(n14312), .ZN(n14314) );
  OAI21_X1 U17670 ( .B1(n14304), .B2(n15623), .A(n14314), .ZN(P1_U2811) );
  AOI21_X1 U17671 ( .B1(n14315), .B2(n9860), .A(n10233), .ZN(n14527) );
  INV_X1 U17672 ( .A(n14527), .ZN(n14450) );
  NOR2_X1 U17673 ( .A1(n14331), .A2(n14316), .ZN(n14317) );
  NOR2_X1 U17674 ( .A1(n14318), .A2(n14317), .ZN(n14663) );
  INV_X1 U17675 ( .A(n14319), .ZN(n14322) );
  NOR2_X1 U17676 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(n14320), .ZN(n14321) );
  NOR2_X1 U17677 ( .A1(n14322), .A2(n14321), .ZN(n14325) );
  AOI22_X1 U17678 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n20046), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n14323) );
  OAI21_X1 U17679 ( .B1(n20063), .B2(n14525), .A(n14323), .ZN(n14324) );
  AOI211_X1 U17680 ( .C1(n14663), .C2(n20067), .A(n14325), .B(n14324), .ZN(
        n14326) );
  OAI21_X1 U17681 ( .B1(n14450), .B2(n15623), .A(n14326), .ZN(P1_U2812) );
  NAND2_X1 U17682 ( .A1(n14339), .A2(n14327), .ZN(n14328) );
  NOR2_X1 U17683 ( .A1(n14341), .A2(n14329), .ZN(n14330) );
  OR2_X1 U17684 ( .A1(n14331), .A2(n14330), .ZN(n14672) );
  INV_X1 U17685 ( .A(n14672), .ZN(n14337) );
  AOI21_X1 U17686 ( .B1(n15644), .B2(n14347), .A(n14332), .ZN(n14345) );
  NOR3_X1 U17687 ( .A1(n15630), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14347), 
        .ZN(n14333) );
  AOI21_X1 U17688 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n20061), .A(n14333), .ZN(
        n14335) );
  AOI22_X1 U17689 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n20024), .B1(
        n20053), .B2(n14532), .ZN(n14334) );
  OAI211_X1 U17690 ( .C1(n14345), .C2(n21027), .A(n14335), .B(n14334), .ZN(
        n14336) );
  AOI21_X1 U17691 ( .B1(n14337), .B2(n20067), .A(n14336), .ZN(n14338) );
  OAI21_X1 U17692 ( .B1(n14454), .B2(n15623), .A(n14338), .ZN(P1_U2813) );
  OAI21_X1 U17693 ( .B1(n14353), .B2(n14340), .A(n14339), .ZN(n14541) );
  AOI21_X1 U17694 ( .B1(n14342), .B2(n14357), .A(n14341), .ZN(n15791) );
  INV_X1 U17695 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14344) );
  OAI22_X1 U17696 ( .A1(n14345), .A2(n14344), .B1(n14343), .B2(n20064), .ZN(
        n14351) );
  NAND2_X1 U17697 ( .A1(n20061), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n14349) );
  NAND3_X1 U17698 ( .A1(n14347), .A2(n14346), .A3(n15644), .ZN(n14348) );
  OAI211_X1 U17699 ( .C1(n20063), .C2(n14543), .A(n14349), .B(n14348), .ZN(
        n14350) );
  AOI211_X1 U17700 ( .C1(n15791), .C2(n20067), .A(n14351), .B(n14350), .ZN(
        n14352) );
  OAI21_X1 U17701 ( .B1(n14541), .B2(n15623), .A(n14352), .ZN(P1_U2814) );
  INV_X1 U17702 ( .A(n14353), .ZN(n14354) );
  OAI21_X1 U17703 ( .B1(n14355), .B2(n9837), .A(n14354), .ZN(n14561) );
  INV_X1 U17704 ( .A(n14356), .ZN(n14370) );
  OAI21_X1 U17705 ( .B1(n14370), .B2(n14358), .A(n14357), .ZN(n14684) );
  INV_X1 U17706 ( .A(n14684), .ZN(n14366) );
  INV_X1 U17707 ( .A(n14559), .ZN(n14364) );
  NOR3_X1 U17708 ( .A1(n15630), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n14359), 
        .ZN(n14361) );
  NOR2_X1 U17709 ( .A1(n20064), .A2(n14554), .ZN(n14360) );
  AOI211_X1 U17710 ( .C1(n20046), .C2(P1_EBX_REG_25__SCAN_IN), .A(n14361), .B(
        n14360), .ZN(n14363) );
  OAI21_X1 U17711 ( .B1(n14374), .B2(n15630), .A(n15629), .ZN(n15602) );
  NOR2_X1 U17712 ( .A1(n15630), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14373) );
  OAI21_X1 U17713 ( .B1(n15602), .B2(n14373), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14362) );
  OAI211_X1 U17714 ( .C1(n20063), .C2(n14364), .A(n14363), .B(n14362), .ZN(
        n14365) );
  AOI21_X1 U17715 ( .B1(n14366), .B2(n20067), .A(n14365), .ZN(n14367) );
  OAI21_X1 U17716 ( .B1(n14561), .B2(n15623), .A(n14367), .ZN(P1_U2815) );
  INV_X1 U17717 ( .A(n14368), .ZN(n14417) );
  AOI21_X1 U17718 ( .B1(n14369), .B2(n14417), .A(n9837), .ZN(n14569) );
  INV_X1 U17719 ( .A(n14569), .ZN(n14468) );
  AOI21_X1 U17720 ( .B1(n14371), .B2(n14421), .A(n14370), .ZN(n14686) );
  INV_X1 U17721 ( .A(n14372), .ZN(n14567) );
  NOR2_X1 U17722 ( .A1(n20063), .A2(n14567), .ZN(n14379) );
  AOI22_X1 U17723 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15602), .B1(n14374), 
        .B2(n14373), .ZN(n14376) );
  NAND2_X1 U17724 ( .A1(n20046), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14375) );
  OAI211_X1 U17725 ( .C1(n20064), .C2(n14377), .A(n14376), .B(n14375), .ZN(
        n14378) );
  AOI211_X1 U17726 ( .C1(n14686), .C2(n20067), .A(n14379), .B(n14378), .ZN(
        n14380) );
  OAI21_X1 U17727 ( .B1(n14468), .B2(n15623), .A(n14380), .ZN(P1_U2816) );
  AOI21_X1 U17728 ( .B1(n14383), .B2(n14381), .A(n14382), .ZN(n15729) );
  INV_X1 U17729 ( .A(n15729), .ZN(n14486) );
  OAI21_X1 U17730 ( .B1(n15619), .B2(n15630), .A(n15629), .ZN(n15620) );
  INV_X1 U17731 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20891) );
  NAND3_X1 U17732 ( .A1(n15644), .A2(P1_REIP_REG_18__SCAN_IN), .A3(n15643), 
        .ZN(n15633) );
  INV_X1 U17733 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n21026) );
  OAI21_X1 U17734 ( .B1(n20891), .B2(n15633), .A(n21026), .ZN(n14389) );
  OR2_X1 U17735 ( .A1(n14436), .A2(n14384), .ZN(n14385) );
  AND2_X1 U17736 ( .A1(n9894), .A2(n14385), .ZN(n15571) );
  AOI22_X1 U17737 ( .A1(n15571), .A2(n20067), .B1(n20046), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14387) );
  NAND2_X1 U17738 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14386) );
  OAI211_X1 U17739 ( .C1(n20063), .C2(n15727), .A(n14387), .B(n14386), .ZN(
        n14388) );
  AOI21_X1 U17740 ( .B1(n15620), .B2(n14389), .A(n14388), .ZN(n14390) );
  OAI21_X1 U17741 ( .B1(n14486), .B2(n15623), .A(n14390), .ZN(P1_U2820) );
  INV_X1 U17742 ( .A(n14391), .ZN(n14394) );
  INV_X1 U17743 ( .A(n14392), .ZN(n14393) );
  AOI21_X1 U17744 ( .B1(n14395), .B2(n14394), .A(n14393), .ZN(n14633) );
  INV_X1 U17745 ( .A(n14633), .ZN(n14506) );
  INV_X1 U17746 ( .A(n14631), .ZN(n14406) );
  AOI21_X1 U17747 ( .B1(n14396), .B2(n15686), .A(n15674), .ZN(n15870) );
  AOI22_X1 U17748 ( .A1(n15870), .A2(n20067), .B1(n20046), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14397) );
  OAI211_X1 U17749 ( .C1(n20064), .C2(n14398), .A(n14397), .B(n20135), .ZN(
        n14405) );
  NAND2_X1 U17750 ( .A1(n14400), .A2(n14399), .ZN(n15684) );
  NOR2_X1 U17751 ( .A1(n14401), .A2(n15684), .ZN(n14403) );
  AOI21_X1 U17752 ( .B1(n14401), .B2(n20062), .A(n15702), .ZN(n15695) );
  INV_X1 U17753 ( .A(n15695), .ZN(n14402) );
  MUX2_X1 U17754 ( .A(n14403), .B(n14402), .S(P1_REIP_REG_13__SCAN_IN), .Z(
        n14404) );
  AOI211_X1 U17755 ( .C1(n20053), .C2(n14406), .A(n14405), .B(n14404), .ZN(
        n14407) );
  OAI21_X1 U17756 ( .B1(n14506), .B2(n15623), .A(n14407), .ZN(P1_U2827) );
  INV_X1 U17757 ( .A(n14408), .ZN(n14410) );
  INV_X1 U17758 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14409) );
  OAI22_X1 U17759 ( .A1(n14410), .A2(n15712), .B1(n14409), .B2(n20078), .ZN(
        P1_U2841) );
  INV_X1 U17760 ( .A(n14646), .ZN(n14411) );
  INV_X1 U17761 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n21128) );
  OAI222_X1 U17762 ( .A1(n14439), .A2(n14443), .B1(n15712), .B2(n14411), .C1(
        n21128), .C2(n20078), .ZN(P1_U2842) );
  OAI222_X1 U17763 ( .A1(n20990), .A2(n20078), .B1(n15712), .B2(n14654), .C1(
        n14439), .C2(n14304), .ZN(P1_U2843) );
  INV_X1 U17764 ( .A(n14663), .ZN(n14412) );
  OAI222_X1 U17765 ( .A1(n20945), .A2(n20078), .B1(n15712), .B2(n14412), .C1(
        n14450), .C2(n14439), .ZN(P1_U2844) );
  INV_X1 U17766 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14413) );
  OAI222_X1 U17767 ( .A1(n14413), .A2(n20078), .B1(n15712), .B2(n14672), .C1(
        n14454), .C2(n14439), .ZN(P1_U2845) );
  INV_X1 U17768 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n21167) );
  INV_X1 U17769 ( .A(n15791), .ZN(n14414) );
  OAI222_X1 U17770 ( .A1(n21167), .A2(n20078), .B1(n15712), .B2(n14414), .C1(
        n14541), .C2(n14439), .ZN(P1_U2846) );
  INV_X1 U17771 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n20992) );
  OAI222_X1 U17772 ( .A1(n14684), .A2(n15712), .B1(n20078), .B2(n20992), .C1(
        n14439), .C2(n14561), .ZN(P1_U2847) );
  INV_X1 U17773 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n21121) );
  INV_X1 U17774 ( .A(n14686), .ZN(n14415) );
  OAI222_X1 U17775 ( .A1(n14439), .A2(n14468), .B1(n20078), .B2(n21121), .C1(
        n14415), .C2(n15712), .ZN(P1_U2848) );
  AOI21_X1 U17776 ( .B1(n14418), .B2(n14416), .A(n14368), .ZN(n14573) );
  INV_X1 U17777 ( .A(n14573), .ZN(n15604) );
  INV_X1 U17778 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n21020) );
  OR2_X1 U17779 ( .A1(n15611), .A2(n14419), .ZN(n14420) );
  NAND2_X1 U17780 ( .A1(n14421), .A2(n14420), .ZN(n15603) );
  OAI222_X1 U17781 ( .A1(n14439), .A2(n15604), .B1(n20078), .B2(n21020), .C1(
        n15603), .C2(n15712), .ZN(P1_U2849) );
  INV_X1 U17782 ( .A(n14422), .ZN(n14423) );
  OAI21_X1 U17783 ( .B1(n14424), .B2(n14382), .A(n14423), .ZN(n15624) );
  NAND2_X1 U17784 ( .A1(n9894), .A2(n14425), .ZN(n14426) );
  NAND2_X1 U17785 ( .A1(n9836), .A2(n14426), .ZN(n15628) );
  OAI22_X1 U17786 ( .A1(n15628), .A2(n15712), .B1(n14427), .B2(n20078), .ZN(
        n14428) );
  INV_X1 U17787 ( .A(n14428), .ZN(n14429) );
  OAI21_X1 U17788 ( .B1(n15624), .B2(n14439), .A(n14429), .ZN(P1_U2851) );
  AOI22_X1 U17789 ( .A1(n15571), .A2(n20073), .B1(n14437), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14430) );
  OAI21_X1 U17790 ( .B1(n14486), .B2(n14439), .A(n14430), .ZN(P1_U2852) );
  NAND2_X1 U17791 ( .A1(n14431), .A2(n14432), .ZN(n14433) );
  INV_X1 U17792 ( .A(n15638), .ZN(n14491) );
  INV_X1 U17793 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21125) );
  NOR2_X1 U17794 ( .A1(n15648), .A2(n14434), .ZN(n14435) );
  OR2_X1 U17795 ( .A1(n14436), .A2(n14435), .ZN(n15641) );
  OAI222_X1 U17796 ( .A1(n14439), .A2(n14491), .B1(n20078), .B2(n21125), .C1(
        n15641), .C2(n15712), .ZN(P1_U2853) );
  AOI22_X1 U17797 ( .A1(n15870), .A2(n20073), .B1(n14437), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14438) );
  OAI21_X1 U17798 ( .B1(n14506), .B2(n14439), .A(n14438), .ZN(P1_U2859) );
  AOI22_X1 U17799 ( .A1(n14488), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14487), .ZN(n14442) );
  AOI22_X1 U17800 ( .A1(n14496), .A2(DATAI_30_), .B1(n14495), .B2(n14440), 
        .ZN(n14441) );
  OAI211_X1 U17801 ( .C1(n14443), .C2(n14499), .A(n14442), .B(n14441), .ZN(
        P1_U2874) );
  AOI22_X1 U17802 ( .A1(n14488), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14487), .ZN(n14445) );
  AOI22_X1 U17803 ( .A1(n14496), .A2(DATAI_29_), .B1(n14495), .B2(n14501), 
        .ZN(n14444) );
  OAI211_X1 U17804 ( .C1(n14304), .C2(n14499), .A(n14445), .B(n14444), .ZN(
        P1_U2875) );
  NOR2_X1 U17805 ( .A1(n14493), .A2(n16379), .ZN(n14448) );
  INV_X1 U17806 ( .A(n14496), .ZN(n14458) );
  INV_X1 U17807 ( .A(n14495), .ZN(n14455) );
  OAI22_X1 U17808 ( .A1(n14458), .A2(n21166), .B1(n14446), .B2(n14455), .ZN(
        n14447) );
  AOI211_X1 U17809 ( .C1(n14487), .C2(P1_EAX_REG_28__SCAN_IN), .A(n14448), .B(
        n14447), .ZN(n14449) );
  OAI21_X1 U17810 ( .B1(n14450), .B2(n14499), .A(n14449), .ZN(P1_U2876) );
  AOI22_X1 U17811 ( .A1(n14488), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14487), .ZN(n14453) );
  AOI22_X1 U17812 ( .A1(n14496), .A2(DATAI_27_), .B1(n14495), .B2(n14451), 
        .ZN(n14452) );
  OAI211_X1 U17813 ( .C1(n14454), .C2(n14499), .A(n14453), .B(n14452), .ZN(
        P1_U2877) );
  INV_X1 U17814 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20161) );
  NOR2_X1 U17815 ( .A1(n14493), .A2(n20161), .ZN(n14460) );
  INV_X1 U17816 ( .A(DATAI_26_), .ZN(n14457) );
  OAI22_X1 U17817 ( .A1(n14458), .A2(n14457), .B1(n14456), .B2(n14455), .ZN(
        n14459) );
  AOI211_X1 U17818 ( .C1(n14487), .C2(P1_EAX_REG_26__SCAN_IN), .A(n14460), .B(
        n14459), .ZN(n14461) );
  OAI21_X1 U17819 ( .B1(n14541), .B2(n14499), .A(n14461), .ZN(P1_U2878) );
  AOI22_X1 U17820 ( .A1(n14488), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14487), .ZN(n14464) );
  AOI22_X1 U17821 ( .A1(n14496), .A2(DATAI_25_), .B1(n14495), .B2(n14462), 
        .ZN(n14463) );
  OAI211_X1 U17822 ( .C1(n14561), .C2(n14499), .A(n14464), .B(n14463), .ZN(
        P1_U2879) );
  AOI22_X1 U17823 ( .A1(n14488), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14487), .ZN(n14467) );
  AOI22_X1 U17824 ( .A1(n14496), .A2(DATAI_24_), .B1(n14495), .B2(n14465), 
        .ZN(n14466) );
  OAI211_X1 U17825 ( .C1(n14468), .C2(n14499), .A(n14467), .B(n14466), .ZN(
        P1_U2880) );
  AOI22_X1 U17826 ( .A1(n14488), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14487), .ZN(n14471) );
  AOI22_X1 U17827 ( .A1(n14496), .A2(DATAI_23_), .B1(n14495), .B2(n14469), 
        .ZN(n14470) );
  OAI211_X1 U17828 ( .C1(n15604), .C2(n14499), .A(n14471), .B(n14470), .ZN(
        P1_U2881) );
  OR2_X1 U17829 ( .A1(n14422), .A2(n14472), .ZN(n14473) );
  AND2_X1 U17830 ( .A1(n14473), .A2(n14416), .ZN(n15723) );
  INV_X1 U17831 ( .A(n15723), .ZN(n14478) );
  INV_X1 U17832 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n20185) );
  OAI22_X1 U17833 ( .A1(n14493), .A2(n20185), .B1(n14474), .B2(n14502), .ZN(
        n14475) );
  INV_X1 U17834 ( .A(n14475), .ZN(n14477) );
  AOI22_X1 U17835 ( .A1(n14496), .A2(DATAI_22_), .B1(n14495), .B2(n20183), 
        .ZN(n14476) );
  OAI211_X1 U17836 ( .C1(n14478), .C2(n14499), .A(n14477), .B(n14476), .ZN(
        P1_U2882) );
  AOI22_X1 U17837 ( .A1(n14488), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14487), .ZN(n14480) );
  AOI22_X1 U17838 ( .A1(n14496), .A2(DATAI_21_), .B1(n14495), .B2(n20175), 
        .ZN(n14479) );
  OAI211_X1 U17839 ( .C1(n15624), .C2(n14499), .A(n14480), .B(n14479), .ZN(
        P1_U2883) );
  OAI22_X1 U17840 ( .A1(n14493), .A2(n16389), .B1(n14481), .B2(n14502), .ZN(
        n14482) );
  INV_X1 U17841 ( .A(n14482), .ZN(n14485) );
  AOI22_X1 U17842 ( .A1(n14496), .A2(DATAI_20_), .B1(n14495), .B2(n14483), 
        .ZN(n14484) );
  OAI211_X1 U17843 ( .C1(n14486), .C2(n14499), .A(n14485), .B(n14484), .ZN(
        P1_U2884) );
  AOI22_X1 U17844 ( .A1(n14488), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14487), .ZN(n14490) );
  AOI22_X1 U17845 ( .A1(n14496), .A2(DATAI_19_), .B1(n14495), .B2(n20169), 
        .ZN(n14489) );
  OAI211_X1 U17846 ( .C1(n14491), .C2(n14499), .A(n14490), .B(n14489), .ZN(
        P1_U2885) );
  INV_X1 U17847 ( .A(n14431), .ZN(n14492) );
  INV_X1 U17848 ( .A(n15708), .ZN(n14500) );
  INV_X1 U17849 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20163) );
  OAI22_X1 U17850 ( .A1(n14493), .A2(n20163), .B1(n13170), .B2(n14502), .ZN(
        n14494) );
  INV_X1 U17851 ( .A(n14494), .ZN(n14498) );
  AOI22_X1 U17852 ( .A1(n14496), .A2(DATAI_18_), .B1(n14495), .B2(n20162), 
        .ZN(n14497) );
  OAI211_X1 U17853 ( .C1(n14500), .C2(n14499), .A(n14498), .B(n14497), .ZN(
        P1_U2886) );
  INV_X1 U17854 ( .A(n14501), .ZN(n14505) );
  OAI222_X1 U17855 ( .A1(n14499), .A2(n14506), .B1(n14505), .B2(n14504), .C1(
        n14503), .C2(n14502), .ZN(P1_U2891) );
  NAND2_X1 U17856 ( .A1(n14508), .A2(n14507), .ZN(n14509) );
  XNOR2_X1 U17857 ( .A(n14509), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14652) );
  NOR2_X1 U17858 ( .A1(n20135), .A2(n14510), .ZN(n14645) );
  AOI21_X1 U17859 ( .B1(n20125), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14645), .ZN(n14511) );
  OAI21_X1 U17860 ( .B1(n15782), .B2(n14512), .A(n14511), .ZN(n14513) );
  AOI21_X1 U17861 ( .B1(n14514), .B2(n15786), .A(n14513), .ZN(n14515) );
  OAI21_X1 U17862 ( .B1(n14652), .B2(n19996), .A(n14515), .ZN(P1_U2969) );
  NAND2_X1 U17863 ( .A1(n9820), .A2(n15796), .ZN(n14538) );
  NAND2_X1 U17864 ( .A1(n14572), .A2(n14538), .ZN(n14521) );
  NAND2_X1 U17865 ( .A1(n14516), .A2(n11606), .ZN(n14517) );
  OAI21_X1 U17866 ( .B1(n14518), .B2(n14517), .A(n14521), .ZN(n14520) );
  MUX2_X1 U17867 ( .A(n14675), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9820), .Z(n14519) );
  OAI211_X1 U17868 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14521), .A(
        n14520), .B(n14519), .ZN(n14522) );
  XNOR2_X1 U17869 ( .A(n14522), .B(n14660), .ZN(n14669) );
  NOR2_X1 U17870 ( .A1(n20135), .A2(n14523), .ZN(n14662) );
  AOI21_X1 U17871 ( .B1(n20125), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14662), .ZN(n14524) );
  OAI21_X1 U17872 ( .B1(n15782), .B2(n14525), .A(n14524), .ZN(n14526) );
  AOI21_X1 U17873 ( .B1(n14527), .B2(n15786), .A(n14526), .ZN(n14528) );
  OAI21_X1 U17874 ( .B1(n19996), .B2(n14669), .A(n14528), .ZN(P1_U2971) );
  MUX2_X1 U17875 ( .A(n14530), .B(n14529), .S(n9820), .Z(n14531) );
  XNOR2_X1 U17876 ( .A(n14531), .B(n14675), .ZN(n14678) );
  INV_X1 U17877 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U17878 ( .A1(n15783), .A2(n14532), .ZN(n14533) );
  NAND2_X1 U17879 ( .A1(n15935), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14671) );
  OAI211_X1 U17880 ( .C1(n15790), .C2(n14534), .A(n14533), .B(n14671), .ZN(
        n14535) );
  AOI21_X1 U17881 ( .B1(n14536), .B2(n15786), .A(n14535), .ZN(n14537) );
  OAI21_X1 U17882 ( .B1(n14678), .B2(n19996), .A(n14537), .ZN(P1_U2972) );
  OAI211_X1 U17883 ( .C1(n14587), .C2(n14572), .A(n14539), .B(n14538), .ZN(
        n14540) );
  XNOR2_X1 U17884 ( .A(n14540), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15792) );
  INV_X1 U17885 ( .A(n15792), .ZN(n14547) );
  INV_X1 U17886 ( .A(n14541), .ZN(n14545) );
  AOI22_X1 U17887 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n15899), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n14542) );
  OAI21_X1 U17888 ( .B1(n15782), .B2(n14543), .A(n14542), .ZN(n14544) );
  AOI21_X1 U17889 ( .B1(n14545), .B2(n15786), .A(n14544), .ZN(n14546) );
  OAI21_X1 U17890 ( .B1(n14547), .B2(n19996), .A(n14546), .ZN(P1_U2973) );
  NAND2_X1 U17891 ( .A1(n14548), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14564) );
  NOR2_X1 U17892 ( .A1(n14689), .A2(n14564), .ZN(n14549) );
  XNOR2_X1 U17893 ( .A(n14553), .B(n14552), .ZN(n14681) );
  OR2_X1 U17894 ( .A1(n15790), .A2(n14554), .ZN(n14555) );
  NAND2_X1 U17895 ( .A1(n15935), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14679) );
  AND2_X1 U17896 ( .A1(n14555), .A2(n14679), .ZN(n14556) );
  AOI21_X1 U17897 ( .B1(n14559), .B2(n15783), .A(n14558), .ZN(n14560) );
  OAI21_X1 U17898 ( .B1(n14561), .B2(n20131), .A(n14560), .ZN(P1_U2974) );
  NAND2_X1 U17899 ( .A1(n14562), .A2(n14564), .ZN(n14563) );
  MUX2_X1 U17900 ( .A(n14564), .B(n14563), .S(n14587), .Z(n14565) );
  XNOR2_X1 U17901 ( .A(n14565), .B(n14689), .ZN(n14694) );
  AND2_X1 U17902 ( .A1(n15899), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14685) );
  AOI21_X1 U17903 ( .B1(n20125), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14685), .ZN(n14566) );
  OAI21_X1 U17904 ( .B1(n15782), .B2(n14567), .A(n14566), .ZN(n14568) );
  AOI21_X1 U17905 ( .B1(n14569), .B2(n15786), .A(n14568), .ZN(n14570) );
  OAI21_X1 U17906 ( .B1(n14694), .B2(n19996), .A(n14570), .ZN(P1_U2975) );
  XNOR2_X1 U17907 ( .A(n9820), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14571) );
  XNOR2_X1 U17908 ( .A(n14572), .B(n14571), .ZN(n14701) );
  NAND2_X1 U17909 ( .A1(n14573), .A2(n15786), .ZN(n14576) );
  OAI22_X1 U17910 ( .A1(n15790), .A2(n15609), .B1(n20135), .B2(n20763), .ZN(
        n14574) );
  AOI21_X1 U17911 ( .B1(n15783), .B2(n15606), .A(n14574), .ZN(n14575) );
  OAI211_X1 U17912 ( .C1(n14701), .C2(n19996), .A(n14576), .B(n14575), .ZN(
        P1_U2976) );
  NOR3_X1 U17913 ( .A1(n14577), .A2(n14587), .A3(n14708), .ZN(n14580) );
  NOR3_X1 U17914 ( .A1(n14578), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n14586), .ZN(n14579) );
  NOR2_X1 U17915 ( .A1(n14580), .A2(n14579), .ZN(n15568) );
  NOR2_X1 U17916 ( .A1(n15568), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15567) );
  AOI22_X1 U17917 ( .A1(n15567), .A2(n14587), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14580), .ZN(n14582) );
  XNOR2_X1 U17918 ( .A(n14582), .B(n14581), .ZN(n14706) );
  NAND2_X1 U17919 ( .A1(n15935), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14702) );
  OAI21_X1 U17920 ( .B1(n15790), .B2(n10886), .A(n14702), .ZN(n14584) );
  NOR2_X1 U17921 ( .A1(n15624), .A2(n20131), .ZN(n14583) );
  AOI211_X1 U17922 ( .C1(n15783), .C2(n15626), .A(n14584), .B(n14583), .ZN(
        n14585) );
  OAI21_X1 U17923 ( .B1(n14706), .B2(n19996), .A(n14585), .ZN(P1_U2978) );
  MUX2_X1 U17924 ( .A(n14587), .B(n14586), .S(n14577), .Z(n14588) );
  XNOR2_X1 U17925 ( .A(n14588), .B(n14708), .ZN(n14712) );
  INV_X1 U17926 ( .A(n15632), .ZN(n14590) );
  AOI22_X1 U17927 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n15899), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14589) );
  OAI21_X1 U17928 ( .B1(n15782), .B2(n14590), .A(n14589), .ZN(n14591) );
  AOI21_X1 U17929 ( .B1(n15638), .B2(n15786), .A(n14591), .ZN(n14592) );
  OAI21_X1 U17930 ( .B1(n14712), .B2(n19996), .A(n14592), .ZN(P1_U2980) );
  OAI21_X1 U17931 ( .B1(n14578), .B2(n14593), .A(n14577), .ZN(n15828) );
  AOI22_X1 U17932 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n15899), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n14594) );
  OAI21_X1 U17933 ( .B1(n15782), .B2(n15656), .A(n14594), .ZN(n14595) );
  AOI21_X1 U17934 ( .B1(n15708), .B2(n15786), .A(n14595), .ZN(n14596) );
  OAI21_X1 U17935 ( .B1(n15828), .B2(n19996), .A(n14596), .ZN(P1_U2981) );
  NAND2_X1 U17936 ( .A1(n14587), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15753) );
  NAND2_X1 U17937 ( .A1(n14587), .A2(n14598), .ZN(n14624) );
  NAND3_X1 U17938 ( .A1(n14597), .A2(n15753), .A3(n14624), .ZN(n15745) );
  INV_X1 U17939 ( .A(n14599), .ZN(n14614) );
  AOI21_X1 U17940 ( .B1(n15863), .B2(n15878), .A(n9820), .ZN(n14600) );
  AOI211_X1 U17941 ( .C1(n15745), .C2(n9870), .A(n14614), .B(n14600), .ZN(
        n14602) );
  NOR2_X1 U17942 ( .A1(n14602), .A2(n14601), .ZN(n14604) );
  NOR2_X1 U17943 ( .A1(n14604), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14603) );
  MUX2_X1 U17944 ( .A(n14604), .B(n14603), .S(n14587), .Z(n14606) );
  XNOR2_X1 U17945 ( .A(n14606), .B(n14605), .ZN(n15838) );
  NAND2_X1 U17946 ( .A1(n15838), .A2(n20127), .ZN(n14611) );
  OAI22_X1 U17947 ( .A1(n15790), .A2(n14607), .B1(n20135), .B2(n20754), .ZN(
        n14608) );
  AOI21_X1 U17948 ( .B1(n15783), .B2(n14609), .A(n14608), .ZN(n14610) );
  OAI211_X1 U17949 ( .C1(n20131), .C2(n14612), .A(n14611), .B(n14610), .ZN(
        P1_U2982) );
  INV_X1 U17950 ( .A(n14613), .ZN(n15733) );
  NOR2_X1 U17951 ( .A1(n15733), .A2(n14614), .ZN(n14617) );
  AND2_X1 U17952 ( .A1(n15735), .A2(n14615), .ZN(n14616) );
  XNOR2_X1 U17953 ( .A(n14617), .B(n14616), .ZN(n15857) );
  INV_X1 U17954 ( .A(n15857), .ZN(n14618) );
  NAND2_X1 U17955 ( .A1(n15935), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n15854) );
  OAI21_X1 U17956 ( .B1(n19996), .B2(n14618), .A(n15854), .ZN(n14621) );
  NOR2_X1 U17957 ( .A1(n15782), .A2(n14619), .ZN(n14620) );
  AOI211_X1 U17958 ( .C1(n20125), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n14621), .B(n14620), .ZN(n14622) );
  OAI21_X1 U17959 ( .B1(n14623), .B2(n20131), .A(n14622), .ZN(P1_U2984) );
  INV_X1 U17960 ( .A(n14597), .ZN(n15762) );
  INV_X1 U17961 ( .A(n14624), .ZN(n14625) );
  AOI21_X1 U17962 ( .B1(n15762), .B2(n14626), .A(n14625), .ZN(n15752) );
  OAI211_X1 U17963 ( .C1(n14627), .C2(n9820), .A(n15752), .B(n15754), .ZN(
        n15755) );
  NAND2_X1 U17964 ( .A1(n15755), .A2(n15754), .ZN(n14629) );
  XNOR2_X1 U17965 ( .A(n14629), .B(n14628), .ZN(n15869) );
  AOI22_X1 U17966 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n15899), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14630) );
  OAI21_X1 U17967 ( .B1(n15782), .B2(n14631), .A(n14630), .ZN(n14632) );
  AOI21_X1 U17968 ( .B1(n14633), .B2(n15786), .A(n14632), .ZN(n14634) );
  OAI21_X1 U17969 ( .B1(n15869), .B2(n19996), .A(n14634), .ZN(P1_U2986) );
  INV_X1 U17970 ( .A(n14635), .ZN(n14642) );
  NAND2_X1 U17971 ( .A1(n15899), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n15908) );
  MUX2_X1 U17972 ( .A(n15765), .B(n14597), .S(n9820), .Z(n14637) );
  INV_X1 U17973 ( .A(n14637), .ZN(n14638) );
  XNOR2_X1 U17974 ( .A(n14638), .B(n15763), .ZN(n15911) );
  NAND2_X1 U17975 ( .A1(n20127), .A2(n15911), .ZN(n14639) );
  OAI211_X1 U17976 ( .C1(n15790), .C2(n14640), .A(n15908), .B(n14639), .ZN(
        n14641) );
  AOI21_X1 U17977 ( .B1(n14642), .B2(n15783), .A(n14641), .ZN(n14643) );
  OAI21_X1 U17978 ( .B1(n14644), .B2(n20131), .A(n14643), .ZN(P1_U2989) );
  AOI21_X1 U17979 ( .B1(n14646), .B2(n15932), .A(n14645), .ZN(n14651) );
  INV_X1 U17980 ( .A(n14647), .ZN(n14648) );
  OAI21_X1 U17981 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14649), .A(
        n14648), .ZN(n14650) );
  OAI211_X1 U17982 ( .C1(n14652), .C2(n20138), .A(n14651), .B(n14650), .ZN(
        P1_U3001) );
  OAI21_X1 U17983 ( .B1(n14654), .B2(n20137), .A(n14653), .ZN(n14656) );
  NOR3_X1 U17984 ( .A1(n14664), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14666), .ZN(n14655) );
  AOI211_X1 U17985 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14657), .A(
        n14656), .B(n14655), .ZN(n14658) );
  OAI21_X1 U17986 ( .B1(n14659), .B2(n20138), .A(n14658), .ZN(P1_U3002) );
  NOR2_X1 U17987 ( .A1(n14670), .A2(n14660), .ZN(n14661) );
  AOI211_X1 U17988 ( .C1(n15932), .C2(n14663), .A(n14662), .B(n14661), .ZN(
        n14668) );
  INV_X1 U17989 ( .A(n14664), .ZN(n14676) );
  NAND3_X1 U17990 ( .A1(n14676), .A2(n14666), .A3(n14665), .ZN(n14667) );
  OAI211_X1 U17991 ( .C1(n14669), .C2(n20138), .A(n14668), .B(n14667), .ZN(
        P1_U3003) );
  NOR2_X1 U17992 ( .A1(n14670), .A2(n14675), .ZN(n14674) );
  OAI21_X1 U17993 ( .B1(n14672), .B2(n20137), .A(n14671), .ZN(n14673) );
  AOI211_X1 U17994 ( .C1(n14676), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14677) );
  OAI21_X1 U17995 ( .B1(n14678), .B2(n20138), .A(n14677), .ZN(P1_U3004) );
  NAND2_X1 U17996 ( .A1(n15793), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14683) );
  INV_X1 U17997 ( .A(n14679), .ZN(n14680) );
  NOR3_X1 U17998 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14687), .A3(
        n15795), .ZN(n15794) );
  AOI211_X1 U17999 ( .C1(n15933), .C2(n14681), .A(n14680), .B(n15794), .ZN(
        n14682) );
  OAI211_X1 U18000 ( .C1(n14684), .C2(n20137), .A(n14683), .B(n14682), .ZN(
        P1_U3006) );
  AOI21_X1 U18001 ( .B1(n14686), .B2(n15932), .A(n14685), .ZN(n14693) );
  OAI21_X1 U18002 ( .B1(n20143), .B2(n14688), .A(n14687), .ZN(n14690) );
  AOI22_X1 U18003 ( .A1(n14695), .A2(n14690), .B1(n14689), .B2(n15795), .ZN(
        n14691) );
  OAI21_X1 U18004 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n14691), .ZN(n14692) );
  OAI211_X1 U18005 ( .C1(n14694), .C2(n20138), .A(n14693), .B(n14692), .ZN(
        P1_U3007) );
  INV_X1 U18006 ( .A(n15795), .ZN(n14699) );
  NOR2_X1 U18007 ( .A1(n14695), .A2(n11606), .ZN(n14698) );
  NAND2_X1 U18008 ( .A1(n15899), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14696) );
  OAI21_X1 U18009 ( .B1(n15603), .B2(n20137), .A(n14696), .ZN(n14697) );
  AOI211_X1 U18010 ( .C1(n14699), .C2(n11606), .A(n14698), .B(n14697), .ZN(
        n14700) );
  OAI21_X1 U18011 ( .B1(n14701), .B2(n20138), .A(n14700), .ZN(P1_U3008) );
  NAND2_X1 U18012 ( .A1(n15809), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14703) );
  OAI211_X1 U18013 ( .C1(n20137), .C2(n15628), .A(n14703), .B(n14702), .ZN(
        n14704) );
  AOI21_X1 U18014 ( .B1(n15808), .B2(n14581), .A(n14704), .ZN(n14705) );
  OAI21_X1 U18015 ( .B1(n14706), .B2(n20138), .A(n14705), .ZN(P1_U3010) );
  INV_X1 U18016 ( .A(n15641), .ZN(n14710) );
  NAND2_X1 U18017 ( .A1(n15899), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14707) );
  OAI221_X1 U18018 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15804), 
        .C1(n14708), .C2(n15573), .A(n14707), .ZN(n14709) );
  AOI21_X1 U18019 ( .B1(n14710), .B2(n15932), .A(n14709), .ZN(n14711) );
  OAI21_X1 U18020 ( .B1(n14712), .B2(n20138), .A(n14711), .ZN(P1_U3012) );
  XNOR2_X1 U18021 ( .A(n20220), .B(P1_STATEBS16_REG_SCAN_IN), .ZN(n14713) );
  OAI22_X1 U18022 ( .A1(n14713), .A2(n20651), .B1(n13514), .B2(n14719), .ZN(
        n14714) );
  MUX2_X1 U18023 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14714), .S(
        n20147), .Z(P1_U3477) );
  NAND2_X1 U18024 ( .A1(n20220), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14715) );
  NAND2_X1 U18025 ( .A1(n14715), .A2(n20658), .ZN(n20650) );
  MUX2_X1 U18026 ( .A(n20650), .B(n14717), .S(n14716), .Z(n14718) );
  OAI21_X1 U18027 ( .B1(n14719), .B2(n13310), .A(n14718), .ZN(n14720) );
  MUX2_X1 U18028 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14720), .S(
        n20147), .Z(P1_U3476) );
  OR2_X1 U18029 ( .A1(n13514), .A2(n14721), .ZN(n14728) );
  INV_X1 U18030 ( .A(n13342), .ZN(n14722) );
  NAND3_X1 U18031 ( .A1(n14724), .A2(n14723), .A3(n14722), .ZN(n14725) );
  AND2_X1 U18032 ( .A1(n14726), .A2(n14725), .ZN(n14727) );
  NAND2_X1 U18033 ( .A1(n14728), .A2(n14727), .ZN(n15504) );
  INV_X1 U18034 ( .A(n15504), .ZN(n14734) );
  INV_X1 U18035 ( .A(n15942), .ZN(n20788) );
  AOI22_X1 U18036 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n14730), .B2(n14729), .ZN(
        n14736) );
  INV_X1 U18037 ( .A(n14736), .ZN(n14732) );
  NOR2_X1 U18038 ( .A1(n20717), .A2(n15823), .ZN(n14737) );
  NOR3_X1 U18039 ( .A1(n13342), .A2(n13311), .A3(n20786), .ZN(n14731) );
  AOI21_X1 U18040 ( .B1(n14732), .B2(n14737), .A(n14731), .ZN(n14733) );
  OAI21_X1 U18041 ( .B1(n14734), .B2(n20788), .A(n14733), .ZN(n14735) );
  MUX2_X1 U18042 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14735), .S(
        n20790), .Z(P1_U3473) );
  AOI22_X1 U18043 ( .A1(n14738), .A2(n15551), .B1(n14737), .B2(n14736), .ZN(
        n14739) );
  OAI21_X1 U18044 ( .B1(n14740), .B2(n20788), .A(n14739), .ZN(n14741) );
  MUX2_X1 U18045 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14741), .S(
        n20790), .Z(P1_U3472) );
  INV_X1 U18046 ( .A(n14745), .ZN(n14810) );
  NAND2_X1 U18047 ( .A1(n14747), .A2(n14746), .ZN(n14809) );
  NAND3_X1 U18048 ( .A1(n14810), .A2(n19107), .A3(n14809), .ZN(n14749) );
  NAND2_X1 U18049 ( .A1(n19116), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14748) );
  OAI211_X1 U18050 ( .C1(n19116), .C2(n15989), .A(n14749), .B(n14748), .ZN(
        P2_U2858) );
  NAND2_X1 U18051 ( .A1(n14751), .A2(n14750), .ZN(n14753) );
  XNOR2_X1 U18052 ( .A(n14753), .B(n14752), .ZN(n14824) );
  NOR2_X1 U18053 ( .A1(n16004), .A2(n19116), .ZN(n14754) );
  AOI21_X1 U18054 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19116), .A(n14754), .ZN(
        n14755) );
  OAI21_X1 U18055 ( .B1(n14824), .B2(n19117), .A(n14755), .ZN(P2_U2859) );
  AOI21_X1 U18056 ( .B1(n14758), .B2(n14757), .A(n14756), .ZN(n14759) );
  INV_X1 U18057 ( .A(n14759), .ZN(n14831) );
  NAND2_X1 U18058 ( .A1(n14767), .A2(n14760), .ZN(n14761) );
  NAND2_X1 U18059 ( .A1(n14762), .A2(n14761), .ZN(n16014) );
  NOR2_X1 U18060 ( .A1(n16014), .A2(n19116), .ZN(n14763) );
  AOI21_X1 U18061 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n19116), .A(n14763), .ZN(
        n14764) );
  OAI21_X1 U18062 ( .B1(n14831), .B2(n19117), .A(n14764), .ZN(P2_U2860) );
  NAND2_X1 U18063 ( .A1(n14776), .A2(n14765), .ZN(n14766) );
  NAND2_X1 U18064 ( .A1(n14767), .A2(n14766), .ZN(n16021) );
  AOI21_X1 U18065 ( .B1(n14768), .B2(n14770), .A(n14769), .ZN(n14832) );
  NAND2_X1 U18066 ( .A1(n14832), .A2(n19107), .ZN(n14772) );
  NAND2_X1 U18067 ( .A1(n19116), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14771) );
  OAI211_X1 U18068 ( .C1(n16021), .C2(n19116), .A(n14772), .B(n14771), .ZN(
        P2_U2861) );
  OAI21_X1 U18069 ( .B1(n14775), .B2(n14774), .A(n14773), .ZN(n14849) );
  OAI21_X1 U18070 ( .B1(n14785), .B2(n14777), .A(n14776), .ZN(n15096) );
  MUX2_X1 U18071 ( .A(n14778), .B(n15096), .S(n19121), .Z(n14779) );
  OAI21_X1 U18072 ( .B1(n14849), .B2(n19117), .A(n14779), .ZN(P2_U2862) );
  AOI21_X1 U18073 ( .B1(n14781), .B2(n14780), .A(n9893), .ZN(n14782) );
  XOR2_X1 U18074 ( .A(n14783), .B(n14782), .Z(n14856) );
  AND2_X1 U18075 ( .A1(n14949), .A2(n14784), .ZN(n14786) );
  OR2_X1 U18076 ( .A1(n14786), .A2(n14785), .ZN(n16038) );
  NOR2_X1 U18077 ( .A1(n16038), .A2(n19116), .ZN(n14787) );
  AOI21_X1 U18078 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n19116), .A(n14787), .ZN(
        n14788) );
  OAI21_X1 U18079 ( .B1(n14856), .B2(n19117), .A(n14788), .ZN(P2_U2863) );
  OAI21_X1 U18080 ( .B1(n16068), .B2(n14790), .A(n14789), .ZN(n14880) );
  NAND2_X1 U18081 ( .A1(n14791), .A2(n14792), .ZN(n14794) );
  INV_X1 U18082 ( .A(n14793), .ZN(n15149) );
  INV_X1 U18083 ( .A(n18847), .ZN(n15594) );
  MUX2_X1 U18084 ( .A(n14795), .B(n15594), .S(n19121), .Z(n14796) );
  OAI21_X1 U18085 ( .B1(n14880), .B2(n19117), .A(n14796), .ZN(P2_U2866) );
  OAI21_X1 U18086 ( .B1(n9917), .B2(n14798), .A(n14797), .ZN(n14892) );
  AND2_X1 U18087 ( .A1(n15008), .A2(n14799), .ZN(n14800) );
  OR2_X1 U18088 ( .A1(n14983), .A2(n14800), .ZN(n18866) );
  NOR2_X1 U18089 ( .A1(n18866), .A2(n19116), .ZN(n14801) );
  AOI21_X1 U18090 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19116), .A(n14801), .ZN(
        n14802) );
  OAI21_X1 U18091 ( .B1(n14892), .B2(n19117), .A(n14802), .ZN(P2_U2868) );
  INV_X1 U18092 ( .A(n14804), .ZN(n14805) );
  AOI21_X1 U18093 ( .B1(n10110), .B2(n14805), .A(n9887), .ZN(n18896) );
  INV_X1 U18094 ( .A(n18896), .ZN(n15213) );
  NOR2_X1 U18095 ( .A1(n15213), .A2(n19116), .ZN(n14806) );
  AOI21_X1 U18096 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n19116), .A(n14806), .ZN(
        n14807) );
  OAI21_X1 U18097 ( .B1(n14808), .B2(n19117), .A(n14807), .ZN(P2_U2870) );
  NAND3_X1 U18098 ( .A1(n14810), .A2(n19176), .A3(n14809), .ZN(n14819) );
  OR2_X1 U18099 ( .A1(n14812), .A2(n14811), .ZN(n14813) );
  NAND2_X1 U18100 ( .A1(n14814), .A2(n14813), .ZN(n15993) );
  INV_X1 U18101 ( .A(n15993), .ZN(n15063) );
  OAI22_X1 U18102 ( .A1(n14884), .A2(n19142), .B1(n19162), .B2(n14815), .ZN(
        n14816) );
  AOI21_X1 U18103 ( .B1(n19187), .B2(n15063), .A(n14816), .ZN(n14818) );
  AOI22_X1 U18104 ( .A1(n19127), .A2(BUF1_REG_29__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14817) );
  NAND3_X1 U18105 ( .A1(n14819), .A2(n14818), .A3(n14817), .ZN(P2_U2890) );
  INV_X1 U18106 ( .A(n19145), .ZN(n14820) );
  OAI22_X1 U18107 ( .A1(n14884), .A2(n14820), .B1(n19162), .B2(n12989), .ZN(
        n14821) );
  AOI21_X1 U18108 ( .B1(n19187), .B2(n16002), .A(n14821), .ZN(n14823) );
  AOI22_X1 U18109 ( .A1(n19127), .A2(BUF1_REG_28__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n14822) );
  OAI211_X1 U18110 ( .C1(n14824), .C2(n19191), .A(n14823), .B(n14822), .ZN(
        P2_U2891) );
  NAND2_X1 U18111 ( .A1(n9896), .A2(n14825), .ZN(n14826) );
  NAND2_X1 U18112 ( .A1(n9835), .A2(n14826), .ZN(n16008) );
  INV_X1 U18113 ( .A(n16008), .ZN(n15077) );
  OAI22_X1 U18114 ( .A1(n14884), .A2(n19148), .B1(n19162), .B2(n14827), .ZN(
        n14828) );
  AOI21_X1 U18115 ( .B1(n19187), .B2(n15077), .A(n14828), .ZN(n14830) );
  AOI22_X1 U18116 ( .A1(n19127), .A2(BUF1_REG_27__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n14829) );
  OAI211_X1 U18117 ( .C1(n14831), .C2(n19191), .A(n14830), .B(n14829), .ZN(
        P2_U2892) );
  NAND2_X1 U18118 ( .A1(n14832), .A2(n19176), .ZN(n14839) );
  INV_X1 U18119 ( .A(n14884), .ZN(n19125) );
  AOI22_X1 U18120 ( .A1(n19125), .A2(n19150), .B1(P2_EAX_REG_26__SCAN_IN), 
        .B2(n19186), .ZN(n14838) );
  AOI22_X1 U18121 ( .A1(n19127), .A2(BUF1_REG_26__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n14837) );
  OAI21_X1 U18122 ( .B1(n14833), .B2(n14834), .A(n9896), .ZN(n14835) );
  INV_X1 U18123 ( .A(n14835), .ZN(n16024) );
  NAND2_X1 U18124 ( .A1(n19187), .A2(n16024), .ZN(n14836) );
  NAND4_X1 U18125 ( .A1(n14839), .A2(n14838), .A3(n14837), .A4(n14836), .ZN(
        P2_U2893) );
  NOR2_X1 U18126 ( .A1(n14850), .A2(n14840), .ZN(n14841) );
  OR2_X1 U18127 ( .A1(n14833), .A2(n14841), .ZN(n16033) );
  INV_X1 U18128 ( .A(n16033), .ZN(n14847) );
  OAI22_X1 U18129 ( .A1(n14884), .A2(n19153), .B1(n19162), .B2(n14842), .ZN(
        n14846) );
  INV_X1 U18130 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n14844) );
  INV_X1 U18131 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n14843) );
  OAI22_X1 U18132 ( .A1(n14888), .A2(n14844), .B1(n14886), .B2(n14843), .ZN(
        n14845) );
  AOI211_X1 U18133 ( .C1(n19187), .C2(n14847), .A(n14846), .B(n14845), .ZN(
        n14848) );
  OAI21_X1 U18134 ( .B1(n14849), .B2(n19191), .A(n14848), .ZN(P2_U2894) );
  AOI21_X1 U18135 ( .B1(n14851), .B2(n14864), .A(n14850), .ZN(n16039) );
  INV_X1 U18136 ( .A(n19156), .ZN(n14852) );
  OAI22_X1 U18137 ( .A1(n14884), .A2(n14852), .B1(n19162), .B2(n12986), .ZN(
        n14853) );
  AOI21_X1 U18138 ( .B1(n19187), .B2(n16039), .A(n14853), .ZN(n14855) );
  AOI22_X1 U18139 ( .A1(n19127), .A2(BUF1_REG_24__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n14854) );
  OAI211_X1 U18140 ( .C1(n14856), .C2(n19191), .A(n14855), .B(n14854), .ZN(
        P2_U2895) );
  NOR2_X1 U18141 ( .A1(n14858), .A2(n14857), .ZN(n14860) );
  NOR2_X1 U18142 ( .A1(n14860), .A2(n14859), .ZN(n16062) );
  INV_X1 U18143 ( .A(n16062), .ZN(n14871) );
  NAND2_X1 U18144 ( .A1(n14861), .A2(n14862), .ZN(n14863) );
  NAND2_X1 U18145 ( .A1(n14864), .A2(n14863), .ZN(n16055) );
  INV_X1 U18146 ( .A(n16055), .ZN(n14869) );
  OAI22_X1 U18147 ( .A1(n14884), .A2(n19159), .B1(n19162), .B2(n14865), .ZN(
        n14868) );
  INV_X1 U18148 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14866) );
  OAI22_X1 U18149 ( .A1(n14888), .A2(n16385), .B1(n14886), .B2(n14866), .ZN(
        n14867) );
  AOI211_X1 U18150 ( .C1(n19187), .C2(n14869), .A(n14868), .B(n14867), .ZN(
        n14870) );
  OAI21_X1 U18151 ( .B1(n14871), .B2(n19191), .A(n14870), .ZN(P2_U2896) );
  OR2_X1 U18152 ( .A1(n10237), .A2(n14872), .ZN(n14873) );
  AND2_X1 U18153 ( .A1(n15145), .A2(n14873), .ZN(n18846) );
  OAI22_X1 U18154 ( .A1(n14884), .A2(n19288), .B1(n19162), .B2(n14874), .ZN(
        n14878) );
  INV_X1 U18155 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14876) );
  INV_X1 U18156 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14875) );
  OAI22_X1 U18157 ( .A1(n14888), .A2(n14876), .B1(n14886), .B2(n14875), .ZN(
        n14877) );
  AOI211_X1 U18158 ( .C1(n19187), .C2(n18846), .A(n14878), .B(n14877), .ZN(
        n14879) );
  OAI21_X1 U18159 ( .B1(n14880), .B2(n19191), .A(n14879), .ZN(P2_U2898) );
  NAND2_X1 U18160 ( .A1(n15186), .A2(n14881), .ZN(n14882) );
  NAND2_X1 U18161 ( .A1(n9891), .A2(n14882), .ZN(n18877) );
  INV_X1 U18162 ( .A(n18877), .ZN(n15171) );
  OAI22_X1 U18163 ( .A1(n14884), .A2(n19279), .B1(n19162), .B2(n14883), .ZN(
        n14890) );
  INV_X1 U18164 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14887) );
  INV_X1 U18165 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14885) );
  OAI22_X1 U18166 ( .A1(n14888), .A2(n14887), .B1(n14886), .B2(n14885), .ZN(
        n14889) );
  AOI211_X1 U18167 ( .C1(n19187), .C2(n15171), .A(n14890), .B(n14889), .ZN(
        n14891) );
  OAI21_X1 U18168 ( .B1(n14892), .B2(n19191), .A(n14891), .ZN(P2_U2900) );
  XNOR2_X1 U18169 ( .A(n9923), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15960) );
  NOR2_X1 U18170 ( .A1(n15960), .A2(n19247), .ZN(n14896) );
  NAND2_X1 U18171 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14893) );
  OAI211_X1 U18172 ( .C1(n15983), .C2(n15339), .A(n14894), .B(n14893), .ZN(
        n14895) );
  AOI211_X1 U18173 ( .C1(n14897), .C2(n19242), .A(n14896), .B(n14895), .ZN(
        n14898) );
  OAI21_X1 U18174 ( .B1(n14899), .B2(n16173), .A(n14898), .ZN(P2_U2984) );
  NOR2_X1 U18175 ( .A1(n14901), .A2(n14900), .ZN(n14904) );
  INV_X1 U18176 ( .A(n14902), .ZN(n14903) );
  XOR2_X1 U18177 ( .A(n14904), .B(n14903), .Z(n15072) );
  AOI21_X1 U18178 ( .B1(n14906), .B2(n14905), .A(n9923), .ZN(n15984) );
  NOR2_X1 U18179 ( .A1(n15989), .A2(n15339), .ZN(n14908) );
  NAND2_X1 U18180 ( .A1(n12763), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15062) );
  OAI21_X1 U18181 ( .B1(n16179), .B2(n14906), .A(n15062), .ZN(n14907) );
  AOI211_X1 U18182 ( .C1(n15984), .C2(n16170), .A(n14908), .B(n14907), .ZN(
        n14912) );
  AOI21_X1 U18183 ( .B1(n14910), .B2(n14909), .A(n13962), .ZN(n15069) );
  NAND2_X1 U18184 ( .A1(n15069), .A2(n19242), .ZN(n14911) );
  OAI211_X1 U18185 ( .C1(n15072), .C2(n16173), .A(n14912), .B(n14911), .ZN(
        P2_U2985) );
  INV_X1 U18186 ( .A(n14914), .ZN(n14915) );
  OAI21_X1 U18187 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n10219), .A(
        n14915), .ZN(n15085) );
  NAND3_X1 U18188 ( .A1(n14916), .A2(n19240), .A3(n15073), .ZN(n14923) );
  NOR2_X1 U18189 ( .A1(n14928), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14918) );
  NOR2_X1 U18190 ( .A1(n16232), .A2(n19894), .ZN(n15076) );
  AOI21_X1 U18191 ( .B1(n19239), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n15076), .ZN(n14920) );
  OAI21_X1 U18192 ( .B1(n16014), .B2(n15339), .A(n14920), .ZN(n14921) );
  AOI21_X1 U18193 ( .B1(n9914), .B2(n16170), .A(n14921), .ZN(n14922) );
  OAI211_X1 U18194 ( .C1(n16172), .C2(n15085), .A(n14923), .B(n14922), .ZN(
        P2_U2987) );
  INV_X1 U18195 ( .A(n14933), .ZN(n14924) );
  OAI21_X1 U18196 ( .B1(n9856), .B2(n14924), .A(n14934), .ZN(n14925) );
  XOR2_X1 U18197 ( .A(n14926), .B(n14925), .Z(n15095) );
  NAND2_X1 U18198 ( .A1(n15112), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15105) );
  AOI21_X1 U18199 ( .B1(n15091), .B2(n15105), .A(n10219), .ZN(n15093) );
  NOR2_X1 U18200 ( .A1(n14936), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14927) );
  OR2_X1 U18201 ( .A1(n14928), .A2(n14927), .ZN(n15961) );
  NOR2_X1 U18202 ( .A1(n16232), .A2(n19890), .ZN(n15088) );
  NOR2_X1 U18203 ( .A1(n16021), .A2(n15339), .ZN(n14929) );
  AOI211_X1 U18204 ( .C1(n19239), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15088), .B(n14929), .ZN(n14930) );
  OAI21_X1 U18205 ( .B1(n15961), .B2(n19247), .A(n14930), .ZN(n14931) );
  AOI21_X1 U18206 ( .B1(n15093), .B2(n19242), .A(n14931), .ZN(n14932) );
  OAI21_X1 U18207 ( .B1(n15095), .B2(n16173), .A(n14932), .ZN(P2_U2988) );
  NAND2_X1 U18208 ( .A1(n14934), .A2(n14933), .ZN(n14935) );
  XOR2_X1 U18209 ( .A(n14935), .B(n9856), .Z(n15108) );
  AOI21_X1 U18210 ( .B1(n15962), .B2(n16028), .A(n14936), .ZN(n16027) );
  NAND2_X1 U18211 ( .A1(n19016), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15097) );
  NAND2_X1 U18212 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14937) );
  OAI211_X1 U18213 ( .C1(n15096), .C2(n15339), .A(n15097), .B(n14937), .ZN(
        n14938) );
  AOI21_X1 U18214 ( .B1(n16027), .B2(n16170), .A(n14938), .ZN(n14941) );
  NAND2_X1 U18215 ( .A1(n14939), .A2(n15102), .ZN(n15104) );
  NAND3_X1 U18216 ( .A1(n15105), .A2(n19242), .A3(n15104), .ZN(n14940) );
  OAI211_X1 U18217 ( .C1(n15108), .C2(n16173), .A(n14941), .B(n14940), .ZN(
        P2_U2989) );
  OAI21_X1 U18218 ( .B1(n9838), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9869), .ZN(n15132) );
  NAND2_X1 U18219 ( .A1(n14944), .A2(n14943), .ZN(n15122) );
  NAND3_X1 U18220 ( .A1(n9975), .A2(n19240), .A3(n15122), .ZN(n14955) );
  INV_X1 U18221 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14945) );
  NAND2_X1 U18222 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n9885), .ZN(
        n15481) );
  AOI21_X1 U18223 ( .B1(n14945), .B2(n15481), .A(n15963), .ZN(n16051) );
  OAI22_X1 U18224 ( .A1(n16179), .A2(n14945), .B1(n19885), .B2(n16232), .ZN(
        n14953) );
  INV_X1 U18225 ( .A(n15148), .ZN(n14948) );
  INV_X1 U18226 ( .A(n14946), .ZN(n14947) );
  NAND2_X1 U18227 ( .A1(n14948), .A2(n14947), .ZN(n14950) );
  AND2_X1 U18228 ( .A1(n14950), .A2(n14949), .ZN(n16061) );
  INV_X1 U18229 ( .A(n16061), .ZN(n14951) );
  NOR2_X1 U18230 ( .A1(n14951), .A2(n15339), .ZN(n14952) );
  AOI211_X1 U18231 ( .C1(n16051), .C2(n16170), .A(n14953), .B(n14952), .ZN(
        n14954) );
  OAI211_X1 U18232 ( .C1(n15132), .C2(n16172), .A(n14955), .B(n14954), .ZN(
        P2_U2991) );
  INV_X1 U18233 ( .A(n15233), .ZN(n14956) );
  NAND2_X1 U18234 ( .A1(n16113), .A2(n16111), .ZN(n15042) );
  INV_X1 U18235 ( .A(n15041), .ZN(n14957) );
  INV_X1 U18236 ( .A(n14960), .ZN(n14961) );
  AOI21_X1 U18237 ( .B1(n14977), .B2(n14962), .A(n14976), .ZN(n14966) );
  NOR2_X1 U18238 ( .A1(n14964), .A2(n14963), .ZN(n14965) );
  XNOR2_X1 U18239 ( .A(n14966), .B(n14965), .ZN(n15599) );
  AND2_X1 U18240 ( .A1(n14980), .A2(n15588), .ZN(n14968) );
  OR2_X1 U18241 ( .A1(n14967), .A2(n14968), .ZN(n15595) );
  AOI21_X1 U18242 ( .B1(n14969), .B2(n14986), .A(n9885), .ZN(n18849) );
  OAI22_X1 U18243 ( .A1(n16179), .A2(n14969), .B1(n19882), .B2(n16232), .ZN(
        n14970) );
  AOI21_X1 U18244 ( .B1(n18849), .B2(n16170), .A(n14970), .ZN(n14972) );
  NAND2_X1 U18245 ( .A1(n18847), .A2(n19250), .ZN(n14971) );
  OAI211_X1 U18246 ( .C1(n15595), .C2(n16172), .A(n14972), .B(n14971), .ZN(
        n14973) );
  INV_X1 U18247 ( .A(n14973), .ZN(n14974) );
  OAI21_X1 U18248 ( .B1(n15599), .B2(n16173), .A(n14974), .ZN(P2_U2993) );
  NOR2_X1 U18249 ( .A1(n14976), .A2(n14975), .ZN(n14978) );
  XOR2_X1 U18250 ( .A(n14978), .B(n14977), .Z(n15168) );
  OAI21_X1 U18251 ( .B1(n14979), .B2(n15177), .A(n15164), .ZN(n14981) );
  AND2_X1 U18252 ( .A1(n14981), .A2(n14980), .ZN(n15166) );
  OR2_X1 U18253 ( .A1(n14983), .A2(n14982), .ZN(n14984) );
  NAND2_X1 U18254 ( .A1(n14791), .A2(n14984), .ZN(n18865) );
  NOR2_X1 U18255 ( .A1(n16232), .A2(n19880), .ZN(n15160) );
  OAI21_X1 U18256 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n14985), .A(
        n14986), .ZN(n15495) );
  NOR2_X1 U18257 ( .A1(n15495), .A2(n19247), .ZN(n14987) );
  AOI211_X1 U18258 ( .C1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n19239), .A(
        n15160), .B(n14987), .ZN(n14988) );
  OAI21_X1 U18259 ( .B1(n18865), .B2(n15339), .A(n14988), .ZN(n14989) );
  AOI21_X1 U18260 ( .B1(n15166), .B2(n19242), .A(n14989), .ZN(n14990) );
  OAI21_X1 U18261 ( .B1(n15168), .B2(n16173), .A(n14990), .ZN(P2_U2994) );
  INV_X1 U18262 ( .A(n15001), .ZN(n14991) );
  OAI21_X1 U18263 ( .B1(n15003), .B2(n14991), .A(n15002), .ZN(n14995) );
  NAND2_X1 U18264 ( .A1(n14993), .A2(n14992), .ZN(n14994) );
  XNOR2_X1 U18265 ( .A(n14995), .B(n14994), .ZN(n15181) );
  XNOR2_X1 U18266 ( .A(n14979), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15179) );
  AOI21_X1 U18267 ( .B1(n14996), .B2(n15012), .A(n14985), .ZN(n18869) );
  NAND2_X1 U18268 ( .A1(n19016), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15169) );
  OAI21_X1 U18269 ( .B1(n16179), .B2(n14996), .A(n15169), .ZN(n14997) );
  AOI21_X1 U18270 ( .B1(n18869), .B2(n16170), .A(n14997), .ZN(n14998) );
  OAI21_X1 U18271 ( .B1(n18866), .B2(n15339), .A(n14998), .ZN(n14999) );
  AOI21_X1 U18272 ( .B1(n15179), .B2(n19242), .A(n14999), .ZN(n15000) );
  OAI21_X1 U18273 ( .B1(n15181), .B2(n16173), .A(n15000), .ZN(P2_U2995) );
  NAND2_X1 U18274 ( .A1(n15002), .A2(n15001), .ZN(n15004) );
  XOR2_X1 U18275 ( .A(n15004), .B(n15003), .Z(n15201) );
  INV_X1 U18276 ( .A(n15005), .ZN(n15210) );
  NOR2_X2 U18277 ( .A1(n15035), .A2(n15210), .ZN(n15203) );
  AOI21_X1 U18278 ( .B1(n15203), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15006) );
  NOR2_X1 U18279 ( .A1(n15006), .A2(n12807), .ZN(n15199) );
  INV_X1 U18280 ( .A(n15007), .ZN(n15009) );
  OAI21_X1 U18281 ( .B1(n9887), .B2(n15009), .A(n15008), .ZN(n18888) );
  NOR2_X1 U18282 ( .A1(n16232), .A2(n15010), .ZN(n15190) );
  OR2_X1 U18283 ( .A1(n15022), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15011) );
  NAND2_X1 U18284 ( .A1(n15012), .A2(n15011), .ZN(n18882) );
  NOR2_X1 U18285 ( .A1(n18882), .A2(n19247), .ZN(n15013) );
  AOI211_X1 U18286 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19239), .A(
        n15190), .B(n15013), .ZN(n15014) );
  OAI21_X1 U18287 ( .B1(n18888), .B2(n15339), .A(n15014), .ZN(n15015) );
  AOI21_X1 U18288 ( .B1(n15199), .B2(n19242), .A(n15015), .ZN(n15016) );
  OAI21_X1 U18289 ( .B1(n15201), .B2(n16173), .A(n15016), .ZN(P2_U2996) );
  NAND2_X1 U18290 ( .A1(n15018), .A2(n15017), .ZN(n15021) );
  NAND2_X1 U18291 ( .A1(n15026), .A2(n15019), .ZN(n15020) );
  XOR2_X1 U18292 ( .A(n15021), .B(n15020), .Z(n15218) );
  INV_X1 U18293 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15024) );
  NAND2_X1 U18294 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n9884), .ZN(
        n15029) );
  AOI21_X1 U18295 ( .B1(n15024), .B2(n15029), .A(n15022), .ZN(n18891) );
  NAND2_X1 U18296 ( .A1(n16170), .A2(n18891), .ZN(n15023) );
  NAND2_X1 U18297 ( .A1(n12763), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15212) );
  OAI211_X1 U18298 ( .C1(n15024), .C2(n16179), .A(n15023), .B(n15212), .ZN(
        n15025) );
  OAI21_X1 U18299 ( .B1(n15028), .B2(n15027), .A(n15026), .ZN(n15219) );
  OAI21_X1 U18300 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n9884), .A(
        n15029), .ZN(n18904) );
  OAI22_X1 U18301 ( .A1(n19873), .A2(n16232), .B1(n19247), .B2(n18904), .ZN(
        n15034) );
  AND2_X1 U18302 ( .A1(n15031), .A2(n15030), .ZN(n15032) );
  OR2_X1 U18303 ( .A1(n15032), .A2(n14804), .ZN(n19091) );
  NOR2_X1 U18304 ( .A1(n19091), .A2(n15339), .ZN(n15033) );
  AOI211_X1 U18305 ( .C1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19239), .A(
        n15034), .B(n15033), .ZN(n15039) );
  INV_X1 U18306 ( .A(n15203), .ZN(n15037) );
  OAI21_X1 U18307 ( .B1(n15035), .B2(n16187), .A(n15230), .ZN(n15036) );
  NAND3_X1 U18308 ( .A1(n15037), .A2(n19242), .A3(n15036), .ZN(n15038) );
  OAI211_X1 U18309 ( .C1(n15219), .C2(n16173), .A(n15039), .B(n15038), .ZN(
        P2_U2998) );
  XNOR2_X1 U18310 ( .A(n15035), .B(n16187), .ZN(n16190) );
  NAND2_X1 U18311 ( .A1(n15041), .A2(n15040), .ZN(n15044) );
  NAND2_X1 U18312 ( .A1(n15042), .A2(n16110), .ZN(n15043) );
  XOR2_X1 U18313 ( .A(n15044), .B(n15043), .Z(n16194) );
  INV_X1 U18314 ( .A(n16194), .ZN(n15049) );
  AOI21_X1 U18315 ( .B1(n15045), .B2(n15493), .A(n9884), .ZN(n18914) );
  AOI22_X1 U18316 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n16170), .B2(n18914), .ZN(n15046) );
  NAND2_X1 U18317 ( .A1(n19016), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n16185) );
  OAI211_X1 U18318 ( .C1(n15047), .C2(n15339), .A(n15046), .B(n16185), .ZN(
        n15048) );
  AOI21_X1 U18319 ( .B1(n15049), .B2(n19240), .A(n15048), .ZN(n15050) );
  OAI21_X1 U18320 ( .B1(n16172), .B2(n16190), .A(n15050), .ZN(P2_U2999) );
  NAND2_X1 U18321 ( .A1(n15051), .A2(n15052), .ZN(n16154) );
  INV_X1 U18322 ( .A(n16153), .ZN(n15054) );
  AND2_X1 U18323 ( .A1(n15052), .A2(n16153), .ZN(n15053) );
  OAI22_X1 U18324 ( .A1(n16154), .A2(n15054), .B1(n15053), .B2(n15051), .ZN(
        n15282) );
  OR2_X1 U18325 ( .A1(n15055), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15270) );
  NAND3_X1 U18326 ( .A1(n15270), .A2(n15269), .A3(n19242), .ZN(n15061) );
  AOI21_X1 U18327 ( .B1(n18994), .B2(n15488), .A(n15056), .ZN(n18998) );
  NOR2_X1 U18328 ( .A1(n15057), .A2(n15339), .ZN(n15059) );
  OAI22_X1 U18329 ( .A1(n16179), .A2(n18994), .B1(n19862), .B2(n16232), .ZN(
        n15058) );
  AOI211_X1 U18330 ( .C1(n16170), .C2(n18998), .A(n15059), .B(n15058), .ZN(
        n15060) );
  OAI211_X1 U18331 ( .C1(n16173), .C2(n15282), .A(n15061), .B(n15060), .ZN(
        P2_U3007) );
  INV_X1 U18332 ( .A(n15064), .ZN(n15065) );
  NOR3_X1 U18333 ( .A1(n15074), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15065), .ZN(n15066) );
  NAND2_X1 U18334 ( .A1(n15069), .A2(n19262), .ZN(n15070) );
  OAI211_X1 U18335 ( .C1(n15072), .C2(n16246), .A(n15071), .B(n15070), .ZN(
        P2_U3017) );
  NAND3_X1 U18336 ( .A1(n14916), .A2(n19263), .A3(n15073), .ZN(n15084) );
  INV_X1 U18337 ( .A(n15074), .ZN(n15082) );
  NOR2_X1 U18338 ( .A1(n16014), .A2(n16253), .ZN(n15075) );
  AOI211_X1 U18339 ( .C1(n15077), .C2(n19257), .A(n15076), .B(n15075), .ZN(
        n15078) );
  OAI21_X1 U18340 ( .B1(n15079), .B2(n15081), .A(n15078), .ZN(n15080) );
  AOI21_X1 U18341 ( .B1(n15082), .B2(n15081), .A(n15080), .ZN(n15083) );
  OAI211_X1 U18342 ( .C1(n15085), .C2(n16264), .A(n15084), .B(n15083), .ZN(
        P2_U3019) );
  OAI211_X1 U18343 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15103), .B(n15086), .ZN(
        n15090) );
  NOR2_X1 U18344 ( .A1(n16021), .A2(n16253), .ZN(n15087) );
  AOI211_X1 U18345 ( .C1(n19257), .C2(n16024), .A(n15088), .B(n15087), .ZN(
        n15089) );
  OAI211_X1 U18346 ( .C1(n15100), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        n15092) );
  AOI21_X1 U18347 ( .B1(n15093), .B2(n19262), .A(n15092), .ZN(n15094) );
  OAI21_X1 U18348 ( .B1(n15095), .B2(n16246), .A(n15094), .ZN(P2_U3020) );
  INV_X1 U18349 ( .A(n15096), .ZN(n16036) );
  OAI21_X1 U18350 ( .B1(n16215), .B2(n16033), .A(n15097), .ZN(n15098) );
  AOI21_X1 U18351 ( .B1(n19255), .B2(n16036), .A(n15098), .ZN(n15099) );
  OAI21_X1 U18352 ( .B1(n15100), .B2(n15102), .A(n15099), .ZN(n15101) );
  AOI21_X1 U18353 ( .B1(n15103), .B2(n15102), .A(n15101), .ZN(n15107) );
  NAND3_X1 U18354 ( .A1(n15105), .A2(n19262), .A3(n15104), .ZN(n15106) );
  OAI211_X1 U18355 ( .C1(n15108), .C2(n16246), .A(n15107), .B(n15106), .ZN(
        P2_U3021) );
  NOR2_X1 U18356 ( .A1(n15109), .A2(n9895), .ZN(n15110) );
  XNOR2_X1 U18357 ( .A(n15111), .B(n15110), .ZN(n16089) );
  INV_X1 U18358 ( .A(n16089), .ZN(n15121) );
  AOI21_X1 U18359 ( .B1(n15115), .B2(n9869), .A(n15112), .ZN(n16087) );
  AOI21_X1 U18360 ( .B1(n15115), .B2(n15114), .A(n15113), .ZN(n15117) );
  NOR2_X1 U18361 ( .A1(n16232), .A2(n12755), .ZN(n15116) );
  AOI211_X1 U18362 ( .C1(n19257), .C2(n16039), .A(n15117), .B(n15116), .ZN(
        n15118) );
  OAI21_X1 U18363 ( .B1(n16253), .B2(n16038), .A(n15118), .ZN(n15119) );
  AOI21_X1 U18364 ( .B1(n16087), .B2(n19262), .A(n15119), .ZN(n15120) );
  OAI21_X1 U18365 ( .B1(n15121), .B2(n16246), .A(n15120), .ZN(P2_U3022) );
  NAND3_X1 U18366 ( .A1(n9975), .A2(n19263), .A3(n15122), .ZN(n15131) );
  AOI21_X1 U18367 ( .B1(n15127), .B2(n15141), .A(n15123), .ZN(n15129) );
  NOR2_X1 U18368 ( .A1(n19885), .A2(n16232), .ZN(n15125) );
  NOR2_X1 U18369 ( .A1(n16215), .A2(n16055), .ZN(n15124) );
  AOI211_X1 U18370 ( .C1(n16061), .C2(n19255), .A(n15125), .B(n15124), .ZN(
        n15126) );
  OAI21_X1 U18371 ( .B1(n15140), .B2(n15127), .A(n15126), .ZN(n15128) );
  AOI21_X1 U18372 ( .B1(n15138), .B2(n15129), .A(n15128), .ZN(n15130) );
  OAI211_X1 U18373 ( .C1(n15132), .C2(n16264), .A(n15131), .B(n15130), .ZN(
        P2_U3023) );
  INV_X1 U18374 ( .A(n15133), .ZN(n15134) );
  NOR2_X1 U18375 ( .A1(n15135), .A2(n15134), .ZN(n15136) );
  XNOR2_X1 U18376 ( .A(n15137), .B(n15136), .ZN(n16094) );
  NOR2_X1 U18377 ( .A1(n14967), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16093) );
  NOR3_X1 U18378 ( .A1(n16093), .A2(n9838), .A3(n16264), .ZN(n15155) );
  INV_X1 U18379 ( .A(n15138), .ZN(n15142) );
  NAND2_X1 U18380 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n12763), .ZN(n15139) );
  OAI221_X1 U18381 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15142), 
        .C1(n15141), .C2(n15140), .A(n15139), .ZN(n15154) );
  INV_X1 U18382 ( .A(n15143), .ZN(n15146) );
  INV_X1 U18383 ( .A(n14861), .ZN(n15144) );
  AOI21_X1 U18384 ( .B1(n15146), .B2(n15145), .A(n15144), .ZN(n16073) );
  INV_X1 U18385 ( .A(n16073), .ZN(n15152) );
  INV_X1 U18386 ( .A(n15147), .ZN(n15150) );
  AOI21_X1 U18387 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(n16097) );
  INV_X1 U18388 ( .A(n16097), .ZN(n15151) );
  OAI22_X1 U18389 ( .A1(n16215), .A2(n15152), .B1(n16253), .B2(n15151), .ZN(
        n15153) );
  NOR3_X1 U18390 ( .A1(n15155), .A2(n15154), .A3(n15153), .ZN(n15156) );
  OAI21_X1 U18391 ( .B1(n16094), .B2(n16246), .A(n15156), .ZN(P2_U3024) );
  AND2_X1 U18392 ( .A1(n9891), .A2(n15157), .ZN(n15158) );
  NOR2_X1 U18393 ( .A1(n18865), .A2(n16253), .ZN(n15159) );
  AOI211_X1 U18394 ( .C1(n19257), .C2(n9883), .A(n15160), .B(n15159), .ZN(
        n15163) );
  OAI211_X1 U18395 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n15174), .B(n15161), .ZN(
        n15162) );
  OAI211_X1 U18396 ( .C1(n15176), .C2(n15164), .A(n15163), .B(n15162), .ZN(
        n15165) );
  AOI21_X1 U18397 ( .B1(n15166), .B2(n19262), .A(n15165), .ZN(n15167) );
  OAI21_X1 U18398 ( .B1(n15168), .B2(n16246), .A(n15167), .ZN(P2_U3026) );
  INV_X1 U18399 ( .A(n15169), .ZN(n15170) );
  AOI21_X1 U18400 ( .B1(n19257), .B2(n15171), .A(n15170), .ZN(n15172) );
  OAI21_X1 U18401 ( .B1(n18866), .B2(n16253), .A(n15172), .ZN(n15173) );
  AOI21_X1 U18402 ( .B1(n15174), .B2(n15177), .A(n15173), .ZN(n15175) );
  OAI21_X1 U18403 ( .B1(n15177), .B2(n15176), .A(n15175), .ZN(n15178) );
  AOI21_X1 U18404 ( .B1(n15179), .B2(n19262), .A(n15178), .ZN(n15180) );
  OAI21_X1 U18405 ( .B1(n15181), .B2(n16246), .A(n15180), .ZN(P2_U3027) );
  INV_X1 U18406 ( .A(n15182), .ZN(n15184) );
  AOI21_X1 U18407 ( .B1(n15184), .B2(n15183), .A(n15255), .ZN(n16189) );
  AOI21_X1 U18408 ( .B1(n15192), .B2(n15185), .A(n16189), .ZN(n15197) );
  OAI21_X1 U18409 ( .B1(n13679), .B2(n15187), .A(n15186), .ZN(n15188) );
  INV_X1 U18410 ( .A(n15188), .ZN(n18885) );
  NOR2_X1 U18411 ( .A1(n18888), .A2(n16253), .ZN(n15189) );
  AOI211_X1 U18412 ( .C1(n19257), .C2(n18885), .A(n15190), .B(n15189), .ZN(
        n15195) );
  INV_X1 U18413 ( .A(n15191), .ZN(n16195) );
  NOR2_X1 U18414 ( .A1(n16201), .A2(n16195), .ZN(n16188) );
  INV_X1 U18415 ( .A(n15192), .ZN(n15193) );
  NAND3_X1 U18416 ( .A1(n16188), .A2(n15193), .A3(n15196), .ZN(n15194) );
  OAI211_X1 U18417 ( .C1(n15197), .C2(n15196), .A(n15195), .B(n15194), .ZN(
        n15198) );
  AOI21_X1 U18418 ( .B1(n15199), .B2(n19262), .A(n15198), .ZN(n15200) );
  OAI21_X1 U18419 ( .B1(n15201), .B2(n16246), .A(n15200), .ZN(P2_U3028) );
  INV_X1 U18420 ( .A(n15204), .ZN(n15205) );
  OAI21_X1 U18421 ( .B1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15285), .A(
        n15231), .ZN(n15216) );
  INV_X1 U18422 ( .A(n15035), .ZN(n15209) );
  AOI21_X1 U18423 ( .B1(n15209), .B2(n19262), .A(n16188), .ZN(n15225) );
  NOR3_X1 U18424 ( .A1(n15225), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15210), .ZN(n15215) );
  NAND2_X1 U18425 ( .A1(n19257), .A2(n18895), .ZN(n15211) );
  OAI211_X1 U18426 ( .C1(n15213), .C2(n16253), .A(n15212), .B(n15211), .ZN(
        n15214) );
  AOI211_X1 U18427 ( .C1(n15216), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n15215), .B(n15214), .ZN(n15217) );
  OAI21_X1 U18428 ( .B1(n15218), .B2(n16246), .A(n15217), .ZN(P2_U3029) );
  INV_X1 U18429 ( .A(n15219), .ZN(n15228) );
  INV_X1 U18430 ( .A(n15220), .ZN(n15221) );
  NAND2_X1 U18431 ( .A1(n9888), .A2(n15221), .ZN(n15223) );
  AND2_X1 U18432 ( .A1(n15223), .A2(n15222), .ZN(n19128) );
  AOI22_X1 U18433 ( .A1(n19257), .A2(n19128), .B1(n12763), .B2(
        P2_REIP_REG_16__SCAN_IN), .ZN(n15224) );
  OAI21_X1 U18434 ( .B1(n19091), .B2(n16253), .A(n15224), .ZN(n15227) );
  NOR3_X1 U18435 ( .A1(n15225), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16187), .ZN(n15226) );
  AOI211_X1 U18436 ( .C1(n19263), .C2(n15228), .A(n15227), .B(n15226), .ZN(
        n15229) );
  OAI21_X1 U18437 ( .B1(n15231), .B2(n15230), .A(n15229), .ZN(P2_U3030) );
  NAND2_X1 U18438 ( .A1(n15233), .A2(n15232), .ZN(n15234) );
  XNOR2_X1 U18439 ( .A(n15235), .B(n15234), .ZN(n16118) );
  INV_X1 U18440 ( .A(n9877), .ZN(n15236) );
  OAI21_X1 U18441 ( .B1(n16124), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15236), .ZN(n16119) );
  OR2_X1 U18442 ( .A1(n16119), .A2(n16264), .ZN(n15249) );
  OR2_X1 U18443 ( .A1(n15238), .A2(n15237), .ZN(n15241) );
  INV_X1 U18444 ( .A(n15239), .ZN(n15240) );
  NAND2_X1 U18445 ( .A1(n15241), .A2(n15240), .ZN(n19143) );
  NAND2_X1 U18446 ( .A1(n18935), .A2(n19255), .ZN(n15245) );
  AOI211_X1 U18447 ( .C1(n12512), .C2(n15242), .A(n16196), .B(n16201), .ZN(
        n15243) );
  AOI21_X1 U18448 ( .B1(n19016), .B2(P2_REIP_REG_13__SCAN_IN), .A(n15243), 
        .ZN(n15244) );
  OAI211_X1 U18449 ( .C1(n16215), .C2(n19143), .A(n15245), .B(n15244), .ZN(
        n15246) );
  AOI21_X1 U18450 ( .B1(n15247), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15246), .ZN(n15248) );
  OAI211_X1 U18451 ( .C1(n16118), .C2(n16246), .A(n15249), .B(n15248), .ZN(
        P2_U3033) );
  NOR2_X1 U18452 ( .A1(n16144), .A2(n12506), .ZN(n16143) );
  OAI21_X1 U18453 ( .B1(n16143), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15250), .ZN(n16131) );
  XNOR2_X1 U18454 ( .A(n15251), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15252) );
  XNOR2_X1 U18455 ( .A(n15253), .B(n15252), .ZN(n16130) );
  NOR2_X1 U18456 ( .A1(n15255), .A2(n15254), .ZN(n16218) );
  NAND2_X1 U18457 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15256), .ZN(
        n16214) );
  AOI211_X1 U18458 ( .C1(n12506), .C2(n15258), .A(n15257), .B(n16214), .ZN(
        n15260) );
  NOR2_X1 U18459 ( .A1(n12685), .A2(n16232), .ZN(n15259) );
  AOI211_X1 U18460 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16218), .A(
        n15260), .B(n15259), .ZN(n15266) );
  OR2_X1 U18461 ( .A1(n15262), .A2(n15261), .ZN(n15263) );
  NAND2_X1 U18462 ( .A1(n15263), .A2(n13919), .ZN(n19149) );
  INV_X1 U18463 ( .A(n19149), .ZN(n15264) );
  AOI22_X1 U18464 ( .A1(n18947), .A2(n19255), .B1(n19257), .B2(n15264), .ZN(
        n15265) );
  OAI211_X1 U18465 ( .C1(n16130), .C2(n16246), .A(n15266), .B(n15265), .ZN(
        n15267) );
  INV_X1 U18466 ( .A(n15267), .ZN(n15268) );
  OAI21_X1 U18467 ( .B1(n16131), .B2(n16264), .A(n15268), .ZN(P2_U3035) );
  NAND3_X1 U18468 ( .A1(n15270), .A2(n15269), .A3(n19262), .ZN(n15281) );
  AOI21_X1 U18469 ( .B1(n16257), .B2(n15272), .A(n15271), .ZN(n16226) );
  NOR2_X1 U18470 ( .A1(n19862), .A2(n16232), .ZN(n15277) );
  OR2_X1 U18471 ( .A1(n15274), .A2(n15273), .ZN(n15275) );
  NAND2_X1 U18472 ( .A1(n15275), .A2(n16229), .ZN(n19160) );
  NOR2_X1 U18473 ( .A1(n16215), .A2(n19160), .ZN(n15276) );
  AOI211_X1 U18474 ( .C1(n18999), .C2(n19255), .A(n15277), .B(n15276), .ZN(
        n15278) );
  OAI21_X1 U18475 ( .B1(n16226), .B2(n16225), .A(n15278), .ZN(n15279) );
  AOI21_X1 U18476 ( .B1(n16224), .B2(n16225), .A(n15279), .ZN(n15280) );
  OAI211_X1 U18477 ( .C1(n15282), .C2(n16246), .A(n15281), .B(n15280), .ZN(
        P2_U3039) );
  XNOR2_X1 U18478 ( .A(n15284), .B(n15283), .ZN(n16174) );
  NOR2_X1 U18479 ( .A1(n15285), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n16242) );
  OR2_X1 U18480 ( .A1(n15286), .A2(n16242), .ZN(n19256) );
  XNOR2_X1 U18481 ( .A(n19031), .B(n15287), .ZN(n19171) );
  NOR2_X1 U18482 ( .A1(n13419), .A2(n15288), .ZN(n19260) );
  OAI221_X1 U18483 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n15289), .C2(n19259), .A(
        n19260), .ZN(n15290) );
  OAI21_X1 U18484 ( .B1(n16232), .B2(n15291), .A(n15290), .ZN(n15292) );
  AOI21_X1 U18485 ( .B1(n19020), .B2(n19255), .A(n15292), .ZN(n15293) );
  OAI21_X1 U18486 ( .B1(n19171), .B2(n16215), .A(n15293), .ZN(n15304) );
  OR2_X1 U18487 ( .A1(n15295), .A2(n15294), .ZN(n15302) );
  INV_X1 U18488 ( .A(n15296), .ZN(n15300) );
  NAND2_X1 U18489 ( .A1(n15298), .A2(n15297), .ZN(n15299) );
  NAND2_X1 U18490 ( .A1(n15300), .A2(n15299), .ZN(n15301) );
  NAND2_X1 U18491 ( .A1(n15302), .A2(n15301), .ZN(n16171) );
  NOR2_X1 U18492 ( .A1(n16171), .A2(n16264), .ZN(n15303) );
  AOI211_X1 U18493 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n19256), .A(
        n15304), .B(n15303), .ZN(n15305) );
  OAI21_X1 U18494 ( .B1(n16246), .B2(n16174), .A(n15305), .ZN(P2_U3041) );
  NAND2_X1 U18495 ( .A1(n13099), .A2(n15306), .ZN(n15320) );
  NAND2_X1 U18496 ( .A1(n12041), .A2(n15307), .ZN(n16278) );
  INV_X1 U18497 ( .A(n15314), .ZN(n15308) );
  NAND2_X1 U18498 ( .A1(n15313), .A2(n15308), .ZN(n16279) );
  INV_X1 U18499 ( .A(n15309), .ZN(n15310) );
  NAND2_X1 U18500 ( .A1(n15310), .A2(n11872), .ZN(n16276) );
  NAND2_X1 U18501 ( .A1(n16279), .A2(n16276), .ZN(n15311) );
  AOI21_X1 U18502 ( .B1(n16277), .B2(n16278), .A(n15311), .ZN(n15316) );
  INV_X1 U18503 ( .A(n16269), .ZN(n15312) );
  NAND2_X1 U18504 ( .A1(n16271), .A2(n15312), .ZN(n16287) );
  AOI22_X1 U18505 ( .A1(n16287), .A2(n16276), .B1(n15314), .B2(n15313), .ZN(
        n15315) );
  MUX2_X1 U18506 ( .A(n15316), .B(n15315), .S(n11987), .Z(n15318) );
  AND2_X1 U18507 ( .A1(n15318), .A2(n15317), .ZN(n15319) );
  NAND2_X1 U18508 ( .A1(n15320), .A2(n15319), .ZN(n16297) );
  INV_X1 U18509 ( .A(n16297), .ZN(n15321) );
  OAI22_X1 U18510 ( .A1(n19925), .A2(n19916), .B1(n15321), .B2(n19922), .ZN(
        n15322) );
  MUX2_X1 U18511 ( .A(n15322), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n19918), .Z(P2_U3596) );
  NOR2_X2 U18512 ( .A1(n19683), .A2(n19926), .ZN(n19823) );
  INV_X1 U18513 ( .A(n19352), .ZN(n15323) );
  NAND2_X1 U18514 ( .A1(n19728), .A2(n15323), .ZN(n15324) );
  OR2_X1 U18515 ( .A1(n19823), .A2(n15324), .ZN(n15325) );
  NAND2_X1 U18516 ( .A1(n19728), .A2(n19920), .ZN(n19923) );
  NOR2_X1 U18517 ( .A1(n19933), .A2(n15326), .ZN(n19818) );
  NOR2_X1 U18518 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19357) );
  NAND2_X1 U18519 ( .A1(n19357), .A2(n19949), .ZN(n19311) );
  NOR2_X1 U18520 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19311), .ZN(
        n19292) );
  NOR2_X1 U18521 ( .A1(n19818), .A2(n19292), .ZN(n15330) );
  OAI21_X1 U18522 ( .B1(n12114), .B2(n19292), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15327) );
  INV_X1 U18523 ( .A(n19296), .ZN(n15350) );
  NOR2_X2 U18524 ( .A1(n15328), .A2(n19503), .ZN(n19770) );
  INV_X1 U18525 ( .A(n19770), .ZN(n19307) );
  INV_X1 U18526 ( .A(n15329), .ZN(n15331) );
  NAND2_X1 U18527 ( .A1(n15331), .A2(n15330), .ZN(n15337) );
  NAND2_X1 U18528 ( .A1(n15332), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n15333) );
  NAND2_X1 U18529 ( .A1(n15333), .A2(n19971), .ZN(n15335) );
  INV_X1 U18530 ( .A(n19292), .ZN(n15334) );
  AOI21_X1 U18531 ( .B1(n15335), .B2(n15334), .A(n19503), .ZN(n15336) );
  INV_X1 U18532 ( .A(n19300), .ZN(n15348) );
  AOI22_X1 U18533 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19294), .ZN(n19781) );
  INV_X1 U18534 ( .A(n19823), .ZN(n15346) );
  AOI22_X1 U18535 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19294), .ZN(n19697) );
  AOI22_X1 U18536 ( .A1(n19778), .A2(n19352), .B1(n19769), .B2(n19292), .ZN(
        n15341) );
  OAI21_X1 U18537 ( .B1(n19781), .B2(n15346), .A(n15341), .ZN(n15342) );
  AOI21_X1 U18538 ( .B1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(n15348), .A(
        n15342), .ZN(n15343) );
  OAI21_X1 U18539 ( .B1(n15350), .B2(n19307), .A(n15343), .ZN(P2_U3048) );
  NOR2_X2 U18540 ( .A1(n19159), .A2(n19503), .ZN(n19820) );
  INV_X1 U18541 ( .A(n19820), .ZN(n19349) );
  AOI22_X1 U18542 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19294), .ZN(n19828) );
  AOI22_X1 U18543 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19294), .ZN(n19764) );
  AND2_X1 U18544 ( .A1(n15344), .A2(n19291), .ZN(n19819) );
  AOI22_X1 U18545 ( .A1(n19822), .A2(n19352), .B1(n19292), .B2(n19819), .ZN(
        n15345) );
  OAI21_X1 U18546 ( .B1(n19828), .B2(n15346), .A(n15345), .ZN(n15347) );
  AOI21_X1 U18547 ( .B1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n15348), .A(
        n15347), .ZN(n15349) );
  OAI21_X1 U18548 ( .B1(n15350), .B2(n19349), .A(n15349), .ZN(P2_U3055) );
  NOR3_X1 U18549 ( .A1(n13030), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19453) );
  INV_X1 U18550 ( .A(n19453), .ZN(n19456) );
  NOR2_X1 U18551 ( .A1(n19958), .A2(n19456), .ZN(n19473) );
  NAND2_X1 U18552 ( .A1(n19925), .A2(n19527), .ZN(n19499) );
  NOR2_X2 U18553 ( .A1(n19926), .A2(n19422), .ZN(n19523) );
  AOI21_X1 U18554 ( .B1(n19498), .B2(n19513), .A(n19920), .ZN(n15351) );
  NOR2_X1 U18555 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19504), .ZN(
        n19493) );
  AOI221_X1 U18556 ( .B1(n19473), .B2(n19971), .C1(n15351), .C2(n19971), .A(
        n19493), .ZN(n15356) );
  INV_X1 U18557 ( .A(n19493), .ZN(n15352) );
  NAND2_X1 U18558 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n15352), .ZN(n15353) );
  OR2_X1 U18559 ( .A1(n15354), .A2(n15353), .ZN(n15359) );
  NAND2_X1 U18560 ( .A1(n15359), .A2(n19776), .ZN(n15355) );
  INV_X1 U18561 ( .A(n19495), .ZN(n19481) );
  INV_X1 U18562 ( .A(n19781), .ZN(n19694) );
  AOI22_X1 U18563 ( .A1(n19523), .A2(n19778), .B1(n19490), .B2(n19694), .ZN(
        n15361) );
  NOR2_X1 U18564 ( .A1(n19473), .A2(n19493), .ZN(n15357) );
  OAI21_X1 U18565 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n15357), .A(n19979), 
        .ZN(n15358) );
  AND2_X1 U18566 ( .A1(n15359), .A2(n15358), .ZN(n19494) );
  AOI22_X1 U18567 ( .A1(n19494), .A2(n19770), .B1(n19769), .B2(n19493), .ZN(
        n15360) );
  OAI211_X1 U18568 ( .C1(n19481), .C2(n15362), .A(n15361), .B(n15360), .ZN(
        P2_U3096) );
  AOI22_X1 U18569 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15366) );
  AOI22_X1 U18570 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15365) );
  AOI22_X1 U18571 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n15364) );
  AOI22_X1 U18572 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15363) );
  NAND4_X1 U18573 ( .A1(n15366), .A2(n15365), .A3(n15364), .A4(n15363), .ZN(
        n15373) );
  AOI22_X1 U18574 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15371) );
  AOI22_X1 U18575 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15370) );
  AOI22_X1 U18576 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15369) );
  AOI22_X1 U18577 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15368) );
  NAND4_X1 U18578 ( .A1(n15371), .A2(n15370), .A3(n15369), .A4(n15368), .ZN(
        n15372) );
  NOR2_X1 U18579 ( .A1(n15373), .A2(n15372), .ZN(n16921) );
  AOI22_X1 U18580 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15377) );
  AOI22_X1 U18581 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15376) );
  AOI22_X1 U18582 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15375) );
  AOI22_X1 U18583 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15374) );
  NAND4_X1 U18584 ( .A1(n15377), .A2(n15376), .A3(n15375), .A4(n15374), .ZN(
        n15383) );
  AOI22_X1 U18585 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15381) );
  AOI22_X1 U18586 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15380) );
  AOI22_X1 U18587 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15379) );
  AOI22_X1 U18588 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n15378) );
  NAND4_X1 U18589 ( .A1(n15381), .A2(n15380), .A3(n15379), .A4(n15378), .ZN(
        n15382) );
  NOR2_X1 U18590 ( .A1(n15383), .A2(n15382), .ZN(n16932) );
  AOI22_X1 U18591 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15387) );
  AOI22_X1 U18592 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15386) );
  AOI22_X1 U18593 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15385) );
  AOI22_X1 U18594 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15384) );
  NAND4_X1 U18595 ( .A1(n15387), .A2(n15386), .A3(n15385), .A4(n15384), .ZN(
        n15393) );
  AOI22_X1 U18596 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15391) );
  AOI22_X1 U18597 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15390) );
  AOI22_X1 U18598 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15389) );
  AOI22_X1 U18599 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n15388) );
  NAND4_X1 U18600 ( .A1(n15391), .A2(n15390), .A3(n15389), .A4(n15388), .ZN(
        n15392) );
  NOR2_X1 U18601 ( .A1(n15393), .A2(n15392), .ZN(n16942) );
  AOI22_X1 U18602 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17024), .B1(
        P3_INSTQUEUE_REG_3__7__SCAN_IN), .B2(n17141), .ZN(n15397) );
  AOI22_X1 U18603 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15396) );
  AOI22_X1 U18604 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .B2(n17109), .ZN(n15395) );
  AOI22_X1 U18605 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17143), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15394) );
  NAND4_X1 U18606 ( .A1(n15397), .A2(n15396), .A3(n15395), .A4(n15394), .ZN(
        n15403) );
  AOI22_X1 U18607 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15401) );
  AOI22_X1 U18608 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n15400) );
  AOI22_X1 U18609 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17150), .B1(
        n11223), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15399) );
  AOI22_X1 U18610 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17152), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15398) );
  NAND4_X1 U18611 ( .A1(n15401), .A2(n15400), .A3(n15399), .A4(n15398), .ZN(
        n15402) );
  NOR2_X1 U18612 ( .A1(n15403), .A2(n15402), .ZN(n16943) );
  NOR2_X1 U18613 ( .A1(n16942), .A2(n16943), .ZN(n16941) );
  AOI22_X1 U18614 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15414) );
  AOI22_X1 U18615 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15413) );
  AOI22_X1 U18616 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15404) );
  OAI21_X1 U18617 ( .B1(n15405), .B2(n17192), .A(n15404), .ZN(n15411) );
  AOI22_X1 U18618 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15409) );
  AOI22_X1 U18619 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15408) );
  AOI22_X1 U18620 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n15407) );
  AOI22_X1 U18621 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n15406) );
  NAND4_X1 U18622 ( .A1(n15409), .A2(n15408), .A3(n15407), .A4(n15406), .ZN(
        n15410) );
  AOI211_X1 U18623 ( .C1(n17082), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n15411), .B(n15410), .ZN(n15412) );
  NAND3_X1 U18624 ( .A1(n15414), .A2(n15413), .A3(n15412), .ZN(n16937) );
  NAND2_X1 U18625 ( .A1(n16941), .A2(n16937), .ZN(n16936) );
  NOR2_X1 U18626 ( .A1(n16932), .A2(n16936), .ZN(n16931) );
  AOI22_X1 U18627 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15425) );
  INV_X1 U18628 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n15417) );
  AOI22_X1 U18629 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15416) );
  AOI22_X1 U18630 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15415) );
  OAI211_X1 U18631 ( .C1(n11237), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n15423) );
  AOI22_X1 U18632 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15421) );
  AOI22_X1 U18633 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15420) );
  AOI22_X1 U18634 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n15419) );
  AOI22_X1 U18635 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15418) );
  NAND4_X1 U18636 ( .A1(n15421), .A2(n15420), .A3(n15419), .A4(n15418), .ZN(
        n15422) );
  AOI211_X1 U18637 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15423), .B(n15422), .ZN(n15424) );
  NAND2_X1 U18638 ( .A1(n15425), .A2(n15424), .ZN(n16927) );
  NAND2_X1 U18639 ( .A1(n16931), .A2(n16927), .ZN(n16926) );
  NOR2_X1 U18640 ( .A1(n16921), .A2(n16926), .ZN(n16920) );
  AOI22_X1 U18641 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15436) );
  INV_X1 U18642 ( .A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15428) );
  AOI22_X1 U18643 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15427) );
  AOI22_X1 U18644 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15426) );
  OAI211_X1 U18645 ( .C1(n11237), .C2(n15428), .A(n15427), .B(n15426), .ZN(
        n15434) );
  AOI22_X1 U18646 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15432) );
  AOI22_X1 U18647 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15431) );
  AOI22_X1 U18648 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15430) );
  AOI22_X1 U18649 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15429) );
  NAND4_X1 U18650 ( .A1(n15432), .A2(n15431), .A3(n15430), .A4(n15429), .ZN(
        n15433) );
  AOI211_X1 U18651 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n15434), .B(n15433), .ZN(n15435) );
  NAND2_X1 U18652 ( .A1(n15436), .A2(n15435), .ZN(n15437) );
  NAND2_X1 U18653 ( .A1(n16920), .A2(n15437), .ZN(n16913) );
  OAI21_X1 U18654 ( .B1(n16920), .B2(n15437), .A(n16913), .ZN(n17220) );
  AND3_X1 U18655 ( .A1(n15439), .A2(n16989), .A3(n15438), .ZN(n15440) );
  NOR3_X2 U18656 ( .A1(n18808), .A2(n15442), .A3(n15581), .ZN(n17200) );
  AND2_X1 U18657 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16917) );
  NAND2_X1 U18658 ( .A1(n16989), .A2(n17200), .ZN(n17194) );
  INV_X1 U18659 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16882) );
  INV_X1 U18660 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16593) );
  INV_X1 U18661 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16973) );
  INV_X1 U18662 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16988) );
  INV_X1 U18663 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17017) );
  NAND4_X1 U18664 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(P3_EBX_REG_4__SCAN_IN), .ZN(n15445) );
  NAND4_X1 U18665 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(P3_EBX_REG_9__SCAN_IN), .A4(P3_EBX_REG_8__SCAN_IN), .ZN(n15444) );
  INV_X1 U18666 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16841) );
  NAND3_X1 U18667 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17187) );
  NOR2_X1 U18668 ( .A1(n16841), .A2(n17187), .ZN(n15460) );
  INV_X1 U18669 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n16697) );
  INV_X1 U18670 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16714) );
  INV_X1 U18671 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n15461) );
  NOR3_X1 U18672 ( .A1(n16697), .A2(n16714), .A3(n15461), .ZN(n17049) );
  NAND4_X1 U18673 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_15__SCAN_IN), 
        .A3(n15460), .A4(n17049), .ZN(n15443) );
  NOR3_X1 U18674 ( .A1(n15445), .A2(n15444), .A3(n15443), .ZN(n17031) );
  NAND3_X1 U18675 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17200), .A3(n17031), 
        .ZN(n17006) );
  NAND2_X1 U18676 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17002), .ZN(n17003) );
  NAND2_X1 U18677 ( .A1(n16989), .A2(n16972), .ZN(n16977) );
  NOR2_X1 U18678 ( .A1(n16973), .A2(n16977), .ZN(n16947) );
  NAND2_X1 U18679 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16947), .ZN(n16940) );
  NAND2_X1 U18680 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16946), .ZN(n16930) );
  NAND2_X1 U18681 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16935), .ZN(n16925) );
  NAND2_X1 U18682 ( .A1(n17191), .A2(n16925), .ZN(n16923) );
  OAI21_X1 U18683 ( .B1(n16917), .B2(n17194), .A(n16923), .ZN(n16915) );
  INV_X1 U18684 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16924) );
  NOR3_X1 U18685 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16924), .A3(n16925), .ZN(
        n15446) );
  AOI21_X1 U18686 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16915), .A(n15446), .ZN(
        n15447) );
  OAI21_X1 U18687 ( .B1(n17220), .B2(n17191), .A(n15447), .ZN(P3_U2675) );
  AOI22_X1 U18688 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15452) );
  AOI22_X1 U18689 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9831), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U18690 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15450) );
  AOI22_X1 U18691 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15449) );
  NAND4_X1 U18692 ( .A1(n15452), .A2(n15451), .A3(n15450), .A4(n15449), .ZN(
        n15459) );
  AOI22_X1 U18693 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15457) );
  AOI22_X1 U18694 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U18695 ( .A1(n15453), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15455) );
  AOI22_X1 U18696 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15454) );
  NAND4_X1 U18697 ( .A1(n15457), .A2(n15456), .A3(n15455), .A4(n15454), .ZN(
        n15458) );
  NOR2_X1 U18698 ( .A1(n15459), .A2(n15458), .ZN(n17293) );
  INV_X1 U18699 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16733) );
  INV_X1 U18700 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16762) );
  INV_X1 U18701 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17166) );
  INV_X1 U18702 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17173) );
  INV_X1 U18703 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16821) );
  NAND2_X1 U18704 ( .A1(n17200), .A2(n15460), .ZN(n17177) );
  NAND2_X1 U18705 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17181), .ZN(n17170) );
  NOR3_X1 U18706 ( .A1(n17166), .A2(n17173), .A3(n17170), .ZN(n17165) );
  NAND2_X1 U18707 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17165), .ZN(n17162) );
  NAND2_X1 U18708 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17140), .ZN(n17103) );
  NAND2_X1 U18709 ( .A1(n16989), .A2(n17105), .ZN(n17089) );
  NOR2_X1 U18710 ( .A1(n15461), .A2(n17089), .ZN(n17063) );
  NOR2_X1 U18711 ( .A1(n17197), .A2(n17063), .ZN(n17090) );
  AOI22_X1 U18712 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17090), .B1(n17063), 
        .B2(n16714), .ZN(n15462) );
  OAI21_X1 U18713 ( .B1(n17293), .B2(n17191), .A(n15462), .ZN(P3_U2690) );
  NOR2_X1 U18714 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18758), .ZN(
        n18149) );
  INV_X1 U18715 ( .A(n18149), .ZN(n18197) );
  INV_X1 U18716 ( .A(n15463), .ZN(n15464) );
  AOI211_X1 U18717 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n15464), .A(
        n17130), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18147) );
  INV_X1 U18718 ( .A(n18452), .ZN(n18497) );
  OAI211_X1 U18719 ( .C1(n18756), .C2(n18147), .A(n18497), .B(n15465), .ZN(
        n18154) );
  NAND2_X1 U18720 ( .A1(n18197), .A2(n18154), .ZN(n15468) );
  INV_X1 U18721 ( .A(n15468), .ZN(n15467) );
  INV_X1 U18722 ( .A(n18448), .ZN(n18401) );
  INV_X1 U18723 ( .A(n17791), .ZN(n17625) );
  INV_X1 U18724 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18621) );
  OAI22_X1 U18725 ( .A1(n17625), .A2(n18803), .B1(n18621), .B2(n18758), .ZN(
        n15470) );
  NAND3_X1 U18726 ( .A1(n18623), .A2(n18154), .A3(n15470), .ZN(n15466) );
  OAI221_X1 U18727 ( .B1(n18623), .B2(n15467), .C1(n18623), .C2(n18401), .A(
        n15466), .ZN(P3_U2864) );
  NAND2_X1 U18728 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18328) );
  NOR2_X1 U18729 ( .A1(n17625), .A2(n18803), .ZN(n15469) );
  AOI221_X1 U18730 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18328), .C1(n15469), 
        .C2(n18328), .A(n15468), .ZN(n18153) );
  OAI221_X1 U18731 ( .B1(n18448), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18448), .C2(n15470), .A(n18154), .ZN(n18151) );
  AOI22_X1 U18732 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18153), .B1(
        n18151), .B2(n18628), .ZN(P3_U2865) );
  INV_X1 U18733 ( .A(n18064), .ZN(n15474) );
  INV_X1 U18734 ( .A(n18126), .ZN(n18145) );
  NOR2_X1 U18735 ( .A1(n16364), .A2(n18145), .ZN(n15471) );
  AOI211_X1 U18736 ( .C1(n15474), .C2(n16367), .A(n15472), .B(n15471), .ZN(
        n15558) );
  INV_X1 U18737 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17472) );
  AOI21_X1 U18738 ( .B1(n17982), .B2(n17836), .A(n15473), .ZN(n16366) );
  AOI22_X1 U18739 ( .A1(n18126), .A2(n16326), .B1(n15474), .B2(n16327), .ZN(
        n15561) );
  OAI21_X1 U18740 ( .B1(n9821), .B2(n16366), .A(n15561), .ZN(n15475) );
  AOI21_X1 U18741 ( .B1(n18130), .B2(n17472), .A(n15475), .ZN(n15479) );
  AOI21_X1 U18742 ( .B1(n16342), .B2(n15477), .A(n15476), .ZN(n16346) );
  AOI22_X1 U18743 ( .A1(n9821), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n9811), .B2(
        n16346), .ZN(n15478) );
  OAI221_X1 U18744 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15558), 
        .C1(n16342), .C2(n15479), .A(n15478), .ZN(P3_U2833) );
  AOI22_X1 U18745 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19053), .ZN(n15503) );
  INV_X1 U18746 ( .A(n19072), .ZN(n18991) );
  AOI22_X1 U18747 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19081), .B1(
        n15480), .B2(n18991), .ZN(n15502) );
  AOI22_X1 U18748 ( .A1(n16097), .A2(n19075), .B1(n16073), .B2(n19069), .ZN(
        n15501) );
  OAI21_X1 U18749 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9885), .A(
        n15481), .ZN(n16100) );
  INV_X1 U18750 ( .A(n16100), .ZN(n15498) );
  AOI21_X1 U18751 ( .B1(n18930), .B2(n15492), .A(n15482), .ZN(n18934) );
  AOI21_X1 U18752 ( .B1(n18955), .B2(n15491), .A(n15483), .ZN(n18958) );
  AOI21_X1 U18753 ( .B1(n16178), .B2(n15486), .A(n15489), .ZN(n19019) );
  NOR2_X1 U18754 ( .A1(n15485), .A2(n15484), .ZN(n19040) );
  OAI21_X1 U18755 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n15487), .A(
        n15486), .ZN(n19238) );
  NAND2_X1 U18756 ( .A1(n19040), .A2(n19238), .ZN(n19017) );
  NOR2_X1 U18757 ( .A1(n19019), .A2(n19017), .ZN(n19006) );
  OAI21_X1 U18758 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n15489), .A(
        n15488), .ZN(n19007) );
  NAND2_X1 U18759 ( .A1(n19006), .A2(n19007), .ZN(n18996) );
  NOR2_X1 U18760 ( .A1(n18998), .A2(n18996), .ZN(n18985) );
  OAI21_X1 U18761 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n15056), .A(
        n15490), .ZN(n18986) );
  NAND2_X1 U18762 ( .A1(n18985), .A2(n18986), .ZN(n18974) );
  NOR2_X1 U18763 ( .A1(n18976), .A2(n18974), .ZN(n18964) );
  OAI21_X1 U18764 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13943), .A(
        n15491), .ZN(n18965) );
  NAND2_X1 U18765 ( .A1(n18964), .A2(n18965), .ZN(n18950) );
  NOR2_X1 U18766 ( .A1(n18958), .A2(n18950), .ZN(n18949) );
  OAI21_X1 U18767 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15483), .A(
        n15492), .ZN(n18938) );
  NAND2_X1 U18768 ( .A1(n18949), .A2(n18938), .ZN(n18928) );
  NOR2_X1 U18769 ( .A1(n18934), .A2(n18928), .ZN(n18927) );
  OAI21_X1 U18770 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15482), .A(
        n15493), .ZN(n18922) );
  NAND2_X1 U18771 ( .A1(n18927), .A2(n18922), .ZN(n18912) );
  NOR2_X1 U18772 ( .A1(n18914), .A2(n18912), .ZN(n18903) );
  NAND2_X1 U18773 ( .A1(n18903), .A2(n18904), .ZN(n18889) );
  NOR2_X1 U18774 ( .A1(n18891), .A2(n18889), .ZN(n18881) );
  INV_X1 U18775 ( .A(n15495), .ZN(n18858) );
  OR2_X1 U18776 ( .A1(n18869), .A2(n18858), .ZN(n15496) );
  NAND2_X1 U18777 ( .A1(n10236), .A2(n10235), .ZN(n18856) );
  AOI21_X1 U18778 ( .B1(n15498), .B2(n15497), .A(n15964), .ZN(n15499) );
  NAND2_X1 U18779 ( .A1(n19058), .A2(n15499), .ZN(n15500) );
  NAND4_X1 U18780 ( .A1(n15503), .A2(n15502), .A3(n15501), .A4(n15500), .ZN(
        P2_U2833) );
  NAND2_X1 U18781 ( .A1(n15505), .A2(n15504), .ZN(n15510) );
  AND2_X1 U18782 ( .A1(n15506), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15507) );
  OR3_X1 U18783 ( .A1(n15508), .A2(n15507), .A3(n20570), .ZN(n15511) );
  NAND2_X1 U18784 ( .A1(n15511), .A2(n20531), .ZN(n15509) );
  NAND2_X1 U18785 ( .A1(n15510), .A2(n15509), .ZN(n15513) );
  OR2_X1 U18786 ( .A1(n15511), .A2(n20531), .ZN(n15512) );
  NAND2_X1 U18787 ( .A1(n15513), .A2(n15512), .ZN(n15514) );
  AND2_X1 U18788 ( .A1(n15514), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n15519) );
  INV_X1 U18789 ( .A(n15514), .ZN(n15516) );
  NAND2_X1 U18790 ( .A1(n15516), .A2(n15515), .ZN(n15517) );
  OAI21_X1 U18791 ( .B1(n15519), .B2(n15518), .A(n15517), .ZN(n15521) );
  NAND2_X1 U18792 ( .A1(n15523), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15520) );
  NAND2_X1 U18793 ( .A1(n15521), .A2(n15520), .ZN(n15522) );
  OAI21_X1 U18794 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15523), .A(
        n15522), .ZN(n15524) );
  NAND2_X1 U18795 ( .A1(n15524), .A2(n20148), .ZN(n15536) );
  INV_X1 U18796 ( .A(n15525), .ZN(n15531) );
  INV_X1 U18797 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21005) );
  NAND2_X1 U18798 ( .A1(n15526), .A2(n21005), .ZN(n15527) );
  NAND2_X1 U18799 ( .A1(n15528), .A2(n15527), .ZN(n15529) );
  AND4_X1 U18800 ( .A1(n15532), .A2(n15531), .A3(n15530), .A4(n15529), .ZN(
        n15533) );
  AND2_X1 U18801 ( .A1(n15534), .A2(n15533), .ZN(n15535) );
  INV_X1 U18802 ( .A(n15549), .ZN(n15544) );
  NAND4_X1 U18803 ( .A1(n15539), .A2(n15538), .A3(n15537), .A4(n21127), .ZN(
        n15542) );
  OAI21_X1 U18804 ( .B1(n15540), .B2(n20800), .A(n15548), .ZN(n15541) );
  OAI21_X1 U18805 ( .B1(n15543), .B2(n15542), .A(n15541), .ZN(n15948) );
  AOI221_X1 U18806 ( .B1(n20718), .B2(n20717), .C1(n15544), .C2(n20717), .A(
        n15948), .ZN(n15953) );
  AOI211_X1 U18807 ( .C1(n15563), .C2(n20721), .A(n15546), .B(n15545), .ZN(
        n15547) );
  OAI21_X1 U18808 ( .B1(n15549), .B2(n15548), .A(n15547), .ZN(n15550) );
  NOR2_X1 U18809 ( .A1(n15953), .A2(n15550), .ZN(n15554) );
  NAND2_X1 U18810 ( .A1(n20804), .A2(n15551), .ZN(n15552) );
  NAND2_X1 U18811 ( .A1(n20718), .A2(n15552), .ZN(n15553) );
  OAI22_X1 U18812 ( .A1(n15554), .A2(n20718), .B1(n15953), .B2(n15553), .ZN(
        P1_U3161) );
  NAND2_X1 U18813 ( .A1(n15556), .A2(n15555), .ZN(n15557) );
  INV_X1 U18814 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18742) );
  NOR2_X1 U18815 ( .A1(n18036), .A2(n18742), .ZN(n16329) );
  NOR3_X1 U18816 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15558), .A3(
        n16342), .ZN(n15559) );
  OAI221_X1 U18817 ( .B1(n16336), .B2(n15562), .C1(n16336), .C2(n15561), .A(
        n15560), .ZN(P3_U2832) );
  INV_X1 U18818 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20735) );
  INV_X1 U18819 ( .A(HOLD), .ZN(n20724) );
  NOR2_X1 U18820 ( .A1(n20735), .A2(n20724), .ZN(n20726) );
  AOI22_X1 U18821 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15565) );
  NAND2_X1 U18822 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15563), .ZN(n20723) );
  OAI211_X1 U18823 ( .C1(n20726), .C2(n15565), .A(n15564), .B(n20723), .ZN(
        P1_U3195) );
  AND2_X1 U18824 ( .A1(n15566), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  AOI21_X1 U18825 ( .B1(n15568), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15567), .ZN(n15732) );
  NAND2_X1 U18826 ( .A1(n15570), .A2(n15569), .ZN(n15576) );
  AOI22_X1 U18827 ( .A1(n15571), .A2(n15932), .B1(n15899), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15575) );
  OR2_X1 U18828 ( .A1(n15573), .A2(n15572), .ZN(n15574) );
  OAI211_X1 U18829 ( .C1(n15804), .C2(n15576), .A(n15575), .B(n15574), .ZN(
        n15577) );
  INV_X1 U18830 ( .A(n15577), .ZN(n15578) );
  OAI21_X1 U18831 ( .B1(n15732), .B2(n20138), .A(n15578), .ZN(P1_U3011) );
  NOR2_X1 U18832 ( .A1(n19980), .A2(n13470), .ZN(n19830) );
  AOI21_X1 U18833 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n13470), .A(n19830), 
        .ZN(n15579) );
  INV_X1 U18834 ( .A(n16324), .ZN(n15580) );
  AOI221_X1 U18835 ( .B1(n15579), .B2(n19979), .C1(n13474), .C2(n19979), .A(
        n15580), .ZN(P2_U3178) );
  AOI221_X1 U18836 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15580), .C1(n19962), .C2(
        n15580), .A(n19776), .ZN(n19959) );
  INV_X1 U18837 ( .A(n19959), .ZN(n19956) );
  NOR2_X1 U18838 ( .A1(n16303), .A2(n19956), .ZN(P2_U3047) );
  NOR3_X1 U18839 ( .A1(n18164), .A2(n18157), .A3(n15581), .ZN(n15582) );
  INV_X1 U18840 ( .A(n17342), .ZN(n15587) );
  NAND2_X1 U18841 ( .A1(n16989), .A2(n15587), .ZN(n17335) );
  INV_X1 U18842 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17412) );
  NAND2_X1 U18843 ( .A1(n17283), .A2(n15584), .ZN(n17341) );
  INV_X1 U18844 ( .A(n17341), .ZN(n17343) );
  AOI22_X1 U18845 ( .A1(n17343), .A2(BUF2_REG_0__SCAN_IN), .B1(n17316), .B2(
        n15585), .ZN(n15586) );
  OAI221_X1 U18846 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17335), .C1(n17412), 
        .C2(n15587), .A(n15586), .ZN(P3_U2735) );
  NAND2_X1 U18847 ( .A1(n15589), .A2(n15588), .ZN(n15592) );
  INV_X1 U18848 ( .A(n18846), .ZN(n15590) );
  OAI22_X1 U18849 ( .A1(n16215), .A2(n15590), .B1(n19882), .B2(n16232), .ZN(
        n15591) );
  AOI21_X1 U18850 ( .B1(n15593), .B2(n15592), .A(n15591), .ZN(n15598) );
  OAI22_X1 U18851 ( .A1(n15595), .A2(n16264), .B1(n16253), .B2(n15594), .ZN(
        n15596) );
  INV_X1 U18852 ( .A(n15596), .ZN(n15597) );
  OAI211_X1 U18853 ( .C1(n16246), .C2(n15599), .A(n15598), .B(n15597), .ZN(
        P2_U3025) );
  OAI21_X1 U18854 ( .B1(n15600), .B2(n15630), .A(n20763), .ZN(n15601) );
  AOI22_X1 U18855 ( .A1(n15602), .A2(n15601), .B1(P1_EBX_REG_23__SCAN_IN), 
        .B2(n20061), .ZN(n15608) );
  OAI22_X1 U18856 ( .A1(n15604), .A2(n15623), .B1(n15603), .B2(n20049), .ZN(
        n15605) );
  AOI21_X1 U18857 ( .B1(n15606), .B2(n20053), .A(n15605), .ZN(n15607) );
  OAI211_X1 U18858 ( .C1(n15609), .C2(n20064), .A(n15608), .B(n15607), .ZN(
        P1_U2817) );
  INV_X1 U18859 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n20959) );
  OAI22_X1 U18860 ( .A1(n20063), .A2(n15726), .B1(n20959), .B2(n15688), .ZN(
        n15610) );
  AOI21_X1 U18861 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20024), .A(
        n15610), .ZN(n15617) );
  AOI21_X1 U18862 ( .B1(n15612), .B2(n9836), .A(n15611), .ZN(n15801) );
  AOI22_X1 U18863 ( .A1(n15723), .A2(n20025), .B1(n15801), .B2(n20067), .ZN(
        n15616) );
  NOR2_X1 U18864 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15630), .ZN(n15618) );
  OAI21_X1 U18865 ( .B1(n15620), .B2(n15618), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15615) );
  INV_X1 U18866 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n21144) );
  NAND3_X1 U18867 ( .A1(n15644), .A2(n15613), .A3(n21144), .ZN(n15614) );
  NAND4_X1 U18868 ( .A1(n15617), .A2(n15616), .A3(n15615), .A4(n15614), .ZN(
        P1_U2818) );
  AOI22_X1 U18869 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15620), .B1(n15619), 
        .B2(n15618), .ZN(n15622) );
  AOI22_X1 U18870 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20046), .B2(P1_EBX_REG_21__SCAN_IN), .ZN(n15621) );
  OAI211_X1 U18871 ( .C1(n15624), .C2(n15623), .A(n15622), .B(n15621), .ZN(
        n15625) );
  AOI21_X1 U18872 ( .B1(n15626), .B2(n20053), .A(n15625), .ZN(n15627) );
  OAI21_X1 U18873 ( .B1(n15628), .B2(n20049), .A(n15627), .ZN(P1_U2819) );
  OAI221_X1 U18874 ( .B1(n15630), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n15630), 
        .C2(n15643), .A(n15629), .ZN(n15631) );
  AOI22_X1 U18875 ( .A1(n15632), .A2(n20053), .B1(P1_REIP_REG_19__SCAN_IN), 
        .B2(n15631), .ZN(n15640) );
  NAND2_X1 U18876 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15636) );
  OAI21_X1 U18877 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15633), .A(n20135), 
        .ZN(n15634) );
  AOI21_X1 U18878 ( .B1(n20046), .B2(P1_EBX_REG_19__SCAN_IN), .A(n15634), .ZN(
        n15635) );
  NAND2_X1 U18879 ( .A1(n15636), .A2(n15635), .ZN(n15637) );
  AOI21_X1 U18880 ( .B1(n15638), .B2(n20025), .A(n15637), .ZN(n15639) );
  OAI211_X1 U18881 ( .C1(n20049), .C2(n15641), .A(n15640), .B(n15639), .ZN(
        P1_U2821) );
  AOI22_X1 U18882 ( .A1(n15642), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_EBX_REG_18__SCAN_IN), .B2(n20061), .ZN(n15646) );
  INV_X1 U18883 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20933) );
  NAND3_X1 U18884 ( .A1(n15644), .A2(n15643), .A3(n20933), .ZN(n15645) );
  NAND2_X1 U18885 ( .A1(n15646), .A2(n15645), .ZN(n15647) );
  AOI211_X1 U18886 ( .C1(n20024), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15899), .B(n15647), .ZN(n15655) );
  INV_X1 U18887 ( .A(n15648), .ZN(n15653) );
  INV_X1 U18888 ( .A(n15649), .ZN(n15651) );
  OAI21_X1 U18889 ( .B1(n15668), .B2(n15651), .A(n15650), .ZN(n15652) );
  NAND2_X1 U18890 ( .A1(n15653), .A2(n15652), .ZN(n15831) );
  INV_X1 U18891 ( .A(n15831), .ZN(n15707) );
  AOI22_X1 U18892 ( .A1(n15708), .A2(n20025), .B1(n15707), .B2(n20067), .ZN(
        n15654) );
  OAI211_X1 U18893 ( .C1(n15656), .C2(n20063), .A(n15655), .B(n15654), .ZN(
        P1_U2822) );
  AOI21_X1 U18894 ( .B1(n15657), .B2(n21124), .A(n15678), .ZN(n15672) );
  NAND2_X1 U18895 ( .A1(n20061), .A2(P1_EBX_REG_16__SCAN_IN), .ZN(n15658) );
  OAI211_X1 U18896 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(n15659), .A(n15658), 
        .B(n20135), .ZN(n15662) );
  INV_X1 U18897 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15660) );
  NOR2_X1 U18898 ( .A1(n20064), .A2(n15660), .ZN(n15661) );
  AOI211_X1 U18899 ( .C1(n20053), .C2(n15663), .A(n15662), .B(n15661), .ZN(
        n15671) );
  INV_X1 U18900 ( .A(n15665), .ZN(n15666) );
  OAI21_X1 U18901 ( .B1(n15676), .B2(n15667), .A(n15666), .ZN(n15669) );
  AND2_X1 U18902 ( .A1(n15669), .A2(n15668), .ZN(n15847) );
  AOI22_X1 U18903 ( .A1(n15738), .A2(n20025), .B1(n15847), .B2(n20067), .ZN(
        n15670) );
  OAI211_X1 U18904 ( .C1(n15672), .C2(n20752), .A(n15671), .B(n15670), .ZN(
        P1_U2824) );
  AOI22_X1 U18905 ( .A1(n20024), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P1_EBX_REG_14__SCAN_IN), .B2(n20061), .ZN(n15683) );
  OR2_X1 U18906 ( .A1(n15674), .A2(n15673), .ZN(n15675) );
  AND2_X1 U18907 ( .A1(n15676), .A2(n15675), .ZN(n15862) );
  AOI21_X1 U18908 ( .B1(n15862), .B2(n20067), .A(n15899), .ZN(n15682) );
  INV_X1 U18909 ( .A(n15713), .ZN(n15749) );
  AOI22_X1 U18910 ( .A1(n15749), .A2(n20025), .B1(n20053), .B2(n15748), .ZN(
        n15681) );
  INV_X1 U18911 ( .A(n15677), .ZN(n20037) );
  OAI221_X1 U18912 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(n15679), .C1(
        P1_REIP_REG_14__SCAN_IN), .C2(n20037), .A(n15678), .ZN(n15680) );
  NAND4_X1 U18913 ( .A1(n15683), .A2(n15682), .A3(n15681), .A4(n15680), .ZN(
        P1_U2826) );
  INV_X1 U18914 ( .A(n15684), .ZN(n15701) );
  AOI21_X1 U18915 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n15701), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n15694) );
  OAI21_X1 U18916 ( .B1(n15696), .B2(n15697), .A(n15685), .ZN(n15687) );
  AND2_X1 U18917 ( .A1(n15687), .A2(n15686), .ZN(n15892) );
  INV_X1 U18918 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15717) );
  OAI22_X1 U18919 ( .A1(n20064), .A2(n15689), .B1(n15717), .B2(n15688), .ZN(
        n15690) );
  AOI211_X1 U18920 ( .C1(n15892), .C2(n20067), .A(n15899), .B(n15690), .ZN(
        n15693) );
  INV_X1 U18921 ( .A(n15691), .ZN(n15758) );
  AOI22_X1 U18922 ( .A1(n15759), .A2(n20053), .B1(n20025), .B2(n15758), .ZN(
        n15692) );
  OAI211_X1 U18923 ( .C1(n15695), .C2(n15694), .A(n15693), .B(n15692), .ZN(
        P1_U2828) );
  INV_X1 U18924 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20987) );
  INV_X1 U18925 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15699) );
  XOR2_X1 U18926 ( .A(n15697), .B(n15696), .Z(n15900) );
  AOI22_X1 U18927 ( .A1(n15900), .A2(n20067), .B1(n20046), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n15698) );
  OAI211_X1 U18928 ( .C1(n20064), .C2(n15699), .A(n15698), .B(n20135), .ZN(
        n15700) );
  AOI221_X1 U18929 ( .B1(n15702), .B2(P1_REIP_REG_11__SCAN_IN), .C1(n15701), 
        .C2(n20987), .A(n15700), .ZN(n15705) );
  INV_X1 U18930 ( .A(n15703), .ZN(n15769) );
  NAND2_X1 U18931 ( .A1(n20025), .A2(n15769), .ZN(n15704) );
  OAI211_X1 U18932 ( .C1(n20063), .C2(n15772), .A(n15705), .B(n15704), .ZN(
        P1_U2829) );
  AOI22_X1 U18933 ( .A1(n15723), .A2(n20074), .B1(n15801), .B2(n20073), .ZN(
        n15706) );
  OAI21_X1 U18934 ( .B1(n20078), .B2(n20959), .A(n15706), .ZN(P1_U2850) );
  INV_X1 U18935 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21059) );
  AOI22_X1 U18936 ( .A1(n15708), .A2(n20074), .B1(n15707), .B2(n20073), .ZN(
        n15709) );
  OAI21_X1 U18937 ( .B1(n20078), .B2(n21059), .A(n15709), .ZN(P1_U2854) );
  AOI22_X1 U18938 ( .A1(n15738), .A2(n20074), .B1(n15847), .B2(n20073), .ZN(
        n15710) );
  OAI21_X1 U18939 ( .B1(n20078), .B2(n21134), .A(n15710), .ZN(P1_U2856) );
  INV_X1 U18940 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n20907) );
  INV_X1 U18941 ( .A(n15862), .ZN(n15711) );
  OAI22_X1 U18942 ( .A1(n15713), .A2(n14439), .B1(n15712), .B2(n15711), .ZN(
        n15714) );
  INV_X1 U18943 ( .A(n15714), .ZN(n15715) );
  OAI21_X1 U18944 ( .B1(n20078), .B2(n20907), .A(n15715), .ZN(P1_U2858) );
  AOI22_X1 U18945 ( .A1(n15758), .A2(n20074), .B1(n20073), .B2(n15892), .ZN(
        n15716) );
  OAI21_X1 U18946 ( .B1(n20078), .B2(n15717), .A(n15716), .ZN(P1_U2860) );
  AOI22_X1 U18947 ( .A1(n15769), .A2(n20074), .B1(n20073), .B2(n15900), .ZN(
        n15718) );
  OAI21_X1 U18948 ( .B1(n20078), .B2(n15719), .A(n15718), .ZN(P1_U2861) );
  AOI22_X1 U18949 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15725) );
  NAND2_X1 U18950 ( .A1(n15721), .A2(n15720), .ZN(n15722) );
  XNOR2_X1 U18951 ( .A(n15722), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15802) );
  AOI22_X1 U18952 ( .A1(n15802), .A2(n20127), .B1(n15786), .B2(n15723), .ZN(
        n15724) );
  OAI211_X1 U18953 ( .C1(n15782), .C2(n15726), .A(n15725), .B(n15724), .ZN(
        P1_U2977) );
  AOI22_X1 U18954 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15899), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15731) );
  INV_X1 U18955 ( .A(n15727), .ZN(n15728) );
  AOI22_X1 U18956 ( .A1(n15729), .A2(n15786), .B1(n15728), .B2(n15783), .ZN(
        n15730) );
  OAI211_X1 U18957 ( .C1(n15732), .C2(n19996), .A(n15731), .B(n15730), .ZN(
        P1_U2979) );
  AOI22_X1 U18958 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15740) );
  AOI21_X1 U18959 ( .B1(n15735), .B2(n15734), .A(n15733), .ZN(n15736) );
  XOR2_X1 U18960 ( .A(n15737), .B(n15736), .Z(n15848) );
  AOI22_X1 U18961 ( .A1(n15848), .A2(n20127), .B1(n15786), .B2(n15738), .ZN(
        n15739) );
  OAI211_X1 U18962 ( .C1(n15782), .C2(n15741), .A(n15740), .B(n15739), .ZN(
        P1_U2983) );
  INV_X1 U18963 ( .A(n15742), .ZN(n15743) );
  AOI21_X1 U18964 ( .B1(n15745), .B2(n15744), .A(n15743), .ZN(n15747) );
  XNOR2_X1 U18965 ( .A(n9820), .B(n15863), .ZN(n15746) );
  XNOR2_X1 U18966 ( .A(n15747), .B(n15746), .ZN(n15868) );
  AOI22_X1 U18967 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n15899), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15751) );
  AOI22_X1 U18968 ( .A1(n15749), .A2(n15786), .B1(n15783), .B2(n15748), .ZN(
        n15750) );
  OAI211_X1 U18969 ( .C1(n15868), .C2(n19996), .A(n15751), .B(n15750), .ZN(
        P1_U2985) );
  AOI21_X1 U18970 ( .B1(n15754), .B2(n15753), .A(n15752), .ZN(n15757) );
  INV_X1 U18971 ( .A(n15755), .ZN(n15756) );
  NOR2_X1 U18972 ( .A1(n15757), .A2(n15756), .ZN(n15897) );
  AOI22_X1 U18973 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15761) );
  AOI22_X1 U18974 ( .A1(n15783), .A2(n15759), .B1(n15786), .B2(n15758), .ZN(
        n15760) );
  OAI211_X1 U18975 ( .C1(n15897), .C2(n19996), .A(n15761), .B(n15760), .ZN(
        P1_U2987) );
  AOI22_X1 U18976 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15771) );
  NAND2_X1 U18977 ( .A1(n9820), .A2(n15762), .ZN(n15766) );
  NAND2_X1 U18978 ( .A1(n14587), .A2(n15763), .ZN(n15764) );
  OAI22_X1 U18979 ( .A1(n15766), .A2(n15763), .B1(n15765), .B2(n15764), .ZN(
        n15767) );
  XNOR2_X1 U18980 ( .A(n15768), .B(n15767), .ZN(n15901) );
  AOI22_X1 U18981 ( .A1(n20127), .A2(n15901), .B1(n15786), .B2(n15769), .ZN(
        n15770) );
  OAI211_X1 U18982 ( .C1(n15782), .C2(n15772), .A(n15771), .B(n15770), .ZN(
        P1_U2988) );
  AOI22_X1 U18983 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15775) );
  AOI22_X1 U18984 ( .A1(n15773), .A2(n20127), .B1(n15786), .B2(n20017), .ZN(
        n15774) );
  OAI211_X1 U18985 ( .C1(n15782), .C2(n20020), .A(n15775), .B(n15774), .ZN(
        P1_U2992) );
  AOI22_X1 U18986 ( .A1(n20125), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n15935), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15781) );
  NAND2_X1 U18987 ( .A1(n15778), .A2(n15777), .ZN(n15779) );
  XNOR2_X1 U18988 ( .A(n15776), .B(n15779), .ZN(n15934) );
  AOI22_X1 U18989 ( .A1(n15934), .A2(n20127), .B1(n15786), .B2(n20075), .ZN(
        n15780) );
  OAI211_X1 U18990 ( .C1(n15782), .C2(n20029), .A(n15781), .B(n15780), .ZN(
        P1_U2993) );
  INV_X1 U18991 ( .A(n20039), .ZN(n15784) );
  AOI222_X1 U18992 ( .A1(n15787), .A2(n20127), .B1(n15786), .B2(n15785), .C1(
        n15784), .C2(n15783), .ZN(n15789) );
  OAI211_X1 U18993 ( .C1(n20033), .C2(n15790), .A(n15789), .B(n15788), .ZN(
        P1_U2994) );
  AOI22_X1 U18994 ( .A1(n15792), .A2(n15933), .B1(n15932), .B2(n15791), .ZN(
        n15800) );
  NAND2_X1 U18995 ( .A1(n15935), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15799) );
  OAI21_X1 U18996 ( .B1(n15794), .B2(n15793), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15798) );
  OR3_X1 U18997 ( .A1(n15796), .A2(n15795), .A3(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15797) );
  NAND4_X1 U18998 ( .A1(n15800), .A2(n15799), .A3(n15798), .A4(n15797), .ZN(
        P1_U3005) );
  AOI22_X1 U18999 ( .A1(n15802), .A2(n15933), .B1(n15932), .B2(n15801), .ZN(
        n15811) );
  INV_X1 U19000 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15803) );
  OAI21_X1 U19001 ( .B1(n15805), .B2(n15804), .A(n15803), .ZN(n15806) );
  OAI221_X1 U19002 ( .B1(n15809), .B2(n15808), .C1(n15809), .C2(n15807), .A(
        n15806), .ZN(n15810) );
  OAI211_X1 U19003 ( .C1(n21144), .C2(n20135), .A(n15811), .B(n15810), .ZN(
        P1_U3009) );
  NAND2_X1 U19004 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15812), .ZN(
        n15820) );
  INV_X1 U19005 ( .A(n15813), .ZN(n15824) );
  INV_X1 U19006 ( .A(n15814), .ZN(n15815) );
  NAND2_X1 U19007 ( .A1(n15816), .A2(n15815), .ZN(n15872) );
  OAI221_X1 U19008 ( .B1(n15886), .B2(n15817), .C1(n15886), .C2(n15824), .A(
        n15872), .ZN(n15818) );
  AOI211_X1 U19009 ( .C1(n15821), .C2(n15820), .A(n15819), .B(n15818), .ZN(
        n15879) );
  NOR3_X1 U19010 ( .A1(n15823), .A2(n15822), .A3(n15873), .ZN(n15826) );
  OAI211_X1 U19011 ( .C1(n15826), .C2(n15825), .A(n15824), .B(n15878), .ZN(
        n15876) );
  NAND2_X1 U19012 ( .A1(n15879), .A2(n15876), .ZN(n15865) );
  AOI21_X1 U19013 ( .B1(n15829), .B2(n15827), .A(n15865), .ZN(n15842) );
  NAND2_X1 U19014 ( .A1(n15864), .A2(n15835), .ZN(n15830) );
  OAI222_X1 U19015 ( .A1(n15831), .A2(n20137), .B1(n15830), .B2(n15829), .C1(
        n20138), .C2(n15828), .ZN(n15832) );
  INV_X1 U19016 ( .A(n15832), .ZN(n15834) );
  NAND2_X1 U19017 ( .A1(n15935), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15833) );
  OAI211_X1 U19018 ( .C1(n15842), .C2(n15835), .A(n15834), .B(n15833), .ZN(
        P1_U3013) );
  INV_X1 U19019 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15843) );
  NOR3_X1 U19020 ( .A1(n15863), .A2(n15844), .A3(n15843), .ZN(n15836) );
  AOI21_X1 U19021 ( .B1(n15864), .B2(n15836), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15841) );
  AOI22_X1 U19022 ( .A1(n15838), .A2(n15933), .B1(n15932), .B2(n15837), .ZN(
        n15840) );
  NAND2_X1 U19023 ( .A1(n15935), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15839) );
  OAI211_X1 U19024 ( .C1(n15842), .C2(n15841), .A(n15840), .B(n15839), .ZN(
        P1_U3014) );
  NOR2_X1 U19025 ( .A1(n15844), .A2(n15843), .ZN(n15852) );
  OAI211_X1 U19026 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n15864), .ZN(n15851) );
  INV_X1 U19027 ( .A(n15865), .ZN(n15845) );
  OAI21_X1 U19028 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15846), .A(
        n15845), .ZN(n15858) );
  AOI22_X1 U19029 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15858), .B1(
        n15899), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15850) );
  AOI22_X1 U19030 ( .A1(n15848), .A2(n15933), .B1(n15932), .B2(n15847), .ZN(
        n15849) );
  OAI211_X1 U19031 ( .C1(n15852), .C2(n15851), .A(n15850), .B(n15849), .ZN(
        P1_U3015) );
  NAND2_X1 U19032 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15864), .ZN(
        n15861) );
  INV_X1 U19033 ( .A(n15853), .ZN(n15856) );
  INV_X1 U19034 ( .A(n15854), .ZN(n15855) );
  AOI21_X1 U19035 ( .B1(n15856), .B2(n15932), .A(n15855), .ZN(n15860) );
  AOI22_X1 U19036 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15858), .B1(
        n15933), .B2(n15857), .ZN(n15859) );
  OAI211_X1 U19037 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15861), .A(
        n15860), .B(n15859), .ZN(P1_U3016) );
  AOI22_X1 U19038 ( .A1(n15932), .A2(n15862), .B1(n15899), .B2(
        P1_REIP_REG_14__SCAN_IN), .ZN(n15867) );
  AOI22_X1 U19039 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15865), .B1(
        n15864), .B2(n15863), .ZN(n15866) );
  OAI211_X1 U19040 ( .C1(n15868), .C2(n20138), .A(n15867), .B(n15866), .ZN(
        P1_U3017) );
  INV_X1 U19041 ( .A(n15869), .ZN(n15875) );
  AOI22_X1 U19042 ( .A1(n15870), .A2(n15932), .B1(n15899), .B2(
        P1_REIP_REG_13__SCAN_IN), .ZN(n15871) );
  OAI21_X1 U19043 ( .B1(n15873), .B2(n15872), .A(n15871), .ZN(n15874) );
  AOI21_X1 U19044 ( .B1(n15875), .B2(n15933), .A(n15874), .ZN(n15877) );
  OAI211_X1 U19045 ( .C1(n15879), .C2(n15878), .A(n15877), .B(n15876), .ZN(
        P1_U3018) );
  INV_X1 U19046 ( .A(n15887), .ZN(n15880) );
  NOR2_X1 U19047 ( .A1(n15906), .A2(n15880), .ZN(n15891) );
  NOR2_X1 U19048 ( .A1(n15883), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15898) );
  OAI21_X1 U19049 ( .B1(n15883), .B2(n15882), .A(n15881), .ZN(n15884) );
  OAI211_X1 U19050 ( .C1(n15887), .C2(n15886), .A(n15885), .B(n15884), .ZN(
        n15902) );
  AOI21_X1 U19051 ( .B1(n15888), .B2(n15898), .A(n15902), .ZN(n15889) );
  INV_X1 U19052 ( .A(n15889), .ZN(n15890) );
  MUX2_X1 U19053 ( .A(n15891), .B(n15890), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n15895) );
  INV_X1 U19054 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21154) );
  NAND2_X1 U19055 ( .A1(n15932), .A2(n15892), .ZN(n15893) );
  OAI21_X1 U19056 ( .B1(n21154), .B2(n20135), .A(n15893), .ZN(n15894) );
  NOR2_X1 U19057 ( .A1(n15895), .A2(n15894), .ZN(n15896) );
  OAI21_X1 U19058 ( .B1(n15897), .B2(n20138), .A(n15896), .ZN(P1_U3019) );
  INV_X1 U19059 ( .A(n15898), .ZN(n15905) );
  AOI22_X1 U19060 ( .A1(n15932), .A2(n15900), .B1(n15899), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15904) );
  AOI22_X1 U19061 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n15902), .B1(
        n15933), .B2(n15901), .ZN(n15903) );
  OAI211_X1 U19062 ( .C1(n15906), .C2(n15905), .A(n15904), .B(n15903), .ZN(
        P1_U3020) );
  AOI22_X1 U19063 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15907), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n15763), .ZN(n15915) );
  INV_X1 U19064 ( .A(n15908), .ZN(n15909) );
  AOI21_X1 U19065 ( .B1(n15932), .B2(n15910), .A(n15909), .ZN(n15914) );
  AOI22_X1 U19066 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n15912), .B1(
        n15933), .B2(n15911), .ZN(n15913) );
  OAI211_X1 U19067 ( .C1(n15916), .C2(n15915), .A(n15914), .B(n15913), .ZN(
        P1_U3021) );
  AOI21_X1 U19068 ( .B1(n15932), .B2(n15918), .A(n15917), .ZN(n15926) );
  AOI22_X1 U19069 ( .A1(n15920), .A2(n15933), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15919), .ZN(n15925) );
  OAI221_X1 U19070 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n15923), .C2(n15922), .A(
        n15921), .ZN(n15924) );
  NAND3_X1 U19071 ( .A1(n15926), .A2(n15925), .A3(n15924), .ZN(P1_U3023) );
  NOR2_X1 U19072 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15927), .ZN(
        n15938) );
  OAI21_X1 U19073 ( .B1(n15930), .B2(n15929), .A(n15928), .ZN(n15931) );
  INV_X1 U19074 ( .A(n15931), .ZN(n20072) );
  AOI22_X1 U19075 ( .A1(n15934), .A2(n15933), .B1(n15932), .B2(n20072), .ZN(
        n15937) );
  NAND2_X1 U19076 ( .A1(n15935), .A2(P1_REIP_REG_6__SCAN_IN), .ZN(n15936) );
  OAI211_X1 U19077 ( .C1(n15939), .C2(n15938), .A(n15937), .B(n15936), .ZN(
        P1_U3025) );
  INV_X1 U19078 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15945) );
  INV_X1 U19079 ( .A(n15940), .ZN(n15943) );
  NAND4_X1 U19080 ( .A1(n15943), .A2(n15942), .A3(n15941), .A4(n20045), .ZN(
        n15944) );
  OAI21_X1 U19081 ( .B1(n20790), .B2(n15945), .A(n15944), .ZN(P1_U3468) );
  NAND4_X1 U19082 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20721), .A4(n20800), .ZN(n15946) );
  NAND2_X1 U19083 ( .A1(n15947), .A2(n15946), .ZN(n20719) );
  OAI21_X1 U19084 ( .B1(n15949), .B2(n20719), .A(n15948), .ZN(n15950) );
  OAI221_X1 U19085 ( .B1(n15951), .B2(n20537), .C1(n15951), .C2(n20800), .A(
        n15950), .ZN(n15952) );
  AOI221_X1 U19086 ( .B1(n15953), .B2(n20717), .C1(n20718), .C2(n20717), .A(
        n15952), .ZN(P1_U3162) );
  NOR2_X1 U19087 ( .A1(n15953), .A2(n20718), .ZN(n15955) );
  OAI22_X1 U19088 ( .A1(n20537), .A2(n15955), .B1(n15954), .B2(n20718), .ZN(
        P1_U3466) );
  INV_X1 U19089 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n15958) );
  INV_X1 U19090 ( .A(n15956), .ZN(n15957) );
  INV_X1 U19091 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16059) );
  OAI222_X1 U19092 ( .A1(n19067), .A2(n15958), .B1(n19072), .B2(n15957), .C1(
        n16059), .C2(n19065), .ZN(n15959) );
  AOI21_X1 U19093 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19081), .A(
        n15959), .ZN(n15971) );
  INV_X1 U19094 ( .A(n15960), .ZN(n15972) );
  INV_X1 U19095 ( .A(n15961), .ZN(n16017) );
  OAI21_X1 U19096 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15963), .A(
        n15962), .ZN(n16092) );
  INV_X1 U19097 ( .A(n16092), .ZN(n16042) );
  NOR2_X1 U19098 ( .A1(n10004), .A2(n15964), .ZN(n16050) );
  NOR2_X1 U19099 ( .A1(n16050), .A2(n16051), .ZN(n16049) );
  NOR2_X1 U19100 ( .A1(n16049), .A2(n10004), .ZN(n16041) );
  NOR2_X1 U19101 ( .A1(n16017), .A2(n16016), .ZN(n16015) );
  NOR2_X1 U19102 ( .A1(n10004), .A2(n16015), .ZN(n16010) );
  OR2_X1 U19103 ( .A1(n9914), .A2(n15996), .ZN(n15966) );
  OAI21_X1 U19104 ( .B1(n16010), .B2(n15966), .A(n9918), .ZN(n15994) );
  NOR2_X1 U19105 ( .A1(n10004), .A2(n15994), .ZN(n15985) );
  AND2_X1 U19106 ( .A1(n15967), .A2(n15984), .ZN(n15968) );
  INV_X1 U19107 ( .A(n19058), .ZN(n19834) );
  NOR2_X1 U19108 ( .A1(n10004), .A2(n19834), .ZN(n19079) );
  AOI22_X1 U19109 ( .A1(n15974), .A2(n19079), .B1(n19069), .B2(n15969), .ZN(
        n15970) );
  OAI211_X1 U19110 ( .C1(n16060), .C2(n19046), .A(n15971), .B(n15970), .ZN(
        P2_U2824) );
  AOI22_X1 U19111 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19053), .ZN(n15976) );
  NAND2_X1 U19112 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19081), .ZN(
        n15975) );
  OAI211_X1 U19113 ( .C1(n19072), .C2(n15977), .A(n15976), .B(n15975), .ZN(
        n15978) );
  AOI21_X1 U19114 ( .B1(n15985), .B2(n15984), .A(n19834), .ZN(n15991) );
  AOI22_X1 U19115 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19047), .B1(n15986), 
        .B2(n18991), .ZN(n15988) );
  AOI22_X1 U19116 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19053), .ZN(n15987) );
  OAI211_X1 U19117 ( .C1(n15989), .C2(n19046), .A(n15988), .B(n15987), .ZN(
        n15990) );
  AOI21_X1 U19118 ( .B1(n10227), .B2(n15991), .A(n15990), .ZN(n15992) );
  OAI21_X1 U19119 ( .B1(n15993), .B2(n19055), .A(n15992), .ZN(P2_U2826) );
  NOR2_X1 U19120 ( .A1(n9914), .A2(n16010), .ZN(n16009) );
  NOR2_X1 U19121 ( .A1(n10004), .A2(n16009), .ZN(n15995) );
  AOI211_X1 U19122 ( .C1(n15996), .C2(n15995), .A(n15994), .B(n19834), .ZN(
        n16001) );
  AOI22_X1 U19123 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19053), .ZN(n15998) );
  NAND2_X1 U19124 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19081), .ZN(
        n15997) );
  OAI211_X1 U19125 ( .C1(n19072), .C2(n15999), .A(n15998), .B(n15997), .ZN(
        n16000) );
  AOI211_X1 U19126 ( .C1(n19069), .C2(n16002), .A(n16001), .B(n16000), .ZN(
        n16003) );
  OAI21_X1 U19127 ( .B1(n16004), .B2(n19046), .A(n16003), .ZN(P2_U2827) );
  AOI22_X1 U19128 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19053), .ZN(n16007) );
  AOI22_X1 U19129 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19081), .B1(
        n16005), .B2(n18991), .ZN(n16006) );
  OAI211_X1 U19130 ( .C1(n16008), .C2(n19055), .A(n16007), .B(n16006), .ZN(
        n16012) );
  AOI211_X1 U19131 ( .C1(n9914), .C2(n16010), .A(n16009), .B(n19834), .ZN(
        n16011) );
  NOR2_X1 U19132 ( .A1(n16012), .A2(n16011), .ZN(n16013) );
  OAI21_X1 U19133 ( .B1(n16014), .B2(n19046), .A(n16013), .ZN(P2_U2828) );
  AOI211_X1 U19134 ( .C1(n16017), .C2(n16016), .A(n16015), .B(n19834), .ZN(
        n16023) );
  AOI22_X1 U19135 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19053), .ZN(n16020) );
  AOI22_X1 U19136 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19081), .B1(
        n16018), .B2(n18991), .ZN(n16019) );
  OAI211_X1 U19137 ( .C1(n16021), .C2(n19046), .A(n16020), .B(n16019), .ZN(
        n16022) );
  AOI211_X1 U19138 ( .C1(n19069), .C2(n16024), .A(n16023), .B(n16022), .ZN(
        n16025) );
  INV_X1 U19139 ( .A(n16025), .ZN(P2_U2829) );
  AOI211_X1 U19140 ( .C1(n16027), .C2(n16026), .A(n10007), .B(n19834), .ZN(
        n16035) );
  AOI22_X1 U19141 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19053), .ZN(n16032) );
  OAI22_X1 U19142 ( .A1(n16029), .A2(n19072), .B1(n16028), .B2(n19049), .ZN(
        n16030) );
  INV_X1 U19143 ( .A(n16030), .ZN(n16031) );
  OAI211_X1 U19144 ( .C1(n16033), .C2(n19055), .A(n16032), .B(n16031), .ZN(
        n16034) );
  AOI211_X1 U19145 ( .C1(n19075), .C2(n16036), .A(n16035), .B(n16034), .ZN(
        n16037) );
  INV_X1 U19146 ( .A(n16037), .ZN(P2_U2830) );
  INV_X1 U19147 ( .A(n16038), .ZN(n16088) );
  AOI22_X1 U19148 ( .A1(n16088), .A2(n19075), .B1(n16039), .B2(n19069), .ZN(
        n16048) );
  AOI211_X1 U19149 ( .C1(n16042), .C2(n16041), .A(n16040), .B(n19834), .ZN(
        n16046) );
  AOI22_X1 U19150 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19053), .ZN(n16043) );
  OAI21_X1 U19151 ( .B1(n16044), .B2(n19072), .A(n16043), .ZN(n16045) );
  AOI211_X1 U19152 ( .C1(n19081), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16046), .B(n16045), .ZN(n16047) );
  NAND2_X1 U19153 ( .A1(n16048), .A2(n16047), .ZN(P2_U2831) );
  AOI211_X1 U19154 ( .C1(n16051), .C2(n16050), .A(n16049), .B(n19834), .ZN(
        n16057) );
  AOI22_X1 U19155 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19053), .ZN(n16054) );
  AOI22_X1 U19156 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n19081), .B1(
        n16052), .B2(n18991), .ZN(n16053) );
  OAI211_X1 U19157 ( .C1(n16055), .C2(n19055), .A(n16054), .B(n16053), .ZN(
        n16056) );
  AOI211_X1 U19158 ( .C1(n19075), .C2(n16061), .A(n16057), .B(n16056), .ZN(
        n16058) );
  INV_X1 U19159 ( .A(n16058), .ZN(P2_U2832) );
  AOI22_X1 U19160 ( .A1(n19121), .A2(n16060), .B1(n16059), .B2(n19116), .ZN(
        P2_U2856) );
  AOI22_X1 U19161 ( .A1(n16062), .A2(n19107), .B1(n19121), .B2(n16061), .ZN(
        n16063) );
  OAI21_X1 U19162 ( .B1(n19121), .B2(n12558), .A(n16063), .ZN(P2_U2864) );
  INV_X1 U19163 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n16067) );
  AOI21_X1 U19164 ( .B1(n16065), .B2(n14789), .A(n16064), .ZN(n16074) );
  AOI22_X1 U19165 ( .A1(n16074), .A2(n19107), .B1(n19121), .B2(n16097), .ZN(
        n16066) );
  OAI21_X1 U19166 ( .B1(n19121), .B2(n16067), .A(n16066), .ZN(P2_U2865) );
  AOI21_X1 U19167 ( .B1(n16069), .B2(n14797), .A(n16068), .ZN(n16078) );
  AOI22_X1 U19168 ( .A1(n16078), .A2(n19107), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19116), .ZN(n16070) );
  OAI21_X1 U19169 ( .B1(n19116), .B2(n18865), .A(n16070), .ZN(P2_U2867) );
  AOI21_X1 U19170 ( .B1(n16071), .B2(n14000), .A(n9917), .ZN(n16083) );
  AOI22_X1 U19171 ( .A1(n16083), .A2(n19107), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n19116), .ZN(n16072) );
  OAI21_X1 U19172 ( .B1(n19116), .B2(n18888), .A(n16072), .ZN(P2_U2869) );
  AOI22_X1 U19173 ( .A1(n19125), .A2(n19161), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19186), .ZN(n16077) );
  AOI22_X1 U19174 ( .A1(n19127), .A2(BUF1_REG_22__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16076) );
  AOI22_X1 U19175 ( .A1(n16074), .A2(n19176), .B1(n19187), .B2(n16073), .ZN(
        n16075) );
  NAND3_X1 U19176 ( .A1(n16077), .A2(n16076), .A3(n16075), .ZN(P2_U2897) );
  AOI22_X1 U19177 ( .A1(n19125), .A2(n19173), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19186), .ZN(n16081) );
  AOI22_X1 U19178 ( .A1(n19127), .A2(BUF1_REG_20__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16080) );
  AOI22_X1 U19179 ( .A1(n16078), .A2(n19176), .B1(n19187), .B2(n9883), .ZN(
        n16079) );
  NAND3_X1 U19180 ( .A1(n16081), .A2(n16080), .A3(n16079), .ZN(P2_U2899) );
  AOI22_X1 U19181 ( .A1(n19125), .A2(n16082), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19186), .ZN(n16086) );
  AOI22_X1 U19182 ( .A1(n19127), .A2(BUF1_REG_18__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16085) );
  AOI22_X1 U19183 ( .A1(n16083), .A2(n19176), .B1(n19187), .B2(n18885), .ZN(
        n16084) );
  NAND3_X1 U19184 ( .A1(n16086), .A2(n16085), .A3(n16084), .ZN(P2_U2901) );
  AOI22_X1 U19185 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n12763), .ZN(n16091) );
  AOI222_X1 U19186 ( .A1(n16089), .A2(n19240), .B1(n19250), .B2(n16088), .C1(
        n19242), .C2(n16087), .ZN(n16090) );
  OAI211_X1 U19187 ( .C1(n19247), .C2(n16092), .A(n16091), .B(n16090), .ZN(
        P2_U2990) );
  AOI22_X1 U19188 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n12763), .ZN(n16099) );
  NOR3_X1 U19189 ( .A1(n16093), .A2(n9838), .A3(n16172), .ZN(n16096) );
  NOR2_X1 U19190 ( .A1(n16094), .A2(n16173), .ZN(n16095) );
  AOI211_X1 U19191 ( .C1(n19250), .C2(n16097), .A(n16096), .B(n16095), .ZN(
        n16098) );
  OAI211_X1 U19192 ( .C1(n19247), .C2(n16100), .A(n16099), .B(n16098), .ZN(
        P2_U2992) );
  AOI22_X1 U19193 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n12763), .ZN(n16117) );
  OR2_X1 U19194 ( .A1(n9877), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16101) );
  AND2_X1 U19195 ( .A1(n15035), .A2(n16101), .ZN(n16203) );
  INV_X1 U19196 ( .A(n16102), .ZN(n16108) );
  INV_X1 U19197 ( .A(n16103), .ZN(n16106) );
  INV_X1 U19198 ( .A(n16104), .ZN(n16105) );
  NAND2_X1 U19199 ( .A1(n16106), .A2(n16105), .ZN(n16107) );
  NAND2_X1 U19200 ( .A1(n16108), .A2(n16107), .ZN(n19096) );
  NOR2_X1 U19201 ( .A1(n19096), .A2(n15339), .ZN(n16109) );
  AOI21_X1 U19202 ( .B1(n16203), .B2(n19242), .A(n16109), .ZN(n16115) );
  NAND2_X1 U19203 ( .A1(n16111), .A2(n16110), .ZN(n16112) );
  XNOR2_X1 U19204 ( .A(n16113), .B(n16112), .ZN(n16206) );
  NAND2_X1 U19205 ( .A1(n16206), .A2(n19240), .ZN(n16114) );
  AND2_X1 U19206 ( .A1(n16115), .A2(n16114), .ZN(n16116) );
  OAI211_X1 U19207 ( .C1(n19247), .C2(n18922), .A(n16117), .B(n16116), .ZN(
        P2_U3000) );
  AOI22_X1 U19208 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n12763), .B1(n16170), 
        .B2(n18934), .ZN(n16122) );
  OAI22_X1 U19209 ( .A1(n16119), .A2(n16172), .B1(n16118), .B2(n16173), .ZN(
        n16120) );
  AOI21_X1 U19210 ( .B1(n19250), .B2(n18935), .A(n16120), .ZN(n16121) );
  OAI211_X1 U19211 ( .C1(n16179), .C2(n18930), .A(n16122), .B(n16121), .ZN(
        P2_U3001) );
  AOI22_X1 U19212 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n12763), .ZN(n16129) );
  NOR3_X1 U19213 ( .A1(n16124), .A2(n16123), .A3(n16172), .ZN(n16127) );
  OAI22_X1 U19214 ( .A1(n16125), .A2(n16173), .B1(n15339), .B2(n19101), .ZN(
        n16126) );
  NOR2_X1 U19215 ( .A1(n16127), .A2(n16126), .ZN(n16128) );
  OAI211_X1 U19216 ( .C1(n19247), .C2(n18938), .A(n16129), .B(n16128), .ZN(
        P2_U3002) );
  AOI22_X1 U19217 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19016), .B1(n16170), 
        .B2(n18958), .ZN(n16134) );
  OAI22_X1 U19218 ( .A1(n16131), .A2(n16172), .B1(n16130), .B2(n16173), .ZN(
        n16132) );
  AOI21_X1 U19219 ( .B1(n19250), .B2(n18947), .A(n16132), .ZN(n16133) );
  OAI211_X1 U19220 ( .C1(n16179), .C2(n18955), .A(n16134), .B(n16133), .ZN(
        P2_U3003) );
  AOI22_X1 U19221 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n12763), .ZN(n16147) );
  NOR2_X1 U19222 ( .A1(n16136), .A2(n16135), .ZN(n16140) );
  NAND2_X1 U19223 ( .A1(n16138), .A2(n16137), .ZN(n16139) );
  XNOR2_X1 U19224 ( .A(n16140), .B(n16139), .ZN(n16222) );
  INV_X1 U19225 ( .A(n16222), .ZN(n16145) );
  NOR2_X1 U19226 ( .A1(n13357), .A2(n16141), .ZN(n16142) );
  NOR2_X1 U19227 ( .A1(n13394), .A2(n16142), .ZN(n19104) );
  AOI21_X1 U19228 ( .B1(n12506), .B2(n16144), .A(n16143), .ZN(n16219) );
  AOI222_X1 U19229 ( .A1(n16145), .A2(n19240), .B1(n19250), .B2(n19104), .C1(
        n19242), .C2(n16219), .ZN(n16146) );
  OAI211_X1 U19230 ( .C1(n19247), .C2(n18965), .A(n16147), .B(n16146), .ZN(
        P2_U3004) );
  AOI22_X1 U19231 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n12763), .ZN(n16162) );
  INV_X1 U19232 ( .A(n13356), .ZN(n16148) );
  OAI21_X1 U19233 ( .B1(n16150), .B2(n16149), .A(n16148), .ZN(n19115) );
  NAND2_X1 U19234 ( .A1(n16152), .A2(n16151), .ZN(n16156) );
  NAND2_X1 U19235 ( .A1(n16154), .A2(n16153), .ZN(n16155) );
  XOR2_X1 U19236 ( .A(n16156), .B(n16155), .Z(n16240) );
  OAI21_X1 U19237 ( .B1(n16159), .B2(n16158), .A(n16157), .ZN(n16235) );
  OAI222_X1 U19238 ( .A1(n19115), .A2(n15339), .B1(n16173), .B2(n16240), .C1(
        n16172), .C2(n16235), .ZN(n16160) );
  INV_X1 U19239 ( .A(n16160), .ZN(n16161) );
  OAI211_X1 U19240 ( .C1(n19247), .C2(n18986), .A(n16162), .B(n16161), .ZN(
        P2_U3006) );
  AOI22_X1 U19241 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n12763), .ZN(n16169) );
  OR2_X1 U19242 ( .A1(n16163), .A2(n16172), .ZN(n16165) );
  NAND2_X1 U19243 ( .A1(n19009), .A2(n19250), .ZN(n16164) );
  OAI211_X1 U19244 ( .C1(n16166), .C2(n16173), .A(n16165), .B(n16164), .ZN(
        n16167) );
  INV_X1 U19245 ( .A(n16167), .ZN(n16168) );
  OAI211_X1 U19246 ( .C1(n19247), .C2(n19007), .A(n16169), .B(n16168), .ZN(
        P2_U3008) );
  AOI22_X1 U19247 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19016), .B1(n16170), 
        .B2(n19019), .ZN(n16177) );
  OAI22_X1 U19248 ( .A1(n16174), .A2(n16173), .B1(n16172), .B2(n16171), .ZN(
        n16175) );
  AOI21_X1 U19249 ( .B1(n19250), .B2(n19020), .A(n16175), .ZN(n16176) );
  OAI211_X1 U19250 ( .C1(n16179), .C2(n16178), .A(n16177), .B(n16176), .ZN(
        P2_U3009) );
  INV_X1 U19251 ( .A(n16180), .ZN(n16183) );
  INV_X1 U19252 ( .A(n16181), .ZN(n16182) );
  NAND2_X1 U19253 ( .A1(n16183), .A2(n16182), .ZN(n16184) );
  NAND2_X1 U19254 ( .A1(n9888), .A2(n16184), .ZN(n19137) );
  OAI21_X1 U19255 ( .B1(n16215), .B2(n19137), .A(n16185), .ZN(n16186) );
  AOI221_X1 U19256 ( .B1(n16189), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), 
        .C1(n16188), .C2(n16187), .A(n16186), .ZN(n16193) );
  INV_X1 U19257 ( .A(n16190), .ZN(n16191) );
  AOI22_X1 U19258 ( .A1(n16191), .A2(n19262), .B1(n19255), .B2(n18916), .ZN(
        n16192) );
  OAI211_X1 U19259 ( .C1(n16194), .C2(n16246), .A(n16193), .B(n16192), .ZN(
        P2_U3031) );
  OAI21_X1 U19260 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16196), .A(
        n16195), .ZN(n16200) );
  NOR2_X1 U19261 ( .A1(n16197), .A2(n15239), .ZN(n16198) );
  NOR2_X1 U19262 ( .A1(n16198), .A2(n16180), .ZN(n19138) );
  AOI22_X1 U19263 ( .A1(n19257), .A2(n19138), .B1(n19016), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n16199) );
  OAI21_X1 U19264 ( .B1(n16201), .B2(n16200), .A(n16199), .ZN(n16202) );
  INV_X1 U19265 ( .A(n16202), .ZN(n16208) );
  INV_X1 U19266 ( .A(n16203), .ZN(n16204) );
  OAI22_X1 U19267 ( .A1(n16204), .A2(n16264), .B1(n16253), .B2(n19096), .ZN(
        n16205) );
  AOI21_X1 U19268 ( .B1(n19263), .B2(n16206), .A(n16205), .ZN(n16207) );
  OAI211_X1 U19269 ( .C1(n16210), .C2(n16209), .A(n16208), .B(n16207), .ZN(
        P2_U3032) );
  NOR2_X1 U19270 ( .A1(n12671), .A2(n16232), .ZN(n16217) );
  INV_X1 U19271 ( .A(n16211), .ZN(n16212) );
  XNOR2_X1 U19272 ( .A(n16213), .B(n16212), .ZN(n19152) );
  OAI22_X1 U19273 ( .A1(n16215), .A2(n19152), .B1(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16214), .ZN(n16216) );
  AOI211_X1 U19274 ( .C1(n16218), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16217), .B(n16216), .ZN(n16221) );
  AOI22_X1 U19275 ( .A1(n16219), .A2(n19262), .B1(n19255), .B2(n19104), .ZN(
        n16220) );
  OAI211_X1 U19276 ( .C1(n16222), .C2(n16246), .A(n16221), .B(n16220), .ZN(
        P2_U3036) );
  NAND2_X1 U19277 ( .A1(n16224), .A2(n16223), .ZN(n16228) );
  AOI222_X1 U19278 ( .A1(n16228), .A2(n16227), .B1(n16228), .B2(n16226), .C1(
        n16227), .C2(n16225), .ZN(n16234) );
  AOI21_X1 U19279 ( .B1(n16230), .B2(n16229), .A(n13933), .ZN(n19155) );
  NAND2_X1 U19280 ( .A1(n19257), .A2(n19155), .ZN(n16231) );
  OAI21_X1 U19281 ( .B1(n12644), .B2(n16232), .A(n16231), .ZN(n16233) );
  NOR2_X1 U19282 ( .A1(n16234), .A2(n16233), .ZN(n16239) );
  INV_X1 U19283 ( .A(n16235), .ZN(n16237) );
  INV_X1 U19284 ( .A(n19115), .ZN(n16236) );
  AOI22_X1 U19285 ( .A1(n16237), .A2(n19262), .B1(n19255), .B2(n16236), .ZN(
        n16238) );
  OAI211_X1 U19286 ( .C1(n16240), .C2(n16246), .A(n16239), .B(n16238), .ZN(
        P2_U3038) );
  INV_X1 U19287 ( .A(n19167), .ZN(n19931) );
  AOI22_X1 U19288 ( .A1(n16242), .A2(n16241), .B1(n19257), .B2(n19931), .ZN(
        n16243) );
  OAI21_X1 U19289 ( .B1(n16244), .B2(n16253), .A(n16243), .ZN(n16249) );
  OAI22_X1 U19290 ( .A1(n16247), .A2(n16246), .B1(n16264), .B2(n16245), .ZN(
        n16248) );
  AOI211_X1 U19291 ( .C1(P2_REIP_REG_3__SCAN_IN), .C2(n12763), .A(n16249), .B(
        n16248), .ZN(n16250) );
  OAI21_X1 U19292 ( .B1(n16251), .B2(n13419), .A(n16250), .ZN(P2_U3043) );
  OAI22_X1 U19293 ( .A1(n16254), .A2(n12056), .B1(n16253), .B2(n16252), .ZN(
        n16255) );
  INV_X1 U19294 ( .A(n16255), .ZN(n16260) );
  AOI22_X1 U19295 ( .A1(n19263), .A2(n16256), .B1(n19257), .B2(n19070), .ZN(
        n16259) );
  NAND2_X1 U19296 ( .A1(n16257), .A2(n12056), .ZN(n16258) );
  AND3_X1 U19297 ( .A1(n16260), .A2(n16259), .A3(n16258), .ZN(n16262) );
  OAI211_X1 U19298 ( .C1(n16264), .C2(n16263), .A(n16262), .B(n16261), .ZN(
        P2_U3046) );
  NOR2_X1 U19299 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13470), .ZN(n19832) );
  AOI21_X1 U19300 ( .B1(n19980), .B2(n19832), .A(n16265), .ZN(n16323) );
  INV_X1 U19301 ( .A(n12423), .ZN(n16275) );
  INV_X1 U19302 ( .A(n16266), .ZN(n16268) );
  AOI22_X1 U19303 ( .A1(n16272), .A2(n16269), .B1(n16268), .B2(n16267), .ZN(
        n16270) );
  OAI21_X1 U19304 ( .B1(n16272), .B2(n16271), .A(n16270), .ZN(n19966) );
  AOI211_X1 U19305 ( .C1(n16275), .C2(n16274), .A(n16273), .B(n19966), .ZN(
        n16310) );
  NAND2_X1 U19306 ( .A1(n16277), .A2(n16276), .ZN(n16286) );
  INV_X1 U19307 ( .A(n16278), .ZN(n16281) );
  OAI22_X1 U19308 ( .A1(n16281), .A2(n16286), .B1(n16280), .B2(n16279), .ZN(
        n16285) );
  NOR2_X1 U19309 ( .A1(n16283), .A2(n16282), .ZN(n16284) );
  AOI211_X1 U19310 ( .C1(n16287), .C2(n16286), .A(n16285), .B(n16284), .ZN(
        n19915) );
  INV_X1 U19311 ( .A(n16293), .ZN(n16289) );
  NOR2_X1 U19312 ( .A1(n16289), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16288) );
  AOI21_X1 U19313 ( .B1(n19915), .B2(n16289), .A(n16288), .ZN(n16298) );
  MUX2_X1 U19314 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n16297), .S(
        n16289), .Z(n16300) );
  AOI22_X1 U19315 ( .A1(n16298), .A2(n16300), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n16293), .ZN(n16309) );
  NAND2_X1 U19316 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n16290), .ZN(
        n16291) );
  OAI21_X1 U19317 ( .B1(n16292), .B2(n16291), .A(n19949), .ZN(n16295) );
  NAND2_X1 U19318 ( .A1(n16292), .A2(n16291), .ZN(n16294) );
  AOI21_X1 U19319 ( .B1(n16295), .B2(n16294), .A(n16293), .ZN(n16296) );
  OAI21_X1 U19320 ( .B1(n19933), .B2(n16297), .A(n16296), .ZN(n16301) );
  INV_X1 U19321 ( .A(n16298), .ZN(n16299) );
  AOI211_X1 U19322 ( .C1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n16301), .A(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16299), .ZN(n16305) );
  INV_X1 U19323 ( .A(n16300), .ZN(n16302) );
  OAI22_X1 U19324 ( .A1(n16302), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16301), .ZN(n16304) );
  OAI21_X1 U19325 ( .B1(n16305), .B2(n16304), .A(n16303), .ZN(n16308) );
  OAI21_X1 U19326 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n16306), .ZN(n16307) );
  NAND4_X1 U19327 ( .A1(n16310), .A2(n16309), .A3(n16308), .A4(n16307), .ZN(
        n16321) );
  AOI21_X1 U19328 ( .B1(n13470), .B2(n19916), .A(n19982), .ZN(n16319) );
  OAI21_X1 U19329 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(n16321), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n16317) );
  NAND2_X1 U19330 ( .A1(n16312), .A2(n16311), .ZN(n16314) );
  OAI211_X1 U19331 ( .C1(n12413), .C2(n16314), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n16313), .ZN(n16315) );
  INV_X1 U19332 ( .A(n16315), .ZN(n16316) );
  NOR2_X1 U19333 ( .A1(n19838), .A2(n16325), .ZN(n16318) );
  OAI22_X1 U19334 ( .A1(n16319), .A2(n16318), .B1(n13470), .B2(n16325), .ZN(
        n16320) );
  AOI21_X1 U19335 ( .B1(n19829), .B2(n16321), .A(n16320), .ZN(n16322) );
  OAI211_X1 U19336 ( .C1(n19962), .C2(n16324), .A(n16323), .B(n16322), .ZN(
        P2_U3176) );
  OAI221_X1 U19337 ( .B1(n19971), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19971), 
        .C2(n16325), .A(n16324), .ZN(P2_U3593) );
  NAND2_X1 U19338 ( .A1(n17818), .A2(n16326), .ZN(n16340) );
  NAND2_X1 U19339 ( .A1(n17528), .A2(n16327), .ZN(n16341) );
  NAND3_X1 U19340 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n17860), .ZN(n17835) );
  NAND2_X1 U19341 ( .A1(n17895), .A2(n17616), .ZN(n17557) );
  NOR2_X1 U19342 ( .A1(n17835), .A2(n17557), .ZN(n17503) );
  NAND2_X1 U19343 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17503), .ZN(
        n17492) );
  NOR3_X1 U19344 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16328), .A3(
        n17492), .ZN(n16334) );
  XOR2_X1 U19345 ( .A(n9924), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Z(n16516) );
  AOI21_X1 U19346 ( .B1(n17685), .B2(n16516), .A(n16329), .ZN(n16330) );
  OAI221_X1 U19347 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16332), .C1(
        n10053), .C2(n16331), .A(n16330), .ZN(n16333) );
  OAI221_X1 U19348 ( .B1(n16336), .B2(n16340), .C1(n16336), .C2(n16341), .A(
        n16335), .ZN(P3_U2800) );
  AOI22_X1 U19349 ( .A1(n16339), .A2(n16338), .B1(
        P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16337), .ZN(n16351) );
  AOI21_X1 U19350 ( .B1(n16342), .B2(n16364), .A(n16340), .ZN(n16345) );
  AOI21_X1 U19351 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n16344) );
  AOI211_X1 U19352 ( .C1(n16346), .C2(n17739), .A(n16345), .B(n16344), .ZN(
        n16350) );
  NAND2_X1 U19353 ( .A1(n9821), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16349) );
  AOI21_X1 U19354 ( .B1(n10051), .B2(n16493), .A(n9924), .ZN(n16525) );
  OAI21_X1 U19355 ( .B1(n17685), .B2(n16347), .A(n16525), .ZN(n16348) );
  NAND4_X1 U19356 ( .A1(n16351), .A2(n16350), .A3(n16349), .A4(n16348), .ZN(
        P3_U2801) );
  AOI22_X1 U19357 ( .A1(n17734), .A2(n17472), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n17702), .ZN(n17470) );
  NAND2_X1 U19358 ( .A1(n9811), .A2(n17470), .ZN(n16371) );
  NAND2_X1 U19359 ( .A1(n17734), .A2(n18136), .ZN(n16360) );
  NOR2_X1 U19360 ( .A1(n16353), .A2(n16352), .ZN(n16358) );
  NAND2_X1 U19361 ( .A1(n18113), .A2(n18114), .ZN(n17935) );
  INV_X1 U19362 ( .A(n18017), .ZN(n18581) );
  NOR2_X1 U19363 ( .A1(n16354), .A2(n18588), .ZN(n18022) );
  AOI22_X1 U19364 ( .A1(n18581), .A2(n18018), .B1(n17997), .B2(n18022), .ZN(
        n17938) );
  OAI21_X1 U19365 ( .B1(n16355), .B2(n17935), .A(n17938), .ZN(n16357) );
  AOI21_X1 U19366 ( .B1(n16358), .B2(n16357), .A(n16356), .ZN(n17901) );
  NOR2_X1 U19367 ( .A1(n17901), .A2(n18127), .ZN(n17910) );
  NAND2_X1 U19368 ( .A1(n17884), .A2(n17910), .ZN(n17870) );
  OAI22_X1 U19369 ( .A1(n17469), .A2(n16360), .B1(n16359), .B2(n17870), .ZN(
        n16361) );
  AOI22_X1 U19370 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n18042), .B1(n17472), 
        .B2(n16361), .ZN(n16370) );
  INV_X1 U19371 ( .A(n18022), .ZN(n17996) );
  AOI21_X1 U19372 ( .B1(n18581), .B2(n16364), .A(n16363), .ZN(n16365) );
  OAI211_X1 U19373 ( .C1(n16367), .C2(n17996), .A(n16366), .B(n16365), .ZN(
        n16368) );
  NAND3_X1 U19374 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18036), .A3(
        n16368), .ZN(n16369) );
  OAI211_X1 U19375 ( .C1(n17483), .C2(n16371), .A(n16370), .B(n16369), .ZN(
        P3_U2834) );
  NOR3_X1 U19376 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16373) );
  NOR4_X1 U19377 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16372) );
  NAND4_X1 U19378 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16373), .A3(n16372), .A4(
        U215), .ZN(U213) );
  INV_X1 U19379 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16463) );
  INV_X2 U19380 ( .A(U214), .ZN(n16423) );
  INV_X1 U19381 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16462) );
  OAI222_X1 U19382 ( .A1(U212), .A2(n16463), .B1(n16426), .B2(n16375), .C1(
        U214), .C2(n16462), .ZN(U216) );
  INV_X1 U19383 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20181) );
  INV_X2 U19384 ( .A(U212), .ZN(n16424) );
  AOI22_X1 U19385 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16423), .ZN(n16376) );
  OAI21_X1 U19386 ( .B1(n20181), .B2(n16426), .A(n16376), .ZN(U217) );
  INV_X1 U19387 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20174) );
  AOI22_X1 U19388 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n16423), .ZN(n16377) );
  OAI21_X1 U19389 ( .B1(n20174), .B2(n16426), .A(n16377), .ZN(U218) );
  AOI22_X1 U19390 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16423), .ZN(n16378) );
  OAI21_X1 U19391 ( .B1(n16379), .B2(n16426), .A(n16378), .ZN(U219) );
  INV_X1 U19392 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20168) );
  AOI22_X1 U19393 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16423), .ZN(n16380) );
  OAI21_X1 U19394 ( .B1(n20168), .B2(n16426), .A(n16380), .ZN(U220) );
  AOI22_X1 U19395 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16423), .ZN(n16381) );
  OAI21_X1 U19396 ( .B1(n20161), .B2(n16426), .A(n16381), .ZN(U221) );
  AOI22_X1 U19397 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n16423), .ZN(n16382) );
  OAI21_X1 U19398 ( .B1(n14844), .B2(n16426), .A(n16382), .ZN(U222) );
  INV_X1 U19399 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20150) );
  AOI22_X1 U19400 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16423), .ZN(n16383) );
  OAI21_X1 U19401 ( .B1(n20150), .B2(n16426), .A(n16383), .ZN(U223) );
  AOI22_X1 U19402 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16423), .ZN(n16384) );
  OAI21_X1 U19403 ( .B1(n16385), .B2(n16426), .A(n16384), .ZN(U224) );
  AOI22_X1 U19404 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16423), .ZN(n16386) );
  OAI21_X1 U19405 ( .B1(n20185), .B2(n16426), .A(n16386), .ZN(U225) );
  AOI22_X1 U19406 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16423), .ZN(n16387) );
  OAI21_X1 U19407 ( .B1(n14876), .B2(n16426), .A(n16387), .ZN(U226) );
  AOI22_X1 U19408 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16423), .ZN(n16388) );
  OAI21_X1 U19409 ( .B1(n16389), .B2(n16426), .A(n16388), .ZN(U227) );
  AOI22_X1 U19410 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16423), .ZN(n16390) );
  OAI21_X1 U19411 ( .B1(n14887), .B2(n16426), .A(n16390), .ZN(U228) );
  AOI22_X1 U19412 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16423), .ZN(n16391) );
  OAI21_X1 U19413 ( .B1(n20163), .B2(n16426), .A(n16391), .ZN(U229) );
  AOI22_X1 U19414 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16423), .ZN(n16392) );
  OAI21_X1 U19415 ( .B1(n13685), .B2(n16426), .A(n16392), .ZN(U230) );
  AOI22_X1 U19416 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n16423), .ZN(n16393) );
  OAI21_X1 U19417 ( .B1(n20152), .B2(n16426), .A(n16393), .ZN(U231) );
  INV_X1 U19418 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16395) );
  AOI22_X1 U19419 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16423), .ZN(n16394) );
  OAI21_X1 U19420 ( .B1(n16395), .B2(n16426), .A(n16394), .ZN(U232) );
  AOI22_X1 U19421 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16423), .ZN(n16396) );
  OAI21_X1 U19422 ( .B1(n16397), .B2(n16426), .A(n16396), .ZN(U233) );
  AOI22_X1 U19423 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16423), .ZN(n16398) );
  OAI21_X1 U19424 ( .B1(n16399), .B2(n16426), .A(n16398), .ZN(U234) );
  AOI22_X1 U19425 ( .A1(P2_DATAO_REG_12__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16423), .ZN(n16400) );
  OAI21_X1 U19426 ( .B1(n16401), .B2(n16426), .A(n16400), .ZN(U235) );
  AOI22_X1 U19427 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16423), .ZN(n16402) );
  OAI21_X1 U19428 ( .B1(n16403), .B2(n16426), .A(n16402), .ZN(U236) );
  AOI22_X1 U19429 ( .A1(P2_DATAO_REG_10__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16423), .ZN(n16404) );
  OAI21_X1 U19430 ( .B1(n16405), .B2(n16426), .A(n16404), .ZN(U237) );
  AOI22_X1 U19431 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16423), .ZN(n16406) );
  OAI21_X1 U19432 ( .B1(n12897), .B2(n16426), .A(n16406), .ZN(U238) );
  AOI22_X1 U19433 ( .A1(P2_DATAO_REG_8__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(n16423), .ZN(n16407) );
  OAI21_X1 U19434 ( .B1(n16408), .B2(n16426), .A(n16407), .ZN(U239) );
  AOI22_X1 U19435 ( .A1(P2_DATAO_REG_7__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16423), .ZN(n16409) );
  OAI21_X1 U19436 ( .B1(n16410), .B2(n16426), .A(n16409), .ZN(U240) );
  AOI22_X1 U19437 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16423), .ZN(n16411) );
  OAI21_X1 U19438 ( .B1(n16412), .B2(n16426), .A(n16411), .ZN(U241) );
  AOI22_X1 U19439 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16423), .ZN(n16413) );
  OAI21_X1 U19440 ( .B1(n16414), .B2(n16426), .A(n16413), .ZN(U242) );
  AOI22_X1 U19441 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n16423), .ZN(n16415) );
  OAI21_X1 U19442 ( .B1(n16416), .B2(n16426), .A(n16415), .ZN(U243) );
  AOI22_X1 U19443 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16423), .ZN(n16417) );
  OAI21_X1 U19444 ( .B1(n16418), .B2(n16426), .A(n16417), .ZN(U244) );
  AOI22_X1 U19445 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16423), .ZN(n16419) );
  OAI21_X1 U19446 ( .B1(n16420), .B2(n16426), .A(n16419), .ZN(U245) );
  INV_X1 U19447 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16422) );
  AOI22_X1 U19448 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16423), .ZN(n16421) );
  OAI21_X1 U19449 ( .B1(n16422), .B2(n16426), .A(n16421), .ZN(U246) );
  AOI22_X1 U19450 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16424), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16423), .ZN(n16425) );
  OAI21_X1 U19451 ( .B1(n16427), .B2(n16426), .A(n16425), .ZN(U247) );
  INV_X1 U19452 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16428) );
  AOI22_X1 U19453 ( .A1(n16454), .A2(n16428), .B1(n18158), .B2(U215), .ZN(U251) );
  OAI22_X1 U19454 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16454), .ZN(n16429) );
  INV_X1 U19455 ( .A(n16429), .ZN(U252) );
  INV_X1 U19456 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16430) );
  AOI22_X1 U19457 ( .A1(n16454), .A2(n16430), .B1(n18168), .B2(U215), .ZN(U253) );
  INV_X1 U19458 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16431) );
  INV_X1 U19459 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18173) );
  AOI22_X1 U19460 ( .A1(n16454), .A2(n16431), .B1(n18173), .B2(U215), .ZN(U254) );
  INV_X1 U19461 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n16432) );
  AOI22_X1 U19462 ( .A1(n16454), .A2(n16432), .B1(n18177), .B2(U215), .ZN(U255) );
  INV_X1 U19463 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16433) );
  INV_X1 U19464 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18181) );
  AOI22_X1 U19465 ( .A1(n16454), .A2(n16433), .B1(n18181), .B2(U215), .ZN(U256) );
  INV_X1 U19466 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19467 ( .A1(n16454), .A2(n16434), .B1(n18185), .B2(U215), .ZN(U257) );
  INV_X1 U19468 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16435) );
  INV_X1 U19469 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U19470 ( .A1(n16454), .A2(n16435), .B1(n18191), .B2(U215), .ZN(U258) );
  INV_X1 U19471 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16436) );
  INV_X1 U19472 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17445) );
  AOI22_X1 U19473 ( .A1(n16460), .A2(n16436), .B1(n17445), .B2(U215), .ZN(U259) );
  INV_X1 U19474 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16437) );
  INV_X1 U19475 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17447) );
  AOI22_X1 U19476 ( .A1(n16454), .A2(n16437), .B1(n17447), .B2(U215), .ZN(U260) );
  INV_X1 U19477 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16438) );
  INV_X1 U19478 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U19479 ( .A1(n16460), .A2(n16438), .B1(n17449), .B2(U215), .ZN(U261) );
  INV_X1 U19480 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16439) );
  INV_X1 U19481 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17452) );
  AOI22_X1 U19482 ( .A1(n16454), .A2(n16439), .B1(n17452), .B2(U215), .ZN(U262) );
  INV_X1 U19483 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16440) );
  INV_X1 U19484 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U19485 ( .A1(n16454), .A2(n16440), .B1(n17454), .B2(U215), .ZN(U263) );
  INV_X1 U19486 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16441) );
  INV_X1 U19487 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U19488 ( .A1(n16460), .A2(n16441), .B1(n17458), .B2(U215), .ZN(U264) );
  OAI22_X1 U19489 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16454), .ZN(n16442) );
  INV_X1 U19490 ( .A(n16442), .ZN(U265) );
  OAI22_X1 U19491 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16454), .ZN(n16443) );
  INV_X1 U19492 ( .A(n16443), .ZN(U266) );
  OAI22_X1 U19493 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16454), .ZN(n16444) );
  INV_X1 U19494 ( .A(n16444), .ZN(U267) );
  OAI22_X1 U19495 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16454), .ZN(n16445) );
  INV_X1 U19496 ( .A(n16445), .ZN(U268) );
  OAI22_X1 U19497 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16454), .ZN(n16446) );
  INV_X1 U19498 ( .A(n16446), .ZN(U269) );
  OAI22_X1 U19499 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16454), .ZN(n16447) );
  INV_X1 U19500 ( .A(n16447), .ZN(U270) );
  OAI22_X1 U19501 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16454), .ZN(n16448) );
  INV_X1 U19502 ( .A(n16448), .ZN(U271) );
  INV_X1 U19503 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16449) );
  AOI22_X1 U19504 ( .A1(n16454), .A2(n16449), .B1(n14875), .B2(U215), .ZN(U272) );
  OAI22_X1 U19505 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16454), .ZN(n16450) );
  INV_X1 U19506 ( .A(n16450), .ZN(U273) );
  INV_X1 U19507 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n16451) );
  AOI22_X1 U19508 ( .A1(n16454), .A2(n16451), .B1(n14866), .B2(U215), .ZN(U274) );
  OAI22_X1 U19509 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16460), .ZN(n16452) );
  INV_X1 U19510 ( .A(n16452), .ZN(U275) );
  INV_X1 U19511 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n16453) );
  AOI22_X1 U19512 ( .A1(n16454), .A2(n16453), .B1(n14843), .B2(U215), .ZN(U276) );
  OAI22_X1 U19513 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16460), .ZN(n16455) );
  INV_X1 U19514 ( .A(n16455), .ZN(U277) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16460), .ZN(n16456) );
  INV_X1 U19516 ( .A(n16456), .ZN(U278) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16460), .ZN(n16457) );
  INV_X1 U19518 ( .A(n16457), .ZN(U279) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16460), .ZN(n16458) );
  INV_X1 U19520 ( .A(n16458), .ZN(U280) );
  OAI22_X1 U19521 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16460), .ZN(n16459) );
  INV_X1 U19522 ( .A(n16459), .ZN(U281) );
  INV_X1 U19523 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18190) );
  AOI22_X1 U19524 ( .A1(n16460), .A2(n16463), .B1(n18190), .B2(U215), .ZN(U282) );
  INV_X1 U19525 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16461) );
  AOI222_X1 U19526 ( .A1(n16463), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16462), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n16461), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16464) );
  INV_X2 U19527 ( .A(n16466), .ZN(n16465) );
  INV_X1 U19528 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18698) );
  INV_X1 U19529 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19867) );
  AOI22_X1 U19530 ( .A1(n16465), .A2(n18698), .B1(n19867), .B2(n16466), .ZN(
        U347) );
  INV_X1 U19531 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18696) );
  INV_X1 U19532 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19866) );
  AOI22_X1 U19533 ( .A1(n16465), .A2(n18696), .B1(n19866), .B2(n16466), .ZN(
        U348) );
  INV_X1 U19534 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18693) );
  INV_X1 U19535 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19864) );
  AOI22_X1 U19536 ( .A1(n16465), .A2(n18693), .B1(n19864), .B2(n16466), .ZN(
        U349) );
  INV_X1 U19537 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18692) );
  INV_X1 U19538 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19863) );
  AOI22_X1 U19539 ( .A1(n16465), .A2(n18692), .B1(n19863), .B2(n16466), .ZN(
        U350) );
  INV_X1 U19540 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18690) );
  INV_X1 U19541 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19861) );
  AOI22_X1 U19542 ( .A1(n16465), .A2(n18690), .B1(n19861), .B2(n16466), .ZN(
        U351) );
  INV_X1 U19543 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18687) );
  INV_X1 U19544 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19860) );
  AOI22_X1 U19545 ( .A1(n16465), .A2(n18687), .B1(n19860), .B2(n16466), .ZN(
        U352) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18686) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19859) );
  AOI22_X1 U19548 ( .A1(n16465), .A2(n18686), .B1(n19859), .B2(n16466), .ZN(
        U353) );
  INV_X1 U19549 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18684) );
  AOI22_X1 U19550 ( .A1(n16465), .A2(n18684), .B1(n19858), .B2(n16466), .ZN(
        U354) );
  INV_X1 U19551 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18737) );
  INV_X1 U19552 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19897) );
  AOI22_X1 U19553 ( .A1(n16465), .A2(n18737), .B1(n19897), .B2(n16466), .ZN(
        U356) );
  INV_X1 U19554 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18734) );
  INV_X1 U19555 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19895) );
  AOI22_X1 U19556 ( .A1(n16465), .A2(n18734), .B1(n19895), .B2(n16466), .ZN(
        U357) );
  INV_X1 U19557 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18732) );
  INV_X1 U19558 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19893) );
  AOI22_X1 U19559 ( .A1(n16465), .A2(n18732), .B1(n19893), .B2(n16466), .ZN(
        U358) );
  INV_X1 U19560 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18730) );
  INV_X1 U19561 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19891) );
  AOI22_X1 U19562 ( .A1(n16465), .A2(n18730), .B1(n19891), .B2(n16466), .ZN(
        U359) );
  INV_X1 U19563 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18728) );
  INV_X1 U19564 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19889) );
  AOI22_X1 U19565 ( .A1(n16465), .A2(n18728), .B1(n19889), .B2(n16466), .ZN(
        U360) );
  INV_X1 U19566 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18726) );
  INV_X1 U19567 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19887) );
  AOI22_X1 U19568 ( .A1(n16465), .A2(n18726), .B1(n19887), .B2(n16466), .ZN(
        U361) );
  INV_X1 U19569 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18723) );
  INV_X1 U19570 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19886) );
  AOI22_X1 U19571 ( .A1(n16465), .A2(n18723), .B1(n19886), .B2(n16466), .ZN(
        U362) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18722) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19884) );
  AOI22_X1 U19574 ( .A1(n16465), .A2(n18722), .B1(n19884), .B2(n16466), .ZN(
        U363) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18719) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19883) );
  AOI22_X1 U19577 ( .A1(n16465), .A2(n18719), .B1(n19883), .B2(n16466), .ZN(
        U364) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18682) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19857) );
  AOI22_X1 U19580 ( .A1(n16465), .A2(n18682), .B1(n19857), .B2(n16466), .ZN(
        U365) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18718) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19881) );
  AOI22_X1 U19583 ( .A1(n16465), .A2(n18718), .B1(n19881), .B2(n16466), .ZN(
        U366) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18715) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19879) );
  AOI22_X1 U19586 ( .A1(n16465), .A2(n18715), .B1(n19879), .B2(n16466), .ZN(
        U367) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18714) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19877) );
  AOI22_X1 U19589 ( .A1(n16465), .A2(n18714), .B1(n19877), .B2(n16466), .ZN(
        U368) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18711) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19876) );
  AOI22_X1 U19592 ( .A1(n16465), .A2(n18711), .B1(n19876), .B2(n16466), .ZN(
        U369) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18710) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19874) );
  AOI22_X1 U19595 ( .A1(n16465), .A2(n18710), .B1(n19874), .B2(n16466), .ZN(
        U370) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18707) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19872) );
  AOI22_X1 U19598 ( .A1(n16465), .A2(n18707), .B1(n19872), .B2(n16466), .ZN(
        U371) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18706) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19871) );
  AOI22_X1 U19601 ( .A1(n16465), .A2(n18706), .B1(n19871), .B2(n16466), .ZN(
        U372) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18704) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19870) );
  AOI22_X1 U19604 ( .A1(n16465), .A2(n18704), .B1(n19870), .B2(n16466), .ZN(
        U373) );
  INV_X1 U19605 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18702) );
  INV_X1 U19606 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19869) );
  AOI22_X1 U19607 ( .A1(n16465), .A2(n18702), .B1(n19869), .B2(n16466), .ZN(
        U374) );
  INV_X1 U19608 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18700) );
  INV_X1 U19609 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19868) );
  AOI22_X1 U19610 ( .A1(n16465), .A2(n18700), .B1(n19868), .B2(n16466), .ZN(
        U375) );
  INV_X1 U19611 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18680) );
  INV_X1 U19612 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19856) );
  AOI22_X1 U19613 ( .A1(n16465), .A2(n18680), .B1(n19856), .B2(n16466), .ZN(
        U376) );
  INV_X1 U19614 ( .A(P3_ADS_N_REG_SCAN_IN), .ZN(n16467) );
  NAND2_X1 U19615 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18679), .ZN(n18666) );
  AOI22_X1 U19616 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18666), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18677), .ZN(n18755) );
  INV_X1 U19617 ( .A(n18755), .ZN(n18660) );
  CLKBUF_X1 U19618 ( .A(n18660), .Z(n18752) );
  OAI21_X1 U19619 ( .B1(n18677), .B2(n16467), .A(n18752), .ZN(P3_U2633) );
  INV_X1 U19620 ( .A(n18821), .ZN(n16469) );
  OAI21_X1 U19621 ( .B1(n16473), .B2(n17414), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16468) );
  OAI21_X1 U19622 ( .B1(n16469), .B2(n18652), .A(n16468), .ZN(P3_U2634) );
  AOI21_X1 U19623 ( .B1(n18677), .B2(n18679), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16470) );
  AOI22_X1 U19624 ( .A1(n18733), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16470), 
        .B2(n18799), .ZN(P3_U2635) );
  INV_X1 U19625 ( .A(BS16), .ZN(n20943) );
  AOI21_X1 U19626 ( .B1(n18661), .B2(n20943), .A(n18752), .ZN(n18750) );
  INV_X1 U19627 ( .A(n18750), .ZN(n18753) );
  OAI21_X1 U19628 ( .B1(n18755), .B2(n18807), .A(n18753), .ZN(P3_U2636) );
  NOR3_X1 U19629 ( .A1(n16473), .A2(n16472), .A3(n16471), .ZN(n18589) );
  NOR2_X1 U19630 ( .A1(n18589), .A2(n18649), .ZN(n18801) );
  OAI21_X1 U19631 ( .B1(n18801), .B2(n16475), .A(n16474), .ZN(P3_U2637) );
  NOR4_X1 U19632 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16479) );
  NOR4_X1 U19633 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16478) );
  NOR4_X1 U19634 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16477) );
  NOR4_X1 U19635 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16476) );
  NAND4_X1 U19636 ( .A1(n16479), .A2(n16478), .A3(n16477), .A4(n16476), .ZN(
        n16485) );
  NOR4_X1 U19637 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16483) );
  AOI211_X1 U19638 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16482) );
  NOR4_X1 U19639 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16481) );
  NOR4_X1 U19640 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16480) );
  NAND4_X1 U19641 ( .A1(n16483), .A2(n16482), .A3(n16481), .A4(n16480), .ZN(
        n16484) );
  NOR2_X1 U19642 ( .A1(n16485), .A2(n16484), .ZN(n18798) );
  INV_X1 U19643 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18748) );
  NOR3_X1 U19644 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16487) );
  OAI21_X1 U19645 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16487), .A(n18798), .ZN(
        n16486) );
  OAI21_X1 U19646 ( .B1(n18798), .B2(n18748), .A(n16486), .ZN(P3_U2638) );
  INV_X1 U19647 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18791) );
  INV_X1 U19648 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18754) );
  AOI21_X1 U19649 ( .B1(n18791), .B2(n18754), .A(n16487), .ZN(n16488) );
  INV_X1 U19650 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18745) );
  INV_X1 U19651 ( .A(n18798), .ZN(n18793) );
  AOI22_X1 U19652 ( .A1(n18798), .A2(n16488), .B1(n18745), .B2(n18793), .ZN(
        P3_U2639) );
  NOR2_X2 U19653 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18758), .ZN(n18523) );
  NAND2_X1 U19654 ( .A1(n18523), .A2(n18813), .ZN(n18645) );
  NOR2_X1 U19655 ( .A1(n18042), .A2(n18653), .ZN(n16823) );
  INV_X1 U19656 ( .A(n18824), .ZN(n18819) );
  AOI211_X1 U19657 ( .C1(n18808), .C2(n18806), .A(n18669), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16490) );
  AOI211_X4 U19658 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18164), .A(n16490), .B(
        n18822), .ZN(n16873) );
  INV_X1 U19659 ( .A(n16490), .ZN(n18644) );
  INV_X1 U19660 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18727) );
  INV_X1 U19661 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18724) );
  INV_X1 U19662 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18720) );
  INV_X1 U19663 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18705) );
  INV_X1 U19664 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18701) );
  INV_X1 U19665 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18685) );
  NAND3_X1 U19666 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16813) );
  NOR2_X1 U19667 ( .A1(n18685), .A2(n16813), .ZN(n16802) );
  NAND2_X1 U19668 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16802), .ZN(n16800) );
  NAND3_X1 U19669 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_7__SCAN_IN), 
        .A3(P3_REIP_REG_6__SCAN_IN), .ZN(n16725) );
  NOR2_X1 U19670 ( .A1(n16800), .A2(n16725), .ZN(n16737) );
  NAND4_X1 U19671 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16737), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16719) );
  NOR2_X1 U19672 ( .A1(n18701), .A2(n16719), .ZN(n16701) );
  NAND2_X1 U19673 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16701), .ZN(n16688) );
  NOR2_X1 U19674 ( .A1(n18705), .A2(n16688), .ZN(n16687) );
  NAND2_X1 U19675 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16687), .ZN(n16629) );
  NAND2_X1 U19676 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16628) );
  NAND2_X1 U19677 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16636) );
  NOR3_X1 U19678 ( .A1(n16629), .A2(n16628), .A3(n16636), .ZN(n16618) );
  NAND2_X1 U19679 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16618), .ZN(n16613) );
  NOR2_X1 U19680 ( .A1(n18720), .A2(n16613), .ZN(n16603) );
  NAND2_X1 U19681 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16603), .ZN(n16586) );
  NOR2_X1 U19682 ( .A1(n18724), .A2(n16586), .ZN(n16578) );
  NAND2_X1 U19683 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16578), .ZN(n16569) );
  NOR2_X1 U19684 ( .A1(n18727), .A2(n16569), .ZN(n16554) );
  NAND2_X1 U19685 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16554), .ZN(n16506) );
  NOR2_X1 U19686 ( .A1(n16864), .A2(n16506), .ZN(n16534) );
  NAND4_X1 U19687 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16534), .ZN(n16508) );
  NOR3_X1 U19688 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18742), .A3(n16508), 
        .ZN(n16491) );
  AOI21_X1 U19689 ( .B1(n16873), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16491), .ZN(
        n16513) );
  NAND2_X1 U19690 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18164), .ZN(n16492) );
  AOI211_X4 U19691 ( .C1(n18807), .C2(n18809), .A(n18822), .B(n16492), .ZN(
        n16872) );
  NOR3_X1 U19692 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16842) );
  NAND2_X1 U19693 ( .A1(n16842), .A2(n16841), .ZN(n16838) );
  NOR2_X1 U19694 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16838), .ZN(n16811) );
  INV_X1 U19695 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16806) );
  NAND2_X1 U19696 ( .A1(n16811), .A2(n16806), .ZN(n16803) );
  NAND2_X1 U19697 ( .A1(n16787), .A2(n17166), .ZN(n16784) );
  NAND2_X1 U19698 ( .A1(n16763), .A2(n16762), .ZN(n16759) );
  NAND2_X1 U19699 ( .A1(n16738), .A2(n16733), .ZN(n16732) );
  NAND2_X1 U19700 ( .A1(n16715), .A2(n16714), .ZN(n16711) );
  INV_X1 U19701 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16683) );
  NAND2_X1 U19702 ( .A1(n16693), .A2(n16683), .ZN(n16682) );
  INV_X1 U19703 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16655) );
  NAND2_X1 U19704 ( .A1(n16667), .A2(n16655), .ZN(n16654) );
  INV_X1 U19705 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16638) );
  NAND2_X1 U19706 ( .A1(n16643), .A2(n16638), .ZN(n16637) );
  NAND2_X1 U19707 ( .A1(n16621), .A2(n16973), .ZN(n16614) );
  NAND2_X1 U19708 ( .A1(n16597), .A2(n16593), .ZN(n16592) );
  NOR2_X1 U19709 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16592), .ZN(n16565) );
  NAND2_X1 U19710 ( .A1(n16565), .A2(n16882), .ZN(n16556) );
  NOR2_X1 U19711 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16556), .ZN(n16555) );
  NAND2_X1 U19712 ( .A1(n16555), .A2(n16924), .ZN(n16549) );
  NOR2_X1 U19713 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16549), .ZN(n16535) );
  INV_X1 U19714 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16916) );
  NAND2_X1 U19715 ( .A1(n16535), .A2(n16916), .ZN(n16514) );
  NOR2_X1 U19716 ( .A1(n16863), .A2(n16514), .ZN(n16520) );
  INV_X1 U19717 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16909) );
  OAI21_X1 U19718 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16495), .A(
        n16493), .ZN(n16494) );
  INV_X1 U19719 ( .A(n16494), .ZN(n17468) );
  AOI21_X1 U19720 ( .B1(n17489), .B2(n16496), .A(n16495), .ZN(n17486) );
  AOI21_X1 U19721 ( .B1(n16564), .B2(n17467), .A(n16497), .ZN(n17497) );
  INV_X1 U19722 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17522) );
  INV_X1 U19723 ( .A(n16500), .ZN(n16499) );
  NOR2_X1 U19724 ( .A1(n17522), .A2(n16499), .ZN(n16498) );
  OAI21_X1 U19725 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16498), .A(
        n17467), .ZN(n17511) );
  INV_X1 U19726 ( .A(n17511), .ZN(n16568) );
  AOI21_X1 U19727 ( .B1(n17522), .B2(n16499), .A(n16498), .ZN(n17520) );
  INV_X1 U19728 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17541) );
  INV_X1 U19729 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16502) );
  NOR2_X1 U19730 ( .A1(n17825), .A2(n17589), .ZN(n17588) );
  INV_X1 U19731 ( .A(n17588), .ZN(n16652) );
  NOR2_X1 U19732 ( .A1(n17591), .A2(n16652), .ZN(n17551) );
  INV_X1 U19733 ( .A(n17551), .ZN(n16631) );
  NOR2_X1 U19734 ( .A1(n10038), .A2(n16631), .ZN(n16504) );
  NAND2_X1 U19735 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16504), .ZN(
        n16503) );
  NOR2_X1 U19736 ( .A1(n16502), .A2(n16503), .ZN(n16501) );
  INV_X1 U19737 ( .A(n16501), .ZN(n17506) );
  AOI21_X1 U19738 ( .B1(n17541), .B2(n17506), .A(n16500), .ZN(n17538) );
  AOI21_X1 U19739 ( .B1(n16502), .B2(n16503), .A(n16501), .ZN(n17553) );
  OAI21_X1 U19740 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16504), .A(
        n16503), .ZN(n17568) );
  INV_X1 U19741 ( .A(n17568), .ZN(n16609) );
  AOI21_X1 U19742 ( .B1(n10038), .B2(n16631), .A(n16504), .ZN(n17581) );
  NOR2_X1 U19743 ( .A1(n17825), .A2(n17624), .ZN(n17626) );
  NAND2_X1 U19744 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17626), .ZN(
        n16674) );
  NOR2_X1 U19745 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16674), .ZN(
        n16664) );
  AND2_X1 U19746 ( .A1(n17551), .A2(n16664), .ZN(n16505) );
  NOR2_X1 U19747 ( .A1(n17581), .A2(n16620), .ZN(n16619) );
  NOR2_X1 U19748 ( .A1(n16619), .A2(n16798), .ZN(n16608) );
  NOR2_X1 U19749 ( .A1(n16607), .A2(n16798), .ZN(n16599) );
  NOR2_X1 U19750 ( .A1(n17553), .A2(n16599), .ZN(n16598) );
  NOR2_X1 U19751 ( .A1(n16598), .A2(n16798), .ZN(n16588) );
  NOR2_X1 U19752 ( .A1(n16587), .A2(n16798), .ZN(n16581) );
  NOR2_X1 U19753 ( .A1(n17520), .A2(n16581), .ZN(n16580) );
  NOR2_X1 U19754 ( .A1(n16580), .A2(n16798), .ZN(n16567) );
  NOR2_X1 U19755 ( .A1(n16566), .A2(n16798), .ZN(n16558) );
  NOR2_X1 U19756 ( .A1(n17497), .A2(n16558), .ZN(n16557) );
  NOR2_X1 U19757 ( .A1(n16557), .A2(n16798), .ZN(n16545) );
  NOR2_X1 U19758 ( .A1(n16544), .A2(n16798), .ZN(n16537) );
  NOR2_X1 U19759 ( .A1(n17468), .A2(n16537), .ZN(n16536) );
  NOR2_X1 U19760 ( .A1(n16536), .A2(n16798), .ZN(n16524) );
  NOR2_X1 U19761 ( .A1(n16523), .A2(n16798), .ZN(n16515) );
  NAND2_X1 U19762 ( .A1(n16818), .A2(n18653), .ZN(n16858) );
  NOR3_X1 U19763 ( .A1(n16516), .A2(n16515), .A3(n16858), .ZN(n16511) );
  NAND3_X1 U19764 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16507) );
  AND2_X1 U19765 ( .A1(n16828), .A2(n16506), .ZN(n16553) );
  NOR2_X1 U19766 ( .A1(n16868), .A2(n16553), .ZN(n16552) );
  INV_X1 U19767 ( .A(n16552), .ZN(n16561) );
  AOI21_X1 U19768 ( .B1(n16828), .B2(n16507), .A(n16561), .ZN(n16533) );
  NOR2_X1 U19769 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16508), .ZN(n16518) );
  INV_X1 U19770 ( .A(n16518), .ZN(n16509) );
  AOI21_X1 U19771 ( .B1(n16533), .B2(n16509), .A(n18740), .ZN(n16510) );
  AOI211_X1 U19772 ( .C1(n16520), .C2(n16909), .A(n16511), .B(n16510), .ZN(
        n16512) );
  OAI211_X1 U19773 ( .C1(n10052), .C2(n16857), .A(n16513), .B(n16512), .ZN(
        P3_U2640) );
  NAND2_X1 U19774 ( .A1(n16872), .A2(n16514), .ZN(n16529) );
  XOR2_X1 U19775 ( .A(n16516), .B(n16515), .Z(n16519) );
  OAI22_X1 U19776 ( .A1(n16533), .A2(n18742), .B1(n10053), .B2(n16857), .ZN(
        n16517) );
  AOI211_X1 U19777 ( .C1(n16519), .C2(n18653), .A(n16518), .B(n16517), .ZN(
        n16522) );
  OAI21_X1 U19778 ( .B1(n16873), .B2(n16520), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16521) );
  OAI211_X1 U19779 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16529), .A(n16522), .B(
        n16521), .ZN(P3_U2641) );
  INV_X1 U19780 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18736) );
  INV_X1 U19781 ( .A(n18653), .ZN(n16775) );
  AOI211_X1 U19782 ( .C1(n16525), .C2(n16524), .A(n16523), .B(n16775), .ZN(
        n16528) );
  NAND3_X1 U19783 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16534), .ZN(n16526) );
  OAI22_X1 U19784 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16526), .B1(n10051), 
        .B2(n16857), .ZN(n16527) );
  AOI211_X1 U19785 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16873), .A(n16528), .B(
        n16527), .ZN(n16532) );
  INV_X1 U19786 ( .A(n16529), .ZN(n16530) );
  OAI21_X1 U19787 ( .B1(n16535), .B2(n16916), .A(n16530), .ZN(n16531) );
  OAI211_X1 U19788 ( .C1(n16533), .C2(n18736), .A(n16532), .B(n16531), .ZN(
        P3_U2642) );
  NAND2_X1 U19789 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16534), .ZN(n16543) );
  AOI22_X1 U19790 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16851), .B1(
        n16873), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16542) );
  INV_X1 U19791 ( .A(n16534), .ZN(n16546) );
  OAI21_X1 U19792 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16546), .A(n16552), 
        .ZN(n16540) );
  AOI211_X1 U19793 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16549), .A(n16535), .B(
        n16863), .ZN(n16539) );
  AOI211_X1 U19794 ( .C1(n17468), .C2(n16537), .A(n16536), .B(n16775), .ZN(
        n16538) );
  AOI211_X1 U19795 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16540), .A(n16539), 
        .B(n16538), .ZN(n16541) );
  OAI211_X1 U19796 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16543), .A(n16542), 
        .B(n16541), .ZN(P3_U2643) );
  INV_X1 U19797 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18731) );
  AOI211_X1 U19798 ( .C1(n17486), .C2(n16545), .A(n16544), .B(n16775), .ZN(
        n16548) );
  OAI22_X1 U19799 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16546), .B1(n17489), 
        .B2(n16857), .ZN(n16547) );
  AOI211_X1 U19800 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16873), .A(n16548), .B(
        n16547), .ZN(n16551) );
  OAI211_X1 U19801 ( .C1(n16555), .C2(n16924), .A(n16872), .B(n16549), .ZN(
        n16550) );
  OAI211_X1 U19802 ( .C1(n16552), .C2(n18731), .A(n16551), .B(n16550), .ZN(
        P3_U2644) );
  AOI22_X1 U19803 ( .A1(n16873), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16554), 
        .B2(n16553), .ZN(n16563) );
  AOI211_X1 U19804 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16556), .A(n16555), .B(
        n16863), .ZN(n16560) );
  AOI211_X1 U19805 ( .C1(n17497), .C2(n16558), .A(n16557), .B(n16775), .ZN(
        n16559) );
  AOI211_X1 U19806 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16561), .A(n16560), 
        .B(n16559), .ZN(n16562) );
  OAI211_X1 U19807 ( .C1(n16564), .C2(n16857), .A(n16563), .B(n16562), .ZN(
        P3_U2645) );
  OR2_X1 U19808 ( .A1(n16863), .A2(n16565), .ZN(n16579) );
  AOI21_X1 U19809 ( .B1(n16872), .B2(n16565), .A(n16873), .ZN(n16576) );
  AOI211_X1 U19810 ( .C1(n16568), .C2(n16567), .A(n16566), .B(n16775), .ZN(
        n16574) );
  NOR2_X1 U19811 ( .A1(n16864), .A2(n16569), .ZN(n16572) );
  INV_X1 U19812 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18725) );
  OAI21_X1 U19813 ( .B1(n16578), .B2(n16864), .A(n16877), .ZN(n16591) );
  AOI21_X1 U19814 ( .B1(n16828), .B2(n18725), .A(n16591), .ZN(n16570) );
  INV_X1 U19815 ( .A(n16570), .ZN(n16571) );
  MUX2_X1 U19816 ( .A(n16572), .B(n16571), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16573) );
  AOI211_X1 U19817 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16574), .B(n16573), .ZN(n16575) );
  OAI221_X1 U19818 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16579), .C1(n16882), 
        .C2(n16576), .A(n16575), .ZN(P3_U2646) );
  NOR2_X1 U19819 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16864), .ZN(n16577) );
  AOI22_X1 U19820 ( .A1(n16873), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16578), 
        .B2(n16577), .ZN(n16585) );
  AOI21_X1 U19821 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16592), .A(n16579), .ZN(
        n16583) );
  AOI211_X1 U19822 ( .C1(n17520), .C2(n16581), .A(n16580), .B(n16775), .ZN(
        n16582) );
  AOI211_X1 U19823 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16591), .A(n16583), 
        .B(n16582), .ZN(n16584) );
  OAI211_X1 U19824 ( .C1(n17522), .C2(n16857), .A(n16585), .B(n16584), .ZN(
        P3_U2647) );
  AOI22_X1 U19825 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16851), .B1(
        n16873), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16596) );
  OAI21_X1 U19826 ( .B1(n16864), .B2(n16586), .A(n18724), .ZN(n16590) );
  AOI211_X1 U19827 ( .C1(n17538), .C2(n16588), .A(n16587), .B(n16775), .ZN(
        n16589) );
  AOI21_X1 U19828 ( .B1(n16591), .B2(n16590), .A(n16589), .ZN(n16595) );
  OAI211_X1 U19829 ( .C1(n16597), .C2(n16593), .A(n16872), .B(n16592), .ZN(
        n16594) );
  NAND3_X1 U19830 ( .A1(n16596), .A2(n16595), .A3(n16594), .ZN(P3_U2648) );
  AOI221_X1 U19831 ( .B1(n18720), .B2(n16828), .C1(n16613), .C2(n16828), .A(
        n16868), .ZN(n16606) );
  INV_X1 U19832 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18721) );
  AOI22_X1 U19833 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16851), .B1(
        n16873), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16605) );
  NOR2_X1 U19834 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16864), .ZN(n16602) );
  AOI211_X1 U19835 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16614), .A(n16597), .B(
        n16863), .ZN(n16601) );
  AOI211_X1 U19836 ( .C1(n17553), .C2(n16599), .A(n16598), .B(n16775), .ZN(
        n16600) );
  AOI211_X1 U19837 ( .C1(n16603), .C2(n16602), .A(n16601), .B(n16600), .ZN(
        n16604) );
  OAI211_X1 U19838 ( .C1(n16606), .C2(n18721), .A(n16605), .B(n16604), .ZN(
        P3_U2649) );
  AOI21_X1 U19839 ( .B1(n16613), .B2(n16828), .A(n16868), .ZN(n16626) );
  INV_X1 U19840 ( .A(n16626), .ZN(n16612) );
  AOI211_X1 U19841 ( .C1(n16609), .C2(n16608), .A(n16607), .B(n16775), .ZN(
        n16611) );
  INV_X1 U19842 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17571) );
  OAI22_X1 U19843 ( .A1(n17571), .A2(n16857), .B1(n16860), .B2(n16973), .ZN(
        n16610) );
  AOI211_X1 U19844 ( .C1(n16612), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16611), 
        .B(n16610), .ZN(n16617) );
  OR3_X1 U19845 ( .A1(n16864), .A2(n16613), .A3(P3_REIP_REG_21__SCAN_IN), .ZN(
        n16616) );
  OAI211_X1 U19846 ( .C1(n16621), .C2(n16973), .A(n16872), .B(n16614), .ZN(
        n16615) );
  NAND3_X1 U19847 ( .A1(n16617), .A2(n16616), .A3(n16615), .ZN(P3_U2650) );
  AOI21_X1 U19848 ( .B1(n16828), .B2(n16618), .A(P3_REIP_REG_20__SCAN_IN), 
        .ZN(n16627) );
  AOI211_X1 U19849 ( .C1(n17581), .C2(n16620), .A(n16619), .B(n16775), .ZN(
        n16624) );
  AOI211_X1 U19850 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16637), .A(n16621), .B(
        n16863), .ZN(n16623) );
  OAI22_X1 U19851 ( .A1(n10038), .A2(n16857), .B1(n16860), .B2(n16988), .ZN(
        n16622) );
  NOR3_X1 U19852 ( .A1(n16624), .A2(n16623), .A3(n16622), .ZN(n16625) );
  OAI21_X1 U19853 ( .B1(n16627), .B2(n16626), .A(n16625), .ZN(P3_U2651) );
  INV_X1 U19854 ( .A(n16628), .ZN(n16630) );
  NOR2_X1 U19855 ( .A1(n16868), .A2(n16828), .ZN(n16874) );
  AOI21_X1 U19856 ( .B1(n16828), .B2(n16629), .A(n16868), .ZN(n16675) );
  OAI21_X1 U19857 ( .B1(n16630), .B2(n16874), .A(n16675), .ZN(n16659) );
  INV_X1 U19858 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17602) );
  NOR2_X1 U19859 ( .A1(n17602), .A2(n16652), .ZN(n16632) );
  OAI21_X1 U19860 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16632), .A(
        n16631), .ZN(n17594) );
  NAND2_X1 U19861 ( .A1(n17588), .A2(n16664), .ZN(n16645) );
  OAI21_X1 U19862 ( .B1(n17602), .B2(n16645), .A(n16818), .ZN(n16633) );
  XNOR2_X1 U19863 ( .A(n17594), .B(n16633), .ZN(n16634) );
  OAI22_X1 U19864 ( .A1(n16860), .A2(n16638), .B1(n16775), .B2(n16634), .ZN(
        n16635) );
  AOI211_X1 U19865 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16659), .A(n18042), 
        .B(n16635), .ZN(n16642) );
  INV_X1 U19866 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18712) );
  NAND4_X1 U19867 ( .A1(n16828), .A2(P3_REIP_REG_15__SCAN_IN), .A3(n16687), 
        .A4(P3_REIP_REG_16__SCAN_IN), .ZN(n16662) );
  NOR2_X1 U19868 ( .A1(n18712), .A2(n16662), .ZN(n16648) );
  OAI211_X1 U19869 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16648), .B(n16636), .ZN(n16641) );
  OAI211_X1 U19870 ( .C1(n16643), .C2(n16638), .A(n16872), .B(n16637), .ZN(
        n16640) );
  NAND2_X1 U19871 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16851), .ZN(
        n16639) );
  NAND4_X1 U19872 ( .A1(n16642), .A2(n16641), .A3(n16640), .A4(n16639), .ZN(
        P3_U2652) );
  AOI211_X1 U19873 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16654), .A(n16643), .B(
        n16863), .ZN(n16644) );
  AOI21_X1 U19874 ( .B1(n16851), .B2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16644), .ZN(n16651) );
  AOI22_X1 U19875 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n16652), .B1(
        n17588), .B2(n17602), .ZN(n17599) );
  NAND2_X1 U19876 ( .A1(n16818), .A2(n16645), .ZN(n16646) );
  XOR2_X1 U19877 ( .A(n17599), .B(n16646), .Z(n16647) );
  AOI22_X1 U19878 ( .A1(n16873), .A2(P3_EBX_REG_18__SCAN_IN), .B1(n18653), 
        .B2(n16647), .ZN(n16650) );
  INV_X1 U19879 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18713) );
  AOI22_X1 U19880 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16659), .B1(n16648), 
        .B2(n18713), .ZN(n16649) );
  NAND4_X1 U19881 ( .A1(n16651), .A2(n16650), .A3(n16649), .A4(n18036), .ZN(
        P3_U2653) );
  AOI22_X1 U19882 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16851), .B1(
        n16873), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16661) );
  AND2_X1 U19883 ( .A1(n17611), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16663) );
  INV_X1 U19884 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16859) );
  AOI21_X1 U19885 ( .B1(n16663), .B2(n16859), .A(n16798), .ZN(n16653) );
  OAI21_X1 U19886 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16663), .A(
        n16652), .ZN(n17619) );
  XOR2_X1 U19887 ( .A(n16653), .B(n17619), .Z(n16657) );
  OAI211_X1 U19888 ( .C1(n16667), .C2(n16655), .A(n16872), .B(n16654), .ZN(
        n16656) );
  OAI211_X1 U19889 ( .C1(n16775), .C2(n16657), .A(n18036), .B(n16656), .ZN(
        n16658) );
  AOI21_X1 U19890 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(n16659), .A(n16658), 
        .ZN(n16660) );
  OAI211_X1 U19891 ( .C1(P3_REIP_REG_17__SCAN_IN), .C2(n16662), .A(n16661), 
        .B(n16660), .ZN(P3_U2654) );
  NAND3_X1 U19892 ( .A1(n16828), .A2(P3_REIP_REG_15__SCAN_IN), .A3(n16687), 
        .ZN(n16673) );
  INV_X1 U19893 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18709) );
  INV_X1 U19894 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16668) );
  AOI21_X1 U19895 ( .B1(n16668), .B2(n16674), .A(n16663), .ZN(n17627) );
  NOR2_X1 U19896 ( .A1(n16664), .A2(n16798), .ZN(n16681) );
  INV_X1 U19897 ( .A(n17627), .ZN(n16666) );
  INV_X1 U19898 ( .A(n16681), .ZN(n16665) );
  AOI221_X1 U19899 ( .B1(n17627), .B2(n16681), .C1(n16666), .C2(n16665), .A(
        n16775), .ZN(n16671) );
  AOI211_X1 U19900 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16682), .A(n16667), .B(
        n16863), .ZN(n16670) );
  INV_X1 U19901 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17046) );
  OAI22_X1 U19902 ( .A1(n16668), .A2(n16857), .B1(n16860), .B2(n17046), .ZN(
        n16669) );
  NOR4_X1 U19903 ( .A1(n9821), .A2(n16671), .A3(n16670), .A4(n16669), .ZN(
        n16672) );
  OAI221_X1 U19904 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16673), .C1(n18709), 
        .C2(n16675), .A(n16672), .ZN(P3_U2655) );
  NOR2_X1 U19905 ( .A1(n16818), .A2(n16775), .ZN(n16777) );
  INV_X1 U19906 ( .A(n16777), .ZN(n16844) );
  OAI21_X1 U19907 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17626), .A(
        n16674), .ZN(n17634) );
  OAI21_X1 U19908 ( .B1(n16798), .B2(n16859), .A(n18653), .ZN(n16861) );
  AOI211_X1 U19909 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16844), .A(
        n17634), .B(n16861), .ZN(n16680) );
  INV_X1 U19910 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18708) );
  NAND2_X1 U19911 ( .A1(n16828), .A2(n16687), .ZN(n16676) );
  AOI21_X1 U19912 ( .B1(n18708), .B2(n16676), .A(n16675), .ZN(n16679) );
  INV_X1 U19913 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16677) );
  OAI22_X1 U19914 ( .A1(n16677), .A2(n16857), .B1(n16860), .B2(n16683), .ZN(
        n16678) );
  NOR3_X1 U19915 ( .A1(n16680), .A2(n16679), .A3(n16678), .ZN(n16686) );
  NAND3_X1 U19916 ( .A1(n18653), .A2(n16681), .A3(n17634), .ZN(n16685) );
  OAI211_X1 U19917 ( .C1(n16693), .C2(n16683), .A(n16872), .B(n16682), .ZN(
        n16684) );
  NAND4_X1 U19918 ( .A1(n16686), .A2(n18036), .A3(n16685), .A4(n16684), .ZN(
        P3_U2656) );
  AOI211_X1 U19919 ( .C1(n18705), .C2(n16688), .A(n16687), .B(n16864), .ZN(
        n16699) );
  INV_X1 U19920 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16689) );
  NAND3_X1 U19921 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17768), .A3(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16788) );
  NOR2_X1 U19922 ( .A1(n16690), .A2(n16788), .ZN(n17665) );
  NAND2_X1 U19923 ( .A1(n17664), .A2(n17665), .ZN(n16703) );
  AOI21_X1 U19924 ( .B1(n16689), .B2(n16703), .A(n17626), .ZN(n17659) );
  INV_X1 U19925 ( .A(n17691), .ZN(n17731) );
  NOR2_X1 U19926 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17825), .ZN(
        n16853) );
  NAND2_X1 U19927 ( .A1(n17731), .A2(n16853), .ZN(n16790) );
  OAI21_X1 U19928 ( .B1(n16690), .B2(n16790), .A(n16818), .ZN(n16717) );
  OAI21_X1 U19929 ( .B1(n17664), .B2(n16798), .A(n16717), .ZN(n16705) );
  INV_X1 U19930 ( .A(n17659), .ZN(n16692) );
  INV_X1 U19931 ( .A(n16705), .ZN(n16691) );
  OAI221_X1 U19932 ( .B1(n17659), .B2(n16705), .C1(n16692), .C2(n16691), .A(
        n18653), .ZN(n16696) );
  AOI211_X1 U19933 ( .C1(n16711), .C2(P3_EBX_REG_14__SCAN_IN), .A(n16863), .B(
        n16693), .ZN(n16694) );
  INV_X1 U19934 ( .A(n16694), .ZN(n16695) );
  OAI211_X1 U19935 ( .C1(n16697), .C2(n16860), .A(n16696), .B(n16695), .ZN(
        n16698) );
  AOI211_X1 U19936 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16699), .B(n16698), .ZN(n16700) );
  OAI211_X1 U19937 ( .C1(n16877), .C2(n18705), .A(n16700), .B(n18036), .ZN(
        P3_U2657) );
  AOI21_X1 U19938 ( .B1(n16828), .B2(n16719), .A(n16868), .ZN(n16729) );
  OAI21_X1 U19939 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16864), .A(n16729), 
        .ZN(n16710) );
  NAND2_X1 U19940 ( .A1(n16828), .A2(n16701), .ZN(n16702) );
  OAI22_X1 U19941 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16702), .B1(n17670), 
        .B2(n16857), .ZN(n16709) );
  INV_X1 U19942 ( .A(n17665), .ZN(n16726) );
  NOR2_X1 U19943 ( .A1(n17681), .A2(n16726), .ZN(n16716) );
  OAI21_X1 U19944 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16716), .A(
        n16703), .ZN(n17668) );
  INV_X1 U19945 ( .A(n16861), .ZN(n16704) );
  OAI21_X1 U19946 ( .B1(n16777), .B2(n17670), .A(n16704), .ZN(n16707) );
  NAND3_X1 U19947 ( .A1(n18653), .A2(n17668), .A3(n16705), .ZN(n16706) );
  OAI211_X1 U19948 ( .C1(n17668), .C2(n16707), .A(n18036), .B(n16706), .ZN(
        n16708) );
  AOI211_X1 U19949 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16710), .A(n16709), 
        .B(n16708), .ZN(n16713) );
  OAI211_X1 U19950 ( .C1(n16715), .C2(n16714), .A(n16872), .B(n16711), .ZN(
        n16712) );
  OAI211_X1 U19951 ( .C1(n16714), .C2(n16860), .A(n16713), .B(n16712), .ZN(
        P3_U2658) );
  AOI21_X1 U19952 ( .B1(n16873), .B2(P3_EBX_REG_12__SCAN_IN), .A(n18042), .ZN(
        n16724) );
  AOI211_X1 U19953 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16732), .A(n16715), .B(
        n16863), .ZN(n16722) );
  AOI21_X1 U19954 ( .B1(n17681), .B2(n16726), .A(n16716), .ZN(n17684) );
  XOR2_X1 U19955 ( .A(n17684), .B(n16717), .Z(n16720) );
  NAND2_X1 U19956 ( .A1(n16828), .A2(n18701), .ZN(n16718) );
  OAI22_X1 U19957 ( .A1(n16775), .A2(n16720), .B1(n16719), .B2(n16718), .ZN(
        n16721) );
  AOI211_X1 U19958 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16722), .B(n16721), .ZN(n16723) );
  OAI211_X1 U19959 ( .C1(n18701), .C2(n16729), .A(n16724), .B(n16723), .ZN(
        P3_U2659) );
  INV_X1 U19960 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16736) );
  INV_X1 U19961 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18697) );
  INV_X1 U19962 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18695) );
  NOR2_X1 U19963 ( .A1(n18697), .A2(n18695), .ZN(n16746) );
  NOR3_X1 U19964 ( .A1(n16864), .A2(n16800), .A3(n16725), .ZN(n16757) );
  AOI21_X1 U19965 ( .B1(n16746), .B2(n16757), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16730) );
  INV_X1 U19966 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16771) );
  INV_X1 U19967 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17746) );
  NOR2_X1 U19968 ( .A1(n17691), .A2(n17746), .ZN(n17741) );
  NAND2_X1 U19969 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17741), .ZN(
        n16773) );
  NOR2_X1 U19970 ( .A1(n16771), .A2(n16773), .ZN(n16764) );
  NAND2_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16764), .ZN(
        n16740) );
  NOR2_X1 U19972 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16740), .ZN(
        n16741) );
  AOI21_X1 U19973 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16741), .A(
        n16798), .ZN(n16727) );
  INV_X1 U19974 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17709) );
  NOR2_X1 U19975 ( .A1(n17709), .A2(n16740), .ZN(n16739) );
  OAI21_X1 U19976 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16739), .A(
        n16726), .ZN(n17693) );
  XOR2_X1 U19977 ( .A(n16727), .B(n17693), .Z(n16728) );
  OAI22_X1 U19978 ( .A1(n16730), .A2(n16729), .B1(n16775), .B2(n16728), .ZN(
        n16731) );
  AOI211_X1 U19979 ( .C1(n16873), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18042), .B(
        n16731), .ZN(n16735) );
  OAI211_X1 U19980 ( .C1(n16738), .C2(n16733), .A(n16872), .B(n16732), .ZN(
        n16734) );
  OAI211_X1 U19981 ( .C1(n16857), .C2(n16736), .A(n16735), .B(n16734), .ZN(
        P3_U2660) );
  OAI21_X1 U19982 ( .B1(n16864), .B2(n16737), .A(n16877), .ZN(n16758) );
  INV_X1 U19983 ( .A(n16758), .ZN(n16766) );
  AOI211_X1 U19984 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16759), .A(n16738), .B(
        n16863), .ZN(n16745) );
  AOI21_X1 U19985 ( .B1(n17709), .B2(n16740), .A(n16739), .ZN(n17712) );
  NOR2_X1 U19986 ( .A1(n16741), .A2(n16798), .ZN(n16753) );
  AOI21_X1 U19987 ( .B1(n17712), .B2(n16753), .A(n16775), .ZN(n16742) );
  OAI21_X1 U19988 ( .B1(n17712), .B2(n16753), .A(n16742), .ZN(n16743) );
  OAI211_X1 U19989 ( .C1(n17709), .C2(n16857), .A(n18036), .B(n16743), .ZN(
        n16744) );
  AOI211_X1 U19990 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16873), .A(n16745), .B(
        n16744), .ZN(n16749) );
  INV_X1 U19991 ( .A(n16746), .ZN(n16747) );
  OAI211_X1 U19992 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16757), .B(n16747), .ZN(n16748) );
  OAI211_X1 U19993 ( .C1(n16766), .C2(n18697), .A(n16749), .B(n16748), .ZN(
        P3_U2661) );
  INV_X1 U19994 ( .A(n16764), .ZN(n16750) );
  AOI22_X1 U19995 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16764), .B1(
        n16750), .B2(n17719), .ZN(n17722) );
  INV_X1 U19996 ( .A(n17722), .ZN(n16752) );
  NOR2_X1 U19997 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16750), .ZN(
        n16751) );
  AOI22_X1 U19998 ( .A1(n16753), .A2(n16752), .B1(n16751), .B2(n16859), .ZN(
        n16755) );
  AOI22_X1 U19999 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16851), .B1(
        n16777), .B2(n17722), .ZN(n16754) );
  OAI211_X1 U20000 ( .C1(n16755), .C2(n16775), .A(n16754), .B(n18036), .ZN(
        n16756) );
  AOI221_X1 U20001 ( .B1(n16758), .B2(P3_REIP_REG_9__SCAN_IN), .C1(n16757), 
        .C2(n18695), .A(n16756), .ZN(n16761) );
  OAI211_X1 U20002 ( .C1(n16763), .C2(n16762), .A(n16872), .B(n16759), .ZN(
        n16760) );
  OAI211_X1 U20003 ( .C1(n16762), .C2(n16860), .A(n16761), .B(n16760), .ZN(
        P3_U2662) );
  AOI211_X1 U20004 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16784), .A(n16763), .B(
        n16863), .ZN(n16769) );
  INV_X1 U20005 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18689) );
  NOR3_X1 U20006 ( .A1(n16864), .A2(n16800), .A3(n18689), .ZN(n16783) );
  AOI21_X1 U20007 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16783), .A(
        P3_REIP_REG_8__SCAN_IN), .ZN(n16767) );
  AOI21_X1 U20008 ( .B1(n16771), .B2(n16773), .A(n16764), .ZN(n17732) );
  AOI21_X1 U20009 ( .B1(n17741), .B2(n16853), .A(n16798), .ZN(n16778) );
  XNOR2_X1 U20010 ( .A(n17732), .B(n16778), .ZN(n16765) );
  OAI22_X1 U20011 ( .A1(n16767), .A2(n16766), .B1(n16775), .B2(n16765), .ZN(
        n16768) );
  AOI211_X1 U20012 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16873), .A(n16769), .B(
        n16768), .ZN(n16770) );
  OAI211_X1 U20013 ( .C1(n16771), .C2(n16857), .A(n16770), .B(n18036), .ZN(
        P3_U2663) );
  INV_X1 U20014 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18691) );
  AOI21_X1 U20015 ( .B1(n16828), .B2(n16800), .A(n16868), .ZN(n16810) );
  NOR2_X1 U20016 ( .A1(n16864), .A2(n16800), .ZN(n16772) );
  NAND2_X1 U20017 ( .A1(n16772), .A2(n18689), .ZN(n16792) );
  NAND2_X1 U20018 ( .A1(n16810), .A2(n16792), .ZN(n16782) );
  INV_X1 U20019 ( .A(n16788), .ZN(n16774) );
  OAI21_X1 U20020 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16774), .A(
        n16773), .ZN(n17755) );
  INV_X1 U20021 ( .A(n17755), .ZN(n16779) );
  AOI21_X1 U20022 ( .B1(n16779), .B2(n16790), .A(n16775), .ZN(n16776) );
  OAI22_X1 U20023 ( .A1(n16779), .A2(n16778), .B1(n16777), .B2(n16776), .ZN(
        n16780) );
  OAI211_X1 U20024 ( .C1(n16860), .C2(n17166), .A(n18036), .B(n16780), .ZN(
        n16781) );
  AOI221_X1 U20025 ( .B1(n16783), .B2(n18691), .C1(n16782), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n16781), .ZN(n16786) );
  OAI211_X1 U20026 ( .C1(n16787), .C2(n17166), .A(n16872), .B(n16784), .ZN(
        n16785) );
  OAI211_X1 U20027 ( .C1(n16857), .C2(n17746), .A(n16786), .B(n16785), .ZN(
        P3_U2664) );
  AOI211_X1 U20028 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16803), .A(n16787), .B(
        n16863), .ZN(n16796) );
  NAND2_X1 U20029 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17768), .ZN(
        n16799) );
  INV_X1 U20030 ( .A(n16799), .ZN(n16789) );
  OAI21_X1 U20031 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16789), .A(
        n16788), .ZN(n17771) );
  NAND2_X1 U20032 ( .A1(n17771), .A2(n16790), .ZN(n16794) );
  AOI211_X1 U20033 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16818), .A(
        n17771), .B(n16861), .ZN(n16791) );
  AOI211_X1 U20034 ( .C1(n16873), .C2(P3_EBX_REG_6__SCAN_IN), .A(n18042), .B(
        n16791), .ZN(n16793) );
  OAI211_X1 U20035 ( .C1(n16858), .C2(n16794), .A(n16793), .B(n16792), .ZN(
        n16795) );
  AOI211_X1 U20036 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16796), .B(n16795), .ZN(n16797) );
  OAI21_X1 U20037 ( .B1(n16810), .B2(n18689), .A(n16797), .ZN(P3_U2665) );
  INV_X1 U20038 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18688) );
  NOR2_X1 U20039 ( .A1(n17825), .A2(n17777), .ZN(n16814) );
  AOI21_X1 U20040 ( .B1(n16814), .B2(n16859), .A(n16798), .ZN(n16820) );
  OAI21_X1 U20041 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16814), .A(
        n16799), .ZN(n17782) );
  XNOR2_X1 U20042 ( .A(n16820), .B(n17782), .ZN(n16808) );
  AND2_X1 U20043 ( .A1(n16800), .A2(n16828), .ZN(n16801) );
  AOI22_X1 U20044 ( .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n16851), .B1(
        n16802), .B2(n16801), .ZN(n16805) );
  OAI211_X1 U20045 ( .C1(n16811), .C2(n16806), .A(n16872), .B(n16803), .ZN(
        n16804) );
  OAI211_X1 U20046 ( .C1(n16806), .C2(n16860), .A(n16805), .B(n16804), .ZN(
        n16807) );
  AOI211_X1 U20047 ( .C1(n18653), .C2(n16808), .A(n18042), .B(n16807), .ZN(
        n16809) );
  OAI21_X1 U20048 ( .B1(n16810), .B2(n18688), .A(n16809), .ZN(P3_U2666) );
  AOI21_X1 U20049 ( .B1(n16828), .B2(n16813), .A(n16868), .ZN(n16835) );
  NOR2_X1 U20050 ( .A1(n18157), .A2(n18819), .ZN(n16875) );
  AOI211_X1 U20051 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16838), .A(n16811), .B(
        n16863), .ZN(n16812) );
  AOI221_X1 U20052 ( .B1(n17082), .B2(n16875), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n16875), .A(n16812), .ZN(
        n16827) );
  NOR3_X1 U20053 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16864), .A3(n16813), .ZN(
        n16825) );
  INV_X1 U20054 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16816) );
  NAND2_X1 U20055 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17792), .ZN(
        n16830) );
  AOI21_X1 U20056 ( .B1(n16816), .B2(n16830), .A(n16814), .ZN(n16815) );
  INV_X1 U20057 ( .A(n16815), .ZN(n17795) );
  INV_X1 U20058 ( .A(n16853), .ZN(n16817) );
  NAND2_X1 U20059 ( .A1(n17792), .A2(n16816), .ZN(n17786) );
  OAI22_X1 U20060 ( .A1(n16818), .A2(n17795), .B1(n16817), .B2(n17786), .ZN(
        n16819) );
  AOI211_X1 U20061 ( .C1(n16820), .C2(n17795), .A(n18042), .B(n16819), .ZN(
        n16822) );
  OAI22_X1 U20062 ( .A1(n16823), .A2(n16822), .B1(n16860), .B2(n16821), .ZN(
        n16824) );
  AOI211_X1 U20063 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16825), .B(n16824), .ZN(n16826) );
  OAI211_X1 U20064 ( .C1(n18685), .C2(n16835), .A(n16827), .B(n16826), .ZN(
        P3_U2667) );
  INV_X1 U20065 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18683) );
  INV_X1 U20066 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18681) );
  NOR2_X1 U20067 ( .A1(n18791), .A2(n18681), .ZN(n16845) );
  AND3_X1 U20068 ( .A1(n18683), .A2(n16828), .A3(n16845), .ZN(n16837) );
  NOR2_X1 U20069 ( .A1(n11412), .A2(n18782), .ZN(n18602) );
  NAND2_X1 U20070 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18602), .ZN(
        n18597) );
  AOI21_X1 U20071 ( .B1(n18597), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17077), .ZN(n16829) );
  INV_X1 U20072 ( .A(n16829), .ZN(n18761) );
  AOI21_X1 U20073 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16853), .A(
        n16858), .ZN(n16852) );
  NOR2_X1 U20074 ( .A1(n17825), .A2(n17816), .ZN(n16831) );
  OAI21_X1 U20075 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16831), .A(
        n16830), .ZN(n17806) );
  AOI22_X1 U20076 ( .A1(n16875), .A2(n18761), .B1(n16852), .B2(n17806), .ZN(
        n16834) );
  INV_X1 U20077 ( .A(n16831), .ZN(n16843) );
  AOI211_X1 U20078 ( .C1(n16843), .C2(n16844), .A(n17806), .B(n16861), .ZN(
        n16832) );
  INV_X1 U20079 ( .A(n16832), .ZN(n16833) );
  OAI211_X1 U20080 ( .C1(n16835), .C2(n18683), .A(n16834), .B(n16833), .ZN(
        n16836) );
  AOI211_X1 U20081 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16837), .B(n16836), .ZN(n16840) );
  OAI211_X1 U20082 ( .C1(n16842), .C2(n16841), .A(n16872), .B(n16838), .ZN(
        n16839) );
  OAI211_X1 U20083 ( .C1(n16841), .C2(n16860), .A(n16840), .B(n16839), .ZN(
        P3_U2668) );
  INV_X1 U20084 ( .A(n16875), .ZN(n16871) );
  NAND2_X1 U20085 ( .A1(n11412), .A2(n18601), .ZN(n18595) );
  NAND2_X1 U20086 ( .A1(n18597), .A2(n18595), .ZN(n18769) );
  INV_X1 U20087 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17199) );
  INV_X1 U20088 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17193) );
  NAND2_X1 U20089 ( .A1(n17199), .A2(n17193), .ZN(n16862) );
  AOI211_X1 U20090 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16862), .A(n16842), .B(
        n16863), .ZN(n16850) );
  OAI21_X1 U20091 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16843), .ZN(n17812) );
  OAI22_X1 U20092 ( .A1(n16877), .A2(n18681), .B1(n17812), .B2(n16844), .ZN(
        n16847) );
  AOI211_X1 U20093 ( .C1(n18791), .C2(n18681), .A(n16864), .B(n16845), .ZN(
        n16846) );
  AOI211_X1 U20094 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16873), .A(n16847), .B(
        n16846), .ZN(n16848) );
  INV_X1 U20095 ( .A(n16848), .ZN(n16849) );
  AOI211_X1 U20096 ( .C1(n16851), .C2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n16850), .B(n16849), .ZN(n16855) );
  OAI21_X1 U20097 ( .B1(n16853), .B2(n17812), .A(n16852), .ZN(n16854) );
  OAI211_X1 U20098 ( .C1(n16871), .C2(n18769), .A(n16855), .B(n16854), .ZN(
        P3_U2669) );
  NAND2_X1 U20099 ( .A1(n18601), .A2(n16856), .ZN(n18775) );
  OAI21_X1 U20100 ( .B1(n16859), .B2(n16858), .A(n16857), .ZN(n16867) );
  OAI22_X1 U20101 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16861), .B1(
        n17193), .B2(n16860), .ZN(n16866) );
  NAND2_X1 U20102 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17185) );
  NAND2_X1 U20103 ( .A1(n16862), .A2(n17185), .ZN(n17195) );
  OAI22_X1 U20104 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16864), .B1(n16863), 
        .B2(n17195), .ZN(n16865) );
  AOI211_X1 U20105 ( .C1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n16867), .A(
        n16866), .B(n16865), .ZN(n16870) );
  NAND2_X1 U20106 ( .A1(n16868), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n16869) );
  OAI211_X1 U20107 ( .C1(n16871), .C2(n18775), .A(n16870), .B(n16869), .ZN(
        P3_U2670) );
  NOR2_X1 U20108 ( .A1(n16873), .A2(n16872), .ZN(n16880) );
  INV_X1 U20109 ( .A(n16874), .ZN(n16876) );
  AOI22_X1 U20110 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16876), .B1(n16875), 
        .B2(n18789), .ZN(n16879) );
  NAND3_X1 U20111 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18771), .A3(
        n16877), .ZN(n16878) );
  OAI211_X1 U20112 ( .C1(n16880), .C2(n17199), .A(n16879), .B(n16878), .ZN(
        P3_U2671) );
  NAND4_X1 U20113 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16881)
         );
  NOR3_X1 U20114 ( .A1(n16916), .A2(n16882), .A3(n16881), .ZN(n16883) );
  NAND4_X1 U20115 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16972), .A3(n16917), 
        .A4(n16883), .ZN(n16908) );
  NOR2_X1 U20116 ( .A1(n16909), .A2(n16908), .ZN(n16907) );
  NAND2_X1 U20117 ( .A1(n17191), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16885) );
  NAND2_X1 U20118 ( .A1(n16907), .A2(n16989), .ZN(n16884) );
  OAI22_X1 U20119 ( .A1(n16907), .A2(n16885), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16884), .ZN(P3_U2672) );
  AOI22_X1 U20120 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20121 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17149), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20122 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17082), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20123 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17132), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17152), .ZN(n16886) );
  NAND4_X1 U20124 ( .A1(n16889), .A2(n16888), .A3(n16887), .A4(n16886), .ZN(
        n16895) );
  AOI22_X1 U20125 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17143), .ZN(n16893) );
  AOI22_X1 U20126 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17141), .ZN(n16892) );
  AOI22_X1 U20127 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17150), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17109), .ZN(n16891) );
  AOI22_X1 U20128 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17116), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16890) );
  NAND4_X1 U20129 ( .A1(n16893), .A2(n16892), .A3(n16891), .A4(n16890), .ZN(
        n16894) );
  NOR2_X1 U20130 ( .A1(n16895), .A2(n16894), .ZN(n16906) );
  AOI22_X1 U20131 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20132 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16898) );
  AOI22_X1 U20133 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16897) );
  AOI22_X1 U20134 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16896) );
  NAND4_X1 U20135 ( .A1(n16899), .A2(n16898), .A3(n16897), .A4(n16896), .ZN(
        n16905) );
  AOI22_X1 U20136 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20137 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20138 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20139 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16900) );
  NAND4_X1 U20140 ( .A1(n16903), .A2(n16902), .A3(n16901), .A4(n16900), .ZN(
        n16904) );
  NOR2_X1 U20141 ( .A1(n16905), .A2(n16904), .ZN(n16914) );
  NOR2_X1 U20142 ( .A1(n16914), .A2(n16913), .ZN(n16912) );
  XNOR2_X1 U20143 ( .A(n16906), .B(n16912), .ZN(n17207) );
  AOI211_X1 U20144 ( .C1(n16909), .C2(n16908), .A(n16907), .B(n17197), .ZN(
        n16910) );
  AOI21_X1 U20145 ( .B1(n17197), .B2(n17207), .A(n16910), .ZN(n16911) );
  INV_X1 U20146 ( .A(n16911), .ZN(P3_U2673) );
  AOI21_X1 U20147 ( .B1(n16914), .B2(n16913), .A(n16912), .ZN(n17214) );
  AOI22_X1 U20148 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16915), .B1(n17214), 
        .B2(n17197), .ZN(n16919) );
  NAND4_X1 U20149 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16935), .A3(n16917), 
        .A4(n16916), .ZN(n16918) );
  NAND2_X1 U20150 ( .A1(n16919), .A2(n16918), .ZN(P3_U2674) );
  AOI21_X1 U20151 ( .B1(n16921), .B2(n16926), .A(n16920), .ZN(n17224) );
  NAND2_X1 U20152 ( .A1(n17224), .A2(n17197), .ZN(n16922) );
  OAI221_X1 U20153 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16925), .C1(n16924), 
        .C2(n16923), .A(n16922), .ZN(P3_U2676) );
  INV_X1 U20154 ( .A(n16925), .ZN(n16929) );
  AOI21_X1 U20155 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17191), .A(n16935), .ZN(
        n16928) );
  OAI21_X1 U20156 ( .B1(n16931), .B2(n16927), .A(n16926), .ZN(n17230) );
  OAI22_X1 U20157 ( .A1(n16929), .A2(n16928), .B1(n17191), .B2(n17230), .ZN(
        P3_U2677) );
  INV_X1 U20158 ( .A(n16930), .ZN(n16939) );
  AOI21_X1 U20159 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17191), .A(n16939), .ZN(
        n16934) );
  AOI21_X1 U20160 ( .B1(n16932), .B2(n16936), .A(n16931), .ZN(n17231) );
  INV_X1 U20161 ( .A(n17231), .ZN(n16933) );
  OAI22_X1 U20162 ( .A1(n16935), .A2(n16934), .B1(n17191), .B2(n16933), .ZN(
        P3_U2678) );
  AOI21_X1 U20163 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17191), .A(n16946), .ZN(
        n16938) );
  OAI21_X1 U20164 ( .B1(n16941), .B2(n16937), .A(n16936), .ZN(n17240) );
  OAI22_X1 U20165 ( .A1(n16939), .A2(n16938), .B1(n17191), .B2(n17240), .ZN(
        P3_U2679) );
  INV_X1 U20166 ( .A(n16940), .ZN(n16961) );
  AOI21_X1 U20167 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17191), .A(n16961), .ZN(
        n16945) );
  AOI21_X1 U20168 ( .B1(n16943), .B2(n16942), .A(n16941), .ZN(n17241) );
  INV_X1 U20169 ( .A(n17241), .ZN(n16944) );
  OAI22_X1 U20170 ( .A1(n16946), .A2(n16945), .B1(n17191), .B2(n16944), .ZN(
        P3_U2680) );
  AOI21_X1 U20171 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17191), .A(n16947), .ZN(
        n16960) );
  AOI22_X1 U20172 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16958) );
  INV_X1 U20173 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16950) );
  AOI22_X1 U20174 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16949) );
  AOI22_X1 U20175 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16948) );
  OAI211_X1 U20176 ( .C1(n11237), .C2(n16950), .A(n16949), .B(n16948), .ZN(
        n16956) );
  AOI22_X1 U20177 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16954) );
  AOI22_X1 U20178 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20179 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16952) );
  AOI22_X1 U20180 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16951) );
  NAND4_X1 U20181 ( .A1(n16954), .A2(n16953), .A3(n16952), .A4(n16951), .ZN(
        n16955) );
  AOI211_X1 U20182 ( .C1(n17152), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n16956), .B(n16955), .ZN(n16957) );
  NAND2_X1 U20183 ( .A1(n16958), .A2(n16957), .ZN(n17246) );
  INV_X1 U20184 ( .A(n17246), .ZN(n16959) );
  OAI22_X1 U20185 ( .A1(n16961), .A2(n16960), .B1(n16959), .B2(n17191), .ZN(
        P3_U2681) );
  AOI22_X1 U20186 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20187 ( .A1(n17141), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20188 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16963) );
  AOI22_X1 U20189 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16962) );
  NAND4_X1 U20190 ( .A1(n16965), .A2(n16964), .A3(n16963), .A4(n16962), .ZN(
        n16971) );
  AOI22_X1 U20191 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20192 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20193 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16967) );
  AOI22_X1 U20194 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16966) );
  NAND4_X1 U20195 ( .A1(n16969), .A2(n16968), .A3(n16967), .A4(n16966), .ZN(
        n16970) );
  NOR2_X1 U20196 ( .A1(n16971), .A2(n16970), .ZN(n17253) );
  INV_X1 U20197 ( .A(n17253), .ZN(n16975) );
  OAI21_X1 U20198 ( .B1(n16973), .B2(n16972), .A(n17191), .ZN(n16974) );
  OAI21_X1 U20199 ( .B1(n17191), .B2(n16975), .A(n16974), .ZN(n16976) );
  OAI21_X1 U20200 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16977), .A(n16976), .ZN(
        P3_U2682) );
  AOI22_X1 U20201 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20202 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20203 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16979) );
  AOI22_X1 U20204 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16978) );
  NAND4_X1 U20205 ( .A1(n16981), .A2(n16980), .A3(n16979), .A4(n16978), .ZN(
        n16987) );
  AOI22_X1 U20206 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20207 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16984) );
  AOI22_X1 U20208 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16983) );
  AOI22_X1 U20209 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16982) );
  NAND4_X1 U20210 ( .A1(n16985), .A2(n16984), .A3(n16983), .A4(n16982), .ZN(
        n16986) );
  NOR2_X1 U20211 ( .A1(n16987), .A2(n16986), .ZN(n17260) );
  NAND3_X1 U20212 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17191), .A3(n17003), 
        .ZN(n16991) );
  NAND4_X1 U20213 ( .A1(n16989), .A2(P3_EBX_REG_19__SCAN_IN), .A3(n17002), 
        .A4(n16988), .ZN(n16990) );
  OAI211_X1 U20214 ( .C1(n17260), .C2(n17191), .A(n16991), .B(n16990), .ZN(
        P3_U2683) );
  AOI22_X1 U20215 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20216 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20217 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20218 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16992) );
  NAND4_X1 U20219 ( .A1(n16995), .A2(n16994), .A3(n16993), .A4(n16992), .ZN(
        n17001) );
  AOI22_X1 U20220 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20221 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20222 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20223 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16996) );
  NAND4_X1 U20224 ( .A1(n16999), .A2(n16998), .A3(n16997), .A4(n16996), .ZN(
        n17000) );
  NOR2_X1 U20225 ( .A1(n17001), .A2(n17000), .ZN(n17265) );
  NOR2_X1 U20226 ( .A1(n17002), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n17005) );
  NAND2_X1 U20227 ( .A1(n17191), .A2(n17003), .ZN(n17004) );
  OAI22_X1 U20228 ( .A1(n17265), .A2(n17191), .B1(n17005), .B2(n17004), .ZN(
        P3_U2684) );
  NAND2_X1 U20229 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17006), .ZN(n17019) );
  AOI22_X1 U20230 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20231 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20232 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20233 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17007) );
  NAND4_X1 U20234 ( .A1(n17010), .A2(n17009), .A3(n17008), .A4(n17007), .ZN(
        n17016) );
  AOI22_X1 U20235 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20236 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20237 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20238 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20239 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  NOR2_X1 U20240 ( .A1(n17016), .A2(n17015), .ZN(n17269) );
  INV_X1 U20241 ( .A(n17194), .ZN(n17196) );
  NAND4_X1 U20242 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17031), .A3(n17196), 
        .A4(n17017), .ZN(n17018) );
  OAI221_X1 U20243 ( .B1(n17197), .B2(n17019), .C1(n17191), .C2(n17269), .A(
        n17018), .ZN(P3_U2685) );
  AOI22_X1 U20244 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20245 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20246 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20247 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17020) );
  NAND4_X1 U20248 ( .A1(n17023), .A2(n17022), .A3(n17021), .A4(n17020), .ZN(
        n17030) );
  AOI22_X1 U20249 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20250 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20251 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20252 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17025) );
  NAND4_X1 U20253 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17029) );
  NOR2_X1 U20254 ( .A1(n17030), .A2(n17029), .ZN(n17275) );
  AND2_X1 U20255 ( .A1(n17031), .A2(n17196), .ZN(n17033) );
  NOR2_X1 U20256 ( .A1(n18188), .A2(n17031), .ZN(n17035) );
  NAND2_X1 U20257 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17200), .ZN(n17032) );
  OAI22_X1 U20258 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17033), .B1(n17035), 
        .B2(n17032), .ZN(n17034) );
  OAI21_X1 U20259 ( .B1(n17275), .B2(n17191), .A(n17034), .ZN(P3_U2686) );
  INV_X1 U20260 ( .A(n17035), .ZN(n17048) );
  NAND3_X1 U20261 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17049), .A3(n17105), 
        .ZN(n17047) );
  AOI22_X1 U20262 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20263 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20264 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20265 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20266 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17045) );
  AOI22_X1 U20267 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20268 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20269 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20270 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17040) );
  NAND4_X1 U20271 ( .A1(n17043), .A2(n17042), .A3(n17041), .A4(n17040), .ZN(
        n17044) );
  NOR2_X1 U20272 ( .A1(n17045), .A2(n17044), .ZN(n17281) );
  NAND2_X1 U20273 ( .A1(n17191), .A2(n17047), .ZN(n17061) );
  OAI222_X1 U20274 ( .A1(n17048), .A2(n17047), .B1(n17191), .B2(n17281), .C1(
        n17046), .C2(n17061), .ZN(P3_U2687) );
  AOI21_X1 U20275 ( .B1(n17049), .B2(n17105), .A(P3_EBX_REG_15__SCAN_IN), .ZN(
        n17062) );
  AOI22_X1 U20276 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17109), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17150), .ZN(n17054) );
  AOI22_X1 U20277 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17143), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20278 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20279 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17051) );
  NAND4_X1 U20280 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n17051), .ZN(
        n17060) );
  AOI22_X1 U20281 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20282 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17149), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17141), .ZN(n17057) );
  AOI22_X1 U20283 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17142), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n17124), .ZN(n17056) );
  AOI22_X1 U20284 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17152), .B1(
        n17132), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17055) );
  NAND4_X1 U20285 ( .A1(n17058), .A2(n17057), .A3(n17056), .A4(n17055), .ZN(
        n17059) );
  NOR2_X1 U20286 ( .A1(n17060), .A2(n17059), .ZN(n17286) );
  OAI22_X1 U20287 ( .A1(n17062), .A2(n17061), .B1(n17286), .B2(n17191), .ZN(
        P3_U2688) );
  NAND2_X1 U20288 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17063), .ZN(n17076) );
  AOI22_X1 U20289 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20290 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20291 ( .A1(n17064), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20292 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17065) );
  NAND4_X1 U20293 ( .A1(n17068), .A2(n17067), .A3(n17066), .A4(n17065), .ZN(
        n17074) );
  AOI22_X1 U20294 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20295 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20296 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20297 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17069) );
  NAND4_X1 U20298 ( .A1(n17072), .A2(n17071), .A3(n17070), .A4(n17069), .ZN(
        n17073) );
  NOR2_X1 U20299 ( .A1(n17074), .A2(n17073), .ZN(n17291) );
  NAND3_X1 U20300 ( .A1(n17076), .A2(P3_EBX_REG_14__SCAN_IN), .A3(n17191), 
        .ZN(n17075) );
  OAI221_X1 U20301 ( .B1(n17076), .B2(P3_EBX_REG_14__SCAN_IN), .C1(n17191), 
        .C2(n17291), .A(n17075), .ZN(P3_U2689) );
  AOI22_X1 U20302 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20303 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17077), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20304 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20305 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17078) );
  NAND4_X1 U20306 ( .A1(n17081), .A2(n17080), .A3(n17079), .A4(n17078), .ZN(
        n17088) );
  AOI22_X1 U20307 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20308 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20309 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17082), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20310 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17083) );
  NAND4_X1 U20311 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17087) );
  NOR2_X1 U20312 ( .A1(n17088), .A2(n17087), .ZN(n17296) );
  INV_X1 U20313 ( .A(n17089), .ZN(n17091) );
  OAI21_X1 U20314 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17091), .A(n17090), .ZN(
        n17092) );
  OAI21_X1 U20315 ( .B1(n17296), .B2(n17191), .A(n17092), .ZN(P3_U2691) );
  AOI22_X1 U20316 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20317 ( .A1(n17116), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20318 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20319 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17093) );
  NAND4_X1 U20320 ( .A1(n17096), .A2(n17095), .A3(n17094), .A4(n17093), .ZN(
        n17102) );
  AOI22_X1 U20321 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20322 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20323 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17098) );
  AOI22_X1 U20324 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17097) );
  NAND4_X1 U20325 ( .A1(n17100), .A2(n17099), .A3(n17098), .A4(n17097), .ZN(
        n17101) );
  NOR2_X1 U20326 ( .A1(n17102), .A2(n17101), .ZN(n17300) );
  NAND2_X1 U20327 ( .A1(n17191), .A2(n17103), .ZN(n17120) );
  NOR2_X1 U20328 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17120), .ZN(n17104) );
  AOI221_X1 U20329 ( .B1(n17300), .B2(n17197), .C1(n17105), .C2(n17191), .A(
        n17104), .ZN(P3_U2692) );
  AOI22_X1 U20330 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20331 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17118) );
  AOI22_X1 U20332 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17106) );
  OAI21_X1 U20333 ( .B1(n17108), .B2(n17107), .A(n17106), .ZN(n17115) );
  AOI22_X1 U20334 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20335 ( .A1(n17109), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20336 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20337 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17110) );
  NAND4_X1 U20338 ( .A1(n17113), .A2(n17112), .A3(n17111), .A4(n17110), .ZN(
        n17114) );
  AOI211_X1 U20339 ( .C1(n17116), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17115), .B(n17114), .ZN(n17117) );
  NAND3_X1 U20340 ( .A1(n17119), .A2(n17118), .A3(n17117), .ZN(n17304) );
  INV_X1 U20341 ( .A(n17304), .ZN(n17122) );
  NOR2_X1 U20342 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17140), .ZN(n17121) );
  OAI22_X1 U20343 ( .A1(n17122), .A2(n17191), .B1(n17121), .B2(n17120), .ZN(
        P3_U2693) );
  INV_X1 U20344 ( .A(n17162), .ZN(n17123) );
  OAI21_X1 U20345 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17123), .A(n17191), .ZN(
        n17139) );
  AOI22_X1 U20346 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20347 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17116), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20348 ( .A1(n17082), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20349 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20350 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17138) );
  AOI22_X1 U20351 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17129), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20352 ( .A1(n17131), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20353 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20354 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17133) );
  NAND4_X1 U20355 ( .A1(n17136), .A2(n17135), .A3(n17134), .A4(n17133), .ZN(
        n17137) );
  NOR2_X1 U20356 ( .A1(n17138), .A2(n17137), .ZN(n17309) );
  OAI22_X1 U20357 ( .A1(n17140), .A2(n17139), .B1(n17309), .B2(n17191), .ZN(
        P3_U2694) );
  AOI22_X1 U20358 ( .A1(n17142), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17141), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20359 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17160) );
  AOI22_X1 U20360 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17109), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17145) );
  OAI21_X1 U20361 ( .B1(n17147), .B2(n17146), .A(n17145), .ZN(n17158) );
  AOI22_X1 U20362 ( .A1(n17130), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17148), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20363 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20364 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17150), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20365 ( .A1(n17132), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17153) );
  NAND4_X1 U20366 ( .A1(n17156), .A2(n17155), .A3(n17154), .A4(n17153), .ZN(
        n17157) );
  AOI211_X1 U20367 ( .C1(n17082), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17158), .B(n17157), .ZN(n17159) );
  NAND3_X1 U20368 ( .A1(n17161), .A2(n17160), .A3(n17159), .ZN(n17315) );
  INV_X1 U20369 ( .A(n17315), .ZN(n17164) );
  OAI21_X1 U20370 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17165), .A(n17162), .ZN(
        n17163) );
  AOI22_X1 U20371 ( .A1(n17197), .A2(n17164), .B1(n17163), .B2(n17191), .ZN(
        P3_U2695) );
  OR2_X1 U20372 ( .A1(n17166), .A2(n17165), .ZN(n17169) );
  NOR2_X1 U20373 ( .A1(n18188), .A2(n17170), .ZN(n17171) );
  NAND3_X1 U20374 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17171), .A3(n17166), .ZN(
        n17167) );
  OAI221_X1 U20375 ( .B1(n17197), .B2(n17169), .C1(n17191), .C2(n17168), .A(
        n17167), .ZN(P3_U2696) );
  NAND2_X1 U20376 ( .A1(n17191), .A2(n17170), .ZN(n17175) );
  AOI22_X1 U20377 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17197), .B1(
        n17171), .B2(n17173), .ZN(n17172) );
  OAI21_X1 U20378 ( .B1(n17173), .B2(n17175), .A(n17172), .ZN(P3_U2697) );
  NOR2_X1 U20379 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17181), .ZN(n17176) );
  INV_X1 U20380 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17174) );
  OAI22_X1 U20381 ( .A1(n17176), .A2(n17175), .B1(n17174), .B2(n17191), .ZN(
        P3_U2698) );
  INV_X1 U20382 ( .A(n17177), .ZN(n17178) );
  OAI21_X1 U20383 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17178), .A(n17191), .ZN(
        n17180) );
  INV_X1 U20384 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17179) );
  OAI22_X1 U20385 ( .A1(n17181), .A2(n17180), .B1(n17179), .B2(n17191), .ZN(
        P3_U2699) );
  OR2_X1 U20386 ( .A1(n17187), .A2(n17194), .ZN(n17184) );
  INV_X1 U20387 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17183) );
  NAND3_X1 U20388 ( .A1(n17184), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17191), .ZN(
        n17182) );
  OAI221_X1 U20389 ( .B1(n17184), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17191), 
        .C2(n17183), .A(n17182), .ZN(P3_U2700) );
  INV_X1 U20390 ( .A(n17185), .ZN(n17186) );
  AOI21_X1 U20391 ( .B1(n17200), .B2(n17186), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17190) );
  OAI21_X1 U20392 ( .B1(n17187), .B2(n17194), .A(n17191), .ZN(n17189) );
  INV_X1 U20393 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17188) );
  OAI22_X1 U20394 ( .A1(n17190), .A2(n17189), .B1(n17188), .B2(n17191), .ZN(
        P3_U2701) );
  OAI222_X1 U20395 ( .A1(n17195), .A2(n17194), .B1(n17193), .B2(n17200), .C1(
        n17192), .C2(n17191), .ZN(P3_U2702) );
  AOI22_X1 U20396 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17197), .B1(
        n17196), .B2(n17199), .ZN(n17198) );
  OAI21_X1 U20397 ( .B1(n17200), .B2(n17199), .A(n17198), .ZN(P3_U2703) );
  INV_X1 U20398 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17353) );
  INV_X1 U20399 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17357) );
  INV_X1 U20400 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17361) );
  INV_X1 U20401 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17367) );
  INV_X1 U20402 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17464) );
  NAND2_X1 U20403 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17344) );
  INV_X1 U20404 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17401) );
  INV_X1 U20405 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17403) );
  NAND4_X1 U20406 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17201) );
  NOR4_X1 U20407 ( .A1(n17344), .A2(n17401), .A3(n17403), .A4(n17201), .ZN(
        n17313) );
  INV_X1 U20408 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17395) );
  INV_X1 U20409 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17385) );
  INV_X1 U20410 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17391) );
  INV_X1 U20411 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17393) );
  NAND2_X1 U20412 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(P3_EAX_REG_11__SCAN_IN), 
        .ZN(n17292) );
  NOR4_X1 U20413 ( .A1(n17385), .A2(n17391), .A3(n17393), .A4(n17292), .ZN(
        n17287) );
  NAND4_X1 U20414 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17313), .A3(n17312), 
        .A4(n17287), .ZN(n17288) );
  INV_X1 U20415 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17369) );
  INV_X1 U20416 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17371) );
  NOR2_X1 U20417 ( .A1(n17369), .A2(n17371), .ZN(n17202) );
  NAND4_X1 U20418 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .A4(n17202), .ZN(n17251) );
  NAND2_X1 U20419 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17243), .ZN(n17242) );
  NOR2_X2 U20420 ( .A1(n18188), .A2(n17242), .ZN(n17237) );
  NOR2_X2 U20421 ( .A1(n17361), .A2(n17236), .ZN(n17232) );
  NAND2_X1 U20422 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17232), .ZN(n17227) );
  NAND2_X1 U20423 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17221), .ZN(n17217) );
  NOR2_X2 U20424 ( .A1(n17353), .A2(n17217), .ZN(n17208) );
  NAND2_X1 U20425 ( .A1(n17208), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17206) );
  NOR2_X2 U20426 ( .A1(n17203), .A2(n17337), .ZN(n17276) );
  INV_X1 U20427 ( .A(n17208), .ZN(n17213) );
  NAND2_X1 U20428 ( .A1(n17337), .A2(n17213), .ZN(n17211) );
  OAI21_X1 U20429 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17335), .A(n17211), .ZN(
        n17204) );
  AOI22_X1 U20430 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17276), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17204), .ZN(n17205) );
  OAI21_X1 U20431 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17206), .A(n17205), .ZN(
        P3_U2704) );
  INV_X1 U20432 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20433 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n17276), .B1(n17316), .B2(
        n17207), .ZN(n17210) );
  NOR2_X2 U20434 ( .A1(n18180), .A2(n17337), .ZN(n17277) );
  AOI22_X1 U20435 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17277), .B1(n17208), .B2(
        n17433), .ZN(n17209) );
  OAI211_X1 U20436 ( .C1(n17211), .C2(n17433), .A(n17210), .B(n17209), .ZN(
        P3_U2705) );
  OAI21_X1 U20437 ( .B1(n17283), .B2(n17353), .A(n17217), .ZN(n17212) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n17276), .B1(n17213), .B2(
        n17212), .ZN(n17216) );
  AOI22_X1 U20439 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17277), .B1(n17316), .B2(
        n17214), .ZN(n17215) );
  NAND2_X1 U20440 ( .A1(n17216), .A2(n17215), .ZN(P3_U2706) );
  AOI22_X1 U20441 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17276), .ZN(n17219) );
  OAI211_X1 U20442 ( .C1(n17221), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17337), .B(
        n17217), .ZN(n17218) );
  OAI211_X1 U20443 ( .C1(n17220), .C2(n17348), .A(n17219), .B(n17218), .ZN(
        P3_U2707) );
  INV_X1 U20444 ( .A(n17221), .ZN(n17223) );
  OAI21_X1 U20445 ( .B1(n17283), .B2(n17357), .A(n17227), .ZN(n17222) );
  AOI22_X1 U20446 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17276), .B1(n17223), .B2(
        n17222), .ZN(n17226) );
  AOI22_X1 U20447 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17277), .B1(n17316), .B2(
        n17224), .ZN(n17225) );
  NAND2_X1 U20448 ( .A1(n17226), .A2(n17225), .ZN(P3_U2708) );
  AOI22_X1 U20449 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17276), .ZN(n17229) );
  OAI211_X1 U20450 ( .C1(n17232), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17337), .B(
        n17227), .ZN(n17228) );
  OAI211_X1 U20451 ( .C1(n17230), .C2(n17348), .A(n17229), .B(n17228), .ZN(
        P3_U2709) );
  INV_X1 U20452 ( .A(n17276), .ZN(n17252) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17277), .B1(n17316), .B2(
        n17231), .ZN(n17235) );
  AOI211_X1 U20454 ( .C1(n17361), .C2(n17236), .A(n17232), .B(n17283), .ZN(
        n17233) );
  INV_X1 U20455 ( .A(n17233), .ZN(n17234) );
  OAI211_X1 U20456 ( .C1(n17252), .C2(n14843), .A(n17235), .B(n17234), .ZN(
        P3_U2710) );
  AOI22_X1 U20457 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17276), .ZN(n17239) );
  OAI211_X1 U20458 ( .C1(n17237), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17337), .B(
        n17236), .ZN(n17238) );
  OAI211_X1 U20459 ( .C1(n17240), .C2(n17348), .A(n17239), .B(n17238), .ZN(
        P3_U2711) );
  AOI22_X1 U20460 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17277), .B1(n17316), .B2(
        n17241), .ZN(n17245) );
  OAI211_X1 U20461 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17243), .A(n17337), .B(
        n17242), .ZN(n17244) );
  OAI211_X1 U20462 ( .C1(n17252), .C2(n14866), .A(n17245), .B(n17244), .ZN(
        P3_U2712) );
  NOR2_X1 U20463 ( .A1(n18188), .A2(n17278), .ZN(n17272) );
  NAND2_X1 U20464 ( .A1(n17272), .A2(n17367), .ZN(n17250) );
  AOI22_X1 U20465 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17276), .B1(n17316), .B2(
        n17246), .ZN(n17249) );
  INV_X1 U20466 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17373) );
  INV_X1 U20467 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17419) );
  NAND2_X1 U20468 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17270), .ZN(n17266) );
  NAND2_X1 U20469 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17261), .ZN(n17257) );
  NAND2_X1 U20470 ( .A1(n17337), .A2(n17257), .ZN(n17256) );
  OAI21_X1 U20471 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17335), .A(n17256), .ZN(
        n17247) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17277), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17247), .ZN(n17248) );
  OAI211_X1 U20473 ( .C1(n17251), .C2(n17250), .A(n17249), .B(n17248), .ZN(
        P3_U2713) );
  OAI22_X1 U20474 ( .A1(n17253), .A2(n17348), .B1(n14875), .B2(n17252), .ZN(
        n17254) );
  AOI21_X1 U20475 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17277), .A(n17254), .ZN(
        n17255) );
  OAI221_X1 U20476 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17257), .C1(n17369), 
        .C2(n17256), .A(n17255), .ZN(P3_U2714) );
  AOI22_X1 U20477 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17276), .ZN(n17259) );
  OAI211_X1 U20478 ( .C1(n17261), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17337), .B(
        n17257), .ZN(n17258) );
  OAI211_X1 U20479 ( .C1(n17260), .C2(n17348), .A(n17259), .B(n17258), .ZN(
        P3_U2715) );
  AOI22_X1 U20480 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17276), .ZN(n17264) );
  AOI211_X1 U20481 ( .C1(n17373), .C2(n17266), .A(n17261), .B(n17283), .ZN(
        n17262) );
  INV_X1 U20482 ( .A(n17262), .ZN(n17263) );
  OAI211_X1 U20483 ( .C1(n17265), .C2(n17348), .A(n17264), .B(n17263), .ZN(
        P3_U2716) );
  AOI22_X1 U20484 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17276), .ZN(n17268) );
  OAI211_X1 U20485 ( .C1(n17270), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17337), .B(
        n17266), .ZN(n17267) );
  OAI211_X1 U20486 ( .C1(n17269), .C2(n17348), .A(n17268), .B(n17267), .ZN(
        P3_U2717) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17276), .ZN(n17274) );
  INV_X1 U20488 ( .A(n17270), .ZN(n17271) );
  OAI211_X1 U20489 ( .C1(n17272), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17337), .B(
        n17271), .ZN(n17273) );
  OAI211_X1 U20490 ( .C1(n17275), .C2(n17348), .A(n17274), .B(n17273), .ZN(
        P3_U2718) );
  AOI22_X1 U20491 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17277), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17276), .ZN(n17280) );
  OAI211_X1 U20492 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17282), .A(n17337), .B(
        n17278), .ZN(n17279) );
  OAI211_X1 U20493 ( .C1(n17281), .C2(n17348), .A(n17280), .B(n17279), .ZN(
        P3_U2719) );
  AOI211_X1 U20494 ( .C1(n17464), .C2(n17288), .A(n17283), .B(n17282), .ZN(
        n17284) );
  AOI21_X1 U20495 ( .B1(n17343), .B2(BUF2_REG_15__SCAN_IN), .A(n17284), .ZN(
        n17285) );
  OAI21_X1 U20496 ( .B1(n17286), .B2(n17348), .A(n17285), .ZN(P3_U2720) );
  INV_X1 U20497 ( .A(n17335), .ZN(n17345) );
  AND3_X1 U20498 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17287), .A3(n17321), .ZN(
        n17295) );
  INV_X1 U20499 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17460) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17343), .B1(n17295), .B2(
        n17460), .ZN(n17290) );
  NAND3_X1 U20501 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17337), .A3(n17288), 
        .ZN(n17289) );
  OAI211_X1 U20502 ( .C1(n17291), .C2(n17348), .A(n17290), .B(n17289), .ZN(
        P3_U2721) );
  NAND2_X1 U20503 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17321), .ZN(n17307) );
  NOR2_X1 U20504 ( .A1(n17393), .A2(n17307), .ZN(n17311) );
  NAND2_X1 U20505 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17311), .ZN(n17303) );
  NOR2_X1 U20506 ( .A1(n17292), .A2(n17303), .ZN(n17298) );
  AOI21_X1 U20507 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17337), .A(n17298), .ZN(
        n17294) );
  OAI222_X1 U20508 ( .A1(n17341), .A2(n17458), .B1(n17295), .B2(n17294), .C1(
        n17348), .C2(n17293), .ZN(P3_U2722) );
  INV_X1 U20509 ( .A(n17303), .ZN(n17299) );
  AOI22_X1 U20510 ( .A1(n17299), .A2(P3_EAX_REG_11__SCAN_IN), .B1(
        P3_EAX_REG_12__SCAN_IN), .B2(n17337), .ZN(n17297) );
  OAI222_X1 U20511 ( .A1(n17341), .A2(n17454), .B1(n17298), .B2(n17297), .C1(
        n17348), .C2(n17296), .ZN(P3_U2723) );
  INV_X1 U20512 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17389) );
  NOR2_X1 U20513 ( .A1(n17389), .A2(n17303), .ZN(n17302) );
  AOI21_X1 U20514 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17337), .A(n17299), .ZN(
        n17301) );
  OAI222_X1 U20515 ( .A1(n17341), .A2(n17452), .B1(n17302), .B2(n17301), .C1(
        n17348), .C2(n17300), .ZN(P3_U2724) );
  OAI211_X1 U20516 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17311), .A(n17337), .B(
        n17303), .ZN(n17306) );
  NAND2_X1 U20517 ( .A1(n17316), .A2(n17304), .ZN(n17305) );
  OAI211_X1 U20518 ( .C1(n17341), .C2(n17449), .A(n17306), .B(n17305), .ZN(
        P3_U2725) );
  INV_X1 U20519 ( .A(n17307), .ZN(n17308) );
  AOI21_X1 U20520 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17337), .A(n17308), .ZN(
        n17310) );
  OAI222_X1 U20521 ( .A1(n17341), .A2(n17447), .B1(n17311), .B2(n17310), .C1(
        n17348), .C2(n17309), .ZN(P3_U2726) );
  OAI21_X1 U20522 ( .B1(n17313), .B2(n18188), .A(n17312), .ZN(n17314) );
  OAI21_X1 U20523 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(n17321), .A(n17314), .ZN(
        n17318) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17343), .B1(n17316), .B2(
        n17315), .ZN(n17317) );
  NAND2_X1 U20525 ( .A1(n17318), .A2(n17317), .ZN(P3_U2727) );
  INV_X1 U20526 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17399) );
  INV_X1 U20527 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17407) );
  NOR3_X1 U20528 ( .A1(n17344), .A2(n17407), .A3(n17335), .ZN(n17340) );
  NAND2_X1 U20529 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17340), .ZN(n17328) );
  NOR2_X1 U20530 ( .A1(n17403), .A2(n17328), .ZN(n17331) );
  NAND2_X1 U20531 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17331), .ZN(n17322) );
  NOR2_X1 U20532 ( .A1(n17399), .A2(n17322), .ZN(n17324) );
  AOI21_X1 U20533 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17337), .A(n17324), .ZN(
        n17320) );
  OAI222_X1 U20534 ( .A1(n17341), .A2(n18191), .B1(n17321), .B2(n17320), .C1(
        n17348), .C2(n17319), .ZN(P3_U2728) );
  INV_X1 U20535 ( .A(n17322), .ZN(n17327) );
  AOI21_X1 U20536 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17337), .A(n17327), .ZN(
        n17323) );
  OAI222_X1 U20537 ( .A1(n18185), .A2(n17341), .B1(n17324), .B2(n17323), .C1(
        n17348), .C2(n17761), .ZN(P3_U2729) );
  AOI21_X1 U20538 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17337), .A(n17331), .ZN(
        n17326) );
  OAI222_X1 U20539 ( .A1(n18181), .A2(n17341), .B1(n17327), .B2(n17326), .C1(
        n17348), .C2(n17325), .ZN(P3_U2730) );
  INV_X1 U20540 ( .A(n17328), .ZN(n17334) );
  AOI21_X1 U20541 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17337), .A(n17334), .ZN(
        n17330) );
  OAI222_X1 U20542 ( .A1(n18177), .A2(n17341), .B1(n17331), .B2(n17330), .C1(
        n17348), .C2(n17329), .ZN(P3_U2731) );
  AOI21_X1 U20543 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17337), .A(n17340), .ZN(
        n17333) );
  OAI222_X1 U20544 ( .A1(n18173), .A2(n17341), .B1(n17334), .B2(n17333), .C1(
        n17348), .C2(n17332), .ZN(P3_U2732) );
  NOR2_X1 U20545 ( .A1(n17344), .A2(n17335), .ZN(n17336) );
  AOI21_X1 U20546 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17337), .A(n17336), .ZN(
        n17339) );
  OAI222_X1 U20547 ( .A1(n18168), .A2(n17341), .B1(n17340), .B2(n17339), .C1(
        n17348), .C2(n17338), .ZN(P3_U2733) );
  AOI22_X1 U20548 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17343), .B1(n17342), .B2(
        P3_EAX_REG_1__SCAN_IN), .ZN(n17347) );
  OAI211_X1 U20549 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17345), .B(n17344), .ZN(n17346) );
  OAI211_X1 U20550 ( .C1(n17349), .C2(n17348), .A(n17347), .B(n17346), .ZN(
        P3_U2734) );
  INV_X1 U20551 ( .A(n17507), .ZN(n18659) );
  NOR2_X1 U20552 ( .A1(n18813), .A2(n18659), .ZN(n18805) );
  AND2_X1 U20553 ( .A1(n17377), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20554 ( .A1(n17381), .A2(n18157), .ZN(n17379) );
  AOI22_X1 U20555 ( .A1(n18805), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17409), .ZN(n17351) );
  OAI21_X1 U20556 ( .B1(n17433), .B2(n17379), .A(n17351), .ZN(P3_U2737) );
  AOI22_X1 U20557 ( .A1(n18805), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17352) );
  OAI21_X1 U20558 ( .B1(n17353), .B2(n17379), .A(n17352), .ZN(P3_U2738) );
  INV_X1 U20559 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17355) );
  AOI22_X1 U20560 ( .A1(n18805), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17354) );
  OAI21_X1 U20561 ( .B1(n17355), .B2(n17379), .A(n17354), .ZN(P3_U2739) );
  AOI22_X1 U20562 ( .A1(n18805), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17356) );
  OAI21_X1 U20563 ( .B1(n17357), .B2(n17379), .A(n17356), .ZN(P3_U2740) );
  INV_X1 U20564 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U20565 ( .A1(n18805), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17358) );
  OAI21_X1 U20566 ( .B1(n17359), .B2(n17379), .A(n17358), .ZN(P3_U2741) );
  AOI22_X1 U20567 ( .A1(n18805), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17360) );
  OAI21_X1 U20568 ( .B1(n17361), .B2(n17379), .A(n17360), .ZN(P3_U2742) );
  INV_X1 U20569 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U20570 ( .A1(n18805), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17362) );
  OAI21_X1 U20571 ( .B1(n17363), .B2(n17379), .A(n17362), .ZN(P3_U2743) );
  INV_X1 U20572 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U20573 ( .A1(n18805), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20574 ( .B1(n17365), .B2(n17379), .A(n17364), .ZN(P3_U2744) );
  CLKBUF_X1 U20575 ( .A(n18805), .Z(n18641) );
  AOI22_X1 U20576 ( .A1(n18641), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17366) );
  OAI21_X1 U20577 ( .B1(n17367), .B2(n17379), .A(n17366), .ZN(P3_U2745) );
  AOI22_X1 U20578 ( .A1(n18641), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17368) );
  OAI21_X1 U20579 ( .B1(n17369), .B2(n17379), .A(n17368), .ZN(P3_U2746) );
  AOI22_X1 U20580 ( .A1(n18641), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17370) );
  OAI21_X1 U20581 ( .B1(n17371), .B2(n17379), .A(n17370), .ZN(P3_U2747) );
  AOI22_X1 U20582 ( .A1(n18641), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17372) );
  OAI21_X1 U20583 ( .B1(n17373), .B2(n17379), .A(n17372), .ZN(P3_U2748) );
  INV_X1 U20584 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U20585 ( .A1(n18641), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17374) );
  OAI21_X1 U20586 ( .B1(n17375), .B2(n17379), .A(n17374), .ZN(P3_U2749) );
  AOI22_X1 U20587 ( .A1(n18641), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17376) );
  OAI21_X1 U20588 ( .B1(n17419), .B2(n17379), .A(n17376), .ZN(P3_U2750) );
  INV_X1 U20589 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17380) );
  AOI22_X1 U20590 ( .A1(n18641), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17377), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17378) );
  OAI21_X1 U20591 ( .B1(n17380), .B2(n17379), .A(n17378), .ZN(P3_U2751) );
  AOI22_X1 U20592 ( .A1(n18641), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U20593 ( .B1(n17464), .B2(n17411), .A(n17382), .ZN(P3_U2752) );
  AOI22_X1 U20594 ( .A1(n18641), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20595 ( .B1(n17460), .B2(n17411), .A(n17383), .ZN(P3_U2753) );
  AOI22_X1 U20596 ( .A1(n18641), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20597 ( .B1(n17385), .B2(n17411), .A(n17384), .ZN(P3_U2754) );
  INV_X1 U20598 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20599 ( .A1(n18641), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17386) );
  OAI21_X1 U20600 ( .B1(n17387), .B2(n17411), .A(n17386), .ZN(P3_U2755) );
  AOI22_X1 U20601 ( .A1(n18641), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20602 ( .B1(n17389), .B2(n17411), .A(n17388), .ZN(P3_U2756) );
  AOI22_X1 U20603 ( .A1(n18641), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20604 ( .B1(n17391), .B2(n17411), .A(n17390), .ZN(P3_U2757) );
  AOI22_X1 U20605 ( .A1(n18641), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20606 ( .B1(n17393), .B2(n17411), .A(n17392), .ZN(P3_U2758) );
  AOI22_X1 U20607 ( .A1(n18641), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17394) );
  OAI21_X1 U20608 ( .B1(n17395), .B2(n17411), .A(n17394), .ZN(P3_U2759) );
  INV_X1 U20609 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20610 ( .A1(n18641), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20611 ( .B1(n17397), .B2(n17411), .A(n17396), .ZN(P3_U2760) );
  AOI22_X1 U20612 ( .A1(n18641), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20613 ( .B1(n17399), .B2(n17411), .A(n17398), .ZN(P3_U2761) );
  AOI22_X1 U20614 ( .A1(n18641), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20615 ( .B1(n17401), .B2(n17411), .A(n17400), .ZN(P3_U2762) );
  AOI22_X1 U20616 ( .A1(n18641), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20617 ( .B1(n17403), .B2(n17411), .A(n17402), .ZN(P3_U2763) );
  INV_X1 U20618 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20619 ( .A1(n18641), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20620 ( .B1(n17405), .B2(n17411), .A(n17404), .ZN(P3_U2764) );
  AOI22_X1 U20621 ( .A1(n18641), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17406) );
  OAI21_X1 U20622 ( .B1(n17407), .B2(n17411), .A(n17406), .ZN(P3_U2765) );
  INV_X1 U20623 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20624 ( .A1(n18641), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20625 ( .B1(n17436), .B2(n17411), .A(n17408), .ZN(P3_U2766) );
  AOI22_X1 U20626 ( .A1(n18641), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17409), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20627 ( .B1(n17412), .B2(n17411), .A(n17410), .ZN(P3_U2767) );
  AOI21_X1 U20628 ( .B1(n18669), .B2(n18164), .A(n17414), .ZN(n17415) );
  NAND2_X1 U20629 ( .A1(n17413), .A2(n17415), .ZN(n17457) );
  NAND2_X1 U20630 ( .A1(n18808), .A2(n17416), .ZN(n18643) );
  AOI22_X1 U20631 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17443), .ZN(n17417) );
  OAI21_X1 U20632 ( .B1(n18158), .B2(n17457), .A(n17417), .ZN(P3_U2768) );
  INV_X1 U20633 ( .A(n17457), .ZN(n17461) );
  AOI22_X1 U20634 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17461), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17443), .ZN(n17418) );
  OAI21_X1 U20635 ( .B1(n17419), .B2(n17463), .A(n17418), .ZN(P3_U2769) );
  AOI22_X1 U20636 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17443), .ZN(n17420) );
  OAI21_X1 U20637 ( .B1(n18168), .B2(n17457), .A(n17420), .ZN(P3_U2770) );
  AOI22_X1 U20638 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17443), .ZN(n17421) );
  OAI21_X1 U20639 ( .B1(n18173), .B2(n17457), .A(n17421), .ZN(P3_U2771) );
  AOI22_X1 U20640 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17443), .ZN(n17422) );
  OAI21_X1 U20641 ( .B1(n18177), .B2(n17457), .A(n17422), .ZN(P3_U2772) );
  AOI22_X1 U20642 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17443), .ZN(n17423) );
  OAI21_X1 U20643 ( .B1(n18181), .B2(n17457), .A(n17423), .ZN(P3_U2773) );
  AOI22_X1 U20644 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17443), .ZN(n17424) );
  OAI21_X1 U20645 ( .B1(n18185), .B2(n17457), .A(n17424), .ZN(P3_U2774) );
  AOI22_X1 U20646 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17443), .ZN(n17425) );
  OAI21_X1 U20647 ( .B1(n18191), .B2(n17457), .A(n17425), .ZN(P3_U2775) );
  AOI22_X1 U20648 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17443), .ZN(n17426) );
  OAI21_X1 U20649 ( .B1(n17445), .B2(n17457), .A(n17426), .ZN(P3_U2776) );
  AOI22_X1 U20650 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17443), .ZN(n17427) );
  OAI21_X1 U20651 ( .B1(n17447), .B2(n17457), .A(n17427), .ZN(P3_U2777) );
  AOI22_X1 U20652 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17443), .ZN(n17428) );
  OAI21_X1 U20653 ( .B1(n17449), .B2(n17457), .A(n17428), .ZN(P3_U2778) );
  AOI22_X1 U20654 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17443), .ZN(n17429) );
  OAI21_X1 U20655 ( .B1(n17452), .B2(n17457), .A(n17429), .ZN(P3_U2779) );
  AOI22_X1 U20656 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17443), .ZN(n17430) );
  OAI21_X1 U20657 ( .B1(n17454), .B2(n17457), .A(n17430), .ZN(P3_U2780) );
  INV_X2 U20658 ( .A(n17463), .ZN(n17455) );
  AOI22_X1 U20659 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17455), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17443), .ZN(n17431) );
  OAI21_X1 U20660 ( .B1(n17458), .B2(n17451), .A(n17431), .ZN(P3_U2781) );
  AOI22_X1 U20661 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17461), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17443), .ZN(n17432) );
  OAI21_X1 U20662 ( .B1(n17433), .B2(n17463), .A(n17432), .ZN(P3_U2782) );
  AOI22_X1 U20663 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17443), .ZN(n17434) );
  OAI21_X1 U20664 ( .B1(n18158), .B2(n17451), .A(n17434), .ZN(P3_U2783) );
  AOI22_X1 U20665 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17461), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17443), .ZN(n17435) );
  OAI21_X1 U20666 ( .B1(n17436), .B2(n17463), .A(n17435), .ZN(P3_U2784) );
  AOI22_X1 U20667 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17443), .ZN(n17437) );
  OAI21_X1 U20668 ( .B1(n18168), .B2(n17451), .A(n17437), .ZN(P3_U2785) );
  AOI22_X1 U20669 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17443), .ZN(n17438) );
  OAI21_X1 U20670 ( .B1(n18173), .B2(n17451), .A(n17438), .ZN(P3_U2786) );
  AOI22_X1 U20671 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17443), .ZN(n17439) );
  OAI21_X1 U20672 ( .B1(n18177), .B2(n17451), .A(n17439), .ZN(P3_U2787) );
  AOI22_X1 U20673 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17443), .ZN(n17440) );
  OAI21_X1 U20674 ( .B1(n18181), .B2(n17451), .A(n17440), .ZN(P3_U2788) );
  AOI22_X1 U20675 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17443), .ZN(n17441) );
  OAI21_X1 U20676 ( .B1(n18185), .B2(n17451), .A(n17441), .ZN(P3_U2789) );
  AOI22_X1 U20677 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17443), .ZN(n17442) );
  OAI21_X1 U20678 ( .B1(n18191), .B2(n17451), .A(n17442), .ZN(P3_U2790) );
  AOI22_X1 U20679 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17443), .ZN(n17444) );
  OAI21_X1 U20680 ( .B1(n17445), .B2(n17451), .A(n17444), .ZN(P3_U2791) );
  AOI22_X1 U20681 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17443), .ZN(n17446) );
  OAI21_X1 U20682 ( .B1(n17447), .B2(n17451), .A(n17446), .ZN(P3_U2792) );
  AOI22_X1 U20683 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17443), .ZN(n17448) );
  OAI21_X1 U20684 ( .B1(n17449), .B2(n17451), .A(n17448), .ZN(P3_U2793) );
  AOI22_X1 U20685 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17443), .ZN(n17450) );
  OAI21_X1 U20686 ( .B1(n17452), .B2(n17451), .A(n17450), .ZN(P3_U2794) );
  AOI22_X1 U20687 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17443), .ZN(n17453) );
  OAI21_X1 U20688 ( .B1(n17454), .B2(n17457), .A(n17453), .ZN(P3_U2795) );
  AOI22_X1 U20689 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17455), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17443), .ZN(n17456) );
  OAI21_X1 U20690 ( .B1(n17458), .B2(n17457), .A(n17456), .ZN(P3_U2796) );
  AOI22_X1 U20691 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17461), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17443), .ZN(n17459) );
  OAI21_X1 U20692 ( .B1(n17460), .B2(n17463), .A(n17459), .ZN(P3_U2797) );
  AOI22_X1 U20693 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17461), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17443), .ZN(n17462) );
  OAI21_X1 U20694 ( .B1(n17464), .B2(n17463), .A(n17462), .ZN(P3_U2798) );
  INV_X1 U20695 ( .A(n17476), .ZN(n17465) );
  OAI21_X1 U20696 ( .B1(n17465), .B2(n17791), .A(n17830), .ZN(n17466) );
  AOI21_X1 U20697 ( .B1(n17507), .B2(n17467), .A(n17466), .ZN(n17500) );
  OAI21_X1 U20698 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17608), .A(
        n17500), .ZN(n17485) );
  AOI22_X1 U20699 ( .A1(n17685), .A2(n17468), .B1(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n17485), .ZN(n17481) );
  AOI21_X1 U20700 ( .B1(n17471), .B2(n17470), .A(n17469), .ZN(n17475) );
  NOR3_X1 U20701 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17836), .A3(
        n17492), .ZN(n17474) );
  NOR2_X1 U20702 ( .A1(n17528), .A2(n17818), .ZN(n17582) );
  OAI22_X1 U20703 ( .A1(n17843), .A2(n17737), .B1(n17842), .B2(n17834), .ZN(
        n17502) );
  NOR2_X1 U20704 ( .A1(n17836), .A2(n17502), .ZN(n17493) );
  NOR3_X1 U20705 ( .A1(n17582), .A2(n17493), .A3(n17472), .ZN(n17473) );
  AOI211_X1 U20706 ( .C1(n17739), .C2(n17475), .A(n17474), .B(n17473), .ZN(
        n17480) );
  NAND2_X1 U20707 ( .A1(n9821), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17479) );
  INV_X1 U20708 ( .A(n17663), .ZN(n17590) );
  NOR2_X1 U20709 ( .A1(n17590), .A2(n17476), .ZN(n17490) );
  OAI211_X1 U20710 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17490), .B(n17477), .ZN(n17478) );
  NAND4_X1 U20711 ( .A1(n17481), .A2(n17480), .A3(n17479), .A4(n17478), .ZN(
        P3_U2802) );
  NAND2_X1 U20712 ( .A1(n17483), .A2(n17482), .ZN(n17484) );
  XNOR2_X1 U20713 ( .A(n17484), .B(n17734), .ZN(n17850) );
  AOI22_X1 U20714 ( .A1(n17685), .A2(n17486), .B1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n17485), .ZN(n17487) );
  NAND2_X1 U20715 ( .A1(n9821), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17848) );
  OAI211_X1 U20716 ( .C1(n17850), .C2(n17717), .A(n17487), .B(n17848), .ZN(
        n17488) );
  AOI21_X1 U20717 ( .B1(n17490), .B2(n17489), .A(n17488), .ZN(n17491) );
  OAI221_X1 U20718 ( .B1(n17493), .B2(n17836), .C1(n17493), .C2(n17492), .A(
        n17491), .ZN(P3_U2803) );
  AOI21_X1 U20719 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17495), .A(
        n17494), .ZN(n17857) );
  AOI21_X1 U20720 ( .B1(n17496), .B2(n18529), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17499) );
  OAI21_X1 U20721 ( .B1(n17685), .B2(n17539), .A(n17497), .ZN(n17498) );
  NAND2_X1 U20722 ( .A1(n9821), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17855) );
  OAI211_X1 U20723 ( .C1(n17500), .C2(n17499), .A(n17498), .B(n17855), .ZN(
        n17501) );
  AOI221_X1 U20724 ( .B1(n17503), .B2(n17851), .C1(n17502), .C2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n17501), .ZN(n17504) );
  OAI21_X1 U20725 ( .B1(n17857), .B2(n17717), .A(n17504), .ZN(P3_U2804) );
  XNOR2_X1 U20726 ( .A(n17515), .B(n17505), .ZN(n17865) );
  AND2_X1 U20727 ( .A1(n17508), .A2(n18529), .ZN(n17548) );
  AOI211_X1 U20728 ( .C1(n17507), .C2(n17506), .A(n17801), .B(n17548), .ZN(
        n17542) );
  OAI21_X1 U20729 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17608), .A(
        n17542), .ZN(n17521) );
  NOR2_X1 U20730 ( .A1(n17590), .A2(n17508), .ZN(n17523) );
  OAI211_X1 U20731 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17523), .B(n17509), .ZN(n17510) );
  NAND2_X1 U20732 ( .A1(n9821), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17862) );
  OAI211_X1 U20733 ( .C1(n17669), .C2(n17511), .A(n17510), .B(n17862), .ZN(
        n17518) );
  XNOR2_X1 U20734 ( .A(n17512), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17869) );
  OAI21_X1 U20735 ( .B1(n17702), .B2(n17514), .A(n17513), .ZN(n17516) );
  XNOR2_X1 U20736 ( .A(n17516), .B(n17515), .ZN(n17864) );
  OAI22_X1 U20737 ( .A1(n17737), .A2(n17869), .B1(n17717), .B2(n17864), .ZN(
        n17517) );
  AOI211_X1 U20738 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17521), .A(
        n17518), .B(n17517), .ZN(n17519) );
  OAI21_X1 U20739 ( .B1(n17834), .B2(n17865), .A(n17519), .ZN(P3_U2805) );
  INV_X1 U20740 ( .A(n17520), .ZN(n17534) );
  NOR2_X1 U20741 ( .A1(n18036), .A2(n18725), .ZN(n17872) );
  AOI221_X1 U20742 ( .B1(n17523), .B2(n17522), .C1(n17521), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17872), .ZN(n17533) );
  OAI21_X1 U20743 ( .B1(n17525), .B2(n17524), .A(n11313), .ZN(n17873) );
  NOR2_X1 U20744 ( .A1(n17526), .A2(n17633), .ZN(n17530) );
  INV_X1 U20745 ( .A(n17527), .ZN(n17875) );
  AOI22_X1 U20746 ( .A1(n17528), .A2(n17874), .B1(n17818), .B2(n17875), .ZN(
        n17529) );
  INV_X1 U20747 ( .A(n17529), .ZN(n17544) );
  MUX2_X1 U20748 ( .A(n17530), .B(n17544), .S(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n17531) );
  AOI21_X1 U20749 ( .B1(n17739), .B2(n17873), .A(n17531), .ZN(n17532) );
  OAI211_X1 U20750 ( .C1(n17669), .C2(n17534), .A(n17533), .B(n17532), .ZN(
        P3_U2806) );
  AOI22_X1 U20751 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17702), .B1(
        n17535), .B2(n17555), .ZN(n17536) );
  NAND2_X1 U20752 ( .A1(n17576), .A2(n17536), .ZN(n17537) );
  XNOR2_X1 U20753 ( .A(n17537), .B(n17878), .ZN(n17890) );
  NAND2_X1 U20754 ( .A1(n9821), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17889) );
  INV_X1 U20755 ( .A(n17608), .ZN(n17539) );
  OAI21_X1 U20756 ( .B1(n17685), .B2(n17539), .A(n17538), .ZN(n17540) );
  OAI211_X1 U20757 ( .C1(n17542), .C2(n17541), .A(n17889), .B(n17540), .ZN(
        n17547) );
  NOR2_X1 U20758 ( .A1(n17543), .A2(n17557), .ZN(n17545) );
  MUX2_X1 U20759 ( .A(n17545), .B(n17544), .S(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(n17546) );
  AOI211_X1 U20760 ( .C1(n17549), .C2(n17548), .A(n17547), .B(n17546), .ZN(
        n17550) );
  OAI21_X1 U20761 ( .B1(n17717), .B2(n17890), .A(n17550), .ZN(P3_U2807) );
  OAI21_X1 U20762 ( .B1(n17551), .B2(n18659), .A(n17830), .ZN(n17552) );
  AOI21_X1 U20763 ( .B1(n17625), .B2(n17559), .A(n17552), .ZN(n17579) );
  OAI21_X1 U20764 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17608), .A(
        n17579), .ZN(n17570) );
  AOI22_X1 U20765 ( .A1(n17685), .A2(n17553), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17570), .ZN(n17563) );
  NOR2_X1 U20766 ( .A1(n17891), .A2(n17737), .ZN(n17644) );
  AOI21_X1 U20767 ( .B1(n17818), .B2(n17970), .A(n17644), .ZN(n17632) );
  OAI21_X1 U20768 ( .B1(n17895), .B2(n17582), .A(n17632), .ZN(n17573) );
  INV_X1 U20769 ( .A(n17576), .ZN(n17554) );
  AOI221_X1 U20770 ( .B1(n17900), .B2(n17555), .C1(n17564), .C2(n17555), .A(
        n17554), .ZN(n17556) );
  XNOR2_X1 U20771 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n17556), .ZN(
        n17905) );
  OAI22_X1 U20772 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17557), .B1(
        n17905), .B2(n17717), .ZN(n17558) );
  AOI21_X1 U20773 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17573), .A(
        n17558), .ZN(n17562) );
  NAND2_X1 U20774 ( .A1(n9821), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17907) );
  NOR2_X1 U20775 ( .A1(n17590), .A2(n17559), .ZN(n17572) );
  OAI211_X1 U20776 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17572), .B(n17560), .ZN(n17561) );
  NAND4_X1 U20777 ( .A1(n17563), .A2(n17562), .A3(n17907), .A4(n17561), .ZN(
        P3_U2808) );
  INV_X1 U20778 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17894) );
  NOR3_X1 U20779 ( .A1(n17702), .A2(n17894), .A3(n17564), .ZN(n17585) );
  INV_X1 U20780 ( .A(n17565), .ZN(n17586) );
  AOI22_X1 U20781 ( .A1(n17916), .A2(n17585), .B1(n17586), .B2(n17566), .ZN(
        n17567) );
  XNOR2_X1 U20782 ( .A(n17567), .B(n17897), .ZN(n17920) );
  OAI22_X1 U20783 ( .A1(n18036), .A2(n18720), .B1(n17669), .B2(n17568), .ZN(
        n17569) );
  AOI221_X1 U20784 ( .B1(n17572), .B2(n17571), .C1(n17570), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17569), .ZN(n17575) );
  NOR2_X1 U20785 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17898), .ZN(
        n17911) );
  NAND2_X1 U20786 ( .A1(n17940), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17912) );
  NOR2_X1 U20787 ( .A1(n17633), .A2(n17912), .ZN(n17597) );
  AOI22_X1 U20788 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17573), .B1(
        n17911), .B2(n17597), .ZN(n17574) );
  OAI211_X1 U20789 ( .C1(n17920), .C2(n17717), .A(n17575), .B(n17574), .ZN(
        P3_U2809) );
  OAI221_X1 U20790 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17604), 
        .C1(n17929), .C2(n17585), .A(n17576), .ZN(n17577) );
  XOR2_X1 U20791 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17577), .Z(
        n17928) );
  AOI21_X1 U20792 ( .B1(n9928), .B2(n18529), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17578) );
  INV_X1 U20793 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18717) );
  OAI22_X1 U20794 ( .A1(n17579), .A2(n17578), .B1(n18036), .B2(n18717), .ZN(
        n17580) );
  AOI221_X1 U20795 ( .B1(n17685), .B2(n17581), .C1(n17539), .C2(n17581), .A(
        n17580), .ZN(n17584) );
  NOR2_X1 U20796 ( .A1(n17929), .A2(n17912), .ZN(n17924) );
  OAI21_X1 U20797 ( .B1(n17582), .B2(n17924), .A(n17632), .ZN(n17596) );
  NOR2_X1 U20798 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17929), .ZN(
        n17921) );
  AOI22_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17596), .B1(
        n17597), .B2(n17921), .ZN(n17583) );
  OAI211_X1 U20800 ( .C1(n17717), .C2(n17928), .A(n17584), .B(n17583), .ZN(
        P3_U2810) );
  AOI21_X1 U20801 ( .B1(n17586), .B2(n17604), .A(n17585), .ZN(n17587) );
  XNOR2_X1 U20802 ( .A(n17587), .B(n17929), .ZN(n17934) );
  AOI21_X1 U20803 ( .B1(n17625), .B2(n17589), .A(n17801), .ZN(n17612) );
  OAI21_X1 U20804 ( .B1(n17588), .B2(n18659), .A(n17612), .ZN(n17601) );
  AOI22_X1 U20805 ( .A1(n9821), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17601), .ZN(n17593) );
  NOR2_X1 U20806 ( .A1(n17590), .A2(n17589), .ZN(n17603) );
  OAI211_X1 U20807 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17603), .B(n17591), .ZN(n17592) );
  OAI211_X1 U20808 ( .C1(n17669), .C2(n17594), .A(n17593), .B(n17592), .ZN(
        n17595) );
  AOI221_X1 U20809 ( .B1(n17597), .B2(n17929), .C1(n17596), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17595), .ZN(n17598) );
  OAI21_X1 U20810 ( .B1(n17934), .B2(n17717), .A(n17598), .ZN(P3_U2811) );
  NAND2_X1 U20811 ( .A1(n17940), .A2(n17894), .ZN(n17949) );
  OAI22_X1 U20812 ( .A1(n18036), .A2(n18713), .B1(n17669), .B2(n17599), .ZN(
        n17600) );
  AOI221_X1 U20813 ( .B1(n17603), .B2(n17602), .C1(n17601), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17600), .ZN(n17607) );
  OAI21_X1 U20814 ( .B1(n17940), .B2(n17633), .A(n17632), .ZN(n17615) );
  AOI21_X1 U20815 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17734), .A(
        n17604), .ZN(n17605) );
  XNOR2_X1 U20816 ( .A(n17605), .B(n17565), .ZN(n17945) );
  AOI22_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17615), .B1(
        n17739), .B2(n17945), .ZN(n17606) );
  OAI211_X1 U20818 ( .C1(n17633), .C2(n17949), .A(n17607), .B(n17606), .ZN(
        P3_U2812) );
  OAI21_X1 U20819 ( .B1(n17610), .B2(n17950), .A(n17609), .ZN(n17954) );
  AOI21_X1 U20820 ( .B1(n17611), .B2(n18529), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17613) );
  OAI22_X1 U20821 ( .A1(n17613), .A2(n17612), .B1(n18036), .B2(n18712), .ZN(
        n17614) );
  AOI21_X1 U20822 ( .B1(n17739), .B2(n17954), .A(n17614), .ZN(n17618) );
  OAI221_X1 U20823 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17616), .A(n17615), .ZN(
        n17617) );
  OAI211_X1 U20824 ( .C1(n17813), .C2(n17619), .A(n17618), .B(n17617), .ZN(
        P3_U2813) );
  AOI21_X1 U20825 ( .B1(n17734), .B2(n17621), .A(n17620), .ZN(n17622) );
  XNOR2_X1 U20826 ( .A(n17622), .B(n17960), .ZN(n17964) );
  NAND4_X1 U20827 ( .A1(n17664), .A2(n17666), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A4(n17663), .ZN(n17635) );
  OAI21_X1 U20828 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17623), .ZN(n17629) );
  AOI21_X1 U20829 ( .B1(n17625), .B2(n17624), .A(n17801), .ZN(n17650) );
  OAI21_X1 U20830 ( .B1(n17626), .B2(n18659), .A(n17650), .ZN(n17637) );
  AOI22_X1 U20831 ( .A1(n17685), .A2(n17627), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17637), .ZN(n17628) );
  NAND2_X1 U20832 ( .A1(n9821), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17965) );
  OAI211_X1 U20833 ( .C1(n17635), .C2(n17629), .A(n17628), .B(n17965), .ZN(
        n17630) );
  AOI21_X1 U20834 ( .B1(n17739), .B2(n17964), .A(n17630), .ZN(n17631) );
  OAI221_X1 U20835 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17633), 
        .C1(n17960), .C2(n17632), .A(n17631), .ZN(P3_U2814) );
  OAI22_X1 U20836 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17635), .B1(
        n17669), .B2(n17634), .ZN(n17636) );
  AOI21_X1 U20837 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17637), .A(
        n17636), .ZN(n17647) );
  INV_X1 U20838 ( .A(n17638), .ZN(n17640) );
  OR2_X1 U20839 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17639), .ZN(
        n17723) );
  NOR2_X1 U20840 ( .A1(n17640), .A2(n17723), .ZN(n17655) );
  NOR4_X1 U20841 ( .A1(n17702), .A2(n17642), .A3(n18071), .A4(n17641), .ZN(
        n17678) );
  INV_X1 U20842 ( .A(n17678), .ZN(n17724) );
  NOR3_X1 U20843 ( .A1(n18010), .A2(n18009), .A3(n17724), .ZN(n17661) );
  INV_X1 U20844 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17651) );
  NAND2_X1 U20845 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17651), .ZN(
        n17654) );
  OAI221_X1 U20846 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17655), 
        .C1(n17987), .C2(n17661), .A(n17654), .ZN(n17643) );
  XNOR2_X1 U20847 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17643), .ZN(
        n17977) );
  NAND2_X1 U20848 ( .A1(n17997), .A2(n17968), .ZN(n17648) );
  NAND2_X1 U20849 ( .A1(n11303), .A2(n17648), .ZN(n17972) );
  AOI22_X1 U20850 ( .A1(n17739), .A2(n17977), .B1(n17644), .B2(n17972), .ZN(
        n17646) );
  NAND2_X1 U20851 ( .A1(n9821), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17978) );
  NAND2_X1 U20852 ( .A1(n18006), .A2(n18018), .ZN(n18000) );
  INV_X1 U20853 ( .A(n18000), .ZN(n17673) );
  NAND3_X1 U20854 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n17673), .ZN(n17652) );
  NAND2_X1 U20855 ( .A1(n11303), .A2(n17652), .ZN(n17974) );
  NAND3_X1 U20856 ( .A1(n17818), .A2(n17970), .A3(n17974), .ZN(n17645) );
  NAND4_X1 U20857 ( .A1(n17647), .A2(n17646), .A3(n17978), .A4(n17645), .ZN(
        P3_U2815) );
  AND2_X1 U20858 ( .A1(n17997), .A2(n18006), .ZN(n17674) );
  OAI221_X1 U20859 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n17674), .A(n17648), .ZN(
        n17994) );
  INV_X1 U20860 ( .A(n17813), .ZN(n17821) );
  AND2_X1 U20861 ( .A1(n17666), .A2(n18529), .ZN(n17695) );
  AOI21_X1 U20862 ( .B1(n17664), .B2(n17695), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17649) );
  OAI22_X1 U20863 ( .A1(n17650), .A2(n17649), .B1(n18036), .B2(n18705), .ZN(
        n17658) );
  NOR2_X1 U20864 ( .A1(n17651), .A2(n18000), .ZN(n17653) );
  OAI21_X1 U20865 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17653), .A(
        n17652), .ZN(n17989) );
  OAI21_X1 U20866 ( .B1(n17661), .B2(n17655), .A(n17654), .ZN(n17656) );
  XNOR2_X1 U20867 ( .A(n17656), .B(n17987), .ZN(n17988) );
  OAI22_X1 U20868 ( .A1(n17834), .A2(n17989), .B1(n17717), .B2(n17988), .ZN(
        n17657) );
  AOI211_X1 U20869 ( .C1(n17659), .C2(n17821), .A(n17658), .B(n17657), .ZN(
        n17660) );
  OAI21_X1 U20870 ( .B1(n17737), .B2(n17994), .A(n17660), .ZN(P3_U2816) );
  NOR3_X1 U20871 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17713), .A3(
        n17723), .ZN(n17677) );
  AOI21_X1 U20872 ( .B1(n17677), .B2(n18009), .A(n17661), .ZN(n17662) );
  XOR2_X1 U20873 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n17662), .Z(
        n18005) );
  NAND2_X1 U20874 ( .A1(n17666), .A2(n17663), .ZN(n17682) );
  AOI211_X1 U20875 ( .C1(n17681), .C2(n17670), .A(n17664), .B(n17682), .ZN(
        n17672) );
  OAI22_X1 U20876 ( .A1(n17666), .A2(n17791), .B1(n17665), .B2(n18659), .ZN(
        n17667) );
  NOR2_X1 U20877 ( .A1(n17801), .A2(n17667), .ZN(n17680) );
  OAI22_X1 U20878 ( .A1(n17680), .A2(n17670), .B1(n17669), .B2(n17668), .ZN(
        n17671) );
  AOI211_X1 U20879 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n9821), .A(n17672), .B(
        n17671), .ZN(n17676) );
  OAI22_X1 U20880 ( .A1(n17674), .A2(n17737), .B1(n17673), .B2(n17834), .ZN(
        n17686) );
  NOR3_X1 U20881 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18009), .A3(
        n18010), .ZN(n17995) );
  INV_X1 U20882 ( .A(n17700), .ZN(n17726) );
  AOI22_X1 U20883 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17686), .B1(
        n17995), .B2(n17726), .ZN(n17675) );
  OAI211_X1 U20884 ( .C1(n18005), .C2(n17717), .A(n17676), .B(n17675), .ZN(
        P3_U2817) );
  INV_X1 U20885 ( .A(n18010), .ZN(n17998) );
  AOI21_X1 U20886 ( .B1(n17678), .B2(n17998), .A(n17677), .ZN(n17679) );
  XNOR2_X1 U20887 ( .A(n17679), .B(n18009), .ZN(n18015) );
  NAND2_X1 U20888 ( .A1(n9821), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18013) );
  OAI221_X1 U20889 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17682), .C1(
        n17681), .C2(n17680), .A(n18013), .ZN(n17683) );
  AOI21_X1 U20890 ( .B1(n17685), .B2(n17684), .A(n17683), .ZN(n17689) );
  OAI21_X1 U20891 ( .B1(n18010), .B2(n17700), .A(n18009), .ZN(n17687) );
  NAND2_X1 U20892 ( .A1(n17687), .A2(n17686), .ZN(n17688) );
  OAI211_X1 U20893 ( .C1(n18015), .C2(n17717), .A(n17689), .B(n17688), .ZN(
        P3_U2818) );
  INV_X1 U20894 ( .A(n18024), .ZN(n17706) );
  OR2_X1 U20895 ( .A1(n17706), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18030) );
  OAI22_X1 U20896 ( .A1(n17706), .A2(n17724), .B1(n17713), .B2(n17723), .ZN(
        n17690) );
  XOR2_X1 U20897 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17690), .Z(
        n18016) );
  INV_X1 U20898 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18699) );
  NOR2_X1 U20899 ( .A1(n18036), .A2(n18699), .ZN(n17697) );
  NOR2_X1 U20900 ( .A1(n17691), .A2(n18498), .ZN(n17747) );
  NAND2_X1 U20901 ( .A1(n17692), .A2(n17747), .ZN(n17721) );
  NOR2_X1 U20902 ( .A1(n17709), .A2(n17721), .ZN(n17708) );
  AOI21_X1 U20903 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17707), .A(
        n17708), .ZN(n17694) );
  OAI22_X1 U20904 ( .A1(n17695), .A2(n17694), .B1(n17813), .B2(n17693), .ZN(
        n17696) );
  AOI211_X1 U20905 ( .C1(n17739), .C2(n18016), .A(n17697), .B(n17696), .ZN(
        n17699) );
  NOR2_X1 U20906 ( .A1(n18024), .A2(n17700), .ZN(n17714) );
  OAI22_X1 U20907 ( .A1(n17997), .A2(n17737), .B1(n17834), .B2(n18018), .ZN(
        n17727) );
  OAI21_X1 U20908 ( .B1(n17714), .B2(n17727), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17698) );
  OAI211_X1 U20909 ( .C1(n17700), .C2(n18030), .A(n17699), .B(n17698), .ZN(
        P3_U2819) );
  OAI221_X1 U20910 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17723), .C1(
        n18041), .C2(n17724), .A(n17701), .ZN(n17705) );
  NAND4_X1 U20911 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17703), .A3(
        n17702), .A4(n18041), .ZN(n17704) );
  OAI211_X1 U20912 ( .C1(n17724), .C2(n17706), .A(n17705), .B(n17704), .ZN(
        n18040) );
  INV_X1 U20913 ( .A(n17707), .ZN(n17826) );
  AOI211_X1 U20914 ( .C1(n17721), .C2(n17709), .A(n17826), .B(n17708), .ZN(
        n17711) );
  NOR2_X1 U20915 ( .A1(n18036), .A2(n18697), .ZN(n17710) );
  AOI211_X1 U20916 ( .C1(n17712), .C2(n17821), .A(n17711), .B(n17710), .ZN(
        n17716) );
  AOI22_X1 U20917 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17727), .B1(
        n17714), .B2(n17713), .ZN(n17715) );
  OAI211_X1 U20918 ( .C1(n17717), .C2(n18040), .A(n17716), .B(n17715), .ZN(
        P3_U2820) );
  INV_X1 U20919 ( .A(n17747), .ZN(n17718) );
  OAI22_X1 U20920 ( .A1(n17826), .A2(n17719), .B1(n17718), .B2(n17740), .ZN(
        n17720) );
  AOI22_X1 U20921 ( .A1(n17821), .A2(n17722), .B1(n17721), .B2(n17720), .ZN(
        n17730) );
  NAND2_X1 U20922 ( .A1(n17724), .A2(n17723), .ZN(n17725) );
  XNOR2_X1 U20923 ( .A(n17725), .B(n18041), .ZN(n18046) );
  AOI22_X1 U20924 ( .A1(n17739), .A2(n18046), .B1(n18041), .B2(n17726), .ZN(
        n17729) );
  NAND2_X1 U20925 ( .A1(n9821), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18047) );
  NAND2_X1 U20926 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17727), .ZN(
        n17728) );
  NAND4_X1 U20927 ( .A1(n17730), .A2(n17729), .A3(n18047), .A4(n17728), .ZN(
        P3_U2821) );
  OAI21_X1 U20928 ( .B1(n17731), .B2(n17791), .A(n17830), .ZN(n17745) );
  AOI22_X1 U20929 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17745), .B1(
        n17732), .B2(n17821), .ZN(n17744) );
  AOI21_X1 U20930 ( .B1(n17734), .B2(n18065), .A(n17733), .ZN(n18061) );
  OAI21_X1 U20931 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17736), .A(
        n17735), .ZN(n18059) );
  OAI22_X1 U20932 ( .A1(n17737), .A2(n18065), .B1(n17834), .B2(n18059), .ZN(
        n17738) );
  AOI21_X1 U20933 ( .B1(n17739), .B2(n18061), .A(n17738), .ZN(n17743) );
  NAND2_X1 U20934 ( .A1(n9821), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18057) );
  OAI211_X1 U20935 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17741), .A(
        n18529), .B(n17740), .ZN(n17742) );
  NAND4_X1 U20936 ( .A1(n17744), .A2(n17743), .A3(n18057), .A4(n17742), .ZN(
        P3_U2822) );
  NOR2_X1 U20937 ( .A1(n18036), .A2(n18691), .ZN(n18073) );
  AOI221_X1 U20938 ( .B1(n17747), .B2(n17746), .C1(n17745), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18073), .ZN(n17754) );
  AOI21_X1 U20939 ( .B1(n18071), .B2(n17749), .A(n17748), .ZN(n18066) );
  NOR2_X1 U20940 ( .A1(n17751), .A2(n17750), .ZN(n17752) );
  XNOR2_X1 U20941 ( .A(n17752), .B(n18071), .ZN(n18067) );
  AOI22_X1 U20942 ( .A1(n17822), .A2(n18066), .B1(n17818), .B2(n18067), .ZN(
        n17753) );
  OAI211_X1 U20943 ( .C1(n17813), .C2(n17755), .A(n17754), .B(n17753), .ZN(
        P3_U2823) );
  NAND2_X1 U20944 ( .A1(n17768), .A2(n18529), .ZN(n17764) );
  INV_X1 U20945 ( .A(n17758), .ZN(n17756) );
  AOI22_X1 U20946 ( .A1(n17758), .A2(n17773), .B1(n17757), .B2(n17756), .ZN(
        n17763) );
  AOI22_X1 U20947 ( .A1(n17761), .A2(n17760), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17759), .ZN(n17762) );
  XNOR2_X1 U20948 ( .A(n17763), .B(n17762), .ZN(n18083) );
  OAI22_X1 U20949 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17764), .B1(
        n18083), .B2(n17834), .ZN(n17765) );
  AOI21_X1 U20950 ( .B1(n9821), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17765), .ZN(
        n17770) );
  AOI21_X1 U20951 ( .B1(n17767), .B2(n17766), .A(n9920), .ZN(n18080) );
  AOI21_X1 U20952 ( .B1(n17768), .B2(n18529), .A(n17826), .ZN(n17779) );
  AOI22_X1 U20953 ( .A1(n17822), .A2(n18080), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17779), .ZN(n17769) );
  OAI211_X1 U20954 ( .C1(n17813), .C2(n17771), .A(n17770), .B(n17769), .ZN(
        P3_U2824) );
  AOI21_X1 U20955 ( .B1(n18084), .B2(n17772), .A(n9857), .ZN(n18086) );
  AOI22_X1 U20956 ( .A1(n17822), .A2(n18086), .B1(n9821), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17781) );
  AOI21_X1 U20957 ( .B1(n17775), .B2(n17774), .A(n17773), .ZN(n18085) );
  OAI21_X1 U20958 ( .B1(n17801), .B2(n17777), .A(n17776), .ZN(n17778) );
  AOI22_X1 U20959 ( .A1(n17818), .A2(n18085), .B1(n17779), .B2(n17778), .ZN(
        n17780) );
  OAI211_X1 U20960 ( .C1(n17813), .C2(n17782), .A(n17781), .B(n17780), .ZN(
        P3_U2825) );
  AOI21_X1 U20961 ( .B1(n17785), .B2(n17784), .A(n17783), .ZN(n18094) );
  OAI22_X1 U20962 ( .A1(n18036), .A2(n18685), .B1(n18498), .B2(n17786), .ZN(
        n17787) );
  AOI21_X1 U20963 ( .B1(n17818), .B2(n18094), .A(n17787), .ZN(n17794) );
  AOI21_X1 U20964 ( .B1(n17790), .B2(n17789), .A(n17788), .ZN(n18091) );
  OAI21_X1 U20965 ( .B1(n17792), .B2(n17791), .A(n17830), .ZN(n17803) );
  AOI22_X1 U20966 ( .A1(n17822), .A2(n18091), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17803), .ZN(n17793) );
  OAI211_X1 U20967 ( .C1(n17813), .C2(n17795), .A(n17794), .B(n17793), .ZN(
        P3_U2826) );
  AOI22_X1 U20968 ( .A1(n17822), .A2(n18099), .B1(n9821), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17805) );
  AOI21_X1 U20969 ( .B1(n17799), .B2(n17798), .A(n17797), .ZN(n18100) );
  OAI21_X1 U20970 ( .B1(n17801), .B2(n17816), .A(n17800), .ZN(n17802) );
  AOI22_X1 U20971 ( .A1(n17818), .A2(n18100), .B1(n17803), .B2(n17802), .ZN(
        n17804) );
  OAI211_X1 U20972 ( .C1(n17813), .C2(n17806), .A(n17805), .B(n17804), .ZN(
        P3_U2827) );
  AOI21_X1 U20973 ( .B1(n17809), .B2(n17808), .A(n17807), .ZN(n18111) );
  NOR2_X1 U20974 ( .A1(n18036), .A2(n18681), .ZN(n18120) );
  XNOR2_X1 U20975 ( .A(n17811), .B(n17810), .ZN(n18123) );
  OAI22_X1 U20976 ( .A1(n17813), .A2(n17812), .B1(n17834), .B2(n18123), .ZN(
        n17814) );
  AOI211_X1 U20977 ( .C1(n17822), .C2(n18111), .A(n18120), .B(n17814), .ZN(
        n17815) );
  OAI221_X1 U20978 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18498), .C1(
        n17816), .C2(n17830), .A(n17815), .ZN(P3_U2828) );
  OAI21_X1 U20979 ( .B1(n17827), .B2(n17820), .A(n17817), .ZN(n18125) );
  AOI22_X1 U20980 ( .A1(n17818), .A2(n18125), .B1(n9821), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17824) );
  AOI21_X1 U20981 ( .B1(n17829), .B2(n17820), .A(n17819), .ZN(n18124) );
  AOI22_X1 U20982 ( .A1(n17822), .A2(n18124), .B1(n17825), .B2(n17821), .ZN(
        n17823) );
  OAI211_X1 U20983 ( .C1(n17826), .C2(n17825), .A(n17824), .B(n17823), .ZN(
        P3_U2829) );
  INV_X1 U20984 ( .A(n17827), .ZN(n17828) );
  NAND2_X1 U20985 ( .A1(n17829), .A2(n17828), .ZN(n18144) );
  INV_X1 U20986 ( .A(n18144), .ZN(n18146) );
  NAND3_X1 U20987 ( .A1(n18813), .A2(n17830), .A3(n18659), .ZN(n17831) );
  AOI22_X1 U20988 ( .A1(n9821), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17831), .ZN(n17832) );
  OAI221_X1 U20989 ( .B1(n18146), .B2(n17834), .C1(n18144), .C2(n17833), .A(
        n17832), .ZN(P3_U2830) );
  OR3_X1 U20990 ( .A1(n17901), .A2(n17835), .A3(n17900), .ZN(n17852) );
  AOI221_X1 U20991 ( .B1(n17851), .B2(n17836), .C1(n17852), .C2(n17836), .A(
        n18127), .ZN(n17847) );
  NAND2_X1 U20992 ( .A1(n18613), .A2(n17837), .ZN(n17879) );
  INV_X1 U20993 ( .A(n17838), .ZN(n17839) );
  AOI21_X1 U20994 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18605), .A(
        n17839), .ZN(n17904) );
  NAND2_X1 U20995 ( .A1(n18617), .A2(n18605), .ZN(n17944) );
  OAI21_X1 U20996 ( .B1(n17904), .B2(n17840), .A(n17944), .ZN(n17876) );
  OAI211_X1 U20997 ( .C1(n18053), .C2(n17860), .A(n17879), .B(n17876), .ZN(
        n17861) );
  NOR2_X1 U20998 ( .A1(n18613), .A2(n18615), .ZN(n18128) );
  OAI22_X1 U20999 ( .A1(n18617), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17841), .B2(n18128), .ZN(n17845) );
  OAI22_X1 U21000 ( .A1(n17843), .A2(n17996), .B1(n17842), .B2(n18017), .ZN(
        n17844) );
  NOR3_X1 U21001 ( .A1(n17861), .A2(n17845), .A3(n17844), .ZN(n17853) );
  OAI211_X1 U21002 ( .C1(n18617), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17853), .ZN(n17846) );
  AOI22_X1 U21003 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18129), .B1(
        n17847), .B2(n17846), .ZN(n17849) );
  OAI211_X1 U21004 ( .C1(n17850), .C2(n18039), .A(n17849), .B(n17848), .ZN(
        P3_U2835) );
  AOI221_X1 U21005 ( .B1(n17853), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), 
        .C1(n17852), .C2(n17851), .A(n18127), .ZN(n17854) );
  AOI21_X1 U21006 ( .B1(n18129), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17854), .ZN(n17856) );
  OAI211_X1 U21007 ( .C1(n17857), .C2(n18039), .A(n17856), .B(n17855), .ZN(
        P3_U2836) );
  NOR2_X1 U21008 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17858), .ZN(
        n17859) );
  AOI22_X1 U21009 ( .A1(n17861), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n17860), .B2(n17859), .ZN(n17863) );
  OAI21_X1 U21010 ( .B1(n18127), .B2(n17863), .A(n17862), .ZN(n17867) );
  OAI22_X1 U21011 ( .A1(n18145), .A2(n17865), .B1(n18039), .B2(n17864), .ZN(
        n17866) );
  AOI211_X1 U21012 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18129), .A(
        n17867), .B(n17866), .ZN(n17868) );
  OAI21_X1 U21013 ( .B1(n18064), .B2(n17869), .A(n17868), .ZN(P3_U2837) );
  NOR3_X1 U21014 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17878), .A3(
        n17870), .ZN(n17871) );
  AOI211_X1 U21015 ( .C1(n9811), .C2(n17873), .A(n17872), .B(n17871), .ZN(
        n17883) );
  INV_X1 U21016 ( .A(n18053), .ZN(n18052) );
  AOI22_X1 U21017 ( .A1(n18581), .A2(n17875), .B1(n18022), .B2(n17874), .ZN(
        n17877) );
  NAND3_X1 U21018 ( .A1(n17877), .A2(n17986), .A3(n17876), .ZN(n17881) );
  NOR2_X1 U21019 ( .A1(n17878), .A2(n17881), .ZN(n17880) );
  AOI21_X1 U21020 ( .B1(n17880), .B2(n17879), .A(n18042), .ZN(n17886) );
  OAI211_X1 U21021 ( .C1(n18052), .C2(n17881), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17886), .ZN(n17882) );
  NAND2_X1 U21022 ( .A1(n17883), .A2(n17882), .ZN(P3_U2838) );
  INV_X1 U21023 ( .A(n17884), .ZN(n17885) );
  NOR3_X1 U21024 ( .A1(n18129), .A2(n17901), .A3(n17885), .ZN(n17887) );
  OAI21_X1 U21025 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17887), .A(
        n17886), .ZN(n17888) );
  OAI211_X1 U21026 ( .C1(n17890), .C2(n18039), .A(n17889), .B(n17888), .ZN(
        P3_U2839) );
  AOI21_X1 U21027 ( .B1(n17939), .B2(n17924), .A(n18617), .ZN(n17893) );
  NOR2_X1 U21028 ( .A1(n17891), .A2(n17996), .ZN(n17971) );
  AOI21_X1 U21029 ( .B1(n18581), .B2(n17970), .A(n17971), .ZN(n17962) );
  OAI21_X1 U21030 ( .B1(n17892), .B2(n17936), .A(n17962), .ZN(n17942) );
  AOI211_X1 U21031 ( .C1(n18613), .C2(n17894), .A(n17893), .B(n17942), .ZN(
        n17914) );
  NOR2_X1 U21032 ( .A1(n18581), .A2(n18022), .ZN(n18023) );
  OAI22_X1 U21033 ( .A1(n18617), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17895), .B2(n18023), .ZN(n17896) );
  INV_X1 U21034 ( .A(n17896), .ZN(n17915) );
  AOI22_X1 U21035 ( .A1(n18613), .A2(n17898), .B1(n17982), .B2(n17897), .ZN(
        n17899) );
  NAND3_X1 U21036 ( .A1(n17914), .A2(n17915), .A3(n17899), .ZN(n17903) );
  NOR2_X1 U21037 ( .A1(n17901), .A2(n17900), .ZN(n17902) );
  OAI22_X1 U21038 ( .A1(n17904), .A2(n17903), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17902), .ZN(n17909) );
  INV_X1 U21039 ( .A(n17905), .ZN(n17906) );
  AOI22_X1 U21040 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18129), .B1(
        n9811), .B2(n17906), .ZN(n17908) );
  OAI211_X1 U21041 ( .C1(n18127), .C2(n17909), .A(n17908), .B(n17907), .ZN(
        P3_U2840) );
  AND2_X1 U21042 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17910), .ZN(
        n17930) );
  AOI22_X1 U21043 ( .A1(n9821), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n17911), 
        .B2(n17930), .ZN(n17919) );
  NOR2_X1 U21044 ( .A1(n18786), .A2(n17956), .ZN(n18019) );
  NAND2_X1 U21045 ( .A1(n9943), .A2(n18019), .ZN(n17958) );
  OAI21_X1 U21046 ( .B1(n17912), .B2(n17958), .A(n18615), .ZN(n17913) );
  NAND3_X1 U21047 ( .A1(n17914), .A2(n18137), .A3(n17913), .ZN(n17922) );
  OAI21_X1 U21048 ( .B1(n17916), .B2(n18128), .A(n17915), .ZN(n17917) );
  OAI211_X1 U21049 ( .C1(n17922), .C2(n17917), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18036), .ZN(n17918) );
  OAI211_X1 U21050 ( .C1(n17920), .C2(n18039), .A(n17919), .B(n17918), .ZN(
        P3_U2841) );
  AOI22_X1 U21051 ( .A1(n9821), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17930), 
        .B2(n17921), .ZN(n17927) );
  INV_X1 U21052 ( .A(n17922), .ZN(n17923) );
  AOI221_X1 U21053 ( .B1(n17924), .B2(n17923), .C1(n18023), .C2(n17923), .A(
        n9821), .ZN(n17931) );
  NOR3_X1 U21054 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18128), .A3(
        n18812), .ZN(n17925) );
  OAI21_X1 U21055 ( .B1(n17931), .B2(n17925), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17926) );
  OAI211_X1 U21056 ( .C1(n18039), .C2(n17928), .A(n17927), .B(n17926), .ZN(
        P3_U2842) );
  AOI22_X1 U21057 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17931), .B1(
        n17930), .B2(n17929), .ZN(n17933) );
  NAND2_X1 U21058 ( .A1(n9821), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17932) );
  OAI211_X1 U21059 ( .C1(n17934), .C2(n18039), .A(n17933), .B(n17932), .ZN(
        P3_U2843) );
  OAI21_X1 U21060 ( .B1(n18050), .B2(n17936), .A(n17935), .ZN(n18103) );
  NAND2_X1 U21061 ( .A1(n17937), .A2(n18103), .ZN(n17984) );
  AOI21_X1 U21062 ( .B1(n17938), .B2(n17984), .A(n18127), .ZN(n18032) );
  NAND2_X1 U21063 ( .A1(n9943), .A2(n18032), .ZN(n17967) );
  NAND2_X1 U21064 ( .A1(n18615), .A2(n18786), .ZN(n18108) );
  NAND3_X1 U21065 ( .A1(n17939), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18108), .ZN(n17943) );
  OAI21_X1 U21066 ( .B1(n17940), .B2(n18023), .A(n18137), .ZN(n17941) );
  AOI211_X1 U21067 ( .C1(n17944), .C2(n17943), .A(n17942), .B(n17941), .ZN(
        n17951) );
  INV_X1 U21068 ( .A(n17944), .ZN(n18107) );
  AOI221_X1 U21069 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17951), 
        .C1(n18107), .C2(n17951), .A(n9821), .ZN(n17946) );
  AOI22_X1 U21070 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17946), .B1(
        n9811), .B2(n17945), .ZN(n17948) );
  NAND2_X1 U21071 ( .A1(n9821), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17947) );
  OAI211_X1 U21072 ( .C1(n17949), .C2(n17967), .A(n17948), .B(n17947), .ZN(
        P3_U2844) );
  NOR3_X1 U21073 ( .A1(n18042), .A2(n17951), .A3(n17950), .ZN(n17953) );
  NOR3_X1 U21074 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17960), .A3(
        n17967), .ZN(n17952) );
  AOI211_X1 U21075 ( .C1(n9811), .C2(n17954), .A(n17953), .B(n17952), .ZN(
        n17955) );
  OAI21_X1 U21076 ( .B1(n18036), .B2(n18712), .A(n17955), .ZN(P3_U2845) );
  INV_X1 U21077 ( .A(n17982), .ZN(n18034) );
  AOI22_X1 U21078 ( .A1(n18613), .A2(n17957), .B1(n18131), .B2(n17956), .ZN(
        n18044) );
  OAI21_X1 U21079 ( .B1(n11303), .B2(n18615), .A(n17958), .ZN(n17959) );
  OAI211_X1 U21080 ( .C1(n18034), .C2(n17968), .A(n18044), .B(n17959), .ZN(
        n17975) );
  AOI21_X1 U21081 ( .B1(n18052), .B2(n17975), .A(n18127), .ZN(n17961) );
  AOI211_X1 U21082 ( .C1(n17962), .C2(n17961), .A(n18042), .B(n17960), .ZN(
        n17963) );
  AOI21_X1 U21083 ( .B1(n17964), .B2(n9811), .A(n17963), .ZN(n17966) );
  OAI211_X1 U21084 ( .C1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n17967), .A(
        n17966), .B(n17965), .ZN(P3_U2846) );
  INV_X1 U21085 ( .A(n17968), .ZN(n17969) );
  OAI21_X1 U21086 ( .B1(n17969), .B2(n17984), .A(n11303), .ZN(n17976) );
  AND2_X1 U21087 ( .A1(n17970), .A2(n18581), .ZN(n17973) );
  AOI222_X1 U21088 ( .A1(n17976), .A2(n17975), .B1(n17974), .B2(n17973), .C1(
        n17972), .C2(n17971), .ZN(n17980) );
  AOI22_X1 U21089 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18129), .B1(
        n9811), .B2(n17977), .ZN(n17979) );
  OAI211_X1 U21090 ( .C1(n17980), .C2(n18127), .A(n17979), .B(n17978), .ZN(
        P3_U2847) );
  AOI21_X1 U21091 ( .B1(n18006), .B2(n18019), .A(n18605), .ZN(n18002) );
  OAI211_X1 U21092 ( .C1(n18605), .C2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18044), .ZN(n17981) );
  AOI211_X1 U21093 ( .C1(n17982), .C2(n17985), .A(n18002), .B(n17981), .ZN(
        n17983) );
  AOI221_X1 U21094 ( .B1(n17985), .B2(n17987), .C1(n17984), .C2(n17987), .A(
        n17983), .ZN(n17992) );
  OAI22_X1 U21095 ( .A1(n17987), .A2(n17986), .B1(n18036), .B2(n18705), .ZN(
        n17991) );
  OAI22_X1 U21096 ( .A1(n18145), .A2(n17989), .B1(n18039), .B2(n17988), .ZN(
        n17990) );
  AOI211_X1 U21097 ( .C1(n18137), .C2(n17992), .A(n17991), .B(n17990), .ZN(
        n17993) );
  OAI21_X1 U21098 ( .B1(n18064), .B2(n17994), .A(n17993), .ZN(P3_U2848) );
  AOI22_X1 U21099 ( .A1(n9821), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18032), 
        .B2(n17995), .ZN(n18004) );
  AOI21_X1 U21100 ( .B1(n17997), .B2(n18006), .A(n17996), .ZN(n17999) );
  AOI21_X1 U21101 ( .B1(n17998), .B2(n18044), .A(n18034), .ZN(n18027) );
  AOI211_X1 U21102 ( .C1(n18581), .C2(n18000), .A(n17999), .B(n18027), .ZN(
        n18007) );
  OAI211_X1 U21103 ( .C1(n18034), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18137), .B(n18007), .ZN(n18001) );
  OAI211_X1 U21104 ( .C1(n18002), .C2(n18001), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18036), .ZN(n18003) );
  OAI211_X1 U21105 ( .C1(n18005), .C2(n18039), .A(n18004), .B(n18003), .ZN(
        P3_U2849) );
  AND2_X1 U21106 ( .A1(n18006), .A2(n18019), .ZN(n18008) );
  OAI211_X1 U21107 ( .C1(n18008), .C2(n18605), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18007), .ZN(n18012) );
  INV_X1 U21108 ( .A(n18032), .ZN(n18049) );
  OAI22_X1 U21109 ( .A1(n18010), .A2(n18049), .B1(n18009), .B2(n18127), .ZN(
        n18011) );
  AOI22_X1 U21110 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18129), .B1(
        n18012), .B2(n18011), .ZN(n18014) );
  OAI211_X1 U21111 ( .C1(n18015), .C2(n18039), .A(n18014), .B(n18013), .ZN(
        P3_U2850) );
  AOI22_X1 U21112 ( .A1(n9821), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n9811), .B2(
        n18016), .ZN(n18029) );
  OAI22_X1 U21113 ( .A1(n18605), .A2(n18019), .B1(n18018), .B2(n18017), .ZN(
        n18020) );
  AOI211_X1 U21114 ( .C1(n18022), .C2(n18021), .A(n18129), .B(n18020), .ZN(
        n18043) );
  OAI21_X1 U21115 ( .B1(n18024), .B2(n18023), .A(n18043), .ZN(n18025) );
  AOI21_X1 U21116 ( .B1(n18615), .B2(n18041), .A(n18025), .ZN(n18033) );
  OAI21_X1 U21117 ( .B1(n18605), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18033), .ZN(n18026) );
  OAI211_X1 U21118 ( .C1(n18027), .C2(n18026), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18036), .ZN(n18028) );
  OAI211_X1 U21119 ( .C1(n18049), .C2(n18030), .A(n18029), .B(n18028), .ZN(
        P3_U2851) );
  NOR2_X1 U21120 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18041), .ZN(
        n18031) );
  AOI22_X1 U21121 ( .A1(n9821), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18032), 
        .B2(n18031), .ZN(n18038) );
  OAI211_X1 U21122 ( .C1(n18034), .C2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18044), .B(n18033), .ZN(n18035) );
  NAND3_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18036), .A3(
        n18035), .ZN(n18037) );
  OAI211_X1 U21124 ( .C1(n18040), .C2(n18039), .A(n18038), .B(n18037), .ZN(
        P3_U2852) );
  AOI211_X1 U21125 ( .C1(n18044), .C2(n18043), .A(n18042), .B(n18041), .ZN(
        n18045) );
  AOI21_X1 U21126 ( .B1(n9811), .B2(n18046), .A(n18045), .ZN(n18048) );
  OAI211_X1 U21127 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18049), .A(
        n18048), .B(n18047), .ZN(P3_U2853) );
  AND3_X1 U21128 ( .A1(n18068), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        n18103), .ZN(n18055) );
  INV_X1 U21129 ( .A(n18068), .ZN(n18051) );
  NAND2_X1 U21130 ( .A1(n18613), .A2(n18050), .ZN(n18117) );
  OAI211_X1 U21131 ( .C1(n18107), .C2(n18114), .A(n18108), .B(n18117), .ZN(
        n18101) );
  AOI211_X1 U21132 ( .C1(n18052), .C2(n18051), .A(n18071), .B(n18101), .ZN(
        n18069) );
  NOR2_X1 U21133 ( .A1(n18053), .A2(n18069), .ZN(n18054) );
  MUX2_X1 U21134 ( .A(n18055), .B(n18054), .S(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Z(n18056) );
  AOI22_X1 U21135 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18129), .B1(
        n18137), .B2(n18056), .ZN(n18058) );
  OAI211_X1 U21136 ( .C1(n18059), .C2(n18145), .A(n18058), .B(n18057), .ZN(
        n18060) );
  AOI21_X1 U21137 ( .B1(n9811), .B2(n18061), .A(n18060), .ZN(n18063) );
  OAI21_X1 U21138 ( .B1(n18065), .B2(n18064), .A(n18063), .ZN(P3_U2854) );
  AOI22_X1 U21139 ( .A1(n18126), .A2(n18067), .B1(n18136), .B2(n18066), .ZN(
        n18075) );
  NAND2_X1 U21140 ( .A1(n18068), .A2(n18103), .ZN(n18070) );
  AOI211_X1 U21141 ( .C1(n18071), .C2(n18070), .A(n18069), .B(n18127), .ZN(
        n18072) );
  AOI211_X1 U21142 ( .C1(n18129), .C2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18073), .B(n18072), .ZN(n18074) );
  NAND2_X1 U21143 ( .A1(n18075), .A2(n18074), .ZN(P3_U2855) );
  NAND3_X1 U21144 ( .A1(n18137), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18103), .ZN(n18092) );
  NOR3_X1 U21145 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18077), .A3(
        n18092), .ZN(n18076) );
  AOI21_X1 U21146 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n9821), .A(n18076), .ZN(
        n18082) );
  INV_X1 U21147 ( .A(n18077), .ZN(n18079) );
  AOI221_X1 U21148 ( .B1(n18102), .B2(n18130), .C1(n18101), .C2(n18130), .A(
        n18129), .ZN(n18098) );
  OAI21_X1 U21149 ( .B1(n18079), .B2(n18078), .A(n18098), .ZN(n18087) );
  AOI22_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18087), .B1(
        n18136), .B2(n18080), .ZN(n18081) );
  OAI211_X1 U21151 ( .C1(n18083), .C2(n18145), .A(n18082), .B(n18081), .ZN(
        P3_U2856) );
  NAND2_X1 U21152 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18084), .ZN(
        n18090) );
  AOI22_X1 U21153 ( .A1(n9821), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18126), .B2(
        n18085), .ZN(n18089) );
  AOI22_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18087), .B1(
        n18136), .B2(n18086), .ZN(n18088) );
  OAI211_X1 U21155 ( .C1(n18092), .C2(n18090), .A(n18089), .B(n18088), .ZN(
        P3_U2857) );
  INV_X1 U21156 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18097) );
  AOI22_X1 U21157 ( .A1(n9821), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18136), .B2(
        n18091), .ZN(n18096) );
  INV_X1 U21158 ( .A(n18092), .ZN(n18093) );
  AOI22_X1 U21159 ( .A1(n18094), .A2(n18126), .B1(n18093), .B2(n18097), .ZN(
        n18095) );
  OAI211_X1 U21160 ( .C1(n18098), .C2(n18097), .A(n18096), .B(n18095), .ZN(
        P3_U2858) );
  AOI22_X1 U21161 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18129), .B1(
        n9821), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18106) );
  AOI22_X1 U21162 ( .A1(n18126), .A2(n18100), .B1(n18136), .B2(n18099), .ZN(
        n18105) );
  OAI221_X1 U21163 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18103), .C1(
        n18102), .C2(n18101), .A(n18137), .ZN(n18104) );
  NAND3_X1 U21164 ( .A1(n18106), .A2(n18105), .A3(n18104), .ZN(P3_U2859) );
  INV_X1 U21165 ( .A(n18588), .ZN(n18110) );
  AOI211_X1 U21166 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n18108), .A(
        n18107), .B(n18112), .ZN(n18109) );
  AOI21_X1 U21167 ( .B1(n18111), .B2(n18110), .A(n18109), .ZN(n18118) );
  NAND3_X1 U21168 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18113), .A3(
        n18112), .ZN(n18116) );
  NAND3_X1 U21169 ( .A1(n18613), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18114), .ZN(n18115) );
  NAND4_X1 U21170 ( .A1(n18118), .A2(n18117), .A3(n18116), .A4(n18115), .ZN(
        n18119) );
  AOI22_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18129), .B1(
        n18137), .B2(n18119), .ZN(n18122) );
  INV_X1 U21172 ( .A(n18120), .ZN(n18121) );
  OAI211_X1 U21173 ( .C1(n18123), .C2(n18145), .A(n18122), .B(n18121), .ZN(
        P3_U2860) );
  AOI22_X1 U21174 ( .A1(n18126), .A2(n18125), .B1(n18136), .B2(n18124), .ZN(
        n18135) );
  NAND2_X1 U21175 ( .A1(n9821), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18134) );
  NOR3_X1 U21176 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18128), .A3(
        n18127), .ZN(n18139) );
  OAI21_X1 U21177 ( .B1(n18129), .B2(n18139), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18133) );
  OAI211_X1 U21178 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18131), .A(
        n18130), .B(n18767), .ZN(n18132) );
  NAND4_X1 U21179 ( .A1(n18135), .A2(n18134), .A3(n18133), .A4(n18132), .ZN(
        P3_U2861) );
  INV_X1 U21180 ( .A(n18136), .ZN(n18143) );
  AOI21_X1 U21181 ( .B1(n18617), .B2(n18137), .A(n18786), .ZN(n18138) );
  NOR2_X1 U21182 ( .A1(n18139), .A2(n18138), .ZN(n18141) );
  INV_X1 U21183 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18140) );
  MUX2_X1 U21184 ( .A(n18141), .B(n18140), .S(n9821), .Z(n18142) );
  OAI221_X1 U21185 ( .B1(n18146), .B2(n18145), .C1(n18144), .C2(n18143), .A(
        n18142), .ZN(P3_U2862) );
  OAI211_X1 U21186 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18147), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18148)
         );
  INV_X1 U21187 ( .A(n18148), .ZN(n18646) );
  OAI21_X1 U21188 ( .B1(n18646), .B2(n18149), .A(n18154), .ZN(n18150) );
  OAI221_X1 U21189 ( .B1(n18621), .B2(n18803), .C1(n18621), .C2(n18154), .A(
        n18150), .ZN(P3_U2863) );
  INV_X1 U21190 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18631) );
  NOR2_X1 U21191 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18631), .ZN(
        n18447) );
  NOR2_X1 U21192 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18628), .ZN(
        n18330) );
  NOR2_X1 U21193 ( .A1(n18447), .A2(n18330), .ZN(n18152) );
  OAI22_X1 U21194 ( .A1(n18153), .A2(n18631), .B1(n18152), .B2(n18151), .ZN(
        P3_U2866) );
  NOR2_X1 U21195 ( .A1(n18632), .A2(n18154), .ZN(P3_U2867) );
  NOR2_X1 U21196 ( .A1(n18156), .A2(n18155), .ZN(n18189) );
  NAND2_X1 U21197 ( .A1(n18189), .A2(n18157), .ZN(n18533) );
  NAND2_X1 U21198 ( .A1(n18623), .A2(n18621), .ZN(n18624) );
  INV_X1 U21199 ( .A(n18624), .ZN(n18350) );
  NOR2_X1 U21200 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18240) );
  NAND2_X1 U21201 ( .A1(n18350), .A2(n18240), .ZN(n18216) );
  NOR2_X2 U21202 ( .A1(n18497), .A2(n18158), .ZN(n18525) );
  NOR2_X1 U21203 ( .A1(n18631), .A2(n18328), .ZN(n18527) );
  NAND2_X1 U21204 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18527), .ZN(
        n18579) );
  AOI21_X1 U21205 ( .B1(n18579), .B2(n18216), .A(n18523), .ZN(n18192) );
  AND2_X1 U21206 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18529), .ZN(n18524) );
  NAND2_X1 U21207 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18160) );
  NOR2_X1 U21208 ( .A1(n18160), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18528) );
  INV_X1 U21209 ( .A(n18528), .ZN(n18473) );
  NOR2_X2 U21210 ( .A1(n18621), .A2(n18473), .ZN(n18570) );
  AOI22_X1 U21211 ( .A1(n18525), .A2(n18192), .B1(n18524), .B2(n18570), .ZN(
        n18163) );
  NOR2_X1 U21212 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18623), .ZN(
        n18397) );
  NOR2_X1 U21213 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18621), .ZN(
        n18374) );
  NOR2_X1 U21214 ( .A1(n18397), .A2(n18374), .ZN(n18450) );
  NOR2_X1 U21215 ( .A1(n18450), .A2(n18160), .ZN(n18495) );
  AOI21_X1 U21216 ( .B1(n18579), .B2(n18216), .A(n18497), .ZN(n18217) );
  NAND2_X1 U21217 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18159) );
  AOI22_X1 U21218 ( .A1(n18529), .A2(n18495), .B1(n18217), .B2(n18159), .ZN(
        n18193) );
  AND2_X1 U21219 ( .A1(n18529), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18530) );
  INV_X1 U21220 ( .A(n18397), .ZN(n18161) );
  NOR2_X2 U21221 ( .A1(n18161), .A2(n18160), .ZN(n18501) );
  AOI22_X1 U21222 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18193), .B1(
        n18530), .B2(n18501), .ZN(n18162) );
  OAI211_X1 U21223 ( .C1(n18533), .C2(n18216), .A(n18163), .B(n18162), .ZN(
        P3_U2868) );
  NAND2_X1 U21224 ( .A1(n18189), .A2(n18164), .ZN(n18539) );
  NOR2_X2 U21225 ( .A1(n14843), .A2(n18498), .ZN(n18536) );
  AND2_X1 U21226 ( .A1(n18452), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18534) );
  AOI22_X1 U21227 ( .A1(n18536), .A2(n18570), .B1(n18534), .B2(n18192), .ZN(
        n18166) );
  AND2_X1 U21228 ( .A1(n18529), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18535) );
  AOI22_X1 U21229 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18193), .B1(
        n18535), .B2(n18501), .ZN(n18165) );
  OAI211_X1 U21230 ( .C1(n18539), .C2(n18216), .A(n18166), .B(n18165), .ZN(
        P3_U2869) );
  NAND2_X1 U21231 ( .A1(n18189), .A2(n18167), .ZN(n18545) );
  AND2_X1 U21232 ( .A1(n18529), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18541) );
  NOR2_X2 U21233 ( .A1(n18497), .A2(n18168), .ZN(n18540) );
  AOI22_X1 U21234 ( .A1(n18541), .A2(n18501), .B1(n18540), .B2(n18192), .ZN(
        n18170) );
  AND2_X1 U21235 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18529), .ZN(n18542) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18193), .B1(
        n18542), .B2(n18570), .ZN(n18169) );
  OAI211_X1 U21237 ( .C1(n18545), .C2(n18216), .A(n18170), .B(n18169), .ZN(
        P3_U2870) );
  INV_X1 U21238 ( .A(n18171), .ZN(n18172) );
  NAND2_X1 U21239 ( .A1(n18189), .A2(n18172), .ZN(n18551) );
  AND2_X1 U21240 ( .A1(n18529), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18547) );
  NOR2_X2 U21241 ( .A1(n18497), .A2(n18173), .ZN(n18546) );
  AOI22_X1 U21242 ( .A1(n18547), .A2(n18501), .B1(n18546), .B2(n18192), .ZN(
        n18175) );
  AND2_X1 U21243 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18529), .ZN(n18548) );
  AOI22_X1 U21244 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18193), .B1(
        n18548), .B2(n18570), .ZN(n18174) );
  OAI211_X1 U21245 ( .C1(n18551), .C2(n18216), .A(n18175), .B(n18174), .ZN(
        P3_U2871) );
  NAND2_X1 U21246 ( .A1(n18189), .A2(n18176), .ZN(n18557) );
  NOR2_X2 U21247 ( .A1(n18497), .A2(n18177), .ZN(n18553) );
  AND2_X1 U21248 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18529), .ZN(n18552) );
  AOI22_X1 U21249 ( .A1(n18553), .A2(n18192), .B1(n18552), .B2(n18570), .ZN(
        n18179) );
  AND2_X1 U21250 ( .A1(n18529), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18554) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18193), .B1(
        n18554), .B2(n18501), .ZN(n18178) );
  OAI211_X1 U21252 ( .C1(n18557), .C2(n18216), .A(n18179), .B(n18178), .ZN(
        P3_U2872) );
  NAND2_X1 U21253 ( .A1(n18189), .A2(n18180), .ZN(n18563) );
  AND2_X1 U21254 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18529), .ZN(n18560) );
  NOR2_X2 U21255 ( .A1(n18497), .A2(n18181), .ZN(n18559) );
  AOI22_X1 U21256 ( .A1(n18560), .A2(n18570), .B1(n18559), .B2(n18192), .ZN(
        n18183) );
  NOR2_X2 U21257 ( .A1(n18498), .A2(n14875), .ZN(n18558) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18193), .B1(
        n18558), .B2(n18501), .ZN(n18182) );
  OAI211_X1 U21259 ( .C1(n18563), .C2(n18216), .A(n18183), .B(n18182), .ZN(
        P3_U2873) );
  NAND2_X1 U21260 ( .A1(n18189), .A2(n18184), .ZN(n18569) );
  NOR2_X2 U21261 ( .A1(n18497), .A2(n18185), .ZN(n18565) );
  AND2_X1 U21262 ( .A1(n18529), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18564) );
  AOI22_X1 U21263 ( .A1(n18565), .A2(n18192), .B1(n18564), .B2(n18501), .ZN(
        n18187) );
  AND2_X1 U21264 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18529), .ZN(n18566) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18193), .B1(
        n18566), .B2(n18570), .ZN(n18186) );
  OAI211_X1 U21266 ( .C1(n18569), .C2(n18216), .A(n18187), .B(n18186), .ZN(
        P3_U2874) );
  NAND2_X1 U21267 ( .A1(n18189), .A2(n18188), .ZN(n18580) );
  NOR2_X2 U21268 ( .A1(n18498), .A2(n18190), .ZN(n18575) );
  NOR2_X2 U21269 ( .A1(n18191), .A2(n18497), .ZN(n18573) );
  AOI22_X1 U21270 ( .A1(n18575), .A2(n18570), .B1(n18573), .B2(n18192), .ZN(
        n18195) );
  NOR2_X2 U21271 ( .A1(n14866), .A2(n18498), .ZN(n18571) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18193), .B1(
        n18571), .B2(n18501), .ZN(n18194) );
  OAI211_X1 U21273 ( .C1(n18580), .C2(n18216), .A(n18195), .B(n18194), .ZN(
        P3_U2875) );
  NAND2_X1 U21274 ( .A1(n18374), .A2(n18240), .ZN(n18239) );
  INV_X1 U21275 ( .A(n18240), .ZN(n18196) );
  AOI22_X1 U21276 ( .A1(n18525), .A2(n18212), .B1(n18524), .B2(n18501), .ZN(
        n18199) );
  NAND2_X1 U21277 ( .A1(n18452), .A2(n18197), .ZN(n18376) );
  NOR2_X1 U21278 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18376), .ZN(
        n18286) );
  AOI22_X1 U21279 ( .A1(n18529), .A2(n18527), .B1(n18240), .B2(n18286), .ZN(
        n18213) );
  INV_X1 U21280 ( .A(n18579), .ZN(n18234) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18213), .B1(
        n18530), .B2(n18234), .ZN(n18198) );
  OAI211_X1 U21282 ( .C1(n18533), .C2(n18239), .A(n18199), .B(n18198), .ZN(
        P3_U2876) );
  AOI22_X1 U21283 ( .A1(n18535), .A2(n18234), .B1(n18534), .B2(n18212), .ZN(
        n18201) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18213), .B1(
        n18536), .B2(n18501), .ZN(n18200) );
  OAI211_X1 U21285 ( .C1(n18539), .C2(n18239), .A(n18201), .B(n18200), .ZN(
        P3_U2877) );
  AOI22_X1 U21286 ( .A1(n18540), .A2(n18212), .B1(n18542), .B2(n18501), .ZN(
        n18203) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18213), .B1(
        n18541), .B2(n18234), .ZN(n18202) );
  OAI211_X1 U21288 ( .C1(n18545), .C2(n18239), .A(n18203), .B(n18202), .ZN(
        P3_U2878) );
  AOI22_X1 U21289 ( .A1(n18546), .A2(n18212), .B1(n18548), .B2(n18501), .ZN(
        n18205) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18213), .B1(
        n18547), .B2(n18234), .ZN(n18204) );
  OAI211_X1 U21291 ( .C1(n18551), .C2(n18239), .A(n18205), .B(n18204), .ZN(
        P3_U2879) );
  AOI22_X1 U21292 ( .A1(n18554), .A2(n18234), .B1(n18553), .B2(n18212), .ZN(
        n18207) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18213), .B1(
        n18552), .B2(n18501), .ZN(n18206) );
  OAI211_X1 U21294 ( .C1(n18557), .C2(n18239), .A(n18207), .B(n18206), .ZN(
        P3_U2880) );
  AOI22_X1 U21295 ( .A1(n18560), .A2(n18501), .B1(n18559), .B2(n18212), .ZN(
        n18209) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18213), .B1(
        n18558), .B2(n18234), .ZN(n18208) );
  OAI211_X1 U21297 ( .C1(n18563), .C2(n18239), .A(n18209), .B(n18208), .ZN(
        P3_U2881) );
  AOI22_X1 U21298 ( .A1(n18565), .A2(n18212), .B1(n18564), .B2(n18234), .ZN(
        n18211) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18213), .B1(
        n18566), .B2(n18501), .ZN(n18210) );
  OAI211_X1 U21300 ( .C1(n18569), .C2(n18239), .A(n18211), .B(n18210), .ZN(
        P3_U2882) );
  AOI22_X1 U21301 ( .A1(n18573), .A2(n18212), .B1(n18571), .B2(n18234), .ZN(
        n18215) );
  AOI22_X1 U21302 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18213), .B1(
        n18575), .B2(n18501), .ZN(n18214) );
  OAI211_X1 U21303 ( .C1(n18580), .C2(n18239), .A(n18215), .B(n18214), .ZN(
        P3_U2883) );
  NAND2_X1 U21304 ( .A1(n18397), .A2(n18240), .ZN(n18238) );
  INV_X1 U21305 ( .A(n18216), .ZN(n18256) );
  AOI21_X1 U21306 ( .B1(n18239), .B2(n18238), .A(n18523), .ZN(n18233) );
  AOI22_X1 U21307 ( .A1(n18530), .A2(n18256), .B1(n18525), .B2(n18233), .ZN(
        n18220) );
  INV_X1 U21308 ( .A(n18238), .ZN(n18303) );
  AOI21_X1 U21309 ( .B1(n18239), .B2(n18238), .A(n18497), .ZN(n18261) );
  AND2_X1 U21310 ( .A1(n18448), .A2(n18217), .ZN(n18218) );
  OAI22_X1 U21311 ( .A1(n18303), .A2(n18758), .B1(n18261), .B2(n18218), .ZN(
        n18235) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18235), .B1(
        n18524), .B2(n18234), .ZN(n18219) );
  OAI211_X1 U21313 ( .C1(n18533), .C2(n18238), .A(n18220), .B(n18219), .ZN(
        P3_U2884) );
  AOI22_X1 U21314 ( .A1(n18535), .A2(n18256), .B1(n18534), .B2(n18233), .ZN(
        n18222) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18235), .B1(
        n18536), .B2(n18234), .ZN(n18221) );
  OAI211_X1 U21316 ( .C1(n18539), .C2(n18238), .A(n18222), .B(n18221), .ZN(
        P3_U2885) );
  AOI22_X1 U21317 ( .A1(n18540), .A2(n18233), .B1(n18542), .B2(n18234), .ZN(
        n18224) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18235), .B1(
        n18541), .B2(n18256), .ZN(n18223) );
  OAI211_X1 U21319 ( .C1(n18545), .C2(n18238), .A(n18224), .B(n18223), .ZN(
        P3_U2886) );
  AOI22_X1 U21320 ( .A1(n18546), .A2(n18233), .B1(n18548), .B2(n18234), .ZN(
        n18226) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18235), .B1(
        n18547), .B2(n18256), .ZN(n18225) );
  OAI211_X1 U21322 ( .C1(n18551), .C2(n18238), .A(n18226), .B(n18225), .ZN(
        P3_U2887) );
  AOI22_X1 U21323 ( .A1(n18554), .A2(n18256), .B1(n18553), .B2(n18233), .ZN(
        n18228) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18235), .B1(
        n18552), .B2(n18234), .ZN(n18227) );
  OAI211_X1 U21325 ( .C1(n18557), .C2(n18238), .A(n18228), .B(n18227), .ZN(
        P3_U2888) );
  AOI22_X1 U21326 ( .A1(n18559), .A2(n18233), .B1(n18558), .B2(n18256), .ZN(
        n18230) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18235), .B1(
        n18560), .B2(n18234), .ZN(n18229) );
  OAI211_X1 U21328 ( .C1(n18563), .C2(n18238), .A(n18230), .B(n18229), .ZN(
        P3_U2889) );
  AOI22_X1 U21329 ( .A1(n18566), .A2(n18234), .B1(n18565), .B2(n18233), .ZN(
        n18232) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18235), .B1(
        n18564), .B2(n18256), .ZN(n18231) );
  OAI211_X1 U21331 ( .C1(n18569), .C2(n18238), .A(n18232), .B(n18231), .ZN(
        P3_U2890) );
  AOI22_X1 U21332 ( .A1(n18573), .A2(n18233), .B1(n18571), .B2(n18256), .ZN(
        n18237) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18235), .B1(
        n18575), .B2(n18234), .ZN(n18236) );
  OAI211_X1 U21334 ( .C1(n18580), .C2(n18238), .A(n18237), .B(n18236), .ZN(
        P3_U2891) );
  NAND2_X1 U21335 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18240), .ZN(
        n18285) );
  NOR2_X2 U21336 ( .A1(n18621), .A2(n18285), .ZN(n18324) );
  INV_X1 U21337 ( .A(n18324), .ZN(n18260) );
  INV_X1 U21338 ( .A(n18239), .ZN(n18279) );
  NOR2_X1 U21339 ( .A1(n18523), .A2(n18285), .ZN(n18255) );
  AOI22_X1 U21340 ( .A1(n18530), .A2(n18279), .B1(n18525), .B2(n18255), .ZN(
        n18242) );
  AOI21_X1 U21341 ( .B1(n18623), .B2(n18401), .A(n18376), .ZN(n18329) );
  NAND2_X1 U21342 ( .A1(n18240), .A2(n18329), .ZN(n18257) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18257), .B1(
        n18524), .B2(n18256), .ZN(n18241) );
  OAI211_X1 U21344 ( .C1(n18260), .C2(n18533), .A(n18242), .B(n18241), .ZN(
        P3_U2892) );
  AOI22_X1 U21345 ( .A1(n18536), .A2(n18256), .B1(n18534), .B2(n18255), .ZN(
        n18244) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18257), .B1(
        n18535), .B2(n18279), .ZN(n18243) );
  OAI211_X1 U21347 ( .C1(n18260), .C2(n18539), .A(n18244), .B(n18243), .ZN(
        P3_U2893) );
  AOI22_X1 U21348 ( .A1(n18540), .A2(n18255), .B1(n18542), .B2(n18256), .ZN(
        n18246) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18257), .B1(
        n18541), .B2(n18279), .ZN(n18245) );
  OAI211_X1 U21350 ( .C1(n18260), .C2(n18545), .A(n18246), .B(n18245), .ZN(
        P3_U2894) );
  AOI22_X1 U21351 ( .A1(n18547), .A2(n18279), .B1(n18546), .B2(n18255), .ZN(
        n18248) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18257), .B1(
        n18548), .B2(n18256), .ZN(n18247) );
  OAI211_X1 U21353 ( .C1(n18260), .C2(n18551), .A(n18248), .B(n18247), .ZN(
        P3_U2895) );
  AOI22_X1 U21354 ( .A1(n18553), .A2(n18255), .B1(n18552), .B2(n18256), .ZN(
        n18250) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18257), .B1(
        n18554), .B2(n18279), .ZN(n18249) );
  OAI211_X1 U21356 ( .C1(n18260), .C2(n18557), .A(n18250), .B(n18249), .ZN(
        P3_U2896) );
  AOI22_X1 U21357 ( .A1(n18559), .A2(n18255), .B1(n18558), .B2(n18279), .ZN(
        n18252) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18257), .B1(
        n18560), .B2(n18256), .ZN(n18251) );
  OAI211_X1 U21359 ( .C1(n18260), .C2(n18563), .A(n18252), .B(n18251), .ZN(
        P3_U2897) );
  AOI22_X1 U21360 ( .A1(n18565), .A2(n18255), .B1(n18564), .B2(n18279), .ZN(
        n18254) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18257), .B1(
        n18566), .B2(n18256), .ZN(n18253) );
  OAI211_X1 U21362 ( .C1(n18260), .C2(n18569), .A(n18254), .B(n18253), .ZN(
        P3_U2898) );
  AOI22_X1 U21363 ( .A1(n18573), .A2(n18255), .B1(n18571), .B2(n18279), .ZN(
        n18259) );
  AOI22_X1 U21364 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18257), .B1(
        n18575), .B2(n18256), .ZN(n18258) );
  OAI211_X1 U21365 ( .C1(n18260), .C2(n18580), .A(n18259), .B(n18258), .ZN(
        P3_U2899) );
  INV_X1 U21366 ( .A(n18330), .ZN(n18284) );
  NOR2_X2 U21367 ( .A1(n18624), .A2(n18284), .ZN(n18346) );
  INV_X1 U21368 ( .A(n18346), .ZN(n18283) );
  NOR2_X1 U21369 ( .A1(n18346), .A2(n18324), .ZN(n18307) );
  NOR2_X1 U21370 ( .A1(n18523), .A2(n18307), .ZN(n18278) );
  AOI22_X1 U21371 ( .A1(n18525), .A2(n18278), .B1(n18524), .B2(n18279), .ZN(
        n18265) );
  INV_X1 U21372 ( .A(n18261), .ZN(n18262) );
  OAI22_X1 U21373 ( .A1(n18307), .A2(n18497), .B1(n18401), .B2(n18262), .ZN(
        n18263) );
  OAI21_X1 U21374 ( .B1(n18346), .B2(n18758), .A(n18263), .ZN(n18280) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18280), .B1(
        n18530), .B2(n18303), .ZN(n18264) );
  OAI211_X1 U21376 ( .C1(n18283), .C2(n18533), .A(n18265), .B(n18264), .ZN(
        P3_U2900) );
  AOI22_X1 U21377 ( .A1(n18536), .A2(n18279), .B1(n18534), .B2(n18278), .ZN(
        n18267) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18280), .B1(
        n18535), .B2(n18303), .ZN(n18266) );
  OAI211_X1 U21379 ( .C1(n18283), .C2(n18539), .A(n18267), .B(n18266), .ZN(
        P3_U2901) );
  AOI22_X1 U21380 ( .A1(n18540), .A2(n18278), .B1(n18542), .B2(n18279), .ZN(
        n18269) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18280), .B1(
        n18541), .B2(n18303), .ZN(n18268) );
  OAI211_X1 U21382 ( .C1(n18283), .C2(n18545), .A(n18269), .B(n18268), .ZN(
        P3_U2902) );
  AOI22_X1 U21383 ( .A1(n18547), .A2(n18303), .B1(n18546), .B2(n18278), .ZN(
        n18271) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18280), .B1(
        n18548), .B2(n18279), .ZN(n18270) );
  OAI211_X1 U21385 ( .C1(n18283), .C2(n18551), .A(n18271), .B(n18270), .ZN(
        P3_U2903) );
  AOI22_X1 U21386 ( .A1(n18554), .A2(n18303), .B1(n18553), .B2(n18278), .ZN(
        n18273) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18280), .B1(
        n18552), .B2(n18279), .ZN(n18272) );
  OAI211_X1 U21388 ( .C1(n18283), .C2(n18557), .A(n18273), .B(n18272), .ZN(
        P3_U2904) );
  AOI22_X1 U21389 ( .A1(n18559), .A2(n18278), .B1(n18558), .B2(n18303), .ZN(
        n18275) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18280), .B1(
        n18560), .B2(n18279), .ZN(n18274) );
  OAI211_X1 U21391 ( .C1(n18283), .C2(n18563), .A(n18275), .B(n18274), .ZN(
        P3_U2905) );
  AOI22_X1 U21392 ( .A1(n18565), .A2(n18278), .B1(n18564), .B2(n18303), .ZN(
        n18277) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18280), .B1(
        n18566), .B2(n18279), .ZN(n18276) );
  OAI211_X1 U21394 ( .C1(n18283), .C2(n18569), .A(n18277), .B(n18276), .ZN(
        P3_U2906) );
  AOI22_X1 U21395 ( .A1(n18575), .A2(n18279), .B1(n18573), .B2(n18278), .ZN(
        n18282) );
  AOI22_X1 U21396 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18280), .B1(
        n18571), .B2(n18303), .ZN(n18281) );
  OAI211_X1 U21397 ( .C1(n18283), .C2(n18580), .A(n18282), .B(n18281), .ZN(
        P3_U2907) );
  NAND2_X1 U21398 ( .A1(n18330), .A2(n18374), .ZN(n18351) );
  AOI22_X1 U21399 ( .A1(n18530), .A2(n18324), .B1(n18525), .B2(n18302), .ZN(
        n18289) );
  INV_X1 U21400 ( .A(n18285), .ZN(n18287) );
  AOI22_X1 U21401 ( .A1(n18529), .A2(n18287), .B1(n18330), .B2(n18286), .ZN(
        n18304) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18304), .B1(
        n18524), .B2(n18303), .ZN(n18288) );
  OAI211_X1 U21403 ( .C1(n18351), .C2(n18533), .A(n18289), .B(n18288), .ZN(
        P3_U2908) );
  AOI22_X1 U21404 ( .A1(n18324), .A2(n18535), .B1(n18534), .B2(n18302), .ZN(
        n18291) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18304), .B1(
        n18536), .B2(n18303), .ZN(n18290) );
  OAI211_X1 U21406 ( .C1(n18351), .C2(n18539), .A(n18291), .B(n18290), .ZN(
        P3_U2909) );
  AOI22_X1 U21407 ( .A1(n18540), .A2(n18302), .B1(n18542), .B2(n18303), .ZN(
        n18293) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18541), .ZN(n18292) );
  OAI211_X1 U21409 ( .C1(n18351), .C2(n18545), .A(n18293), .B(n18292), .ZN(
        P3_U2910) );
  AOI22_X1 U21410 ( .A1(n18546), .A2(n18302), .B1(n18548), .B2(n18303), .ZN(
        n18295) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18547), .ZN(n18294) );
  OAI211_X1 U21412 ( .C1(n18351), .C2(n18551), .A(n18295), .B(n18294), .ZN(
        P3_U2911) );
  AOI22_X1 U21413 ( .A1(n18553), .A2(n18302), .B1(n18552), .B2(n18303), .ZN(
        n18297) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18554), .ZN(n18296) );
  OAI211_X1 U21415 ( .C1(n18351), .C2(n18557), .A(n18297), .B(n18296), .ZN(
        P3_U2912) );
  AOI22_X1 U21416 ( .A1(n18560), .A2(n18303), .B1(n18559), .B2(n18302), .ZN(
        n18299) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18558), .ZN(n18298) );
  OAI211_X1 U21418 ( .C1(n18351), .C2(n18563), .A(n18299), .B(n18298), .ZN(
        P3_U2913) );
  AOI22_X1 U21419 ( .A1(n18566), .A2(n18303), .B1(n18565), .B2(n18302), .ZN(
        n18301) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18564), .ZN(n18300) );
  OAI211_X1 U21421 ( .C1(n18351), .C2(n18569), .A(n18301), .B(n18300), .ZN(
        P3_U2914) );
  AOI22_X1 U21422 ( .A1(n18575), .A2(n18303), .B1(n18573), .B2(n18302), .ZN(
        n18306) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18304), .B1(
        n18324), .B2(n18571), .ZN(n18305) );
  OAI211_X1 U21424 ( .C1(n18351), .C2(n18580), .A(n18306), .B(n18305), .ZN(
        P3_U2915) );
  NAND2_X1 U21425 ( .A1(n18330), .A2(n18397), .ZN(n18352) );
  AOI21_X1 U21426 ( .B1(n18352), .B2(n18351), .A(n18523), .ZN(n18323) );
  AOI22_X1 U21427 ( .A1(n18324), .A2(n18524), .B1(n18525), .B2(n18323), .ZN(
        n18310) );
  INV_X1 U21428 ( .A(n18352), .ZN(n18393) );
  AOI221_X1 U21429 ( .B1(n18307), .B2(n18351), .C1(n18401), .C2(n18351), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18308) );
  OAI21_X1 U21430 ( .B1(n18393), .B2(n18308), .A(n18452), .ZN(n18325) );
  AOI22_X1 U21431 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18325), .B1(
        n18530), .B2(n18346), .ZN(n18309) );
  OAI211_X1 U21432 ( .C1(n18352), .C2(n18533), .A(n18310), .B(n18309), .ZN(
        P3_U2916) );
  AOI22_X1 U21433 ( .A1(n18346), .A2(n18535), .B1(n18323), .B2(n18534), .ZN(
        n18312) );
  AOI22_X1 U21434 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18536), .ZN(n18311) );
  OAI211_X1 U21435 ( .C1(n18352), .C2(n18539), .A(n18312), .B(n18311), .ZN(
        P3_U2917) );
  AOI22_X1 U21436 ( .A1(n18324), .A2(n18542), .B1(n18323), .B2(n18540), .ZN(
        n18314) );
  AOI22_X1 U21437 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18541), .ZN(n18313) );
  OAI211_X1 U21438 ( .C1(n18352), .C2(n18545), .A(n18314), .B(n18313), .ZN(
        P3_U2918) );
  AOI22_X1 U21439 ( .A1(n18324), .A2(n18548), .B1(n18323), .B2(n18546), .ZN(
        n18316) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18547), .ZN(n18315) );
  OAI211_X1 U21441 ( .C1(n18352), .C2(n18551), .A(n18316), .B(n18315), .ZN(
        P3_U2919) );
  AOI22_X1 U21442 ( .A1(n18324), .A2(n18552), .B1(n18323), .B2(n18553), .ZN(
        n18318) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18325), .B1(
        n18346), .B2(n18554), .ZN(n18317) );
  OAI211_X1 U21444 ( .C1(n18352), .C2(n18557), .A(n18318), .B(n18317), .ZN(
        P3_U2920) );
  AOI22_X1 U21445 ( .A1(n18346), .A2(n18558), .B1(n18323), .B2(n18559), .ZN(
        n18320) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18560), .ZN(n18319) );
  OAI211_X1 U21447 ( .C1(n18352), .C2(n18563), .A(n18320), .B(n18319), .ZN(
        P3_U2921) );
  AOI22_X1 U21448 ( .A1(n18346), .A2(n18564), .B1(n18323), .B2(n18565), .ZN(
        n18322) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18566), .ZN(n18321) );
  OAI211_X1 U21450 ( .C1(n18352), .C2(n18569), .A(n18322), .B(n18321), .ZN(
        P3_U2922) );
  AOI22_X1 U21451 ( .A1(n18346), .A2(n18571), .B1(n18323), .B2(n18573), .ZN(
        n18327) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18575), .ZN(n18326) );
  OAI211_X1 U21453 ( .C1(n18352), .C2(n18580), .A(n18327), .B(n18326), .ZN(
        P3_U2923) );
  NOR2_X1 U21454 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18328), .ZN(
        n18377) );
  NAND2_X1 U21455 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18377), .ZN(
        n18375) );
  INV_X1 U21456 ( .A(n18351), .ZN(n18369) );
  AOI22_X1 U21457 ( .A1(n18530), .A2(n18369), .B1(n18525), .B2(n18345), .ZN(
        n18332) );
  NAND2_X1 U21458 ( .A1(n18330), .A2(n18329), .ZN(n18347) );
  AOI22_X1 U21459 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18524), .ZN(n18331) );
  OAI211_X1 U21460 ( .C1(n18533), .C2(n18375), .A(n18332), .B(n18331), .ZN(
        P3_U2924) );
  AOI22_X1 U21461 ( .A1(n18346), .A2(n18536), .B1(n18534), .B2(n18345), .ZN(
        n18334) );
  AOI22_X1 U21462 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18347), .B1(
        n18369), .B2(n18535), .ZN(n18333) );
  OAI211_X1 U21463 ( .C1(n18539), .C2(n18375), .A(n18334), .B(n18333), .ZN(
        P3_U2925) );
  AOI22_X1 U21464 ( .A1(n18369), .A2(n18541), .B1(n18540), .B2(n18345), .ZN(
        n18336) );
  AOI22_X1 U21465 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18542), .ZN(n18335) );
  OAI211_X1 U21466 ( .C1(n18545), .C2(n18375), .A(n18336), .B(n18335), .ZN(
        P3_U2926) );
  AOI22_X1 U21467 ( .A1(n18369), .A2(n18547), .B1(n18546), .B2(n18345), .ZN(
        n18338) );
  AOI22_X1 U21468 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18548), .ZN(n18337) );
  OAI211_X1 U21469 ( .C1(n18551), .C2(n18375), .A(n18338), .B(n18337), .ZN(
        P3_U2927) );
  AOI22_X1 U21470 ( .A1(n18369), .A2(n18554), .B1(n18553), .B2(n18345), .ZN(
        n18340) );
  AOI22_X1 U21471 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18552), .ZN(n18339) );
  OAI211_X1 U21472 ( .C1(n18557), .C2(n18375), .A(n18340), .B(n18339), .ZN(
        P3_U2928) );
  AOI22_X1 U21473 ( .A1(n18346), .A2(n18560), .B1(n18559), .B2(n18345), .ZN(
        n18342) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18347), .B1(
        n18369), .B2(n18558), .ZN(n18341) );
  OAI211_X1 U21475 ( .C1(n18563), .C2(n18375), .A(n18342), .B(n18341), .ZN(
        P3_U2929) );
  AOI22_X1 U21476 ( .A1(n18369), .A2(n18564), .B1(n18565), .B2(n18345), .ZN(
        n18344) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18566), .ZN(n18343) );
  OAI211_X1 U21478 ( .C1(n18569), .C2(n18375), .A(n18344), .B(n18343), .ZN(
        P3_U2930) );
  AOI22_X1 U21479 ( .A1(n18369), .A2(n18571), .B1(n18573), .B2(n18345), .ZN(
        n18349) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18347), .B1(
        n18346), .B2(n18575), .ZN(n18348) );
  OAI211_X1 U21481 ( .C1(n18580), .C2(n18375), .A(n18349), .B(n18348), .ZN(
        P3_U2931) );
  NAND2_X1 U21482 ( .A1(n18350), .A2(n18447), .ZN(n18373) );
  AOI21_X1 U21483 ( .B1(n18375), .B2(n18373), .A(n18523), .ZN(n18368) );
  AOI22_X1 U21484 ( .A1(n18530), .A2(n18393), .B1(n18525), .B2(n18368), .ZN(
        n18355) );
  INV_X1 U21485 ( .A(n18373), .ZN(n18442) );
  AOI21_X1 U21486 ( .B1(n18375), .B2(n18373), .A(n18497), .ZN(n18399) );
  AOI21_X1 U21487 ( .B1(n18352), .B2(n18351), .A(n18498), .ZN(n18353) );
  OAI22_X1 U21488 ( .A1(n18442), .A2(n18758), .B1(n18399), .B2(n18353), .ZN(
        n18370) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18370), .B1(
        n18369), .B2(n18524), .ZN(n18354) );
  OAI211_X1 U21490 ( .C1(n18533), .C2(n18373), .A(n18355), .B(n18354), .ZN(
        P3_U2932) );
  AOI22_X1 U21491 ( .A1(n18393), .A2(n18535), .B1(n18534), .B2(n18368), .ZN(
        n18357) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18370), .B1(
        n18369), .B2(n18536), .ZN(n18356) );
  OAI211_X1 U21493 ( .C1(n18539), .C2(n18373), .A(n18357), .B(n18356), .ZN(
        P3_U2933) );
  AOI22_X1 U21494 ( .A1(n18369), .A2(n18542), .B1(n18540), .B2(n18368), .ZN(
        n18359) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18370), .B1(
        n18393), .B2(n18541), .ZN(n18358) );
  OAI211_X1 U21496 ( .C1(n18545), .C2(n18373), .A(n18359), .B(n18358), .ZN(
        P3_U2934) );
  AOI22_X1 U21497 ( .A1(n18393), .A2(n18547), .B1(n18546), .B2(n18368), .ZN(
        n18361) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18370), .B1(
        n18369), .B2(n18548), .ZN(n18360) );
  OAI211_X1 U21499 ( .C1(n18551), .C2(n18373), .A(n18361), .B(n18360), .ZN(
        P3_U2935) );
  AOI22_X1 U21500 ( .A1(n18393), .A2(n18554), .B1(n18553), .B2(n18368), .ZN(
        n18363) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18370), .B1(
        n18369), .B2(n18552), .ZN(n18362) );
  OAI211_X1 U21502 ( .C1(n18557), .C2(n18373), .A(n18363), .B(n18362), .ZN(
        P3_U2936) );
  AOI22_X1 U21503 ( .A1(n18393), .A2(n18558), .B1(n18559), .B2(n18368), .ZN(
        n18365) );
  AOI22_X1 U21504 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18370), .B1(
        n18369), .B2(n18560), .ZN(n18364) );
  OAI211_X1 U21505 ( .C1(n18563), .C2(n18373), .A(n18365), .B(n18364), .ZN(
        P3_U2937) );
  AOI22_X1 U21506 ( .A1(n18369), .A2(n18566), .B1(n18565), .B2(n18368), .ZN(
        n18367) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18370), .B1(
        n18393), .B2(n18564), .ZN(n18366) );
  OAI211_X1 U21508 ( .C1(n18569), .C2(n18373), .A(n18367), .B(n18366), .ZN(
        P3_U2938) );
  AOI22_X1 U21509 ( .A1(n18369), .A2(n18575), .B1(n18573), .B2(n18368), .ZN(
        n18372) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18370), .B1(
        n18393), .B2(n18571), .ZN(n18371) );
  OAI211_X1 U21511 ( .C1(n18580), .C2(n18373), .A(n18372), .B(n18371), .ZN(
        P3_U2939) );
  NAND2_X1 U21512 ( .A1(n18374), .A2(n18447), .ZN(n18398) );
  INV_X1 U21513 ( .A(n18375), .ZN(n18419) );
  INV_X1 U21514 ( .A(n18447), .ZN(n18424) );
  AOI22_X1 U21515 ( .A1(n18530), .A2(n18419), .B1(n18525), .B2(n18392), .ZN(
        n18379) );
  INV_X1 U21516 ( .A(n18376), .ZN(n18526) );
  NOR2_X1 U21517 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18424), .ZN(
        n18426) );
  AOI22_X1 U21518 ( .A1(n18529), .A2(n18377), .B1(n18526), .B2(n18426), .ZN(
        n18394) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18524), .ZN(n18378) );
  OAI211_X1 U21520 ( .C1(n18533), .C2(n18398), .A(n18379), .B(n18378), .ZN(
        P3_U2940) );
  AOI22_X1 U21521 ( .A1(n18393), .A2(n18536), .B1(n18534), .B2(n18392), .ZN(
        n18381) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18394), .B1(
        n18535), .B2(n18419), .ZN(n18380) );
  OAI211_X1 U21523 ( .C1(n18539), .C2(n18398), .A(n18381), .B(n18380), .ZN(
        P3_U2941) );
  AOI22_X1 U21524 ( .A1(n18393), .A2(n18542), .B1(n18540), .B2(n18392), .ZN(
        n18383) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18394), .B1(
        n18541), .B2(n18419), .ZN(n18382) );
  OAI211_X1 U21526 ( .C1(n18545), .C2(n18398), .A(n18383), .B(n18382), .ZN(
        P3_U2942) );
  AOI22_X1 U21527 ( .A1(n18547), .A2(n18419), .B1(n18546), .B2(n18392), .ZN(
        n18385) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18548), .ZN(n18384) );
  OAI211_X1 U21529 ( .C1(n18551), .C2(n18398), .A(n18385), .B(n18384), .ZN(
        P3_U2943) );
  AOI22_X1 U21530 ( .A1(n18393), .A2(n18552), .B1(n18553), .B2(n18392), .ZN(
        n18387) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18394), .B1(
        n18554), .B2(n18419), .ZN(n18386) );
  OAI211_X1 U21532 ( .C1(n18557), .C2(n18398), .A(n18387), .B(n18386), .ZN(
        P3_U2944) );
  AOI22_X1 U21533 ( .A1(n18559), .A2(n18392), .B1(n18558), .B2(n18419), .ZN(
        n18389) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18560), .ZN(n18388) );
  OAI211_X1 U21535 ( .C1(n18563), .C2(n18398), .A(n18389), .B(n18388), .ZN(
        P3_U2945) );
  AOI22_X1 U21536 ( .A1(n18393), .A2(n18566), .B1(n18565), .B2(n18392), .ZN(
        n18391) );
  AOI22_X1 U21537 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18394), .B1(
        n18564), .B2(n18419), .ZN(n18390) );
  OAI211_X1 U21538 ( .C1(n18569), .C2(n18398), .A(n18391), .B(n18390), .ZN(
        P3_U2946) );
  AOI22_X1 U21539 ( .A1(n18573), .A2(n18392), .B1(n18571), .B2(n18419), .ZN(
        n18396) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18394), .B1(
        n18393), .B2(n18575), .ZN(n18395) );
  OAI211_X1 U21541 ( .C1(n18580), .C2(n18398), .A(n18396), .B(n18395), .ZN(
        P3_U2947) );
  NAND2_X1 U21542 ( .A1(n18397), .A2(n18447), .ZN(n18423) );
  AOI21_X1 U21543 ( .B1(n18398), .B2(n18423), .A(n18523), .ZN(n18418) );
  AOI22_X1 U21544 ( .A1(n18530), .A2(n18442), .B1(n18525), .B2(n18418), .ZN(
        n18405) );
  INV_X1 U21545 ( .A(n18423), .ZN(n18490) );
  INV_X1 U21546 ( .A(n18398), .ZN(n18468) );
  NOR2_X1 U21547 ( .A1(n18468), .A2(n18490), .ZN(n18402) );
  INV_X1 U21548 ( .A(n18399), .ZN(n18400) );
  OAI22_X1 U21549 ( .A1(n18402), .A2(n18497), .B1(n18401), .B2(n18400), .ZN(
        n18403) );
  OAI21_X1 U21550 ( .B1(n18490), .B2(n18758), .A(n18403), .ZN(n18420) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18420), .B1(
        n18524), .B2(n18419), .ZN(n18404) );
  OAI211_X1 U21552 ( .C1(n18533), .C2(n18423), .A(n18405), .B(n18404), .ZN(
        P3_U2948) );
  AOI22_X1 U21553 ( .A1(n18535), .A2(n18442), .B1(n18534), .B2(n18418), .ZN(
        n18407) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18420), .B1(
        n18536), .B2(n18419), .ZN(n18406) );
  OAI211_X1 U21555 ( .C1(n18539), .C2(n18423), .A(n18407), .B(n18406), .ZN(
        P3_U2949) );
  AOI22_X1 U21556 ( .A1(n18540), .A2(n18418), .B1(n18542), .B2(n18419), .ZN(
        n18409) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18420), .B1(
        n18541), .B2(n18442), .ZN(n18408) );
  OAI211_X1 U21558 ( .C1(n18545), .C2(n18423), .A(n18409), .B(n18408), .ZN(
        P3_U2950) );
  AOI22_X1 U21559 ( .A1(n18546), .A2(n18418), .B1(n18548), .B2(n18419), .ZN(
        n18411) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18420), .B1(
        n18547), .B2(n18442), .ZN(n18410) );
  OAI211_X1 U21561 ( .C1(n18551), .C2(n18423), .A(n18411), .B(n18410), .ZN(
        P3_U2951) );
  AOI22_X1 U21562 ( .A1(n18554), .A2(n18442), .B1(n18553), .B2(n18418), .ZN(
        n18413) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18420), .B1(
        n18552), .B2(n18419), .ZN(n18412) );
  OAI211_X1 U21564 ( .C1(n18557), .C2(n18423), .A(n18413), .B(n18412), .ZN(
        P3_U2952) );
  AOI22_X1 U21565 ( .A1(n18560), .A2(n18419), .B1(n18559), .B2(n18418), .ZN(
        n18415) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18420), .B1(
        n18558), .B2(n18442), .ZN(n18414) );
  OAI211_X1 U21567 ( .C1(n18563), .C2(n18423), .A(n18415), .B(n18414), .ZN(
        P3_U2953) );
  AOI22_X1 U21568 ( .A1(n18565), .A2(n18418), .B1(n18564), .B2(n18442), .ZN(
        n18417) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18420), .B1(
        n18566), .B2(n18419), .ZN(n18416) );
  OAI211_X1 U21570 ( .C1(n18569), .C2(n18423), .A(n18417), .B(n18416), .ZN(
        P3_U2954) );
  AOI22_X1 U21571 ( .A1(n18575), .A2(n18419), .B1(n18573), .B2(n18418), .ZN(
        n18422) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18420), .B1(
        n18571), .B2(n18442), .ZN(n18421) );
  OAI211_X1 U21573 ( .C1(n18580), .C2(n18423), .A(n18422), .B(n18421), .ZN(
        P3_U2955) );
  NOR2_X1 U21574 ( .A1(n18623), .A2(n18424), .ZN(n18474) );
  NAND2_X1 U21575 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18474), .ZN(
        n18446) );
  INV_X1 U21576 ( .A(n18474), .ZN(n18425) );
  NOR2_X1 U21577 ( .A1(n18523), .A2(n18425), .ZN(n18441) );
  AOI22_X1 U21578 ( .A1(n18530), .A2(n18468), .B1(n18525), .B2(n18441), .ZN(
        n18428) );
  AOI22_X1 U21579 ( .A1(n18529), .A2(n18426), .B1(n18526), .B2(n18474), .ZN(
        n18443) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18443), .B1(
        n18524), .B2(n18442), .ZN(n18427) );
  OAI211_X1 U21581 ( .C1(n18533), .C2(n18446), .A(n18428), .B(n18427), .ZN(
        P3_U2956) );
  AOI22_X1 U21582 ( .A1(n18536), .A2(n18442), .B1(n18534), .B2(n18441), .ZN(
        n18430) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18443), .B1(
        n18535), .B2(n18468), .ZN(n18429) );
  OAI211_X1 U21584 ( .C1(n18539), .C2(n18446), .A(n18430), .B(n18429), .ZN(
        P3_U2957) );
  AOI22_X1 U21585 ( .A1(n18540), .A2(n18441), .B1(n18542), .B2(n18442), .ZN(
        n18432) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18443), .B1(
        n18541), .B2(n18468), .ZN(n18431) );
  OAI211_X1 U21587 ( .C1(n18545), .C2(n18446), .A(n18432), .B(n18431), .ZN(
        P3_U2958) );
  AOI22_X1 U21588 ( .A1(n18547), .A2(n18468), .B1(n18546), .B2(n18441), .ZN(
        n18434) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18443), .B1(
        n18548), .B2(n18442), .ZN(n18433) );
  OAI211_X1 U21590 ( .C1(n18551), .C2(n18446), .A(n18434), .B(n18433), .ZN(
        P3_U2959) );
  AOI22_X1 U21591 ( .A1(n18553), .A2(n18441), .B1(n18552), .B2(n18442), .ZN(
        n18436) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18443), .B1(
        n18554), .B2(n18468), .ZN(n18435) );
  OAI211_X1 U21593 ( .C1(n18557), .C2(n18446), .A(n18436), .B(n18435), .ZN(
        P3_U2960) );
  AOI22_X1 U21594 ( .A1(n18560), .A2(n18442), .B1(n18559), .B2(n18441), .ZN(
        n18438) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18443), .B1(
        n18558), .B2(n18468), .ZN(n18437) );
  OAI211_X1 U21596 ( .C1(n18563), .C2(n18446), .A(n18438), .B(n18437), .ZN(
        P3_U2961) );
  AOI22_X1 U21597 ( .A1(n18566), .A2(n18442), .B1(n18565), .B2(n18441), .ZN(
        n18440) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18443), .B1(
        n18564), .B2(n18468), .ZN(n18439) );
  OAI211_X1 U21599 ( .C1(n18569), .C2(n18446), .A(n18440), .B(n18439), .ZN(
        P3_U2962) );
  AOI22_X1 U21600 ( .A1(n18575), .A2(n18442), .B1(n18573), .B2(n18441), .ZN(
        n18445) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18443), .B1(
        n18571), .B2(n18468), .ZN(n18444) );
  OAI211_X1 U21602 ( .C1(n18580), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2963) );
  NAND2_X1 U21603 ( .A1(n18528), .A2(n18621), .ZN(n18472) );
  INV_X1 U21604 ( .A(n18472), .ZN(n18574) );
  NOR2_X1 U21605 ( .A1(n18517), .A2(n18574), .ZN(n18499) );
  NOR2_X1 U21606 ( .A1(n18523), .A2(n18499), .ZN(n18467) );
  AOI22_X1 U21607 ( .A1(n18525), .A2(n18467), .B1(n18524), .B2(n18468), .ZN(
        n18454) );
  NAND2_X1 U21608 ( .A1(n18448), .A2(n18447), .ZN(n18449) );
  OAI21_X1 U21609 ( .B1(n18450), .B2(n18449), .A(n18499), .ZN(n18451) );
  OAI211_X1 U21610 ( .C1(n18574), .C2(n18758), .A(n18452), .B(n18451), .ZN(
        n18469) );
  AOI22_X1 U21611 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18469), .B1(
        n18530), .B2(n18490), .ZN(n18453) );
  OAI211_X1 U21612 ( .C1(n18533), .C2(n18472), .A(n18454), .B(n18453), .ZN(
        P3_U2964) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18469), .B1(
        n18534), .B2(n18467), .ZN(n18456) );
  AOI22_X1 U21614 ( .A1(n18536), .A2(n18468), .B1(n18535), .B2(n18490), .ZN(
        n18455) );
  OAI211_X1 U21615 ( .C1(n18539), .C2(n18472), .A(n18456), .B(n18455), .ZN(
        P3_U2965) );
  AOI22_X1 U21616 ( .A1(n18541), .A2(n18490), .B1(n18540), .B2(n18467), .ZN(
        n18458) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18469), .B1(
        n18542), .B2(n18468), .ZN(n18457) );
  OAI211_X1 U21618 ( .C1(n18545), .C2(n18472), .A(n18458), .B(n18457), .ZN(
        P3_U2966) );
  AOI22_X1 U21619 ( .A1(n18546), .A2(n18467), .B1(n18548), .B2(n18468), .ZN(
        n18460) );
  AOI22_X1 U21620 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18469), .B1(
        n18547), .B2(n18490), .ZN(n18459) );
  OAI211_X1 U21621 ( .C1(n18551), .C2(n18472), .A(n18460), .B(n18459), .ZN(
        P3_U2967) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18469), .B1(
        n18553), .B2(n18467), .ZN(n18462) );
  AOI22_X1 U21623 ( .A1(n18554), .A2(n18490), .B1(n18552), .B2(n18468), .ZN(
        n18461) );
  OAI211_X1 U21624 ( .C1(n18557), .C2(n18472), .A(n18462), .B(n18461), .ZN(
        P3_U2968) );
  AOI22_X1 U21625 ( .A1(n18560), .A2(n18468), .B1(n18559), .B2(n18467), .ZN(
        n18464) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18469), .B1(
        n18558), .B2(n18490), .ZN(n18463) );
  OAI211_X1 U21627 ( .C1(n18563), .C2(n18472), .A(n18464), .B(n18463), .ZN(
        P3_U2969) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18469), .B1(
        n18565), .B2(n18467), .ZN(n18466) );
  AOI22_X1 U21629 ( .A1(n18566), .A2(n18468), .B1(n18564), .B2(n18490), .ZN(
        n18465) );
  OAI211_X1 U21630 ( .C1(n18569), .C2(n18472), .A(n18466), .B(n18465), .ZN(
        P3_U2970) );
  AOI22_X1 U21631 ( .A1(n18575), .A2(n18468), .B1(n18573), .B2(n18467), .ZN(
        n18471) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18469), .B1(
        n18571), .B2(n18490), .ZN(n18470) );
  OAI211_X1 U21633 ( .C1(n18580), .C2(n18472), .A(n18471), .B(n18470), .ZN(
        P3_U2971) );
  INV_X1 U21634 ( .A(n18570), .ZN(n18494) );
  NOR2_X1 U21635 ( .A1(n18523), .A2(n18473), .ZN(n18489) );
  AOI22_X1 U21636 ( .A1(n18525), .A2(n18489), .B1(n18524), .B2(n18490), .ZN(
        n18476) );
  AOI22_X1 U21637 ( .A1(n18529), .A2(n18474), .B1(n18528), .B2(n18526), .ZN(
        n18491) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18491), .B1(
        n18530), .B2(n18517), .ZN(n18475) );
  OAI211_X1 U21639 ( .C1(n18533), .C2(n18494), .A(n18476), .B(n18475), .ZN(
        P3_U2972) );
  AOI22_X1 U21640 ( .A1(n18536), .A2(n18490), .B1(n18534), .B2(n18489), .ZN(
        n18478) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18491), .B1(
        n18535), .B2(n18517), .ZN(n18477) );
  OAI211_X1 U21642 ( .C1(n18539), .C2(n18494), .A(n18478), .B(n18477), .ZN(
        P3_U2973) );
  AOI22_X1 U21643 ( .A1(n18541), .A2(n18517), .B1(n18540), .B2(n18489), .ZN(
        n18480) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18491), .B1(
        n18542), .B2(n18490), .ZN(n18479) );
  OAI211_X1 U21645 ( .C1(n18545), .C2(n18494), .A(n18480), .B(n18479), .ZN(
        P3_U2974) );
  AOI22_X1 U21646 ( .A1(n18546), .A2(n18489), .B1(n18548), .B2(n18490), .ZN(
        n18482) );
  AOI22_X1 U21647 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18491), .B1(
        n18547), .B2(n18517), .ZN(n18481) );
  OAI211_X1 U21648 ( .C1(n18551), .C2(n18494), .A(n18482), .B(n18481), .ZN(
        P3_U2975) );
  AOI22_X1 U21649 ( .A1(n18554), .A2(n18517), .B1(n18553), .B2(n18489), .ZN(
        n18484) );
  AOI22_X1 U21650 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18491), .B1(
        n18552), .B2(n18490), .ZN(n18483) );
  OAI211_X1 U21651 ( .C1(n18557), .C2(n18494), .A(n18484), .B(n18483), .ZN(
        P3_U2976) );
  AOI22_X1 U21652 ( .A1(n18560), .A2(n18490), .B1(n18559), .B2(n18489), .ZN(
        n18486) );
  AOI22_X1 U21653 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18491), .B1(
        n18558), .B2(n18517), .ZN(n18485) );
  OAI211_X1 U21654 ( .C1(n18563), .C2(n18494), .A(n18486), .B(n18485), .ZN(
        P3_U2977) );
  AOI22_X1 U21655 ( .A1(n18566), .A2(n18490), .B1(n18565), .B2(n18489), .ZN(
        n18488) );
  AOI22_X1 U21656 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18491), .B1(
        n18564), .B2(n18517), .ZN(n18487) );
  OAI211_X1 U21657 ( .C1(n18569), .C2(n18494), .A(n18488), .B(n18487), .ZN(
        P3_U2978) );
  AOI22_X1 U21658 ( .A1(n18575), .A2(n18490), .B1(n18573), .B2(n18489), .ZN(
        n18493) );
  AOI22_X1 U21659 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18491), .B1(
        n18571), .B2(n18517), .ZN(n18492) );
  OAI211_X1 U21660 ( .C1(n18580), .C2(n18494), .A(n18493), .B(n18492), .ZN(
        P3_U2979) );
  INV_X1 U21661 ( .A(n18501), .ZN(n18521) );
  INV_X1 U21662 ( .A(n18495), .ZN(n18496) );
  NOR2_X1 U21663 ( .A1(n18523), .A2(n18496), .ZN(n18516) );
  AOI22_X1 U21664 ( .A1(n18525), .A2(n18516), .B1(n18524), .B2(n18517), .ZN(
        n18503) );
  OAI22_X1 U21665 ( .A1(n18499), .A2(n18498), .B1(n18497), .B2(n18496), .ZN(
        n18500) );
  OAI21_X1 U21666 ( .B1(n18501), .B2(n18758), .A(n18500), .ZN(n18518) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18518), .B1(
        n18530), .B2(n18574), .ZN(n18502) );
  OAI211_X1 U21668 ( .C1(n18533), .C2(n18521), .A(n18503), .B(n18502), .ZN(
        P3_U2980) );
  AOI22_X1 U21669 ( .A1(n18535), .A2(n18574), .B1(n18534), .B2(n18516), .ZN(
        n18505) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18518), .B1(
        n18536), .B2(n18517), .ZN(n18504) );
  OAI211_X1 U21671 ( .C1(n18539), .C2(n18521), .A(n18505), .B(n18504), .ZN(
        P3_U2981) );
  AOI22_X1 U21672 ( .A1(n18540), .A2(n18516), .B1(n18542), .B2(n18517), .ZN(
        n18507) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18518), .B1(
        n18541), .B2(n18574), .ZN(n18506) );
  OAI211_X1 U21674 ( .C1(n18545), .C2(n18521), .A(n18507), .B(n18506), .ZN(
        P3_U2982) );
  AOI22_X1 U21675 ( .A1(n18547), .A2(n18574), .B1(n18546), .B2(n18516), .ZN(
        n18509) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18518), .B1(
        n18548), .B2(n18517), .ZN(n18508) );
  OAI211_X1 U21677 ( .C1(n18551), .C2(n18521), .A(n18509), .B(n18508), .ZN(
        P3_U2983) );
  AOI22_X1 U21678 ( .A1(n18553), .A2(n18516), .B1(n18552), .B2(n18517), .ZN(
        n18511) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18518), .B1(
        n18554), .B2(n18574), .ZN(n18510) );
  OAI211_X1 U21680 ( .C1(n18557), .C2(n18521), .A(n18511), .B(n18510), .ZN(
        P3_U2984) );
  AOI22_X1 U21681 ( .A1(n18559), .A2(n18516), .B1(n18558), .B2(n18574), .ZN(
        n18513) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18518), .B1(
        n18560), .B2(n18517), .ZN(n18512) );
  OAI211_X1 U21683 ( .C1(n18563), .C2(n18521), .A(n18513), .B(n18512), .ZN(
        P3_U2985) );
  AOI22_X1 U21684 ( .A1(n18565), .A2(n18516), .B1(n18564), .B2(n18574), .ZN(
        n18515) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18518), .B1(
        n18566), .B2(n18517), .ZN(n18514) );
  OAI211_X1 U21686 ( .C1(n18569), .C2(n18521), .A(n18515), .B(n18514), .ZN(
        P3_U2986) );
  AOI22_X1 U21687 ( .A1(n18573), .A2(n18516), .B1(n18571), .B2(n18574), .ZN(
        n18520) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18518), .B1(
        n18575), .B2(n18517), .ZN(n18519) );
  OAI211_X1 U21689 ( .C1(n18580), .C2(n18521), .A(n18520), .B(n18519), .ZN(
        P3_U2987) );
  INV_X1 U21690 ( .A(n18527), .ZN(n18522) );
  NOR2_X1 U21691 ( .A1(n18523), .A2(n18522), .ZN(n18572) );
  AOI22_X1 U21692 ( .A1(n18525), .A2(n18572), .B1(n18524), .B2(n18574), .ZN(
        n18532) );
  AOI22_X1 U21693 ( .A1(n18529), .A2(n18528), .B1(n18527), .B2(n18526), .ZN(
        n18576) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18576), .B1(
        n18530), .B2(n18570), .ZN(n18531) );
  OAI211_X1 U21695 ( .C1(n18533), .C2(n18579), .A(n18532), .B(n18531), .ZN(
        P3_U2988) );
  AOI22_X1 U21696 ( .A1(n18535), .A2(n18570), .B1(n18534), .B2(n18572), .ZN(
        n18538) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18576), .B1(
        n18536), .B2(n18574), .ZN(n18537) );
  OAI211_X1 U21698 ( .C1(n18539), .C2(n18579), .A(n18538), .B(n18537), .ZN(
        P3_U2989) );
  AOI22_X1 U21699 ( .A1(n18541), .A2(n18570), .B1(n18540), .B2(n18572), .ZN(
        n18544) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18576), .B1(
        n18542), .B2(n18574), .ZN(n18543) );
  OAI211_X1 U21701 ( .C1(n18545), .C2(n18579), .A(n18544), .B(n18543), .ZN(
        P3_U2990) );
  AOI22_X1 U21702 ( .A1(n18547), .A2(n18570), .B1(n18546), .B2(n18572), .ZN(
        n18550) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18576), .B1(
        n18548), .B2(n18574), .ZN(n18549) );
  OAI211_X1 U21704 ( .C1(n18551), .C2(n18579), .A(n18550), .B(n18549), .ZN(
        P3_U2991) );
  AOI22_X1 U21705 ( .A1(n18553), .A2(n18572), .B1(n18552), .B2(n18574), .ZN(
        n18556) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18576), .B1(
        n18554), .B2(n18570), .ZN(n18555) );
  OAI211_X1 U21707 ( .C1(n18557), .C2(n18579), .A(n18556), .B(n18555), .ZN(
        P3_U2992) );
  AOI22_X1 U21708 ( .A1(n18559), .A2(n18572), .B1(n18558), .B2(n18570), .ZN(
        n18562) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18576), .B1(
        n18560), .B2(n18574), .ZN(n18561) );
  OAI211_X1 U21710 ( .C1(n18563), .C2(n18579), .A(n18562), .B(n18561), .ZN(
        P3_U2993) );
  AOI22_X1 U21711 ( .A1(n18565), .A2(n18572), .B1(n18564), .B2(n18570), .ZN(
        n18568) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18576), .B1(
        n18566), .B2(n18574), .ZN(n18567) );
  OAI211_X1 U21713 ( .C1(n18569), .C2(n18579), .A(n18568), .B(n18567), .ZN(
        P3_U2994) );
  AOI22_X1 U21714 ( .A1(n18573), .A2(n18572), .B1(n18571), .B2(n18570), .ZN(
        n18578) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18576), .B1(
        n18575), .B2(n18574), .ZN(n18577) );
  OAI211_X1 U21716 ( .C1(n18580), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2995) );
  NOR2_X1 U21717 ( .A1(n18613), .A2(n18581), .ZN(n18584) );
  INV_X1 U21718 ( .A(n18582), .ZN(n18583) );
  OAI222_X1 U21719 ( .A1(n18588), .A2(n18587), .B1(n18586), .B2(n18585), .C1(
        n18584), .C2(n18583), .ZN(n18802) );
  OAI21_X1 U21720 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18589), .ZN(n18590) );
  OAI211_X1 U21721 ( .C1(n18614), .C2(n18639), .A(n18591), .B(n18590), .ZN(
        n18637) );
  NAND2_X1 U21722 ( .A1(n18617), .A2(n18789), .ZN(n18618) );
  AOI22_X1 U21723 ( .A1(n18613), .A2(n18595), .B1(n18602), .B2(n18618), .ZN(
        n18759) );
  NOR2_X1 U21724 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18759), .ZN(
        n18599) );
  OAI21_X1 U21725 ( .B1(n18594), .B2(n18593), .A(n18592), .ZN(n18600) );
  OAI21_X1 U21726 ( .B1(n18617), .B2(n18602), .A(n18595), .ZN(n18596) );
  AOI21_X1 U21727 ( .B1(n18597), .B2(n18600), .A(n18596), .ZN(n18762) );
  NAND2_X1 U21728 ( .A1(n18614), .A2(n18762), .ZN(n18598) );
  AOI22_X1 U21729 ( .A1(n18614), .A2(n18599), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18598), .ZN(n18635) );
  AOI21_X1 U21730 ( .B1(n18782), .B2(n18606), .A(n18600), .ZN(n18611) );
  NAND2_X1 U21731 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18601), .ZN(
        n18610) );
  INV_X1 U21732 ( .A(n18602), .ZN(n18603) );
  OAI211_X1 U21733 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18604), .B(n18603), .ZN(
        n18609) );
  NOR2_X1 U21734 ( .A1(n18605), .A2(n18789), .ZN(n18607) );
  OAI211_X1 U21735 ( .C1(n18607), .C2(n18606), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n11412), .ZN(n18608) );
  OAI211_X1 U21736 ( .C1(n18611), .C2(n18610), .A(n18609), .B(n18608), .ZN(
        n18612) );
  AOI21_X1 U21737 ( .B1(n18613), .B2(n18769), .A(n18612), .ZN(n18772) );
  AOI22_X1 U21738 ( .A1(n18626), .A2(n11412), .B1(n18772), .B2(n18614), .ZN(
        n18630) );
  NOR2_X1 U21739 ( .A1(n18616), .A2(n18615), .ZN(n18620) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18617), .B1(
        n18620), .B2(n18789), .ZN(n18784) );
  INV_X1 U21741 ( .A(n18618), .ZN(n18619) );
  OAI22_X1 U21742 ( .A1(n18620), .A2(n18775), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18619), .ZN(n18780) );
  OR3_X1 U21743 ( .A1(n18784), .A2(n18623), .A3(n18621), .ZN(n18622) );
  AOI22_X1 U21744 ( .A1(n18784), .A2(n18623), .B1(n18780), .B2(n18622), .ZN(
        n18625) );
  OAI21_X1 U21745 ( .B1(n18626), .B2(n18625), .A(n18624), .ZN(n18629) );
  AND2_X1 U21746 ( .A1(n18630), .A2(n18629), .ZN(n18627) );
  OAI221_X1 U21747 ( .B1(n18630), .B2(n18629), .C1(n18628), .C2(n18627), .A(
        n18632), .ZN(n18634) );
  AOI21_X1 U21748 ( .B1(n18632), .B2(n18631), .A(n18630), .ZN(n18633) );
  AOI222_X1 U21749 ( .A1(n18635), .A2(n18634), .B1(n18635), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18634), .C2(n18633), .ZN(
        n18636) );
  NOR4_X1 U21750 ( .A1(n18638), .A2(n18802), .A3(n18637), .A4(n18636), .ZN(
        n18650) );
  INV_X1 U21751 ( .A(n18645), .ZN(n18640) );
  AOI22_X1 U21752 ( .A1(n18641), .A2(n18669), .B1(n18640), .B2(n18639), .ZN(
        n18647) );
  OAI211_X1 U21753 ( .C1(n18644), .C2(n18643), .A(n18642), .B(n18650), .ZN(
        n18757) );
  NAND2_X1 U21754 ( .A1(n18669), .A2(n18812), .ZN(n18651) );
  NAND4_X1 U21755 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18757), .A3(n18645), 
        .A4(n18651), .ZN(n18655) );
  OAI22_X1 U21756 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18647), .B1(n18646), 
        .B2(n18655), .ZN(n18648) );
  OAI21_X1 U21757 ( .B1(n18650), .B2(n18649), .A(n18648), .ZN(P3_U2996) );
  NOR3_X1 U21758 ( .A1(n18813), .A2(n18652), .A3(n18651), .ZN(n18657) );
  AOI211_X1 U21759 ( .C1(n18669), .C2(n18805), .A(n18653), .B(n18657), .ZN(
        n18654) );
  OAI21_X1 U21760 ( .B1(P3_STATE2_REG_1__SCAN_IN), .B2(n18655), .A(n18654), 
        .ZN(P3_U2997) );
  OAI21_X1 U21761 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18656), .ZN(n18658) );
  AOI21_X1 U21762 ( .B1(n18659), .B2(n18658), .A(n18657), .ZN(P3_U2998) );
  AND2_X1 U21763 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18752), .ZN(
        P3_U2999) );
  AND2_X1 U21764 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18660), .ZN(
        P3_U3000) );
  AND2_X1 U21765 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18660), .ZN(
        P3_U3001) );
  AND2_X1 U21766 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18752), .ZN(
        P3_U3002) );
  AND2_X1 U21767 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18752), .ZN(
        P3_U3003) );
  AND2_X1 U21768 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18752), .ZN(
        P3_U3004) );
  AND2_X1 U21769 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18752), .ZN(
        P3_U3005) );
  AND2_X1 U21770 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18752), .ZN(
        P3_U3006) );
  AND2_X1 U21771 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18660), .ZN(
        P3_U3007) );
  AND2_X1 U21772 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18660), .ZN(
        P3_U3008) );
  AND2_X1 U21773 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18660), .ZN(
        P3_U3009) );
  AND2_X1 U21774 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18660), .ZN(
        P3_U3010) );
  AND2_X1 U21775 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18660), .ZN(
        P3_U3011) );
  AND2_X1 U21776 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18660), .ZN(
        P3_U3012) );
  AND2_X1 U21777 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18660), .ZN(
        P3_U3013) );
  AND2_X1 U21778 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18660), .ZN(
        P3_U3014) );
  AND2_X1 U21779 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18660), .ZN(
        P3_U3015) );
  AND2_X1 U21780 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18660), .ZN(
        P3_U3016) );
  AND2_X1 U21781 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18752), .ZN(
        P3_U3017) );
  AND2_X1 U21782 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18752), .ZN(
        P3_U3018) );
  AND2_X1 U21783 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18752), .ZN(
        P3_U3019) );
  AND2_X1 U21784 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18752), .ZN(
        P3_U3020) );
  AND2_X1 U21785 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18660), .ZN(P3_U3021) );
  AND2_X1 U21786 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18752), .ZN(P3_U3022) );
  AND2_X1 U21787 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18752), .ZN(P3_U3023) );
  AND2_X1 U21788 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18752), .ZN(P3_U3024) );
  AND2_X1 U21789 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18752), .ZN(P3_U3025) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18752), .ZN(P3_U3026) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18752), .ZN(P3_U3027) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18752), .ZN(P3_U3028) );
  INV_X1 U21793 ( .A(n18661), .ZN(n18662) );
  OAI21_X1 U21794 ( .B1(n18662), .B2(n20724), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18663) );
  AOI22_X1 U21795 ( .A1(n18677), .A2(n18679), .B1(n18799), .B2(n18663), .ZN(
        n18665) );
  NAND3_X1 U21796 ( .A1(NA), .A2(n18677), .A3(n18671), .ZN(n18664) );
  OAI211_X1 U21797 ( .C1(n18666), .C2(n18809), .A(n18665), .B(n18664), .ZN(
        P3_U3029) );
  AOI21_X1 U21798 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18667) );
  AOI21_X1 U21799 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18667), .ZN(
        n18668) );
  AOI22_X1 U21800 ( .A1(n18669), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18668), .ZN(n18670) );
  NAND2_X1 U21801 ( .A1(n18670), .A2(n18806), .ZN(P3_U3030) );
  INV_X1 U21802 ( .A(NA), .ZN(n21174) );
  NOR2_X1 U21803 ( .A1(n18809), .A2(n18671), .ZN(n18672) );
  AOI221_X1 U21804 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(n18677), .C1(n21174), 
        .C2(n18677), .A(n18672), .ZN(n18678) );
  NOR2_X1 U21805 ( .A1(n18679), .A2(n20724), .ZN(n18675) );
  INV_X1 U21806 ( .A(n18672), .ZN(n18673) );
  OAI22_X1 U21807 ( .A1(NA), .A2(n18673), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18674) );
  OAI22_X1 U21808 ( .A1(n18675), .A2(n18674), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18676) );
  OAI22_X1 U21809 ( .A1(n18678), .A2(n18679), .B1(n18677), .B2(n18676), .ZN(
        P3_U3031) );
  NAND2_X1 U21810 ( .A1(n18733), .A2(n18679), .ZN(n18738) );
  CLKBUF_X1 U21811 ( .A(n18738), .Z(n18739) );
  OAI222_X1 U21812 ( .A1(n18791), .A2(n18743), .B1(n18680), .B2(n18733), .C1(
        n18681), .C2(n18739), .ZN(P3_U3032) );
  OAI222_X1 U21813 ( .A1(n18738), .A2(n18683), .B1(n18682), .B2(n18733), .C1(
        n18681), .C2(n18743), .ZN(P3_U3033) );
  OAI222_X1 U21814 ( .A1(n18738), .A2(n18685), .B1(n18684), .B2(n18733), .C1(
        n18683), .C2(n18743), .ZN(P3_U3034) );
  OAI222_X1 U21815 ( .A1(n18738), .A2(n18688), .B1(n18686), .B2(n18733), .C1(
        n18685), .C2(n18743), .ZN(P3_U3035) );
  OAI222_X1 U21816 ( .A1(n18688), .A2(n18743), .B1(n18687), .B2(n18733), .C1(
        n18689), .C2(n18739), .ZN(P3_U3036) );
  OAI222_X1 U21817 ( .A1(n18738), .A2(n18691), .B1(n18690), .B2(n18733), .C1(
        n18689), .C2(n18743), .ZN(P3_U3037) );
  INV_X1 U21818 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18694) );
  OAI222_X1 U21819 ( .A1(n18738), .A2(n18694), .B1(n18692), .B2(n18733), .C1(
        n18691), .C2(n18743), .ZN(P3_U3038) );
  OAI222_X1 U21820 ( .A1(n18694), .A2(n18743), .B1(n18693), .B2(n18733), .C1(
        n18695), .C2(n18739), .ZN(P3_U3039) );
  OAI222_X1 U21821 ( .A1(n18738), .A2(n18697), .B1(n18696), .B2(n18733), .C1(
        n18695), .C2(n18743), .ZN(P3_U3040) );
  OAI222_X1 U21822 ( .A1(n18739), .A2(n18699), .B1(n18698), .B2(n18733), .C1(
        n18697), .C2(n18743), .ZN(P3_U3041) );
  OAI222_X1 U21823 ( .A1(n18739), .A2(n18701), .B1(n18700), .B2(n18733), .C1(
        n18699), .C2(n18743), .ZN(P3_U3042) );
  INV_X1 U21824 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18703) );
  OAI222_X1 U21825 ( .A1(n18739), .A2(n18703), .B1(n18702), .B2(n18733), .C1(
        n18701), .C2(n18743), .ZN(P3_U3043) );
  OAI222_X1 U21826 ( .A1(n18739), .A2(n18705), .B1(n18704), .B2(n18733), .C1(
        n18703), .C2(n18743), .ZN(P3_U3044) );
  OAI222_X1 U21827 ( .A1(n18739), .A2(n18708), .B1(n18706), .B2(n18733), .C1(
        n18705), .C2(n18743), .ZN(P3_U3045) );
  OAI222_X1 U21828 ( .A1(n18708), .A2(n18743), .B1(n18707), .B2(n18733), .C1(
        n18709), .C2(n18739), .ZN(P3_U3046) );
  OAI222_X1 U21829 ( .A1(n18739), .A2(n18712), .B1(n18710), .B2(n18733), .C1(
        n18709), .C2(n18743), .ZN(P3_U3047) );
  OAI222_X1 U21830 ( .A1(n18712), .A2(n18743), .B1(n18711), .B2(n18733), .C1(
        n18713), .C2(n18739), .ZN(P3_U3048) );
  INV_X1 U21831 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18716) );
  OAI222_X1 U21832 ( .A1(n18738), .A2(n18716), .B1(n18714), .B2(n18733), .C1(
        n18713), .C2(n18743), .ZN(P3_U3049) );
  OAI222_X1 U21833 ( .A1(n18716), .A2(n18743), .B1(n18715), .B2(n18733), .C1(
        n18717), .C2(n18739), .ZN(P3_U3050) );
  OAI222_X1 U21834 ( .A1(n18738), .A2(n18720), .B1(n18718), .B2(n18733), .C1(
        n18717), .C2(n18743), .ZN(P3_U3051) );
  OAI222_X1 U21835 ( .A1(n18720), .A2(n18743), .B1(n18719), .B2(n18733), .C1(
        n18721), .C2(n18739), .ZN(P3_U3052) );
  OAI222_X1 U21836 ( .A1(n18738), .A2(n18724), .B1(n18722), .B2(n18733), .C1(
        n18721), .C2(n18743), .ZN(P3_U3053) );
  OAI222_X1 U21837 ( .A1(n18724), .A2(n18743), .B1(n18723), .B2(n18733), .C1(
        n18725), .C2(n18739), .ZN(P3_U3054) );
  OAI222_X1 U21838 ( .A1(n18738), .A2(n18727), .B1(n18726), .B2(n18733), .C1(
        n18725), .C2(n18743), .ZN(P3_U3055) );
  INV_X1 U21839 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18729) );
  OAI222_X1 U21840 ( .A1(n18738), .A2(n18729), .B1(n18728), .B2(n18733), .C1(
        n18727), .C2(n18743), .ZN(P3_U3056) );
  OAI222_X1 U21841 ( .A1(n18739), .A2(n18731), .B1(n18730), .B2(n18733), .C1(
        n18729), .C2(n18743), .ZN(P3_U3057) );
  INV_X1 U21842 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18735) );
  OAI222_X1 U21843 ( .A1(n18739), .A2(n18735), .B1(n18732), .B2(n18733), .C1(
        n18731), .C2(n18743), .ZN(P3_U3058) );
  OAI222_X1 U21844 ( .A1(n18735), .A2(n18743), .B1(n18734), .B2(n18733), .C1(
        n18736), .C2(n18739), .ZN(P3_U3059) );
  OAI222_X1 U21845 ( .A1(n18738), .A2(n18742), .B1(n18737), .B2(n18733), .C1(
        n18736), .C2(n18743), .ZN(P3_U3060) );
  INV_X1 U21846 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18741) );
  OAI222_X1 U21847 ( .A1(n18743), .A2(n18742), .B1(n18741), .B2(n18733), .C1(
        n18740), .C2(n18739), .ZN(P3_U3061) );
  INV_X1 U21848 ( .A(P3_BE_N_REG_3__SCAN_IN), .ZN(n18744) );
  AOI22_X1 U21849 ( .A1(n18733), .A2(n18745), .B1(n18744), .B2(n18799), .ZN(
        P3_U3274) );
  INV_X1 U21850 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18794) );
  INV_X1 U21851 ( .A(P3_BE_N_REG_2__SCAN_IN), .ZN(n18746) );
  AOI22_X1 U21852 ( .A1(n18733), .A2(n18794), .B1(n18746), .B2(n18799), .ZN(
        P3_U3275) );
  INV_X1 U21853 ( .A(P3_BE_N_REG_1__SCAN_IN), .ZN(n18747) );
  AOI22_X1 U21854 ( .A1(n18733), .A2(n18748), .B1(n18747), .B2(n18799), .ZN(
        P3_U3276) );
  INV_X1 U21855 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18797) );
  INV_X1 U21856 ( .A(P3_BE_N_REG_0__SCAN_IN), .ZN(n18749) );
  AOI22_X1 U21857 ( .A1(n18733), .A2(n18797), .B1(n18749), .B2(n18799), .ZN(
        P3_U3277) );
  INV_X1 U21858 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18751) );
  AOI21_X1 U21859 ( .B1(n18752), .B2(n18751), .A(n18750), .ZN(P3_U3280) );
  OAI21_X1 U21860 ( .B1(n18755), .B2(n18754), .A(n18753), .ZN(P3_U3281) );
  OAI221_X1 U21861 ( .B1(n18758), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18758), 
        .C2(n18757), .A(n18756), .ZN(P3_U3282) );
  NOR3_X1 U21862 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18759), .A3(
        n18771), .ZN(n18760) );
  AOI21_X1 U21863 ( .B1(n18783), .B2(n18761), .A(n18760), .ZN(n18766) );
  INV_X1 U21864 ( .A(n18771), .ZN(n18785) );
  INV_X1 U21865 ( .A(n18762), .ZN(n18763) );
  AOI21_X1 U21866 ( .B1(n18785), .B2(n18763), .A(n18790), .ZN(n18765) );
  OAI22_X1 U21867 ( .A1(n18790), .A2(n18766), .B1(n18765), .B2(n18764), .ZN(
        P3_U3285) );
  AOI22_X1 U21868 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n18768), .B2(n18767), .ZN(
        n18776) );
  NOR2_X1 U21869 ( .A1(n18813), .A2(n18786), .ZN(n18777) );
  INV_X1 U21870 ( .A(n18783), .ZN(n18770) );
  OAI22_X1 U21871 ( .A1(n18772), .A2(n18771), .B1(n18770), .B2(n18769), .ZN(
        n18773) );
  AOI21_X1 U21872 ( .B1(n18776), .B2(n18777), .A(n18773), .ZN(n18774) );
  AOI22_X1 U21873 ( .A1(n18790), .A2(n11412), .B1(n18774), .B2(n18787), .ZN(
        P3_U3288) );
  INV_X1 U21874 ( .A(n18775), .ZN(n18779) );
  INV_X1 U21875 ( .A(n18776), .ZN(n18778) );
  AOI222_X1 U21876 ( .A1(n18780), .A2(n18785), .B1(n18783), .B2(n18779), .C1(
        n18778), .C2(n18777), .ZN(n18781) );
  AOI22_X1 U21877 ( .A1(n18790), .A2(n18782), .B1(n18781), .B2(n18787), .ZN(
        P3_U3289) );
  AOI222_X1 U21878 ( .A1(n18786), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18785), 
        .B2(n18784), .C1(n18789), .C2(n18783), .ZN(n18788) );
  AOI22_X1 U21879 ( .A1(n18790), .A2(n18789), .B1(n18788), .B2(n18787), .ZN(
        P3_U3290) );
  AOI21_X1 U21880 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18792) );
  AOI22_X1 U21881 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18792), .B2(n18791), .ZN(n18795) );
  AOI22_X1 U21882 ( .A1(n18798), .A2(n18795), .B1(n18794), .B2(n18793), .ZN(
        P3_U3292) );
  OAI21_X1 U21883 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18798), .ZN(n18796) );
  OAI21_X1 U21884 ( .B1(n18798), .B2(n18797), .A(n18796), .ZN(P3_U3293) );
  INV_X1 U21885 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18800) );
  AOI22_X1 U21886 ( .A1(n18733), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18800), 
        .B2(n18799), .ZN(P3_U3294) );
  MUX2_X1 U21887 ( .A(P3_MORE_REG_SCAN_IN), .B(n18802), .S(n18801), .Z(
        P3_U3295) );
  AOI21_X1 U21888 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_0__SCAN_IN), .A(n18803), .ZN(n18804) );
  AOI211_X1 U21889 ( .C1(n18805), .C2(n18809), .A(n18804), .B(n18824), .ZN(
        n18817) );
  AOI21_X1 U21890 ( .B1(n18808), .B2(n18807), .A(n18806), .ZN(n18811) );
  OAI211_X1 U21891 ( .C1(n18811), .C2(n18810), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18809), .ZN(n18814) );
  AOI22_X1 U21892 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18814), .B1(n18813), 
        .B2(n18812), .ZN(n18816) );
  NAND2_X1 U21893 ( .A1(n18817), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18815) );
  OAI21_X1 U21894 ( .B1(n18817), .B2(n18816), .A(n18815), .ZN(P3_U3296) );
  MUX2_X1 U21895 ( .A(P3_M_IO_N_REG_SCAN_IN), .B(P3_MEMORYFETCH_REG_SCAN_IN), 
        .S(n18733), .Z(P3_U3297) );
  OAI21_X1 U21896 ( .B1(P3_READREQUEST_REG_SCAN_IN), .B2(n18821), .A(n18819), 
        .ZN(n18818) );
  OAI21_X1 U21897 ( .B1(n18820), .B2(n18819), .A(n18818), .ZN(P3_U3298) );
  NOR2_X1 U21898 ( .A1(n18821), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18823)
         );
  OAI21_X1 U21899 ( .B1(n18824), .B2(n18823), .A(n18822), .ZN(P3_U3299) );
  INV_X1 U21900 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19839) );
  INV_X1 U21901 ( .A(P2_ADS_N_REG_SCAN_IN), .ZN(n18825) );
  INV_X1 U21902 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19855) );
  NAND2_X1 U21903 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19855), .ZN(n19845) );
  AOI22_X1 U21904 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19845), .B1(
        P2_STATE_REG_1__SCAN_IN), .B2(n19839), .ZN(n19911) );
  OAI21_X1 U21905 ( .B1(n19839), .B2(n18825), .A(n19837), .ZN(P2_U2815) );
  AOI22_X1 U21906 ( .A1(n19974), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(
        P2_STATE2_REG_0__SCAN_IN), .B2(n18826), .ZN(n18827) );
  INV_X1 U21907 ( .A(n18827), .ZN(P2_U2816) );
  NAND2_X1 U21908 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19839), .ZN(n19990) );
  AOI21_X1 U21909 ( .B1(n19839), .B2(n19855), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18828) );
  AOI22_X1 U21910 ( .A1(n19892), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18828), 
        .B2(n19990), .ZN(P2_U2817) );
  OAI21_X1 U21911 ( .B1(n19847), .B2(BS16), .A(n19911), .ZN(n19909) );
  OAI21_X1 U21912 ( .B1(n19911), .B2(n19920), .A(n19909), .ZN(P2_U2818) );
  NOR4_X1 U21913 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18832) );
  NOR4_X1 U21914 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18831) );
  NOR4_X1 U21915 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18830) );
  NOR4_X1 U21916 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18829) );
  NAND4_X1 U21917 ( .A1(n18832), .A2(n18831), .A3(n18830), .A4(n18829), .ZN(
        n18838) );
  NOR4_X1 U21918 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18836) );
  AOI211_X1 U21919 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18835) );
  NOR4_X1 U21920 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18834) );
  NOR4_X1 U21921 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18833) );
  NAND4_X1 U21922 ( .A1(n18836), .A2(n18835), .A3(n18834), .A4(n18833), .ZN(
        n18837) );
  NOR2_X1 U21923 ( .A1(n18838), .A2(n18837), .ZN(n18845) );
  INV_X1 U21924 ( .A(n18845), .ZN(n18844) );
  NOR2_X1 U21925 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18844), .ZN(n18839) );
  INV_X1 U21926 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19907) );
  AOI22_X1 U21927 ( .A1(n18839), .A2(n19066), .B1(n18844), .B2(n19907), .ZN(
        P2_U2820) );
  OR3_X1 U21928 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18843) );
  INV_X1 U21929 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19905) );
  AOI22_X1 U21930 ( .A1(n18839), .A2(n18843), .B1(n18844), .B2(n19905), .ZN(
        P2_U2821) );
  INV_X1 U21931 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19910) );
  NAND2_X1 U21932 ( .A1(n18839), .A2(n19910), .ZN(n18842) );
  OAI21_X1 U21933 ( .B1(n12061), .B2(n19066), .A(n18845), .ZN(n18840) );
  OAI21_X1 U21934 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18845), .A(n18840), 
        .ZN(n18841) );
  OAI221_X1 U21935 ( .B1(n18842), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18842), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18841), .ZN(P2_U2822) );
  INV_X1 U21936 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19903) );
  OAI221_X1 U21937 ( .B1(n18845), .B2(n19903), .C1(n18844), .C2(n18843), .A(
        n18842), .ZN(P2_U2823) );
  AOI22_X1 U21938 ( .A1(n18847), .A2(n19075), .B1(n18846), .B2(n19069), .ZN(
        n18855) );
  AOI211_X1 U21939 ( .C1(n18849), .C2(n18848), .A(n9910), .B(n19834), .ZN(
        n18853) );
  AOI22_X1 U21940 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19053), .ZN(n18850) );
  OAI21_X1 U21941 ( .B1(n18851), .B2(n19072), .A(n18850), .ZN(n18852) );
  AOI211_X1 U21942 ( .C1(n19081), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n18853), .B(n18852), .ZN(n18854) );
  NAND2_X1 U21943 ( .A1(n18855), .A2(n18854), .ZN(P2_U2834) );
  NOR2_X1 U21944 ( .A1(n18869), .A2(n18868), .ZN(n18867) );
  NOR2_X1 U21945 ( .A1(n10004), .A2(n18867), .ZN(n18857) );
  AOI211_X1 U21946 ( .C1(n18858), .C2(n18857), .A(n18856), .B(n19834), .ZN(
        n18863) );
  AOI22_X1 U21947 ( .A1(P2_EBX_REG_20__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19053), .ZN(n18860) );
  NAND2_X1 U21948 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19081), .ZN(
        n18859) );
  OAI211_X1 U21949 ( .C1(n19072), .C2(n18861), .A(n18860), .B(n18859), .ZN(
        n18862) );
  AOI211_X1 U21950 ( .C1(n19069), .C2(n9883), .A(n18863), .B(n18862), .ZN(
        n18864) );
  OAI21_X1 U21951 ( .B1(n18865), .B2(n19046), .A(n18864), .ZN(P2_U2835) );
  INV_X1 U21952 ( .A(n18866), .ZN(n18875) );
  AOI211_X1 U21953 ( .C1(n18869), .C2(n18868), .A(n18867), .B(n19834), .ZN(
        n18874) );
  AOI21_X1 U21954 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19047), .A(n19016), .ZN(
        n18871) );
  AOI22_X1 U21955 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_19__SCAN_IN), .B2(n19053), .ZN(n18870) );
  OAI211_X1 U21956 ( .C1(n18872), .C2(n19072), .A(n18871), .B(n18870), .ZN(
        n18873) );
  AOI211_X1 U21957 ( .C1(n19075), .C2(n18875), .A(n18874), .B(n18873), .ZN(
        n18876) );
  OAI21_X1 U21958 ( .B1(n18877), .B2(n19055), .A(n18876), .ZN(P2_U2836) );
  AOI22_X1 U21959 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19053), .ZN(n18878) );
  OAI21_X1 U21960 ( .B1(n18879), .B2(n19072), .A(n18878), .ZN(n18880) );
  AOI211_X1 U21961 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18880), .ZN(n18887) );
  NOR2_X1 U21962 ( .A1(n10004), .A2(n18881), .ZN(n18883) );
  XNOR2_X1 U21963 ( .A(n18883), .B(n18882), .ZN(n18884) );
  AOI22_X1 U21964 ( .A1(n18885), .A2(n19069), .B1(n19058), .B2(n18884), .ZN(
        n18886) );
  OAI211_X1 U21965 ( .C1(n18888), .C2(n19046), .A(n18887), .B(n18886), .ZN(
        P2_U2837) );
  NAND2_X1 U21966 ( .A1(n10005), .A2(n18889), .ZN(n18890) );
  XOR2_X1 U21967 ( .A(n18891), .B(n18890), .Z(n18899) );
  AOI22_X1 U21968 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19053), .ZN(n18892) );
  OAI21_X1 U21969 ( .B1(n18893), .B2(n19072), .A(n18892), .ZN(n18894) );
  AOI211_X1 U21970 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18894), .ZN(n18898) );
  AOI22_X1 U21971 ( .A1(n18896), .A2(n19075), .B1(n18895), .B2(n19069), .ZN(
        n18897) );
  OAI211_X1 U21972 ( .C1(n19834), .C2(n18899), .A(n18898), .B(n18897), .ZN(
        P2_U2838) );
  AOI22_X1 U21973 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19053), .ZN(n18900) );
  OAI21_X1 U21974 ( .B1(n18901), .B2(n19072), .A(n18900), .ZN(n18902) );
  AOI211_X1 U21975 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18902), .ZN(n18908) );
  NOR2_X1 U21976 ( .A1(n10004), .A2(n18903), .ZN(n18905) );
  XNOR2_X1 U21977 ( .A(n18905), .B(n18904), .ZN(n18906) );
  AOI22_X1 U21978 ( .A1(n19128), .A2(n19069), .B1(n19058), .B2(n18906), .ZN(
        n18907) );
  OAI211_X1 U21979 ( .C1(n19091), .C2(n19046), .A(n18908), .B(n18907), .ZN(
        P2_U2839) );
  AOI22_X1 U21980 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19053), .ZN(n18909) );
  OAI21_X1 U21981 ( .B1(n18910), .B2(n19072), .A(n18909), .ZN(n18911) );
  AOI211_X1 U21982 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18911), .ZN(n18918) );
  NAND2_X1 U21983 ( .A1(n10005), .A2(n18912), .ZN(n18913) );
  XNOR2_X1 U21984 ( .A(n18914), .B(n18913), .ZN(n18915) );
  AOI22_X1 U21985 ( .A1(n18916), .A2(n19075), .B1(n19058), .B2(n18915), .ZN(
        n18917) );
  OAI211_X1 U21986 ( .C1(n19137), .C2(n19055), .A(n18918), .B(n18917), .ZN(
        P2_U2840) );
  AOI22_X1 U21987 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19053), .ZN(n18919) );
  OAI21_X1 U21988 ( .B1(n18920), .B2(n19072), .A(n18919), .ZN(n18921) );
  AOI211_X1 U21989 ( .C1(P2_EBX_REG_14__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18921), .ZN(n18926) );
  NOR2_X1 U21990 ( .A1(n10004), .A2(n18927), .ZN(n18923) );
  XNOR2_X1 U21991 ( .A(n18923), .B(n18922), .ZN(n18924) );
  AOI22_X1 U21992 ( .A1(n19138), .A2(n19069), .B1(n19058), .B2(n18924), .ZN(
        n18925) );
  OAI211_X1 U21993 ( .C1(n19096), .C2(n19046), .A(n18926), .B(n18925), .ZN(
        P2_U2841) );
  INV_X1 U21994 ( .A(n19079), .ZN(n18948) );
  AOI211_X1 U21995 ( .C1(n18934), .C2(n18928), .A(n18927), .B(n18948), .ZN(
        n18932) );
  AOI22_X1 U21996 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_13__SCAN_IN), .B2(n19053), .ZN(n18929) );
  OAI211_X1 U21997 ( .C1(n18930), .C2(n19049), .A(n18929), .B(n16232), .ZN(
        n18931) );
  AOI211_X1 U21998 ( .C1(n18991), .C2(n18933), .A(n18932), .B(n18931), .ZN(
        n18937) );
  NOR2_X1 U21999 ( .A1(n10005), .A2(n19834), .ZN(n19080) );
  AOI22_X1 U22000 ( .A1(n18935), .A2(n19075), .B1(n18934), .B2(n19080), .ZN(
        n18936) );
  OAI211_X1 U22001 ( .C1(n19143), .C2(n19055), .A(n18937), .B(n18936), .ZN(
        P2_U2842) );
  NOR2_X1 U22002 ( .A1(n10004), .A2(n18949), .ZN(n18939) );
  XOR2_X1 U22003 ( .A(n18939), .B(n18938), .Z(n18946) );
  AOI22_X1 U22004 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19053), .ZN(n18940) );
  OAI21_X1 U22005 ( .B1(n18941), .B2(n19072), .A(n18940), .ZN(n18942) );
  AOI211_X1 U22006 ( .C1(P2_EBX_REG_12__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18942), .ZN(n18945) );
  AOI22_X1 U22007 ( .A1(n18943), .A2(n19075), .B1(n19144), .B2(n19069), .ZN(
        n18944) );
  OAI211_X1 U22008 ( .C1(n19834), .C2(n18946), .A(n18945), .B(n18944), .ZN(
        P2_U2843) );
  INV_X1 U22009 ( .A(n18947), .ZN(n18960) );
  AOI211_X1 U22010 ( .C1(n18958), .C2(n18950), .A(n18949), .B(n18948), .ZN(
        n18957) );
  AOI22_X1 U22011 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19053), .ZN(n18951) );
  OAI211_X1 U22012 ( .C1(n19149), .C2(n19055), .A(n18951), .B(n16232), .ZN(
        n18952) );
  AOI21_X1 U22013 ( .B1(n18953), .B2(n18991), .A(n18952), .ZN(n18954) );
  OAI21_X1 U22014 ( .B1(n18955), .B2(n19049), .A(n18954), .ZN(n18956) );
  AOI211_X1 U22015 ( .C1(n19080), .C2(n18958), .A(n18957), .B(n18956), .ZN(
        n18959) );
  OAI21_X1 U22016 ( .B1(n18960), .B2(n19046), .A(n18959), .ZN(P2_U2844) );
  AOI22_X1 U22017 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19053), .ZN(n18961) );
  OAI21_X1 U22018 ( .B1(n18962), .B2(n19072), .A(n18961), .ZN(n18963) );
  AOI211_X1 U22019 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18963), .ZN(n18969) );
  NOR2_X1 U22020 ( .A1(n10004), .A2(n18964), .ZN(n18966) );
  XNOR2_X1 U22021 ( .A(n18966), .B(n18965), .ZN(n18967) );
  AOI22_X1 U22022 ( .A1(n19104), .A2(n19075), .B1(n19058), .B2(n18967), .ZN(
        n18968) );
  OAI211_X1 U22023 ( .C1(n19152), .C2(n19055), .A(n18969), .B(n18968), .ZN(
        P2_U2845) );
  AOI22_X1 U22024 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19053), .B1(n18991), 
        .B2(n18970), .ZN(n18971) );
  OAI21_X1 U22025 ( .B1(n18972), .B2(n19049), .A(n18971), .ZN(n18973) );
  AOI211_X1 U22026 ( .C1(P2_EBX_REG_9__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18973), .ZN(n18980) );
  NAND2_X1 U22027 ( .A1(n10005), .A2(n18974), .ZN(n18975) );
  XNOR2_X1 U22028 ( .A(n18976), .B(n18975), .ZN(n18977) );
  AOI22_X1 U22029 ( .A1(n18978), .A2(n19069), .B1(n19058), .B2(n18977), .ZN(
        n18979) );
  OAI211_X1 U22030 ( .C1(n18981), .C2(n19046), .A(n18980), .B(n18979), .ZN(
        P2_U2846) );
  AOI22_X1 U22031 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19053), .ZN(n18982) );
  OAI21_X1 U22032 ( .B1(n18983), .B2(n19072), .A(n18982), .ZN(n18984) );
  AOI211_X1 U22033 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18984), .ZN(n18990) );
  NOR2_X1 U22034 ( .A1(n10004), .A2(n18985), .ZN(n18987) );
  XNOR2_X1 U22035 ( .A(n18987), .B(n18986), .ZN(n18988) );
  AOI22_X1 U22036 ( .A1(n19069), .A2(n19155), .B1(n19058), .B2(n18988), .ZN(
        n18989) );
  OAI211_X1 U22037 ( .C1(n19046), .C2(n19115), .A(n18990), .B(n18989), .ZN(
        P2_U2847) );
  AOI22_X1 U22038 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19053), .B1(n18992), 
        .B2(n18991), .ZN(n18993) );
  OAI21_X1 U22039 ( .B1(n18994), .B2(n19049), .A(n18993), .ZN(n18995) );
  AOI211_X1 U22040 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n18995), .ZN(n19002) );
  NAND2_X1 U22041 ( .A1(n10005), .A2(n18996), .ZN(n18997) );
  XNOR2_X1 U22042 ( .A(n18998), .B(n18997), .ZN(n19000) );
  AOI22_X1 U22043 ( .A1(n19058), .A2(n19000), .B1(n19075), .B2(n18999), .ZN(
        n19001) );
  OAI211_X1 U22044 ( .C1(n19055), .C2(n19160), .A(n19002), .B(n19001), .ZN(
        P2_U2848) );
  AOI22_X1 U22045 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19053), .ZN(n19003) );
  OAI21_X1 U22046 ( .B1(n19004), .B2(n19072), .A(n19003), .ZN(n19005) );
  AOI211_X1 U22047 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n19005), .ZN(n19012) );
  NOR2_X1 U22048 ( .A1(n10004), .A2(n19006), .ZN(n19008) );
  XNOR2_X1 U22049 ( .A(n19008), .B(n19007), .ZN(n19010) );
  AOI22_X1 U22050 ( .A1(n19058), .A2(n19010), .B1(n19075), .B2(n19009), .ZN(
        n19011) );
  OAI211_X1 U22051 ( .C1(n19055), .C2(n19163), .A(n19012), .B(n19011), .ZN(
        P2_U2849) );
  AOI22_X1 U22052 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19081), .B1(
        P2_REIP_REG_5__SCAN_IN), .B2(n19053), .ZN(n19013) );
  OAI21_X1 U22053 ( .B1(n19014), .B2(n19072), .A(n19013), .ZN(n19015) );
  AOI211_X1 U22054 ( .C1(P2_EBX_REG_5__SCAN_IN), .C2(n19047), .A(n19016), .B(
        n19015), .ZN(n19023) );
  NAND2_X1 U22055 ( .A1(n10005), .A2(n19017), .ZN(n19018) );
  XNOR2_X1 U22056 ( .A(n19019), .B(n19018), .ZN(n19021) );
  AOI22_X1 U22057 ( .A1(n19058), .A2(n19021), .B1(n19075), .B2(n19020), .ZN(
        n19022) );
  OAI211_X1 U22058 ( .C1(n19055), .C2(n19171), .A(n19023), .B(n19022), .ZN(
        P2_U2850) );
  OR2_X1 U22059 ( .A1(n19025), .A2(n19024), .ZN(n19026) );
  NAND2_X1 U22060 ( .A1(n19026), .A2(n13223), .ZN(n19232) );
  NAND3_X1 U22061 ( .A1(n19027), .A2(n19029), .A3(n10096), .ZN(n19030) );
  NAND2_X1 U22062 ( .A1(n13258), .A2(n19030), .ZN(n19175) );
  INV_X1 U22063 ( .A(n19175), .ZN(n19039) );
  AOI21_X1 U22064 ( .B1(n19032), .B2(n13500), .A(n19031), .ZN(n19258) );
  INV_X1 U22065 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19034) );
  AOI22_X1 U22066 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n19047), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19053), .ZN(n19033) );
  OAI211_X1 U22067 ( .C1(n19034), .C2(n19049), .A(n16232), .B(n19033), .ZN(
        n19035) );
  AOI21_X1 U22068 ( .B1(n19069), .B2(n19258), .A(n19035), .ZN(n19036) );
  OAI21_X1 U22069 ( .B1(n19037), .B2(n19072), .A(n19036), .ZN(n19038) );
  AOI21_X1 U22070 ( .B1(n19039), .B2(n19077), .A(n19038), .ZN(n19045) );
  INV_X1 U22071 ( .A(n19238), .ZN(n19043) );
  NOR2_X1 U22072 ( .A1(n10004), .A2(n19040), .ZN(n19042) );
  AOI21_X1 U22073 ( .B1(n19043), .B2(n19042), .A(n19834), .ZN(n19041) );
  OAI21_X1 U22074 ( .B1(n19043), .B2(n19042), .A(n19041), .ZN(n19044) );
  OAI211_X1 U22075 ( .C1(n19232), .C2(n19046), .A(n19045), .B(n19044), .ZN(
        P2_U2851) );
  INV_X1 U22076 ( .A(n19080), .ZN(n19062) );
  NAND2_X1 U22077 ( .A1(n19047), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n19048) );
  OAI21_X1 U22078 ( .B1(n19049), .B2(n13908), .A(n19048), .ZN(n19052) );
  NOR2_X1 U22079 ( .A1(n19050), .A2(n19072), .ZN(n19051) );
  AOI211_X1 U22080 ( .C1(n19053), .C2(P2_REIP_REG_1__SCAN_IN), .A(n19052), .B(
        n19051), .ZN(n19054) );
  OAI21_X1 U22081 ( .B1(n19056), .B2(n19055), .A(n19054), .ZN(n19057) );
  AOI21_X1 U22082 ( .B1(n12112), .B2(n19075), .A(n19057), .ZN(n19061) );
  AOI22_X1 U22083 ( .A1(n19059), .A2(n19058), .B1(n19943), .B2(n19077), .ZN(
        n19060) );
  OAI211_X1 U22084 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19062), .A(
        n19061), .B(n19060), .ZN(P2_U2854) );
  INV_X1 U22085 ( .A(n19063), .ZN(n19073) );
  OAI22_X1 U22086 ( .A1(n19067), .A2(n19066), .B1(n19065), .B2(n19064), .ZN(
        n19068) );
  AOI21_X1 U22087 ( .B1(n19070), .B2(n19069), .A(n19068), .ZN(n19071) );
  OAI21_X1 U22088 ( .B1(n19073), .B2(n19072), .A(n19071), .ZN(n19074) );
  AOI21_X1 U22089 ( .B1(n19076), .B2(n19075), .A(n19074), .ZN(n19084) );
  AOI22_X1 U22090 ( .A1(n19079), .A2(n19078), .B1(n19527), .B2(n19077), .ZN(
        n19083) );
  OAI21_X1 U22091 ( .B1(n19081), .B2(n19080), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19082) );
  NAND3_X1 U22092 ( .A1(n19084), .A2(n19083), .A3(n19082), .ZN(P2_U2855) );
  NOR2_X1 U22093 ( .A1(n19086), .A2(n19085), .ZN(n19087) );
  OR2_X1 U22094 ( .A1(n13677), .A2(n19087), .ZN(n19131) );
  INV_X1 U22095 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n19088) );
  OAI22_X1 U22096 ( .A1(n19131), .A2(n19117), .B1(n19121), .B2(n19088), .ZN(
        n19089) );
  INV_X1 U22097 ( .A(n19089), .ZN(n19090) );
  OAI21_X1 U22098 ( .B1(n19116), .B2(n19091), .A(n19090), .ZN(P2_U2871) );
  XOR2_X1 U22099 ( .A(n19093), .B(n19092), .Z(n19094) );
  AOI22_X1 U22100 ( .A1(n19094), .A2(n19107), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19116), .ZN(n19095) );
  OAI21_X1 U22101 ( .B1(n19096), .B2(n19116), .A(n19095), .ZN(P2_U2873) );
  XOR2_X1 U22102 ( .A(n19098), .B(n19097), .Z(n19099) );
  AOI22_X1 U22103 ( .A1(n19099), .A2(n19107), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19116), .ZN(n19100) );
  OAI21_X1 U22104 ( .B1(n19101), .B2(n19116), .A(n19100), .ZN(P2_U2875) );
  XNOR2_X1 U22105 ( .A(n19103), .B(n19102), .ZN(n19105) );
  AOI22_X1 U22106 ( .A1(n19105), .A2(n19107), .B1(n19121), .B2(n19104), .ZN(
        n19106) );
  OAI21_X1 U22107 ( .B1(n19121), .B2(n12509), .A(n19106), .ZN(P2_U2877) );
  OAI21_X1 U22108 ( .B1(n19109), .B2(n19108), .A(n19107), .ZN(n19112) );
  OAI22_X1 U22109 ( .A1(n19112), .A2(n19111), .B1(n19121), .B2(n19110), .ZN(
        n19113) );
  INV_X1 U22110 ( .A(n19113), .ZN(n19114) );
  OAI21_X1 U22111 ( .B1(n19115), .B2(n19116), .A(n19114), .ZN(P2_U2879) );
  OAI22_X1 U22112 ( .A1(n19175), .A2(n19117), .B1(n19116), .B2(n19232), .ZN(
        n19118) );
  INV_X1 U22113 ( .A(n19118), .ZN(n19119) );
  OAI21_X1 U22114 ( .B1(n19121), .B2(n19120), .A(n19119), .ZN(P2_U2883) );
  AOI22_X1 U22115 ( .A1(n15969), .A2(n19187), .B1(n19126), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19123) );
  AOI22_X1 U22116 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19186), .B1(n19127), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19122) );
  NAND2_X1 U22117 ( .A1(n19123), .A2(n19122), .ZN(P2_U2888) );
  AOI22_X1 U22118 ( .A1(n19125), .A2(n19124), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19186), .ZN(n19135) );
  AOI22_X1 U22119 ( .A1(n19127), .A2(BUF1_REG_16__SCAN_IN), .B1(n19126), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19134) );
  INV_X1 U22120 ( .A(n19187), .ZN(n19130) );
  INV_X1 U22121 ( .A(n19128), .ZN(n19129) );
  OAI22_X1 U22122 ( .A1(n19131), .A2(n19191), .B1(n19130), .B2(n19129), .ZN(
        n19132) );
  INV_X1 U22123 ( .A(n19132), .ZN(n19133) );
  NAND3_X1 U22124 ( .A1(n19135), .A2(n19134), .A3(n19133), .ZN(P2_U2903) );
  OAI222_X1 U22125 ( .A1(n19137), .A2(n19172), .B1(n12872), .B2(n19162), .C1(
        n19136), .C2(n19195), .ZN(P2_U2904) );
  INV_X1 U22126 ( .A(n19138), .ZN(n19141) );
  AOI22_X1 U22127 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19186), .B1(n19139), 
        .B2(n19164), .ZN(n19140) );
  OAI21_X1 U22128 ( .B1(n19172), .B2(n19141), .A(n19140), .ZN(P2_U2905) );
  INV_X1 U22129 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19202) );
  OAI222_X1 U22130 ( .A1(n19143), .A2(n19172), .B1(n19202), .B2(n19162), .C1(
        n19195), .C2(n19142), .ZN(P2_U2906) );
  INV_X1 U22131 ( .A(n19144), .ZN(n19147) );
  AOI22_X1 U22132 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19186), .B1(n19145), 
        .B2(n19164), .ZN(n19146) );
  OAI21_X1 U22133 ( .B1(n19172), .B2(n19147), .A(n19146), .ZN(P2_U2907) );
  INV_X1 U22134 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19206) );
  OAI222_X1 U22135 ( .A1(n19149), .A2(n19172), .B1(n19206), .B2(n19162), .C1(
        n19195), .C2(n19148), .ZN(P2_U2908) );
  AOI22_X1 U22136 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19186), .B1(n19150), 
        .B2(n19164), .ZN(n19151) );
  OAI21_X1 U22137 ( .B1(n19172), .B2(n19152), .A(n19151), .ZN(P2_U2909) );
  INV_X1 U22138 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19210) );
  OAI222_X1 U22139 ( .A1(n19154), .A2(n19172), .B1(n19210), .B2(n19162), .C1(
        n19195), .C2(n19153), .ZN(P2_U2910) );
  INV_X1 U22140 ( .A(n19155), .ZN(n19158) );
  AOI22_X1 U22141 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19186), .B1(n19156), .B2(
        n19164), .ZN(n19157) );
  OAI21_X1 U22142 ( .B1(n19172), .B2(n19158), .A(n19157), .ZN(P2_U2911) );
  INV_X1 U22143 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19214) );
  OAI222_X1 U22144 ( .A1(n19160), .A2(n19172), .B1(n19214), .B2(n19162), .C1(
        n19195), .C2(n19159), .ZN(P2_U2912) );
  INV_X1 U22145 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19216) );
  INV_X1 U22146 ( .A(n19161), .ZN(n19293) );
  OAI222_X1 U22147 ( .A1(n19163), .A2(n19172), .B1(n19216), .B2(n19162), .C1(
        n19195), .C2(n19293), .ZN(P2_U2913) );
  AOI22_X1 U22148 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19186), .B1(n19165), .B2(
        n19164), .ZN(n19170) );
  AOI21_X1 U22149 ( .B1(n19935), .B2(n19917), .A(n19166), .ZN(n19182) );
  XNOR2_X1 U22150 ( .A(n19925), .B(n19167), .ZN(n19181) );
  NOR2_X1 U22151 ( .A1(n19182), .A2(n19181), .ZN(n19180) );
  AOI21_X1 U22152 ( .B1(n19925), .B2(n19167), .A(n19180), .ZN(n19168) );
  NOR2_X1 U22153 ( .A1(n19168), .A2(n19258), .ZN(n19174) );
  OR3_X1 U22154 ( .A1(n19174), .A2(n19175), .A3(n19191), .ZN(n19169) );
  OAI211_X1 U22155 ( .C1(n19172), .C2(n19171), .A(n19170), .B(n19169), .ZN(
        P2_U2914) );
  INV_X1 U22156 ( .A(n19173), .ZN(n19284) );
  AOI22_X1 U22157 ( .A1(n19187), .A2(n19258), .B1(n19186), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19179) );
  XOR2_X1 U22158 ( .A(n19175), .B(n19174), .Z(n19177) );
  NAND2_X1 U22159 ( .A1(n19177), .A2(n19176), .ZN(n19178) );
  OAI211_X1 U22160 ( .C1(n19284), .C2(n19195), .A(n19179), .B(n19178), .ZN(
        P2_U2915) );
  AOI22_X1 U22161 ( .A1(n19187), .A2(n19931), .B1(n19186), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19185) );
  AOI21_X1 U22162 ( .B1(n19182), .B2(n19181), .A(n19180), .ZN(n19183) );
  OR2_X1 U22163 ( .A1(n19183), .A2(n19191), .ZN(n19184) );
  OAI211_X1 U22164 ( .C1(n19279), .C2(n19195), .A(n19185), .B(n19184), .ZN(
        P2_U2916) );
  AOI22_X1 U22165 ( .A1(n19187), .A2(n19947), .B1(n19186), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19194) );
  AOI21_X1 U22166 ( .B1(n19190), .B2(n19189), .A(n19188), .ZN(n19192) );
  OR2_X1 U22167 ( .A1(n19192), .A2(n19191), .ZN(n19193) );
  OAI211_X1 U22168 ( .C1(n19269), .C2(n19195), .A(n19194), .B(n19193), .ZN(
        P2_U2918) );
  AND2_X1 U22169 ( .A1(n19196), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22170 ( .A1(n13117), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22171 ( .B1(n12872), .B2(n19229), .A(n19198), .ZN(P2_U2936) );
  AOI22_X1 U22172 ( .A1(n13117), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19199) );
  OAI21_X1 U22173 ( .B1(n19200), .B2(n19229), .A(n19199), .ZN(P2_U2937) );
  AOI22_X1 U22174 ( .A1(n13117), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19201) );
  OAI21_X1 U22175 ( .B1(n19202), .B2(n19229), .A(n19201), .ZN(P2_U2938) );
  AOI22_X1 U22176 ( .A1(n13117), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19203) );
  OAI21_X1 U22177 ( .B1(n19204), .B2(n19229), .A(n19203), .ZN(P2_U2939) );
  AOI22_X1 U22178 ( .A1(n13117), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19205) );
  OAI21_X1 U22179 ( .B1(n19206), .B2(n19229), .A(n19205), .ZN(P2_U2940) );
  AOI22_X1 U22180 ( .A1(n13117), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22181 ( .B1(n19208), .B2(n19229), .A(n19207), .ZN(P2_U2941) );
  AOI22_X1 U22182 ( .A1(n13117), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19209) );
  OAI21_X1 U22183 ( .B1(n19210), .B2(n19229), .A(n19209), .ZN(P2_U2942) );
  AOI22_X1 U22184 ( .A1(n13117), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22185 ( .B1(n19212), .B2(n19229), .A(n19211), .ZN(P2_U2943) );
  AOI22_X1 U22186 ( .A1(n13117), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19213) );
  OAI21_X1 U22187 ( .B1(n19214), .B2(n19229), .A(n19213), .ZN(P2_U2944) );
  AOI22_X1 U22188 ( .A1(n13117), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U22189 ( .B1(n19216), .B2(n19229), .A(n19215), .ZN(P2_U2945) );
  INV_X1 U22190 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19218) );
  AOI22_X1 U22191 ( .A1(n13117), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19217) );
  OAI21_X1 U22192 ( .B1(n19218), .B2(n19229), .A(n19217), .ZN(P2_U2946) );
  INV_X1 U22193 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19220) );
  AOI22_X1 U22194 ( .A1(n13117), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19219) );
  OAI21_X1 U22195 ( .B1(n19220), .B2(n19229), .A(n19219), .ZN(P2_U2947) );
  INV_X1 U22196 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U22197 ( .A1(n13117), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19221) );
  OAI21_X1 U22198 ( .B1(n19222), .B2(n19229), .A(n19221), .ZN(P2_U2948) );
  INV_X1 U22199 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19224) );
  AOI22_X1 U22200 ( .A1(n13117), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19223) );
  OAI21_X1 U22201 ( .B1(n19224), .B2(n19229), .A(n19223), .ZN(P2_U2949) );
  INV_X1 U22202 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19226) );
  AOI22_X1 U22203 ( .A1(n13117), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19225) );
  OAI21_X1 U22204 ( .B1(n19226), .B2(n19229), .A(n19225), .ZN(P2_U2950) );
  AOI22_X1 U22205 ( .A1(n13117), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19227), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19228) );
  OAI21_X1 U22206 ( .B1(n12874), .B2(n19229), .A(n19228), .ZN(P2_U2951) );
  AOI22_X1 U22207 ( .A1(n19239), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n12763), .ZN(n19237) );
  XOR2_X1 U22208 ( .A(n19231), .B(n19230), .Z(n19264) );
  INV_X1 U22209 ( .A(n19232), .ZN(n19254) );
  NAND2_X1 U22210 ( .A1(n19234), .A2(n19233), .ZN(n19235) );
  XNOR2_X1 U22211 ( .A(n19235), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19261) );
  AOI222_X1 U22212 ( .A1(n19264), .A2(n19240), .B1(n19250), .B2(n19254), .C1(
        n19242), .C2(n19261), .ZN(n19236) );
  OAI211_X1 U22213 ( .C1(n19247), .C2(n19238), .A(n19237), .B(n19236), .ZN(
        P2_U3010) );
  AOI22_X1 U22214 ( .A1(n19241), .A2(n19240), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19239), .ZN(n19253) );
  NAND2_X1 U22215 ( .A1(n19243), .A2(n19242), .ZN(n19246) );
  INV_X1 U22216 ( .A(n19244), .ZN(n19245) );
  OAI211_X1 U22217 ( .C1(n19248), .C2(n19247), .A(n19246), .B(n19245), .ZN(
        n19249) );
  AOI21_X1 U22218 ( .B1(n19251), .B2(n19250), .A(n19249), .ZN(n19252) );
  NAND2_X1 U22219 ( .A1(n19253), .A2(n19252), .ZN(P2_U3012) );
  AOI22_X1 U22220 ( .A1(n19256), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n19255), .B2(n19254), .ZN(n19268) );
  AOI22_X1 U22221 ( .A1(n19260), .A2(n19259), .B1(n19258), .B2(n19257), .ZN(
        n19267) );
  AOI22_X1 U22222 ( .A1(n19264), .A2(n19263), .B1(n19262), .B2(n19261), .ZN(
        n19266) );
  NAND2_X1 U22223 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n12763), .ZN(n19265) );
  NAND4_X1 U22224 ( .A1(n19268), .A2(n19267), .A3(n19266), .A4(n19265), .ZN(
        P2_U3042) );
  AOI22_X1 U22225 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19294), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19295), .ZN(n19787) );
  AOI22_X1 U22226 ( .A1(n19741), .A2(n19823), .B1(n19292), .B2(n19782), .ZN(
        n19271) );
  NOR2_X2 U22227 ( .A1(n19269), .A2(n19503), .ZN(n19783) );
  AOI22_X1 U22228 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19294), .ZN(n19744) );
  INV_X1 U22229 ( .A(n19744), .ZN(n19784) );
  AOI22_X1 U22230 ( .A1(n19783), .A2(n19296), .B1(n19352), .B2(n19784), .ZN(
        n19270) );
  OAI211_X1 U22231 ( .C1(n19300), .C2(n19272), .A(n19271), .B(n19270), .ZN(
        P2_U3049) );
  AOI22_X1 U22232 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19294), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19295), .ZN(n19793) );
  INV_X1 U22233 ( .A(n19793), .ZN(n19700) );
  NOR2_X2 U22234 ( .A1(n19273), .A2(n19287), .ZN(n19788) );
  AOI22_X1 U22235 ( .A1(n19700), .A2(n19823), .B1(n19292), .B2(n19788), .ZN(
        n19276) );
  NOR2_X2 U22236 ( .A1(n19274), .A2(n19503), .ZN(n19789) );
  AOI22_X1 U22237 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19294), .ZN(n19703) );
  INV_X1 U22238 ( .A(n19703), .ZN(n19790) );
  AOI22_X1 U22239 ( .A1(n19789), .A2(n19296), .B1(n19352), .B2(n19790), .ZN(
        n19275) );
  OAI211_X1 U22240 ( .C1(n19300), .C2(n19277), .A(n19276), .B(n19275), .ZN(
        P2_U3050) );
  AOI22_X1 U22241 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19294), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19295), .ZN(n19799) );
  INV_X1 U22242 ( .A(n19799), .ZN(n19704) );
  AND2_X1 U22243 ( .A1(n19278), .A2(n19291), .ZN(n19794) );
  AOI22_X1 U22244 ( .A1(n19704), .A2(n19823), .B1(n19292), .B2(n19794), .ZN(
        n19281) );
  NOR2_X2 U22245 ( .A1(n19279), .A2(n19503), .ZN(n19795) );
  AOI22_X1 U22246 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19294), .ZN(n19707) );
  AOI22_X1 U22247 ( .A1(n19795), .A2(n19296), .B1(n19352), .B2(n19796), .ZN(
        n19280) );
  OAI211_X1 U22248 ( .C1(n19300), .C2(n19282), .A(n19281), .B(n19280), .ZN(
        P2_U3051) );
  AOI22_X1 U22249 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19294), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19295), .ZN(n19805) );
  INV_X1 U22250 ( .A(n19805), .ZN(n19708) );
  AOI22_X1 U22251 ( .A1(n19708), .A2(n19823), .B1(n19292), .B2(n19800), .ZN(
        n19286) );
  NOR2_X2 U22252 ( .A1(n19284), .A2(n19503), .ZN(n19801) );
  AOI22_X1 U22253 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19294), .ZN(n19711) );
  AOI22_X1 U22254 ( .A1(n19801), .A2(n19296), .B1(n19352), .B2(n19802), .ZN(
        n19285) );
  OAI211_X1 U22255 ( .C1(n19300), .C2(n14178), .A(n19286), .B(n19285), .ZN(
        P2_U3052) );
  AOI22_X1 U22256 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19294), .ZN(n19811) );
  INV_X1 U22257 ( .A(n19811), .ZN(n19712) );
  NOR2_X2 U22258 ( .A1(n12264), .A2(n19287), .ZN(n19806) );
  AOI22_X1 U22259 ( .A1(n19712), .A2(n19823), .B1(n19292), .B2(n19806), .ZN(
        n19290) );
  NOR2_X2 U22260 ( .A1(n19288), .A2(n19503), .ZN(n19807) );
  AOI22_X1 U22261 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19294), .ZN(n19715) );
  AOI22_X1 U22262 ( .A1(n19807), .A2(n19296), .B1(n19352), .B2(n19808), .ZN(
        n19289) );
  OAI211_X1 U22263 ( .C1(n19300), .C2(n14204), .A(n19290), .B(n19289), .ZN(
        P2_U3053) );
  AOI22_X1 U22264 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19294), .ZN(n19817) );
  INV_X1 U22265 ( .A(n19817), .ZN(n19716) );
  AND2_X1 U22266 ( .A1(n13016), .A2(n19291), .ZN(n19812) );
  AOI22_X1 U22267 ( .A1(n19716), .A2(n19823), .B1(n19292), .B2(n19812), .ZN(
        n19298) );
  NOR2_X2 U22268 ( .A1(n19293), .A2(n19503), .ZN(n19813) );
  AOI22_X1 U22269 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19295), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19294), .ZN(n19719) );
  AOI22_X1 U22270 ( .A1(n19813), .A2(n19296), .B1(n19352), .B2(n19814), .ZN(
        n19297) );
  OAI211_X1 U22271 ( .C1(n19300), .C2(n19299), .A(n19298), .B(n19297), .ZN(
        P2_U3054) );
  NAND2_X1 U22272 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19949), .ZN(
        n19558) );
  INV_X1 U22273 ( .A(n19357), .ZN(n19387) );
  NOR2_X1 U22274 ( .A1(n19558), .A2(n19387), .ZN(n19314) );
  OR2_X1 U22275 ( .A1(n19314), .A2(n19979), .ZN(n19301) );
  NOR2_X1 U22276 ( .A1(n19302), .A2(n19301), .ZN(n19310) );
  INV_X1 U22277 ( .A(n19303), .ZN(n19500) );
  INV_X1 U22278 ( .A(n19311), .ZN(n19304) );
  NOR2_X1 U22279 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19304), .ZN(n19305) );
  INV_X1 U22280 ( .A(n19769), .ZN(n19306) );
  INV_X1 U22281 ( .A(n19314), .ZN(n19347) );
  OAI22_X1 U22282 ( .A1(n19350), .A2(n19307), .B1(n19306), .B2(n19347), .ZN(
        n19308) );
  INV_X1 U22283 ( .A(n19308), .ZN(n19316) );
  NAND2_X1 U22284 ( .A1(n19925), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19928) );
  INV_X1 U22285 ( .A(n19928), .ZN(n19501) );
  INV_X1 U22286 ( .A(n19560), .ZN(n19309) );
  NAND2_X1 U22287 ( .A1(n19501), .A2(n19309), .ZN(n19312) );
  AOI21_X1 U22288 ( .B1(n19312), .B2(n19311), .A(n19310), .ZN(n19313) );
  OAI211_X1 U22289 ( .C1(n19314), .C2(n19971), .A(n19313), .B(n19776), .ZN(
        n19353) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19694), .ZN(n19315) );
  OAI211_X1 U22291 ( .C1(n19697), .C2(n19386), .A(n19316), .B(n19315), .ZN(
        P2_U3056) );
  INV_X1 U22292 ( .A(n19783), .ZN(n19318) );
  INV_X1 U22293 ( .A(n19782), .ZN(n19317) );
  OAI22_X1 U22294 ( .A1(n19350), .A2(n19318), .B1(n19317), .B2(n19347), .ZN(
        n19319) );
  INV_X1 U22295 ( .A(n19319), .ZN(n19321) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19741), .ZN(n19320) );
  OAI211_X1 U22297 ( .C1(n19744), .C2(n19386), .A(n19321), .B(n19320), .ZN(
        P2_U3057) );
  INV_X1 U22298 ( .A(n19789), .ZN(n19323) );
  INV_X1 U22299 ( .A(n19788), .ZN(n19322) );
  OAI22_X1 U22300 ( .A1(n19350), .A2(n19323), .B1(n19322), .B2(n19347), .ZN(
        n19324) );
  INV_X1 U22301 ( .A(n19324), .ZN(n19326) );
  AOI22_X1 U22302 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19700), .ZN(n19325) );
  OAI211_X1 U22303 ( .C1(n19703), .C2(n19386), .A(n19326), .B(n19325), .ZN(
        P2_U3058) );
  INV_X1 U22304 ( .A(n19795), .ZN(n19328) );
  INV_X1 U22305 ( .A(n19794), .ZN(n19327) );
  OAI22_X1 U22306 ( .A1(n19350), .A2(n19328), .B1(n19327), .B2(n19347), .ZN(
        n19329) );
  INV_X1 U22307 ( .A(n19329), .ZN(n19331) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19704), .ZN(n19330) );
  OAI211_X1 U22309 ( .C1(n19707), .C2(n19386), .A(n19331), .B(n19330), .ZN(
        P2_U3059) );
  INV_X1 U22310 ( .A(n19801), .ZN(n19333) );
  INV_X1 U22311 ( .A(n19800), .ZN(n19332) );
  OAI22_X1 U22312 ( .A1(n19350), .A2(n19333), .B1(n19332), .B2(n19347), .ZN(
        n19334) );
  INV_X1 U22313 ( .A(n19334), .ZN(n19336) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19708), .ZN(n19335) );
  OAI211_X1 U22315 ( .C1(n19711), .C2(n19386), .A(n19336), .B(n19335), .ZN(
        P2_U3060) );
  INV_X1 U22316 ( .A(n19807), .ZN(n19338) );
  INV_X1 U22317 ( .A(n19806), .ZN(n19337) );
  OAI22_X1 U22318 ( .A1(n19350), .A2(n19338), .B1(n19337), .B2(n19347), .ZN(
        n19339) );
  INV_X1 U22319 ( .A(n19339), .ZN(n19341) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19712), .ZN(n19340) );
  OAI211_X1 U22321 ( .C1(n19715), .C2(n19386), .A(n19341), .B(n19340), .ZN(
        P2_U3061) );
  INV_X1 U22322 ( .A(n19813), .ZN(n19343) );
  INV_X1 U22323 ( .A(n19812), .ZN(n19342) );
  OAI22_X1 U22324 ( .A1(n19350), .A2(n19343), .B1(n19342), .B2(n19347), .ZN(
        n19344) );
  INV_X1 U22325 ( .A(n19344), .ZN(n19346) );
  AOI22_X1 U22326 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19716), .ZN(n19345) );
  OAI211_X1 U22327 ( .C1(n19719), .C2(n19386), .A(n19346), .B(n19345), .ZN(
        P2_U3062) );
  INV_X1 U22328 ( .A(n19819), .ZN(n19348) );
  OAI22_X1 U22329 ( .A1(n19350), .A2(n19349), .B1(n19348), .B2(n19347), .ZN(
        n19351) );
  INV_X1 U22330 ( .A(n19351), .ZN(n19355) );
  INV_X1 U22331 ( .A(n19828), .ZN(n19759) );
  AOI22_X1 U22332 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19353), .B1(
        n19352), .B2(n19759), .ZN(n19354) );
  OAI211_X1 U22333 ( .C1(n19764), .C2(n19386), .A(n19355), .B(n19354), .ZN(
        P2_U3063) );
  INV_X1 U22334 ( .A(n19356), .ZN(n19360) );
  NOR2_X1 U22335 ( .A1(n19949), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19589) );
  NAND2_X1 U22336 ( .A1(n19589), .A2(n19357), .ZN(n19359) );
  AND2_X1 U22337 ( .A1(n19360), .A2(n19359), .ZN(n19358) );
  INV_X1 U22338 ( .A(n19728), .ZN(n19927) );
  NAND2_X1 U22339 ( .A1(n19417), .A2(n19357), .ZN(n19363) );
  OAI22_X1 U22340 ( .A1(n19358), .A2(n19979), .B1(n19927), .B2(n19363), .ZN(
        n19382) );
  INV_X1 U22341 ( .A(n19359), .ZN(n19381) );
  AOI22_X1 U22342 ( .A1(n19382), .A2(n19770), .B1(n19769), .B2(n19381), .ZN(
        n19367) );
  AOI21_X1 U22343 ( .B1(n19360), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19365) );
  OAI21_X1 U22344 ( .B1(n19370), .B2(n19406), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19362) );
  NAND2_X1 U22345 ( .A1(n19363), .A2(n19362), .ZN(n19364) );
  OAI211_X1 U22346 ( .C1(n19381), .C2(n19365), .A(n19364), .B(n19776), .ZN(
        n19383) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19383), .B1(
        n19406), .B2(n19778), .ZN(n19366) );
  OAI211_X1 U22348 ( .C1(n19781), .C2(n19386), .A(n19367), .B(n19366), .ZN(
        P2_U3064) );
  AOI22_X1 U22349 ( .A1(n19382), .A2(n19783), .B1(n19782), .B2(n19381), .ZN(
        n19369) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19383), .B1(
        n19370), .B2(n19741), .ZN(n19368) );
  OAI211_X1 U22351 ( .C1(n19744), .C2(n19416), .A(n19369), .B(n19368), .ZN(
        P2_U3065) );
  AOI22_X1 U22352 ( .A1(n19382), .A2(n19789), .B1(n19788), .B2(n19381), .ZN(
        n19372) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19383), .B1(
        n19370), .B2(n19700), .ZN(n19371) );
  OAI211_X1 U22354 ( .C1(n19703), .C2(n19416), .A(n19372), .B(n19371), .ZN(
        P2_U3066) );
  AOI22_X1 U22355 ( .A1(n19382), .A2(n19795), .B1(n19794), .B2(n19381), .ZN(
        n19374) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19383), .B1(
        n19406), .B2(n19796), .ZN(n19373) );
  OAI211_X1 U22357 ( .C1(n19799), .C2(n19386), .A(n19374), .B(n19373), .ZN(
        P2_U3067) );
  AOI22_X1 U22358 ( .A1(n19382), .A2(n19801), .B1(n19800), .B2(n19381), .ZN(
        n19376) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19383), .B1(
        n19406), .B2(n19802), .ZN(n19375) );
  OAI211_X1 U22360 ( .C1(n19805), .C2(n19386), .A(n19376), .B(n19375), .ZN(
        P2_U3068) );
  AOI22_X1 U22361 ( .A1(n19382), .A2(n19807), .B1(n19806), .B2(n19381), .ZN(
        n19378) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19383), .B1(
        n19406), .B2(n19808), .ZN(n19377) );
  OAI211_X1 U22363 ( .C1(n19811), .C2(n19386), .A(n19378), .B(n19377), .ZN(
        P2_U3069) );
  AOI22_X1 U22364 ( .A1(n19382), .A2(n19813), .B1(n19812), .B2(n19381), .ZN(
        n19380) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19383), .B1(
        n19406), .B2(n19814), .ZN(n19379) );
  OAI211_X1 U22366 ( .C1(n19817), .C2(n19386), .A(n19380), .B(n19379), .ZN(
        P2_U3070) );
  AOI22_X1 U22367 ( .A1(n19382), .A2(n19820), .B1(n19819), .B2(n19381), .ZN(
        n19385) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19383), .B1(
        n19406), .B2(n19822), .ZN(n19384) );
  OAI211_X1 U22369 ( .C1(n19828), .C2(n19386), .A(n19385), .B(n19384), .ZN(
        P2_U3071) );
  NOR2_X1 U22370 ( .A1(n19622), .A2(n19387), .ZN(n19411) );
  AOI22_X1 U22371 ( .A1(n19694), .A2(n19406), .B1(n19769), .B2(n19411), .ZN(
        n19397) );
  OAI21_X1 U22372 ( .B1(n19928), .B2(n19630), .A(n19728), .ZN(n19395) );
  NOR2_X1 U22373 ( .A1(n19949), .A2(n19387), .ZN(n19391) );
  INV_X1 U22374 ( .A(n19392), .ZN(n19389) );
  INV_X1 U22375 ( .A(n19411), .ZN(n19388) );
  OAI211_X1 U22376 ( .C1(n19389), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19927), 
        .B(n19388), .ZN(n19390) );
  OAI211_X1 U22377 ( .C1(n19395), .C2(n19391), .A(n19776), .B(n19390), .ZN(
        n19413) );
  INV_X1 U22378 ( .A(n19391), .ZN(n19394) );
  OAI21_X1 U22379 ( .B1(n19392), .B2(n19411), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19393) );
  OAI21_X1 U22380 ( .B1(n19395), .B2(n19394), .A(n19393), .ZN(n19412) );
  AOI22_X1 U22381 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19413), .B1(
        n19770), .B2(n19412), .ZN(n19396) );
  OAI211_X1 U22382 ( .C1(n19697), .C2(n19443), .A(n19397), .B(n19396), .ZN(
        P2_U3072) );
  AOI22_X1 U22383 ( .A1(n19741), .A2(n19406), .B1(n19411), .B2(n19782), .ZN(
        n19399) );
  AOI22_X1 U22384 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19413), .B1(
        n19783), .B2(n19412), .ZN(n19398) );
  OAI211_X1 U22385 ( .C1(n19744), .C2(n19443), .A(n19399), .B(n19398), .ZN(
        P2_U3073) );
  AOI22_X1 U22386 ( .A1(n19790), .A2(n19446), .B1(n19411), .B2(n19788), .ZN(
        n19401) );
  AOI22_X1 U22387 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19413), .B1(
        n19789), .B2(n19412), .ZN(n19400) );
  OAI211_X1 U22388 ( .C1(n19793), .C2(n19416), .A(n19401), .B(n19400), .ZN(
        P2_U3074) );
  AOI22_X1 U22389 ( .A1(n19704), .A2(n19406), .B1(n19411), .B2(n19794), .ZN(
        n19403) );
  AOI22_X1 U22390 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19413), .B1(
        n19795), .B2(n19412), .ZN(n19402) );
  OAI211_X1 U22391 ( .C1(n19707), .C2(n19443), .A(n19403), .B(n19402), .ZN(
        P2_U3075) );
  AOI22_X1 U22392 ( .A1(n19708), .A2(n19406), .B1(n19411), .B2(n19800), .ZN(
        n19405) );
  AOI22_X1 U22393 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19413), .B1(
        n19801), .B2(n19412), .ZN(n19404) );
  OAI211_X1 U22394 ( .C1(n19711), .C2(n19443), .A(n19405), .B(n19404), .ZN(
        P2_U3076) );
  AOI22_X1 U22395 ( .A1(n19712), .A2(n19406), .B1(n19411), .B2(n19806), .ZN(
        n19408) );
  AOI22_X1 U22396 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19413), .B1(
        n19807), .B2(n19412), .ZN(n19407) );
  OAI211_X1 U22397 ( .C1(n19715), .C2(n19443), .A(n19408), .B(n19407), .ZN(
        P2_U3077) );
  AOI22_X1 U22398 ( .A1(n19814), .A2(n19446), .B1(n19411), .B2(n19812), .ZN(
        n19410) );
  AOI22_X1 U22399 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19413), .B1(
        n19813), .B2(n19412), .ZN(n19409) );
  OAI211_X1 U22400 ( .C1(n19817), .C2(n19416), .A(n19410), .B(n19409), .ZN(
        P2_U3078) );
  AOI22_X1 U22401 ( .A1(n19822), .A2(n19446), .B1(n19819), .B2(n19411), .ZN(
        n19415) );
  AOI22_X1 U22402 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19413), .B1(
        n19820), .B2(n19412), .ZN(n19414) );
  OAI211_X1 U22403 ( .C1(n19828), .C2(n19416), .A(n19415), .B(n19414), .ZN(
        P2_U3079) );
  INV_X1 U22404 ( .A(n19417), .ZN(n19419) );
  NAND2_X1 U22405 ( .A1(n19419), .A2(n19418), .ZN(n19658) );
  NOR2_X1 U22406 ( .A1(n19658), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19428) );
  INV_X1 U22407 ( .A(n19428), .ZN(n19421) );
  NOR2_X1 U22408 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19456), .ZN(
        n19444) );
  OAI21_X1 U22409 ( .B1(n19423), .B2(n19444), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19420) );
  OAI21_X1 U22410 ( .B1(n19927), .B2(n19421), .A(n19420), .ZN(n19445) );
  AOI22_X1 U22411 ( .A1(n19445), .A2(n19770), .B1(n19769), .B2(n19444), .ZN(
        n19430) );
  AOI21_X1 U22412 ( .B1(n19443), .B2(n19464), .A(n19920), .ZN(n19427) );
  OAI21_X1 U22413 ( .B1(n19423), .B2(n19979), .A(n19971), .ZN(n19425) );
  INV_X1 U22414 ( .A(n19444), .ZN(n19424) );
  NAND2_X1 U22415 ( .A1(n19425), .A2(n19424), .ZN(n19426) );
  OAI211_X1 U22416 ( .C1(n19428), .C2(n19427), .A(n19426), .B(n19776), .ZN(
        n19447) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19447), .B1(
        n19474), .B2(n19778), .ZN(n19429) );
  OAI211_X1 U22418 ( .C1(n19781), .C2(n19443), .A(n19430), .B(n19429), .ZN(
        P2_U3080) );
  AOI22_X1 U22419 ( .A1(n19445), .A2(n19783), .B1(n19782), .B2(n19444), .ZN(
        n19432) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19447), .B1(
        n19446), .B2(n19741), .ZN(n19431) );
  OAI211_X1 U22421 ( .C1(n19744), .C2(n19464), .A(n19432), .B(n19431), .ZN(
        P2_U3081) );
  AOI22_X1 U22422 ( .A1(n19445), .A2(n19789), .B1(n19788), .B2(n19444), .ZN(
        n19434) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19447), .B1(
        n19446), .B2(n19700), .ZN(n19433) );
  OAI211_X1 U22424 ( .C1(n19703), .C2(n19464), .A(n19434), .B(n19433), .ZN(
        P2_U3082) );
  AOI22_X1 U22425 ( .A1(n19445), .A2(n19795), .B1(n19794), .B2(n19444), .ZN(
        n19436) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19447), .B1(
        n19474), .B2(n19796), .ZN(n19435) );
  OAI211_X1 U22427 ( .C1(n19799), .C2(n19443), .A(n19436), .B(n19435), .ZN(
        P2_U3083) );
  AOI22_X1 U22428 ( .A1(n19445), .A2(n19801), .B1(n19800), .B2(n19444), .ZN(
        n19438) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19447), .B1(
        n19474), .B2(n19802), .ZN(n19437) );
  OAI211_X1 U22430 ( .C1(n19805), .C2(n19443), .A(n19438), .B(n19437), .ZN(
        P2_U3084) );
  AOI22_X1 U22431 ( .A1(n19445), .A2(n19807), .B1(n19806), .B2(n19444), .ZN(
        n19440) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19447), .B1(
        n19446), .B2(n19712), .ZN(n19439) );
  OAI211_X1 U22433 ( .C1(n19715), .C2(n19464), .A(n19440), .B(n19439), .ZN(
        P2_U3085) );
  AOI22_X1 U22434 ( .A1(n19445), .A2(n19813), .B1(n19812), .B2(n19444), .ZN(
        n19442) );
  AOI22_X1 U22435 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19447), .B1(
        n19474), .B2(n19814), .ZN(n19441) );
  OAI211_X1 U22436 ( .C1(n19817), .C2(n19443), .A(n19442), .B(n19441), .ZN(
        P2_U3086) );
  AOI22_X1 U22437 ( .A1(n19445), .A2(n19820), .B1(n19819), .B2(n19444), .ZN(
        n19449) );
  AOI22_X1 U22438 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19447), .B1(
        n19446), .B2(n19759), .ZN(n19448) );
  OAI211_X1 U22439 ( .C1(n19764), .C2(n19464), .A(n19449), .B(n19448), .ZN(
        P2_U3087) );
  AOI22_X1 U22440 ( .A1(n19778), .A2(n19490), .B1(n19769), .B2(n19473), .ZN(
        n19459) );
  OAI21_X1 U22441 ( .B1(n19928), .B2(n19684), .A(n19728), .ZN(n19457) );
  INV_X1 U22442 ( .A(n19454), .ZN(n19451) );
  INV_X1 U22443 ( .A(n19473), .ZN(n19450) );
  OAI211_X1 U22444 ( .C1(n19451), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19927), 
        .B(n19450), .ZN(n19452) );
  OAI211_X1 U22445 ( .C1(n19457), .C2(n19453), .A(n19776), .B(n19452), .ZN(
        n19476) );
  OAI21_X1 U22446 ( .B1(n19454), .B2(n19473), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19455) );
  OAI21_X1 U22447 ( .B1(n19457), .B2(n19456), .A(n19455), .ZN(n19475) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19476), .B1(
        n19770), .B2(n19475), .ZN(n19458) );
  OAI211_X1 U22449 ( .C1(n19781), .C2(n19464), .A(n19459), .B(n19458), .ZN(
        P2_U3088) );
  AOI22_X1 U22450 ( .A1(n19784), .A2(n19490), .B1(n19782), .B2(n19473), .ZN(
        n19461) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19476), .B1(
        n19783), .B2(n19475), .ZN(n19460) );
  OAI211_X1 U22452 ( .C1(n19787), .C2(n19464), .A(n19461), .B(n19460), .ZN(
        P2_U3089) );
  AOI22_X1 U22453 ( .A1(n19790), .A2(n19490), .B1(n19788), .B2(n19473), .ZN(
        n19463) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19476), .B1(
        n19789), .B2(n19475), .ZN(n19462) );
  OAI211_X1 U22455 ( .C1(n19793), .C2(n19464), .A(n19463), .B(n19462), .ZN(
        P2_U3090) );
  AOI22_X1 U22456 ( .A1(n19704), .A2(n19474), .B1(n19473), .B2(n19794), .ZN(
        n19466) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19476), .B1(
        n19795), .B2(n19475), .ZN(n19465) );
  OAI211_X1 U22458 ( .C1(n19707), .C2(n19498), .A(n19466), .B(n19465), .ZN(
        P2_U3091) );
  AOI22_X1 U22459 ( .A1(n19708), .A2(n19474), .B1(n19473), .B2(n19800), .ZN(
        n19468) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19476), .B1(
        n19801), .B2(n19475), .ZN(n19467) );
  OAI211_X1 U22461 ( .C1(n19711), .C2(n19498), .A(n19468), .B(n19467), .ZN(
        P2_U3092) );
  AOI22_X1 U22462 ( .A1(n19712), .A2(n19474), .B1(n19473), .B2(n19806), .ZN(
        n19470) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19476), .B1(
        n19807), .B2(n19475), .ZN(n19469) );
  OAI211_X1 U22464 ( .C1(n19715), .C2(n19498), .A(n19470), .B(n19469), .ZN(
        P2_U3093) );
  AOI22_X1 U22465 ( .A1(n19716), .A2(n19474), .B1(n19473), .B2(n19812), .ZN(
        n19472) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19476), .B1(
        n19813), .B2(n19475), .ZN(n19471) );
  OAI211_X1 U22467 ( .C1(n19719), .C2(n19498), .A(n19472), .B(n19471), .ZN(
        P2_U3094) );
  AOI22_X1 U22468 ( .A1(n19759), .A2(n19474), .B1(n19819), .B2(n19473), .ZN(
        n19478) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19476), .B1(
        n19820), .B2(n19475), .ZN(n19477) );
  OAI211_X1 U22470 ( .C1(n19764), .C2(n19498), .A(n19478), .B(n19477), .ZN(
        P2_U3095) );
  AOI22_X1 U22471 ( .A1(n19494), .A2(n19783), .B1(n19493), .B2(n19782), .ZN(
        n19480) );
  AOI22_X1 U22472 ( .A1(n19490), .A2(n19741), .B1(n19523), .B2(n19784), .ZN(
        n19479) );
  OAI211_X1 U22473 ( .C1(n19481), .C2(n14094), .A(n19480), .B(n19479), .ZN(
        P2_U3097) );
  AOI22_X1 U22474 ( .A1(n19494), .A2(n19789), .B1(n19493), .B2(n19788), .ZN(
        n19483) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19495), .B1(
        n19523), .B2(n19790), .ZN(n19482) );
  OAI211_X1 U22476 ( .C1(n19793), .C2(n19498), .A(n19483), .B(n19482), .ZN(
        P2_U3098) );
  AOI22_X1 U22477 ( .A1(n19494), .A2(n19795), .B1(n19493), .B2(n19794), .ZN(
        n19485) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19495), .B1(
        n19523), .B2(n19796), .ZN(n19484) );
  OAI211_X1 U22479 ( .C1(n19799), .C2(n19498), .A(n19485), .B(n19484), .ZN(
        P2_U3099) );
  AOI22_X1 U22480 ( .A1(n19494), .A2(n19801), .B1(n19493), .B2(n19800), .ZN(
        n19487) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19495), .B1(
        n19523), .B2(n19802), .ZN(n19486) );
  OAI211_X1 U22482 ( .C1(n19805), .C2(n19498), .A(n19487), .B(n19486), .ZN(
        P2_U3100) );
  AOI22_X1 U22483 ( .A1(n19494), .A2(n19807), .B1(n19493), .B2(n19806), .ZN(
        n19489) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19495), .B1(
        n19523), .B2(n19808), .ZN(n19488) );
  OAI211_X1 U22485 ( .C1(n19811), .C2(n19498), .A(n19489), .B(n19488), .ZN(
        P2_U3101) );
  AOI22_X1 U22486 ( .A1(n19494), .A2(n19813), .B1(n19493), .B2(n19812), .ZN(
        n19492) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19495), .B1(
        n19490), .B2(n19716), .ZN(n19491) );
  OAI211_X1 U22488 ( .C1(n19719), .C2(n19513), .A(n19492), .B(n19491), .ZN(
        P2_U3102) );
  AOI22_X1 U22489 ( .A1(n19494), .A2(n19820), .B1(n19493), .B2(n19819), .ZN(
        n19497) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19495), .B1(
        n19523), .B2(n19822), .ZN(n19496) );
  OAI211_X1 U22491 ( .C1(n19828), .C2(n19498), .A(n19497), .B(n19496), .ZN(
        P2_U3103) );
  NOR3_X1 U22492 ( .A1(n12192), .A2(n19534), .A3(n19979), .ZN(n19502) );
  AOI211_X2 U22493 ( .C1(n19504), .C2(n19979), .A(n19500), .B(n19502), .ZN(
        n19522) );
  AOI22_X1 U22494 ( .A1(n19522), .A2(n19770), .B1(n19534), .B2(n19769), .ZN(
        n19508) );
  NAND2_X1 U22495 ( .A1(n19501), .A2(n19771), .ZN(n19505) );
  AOI211_X1 U22496 ( .C1(n19505), .C2(n19504), .A(n19503), .B(n19502), .ZN(
        n19506) );
  OAI21_X1 U22497 ( .B1(n19534), .B2(n19971), .A(n19506), .ZN(n19524) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19524), .B1(
        n19523), .B2(n19694), .ZN(n19507) );
  OAI211_X1 U22499 ( .C1(n19697), .C2(n19557), .A(n19508), .B(n19507), .ZN(
        P2_U3104) );
  AOI22_X1 U22500 ( .A1(n19522), .A2(n19783), .B1(n19534), .B2(n19782), .ZN(
        n19510) );
  INV_X1 U22501 ( .A(n19557), .ZN(n19541) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19524), .B1(
        n19541), .B2(n19784), .ZN(n19509) );
  OAI211_X1 U22503 ( .C1(n19787), .C2(n19513), .A(n19510), .B(n19509), .ZN(
        P2_U3105) );
  AOI22_X1 U22504 ( .A1(n19522), .A2(n19789), .B1(n19534), .B2(n19788), .ZN(
        n19512) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19524), .B1(
        n19541), .B2(n19790), .ZN(n19511) );
  OAI211_X1 U22506 ( .C1(n19793), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3106) );
  AOI22_X1 U22507 ( .A1(n19522), .A2(n19795), .B1(n19534), .B2(n19794), .ZN(
        n19515) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19524), .B1(
        n19523), .B2(n19704), .ZN(n19514) );
  OAI211_X1 U22509 ( .C1(n19707), .C2(n19557), .A(n19515), .B(n19514), .ZN(
        P2_U3107) );
  AOI22_X1 U22510 ( .A1(n19522), .A2(n19801), .B1(n19534), .B2(n19800), .ZN(
        n19517) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19524), .B1(
        n19523), .B2(n19708), .ZN(n19516) );
  OAI211_X1 U22512 ( .C1(n19711), .C2(n19557), .A(n19517), .B(n19516), .ZN(
        P2_U3108) );
  AOI22_X1 U22513 ( .A1(n19522), .A2(n19807), .B1(n19534), .B2(n19806), .ZN(
        n19519) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19524), .B1(
        n19523), .B2(n19712), .ZN(n19518) );
  OAI211_X1 U22515 ( .C1(n19715), .C2(n19557), .A(n19519), .B(n19518), .ZN(
        P2_U3109) );
  AOI22_X1 U22516 ( .A1(n19522), .A2(n19813), .B1(n19534), .B2(n19812), .ZN(
        n19521) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19524), .B1(
        n19523), .B2(n19716), .ZN(n19520) );
  OAI211_X1 U22518 ( .C1(n19719), .C2(n19557), .A(n19521), .B(n19520), .ZN(
        P2_U3110) );
  AOI22_X1 U22519 ( .A1(n19522), .A2(n19820), .B1(n19534), .B2(n19819), .ZN(
        n19526) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19524), .B1(
        n19523), .B2(n19759), .ZN(n19525) );
  OAI211_X1 U22521 ( .C1(n19764), .C2(n19557), .A(n19526), .B(n19525), .ZN(
        P2_U3111) );
  NOR2_X1 U22522 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19933), .ZN(
        n19619) );
  NAND2_X1 U22523 ( .A1(n19619), .A2(n19949), .ZN(n19567) );
  NOR2_X1 U22524 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19567), .ZN(
        n19552) );
  AOI22_X1 U22525 ( .A1(n19778), .A2(n19575), .B1(n19769), .B2(n19552), .ZN(
        n19538) );
  NAND2_X1 U22526 ( .A1(n19557), .A2(n19728), .ZN(n19528) );
  OAI21_X1 U22527 ( .B1(n19575), .B2(n19528), .A(n19923), .ZN(n19533) );
  OAI21_X1 U22528 ( .B1(n19529), .B2(n19979), .A(n19971), .ZN(n19530) );
  AOI21_X1 U22529 ( .B1(n19533), .B2(n19531), .A(n19530), .ZN(n19532) );
  OAI21_X1 U22530 ( .B1(n19552), .B2(n19532), .A(n19776), .ZN(n19554) );
  OAI21_X1 U22531 ( .B1(n19534), .B2(n19552), .A(n19533), .ZN(n19536) );
  OAI21_X1 U22532 ( .B1(n19529), .B2(n19552), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19535) );
  NAND2_X1 U22533 ( .A1(n19536), .A2(n19535), .ZN(n19553) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19554), .B1(
        n19770), .B2(n19553), .ZN(n19537) );
  OAI211_X1 U22535 ( .C1(n19781), .C2(n19557), .A(n19538), .B(n19537), .ZN(
        P2_U3112) );
  AOI22_X1 U22536 ( .A1(n19741), .A2(n19541), .B1(n19782), .B2(n19552), .ZN(
        n19540) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19783), .ZN(n19539) );
  OAI211_X1 U22538 ( .C1(n19744), .C2(n19588), .A(n19540), .B(n19539), .ZN(
        P2_U3113) );
  AOI22_X1 U22539 ( .A1(n19700), .A2(n19541), .B1(n19552), .B2(n19788), .ZN(
        n19543) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19789), .ZN(n19542) );
  OAI211_X1 U22541 ( .C1(n19703), .C2(n19588), .A(n19543), .B(n19542), .ZN(
        P2_U3114) );
  AOI22_X1 U22542 ( .A1(n19796), .A2(n19575), .B1(n19552), .B2(n19794), .ZN(
        n19545) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19795), .ZN(n19544) );
  OAI211_X1 U22544 ( .C1(n19799), .C2(n19557), .A(n19545), .B(n19544), .ZN(
        P2_U3115) );
  AOI22_X1 U22545 ( .A1(n19802), .A2(n19575), .B1(n19552), .B2(n19800), .ZN(
        n19547) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19801), .ZN(n19546) );
  OAI211_X1 U22547 ( .C1(n19805), .C2(n19557), .A(n19547), .B(n19546), .ZN(
        P2_U3116) );
  AOI22_X1 U22548 ( .A1(n19808), .A2(n19575), .B1(n19552), .B2(n19806), .ZN(
        n19549) );
  AOI22_X1 U22549 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19807), .ZN(n19548) );
  OAI211_X1 U22550 ( .C1(n19811), .C2(n19557), .A(n19549), .B(n19548), .ZN(
        P2_U3117) );
  AOI22_X1 U22551 ( .A1(n19814), .A2(n19575), .B1(n19552), .B2(n19812), .ZN(
        n19551) );
  AOI22_X1 U22552 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19813), .ZN(n19550) );
  OAI211_X1 U22553 ( .C1(n19817), .C2(n19557), .A(n19551), .B(n19550), .ZN(
        P2_U3118) );
  AOI22_X1 U22554 ( .A1(n19822), .A2(n19575), .B1(n19819), .B2(n19552), .ZN(
        n19556) );
  AOI22_X1 U22555 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19554), .B1(
        n19553), .B2(n19820), .ZN(n19555) );
  OAI211_X1 U22556 ( .C1(n19828), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3119) );
  INV_X1 U22557 ( .A(n19619), .ZN(n19621) );
  NOR2_X1 U22558 ( .A1(n19558), .A2(n19621), .ZN(n19593) );
  AOI22_X1 U22559 ( .A1(n19694), .A2(n19575), .B1(n19769), .B2(n19593), .ZN(
        n19570) );
  INV_X1 U22560 ( .A(n19925), .ZN(n19559) );
  NAND2_X1 U22561 ( .A1(n19559), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19625) );
  OAI21_X1 U22562 ( .B1(n19625), .B2(n19560), .A(n19728), .ZN(n19568) );
  INV_X1 U22563 ( .A(n19567), .ZN(n19563) );
  INV_X1 U22564 ( .A(n19593), .ZN(n19561) );
  OAI211_X1 U22565 ( .C1(n19564), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19927), 
        .B(n19561), .ZN(n19562) );
  OAI211_X1 U22566 ( .C1(n19568), .C2(n19563), .A(n19776), .B(n19562), .ZN(
        n19585) );
  INV_X1 U22567 ( .A(n19564), .ZN(n19565) );
  OAI21_X1 U22568 ( .B1(n19565), .B2(n19593), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19566) );
  OAI21_X1 U22569 ( .B1(n19568), .B2(n19567), .A(n19566), .ZN(n19584) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19585), .B1(
        n19770), .B2(n19584), .ZN(n19569) );
  OAI211_X1 U22571 ( .C1(n19697), .C2(n19618), .A(n19570), .B(n19569), .ZN(
        P2_U3120) );
  AOI22_X1 U22572 ( .A1(n19741), .A2(n19575), .B1(n19782), .B2(n19593), .ZN(
        n19572) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19585), .B1(
        n19783), .B2(n19584), .ZN(n19571) );
  OAI211_X1 U22574 ( .C1(n19744), .C2(n19618), .A(n19572), .B(n19571), .ZN(
        P2_U3121) );
  AOI22_X1 U22575 ( .A1(n19790), .A2(n19602), .B1(n19788), .B2(n19593), .ZN(
        n19574) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19585), .B1(
        n19789), .B2(n19584), .ZN(n19573) );
  OAI211_X1 U22577 ( .C1(n19793), .C2(n19588), .A(n19574), .B(n19573), .ZN(
        P2_U3122) );
  AOI22_X1 U22578 ( .A1(n19704), .A2(n19575), .B1(n19794), .B2(n19593), .ZN(
        n19577) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19585), .B1(
        n19795), .B2(n19584), .ZN(n19576) );
  OAI211_X1 U22580 ( .C1(n19707), .C2(n19618), .A(n19577), .B(n19576), .ZN(
        P2_U3123) );
  AOI22_X1 U22581 ( .A1(n19802), .A2(n19602), .B1(n19800), .B2(n19593), .ZN(
        n19579) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19585), .B1(
        n19801), .B2(n19584), .ZN(n19578) );
  OAI211_X1 U22583 ( .C1(n19805), .C2(n19588), .A(n19579), .B(n19578), .ZN(
        P2_U3124) );
  AOI22_X1 U22584 ( .A1(n19808), .A2(n19602), .B1(n19806), .B2(n19593), .ZN(
        n19581) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19585), .B1(
        n19807), .B2(n19584), .ZN(n19580) );
  OAI211_X1 U22586 ( .C1(n19811), .C2(n19588), .A(n19581), .B(n19580), .ZN(
        P2_U3125) );
  AOI22_X1 U22587 ( .A1(n19814), .A2(n19602), .B1(n19812), .B2(n19593), .ZN(
        n19583) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19585), .B1(
        n19813), .B2(n19584), .ZN(n19582) );
  OAI211_X1 U22589 ( .C1(n19817), .C2(n19588), .A(n19583), .B(n19582), .ZN(
        P2_U3126) );
  AOI22_X1 U22590 ( .A1(n19822), .A2(n19602), .B1(n19819), .B2(n19593), .ZN(
        n19587) );
  AOI22_X1 U22591 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19585), .B1(
        n19820), .B2(n19584), .ZN(n19586) );
  OAI211_X1 U22592 ( .C1(n19828), .C2(n19588), .A(n19587), .B(n19586), .ZN(
        P2_U3127) );
  INV_X1 U22593 ( .A(n19595), .ZN(n19590) );
  AND2_X1 U22594 ( .A1(n19589), .A2(n19619), .ZN(n19613) );
  OAI21_X1 U22595 ( .B1(n19590), .B2(n19613), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19591) );
  OAI21_X1 U22596 ( .B1(n19621), .B2(n19592), .A(n19591), .ZN(n19614) );
  AOI22_X1 U22597 ( .A1(n19614), .A2(n19770), .B1(n19769), .B2(n19613), .ZN(
        n19599) );
  NOR2_X2 U22598 ( .A1(n19725), .A2(n19630), .ZN(n19643) );
  AOI221_X1 U22599 ( .B1(n19602), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19643), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19593), .ZN(n19594) );
  MUX2_X1 U22600 ( .A(n19595), .B(n19594), .S(n19979), .Z(n19596) );
  NOR2_X1 U22601 ( .A1(n19596), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19597) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19615), .B1(
        n19643), .B2(n19778), .ZN(n19598) );
  OAI211_X1 U22603 ( .C1(n19781), .C2(n19618), .A(n19599), .B(n19598), .ZN(
        P2_U3128) );
  INV_X1 U22604 ( .A(n19643), .ZN(n19651) );
  AOI22_X1 U22605 ( .A1(n19614), .A2(n19783), .B1(n19782), .B2(n19613), .ZN(
        n19601) );
  AOI22_X1 U22606 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19615), .B1(
        n19602), .B2(n19741), .ZN(n19600) );
  OAI211_X1 U22607 ( .C1(n19744), .C2(n19651), .A(n19601), .B(n19600), .ZN(
        P2_U3129) );
  AOI22_X1 U22608 ( .A1(n19614), .A2(n19789), .B1(n19788), .B2(n19613), .ZN(
        n19604) );
  AOI22_X1 U22609 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19615), .B1(
        n19602), .B2(n19700), .ZN(n19603) );
  OAI211_X1 U22610 ( .C1(n19703), .C2(n19651), .A(n19604), .B(n19603), .ZN(
        P2_U3130) );
  AOI22_X1 U22611 ( .A1(n19614), .A2(n19795), .B1(n19794), .B2(n19613), .ZN(
        n19606) );
  AOI22_X1 U22612 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19615), .B1(
        n19643), .B2(n19796), .ZN(n19605) );
  OAI211_X1 U22613 ( .C1(n19799), .C2(n19618), .A(n19606), .B(n19605), .ZN(
        P2_U3131) );
  AOI22_X1 U22614 ( .A1(n19614), .A2(n19801), .B1(n19800), .B2(n19613), .ZN(
        n19608) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19615), .B1(
        n19643), .B2(n19802), .ZN(n19607) );
  OAI211_X1 U22616 ( .C1(n19805), .C2(n19618), .A(n19608), .B(n19607), .ZN(
        P2_U3132) );
  AOI22_X1 U22617 ( .A1(n19614), .A2(n19807), .B1(n19806), .B2(n19613), .ZN(
        n19610) );
  AOI22_X1 U22618 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19615), .B1(
        n19643), .B2(n19808), .ZN(n19609) );
  OAI211_X1 U22619 ( .C1(n19811), .C2(n19618), .A(n19610), .B(n19609), .ZN(
        P2_U3133) );
  AOI22_X1 U22620 ( .A1(n19614), .A2(n19813), .B1(n19812), .B2(n19613), .ZN(
        n19612) );
  AOI22_X1 U22621 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19615), .B1(
        n19643), .B2(n19814), .ZN(n19611) );
  OAI211_X1 U22622 ( .C1(n19817), .C2(n19618), .A(n19612), .B(n19611), .ZN(
        P2_U3134) );
  AOI22_X1 U22623 ( .A1(n19614), .A2(n19820), .B1(n19819), .B2(n19613), .ZN(
        n19617) );
  AOI22_X1 U22624 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19615), .B1(
        n19643), .B2(n19822), .ZN(n19616) );
  OAI211_X1 U22625 ( .C1(n19828), .C2(n19618), .A(n19617), .B(n19616), .ZN(
        P2_U3135) );
  NAND2_X1 U22626 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19619), .ZN(
        n19627) );
  OR2_X1 U22627 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19627), .ZN(n19624) );
  INV_X1 U22628 ( .A(n19620), .ZN(n19623) );
  NOR2_X1 U22629 ( .A1(n19622), .A2(n19621), .ZN(n19646) );
  NOR3_X1 U22630 ( .A1(n19623), .A2(n19646), .A3(n19979), .ZN(n19626) );
  AOI21_X1 U22631 ( .B1(n19979), .B2(n19624), .A(n19626), .ZN(n19647) );
  AOI22_X1 U22632 ( .A1(n19647), .A2(n19770), .B1(n19769), .B2(n19646), .ZN(
        n19632) );
  INV_X1 U22633 ( .A(n19625), .ZN(n19772) );
  INV_X1 U22634 ( .A(n19630), .ZN(n19921) );
  NAND2_X1 U22635 ( .A1(n19772), .A2(n19921), .ZN(n19628) );
  AOI21_X1 U22636 ( .B1(n19628), .B2(n19627), .A(n19626), .ZN(n19629) );
  OAI211_X1 U22637 ( .C1(n19646), .C2(n19971), .A(n19629), .B(n19776), .ZN(
        n19648) );
  AOI22_X1 U22638 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19648), .B1(
        n19656), .B2(n19778), .ZN(n19631) );
  OAI211_X1 U22639 ( .C1(n19781), .C2(n19651), .A(n19632), .B(n19631), .ZN(
        P2_U3136) );
  AOI22_X1 U22640 ( .A1(n19647), .A2(n19783), .B1(n19782), .B2(n19646), .ZN(
        n19634) );
  AOI22_X1 U22641 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19648), .B1(
        n19643), .B2(n19741), .ZN(n19633) );
  OAI211_X1 U22642 ( .C1(n19744), .C2(n19682), .A(n19634), .B(n19633), .ZN(
        P2_U3137) );
  AOI22_X1 U22643 ( .A1(n19647), .A2(n19789), .B1(n19788), .B2(n19646), .ZN(
        n19636) );
  AOI22_X1 U22644 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19648), .B1(
        n19643), .B2(n19700), .ZN(n19635) );
  OAI211_X1 U22645 ( .C1(n19703), .C2(n19682), .A(n19636), .B(n19635), .ZN(
        P2_U3138) );
  AOI22_X1 U22646 ( .A1(n19647), .A2(n19795), .B1(n19794), .B2(n19646), .ZN(
        n19638) );
  AOI22_X1 U22647 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19648), .B1(
        n19643), .B2(n19704), .ZN(n19637) );
  OAI211_X1 U22648 ( .C1(n19707), .C2(n19682), .A(n19638), .B(n19637), .ZN(
        P2_U3139) );
  AOI22_X1 U22649 ( .A1(n19647), .A2(n19801), .B1(n19800), .B2(n19646), .ZN(
        n19640) );
  AOI22_X1 U22650 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19648), .B1(
        n19643), .B2(n19708), .ZN(n19639) );
  OAI211_X1 U22651 ( .C1(n19711), .C2(n19682), .A(n19640), .B(n19639), .ZN(
        P2_U3140) );
  AOI22_X1 U22652 ( .A1(n19647), .A2(n19807), .B1(n19806), .B2(n19646), .ZN(
        n19642) );
  AOI22_X1 U22653 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19648), .B1(
        n19643), .B2(n19712), .ZN(n19641) );
  OAI211_X1 U22654 ( .C1(n19715), .C2(n19682), .A(n19642), .B(n19641), .ZN(
        P2_U3141) );
  AOI22_X1 U22655 ( .A1(n19647), .A2(n19813), .B1(n19812), .B2(n19646), .ZN(
        n19645) );
  AOI22_X1 U22656 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19648), .B1(
        n19643), .B2(n19716), .ZN(n19644) );
  OAI211_X1 U22657 ( .C1(n19719), .C2(n19682), .A(n19645), .B(n19644), .ZN(
        P2_U3142) );
  AOI22_X1 U22658 ( .A1(n19647), .A2(n19820), .B1(n19819), .B2(n19646), .ZN(
        n19650) );
  AOI22_X1 U22659 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19648), .B1(
        n19656), .B2(n19822), .ZN(n19649) );
  OAI211_X1 U22660 ( .C1(n19828), .C2(n19651), .A(n19650), .B(n19649), .ZN(
        P2_U3143) );
  INV_X1 U22661 ( .A(n19652), .ZN(n19655) );
  NAND3_X1 U22662 ( .A1(n19949), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19691) );
  NOR2_X1 U22663 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19691), .ZN(
        n19677) );
  OAI21_X1 U22664 ( .B1(n19653), .B2(n19677), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19654) );
  OAI21_X1 U22665 ( .B1(n19655), .B2(n19658), .A(n19654), .ZN(n19678) );
  AOI22_X1 U22666 ( .A1(n19678), .A2(n19770), .B1(n19769), .B2(n19677), .ZN(
        n19664) );
  NOR2_X2 U22667 ( .A1(n19725), .A2(n19684), .ZN(n19721) );
  OAI21_X1 U22668 ( .B1(n19656), .B2(n19721), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19657) );
  OAI21_X1 U22669 ( .B1(n19658), .B2(n19933), .A(n19657), .ZN(n19662) );
  INV_X1 U22670 ( .A(n19677), .ZN(n19659) );
  OAI211_X1 U22671 ( .C1(n19660), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19927), 
        .B(n19659), .ZN(n19661) );
  NAND3_X1 U22672 ( .A1(n19662), .A2(n19776), .A3(n19661), .ZN(n19679) );
  AOI22_X1 U22673 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19778), .ZN(n19663) );
  OAI211_X1 U22674 ( .C1(n19781), .C2(n19682), .A(n19664), .B(n19663), .ZN(
        P2_U3144) );
  AOI22_X1 U22675 ( .A1(n19678), .A2(n19783), .B1(n19782), .B2(n19677), .ZN(
        n19666) );
  AOI22_X1 U22676 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19784), .ZN(n19665) );
  OAI211_X1 U22677 ( .C1(n19787), .C2(n19682), .A(n19666), .B(n19665), .ZN(
        P2_U3145) );
  AOI22_X1 U22678 ( .A1(n19678), .A2(n19789), .B1(n19788), .B2(n19677), .ZN(
        n19668) );
  AOI22_X1 U22679 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19790), .ZN(n19667) );
  OAI211_X1 U22680 ( .C1(n19793), .C2(n19682), .A(n19668), .B(n19667), .ZN(
        P2_U3146) );
  AOI22_X1 U22681 ( .A1(n19678), .A2(n19795), .B1(n19794), .B2(n19677), .ZN(
        n19670) );
  AOI22_X1 U22682 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19796), .ZN(n19669) );
  OAI211_X1 U22683 ( .C1(n19799), .C2(n19682), .A(n19670), .B(n19669), .ZN(
        P2_U3147) );
  AOI22_X1 U22684 ( .A1(n19678), .A2(n19801), .B1(n19800), .B2(n19677), .ZN(
        n19672) );
  AOI22_X1 U22685 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19802), .ZN(n19671) );
  OAI211_X1 U22686 ( .C1(n19805), .C2(n19682), .A(n19672), .B(n19671), .ZN(
        P2_U3148) );
  AOI22_X1 U22687 ( .A1(n19678), .A2(n19807), .B1(n19806), .B2(n19677), .ZN(
        n19674) );
  AOI22_X1 U22688 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19808), .ZN(n19673) );
  OAI211_X1 U22689 ( .C1(n19811), .C2(n19682), .A(n19674), .B(n19673), .ZN(
        P2_U3149) );
  AOI22_X1 U22690 ( .A1(n19678), .A2(n19813), .B1(n19812), .B2(n19677), .ZN(
        n19676) );
  AOI22_X1 U22691 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19814), .ZN(n19675) );
  OAI211_X1 U22692 ( .C1(n19817), .C2(n19682), .A(n19676), .B(n19675), .ZN(
        P2_U3150) );
  AOI22_X1 U22693 ( .A1(n19678), .A2(n19820), .B1(n19819), .B2(n19677), .ZN(
        n19681) );
  AOI22_X1 U22694 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19679), .B1(
        n19721), .B2(n19822), .ZN(n19680) );
  OAI211_X1 U22695 ( .C1(n19828), .C2(n19682), .A(n19681), .B(n19680), .ZN(
        P2_U3151) );
  INV_X1 U22696 ( .A(n19683), .ZN(n19685) );
  INV_X1 U22697 ( .A(n19684), .ZN(n19689) );
  NOR2_X1 U22698 ( .A1(n19958), .A2(n19691), .ZN(n19730) );
  NOR3_X1 U22699 ( .A1(n19686), .A2(n19730), .A3(n19979), .ZN(n19690) );
  INV_X1 U22700 ( .A(n19691), .ZN(n19687) );
  AOI21_X1 U22701 ( .B1(n19971), .B2(n19687), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19688) );
  NOR2_X1 U22702 ( .A1(n19690), .A2(n19688), .ZN(n19720) );
  AOI22_X1 U22703 ( .A1(n19720), .A2(n19770), .B1(n19769), .B2(n19730), .ZN(
        n19696) );
  NAND2_X1 U22704 ( .A1(n19772), .A2(n19689), .ZN(n19692) );
  AOI21_X1 U22705 ( .B1(n19692), .B2(n19691), .A(n19690), .ZN(n19693) );
  OAI211_X1 U22706 ( .C1(n19730), .C2(n19971), .A(n19693), .B(n19776), .ZN(
        n19722) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19694), .ZN(n19695) );
  OAI211_X1 U22708 ( .C1(n19697), .C2(n19756), .A(n19696), .B(n19695), .ZN(
        P2_U3152) );
  AOI22_X1 U22709 ( .A1(n19720), .A2(n19783), .B1(n19782), .B2(n19730), .ZN(
        n19699) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19741), .ZN(n19698) );
  OAI211_X1 U22711 ( .C1(n19744), .C2(n19756), .A(n19699), .B(n19698), .ZN(
        P2_U3153) );
  AOI22_X1 U22712 ( .A1(n19720), .A2(n19789), .B1(n19788), .B2(n19730), .ZN(
        n19702) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19700), .ZN(n19701) );
  OAI211_X1 U22714 ( .C1(n19703), .C2(n19756), .A(n19702), .B(n19701), .ZN(
        P2_U3154) );
  AOI22_X1 U22715 ( .A1(n19720), .A2(n19795), .B1(n19794), .B2(n19730), .ZN(
        n19706) );
  AOI22_X1 U22716 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19704), .ZN(n19705) );
  OAI211_X1 U22717 ( .C1(n19707), .C2(n19756), .A(n19706), .B(n19705), .ZN(
        P2_U3155) );
  AOI22_X1 U22718 ( .A1(n19720), .A2(n19801), .B1(n19800), .B2(n19730), .ZN(
        n19710) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19708), .ZN(n19709) );
  OAI211_X1 U22720 ( .C1(n19711), .C2(n19756), .A(n19710), .B(n19709), .ZN(
        P2_U3156) );
  AOI22_X1 U22721 ( .A1(n19720), .A2(n19807), .B1(n19806), .B2(n19730), .ZN(
        n19714) );
  AOI22_X1 U22722 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19712), .ZN(n19713) );
  OAI211_X1 U22723 ( .C1(n19715), .C2(n19756), .A(n19714), .B(n19713), .ZN(
        P2_U3157) );
  AOI22_X1 U22724 ( .A1(n19720), .A2(n19813), .B1(n19812), .B2(n19730), .ZN(
        n19718) );
  AOI22_X1 U22725 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19716), .ZN(n19717) );
  OAI211_X1 U22726 ( .C1(n19719), .C2(n19756), .A(n19718), .B(n19717), .ZN(
        P2_U3158) );
  AOI22_X1 U22727 ( .A1(n19720), .A2(n19820), .B1(n19819), .B2(n19730), .ZN(
        n19724) );
  AOI22_X1 U22728 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19722), .B1(
        n19721), .B2(n19759), .ZN(n19723) );
  OAI211_X1 U22729 ( .C1(n19764), .C2(n19756), .A(n19724), .B(n19723), .ZN(
        P2_U3159) );
  INV_X1 U22730 ( .A(n19725), .ZN(n19726) );
  NAND2_X1 U22731 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19727), .ZN(
        n19774) );
  NOR2_X1 U22732 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19774), .ZN(
        n19757) );
  AOI22_X1 U22733 ( .A1(n19778), .A2(n19753), .B1(n19769), .B2(n19757), .ZN(
        n19740) );
  NOR2_X1 U22734 ( .A1(n19758), .A2(n19753), .ZN(n19729) );
  OAI21_X1 U22735 ( .B1(n19729), .B2(n19920), .A(n19728), .ZN(n19738) );
  NOR2_X1 U22736 ( .A1(n19757), .A2(n19730), .ZN(n19737) );
  INV_X1 U22737 ( .A(n19737), .ZN(n19733) );
  INV_X1 U22738 ( .A(n19757), .ZN(n19731) );
  OAI211_X1 U22739 ( .C1(n19734), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19927), 
        .B(n19731), .ZN(n19732) );
  OAI211_X1 U22740 ( .C1(n19738), .C2(n19733), .A(n19776), .B(n19732), .ZN(
        n19761) );
  INV_X1 U22741 ( .A(n19734), .ZN(n19735) );
  OAI21_X1 U22742 ( .B1(n19735), .B2(n19757), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19736) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19761), .B1(
        n19770), .B2(n19760), .ZN(n19739) );
  OAI211_X1 U22744 ( .C1(n19781), .C2(n19756), .A(n19740), .B(n19739), .ZN(
        P2_U3160) );
  AOI22_X1 U22745 ( .A1(n19741), .A2(n19758), .B1(n19782), .B2(n19757), .ZN(
        n19743) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19761), .B1(
        n19783), .B2(n19760), .ZN(n19742) );
  OAI211_X1 U22747 ( .C1(n19744), .C2(n19827), .A(n19743), .B(n19742), .ZN(
        P2_U3161) );
  AOI22_X1 U22748 ( .A1(n19790), .A2(n19753), .B1(n19788), .B2(n19757), .ZN(
        n19746) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19761), .B1(
        n19789), .B2(n19760), .ZN(n19745) );
  OAI211_X1 U22750 ( .C1(n19793), .C2(n19756), .A(n19746), .B(n19745), .ZN(
        P2_U3162) );
  AOI22_X1 U22751 ( .A1(n19796), .A2(n19753), .B1(n19794), .B2(n19757), .ZN(
        n19748) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19761), .B1(
        n19795), .B2(n19760), .ZN(n19747) );
  OAI211_X1 U22753 ( .C1(n19799), .C2(n19756), .A(n19748), .B(n19747), .ZN(
        P2_U3163) );
  AOI22_X1 U22754 ( .A1(n19802), .A2(n19753), .B1(n19800), .B2(n19757), .ZN(
        n19750) );
  AOI22_X1 U22755 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19761), .B1(
        n19801), .B2(n19760), .ZN(n19749) );
  OAI211_X1 U22756 ( .C1(n19805), .C2(n19756), .A(n19750), .B(n19749), .ZN(
        P2_U3164) );
  AOI22_X1 U22757 ( .A1(n19808), .A2(n19753), .B1(n19806), .B2(n19757), .ZN(
        n19752) );
  AOI22_X1 U22758 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19761), .B1(
        n19807), .B2(n19760), .ZN(n19751) );
  OAI211_X1 U22759 ( .C1(n19811), .C2(n19756), .A(n19752), .B(n19751), .ZN(
        P2_U3165) );
  AOI22_X1 U22760 ( .A1(n19814), .A2(n19753), .B1(n19812), .B2(n19757), .ZN(
        n19755) );
  AOI22_X1 U22761 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19761), .B1(
        n19813), .B2(n19760), .ZN(n19754) );
  OAI211_X1 U22762 ( .C1(n19817), .C2(n19756), .A(n19755), .B(n19754), .ZN(
        P2_U3166) );
  AOI22_X1 U22763 ( .A1(n19759), .A2(n19758), .B1(n19819), .B2(n19757), .ZN(
        n19763) );
  AOI22_X1 U22764 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19761), .B1(
        n19820), .B2(n19760), .ZN(n19762) );
  OAI211_X1 U22765 ( .C1(n19764), .C2(n19827), .A(n19763), .B(n19762), .ZN(
        P2_U3167) );
  INV_X1 U22766 ( .A(n19765), .ZN(n19766) );
  NOR3_X1 U22767 ( .A1(n19766), .A2(n19818), .A3(n19979), .ZN(n19773) );
  INV_X1 U22768 ( .A(n19774), .ZN(n19767) );
  AOI21_X1 U22769 ( .B1(n19971), .B2(n19767), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19768) );
  NOR2_X1 U22770 ( .A1(n19773), .A2(n19768), .ZN(n19821) );
  AOI22_X1 U22771 ( .A1(n19821), .A2(n19770), .B1(n19769), .B2(n19818), .ZN(
        n19780) );
  NAND2_X1 U22772 ( .A1(n19772), .A2(n19771), .ZN(n19775) );
  AOI21_X1 U22773 ( .B1(n19775), .B2(n19774), .A(n19773), .ZN(n19777) );
  OAI211_X1 U22774 ( .C1(n19818), .C2(n19971), .A(n19777), .B(n19776), .ZN(
        n19824) );
  AOI22_X1 U22775 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19778), .ZN(n19779) );
  OAI211_X1 U22776 ( .C1(n19781), .C2(n19827), .A(n19780), .B(n19779), .ZN(
        P2_U3168) );
  AOI22_X1 U22777 ( .A1(n19821), .A2(n19783), .B1(n19782), .B2(n19818), .ZN(
        n19786) );
  AOI22_X1 U22778 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19784), .ZN(n19785) );
  OAI211_X1 U22779 ( .C1(n19787), .C2(n19827), .A(n19786), .B(n19785), .ZN(
        P2_U3169) );
  AOI22_X1 U22780 ( .A1(n19821), .A2(n19789), .B1(n19788), .B2(n19818), .ZN(
        n19792) );
  AOI22_X1 U22781 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19790), .ZN(n19791) );
  OAI211_X1 U22782 ( .C1(n19793), .C2(n19827), .A(n19792), .B(n19791), .ZN(
        P2_U3170) );
  AOI22_X1 U22783 ( .A1(n19821), .A2(n19795), .B1(n19794), .B2(n19818), .ZN(
        n19798) );
  AOI22_X1 U22784 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19796), .ZN(n19797) );
  OAI211_X1 U22785 ( .C1(n19799), .C2(n19827), .A(n19798), .B(n19797), .ZN(
        P2_U3171) );
  AOI22_X1 U22786 ( .A1(n19821), .A2(n19801), .B1(n19800), .B2(n19818), .ZN(
        n19804) );
  AOI22_X1 U22787 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19802), .ZN(n19803) );
  OAI211_X1 U22788 ( .C1(n19805), .C2(n19827), .A(n19804), .B(n19803), .ZN(
        P2_U3172) );
  AOI22_X1 U22789 ( .A1(n19821), .A2(n19807), .B1(n19806), .B2(n19818), .ZN(
        n19810) );
  AOI22_X1 U22790 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19808), .ZN(n19809) );
  OAI211_X1 U22791 ( .C1(n19811), .C2(n19827), .A(n19810), .B(n19809), .ZN(
        P2_U3173) );
  AOI22_X1 U22792 ( .A1(n19821), .A2(n19813), .B1(n19812), .B2(n19818), .ZN(
        n19816) );
  AOI22_X1 U22793 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19814), .ZN(n19815) );
  OAI211_X1 U22794 ( .C1(n19817), .C2(n19827), .A(n19816), .B(n19815), .ZN(
        P2_U3174) );
  AOI22_X1 U22795 ( .A1(n19821), .A2(n19820), .B1(n19819), .B2(n19818), .ZN(
        n19826) );
  AOI22_X1 U22796 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19824), .B1(
        n19823), .B2(n19822), .ZN(n19825) );
  OAI211_X1 U22797 ( .C1(n19828), .C2(n19827), .A(n19826), .B(n19825), .ZN(
        P2_U3175) );
  AOI21_X1 U22798 ( .B1(n19831), .B2(n19830), .A(n19829), .ZN(n19835) );
  OAI211_X1 U22799 ( .C1(n19836), .C2(n19832), .A(n19980), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19833) );
  OAI211_X1 U22800 ( .C1(n19836), .C2(n19835), .A(n19834), .B(n19833), .ZN(
        P2_U3177) );
  AND2_X1 U22801 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19837), .ZN(
        P2_U3179) );
  AND2_X1 U22802 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19837), .ZN(
        P2_U3180) );
  AND2_X1 U22803 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19837), .ZN(
        P2_U3181) );
  AND2_X1 U22804 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19837), .ZN(
        P2_U3182) );
  AND2_X1 U22805 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19837), .ZN(
        P2_U3183) );
  AND2_X1 U22806 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19837), .ZN(
        P2_U3184) );
  AND2_X1 U22807 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19837), .ZN(
        P2_U3185) );
  AND2_X1 U22808 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19837), .ZN(
        P2_U3186) );
  AND2_X1 U22809 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19837), .ZN(
        P2_U3187) );
  AND2_X1 U22810 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19837), .ZN(
        P2_U3188) );
  AND2_X1 U22811 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19837), .ZN(
        P2_U3189) );
  AND2_X1 U22812 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19837), .ZN(
        P2_U3190) );
  AND2_X1 U22813 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19837), .ZN(
        P2_U3191) );
  AND2_X1 U22814 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19837), .ZN(
        P2_U3192) );
  AND2_X1 U22815 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19837), .ZN(
        P2_U3193) );
  AND2_X1 U22816 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19837), .ZN(
        P2_U3194) );
  AND2_X1 U22817 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19837), .ZN(
        P2_U3195) );
  AND2_X1 U22818 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19837), .ZN(
        P2_U3196) );
  AND2_X1 U22819 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19837), .ZN(
        P2_U3197) );
  AND2_X1 U22820 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19837), .ZN(
        P2_U3198) );
  AND2_X1 U22821 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19837), .ZN(
        P2_U3199) );
  AND2_X1 U22822 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19837), .ZN(
        P2_U3200) );
  AND2_X1 U22823 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19837), .ZN(P2_U3201) );
  AND2_X1 U22824 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19837), .ZN(P2_U3202) );
  AND2_X1 U22825 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19837), .ZN(P2_U3203) );
  AND2_X1 U22826 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19837), .ZN(P2_U3204) );
  AND2_X1 U22827 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19837), .ZN(P2_U3205) );
  AND2_X1 U22828 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19837), .ZN(P2_U3206) );
  AND2_X1 U22829 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19837), .ZN(P2_U3207) );
  AND2_X1 U22830 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19837), .ZN(P2_U3208) );
  INV_X1 U22831 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19848) );
  NOR2_X1 U22832 ( .A1(n19848), .A2(n19838), .ZN(n19846) );
  INV_X1 U22833 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19988) );
  OR3_X1 U22834 ( .A1(n19846), .A2(n19988), .A3(n19839), .ZN(n19841) );
  AOI211_X1 U22835 ( .C1(n20724), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19847), .B(n19892), .ZN(n19840) );
  NOR3_X1 U22836 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .A3(n21174), .ZN(n19852) );
  AOI211_X1 U22837 ( .C1(n19855), .C2(n19841), .A(n19840), .B(n19852), .ZN(
        n19842) );
  INV_X1 U22838 ( .A(n19842), .ZN(P2_U3209) );
  AOI21_X1 U22839 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20724), .A(n19855), 
        .ZN(n19849) );
  NOR3_X1 U22840 ( .A1(n19849), .A2(n19988), .A3(n19839), .ZN(n19843) );
  NOR2_X1 U22841 ( .A1(n19843), .A2(n19846), .ZN(n19844) );
  INV_X1 U22842 ( .A(n19977), .ZN(n19978) );
  OAI211_X1 U22843 ( .C1(n20724), .C2(n19845), .A(n19844), .B(n19978), .ZN(
        P2_U3210) );
  AOI22_X1 U22844 ( .A1(n19847), .A2(n19988), .B1(n19846), .B2(n21174), .ZN(
        n19854) );
  OAI21_X1 U22845 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19853) );
  NOR2_X1 U22846 ( .A1(n19848), .A2(n19855), .ZN(n19850) );
  AOI21_X1 U22847 ( .B1(n19980), .B2(n19850), .A(n19849), .ZN(n19851) );
  OAI22_X1 U22848 ( .A1(n19854), .A2(n19853), .B1(n19852), .B2(n19851), .ZN(
        P2_U3211) );
  NAND2_X1 U22849 ( .A1(n19892), .A2(n19855), .ZN(n19901) );
  CLKBUF_X1 U22850 ( .A(n19901), .Z(n19898) );
  OAI222_X1 U22851 ( .A1(n19898), .A2(n12075), .B1(n19856), .B2(n19892), .C1(
        n12061), .C2(n19899), .ZN(P2_U3212) );
  OAI222_X1 U22852 ( .A1(n19901), .A2(n13425), .B1(n19857), .B2(n19892), .C1(
        n12075), .C2(n19899), .ZN(P2_U3213) );
  OAI222_X1 U22853 ( .A1(n19901), .A2(n12621), .B1(n19858), .B2(n19892), .C1(
        n13425), .C2(n19899), .ZN(P2_U3214) );
  OAI222_X1 U22854 ( .A1(n19901), .A2(n15291), .B1(n19859), .B2(n19892), .C1(
        n12621), .C2(n19899), .ZN(P2_U3215) );
  OAI222_X1 U22855 ( .A1(n19901), .A2(n12495), .B1(n19860), .B2(n19892), .C1(
        n15291), .C2(n19899), .ZN(P2_U3216) );
  OAI222_X1 U22856 ( .A1(n19901), .A2(n19862), .B1(n19861), .B2(n19892), .C1(
        n12495), .C2(n19899), .ZN(P2_U3217) );
  OAI222_X1 U22857 ( .A1(n19898), .A2(n12644), .B1(n19863), .B2(n19892), .C1(
        n19862), .C2(n19899), .ZN(P2_U3218) );
  INV_X1 U22858 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19865) );
  OAI222_X1 U22859 ( .A1(n19898), .A2(n19865), .B1(n19864), .B2(n19892), .C1(
        n12644), .C2(n19899), .ZN(P2_U3219) );
  OAI222_X1 U22860 ( .A1(n19898), .A2(n12671), .B1(n19866), .B2(n19892), .C1(
        n19865), .C2(n19899), .ZN(P2_U3220) );
  OAI222_X1 U22861 ( .A1(n19898), .A2(n12685), .B1(n19867), .B2(n19892), .C1(
        n12671), .C2(n19899), .ZN(P2_U3221) );
  OAI222_X1 U22862 ( .A1(n19898), .A2(n12698), .B1(n19868), .B2(n19892), .C1(
        n12685), .C2(n19899), .ZN(P2_U3222) );
  OAI222_X1 U22863 ( .A1(n19898), .A2(n12712), .B1(n19869), .B2(n19892), .C1(
        n12698), .C2(n19899), .ZN(P2_U3223) );
  OAI222_X1 U22864 ( .A1(n19901), .A2(n12725), .B1(n19870), .B2(n19892), .C1(
        n12712), .C2(n19899), .ZN(P2_U3224) );
  OAI222_X1 U22865 ( .A1(n19901), .A2(n12739), .B1(n19871), .B2(n19892), .C1(
        n12725), .C2(n19899), .ZN(P2_U3225) );
  OAI222_X1 U22866 ( .A1(n19901), .A2(n19873), .B1(n19872), .B2(n19892), .C1(
        n12739), .C2(n19899), .ZN(P2_U3226) );
  OAI222_X1 U22867 ( .A1(n19901), .A2(n19875), .B1(n19874), .B2(n19892), .C1(
        n19873), .C2(n19899), .ZN(P2_U3227) );
  OAI222_X1 U22868 ( .A1(n19901), .A2(n15010), .B1(n19876), .B2(n19892), .C1(
        n19875), .C2(n19899), .ZN(P2_U3228) );
  OAI222_X1 U22869 ( .A1(n19901), .A2(n19878), .B1(n19877), .B2(n19892), .C1(
        n15010), .C2(n19899), .ZN(P2_U3229) );
  OAI222_X1 U22870 ( .A1(n19898), .A2(n19880), .B1(n19879), .B2(n19892), .C1(
        n19878), .C2(n19899), .ZN(P2_U3230) );
  OAI222_X1 U22871 ( .A1(n19898), .A2(n19882), .B1(n19881), .B2(n19892), .C1(
        n19880), .C2(n19899), .ZN(P2_U3231) );
  OAI222_X1 U22872 ( .A1(n19898), .A2(n12750), .B1(n19883), .B2(n19892), .C1(
        n19882), .C2(n19899), .ZN(P2_U3232) );
  OAI222_X1 U22873 ( .A1(n19898), .A2(n19885), .B1(n19884), .B2(n19892), .C1(
        n12750), .C2(n19899), .ZN(P2_U3233) );
  OAI222_X1 U22874 ( .A1(n19898), .A2(n12755), .B1(n19886), .B2(n19892), .C1(
        n19885), .C2(n19899), .ZN(P2_U3234) );
  OAI222_X1 U22875 ( .A1(n19898), .A2(n19888), .B1(n19887), .B2(n19892), .C1(
        n12755), .C2(n19899), .ZN(P2_U3235) );
  OAI222_X1 U22876 ( .A1(n19898), .A2(n19890), .B1(n19889), .B2(n19892), .C1(
        n19888), .C2(n19899), .ZN(P2_U3236) );
  OAI222_X1 U22877 ( .A1(n19898), .A2(n19894), .B1(n19891), .B2(n19892), .C1(
        n19890), .C2(n19899), .ZN(P2_U3237) );
  OAI222_X1 U22878 ( .A1(n19899), .A2(n19894), .B1(n19893), .B2(n19892), .C1(
        n12764), .C2(n19898), .ZN(P2_U3238) );
  OAI222_X1 U22879 ( .A1(n19898), .A2(n19896), .B1(n19895), .B2(n19892), .C1(
        n12764), .C2(n19899), .ZN(P2_U3239) );
  OAI222_X1 U22880 ( .A1(n19898), .A2(n13879), .B1(n19897), .B2(n19892), .C1(
        n19896), .C2(n19899), .ZN(P2_U3240) );
  INV_X1 U22881 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19900) );
  OAI222_X1 U22882 ( .A1(n19901), .A2(n15958), .B1(n19900), .B2(n19892), .C1(
        n13879), .C2(n19899), .ZN(P2_U3241) );
  INV_X1 U22883 ( .A(P2_BE_N_REG_3__SCAN_IN), .ZN(n19902) );
  AOI22_X1 U22884 ( .A1(n19892), .A2(n19903), .B1(n19902), .B2(n19990), .ZN(
        P2_U3585) );
  MUX2_X1 U22885 ( .A(P2_BE_N_REG_2__SCAN_IN), .B(P2_BYTEENABLE_REG_2__SCAN_IN), .S(n19892), .Z(P2_U3586) );
  INV_X1 U22886 ( .A(P2_BE_N_REG_1__SCAN_IN), .ZN(n19904) );
  AOI22_X1 U22887 ( .A1(n19892), .A2(n19905), .B1(n19904), .B2(n19990), .ZN(
        P2_U3587) );
  INV_X1 U22888 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n19906) );
  AOI22_X1 U22889 ( .A1(n19892), .A2(n19907), .B1(n19906), .B2(n19990), .ZN(
        P2_U3588) );
  OAI21_X1 U22890 ( .B1(n19911), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19909), 
        .ZN(n19908) );
  INV_X1 U22891 ( .A(n19908), .ZN(P2_U3591) );
  OAI21_X1 U22892 ( .B1(n19911), .B2(n19910), .A(n19909), .ZN(P2_U3592) );
  INV_X1 U22893 ( .A(n19912), .ZN(n19913) );
  OAI222_X1 U22894 ( .A1(n19917), .A2(n19916), .B1(n19922), .B2(n19915), .C1(
        n19914), .C2(n19913), .ZN(n19919) );
  MUX2_X1 U22895 ( .A(n19919), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n19918), .Z(P2_U3599) );
  NOR2_X1 U22896 ( .A1(n19927), .A2(n19920), .ZN(n19945) );
  NAND2_X1 U22897 ( .A1(n19921), .A2(n19945), .ZN(n19936) );
  OR2_X1 U22898 ( .A1(n19943), .A2(n19927), .ZN(n19924) );
  AND2_X1 U22899 ( .A1(n19923), .A2(n19922), .ZN(n19942) );
  AND2_X1 U22900 ( .A1(n19924), .A2(n19942), .ZN(n19934) );
  AOI21_X1 U22901 ( .B1(n19936), .B2(n19934), .A(n19925), .ZN(n19930) );
  NOR3_X1 U22902 ( .A1(n19928), .A2(n19927), .A3(n19926), .ZN(n19929) );
  AOI211_X1 U22903 ( .C1(n19931), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19930), 
        .B(n19929), .ZN(n19932) );
  AOI22_X1 U22904 ( .A1(n19959), .A2(n19933), .B1(n19932), .B2(n19956), .ZN(
        P2_U3602) );
  INV_X1 U22905 ( .A(n19934), .ZN(n19939) );
  NOR2_X1 U22906 ( .A1(n19935), .A2(n19971), .ZN(n19938) );
  INV_X1 U22907 ( .A(n19936), .ZN(n19937) );
  AOI211_X1 U22908 ( .C1(n19940), .C2(n19939), .A(n19938), .B(n19937), .ZN(
        n19941) );
  AOI22_X1 U22909 ( .A1(n19959), .A2(n13030), .B1(n19941), .B2(n19956), .ZN(
        P2_U3603) );
  INV_X1 U22910 ( .A(n19942), .ZN(n19944) );
  MUX2_X1 U22911 ( .A(n19945), .B(n19944), .S(n19943), .Z(n19946) );
  AOI21_X1 U22912 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19947), .A(n19946), 
        .ZN(n19948) );
  AOI22_X1 U22913 ( .A1(n19959), .A2(n19949), .B1(n19948), .B2(n19956), .ZN(
        P2_U3604) );
  INV_X1 U22914 ( .A(n19950), .ZN(n19951) );
  OAI22_X1 U22915 ( .A1(n19952), .A2(n19951), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19971), .ZN(n19953) );
  AOI21_X1 U22916 ( .B1(n19955), .B2(n19954), .A(n19953), .ZN(n19957) );
  AOI22_X1 U22917 ( .A1(n19959), .A2(n19958), .B1(n19957), .B2(n19956), .ZN(
        P2_U3605) );
  INV_X1 U22918 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19960) );
  AOI22_X1 U22919 ( .A1(n19892), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19960), 
        .B2(n19990), .ZN(P2_U3608) );
  INV_X1 U22920 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19970) );
  INV_X1 U22921 ( .A(n19961), .ZN(n19969) );
  AOI22_X1 U22922 ( .A1(n19965), .A2(n19964), .B1(n19963), .B2(n19962), .ZN(
        n19968) );
  NOR2_X1 U22923 ( .A1(n19969), .A2(n19966), .ZN(n19967) );
  AOI22_X1 U22924 ( .A1(n19970), .A2(n19969), .B1(n19968), .B2(n19967), .ZN(
        P2_U3609) );
  OAI21_X1 U22925 ( .B1(n19972), .B2(n19979), .A(n19971), .ZN(n19973) );
  OAI211_X1 U22926 ( .C1(n19980), .C2(n19975), .A(n19974), .B(n19973), .ZN(
        n19989) );
  AOI211_X1 U22927 ( .C1(P2_STATEBS16_REG_SCAN_IN), .C2(n19977), .A(n19976), 
        .B(n12376), .ZN(n19986) );
  NAND2_X1 U22928 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19978), .ZN(n19983) );
  NOR2_X1 U22929 ( .A1(n19980), .A2(n19979), .ZN(n19981) );
  OAI22_X1 U22930 ( .A1(n19984), .A2(n19983), .B1(n19982), .B2(n19981), .ZN(
        n19985) );
  OAI21_X1 U22931 ( .B1(n19986), .B2(n19985), .A(n19989), .ZN(n19987) );
  OAI21_X1 U22932 ( .B1(n19989), .B2(n19988), .A(n19987), .ZN(P2_U3610) );
  OAI22_X1 U22933 ( .A1(n19990), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19892), .ZN(n19991) );
  INV_X1 U22934 ( .A(n19991), .ZN(P2_U3611) );
  AOI21_X1 U22935 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20735), .A(n11622), 
        .ZN(n19994) );
  INV_X1 U22936 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19992) );
  NAND2_X1 U22937 ( .A1(n11622), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20808) );
  INV_X2 U22938 ( .A(n20808), .ZN(n20772) );
  AOI21_X1 U22939 ( .B1(n19994), .B2(n19992), .A(n20772), .ZN(P1_U2802) );
  INV_X1 U22940 ( .A(P1_D_C_N_REG_SCAN_IN), .ZN(n20930) );
  NOR2_X1 U22941 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19995) );
  NOR2_X1 U22942 ( .A1(n20772), .A2(n19995), .ZN(n19993) );
  AOI22_X1 U22943 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(n20772), .B1(n20930), 
        .B2(n19993), .ZN(P1_U2804) );
  NOR2_X1 U22944 ( .A1(n20772), .A2(n19994), .ZN(n20784) );
  OAI21_X1 U22945 ( .B1(BS16), .B2(n19995), .A(n20784), .ZN(n20782) );
  OAI21_X1 U22946 ( .B1(n20784), .B2(n21127), .A(n20782), .ZN(P1_U2805) );
  OAI21_X1 U22947 ( .B1(n19997), .B2(n21005), .A(n19996), .ZN(P1_U2806) );
  NOR4_X1 U22948 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20001) );
  NOR4_X1 U22949 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20000) );
  NOR4_X1 U22950 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19999) );
  NOR4_X1 U22951 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19998) );
  NAND4_X1 U22952 ( .A1(n20001), .A2(n20000), .A3(n19999), .A4(n19998), .ZN(
        n20007) );
  NOR4_X1 U22953 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20005) );
  AOI211_X1 U22954 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20004) );
  NOR4_X1 U22955 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20003) );
  NOR4_X1 U22956 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20002) );
  NAND4_X1 U22957 ( .A1(n20005), .A2(n20004), .A3(n20003), .A4(n20002), .ZN(
        n20006) );
  NOR2_X1 U22958 ( .A1(n20007), .A2(n20006), .ZN(n20797) );
  INV_X1 U22959 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20989) );
  NOR3_X1 U22960 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20009) );
  OAI21_X1 U22961 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20009), .A(n20797), .ZN(
        n20008) );
  OAI21_X1 U22962 ( .B1(n20797), .B2(n20989), .A(n20008), .ZN(P1_U2807) );
  INV_X1 U22963 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20783) );
  AOI21_X1 U22964 ( .B1(n20904), .B2(n20783), .A(n20009), .ZN(n20010) );
  INV_X1 U22965 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20913) );
  INV_X1 U22966 ( .A(n20797), .ZN(n20793) );
  AOI22_X1 U22967 ( .A1(n20797), .A2(n20010), .B1(n20913), .B2(n20793), .ZN(
        P1_U2808) );
  INV_X1 U22968 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n20905) );
  INV_X1 U22969 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n21141) );
  NOR2_X1 U22970 ( .A1(n20905), .A2(n21141), .ZN(n20015) );
  AND3_X1 U22971 ( .A1(n21008), .A2(n20015), .A3(n20037), .ZN(n20011) );
  AOI211_X1 U22972 ( .C1(n20024), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n15899), .B(n20011), .ZN(n20014) );
  AOI22_X1 U22973 ( .A1(n20012), .A2(n20067), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n20061), .ZN(n20013) );
  AND2_X1 U22974 ( .A1(n20014), .A2(n20013), .ZN(n20019) );
  OAI21_X1 U22975 ( .B1(n20016), .B2(n20015), .A(n20060), .ZN(n20026) );
  AOI22_X1 U22976 ( .A1(n20025), .A2(n20017), .B1(n20026), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n20018) );
  OAI211_X1 U22977 ( .C1(n20020), .C2(n20063), .A(n20019), .B(n20018), .ZN(
        P1_U2833) );
  NAND2_X1 U22978 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n20037), .ZN(n20022) );
  AOI22_X1 U22979 ( .A1(n20072), .A2(n20067), .B1(n20046), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n20021) );
  OAI21_X1 U22980 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n20022), .A(n20021), .ZN(
        n20023) );
  AOI211_X1 U22981 ( .C1(n20024), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n15899), .B(n20023), .ZN(n20028) );
  AOI22_X1 U22982 ( .A1(n20026), .A2(P1_REIP_REG_6__SCAN_IN), .B1(n20025), 
        .B2(n20075), .ZN(n20027) );
  OAI211_X1 U22983 ( .C1(n20029), .C2(n20063), .A(n20028), .B(n20027), .ZN(
        P1_U2834) );
  NOR2_X1 U22984 ( .A1(n20030), .A2(n20049), .ZN(n20031) );
  AOI211_X1 U22985 ( .C1(n20061), .C2(P1_EBX_REG_5__SCAN_IN), .A(n15899), .B(
        n20031), .ZN(n20032) );
  OAI21_X1 U22986 ( .B1(n20064), .B2(n20033), .A(n20032), .ZN(n20036) );
  OAI22_X1 U22987 ( .A1(n20060), .A2(n20905), .B1(n20034), .B2(n20071), .ZN(
        n20035) );
  AOI211_X1 U22988 ( .C1(n20905), .C2(n20037), .A(n20036), .B(n20035), .ZN(
        n20038) );
  OAI21_X1 U22989 ( .B1(n20039), .B2(n20063), .A(n20038), .ZN(P1_U2835) );
  NOR2_X1 U22990 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n20040), .ZN(n20059) );
  INV_X1 U22991 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20056) );
  NAND2_X1 U22992 ( .A1(n20042), .A2(n20041), .ZN(n20055) );
  INV_X1 U22993 ( .A(n20043), .ZN(n20052) );
  INV_X1 U22994 ( .A(n20044), .ZN(n20050) );
  NAND2_X1 U22995 ( .A1(n20045), .A2(n20065), .ZN(n20048) );
  AOI21_X1 U22996 ( .B1(n20046), .B2(P1_EBX_REG_4__SCAN_IN), .A(n15935), .ZN(
        n20047) );
  OAI211_X1 U22997 ( .C1(n20050), .C2(n20049), .A(n20048), .B(n20047), .ZN(
        n20051) );
  AOI21_X1 U22998 ( .B1(n20053), .B2(n20052), .A(n20051), .ZN(n20054) );
  OAI211_X1 U22999 ( .C1(n20064), .C2(n20056), .A(n20055), .B(n20054), .ZN(
        n20057) );
  INV_X1 U23000 ( .A(n20057), .ZN(n20058) );
  OAI21_X1 U23001 ( .B1(n20060), .B2(n20059), .A(n20058), .ZN(P1_U2836) );
  AOI22_X1 U23002 ( .A1(n20062), .A2(P1_REIP_REG_0__SCAN_IN), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(n20061), .ZN(n20070) );
  NAND2_X1 U23003 ( .A1(n20064), .A2(n20063), .ZN(n20068) );
  AOI222_X1 U23004 ( .A1(n20068), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20067), .B2(n20066), .C1(n10503), .C2(n20065), .ZN(n20069) );
  OAI211_X1 U23005 ( .C1(n20071), .C2(n20132), .A(n20070), .B(n20069), .ZN(
        P1_U2840) );
  AOI22_X1 U23006 ( .A1(n20075), .A2(n20074), .B1(n20073), .B2(n20072), .ZN(
        n20076) );
  OAI21_X1 U23007 ( .B1(n20078), .B2(n20077), .A(n20076), .ZN(P1_U2866) );
  AOI22_X1 U23008 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20082), .B1(n15566), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20079) );
  OAI21_X1 U23009 ( .B1(n20081), .B2(n20080), .A(n20079), .ZN(P1_U2921) );
  INV_X1 U23010 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20084) );
  AOI22_X1 U23011 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20083) );
  OAI21_X1 U23012 ( .B1(n20084), .B2(n20108), .A(n20083), .ZN(P1_U2922) );
  AOI22_X1 U23013 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20085) );
  OAI21_X1 U23014 ( .B1(n14503), .B2(n20108), .A(n20085), .ZN(P1_U2923) );
  AOI22_X1 U23015 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20086) );
  OAI21_X1 U23016 ( .B1(n13823), .B2(n20108), .A(n20086), .ZN(P1_U2924) );
  INV_X1 U23017 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20088) );
  AOI22_X1 U23018 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20087) );
  OAI21_X1 U23019 ( .B1(n20088), .B2(n20108), .A(n20087), .ZN(P1_U2925) );
  AOI22_X1 U23020 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20089) );
  OAI21_X1 U23021 ( .B1(n13754), .B2(n20108), .A(n20089), .ZN(P1_U2926) );
  INV_X1 U23022 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20091) );
  AOI22_X1 U23023 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20090) );
  OAI21_X1 U23024 ( .B1(n20091), .B2(n20108), .A(n20090), .ZN(P1_U2927) );
  AOI22_X1 U23025 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20801), .B1(n15566), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20092) );
  OAI21_X1 U23026 ( .B1(n20093), .B2(n20108), .A(n20092), .ZN(P1_U2928) );
  AOI22_X1 U23027 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20094) );
  OAI21_X1 U23028 ( .B1(n10659), .B2(n20108), .A(n20094), .ZN(P1_U2929) );
  AOI22_X1 U23029 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20095) );
  OAI21_X1 U23030 ( .B1(n10651), .B2(n20108), .A(n20095), .ZN(P1_U2930) );
  AOI22_X1 U23031 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20096) );
  OAI21_X1 U23032 ( .B1(n20097), .B2(n20108), .A(n20096), .ZN(P1_U2931) );
  AOI22_X1 U23033 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20098) );
  OAI21_X1 U23034 ( .B1(n20099), .B2(n20108), .A(n20098), .ZN(P1_U2932) );
  AOI22_X1 U23035 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20100) );
  OAI21_X1 U23036 ( .B1(n20101), .B2(n20108), .A(n20100), .ZN(P1_U2933) );
  AOI22_X1 U23037 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20102) );
  OAI21_X1 U23038 ( .B1(n20103), .B2(n20108), .A(n20102), .ZN(P1_U2934) );
  AOI22_X1 U23039 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20104) );
  OAI21_X1 U23040 ( .B1(n20105), .B2(n20108), .A(n20104), .ZN(P1_U2935) );
  AOI22_X1 U23041 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20106), .B1(n15566), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20107) );
  OAI21_X1 U23042 ( .B1(n20109), .B2(n20108), .A(n20107), .ZN(P1_U2936) );
  AOI22_X1 U23043 ( .A1(n20121), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20120), .ZN(n20111) );
  NAND2_X1 U23044 ( .A1(n20111), .A2(n20110), .ZN(P1_U2961) );
  AOI22_X1 U23045 ( .A1(n20121), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20120), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20113) );
  NAND2_X1 U23046 ( .A1(n20113), .A2(n20112), .ZN(P1_U2962) );
  AOI22_X1 U23047 ( .A1(n20121), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20120), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20115) );
  NAND2_X1 U23048 ( .A1(n20115), .A2(n20114), .ZN(P1_U2963) );
  AOI22_X1 U23049 ( .A1(n20121), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20120), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20117) );
  NAND2_X1 U23050 ( .A1(n20117), .A2(n20116), .ZN(P1_U2964) );
  AOI22_X1 U23051 ( .A1(n20121), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20120), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20119) );
  NAND2_X1 U23052 ( .A1(n20119), .A2(n20118), .ZN(P1_U2965) );
  AOI22_X1 U23053 ( .A1(n20121), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20120), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20123) );
  NAND2_X1 U23054 ( .A1(n20123), .A2(n20122), .ZN(P1_U2966) );
  OR2_X1 U23055 ( .A1(n20125), .A2(n20124), .ZN(n20128) );
  AOI22_X1 U23056 ( .A1(n20128), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20127), .B2(n20126), .ZN(n20130) );
  OAI211_X1 U23057 ( .C1(n20132), .C2(n20131), .A(n20130), .B(n20129), .ZN(
        P1_U2999) );
  NAND2_X1 U23058 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20134) );
  OAI21_X1 U23059 ( .B1(n11540), .B2(n20134), .A(n20133), .ZN(n20142) );
  INV_X1 U23060 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n21151) );
  OAI22_X1 U23061 ( .A1(n20137), .A2(n20136), .B1(n21151), .B2(n20135), .ZN(
        n20141) );
  NOR2_X1 U23062 ( .A1(n20139), .A2(n20138), .ZN(n20140) );
  AOI211_X1 U23063 ( .C1(n20143), .C2(n20142), .A(n20141), .B(n20140), .ZN(
        n20144) );
  OAI221_X1 U23064 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20146), .C1(
        n11540), .C2(n20145), .A(n20144), .ZN(P1_U3029) );
  NOR2_X1 U23065 ( .A1(n20148), .A2(n20147), .ZN(P1_U3032) );
  INV_X1 U23066 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20155) );
  NOR2_X2 U23067 ( .A1(n20179), .A2(n20149), .ZN(n20648) );
  INV_X1 U23068 ( .A(DATAI_24_), .ZN(n21015) );
  OAI22_X2 U23069 ( .A1(n20150), .A2(n20184), .B1(n21015), .B2(n20186), .ZN(
        n20608) );
  AOI22_X1 U23070 ( .A1(n20648), .A2(n20182), .B1(n20692), .B2(n20608), .ZN(
        n20154) );
  NAND2_X1 U23071 ( .A1(n20196), .A2(n20151), .ZN(n20540) );
  INV_X1 U23072 ( .A(DATAI_16_), .ZN(n21135) );
  AOI22_X1 U23073 ( .A1(n20647), .A2(n20187), .B1(n20216), .B2(n20660), .ZN(
        n20153) );
  OAI211_X1 U23074 ( .C1(n20191), .C2(n20155), .A(n20154), .B(n20153), .ZN(
        P1_U3033) );
  NOR2_X2 U23075 ( .A1(n20179), .A2(n20156), .ZN(n20665) );
  INV_X1 U23076 ( .A(DATAI_25_), .ZN(n20157) );
  OAI22_X2 U23077 ( .A1(n14844), .A2(n20184), .B1(n20157), .B2(n20186), .ZN(
        n20612) );
  AOI22_X1 U23078 ( .A1(n20665), .A2(n20182), .B1(n20692), .B2(n20612), .ZN(
        n20160) );
  NAND2_X1 U23079 ( .A1(n20196), .A2(n20158), .ZN(n20543) );
  INV_X1 U23080 ( .A(DATAI_17_), .ZN(n21118) );
  AOI22_X1 U23081 ( .A1(n20664), .A2(n20187), .B1(n20216), .B2(n20666), .ZN(
        n20159) );
  OAI211_X1 U23082 ( .C1(n20191), .C2(n10464), .A(n20160), .B(n20159), .ZN(
        P1_U3034) );
  NOR2_X2 U23083 ( .A1(n20179), .A2(n13142), .ZN(n20671) );
  OAI22_X2 U23084 ( .A1(n20161), .A2(n20184), .B1(n14457), .B2(n20186), .ZN(
        n20616) );
  AOI22_X1 U23085 ( .A1(n20671), .A2(n20182), .B1(n20692), .B2(n20616), .ZN(
        n20165) );
  NAND2_X1 U23086 ( .A1(n20196), .A2(n20162), .ZN(n20546) );
  INV_X1 U23087 ( .A(DATAI_18_), .ZN(n21033) );
  AOI22_X1 U23088 ( .A1(n20670), .A2(n20187), .B1(n20216), .B2(n20672), .ZN(
        n20164) );
  OAI211_X1 U23089 ( .C1(n20191), .C2(n20166), .A(n20165), .B(n20164), .ZN(
        P1_U3035) );
  NOR2_X2 U23090 ( .A1(n20179), .A2(n20167), .ZN(n20677) );
  INV_X1 U23091 ( .A(DATAI_27_), .ZN(n21137) );
  OAI22_X2 U23092 ( .A1(n20168), .A2(n20184), .B1(n21137), .B2(n20186), .ZN(
        n20620) );
  AOI22_X1 U23093 ( .A1(n20677), .A2(n20182), .B1(n20692), .B2(n20620), .ZN(
        n20172) );
  NAND2_X1 U23094 ( .A1(n20196), .A2(n20169), .ZN(n20549) );
  INV_X1 U23095 ( .A(DATAI_19_), .ZN(n20170) );
  AOI22_X1 U23096 ( .A1(n20676), .A2(n20187), .B1(n20216), .B2(n20678), .ZN(
        n20171) );
  OAI211_X1 U23097 ( .C1(n20191), .C2(n20173), .A(n20172), .B(n20171), .ZN(
        P1_U3036) );
  NOR2_X2 U23098 ( .A1(n20179), .A2(n11114), .ZN(n20690) );
  INV_X1 U23099 ( .A(DATAI_29_), .ZN(n21160) );
  OAI22_X2 U23100 ( .A1(n20174), .A2(n20184), .B1(n21160), .B2(n20186), .ZN(
        n20628) );
  AOI22_X1 U23101 ( .A1(n20690), .A2(n20182), .B1(n20692), .B2(n20628), .ZN(
        n20177) );
  NAND2_X1 U23102 ( .A1(n20196), .A2(n20175), .ZN(n20555) );
  INV_X1 U23103 ( .A(DATAI_21_), .ZN(n21024) );
  AOI22_X1 U23104 ( .A1(n20689), .A2(n20187), .B1(n20216), .B2(n20691), .ZN(
        n20176) );
  OAI211_X1 U23105 ( .C1(n20191), .C2(n20178), .A(n20177), .B(n20176), .ZN(
        P1_U3038) );
  NOR2_X2 U23106 ( .A1(n20179), .A2(n10416), .ZN(n20700) );
  INV_X1 U23107 ( .A(DATAI_30_), .ZN(n20180) );
  OAI22_X2 U23108 ( .A1(n20181), .A2(n20184), .B1(n20180), .B2(n20186), .ZN(
        n20701) );
  AOI22_X1 U23109 ( .A1(n20700), .A2(n20182), .B1(n20692), .B2(n20701), .ZN(
        n20189) );
  NAND2_X1 U23110 ( .A1(n20196), .A2(n20183), .ZN(n20560) );
  INV_X1 U23111 ( .A(DATAI_22_), .ZN(n20999) );
  OAI22_X1 U23112 ( .A1(n20999), .A2(n20186), .B1(n20185), .B2(n20184), .ZN(
        n20556) );
  AOI22_X1 U23113 ( .A1(n20698), .A2(n20187), .B1(n20216), .B2(n20556), .ZN(
        n20188) );
  OAI211_X1 U23114 ( .C1(n20191), .C2(n20190), .A(n20189), .B(n20188), .ZN(
        P1_U3039) );
  INV_X1 U23115 ( .A(n20660), .ZN(n20611) );
  INV_X1 U23116 ( .A(n20569), .ZN(n20192) );
  NOR2_X1 U23117 ( .A1(n20570), .A2(n20195), .ZN(n20215) );
  INV_X1 U23118 ( .A(n20254), .ZN(n20194) );
  INV_X1 U23119 ( .A(n20193), .ZN(n20571) );
  AOI21_X1 U23120 ( .B1(n20194), .B2(n20571), .A(n20215), .ZN(n20197) );
  OAI22_X1 U23121 ( .A1(n20197), .A2(n20651), .B1(n20195), .B2(n20721), .ZN(
        n20214) );
  AOI22_X1 U23122 ( .A1(n20648), .A2(n20215), .B1(n20647), .B2(n20214), .ZN(
        n20201) );
  INV_X1 U23123 ( .A(n20195), .ZN(n20199) );
  OAI21_X1 U23124 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20537), .A(
        n20196), .ZN(n20257) );
  OAI211_X1 U23125 ( .C1(n20262), .C2(n21127), .A(n20658), .B(n20197), .ZN(
        n20198) );
  OAI211_X1 U23126 ( .C1(n20658), .C2(n20199), .A(n20657), .B(n20198), .ZN(
        n20217) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20608), .ZN(n20200) );
  OAI211_X1 U23128 ( .C1(n20611), .C2(n20244), .A(n20201), .B(n20200), .ZN(
        P1_U3041) );
  INV_X1 U23129 ( .A(n20666), .ZN(n20615) );
  AOI22_X1 U23130 ( .A1(n20665), .A2(n20215), .B1(n20664), .B2(n20214), .ZN(
        n20203) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20612), .ZN(n20202) );
  OAI211_X1 U23132 ( .C1(n20615), .C2(n20244), .A(n20203), .B(n20202), .ZN(
        P1_U3042) );
  INV_X1 U23133 ( .A(n20672), .ZN(n20619) );
  AOI22_X1 U23134 ( .A1(n20671), .A2(n20215), .B1(n20670), .B2(n20214), .ZN(
        n20205) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20616), .ZN(n20204) );
  OAI211_X1 U23136 ( .C1(n20619), .C2(n20244), .A(n20205), .B(n20204), .ZN(
        P1_U3043) );
  INV_X1 U23137 ( .A(n20678), .ZN(n20623) );
  AOI22_X1 U23138 ( .A1(n20677), .A2(n20215), .B1(n20676), .B2(n20214), .ZN(
        n20207) );
  AOI22_X1 U23139 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20620), .ZN(n20206) );
  OAI211_X1 U23140 ( .C1(n20623), .C2(n20244), .A(n20207), .B(n20206), .ZN(
        P1_U3044) );
  INV_X1 U23141 ( .A(n20509), .ZN(n20688) );
  AOI22_X1 U23142 ( .A1(n20625), .A2(n20215), .B1(n20624), .B2(n20214), .ZN(
        n20209) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20685), .ZN(n20208) );
  OAI211_X1 U23144 ( .C1(n20688), .C2(n20244), .A(n20209), .B(n20208), .ZN(
        P1_U3045) );
  INV_X1 U23145 ( .A(n20691), .ZN(n20631) );
  AOI22_X1 U23146 ( .A1(n20690), .A2(n20215), .B1(n20689), .B2(n20214), .ZN(
        n20211) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20628), .ZN(n20210) );
  OAI211_X1 U23148 ( .C1(n20631), .C2(n20244), .A(n20211), .B(n20210), .ZN(
        P1_U3046) );
  INV_X1 U23149 ( .A(n20556), .ZN(n20704) );
  AOI22_X1 U23150 ( .A1(n20700), .A2(n20215), .B1(n20698), .B2(n20214), .ZN(
        n20213) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20701), .ZN(n20212) );
  OAI211_X1 U23152 ( .C1(n20704), .C2(n20244), .A(n20213), .B(n20212), .ZN(
        P1_U3047) );
  INV_X1 U23153 ( .A(n20520), .ZN(n20716) );
  AOI22_X1 U23154 ( .A1(n20637), .A2(n20215), .B1(n20635), .B2(n20214), .ZN(
        n20219) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20217), .B1(
        n20216), .B2(n20710), .ZN(n20218) );
  OAI211_X1 U23156 ( .C1(n20716), .C2(n20244), .A(n20219), .B(n20218), .ZN(
        P1_U3048) );
  NOR3_X1 U23157 ( .A1(n20278), .A2(n20239), .A3(n20651), .ZN(n20221) );
  INV_X1 U23158 ( .A(n20527), .ZN(n20313) );
  NOR2_X1 U23159 ( .A1(n20221), .A2(n20313), .ZN(n20225) );
  INV_X1 U23160 ( .A(n20225), .ZN(n20222) );
  NOR2_X1 U23161 ( .A1(n20254), .A2(n13514), .ZN(n20224) );
  NAND3_X1 U23162 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20489), .A3(
        n15515), .ZN(n20258) );
  NOR2_X1 U23163 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20258), .ZN(
        n20238) );
  AOI22_X1 U23164 ( .A1(n20239), .A2(n20608), .B1(n20648), .B2(n20238), .ZN(
        n20227) );
  INV_X1 U23165 ( .A(n20238), .ZN(n20242) );
  NOR2_X1 U23166 ( .A1(n10223), .A2(n20721), .ZN(n20340) );
  AOI211_X1 U23167 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20242), .A(n20340), 
        .B(n20403), .ZN(n20223) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20246), .B1(
        n20278), .B2(n20660), .ZN(n20226) );
  OAI211_X1 U23169 ( .C1(n20249), .C2(n20540), .A(n20227), .B(n20226), .ZN(
        P1_U3049) );
  AOI22_X1 U23170 ( .A1(n20239), .A2(n20612), .B1(n20665), .B2(n20238), .ZN(
        n20229) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20246), .B1(
        n20278), .B2(n20666), .ZN(n20228) );
  OAI211_X1 U23172 ( .C1(n20249), .C2(n20543), .A(n20229), .B(n20228), .ZN(
        P1_U3050) );
  AOI22_X1 U23173 ( .A1(n20239), .A2(n20616), .B1(n20671), .B2(n20238), .ZN(
        n20231) );
  AOI22_X1 U23174 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20246), .B1(
        n20278), .B2(n20672), .ZN(n20230) );
  OAI211_X1 U23175 ( .C1(n20249), .C2(n20546), .A(n20231), .B(n20230), .ZN(
        P1_U3051) );
  AOI22_X1 U23176 ( .A1(n20278), .A2(n20678), .B1(n20677), .B2(n20238), .ZN(
        n20233) );
  AOI22_X1 U23177 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20246), .B1(
        n20239), .B2(n20620), .ZN(n20232) );
  OAI211_X1 U23178 ( .C1(n20249), .C2(n20549), .A(n20233), .B(n20232), .ZN(
        P1_U3052) );
  AOI22_X1 U23179 ( .A1(n20278), .A2(n20509), .B1(n20625), .B2(n20238), .ZN(
        n20235) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20246), .B1(
        n20239), .B2(n20685), .ZN(n20234) );
  OAI211_X1 U23181 ( .C1(n20249), .C2(n20682), .A(n20235), .B(n20234), .ZN(
        P1_U3053) );
  AOI22_X1 U23182 ( .A1(n20278), .A2(n20691), .B1(n20690), .B2(n20238), .ZN(
        n20237) );
  AOI22_X1 U23183 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20246), .B1(
        n20239), .B2(n20628), .ZN(n20236) );
  OAI211_X1 U23184 ( .C1(n20249), .C2(n20555), .A(n20237), .B(n20236), .ZN(
        P1_U3054) );
  AOI22_X1 U23185 ( .A1(n20278), .A2(n20556), .B1(n20700), .B2(n20238), .ZN(
        n20241) );
  AOI22_X1 U23186 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20246), .B1(
        n20239), .B2(n20701), .ZN(n20240) );
  OAI211_X1 U23187 ( .C1(n20249), .C2(n20560), .A(n20241), .B(n20240), .ZN(
        P1_U3055) );
  OR2_X1 U23188 ( .A1(n20708), .A2(n20242), .ZN(n20243) );
  OAI21_X1 U23189 ( .B1(n20244), .B2(n20525), .A(n20243), .ZN(n20245) );
  INV_X1 U23190 ( .A(n20245), .ZN(n20248) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20246), .B1(
        n20278), .B2(n20520), .ZN(n20247) );
  OAI211_X1 U23192 ( .C1(n20249), .C2(n20706), .A(n20248), .B(n20247), .ZN(
        P1_U3056) );
  INV_X1 U23193 ( .A(n20258), .ZN(n20256) );
  OR2_X1 U23194 ( .A1(n20250), .A2(n20651), .ZN(n20251) );
  AND2_X1 U23195 ( .A1(n20251), .A2(n20650), .ZN(n20261) );
  INV_X1 U23196 ( .A(n20261), .ZN(n20255) );
  AND2_X1 U23197 ( .A1(n20252), .A2(n10503), .ZN(n20491) );
  INV_X1 U23198 ( .A(n20491), .ZN(n20642) );
  NOR2_X1 U23199 ( .A1(n20490), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20277) );
  INV_X1 U23200 ( .A(n20277), .ZN(n20253) );
  OAI21_X1 U23201 ( .B1(n20254), .B2(n20642), .A(n20253), .ZN(n20260) );
  AOI22_X1 U23202 ( .A1(n20278), .A2(n20608), .B1(n20277), .B2(n20648), .ZN(
        n20264) );
  AOI21_X1 U23203 ( .B1(n20651), .B2(n20258), .A(n20257), .ZN(n20259) );
  OAI21_X1 U23204 ( .B1(n20261), .B2(n20260), .A(n20259), .ZN(n20279) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20279), .B1(
        n20307), .B2(n20660), .ZN(n20263) );
  OAI211_X1 U23206 ( .C1(n20282), .C2(n20540), .A(n20264), .B(n20263), .ZN(
        P1_U3057) );
  AOI22_X1 U23207 ( .A1(n20307), .A2(n20666), .B1(n20665), .B2(n20277), .ZN(
        n20266) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20612), .ZN(n20265) );
  OAI211_X1 U23209 ( .C1(n20282), .C2(n20543), .A(n20266), .B(n20265), .ZN(
        P1_U3058) );
  AOI22_X1 U23210 ( .A1(n20278), .A2(n20616), .B1(n20277), .B2(n20671), .ZN(
        n20268) );
  AOI22_X1 U23211 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20279), .B1(
        n20307), .B2(n20672), .ZN(n20267) );
  OAI211_X1 U23212 ( .C1(n20282), .C2(n20546), .A(n20268), .B(n20267), .ZN(
        P1_U3059) );
  AOI22_X1 U23213 ( .A1(n20307), .A2(n20678), .B1(n20277), .B2(n20677), .ZN(
        n20270) );
  AOI22_X1 U23214 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20620), .ZN(n20269) );
  OAI211_X1 U23215 ( .C1(n20282), .C2(n20549), .A(n20270), .B(n20269), .ZN(
        P1_U3060) );
  AOI22_X1 U23216 ( .A1(n20278), .A2(n20685), .B1(n20625), .B2(n20277), .ZN(
        n20272) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20279), .B1(
        n20307), .B2(n20509), .ZN(n20271) );
  OAI211_X1 U23218 ( .C1(n20282), .C2(n20682), .A(n20272), .B(n20271), .ZN(
        P1_U3061) );
  AOI22_X1 U23219 ( .A1(n20307), .A2(n20691), .B1(n20277), .B2(n20690), .ZN(
        n20274) );
  AOI22_X1 U23220 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20628), .ZN(n20273) );
  OAI211_X1 U23221 ( .C1(n20282), .C2(n20555), .A(n20274), .B(n20273), .ZN(
        P1_U3062) );
  AOI22_X1 U23222 ( .A1(n20307), .A2(n20556), .B1(n20277), .B2(n20700), .ZN(
        n20276) );
  AOI22_X1 U23223 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20279), .B1(
        n20278), .B2(n20701), .ZN(n20275) );
  OAI211_X1 U23224 ( .C1(n20282), .C2(n20560), .A(n20276), .B(n20275), .ZN(
        P1_U3063) );
  AOI22_X1 U23225 ( .A1(n20278), .A2(n20710), .B1(n20637), .B2(n20277), .ZN(
        n20281) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20279), .B1(
        n20307), .B2(n20520), .ZN(n20280) );
  OAI211_X1 U23227 ( .C1(n20282), .C2(n20706), .A(n20281), .B(n20280), .ZN(
        P1_U3064) );
  NAND3_X1 U23228 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20489), .A3(
        n20531), .ZN(n20311) );
  NOR2_X1 U23229 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20311), .ZN(
        n20306) );
  NOR2_X1 U23230 ( .A1(n13310), .A2(n20283), .ZN(n20369) );
  NAND3_X1 U23231 ( .A1(n20369), .A2(n20658), .A3(n13514), .ZN(n20284) );
  OAI21_X1 U23232 ( .B1(n20600), .B2(n20285), .A(n20284), .ZN(n20305) );
  AOI22_X1 U23233 ( .A1(n20648), .A2(n20306), .B1(n20647), .B2(n20305), .ZN(
        n20292) );
  INV_X1 U23234 ( .A(n20307), .ZN(n20286) );
  AOI21_X1 U23235 ( .B1(n20286), .B2(n20335), .A(n21127), .ZN(n20287) );
  AOI21_X1 U23236 ( .B1(n20369), .B2(n13514), .A(n20287), .ZN(n20288) );
  NOR2_X1 U23237 ( .A1(n20288), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20290) );
  AOI22_X1 U23238 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20608), .ZN(n20291) );
  OAI211_X1 U23239 ( .C1(n20611), .C2(n20335), .A(n20292), .B(n20291), .ZN(
        P1_U3065) );
  AOI22_X1 U23240 ( .A1(n20665), .A2(n20306), .B1(n20664), .B2(n20305), .ZN(
        n20294) );
  AOI22_X1 U23241 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20612), .ZN(n20293) );
  OAI211_X1 U23242 ( .C1(n20615), .C2(n20335), .A(n20294), .B(n20293), .ZN(
        P1_U3066) );
  AOI22_X1 U23243 ( .A1(n20671), .A2(n20306), .B1(n20670), .B2(n20305), .ZN(
        n20296) );
  AOI22_X1 U23244 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20616), .ZN(n20295) );
  OAI211_X1 U23245 ( .C1(n20619), .C2(n20335), .A(n20296), .B(n20295), .ZN(
        P1_U3067) );
  AOI22_X1 U23246 ( .A1(n20677), .A2(n20306), .B1(n20676), .B2(n20305), .ZN(
        n20298) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20620), .ZN(n20297) );
  OAI211_X1 U23248 ( .C1(n20623), .C2(n20335), .A(n20298), .B(n20297), .ZN(
        P1_U3068) );
  AOI22_X1 U23249 ( .A1(n20625), .A2(n20306), .B1(n20624), .B2(n20305), .ZN(
        n20300) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20685), .ZN(n20299) );
  OAI211_X1 U23251 ( .C1(n20688), .C2(n20335), .A(n20300), .B(n20299), .ZN(
        P1_U3069) );
  AOI22_X1 U23252 ( .A1(n20690), .A2(n20306), .B1(n20689), .B2(n20305), .ZN(
        n20302) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20628), .ZN(n20301) );
  OAI211_X1 U23254 ( .C1(n20631), .C2(n20335), .A(n20302), .B(n20301), .ZN(
        P1_U3070) );
  AOI22_X1 U23255 ( .A1(n20700), .A2(n20306), .B1(n20698), .B2(n20305), .ZN(
        n20304) );
  AOI22_X1 U23256 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20701), .ZN(n20303) );
  OAI211_X1 U23257 ( .C1(n20704), .C2(n20335), .A(n20304), .B(n20303), .ZN(
        P1_U3071) );
  AOI22_X1 U23258 ( .A1(n20637), .A2(n20306), .B1(n20635), .B2(n20305), .ZN(
        n20310) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20710), .ZN(n20309) );
  OAI211_X1 U23260 ( .C1(n20716), .C2(n20335), .A(n20310), .B(n20309), .ZN(
        P1_U3072) );
  INV_X1 U23261 ( .A(n20608), .ZN(n20663) );
  NOR2_X1 U23262 ( .A1(n20570), .A2(n20311), .ZN(n20331) );
  AOI21_X1 U23263 ( .B1(n20369), .B2(n20571), .A(n20331), .ZN(n20312) );
  OAI22_X1 U23264 ( .A1(n20312), .A2(n20651), .B1(n20311), .B2(n20721), .ZN(
        n20330) );
  AOI22_X1 U23265 ( .A1(n20648), .A2(n20331), .B1(n20647), .B2(n20330), .ZN(
        n20317) );
  INV_X1 U23266 ( .A(n20311), .ZN(n20315) );
  OAI21_X1 U23267 ( .B1(n20368), .B2(n20313), .A(n20312), .ZN(n20314) );
  OAI211_X1 U23268 ( .C1(n20658), .C2(n20315), .A(n20657), .B(n20314), .ZN(
        n20332) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20660), .ZN(n20316) );
  OAI211_X1 U23270 ( .C1(n20663), .C2(n20335), .A(n20317), .B(n20316), .ZN(
        P1_U3073) );
  INV_X1 U23271 ( .A(n20612), .ZN(n20669) );
  AOI22_X1 U23272 ( .A1(n20665), .A2(n20331), .B1(n20664), .B2(n20330), .ZN(
        n20319) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20666), .ZN(n20318) );
  OAI211_X1 U23274 ( .C1(n20669), .C2(n20335), .A(n20319), .B(n20318), .ZN(
        P1_U3074) );
  INV_X1 U23275 ( .A(n20616), .ZN(n20675) );
  AOI22_X1 U23276 ( .A1(n20671), .A2(n20331), .B1(n20670), .B2(n20330), .ZN(
        n20321) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20672), .ZN(n20320) );
  OAI211_X1 U23278 ( .C1(n20675), .C2(n20335), .A(n20321), .B(n20320), .ZN(
        P1_U3075) );
  INV_X1 U23279 ( .A(n20620), .ZN(n20681) );
  AOI22_X1 U23280 ( .A1(n20677), .A2(n20331), .B1(n20676), .B2(n20330), .ZN(
        n20323) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20678), .ZN(n20322) );
  OAI211_X1 U23282 ( .C1(n20681), .C2(n20335), .A(n20323), .B(n20322), .ZN(
        P1_U3076) );
  AOI22_X1 U23283 ( .A1(n20625), .A2(n20331), .B1(n20624), .B2(n20330), .ZN(
        n20325) );
  AOI22_X1 U23284 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20509), .ZN(n20324) );
  OAI211_X1 U23285 ( .C1(n20512), .C2(n20335), .A(n20325), .B(n20324), .ZN(
        P1_U3077) );
  INV_X1 U23286 ( .A(n20628), .ZN(n20696) );
  AOI22_X1 U23287 ( .A1(n20690), .A2(n20331), .B1(n20689), .B2(n20330), .ZN(
        n20327) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20691), .ZN(n20326) );
  OAI211_X1 U23289 ( .C1(n20696), .C2(n20335), .A(n20327), .B(n20326), .ZN(
        P1_U3078) );
  INV_X1 U23290 ( .A(n20701), .ZN(n20517) );
  AOI22_X1 U23291 ( .A1(n20700), .A2(n20331), .B1(n20698), .B2(n20330), .ZN(
        n20329) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20556), .ZN(n20328) );
  OAI211_X1 U23293 ( .C1(n20517), .C2(n20335), .A(n20329), .B(n20328), .ZN(
        P1_U3079) );
  AOI22_X1 U23294 ( .A1(n20637), .A2(n20331), .B1(n20635), .B2(n20330), .ZN(
        n20334) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20332), .B1(
        n20363), .B2(n20520), .ZN(n20333) );
  OAI211_X1 U23296 ( .C1(n20525), .C2(n20335), .A(n20334), .B(n20333), .ZN(
        P1_U3080) );
  NAND3_X1 U23297 ( .A1(n20360), .A2(n20336), .A3(n20658), .ZN(n20337) );
  NAND2_X1 U23298 ( .A1(n20337), .A2(n20527), .ZN(n20342) );
  AND2_X1 U23299 ( .A1(n20369), .A2(n20598), .ZN(n20339) );
  INV_X1 U23300 ( .A(n20600), .ZN(n20530) );
  INV_X1 U23301 ( .A(n20375), .ZN(n20338) );
  NOR2_X1 U23302 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20338), .ZN(
        n20357) );
  AOI22_X1 U23303 ( .A1(n20648), .A2(n20357), .B1(n20363), .B2(n20608), .ZN(
        n20345) );
  INV_X1 U23304 ( .A(n20339), .ZN(n20341) );
  AOI21_X1 U23305 ( .B1(n20342), .B2(n20341), .A(n20340), .ZN(n20343) );
  OAI211_X1 U23306 ( .C1(n20357), .C2(n20537), .A(n20606), .B(n20343), .ZN(
        n20364) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20364), .B1(
        n20396), .B2(n20660), .ZN(n20344) );
  OAI211_X1 U23308 ( .C1(n20367), .C2(n20540), .A(n20345), .B(n20344), .ZN(
        P1_U3081) );
  AOI22_X1 U23309 ( .A1(n20665), .A2(n20357), .B1(n20396), .B2(n20666), .ZN(
        n20347) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20364), .B1(
        n20363), .B2(n20612), .ZN(n20346) );
  OAI211_X1 U23311 ( .C1(n20367), .C2(n20543), .A(n20347), .B(n20346), .ZN(
        P1_U3082) );
  AOI22_X1 U23312 ( .A1(n20671), .A2(n20357), .B1(n20363), .B2(n20616), .ZN(
        n20349) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20364), .B1(
        n20396), .B2(n20672), .ZN(n20348) );
  OAI211_X1 U23314 ( .C1(n20367), .C2(n20546), .A(n20349), .B(n20348), .ZN(
        P1_U3083) );
  AOI22_X1 U23315 ( .A1(n20677), .A2(n20357), .B1(n20396), .B2(n20678), .ZN(
        n20351) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20364), .B1(
        n20363), .B2(n20620), .ZN(n20350) );
  OAI211_X1 U23317 ( .C1(n20367), .C2(n20549), .A(n20351), .B(n20350), .ZN(
        P1_U3084) );
  INV_X1 U23318 ( .A(n20357), .ZN(n20361) );
  OAI22_X1 U23319 ( .A1(n20683), .A2(n20361), .B1(n20688), .B2(n20360), .ZN(
        n20352) );
  INV_X1 U23320 ( .A(n20352), .ZN(n20354) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20364), .B1(
        n20363), .B2(n20685), .ZN(n20353) );
  OAI211_X1 U23322 ( .C1(n20367), .C2(n20682), .A(n20354), .B(n20353), .ZN(
        P1_U3085) );
  AOI22_X1 U23323 ( .A1(n20690), .A2(n20357), .B1(n20363), .B2(n20628), .ZN(
        n20356) );
  AOI22_X1 U23324 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20364), .B1(
        n20396), .B2(n20691), .ZN(n20355) );
  OAI211_X1 U23325 ( .C1(n20367), .C2(n20555), .A(n20356), .B(n20355), .ZN(
        P1_U3086) );
  AOI22_X1 U23326 ( .A1(n20700), .A2(n20357), .B1(n20396), .B2(n20556), .ZN(
        n20359) );
  AOI22_X1 U23327 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20364), .B1(
        n20363), .B2(n20701), .ZN(n20358) );
  OAI211_X1 U23328 ( .C1(n20367), .C2(n20560), .A(n20359), .B(n20358), .ZN(
        P1_U3087) );
  OAI22_X1 U23329 ( .A1(n20708), .A2(n20361), .B1(n20716), .B2(n20360), .ZN(
        n20362) );
  INV_X1 U23330 ( .A(n20362), .ZN(n20366) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20364), .B1(
        n20363), .B2(n20710), .ZN(n20365) );
  OAI211_X1 U23332 ( .C1(n20367), .C2(n20706), .A(n20366), .B(n20365), .ZN(
        P1_U3088) );
  INV_X1 U23333 ( .A(n20394), .ZN(n20390) );
  NAND2_X1 U23334 ( .A1(n20369), .A2(n20491), .ZN(n20370) );
  NAND2_X1 U23335 ( .A1(n20370), .A2(n20394), .ZN(n20371) );
  NAND2_X1 U23336 ( .A1(n20371), .A2(n20658), .ZN(n20373) );
  NAND2_X1 U23337 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20375), .ZN(n20372) );
  AND2_X1 U23338 ( .A1(n20373), .A2(n20372), .ZN(n20393) );
  AOI22_X1 U23339 ( .A1(n20648), .A2(n20390), .B1(n20647), .B2(n20389), .ZN(
        n20377) );
  OAI21_X1 U23340 ( .B1(n20375), .B2(n20374), .A(n20657), .ZN(n20397) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20608), .ZN(n20376) );
  OAI211_X1 U23342 ( .C1(n20611), .C2(n20404), .A(n20377), .B(n20376), .ZN(
        P1_U3089) );
  AOI22_X1 U23343 ( .A1(n20665), .A2(n20390), .B1(n20664), .B2(n20389), .ZN(
        n20379) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20612), .ZN(n20378) );
  OAI211_X1 U23345 ( .C1(n20615), .C2(n20404), .A(n20379), .B(n20378), .ZN(
        P1_U3090) );
  AOI22_X1 U23346 ( .A1(n20671), .A2(n20390), .B1(n20670), .B2(n20389), .ZN(
        n20381) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20616), .ZN(n20380) );
  OAI211_X1 U23348 ( .C1(n20619), .C2(n20404), .A(n20381), .B(n20380), .ZN(
        P1_U3091) );
  AOI22_X1 U23349 ( .A1(n20677), .A2(n20390), .B1(n20676), .B2(n20389), .ZN(
        n20383) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20620), .ZN(n20382) );
  OAI211_X1 U23351 ( .C1(n20623), .C2(n20404), .A(n20383), .B(n20382), .ZN(
        P1_U3092) );
  OAI22_X1 U23352 ( .A1(n20683), .A2(n20394), .B1(n20682), .B2(n20393), .ZN(
        n20384) );
  INV_X1 U23353 ( .A(n20384), .ZN(n20386) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20685), .ZN(n20385) );
  OAI211_X1 U23355 ( .C1(n20688), .C2(n20404), .A(n20386), .B(n20385), .ZN(
        P1_U3093) );
  AOI22_X1 U23356 ( .A1(n20690), .A2(n20390), .B1(n20689), .B2(n20389), .ZN(
        n20388) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20628), .ZN(n20387) );
  OAI211_X1 U23358 ( .C1(n20631), .C2(n20404), .A(n20388), .B(n20387), .ZN(
        P1_U3094) );
  AOI22_X1 U23359 ( .A1(n20700), .A2(n20390), .B1(n20698), .B2(n20389), .ZN(
        n20392) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20701), .ZN(n20391) );
  OAI211_X1 U23361 ( .C1(n20704), .C2(n20404), .A(n20392), .B(n20391), .ZN(
        P1_U3095) );
  OAI22_X1 U23362 ( .A1(n20708), .A2(n20394), .B1(n20706), .B2(n20393), .ZN(
        n20395) );
  INV_X1 U23363 ( .A(n20395), .ZN(n20399) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20397), .B1(
        n20396), .B2(n20710), .ZN(n20398) );
  OAI211_X1 U23365 ( .C1(n20716), .C2(n20404), .A(n20399), .B(n20398), .ZN(
        P1_U3096) );
  NAND3_X1 U23366 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n15515), .A3(
        n20531), .ZN(n20429) );
  NOR2_X1 U23367 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20429), .ZN(
        n20424) );
  AOI21_X1 U23368 ( .B1(n20492), .B2(n13514), .A(n20424), .ZN(n20406) );
  AND2_X1 U23369 ( .A1(n20401), .A2(n20456), .ZN(n20529) );
  INV_X1 U23370 ( .A(n20529), .ZN(n20533) );
  OAI22_X1 U23371 ( .A1(n20406), .A2(n20651), .B1(n20402), .B2(n20533), .ZN(
        n20423) );
  AOI22_X1 U23372 ( .A1(n20648), .A2(n20424), .B1(n20647), .B2(n20423), .ZN(
        n20410) );
  INV_X1 U23373 ( .A(n20403), .ZN(n20460) );
  INV_X1 U23374 ( .A(n20452), .ZN(n20405) );
  OAI21_X1 U23375 ( .B1(n20405), .B2(n20425), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20407) );
  NAND2_X1 U23376 ( .A1(n20407), .A2(n20406), .ZN(n20408) );
  AOI22_X1 U23377 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20608), .ZN(n20409) );
  OAI211_X1 U23378 ( .C1(n20611), .C2(n20452), .A(n20410), .B(n20409), .ZN(
        P1_U3097) );
  AOI22_X1 U23379 ( .A1(n20665), .A2(n20424), .B1(n20423), .B2(n20664), .ZN(
        n20412) );
  AOI22_X1 U23380 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20612), .ZN(n20411) );
  OAI211_X1 U23381 ( .C1(n20615), .C2(n20452), .A(n20412), .B(n20411), .ZN(
        P1_U3098) );
  AOI22_X1 U23382 ( .A1(n20671), .A2(n20424), .B1(n20423), .B2(n20670), .ZN(
        n20414) );
  AOI22_X1 U23383 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20616), .ZN(n20413) );
  OAI211_X1 U23384 ( .C1(n20619), .C2(n20452), .A(n20414), .B(n20413), .ZN(
        P1_U3099) );
  AOI22_X1 U23385 ( .A1(n20677), .A2(n20424), .B1(n20423), .B2(n20676), .ZN(
        n20416) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20620), .ZN(n20415) );
  OAI211_X1 U23387 ( .C1(n20623), .C2(n20452), .A(n20416), .B(n20415), .ZN(
        P1_U3100) );
  AOI22_X1 U23388 ( .A1(n20625), .A2(n20424), .B1(n20624), .B2(n20423), .ZN(
        n20418) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20685), .ZN(n20417) );
  OAI211_X1 U23390 ( .C1(n20688), .C2(n20452), .A(n20418), .B(n20417), .ZN(
        P1_U3101) );
  AOI22_X1 U23391 ( .A1(n20690), .A2(n20424), .B1(n20423), .B2(n20689), .ZN(
        n20420) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20628), .ZN(n20419) );
  OAI211_X1 U23393 ( .C1(n20631), .C2(n20452), .A(n20420), .B(n20419), .ZN(
        P1_U3102) );
  AOI22_X1 U23394 ( .A1(n20700), .A2(n20424), .B1(n20423), .B2(n20698), .ZN(
        n20422) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20701), .ZN(n20421) );
  OAI211_X1 U23396 ( .C1(n20704), .C2(n20452), .A(n20422), .B(n20421), .ZN(
        P1_U3103) );
  AOI22_X1 U23397 ( .A1(n20637), .A2(n20424), .B1(n20635), .B2(n20423), .ZN(
        n20428) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20426), .B1(
        n20425), .B2(n20710), .ZN(n20427) );
  OAI211_X1 U23399 ( .C1(n20716), .C2(n20452), .A(n20428), .B(n20427), .ZN(
        P1_U3104) );
  NOR2_X1 U23400 ( .A1(n20570), .A2(n20429), .ZN(n20448) );
  AOI21_X1 U23401 ( .B1(n20492), .B2(n20571), .A(n20448), .ZN(n20430) );
  OAI22_X1 U23402 ( .A1(n20430), .A2(n20651), .B1(n20429), .B2(n20721), .ZN(
        n20447) );
  AOI22_X1 U23403 ( .A1(n20648), .A2(n20448), .B1(n20647), .B2(n20447), .ZN(
        n20434) );
  INV_X1 U23404 ( .A(n20429), .ZN(n20432) );
  OAI211_X1 U23405 ( .C1(n20500), .C2(n21127), .A(n20658), .B(n20430), .ZN(
        n20431) );
  OAI211_X1 U23406 ( .C1(n20658), .C2(n20432), .A(n20657), .B(n20431), .ZN(
        n20449) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20660), .ZN(n20433) );
  OAI211_X1 U23408 ( .C1(n20663), .C2(n20452), .A(n20434), .B(n20433), .ZN(
        P1_U3105) );
  AOI22_X1 U23409 ( .A1(n20665), .A2(n20448), .B1(n20664), .B2(n20447), .ZN(
        n20436) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20666), .ZN(n20435) );
  OAI211_X1 U23411 ( .C1(n20669), .C2(n20452), .A(n20436), .B(n20435), .ZN(
        P1_U3106) );
  AOI22_X1 U23412 ( .A1(n20671), .A2(n20448), .B1(n20670), .B2(n20447), .ZN(
        n20438) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20672), .ZN(n20437) );
  OAI211_X1 U23414 ( .C1(n20675), .C2(n20452), .A(n20438), .B(n20437), .ZN(
        P1_U3107) );
  AOI22_X1 U23415 ( .A1(n20677), .A2(n20448), .B1(n20676), .B2(n20447), .ZN(
        n20440) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20678), .ZN(n20439) );
  OAI211_X1 U23417 ( .C1(n20681), .C2(n20452), .A(n20440), .B(n20439), .ZN(
        P1_U3108) );
  AOI22_X1 U23418 ( .A1(n20625), .A2(n20448), .B1(n20624), .B2(n20447), .ZN(
        n20442) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20509), .ZN(n20441) );
  OAI211_X1 U23420 ( .C1(n20512), .C2(n20452), .A(n20442), .B(n20441), .ZN(
        P1_U3109) );
  AOI22_X1 U23421 ( .A1(n20690), .A2(n20448), .B1(n20689), .B2(n20447), .ZN(
        n20444) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20691), .ZN(n20443) );
  OAI211_X1 U23423 ( .C1(n20696), .C2(n20452), .A(n20444), .B(n20443), .ZN(
        P1_U3110) );
  AOI22_X1 U23424 ( .A1(n20700), .A2(n20448), .B1(n20698), .B2(n20447), .ZN(
        n20446) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20556), .ZN(n20445) );
  OAI211_X1 U23426 ( .C1(n20517), .C2(n20452), .A(n20446), .B(n20445), .ZN(
        P1_U3111) );
  AOI22_X1 U23427 ( .A1(n20637), .A2(n20448), .B1(n20635), .B2(n20447), .ZN(
        n20451) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20449), .B1(
        n20484), .B2(n20520), .ZN(n20450) );
  OAI211_X1 U23429 ( .C1(n20525), .C2(n20452), .A(n20451), .B(n20450), .ZN(
        P1_U3112) );
  INV_X1 U23430 ( .A(n20484), .ZN(n20454) );
  NAND3_X1 U23431 ( .A1(n20454), .A2(n20658), .A3(n20524), .ZN(n20455) );
  NAND2_X1 U23432 ( .A1(n20455), .A2(n20527), .ZN(n20463) );
  AND2_X1 U23433 ( .A1(n20492), .A2(n20598), .ZN(n20459) );
  OR2_X1 U23434 ( .A1(n20456), .A2(n20489), .ZN(n20601) );
  INV_X1 U23435 ( .A(n20601), .ZN(n20457) );
  NAND3_X1 U23436 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n15515), .ZN(n20493) );
  NOR2_X1 U23437 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20493), .ZN(
        n20478) );
  AOI22_X1 U23438 ( .A1(n20479), .A2(n20660), .B1(n20648), .B2(n20478), .ZN(
        n20466) );
  INV_X1 U23439 ( .A(n20459), .ZN(n20462) );
  NAND2_X1 U23440 ( .A1(n20601), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20605) );
  OAI211_X1 U23441 ( .C1(n20537), .C2(n20478), .A(n20605), .B(n20460), .ZN(
        n20461) );
  AOI21_X1 U23442 ( .B1(n20463), .B2(n20462), .A(n20461), .ZN(n20464) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20485), .B1(
        n20484), .B2(n20608), .ZN(n20465) );
  OAI211_X1 U23444 ( .C1(n20488), .C2(n20540), .A(n20466), .B(n20465), .ZN(
        P1_U3113) );
  AOI22_X1 U23445 ( .A1(n20484), .A2(n20612), .B1(n20665), .B2(n20478), .ZN(
        n20468) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20485), .B1(
        n20479), .B2(n20666), .ZN(n20467) );
  OAI211_X1 U23447 ( .C1(n20488), .C2(n20543), .A(n20468), .B(n20467), .ZN(
        P1_U3114) );
  AOI22_X1 U23448 ( .A1(n20479), .A2(n20672), .B1(n20671), .B2(n20478), .ZN(
        n20470) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20485), .B1(
        n20484), .B2(n20616), .ZN(n20469) );
  OAI211_X1 U23450 ( .C1(n20488), .C2(n20546), .A(n20470), .B(n20469), .ZN(
        P1_U3115) );
  AOI22_X1 U23451 ( .A1(n20484), .A2(n20620), .B1(n20677), .B2(n20478), .ZN(
        n20472) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20485), .B1(
        n20479), .B2(n20678), .ZN(n20471) );
  OAI211_X1 U23453 ( .C1(n20488), .C2(n20549), .A(n20472), .B(n20471), .ZN(
        P1_U3116) );
  INV_X1 U23454 ( .A(n20478), .ZN(n20482) );
  OAI22_X1 U23455 ( .A1(n20524), .A2(n20688), .B1(n20683), .B2(n20482), .ZN(
        n20473) );
  INV_X1 U23456 ( .A(n20473), .ZN(n20475) );
  AOI22_X1 U23457 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20485), .B1(
        n20484), .B2(n20685), .ZN(n20474) );
  OAI211_X1 U23458 ( .C1(n20488), .C2(n20682), .A(n20475), .B(n20474), .ZN(
        P1_U3117) );
  AOI22_X1 U23459 ( .A1(n20479), .A2(n20691), .B1(n20690), .B2(n20478), .ZN(
        n20477) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20485), .B1(
        n20484), .B2(n20628), .ZN(n20476) );
  OAI211_X1 U23461 ( .C1(n20488), .C2(n20555), .A(n20477), .B(n20476), .ZN(
        P1_U3118) );
  AOI22_X1 U23462 ( .A1(n20479), .A2(n20556), .B1(n20700), .B2(n20478), .ZN(
        n20481) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20485), .B1(
        n20484), .B2(n20701), .ZN(n20480) );
  OAI211_X1 U23464 ( .C1(n20488), .C2(n20560), .A(n20481), .B(n20480), .ZN(
        P1_U3119) );
  OAI22_X1 U23465 ( .A1(n20524), .A2(n20716), .B1(n20708), .B2(n20482), .ZN(
        n20483) );
  INV_X1 U23466 ( .A(n20483), .ZN(n20487) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20485), .B1(
        n20484), .B2(n20710), .ZN(n20486) );
  OAI211_X1 U23468 ( .C1(n20488), .C2(n20706), .A(n20487), .B(n20486), .ZN(
        P1_U3120) );
  NOR2_X1 U23469 ( .A1(n20490), .A2(n20489), .ZN(n20519) );
  AOI21_X1 U23470 ( .B1(n20492), .B2(n20491), .A(n20519), .ZN(n20495) );
  OAI22_X1 U23471 ( .A1(n20495), .A2(n20651), .B1(n20493), .B2(n20721), .ZN(
        n20518) );
  AOI22_X1 U23472 ( .A1(n20648), .A2(n20519), .B1(n20647), .B2(n20518), .ZN(
        n20502) );
  INV_X1 U23473 ( .A(n20493), .ZN(n20498) );
  OAI21_X1 U23474 ( .B1(n20494), .B2(n20651), .A(n20650), .ZN(n20496) );
  NAND2_X1 U23475 ( .A1(n20496), .A2(n20495), .ZN(n20497) );
  OAI211_X1 U23476 ( .C1(n20658), .C2(n20498), .A(n20497), .B(n20657), .ZN(
        n20521) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20660), .ZN(n20501) );
  OAI211_X1 U23478 ( .C1(n20663), .C2(n20524), .A(n20502), .B(n20501), .ZN(
        P1_U3121) );
  AOI22_X1 U23479 ( .A1(n20665), .A2(n20519), .B1(n20664), .B2(n20518), .ZN(
        n20504) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20666), .ZN(n20503) );
  OAI211_X1 U23481 ( .C1(n20669), .C2(n20524), .A(n20504), .B(n20503), .ZN(
        P1_U3122) );
  AOI22_X1 U23482 ( .A1(n20671), .A2(n20519), .B1(n20670), .B2(n20518), .ZN(
        n20506) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20672), .ZN(n20505) );
  OAI211_X1 U23484 ( .C1(n20675), .C2(n20524), .A(n20506), .B(n20505), .ZN(
        P1_U3123) );
  AOI22_X1 U23485 ( .A1(n20677), .A2(n20519), .B1(n20676), .B2(n20518), .ZN(
        n20508) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20678), .ZN(n20507) );
  OAI211_X1 U23487 ( .C1(n20681), .C2(n20524), .A(n20508), .B(n20507), .ZN(
        P1_U3124) );
  AOI22_X1 U23488 ( .A1(n20625), .A2(n20519), .B1(n20624), .B2(n20518), .ZN(
        n20511) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20509), .ZN(n20510) );
  OAI211_X1 U23490 ( .C1(n20512), .C2(n20524), .A(n20511), .B(n20510), .ZN(
        P1_U3125) );
  AOI22_X1 U23491 ( .A1(n20690), .A2(n20519), .B1(n20689), .B2(n20518), .ZN(
        n20514) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20691), .ZN(n20513) );
  OAI211_X1 U23493 ( .C1(n20696), .C2(n20524), .A(n20514), .B(n20513), .ZN(
        P1_U3126) );
  AOI22_X1 U23494 ( .A1(n20700), .A2(n20519), .B1(n20698), .B2(n20518), .ZN(
        n20516) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20556), .ZN(n20515) );
  OAI211_X1 U23496 ( .C1(n20517), .C2(n20524), .A(n20516), .B(n20515), .ZN(
        P1_U3127) );
  AOI22_X1 U23497 ( .A1(n20637), .A2(n20519), .B1(n20635), .B2(n20518), .ZN(
        n20523) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20521), .B1(
        n20564), .B2(n20520), .ZN(n20522) );
  OAI211_X1 U23499 ( .C1(n20525), .C2(n20524), .A(n20523), .B(n20522), .ZN(
        P1_U3128) );
  NAND2_X1 U23500 ( .A1(n20561), .A2(n20658), .ZN(n20528) );
  OAI21_X1 U23501 ( .B1(n20564), .B2(n20528), .A(n20527), .ZN(n20535) );
  OR2_X1 U23502 ( .A1(n13310), .A2(n9986), .ZN(n20643) );
  NOR2_X1 U23503 ( .A1(n20643), .A2(n20598), .ZN(n20532) );
  NAND3_X1 U23504 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n20531), .ZN(n20573) );
  NOR2_X1 U23505 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20573), .ZN(
        n20557) );
  AOI22_X1 U23506 ( .A1(n20648), .A2(n20557), .B1(n20592), .B2(n20660), .ZN(
        n20539) );
  INV_X1 U23507 ( .A(n20532), .ZN(n20534) );
  AOI22_X1 U23508 ( .A1(n20535), .A2(n20534), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20533), .ZN(n20536) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20608), .ZN(n20538) );
  OAI211_X1 U23510 ( .C1(n20568), .C2(n20540), .A(n20539), .B(n20538), .ZN(
        P1_U3129) );
  AOI22_X1 U23511 ( .A1(n20665), .A2(n20557), .B1(n20592), .B2(n20666), .ZN(
        n20542) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20612), .ZN(n20541) );
  OAI211_X1 U23513 ( .C1(n20568), .C2(n20543), .A(n20542), .B(n20541), .ZN(
        P1_U3130) );
  AOI22_X1 U23514 ( .A1(n20671), .A2(n20557), .B1(n20592), .B2(n20672), .ZN(
        n20545) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20616), .ZN(n20544) );
  OAI211_X1 U23516 ( .C1(n20568), .C2(n20546), .A(n20545), .B(n20544), .ZN(
        P1_U3131) );
  AOI22_X1 U23517 ( .A1(n20677), .A2(n20557), .B1(n20592), .B2(n20678), .ZN(
        n20548) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20620), .ZN(n20547) );
  OAI211_X1 U23519 ( .C1(n20568), .C2(n20549), .A(n20548), .B(n20547), .ZN(
        P1_U3132) );
  INV_X1 U23520 ( .A(n20557), .ZN(n20562) );
  OAI22_X1 U23521 ( .A1(n20683), .A2(n20562), .B1(n20688), .B2(n20561), .ZN(
        n20550) );
  INV_X1 U23522 ( .A(n20550), .ZN(n20552) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20685), .ZN(n20551) );
  OAI211_X1 U23524 ( .C1(n20568), .C2(n20682), .A(n20552), .B(n20551), .ZN(
        P1_U3133) );
  AOI22_X1 U23525 ( .A1(n20690), .A2(n20557), .B1(n20592), .B2(n20691), .ZN(
        n20554) );
  AOI22_X1 U23526 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20628), .ZN(n20553) );
  OAI211_X1 U23527 ( .C1(n20568), .C2(n20555), .A(n20554), .B(n20553), .ZN(
        P1_U3134) );
  AOI22_X1 U23528 ( .A1(n20700), .A2(n20557), .B1(n20592), .B2(n20556), .ZN(
        n20559) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20701), .ZN(n20558) );
  OAI211_X1 U23530 ( .C1(n20568), .C2(n20560), .A(n20559), .B(n20558), .ZN(
        P1_U3135) );
  OAI22_X1 U23531 ( .A1(n20708), .A2(n20562), .B1(n20716), .B2(n20561), .ZN(
        n20563) );
  INV_X1 U23532 ( .A(n20563), .ZN(n20567) );
  AOI22_X1 U23533 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20565), .B1(
        n20564), .B2(n20710), .ZN(n20566) );
  OAI211_X1 U23534 ( .C1(n20568), .C2(n20706), .A(n20567), .B(n20566), .ZN(
        P1_U3136) );
  NOR2_X1 U23535 ( .A1(n20570), .A2(n20573), .ZN(n20591) );
  INV_X1 U23536 ( .A(n20643), .ZN(n20599) );
  AOI21_X1 U23537 ( .B1(n20599), .B2(n20571), .A(n20591), .ZN(n20572) );
  OAI22_X1 U23538 ( .A1(n20572), .A2(n20651), .B1(n20573), .B2(n20721), .ZN(
        n20590) );
  AOI22_X1 U23539 ( .A1(n20648), .A2(n20591), .B1(n20647), .B2(n20590), .ZN(
        n20577) );
  INV_X1 U23540 ( .A(n20573), .ZN(n20575) );
  OAI21_X1 U23541 ( .B1(n20575), .B2(n20574), .A(n20657), .ZN(n20593) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20608), .ZN(n20576) );
  OAI211_X1 U23543 ( .C1(n20611), .C2(n20602), .A(n20577), .B(n20576), .ZN(
        P1_U3137) );
  AOI22_X1 U23544 ( .A1(n20665), .A2(n20591), .B1(n20664), .B2(n20590), .ZN(
        n20579) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20612), .ZN(n20578) );
  OAI211_X1 U23546 ( .C1(n20615), .C2(n20602), .A(n20579), .B(n20578), .ZN(
        P1_U3138) );
  AOI22_X1 U23547 ( .A1(n20671), .A2(n20591), .B1(n20670), .B2(n20590), .ZN(
        n20581) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20616), .ZN(n20580) );
  OAI211_X1 U23549 ( .C1(n20619), .C2(n20602), .A(n20581), .B(n20580), .ZN(
        P1_U3139) );
  AOI22_X1 U23550 ( .A1(n20677), .A2(n20591), .B1(n20676), .B2(n20590), .ZN(
        n20583) );
  AOI22_X1 U23551 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20620), .ZN(n20582) );
  OAI211_X1 U23552 ( .C1(n20623), .C2(n20602), .A(n20583), .B(n20582), .ZN(
        P1_U3140) );
  AOI22_X1 U23553 ( .A1(n20625), .A2(n20591), .B1(n20624), .B2(n20590), .ZN(
        n20585) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20685), .ZN(n20584) );
  OAI211_X1 U23555 ( .C1(n20688), .C2(n20602), .A(n20585), .B(n20584), .ZN(
        P1_U3141) );
  AOI22_X1 U23556 ( .A1(n20690), .A2(n20591), .B1(n20689), .B2(n20590), .ZN(
        n20587) );
  AOI22_X1 U23557 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20628), .ZN(n20586) );
  OAI211_X1 U23558 ( .C1(n20631), .C2(n20602), .A(n20587), .B(n20586), .ZN(
        P1_U3142) );
  AOI22_X1 U23559 ( .A1(n20700), .A2(n20591), .B1(n20698), .B2(n20590), .ZN(
        n20589) );
  AOI22_X1 U23560 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20701), .ZN(n20588) );
  OAI211_X1 U23561 ( .C1(n20704), .C2(n20602), .A(n20589), .B(n20588), .ZN(
        P1_U3143) );
  AOI22_X1 U23562 ( .A1(n20637), .A2(n20591), .B1(n20635), .B2(n20590), .ZN(
        n20595) );
  AOI22_X1 U23563 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20593), .B1(
        n20592), .B2(n20710), .ZN(n20594) );
  OAI211_X1 U23564 ( .C1(n20716), .C2(n20602), .A(n20595), .B(n20594), .ZN(
        P1_U3144) );
  NOR2_X1 U23565 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20597), .ZN(
        n20636) );
  NAND2_X1 U23566 ( .A1(n20599), .A2(n20598), .ZN(n20603) );
  OAI22_X1 U23567 ( .A1(n20603), .A2(n20651), .B1(n20601), .B2(n20600), .ZN(
        n20634) );
  AOI22_X1 U23568 ( .A1(n20648), .A2(n20636), .B1(n20647), .B2(n20634), .ZN(
        n20610) );
  INV_X1 U23569 ( .A(n20695), .ZN(n20711) );
  OAI21_X1 U23570 ( .B1(n20711), .B2(n20638), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20604) );
  AOI21_X1 U23571 ( .B1(n20604), .B2(n20603), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20607) );
  AOI22_X1 U23572 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23573 ( .C1(n20611), .C2(n20695), .A(n20610), .B(n20609), .ZN(
        P1_U3145) );
  AOI22_X1 U23574 ( .A1(n20665), .A2(n20636), .B1(n20664), .B2(n20634), .ZN(
        n20614) );
  AOI22_X1 U23575 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20612), .ZN(n20613) );
  OAI211_X1 U23576 ( .C1(n20615), .C2(n20695), .A(n20614), .B(n20613), .ZN(
        P1_U3146) );
  AOI22_X1 U23577 ( .A1(n20671), .A2(n20636), .B1(n20670), .B2(n20634), .ZN(
        n20618) );
  AOI22_X1 U23578 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20616), .ZN(n20617) );
  OAI211_X1 U23579 ( .C1(n20619), .C2(n20695), .A(n20618), .B(n20617), .ZN(
        P1_U3147) );
  AOI22_X1 U23580 ( .A1(n20677), .A2(n20636), .B1(n20676), .B2(n20634), .ZN(
        n20622) );
  AOI22_X1 U23581 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20620), .ZN(n20621) );
  OAI211_X1 U23582 ( .C1(n20623), .C2(n20695), .A(n20622), .B(n20621), .ZN(
        P1_U3148) );
  AOI22_X1 U23583 ( .A1(n20625), .A2(n20636), .B1(n20624), .B2(n20634), .ZN(
        n20627) );
  AOI22_X1 U23584 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20685), .ZN(n20626) );
  OAI211_X1 U23585 ( .C1(n20688), .C2(n20695), .A(n20627), .B(n20626), .ZN(
        P1_U3149) );
  AOI22_X1 U23586 ( .A1(n20690), .A2(n20636), .B1(n20689), .B2(n20634), .ZN(
        n20630) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20628), .ZN(n20629) );
  OAI211_X1 U23588 ( .C1(n20631), .C2(n20695), .A(n20630), .B(n20629), .ZN(
        P1_U3150) );
  AOI22_X1 U23589 ( .A1(n20700), .A2(n20636), .B1(n20698), .B2(n20634), .ZN(
        n20633) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20701), .ZN(n20632) );
  OAI211_X1 U23591 ( .C1(n20704), .C2(n20695), .A(n20633), .B(n20632), .ZN(
        P1_U3151) );
  AOI22_X1 U23592 ( .A1(n20637), .A2(n20636), .B1(n20635), .B2(n20634), .ZN(
        n20641) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20639), .B1(
        n20638), .B2(n20710), .ZN(n20640) );
  OAI211_X1 U23594 ( .C1(n20716), .C2(n20695), .A(n20641), .B(n20640), .ZN(
        P1_U3152) );
  INV_X1 U23595 ( .A(n20707), .ZN(n20699) );
  OR2_X1 U23596 ( .A1(n20643), .A2(n20642), .ZN(n20644) );
  NAND2_X1 U23597 ( .A1(n20644), .A2(n20707), .ZN(n20653) );
  NAND2_X1 U23598 ( .A1(n20653), .A2(n20658), .ZN(n20646) );
  NAND2_X1 U23599 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20659), .ZN(n20645) );
  AND2_X1 U23600 ( .A1(n20646), .A2(n20645), .ZN(n20705) );
  INV_X1 U23601 ( .A(n20705), .ZN(n20697) );
  AOI22_X1 U23602 ( .A1(n20648), .A2(n20699), .B1(n20647), .B2(n20697), .ZN(
        n20662) );
  INV_X1 U23603 ( .A(n20649), .ZN(n20652) );
  OAI21_X1 U23604 ( .B1(n20652), .B2(n20651), .A(n20650), .ZN(n20655) );
  INV_X1 U23605 ( .A(n20653), .ZN(n20654) );
  NAND2_X1 U23606 ( .A1(n20655), .A2(n20654), .ZN(n20656) );
  OAI211_X1 U23607 ( .C1(n20659), .C2(n20658), .A(n20657), .B(n20656), .ZN(
        n20712) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20712), .B1(
        n20692), .B2(n20660), .ZN(n20661) );
  OAI211_X1 U23609 ( .C1(n20663), .C2(n20695), .A(n20662), .B(n20661), .ZN(
        P1_U3153) );
  AOI22_X1 U23610 ( .A1(n20665), .A2(n20699), .B1(n20664), .B2(n20697), .ZN(
        n20668) );
  AOI22_X1 U23611 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20712), .B1(
        n20692), .B2(n20666), .ZN(n20667) );
  OAI211_X1 U23612 ( .C1(n20669), .C2(n20695), .A(n20668), .B(n20667), .ZN(
        P1_U3154) );
  AOI22_X1 U23613 ( .A1(n20671), .A2(n20699), .B1(n20670), .B2(n20697), .ZN(
        n20674) );
  AOI22_X1 U23614 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20712), .B1(
        n20692), .B2(n20672), .ZN(n20673) );
  OAI211_X1 U23615 ( .C1(n20675), .C2(n20695), .A(n20674), .B(n20673), .ZN(
        P1_U3155) );
  AOI22_X1 U23616 ( .A1(n20677), .A2(n20699), .B1(n20676), .B2(n20697), .ZN(
        n20680) );
  AOI22_X1 U23617 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20712), .B1(
        n20692), .B2(n20678), .ZN(n20679) );
  OAI211_X1 U23618 ( .C1(n20681), .C2(n20695), .A(n20680), .B(n20679), .ZN(
        P1_U3156) );
  OAI22_X1 U23619 ( .A1(n20683), .A2(n20707), .B1(n20682), .B2(n20705), .ZN(
        n20684) );
  INV_X1 U23620 ( .A(n20684), .ZN(n20687) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20712), .B1(
        n20711), .B2(n20685), .ZN(n20686) );
  OAI211_X1 U23622 ( .C1(n20688), .C2(n20715), .A(n20687), .B(n20686), .ZN(
        P1_U3157) );
  AOI22_X1 U23623 ( .A1(n20690), .A2(n20699), .B1(n20689), .B2(n20697), .ZN(
        n20694) );
  AOI22_X1 U23624 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20712), .B1(
        n20692), .B2(n20691), .ZN(n20693) );
  OAI211_X1 U23625 ( .C1(n20696), .C2(n20695), .A(n20694), .B(n20693), .ZN(
        P1_U3158) );
  AOI22_X1 U23626 ( .A1(n20700), .A2(n20699), .B1(n20698), .B2(n20697), .ZN(
        n20703) );
  AOI22_X1 U23627 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20712), .B1(
        n20711), .B2(n20701), .ZN(n20702) );
  OAI211_X1 U23628 ( .C1(n20704), .C2(n20715), .A(n20703), .B(n20702), .ZN(
        P1_U3159) );
  OAI22_X1 U23629 ( .A1(n20708), .A2(n20707), .B1(n20706), .B2(n20705), .ZN(
        n20709) );
  INV_X1 U23630 ( .A(n20709), .ZN(n20714) );
  AOI22_X1 U23631 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20712), .B1(
        n20711), .B2(n20710), .ZN(n20713) );
  OAI211_X1 U23632 ( .C1(n20716), .C2(n20715), .A(n20714), .B(n20713), .ZN(
        P1_U3160) );
  NOR2_X1 U23633 ( .A1(n20718), .A2(n20717), .ZN(n20722) );
  INV_X1 U23634 ( .A(n20719), .ZN(n20720) );
  OAI21_X1 U23635 ( .B1(n20722), .B2(n20721), .A(n20720), .ZN(P1_U3163) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20780), .ZN(
        P1_U3164) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20780), .ZN(
        P1_U3165) );
  AND2_X1 U23638 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20780), .ZN(
        P1_U3166) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20780), .ZN(
        P1_U3167) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20780), .ZN(
        P1_U3168) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20780), .ZN(
        P1_U3169) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20780), .ZN(
        P1_U3170) );
  AND2_X1 U23643 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20780), .ZN(
        P1_U3171) );
  AND2_X1 U23644 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20780), .ZN(
        P1_U3172) );
  AND2_X1 U23645 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20780), .ZN(
        P1_U3173) );
  AND2_X1 U23646 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20780), .ZN(
        P1_U3174) );
  AND2_X1 U23647 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20780), .ZN(
        P1_U3175) );
  AND2_X1 U23648 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20780), .ZN(
        P1_U3176) );
  AND2_X1 U23649 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20780), .ZN(
        P1_U3177) );
  AND2_X1 U23650 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20780), .ZN(
        P1_U3178) );
  AND2_X1 U23651 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20780), .ZN(
        P1_U3179) );
  AND2_X1 U23652 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20780), .ZN(
        P1_U3180) );
  AND2_X1 U23653 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20780), .ZN(
        P1_U3181) );
  AND2_X1 U23654 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20780), .ZN(
        P1_U3182) );
  AND2_X1 U23655 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20780), .ZN(
        P1_U3183) );
  AND2_X1 U23656 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20780), .ZN(
        P1_U3184) );
  AND2_X1 U23657 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20780), .ZN(
        P1_U3185) );
  AND2_X1 U23658 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20780), .ZN(P1_U3186) );
  AND2_X1 U23659 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20780), .ZN(P1_U3187) );
  AND2_X1 U23660 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20780), .ZN(P1_U3188) );
  AND2_X1 U23661 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20780), .ZN(P1_U3189) );
  AND2_X1 U23662 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20780), .ZN(P1_U3190) );
  AND2_X1 U23663 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20780), .ZN(P1_U3191) );
  AND2_X1 U23664 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20780), .ZN(P1_U3192) );
  AND2_X1 U23665 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20780), .ZN(P1_U3193) );
  AND2_X1 U23666 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20723), .ZN(n20734) );
  INV_X1 U23667 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20884) );
  OAI22_X1 U23668 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n21174), .B1(n20728), 
        .B2(n20724), .ZN(n20725) );
  NOR3_X1 U23669 ( .A1(n20726), .A2(n20884), .A3(n20725), .ZN(n20727) );
  OAI22_X1 U23670 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20734), .B1(n20772), 
        .B2(n20727), .ZN(P1_U3194) );
  NOR2_X1 U23671 ( .A1(n20735), .A2(n20728), .ZN(n20730) );
  NOR2_X1 U23672 ( .A1(n11622), .A2(n20884), .ZN(n20729) );
  OAI22_X1 U23673 ( .A1(n20730), .A2(n21174), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20729), .ZN(n20733) );
  OAI211_X1 U23674 ( .C1(NA), .C2(n20800), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20735), .ZN(n20731) );
  OAI211_X1 U23675 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20884), .A(HOLD), .B(
        n20731), .ZN(n20732) );
  OAI22_X1 U23676 ( .A1(n20734), .A2(n20733), .B1(n11622), .B2(n20732), .ZN(
        P1_U3196) );
  AND2_X1 U23677 ( .A1(n20772), .A2(n20735), .ZN(n20759) );
  INV_X1 U23678 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20736) );
  NAND2_X1 U23679 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20772), .ZN(n20774) );
  INV_X1 U23680 ( .A(n20774), .ZN(n20758) );
  OAI222_X1 U23681 ( .A1(n9822), .A2(n21151), .B1(n20736), .B2(n20772), .C1(
        n20904), .C2(n20771), .ZN(P1_U3197) );
  INV_X1 U23682 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20737) );
  INV_X1 U23683 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20934) );
  OAI222_X1 U23684 ( .A1(n20771), .A2(n21151), .B1(n20737), .B2(n20772), .C1(
        n20934), .C2(n9822), .ZN(P1_U3198) );
  INV_X1 U23685 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n21170) );
  OAI222_X1 U23686 ( .A1(n20774), .A2(n20934), .B1(n20738), .B2(n20772), .C1(
        n21170), .C2(n9822), .ZN(P1_U3199) );
  INV_X1 U23687 ( .A(P1_ADDRESS_REG_3__SCAN_IN), .ZN(n20739) );
  OAI222_X1 U23688 ( .A1(n9822), .A2(n20905), .B1(n20739), .B2(n20772), .C1(
        n21170), .C2(n20771), .ZN(P1_U3200) );
  INV_X1 U23689 ( .A(P1_ADDRESS_REG_4__SCAN_IN), .ZN(n20740) );
  OAI222_X1 U23690 ( .A1(n9822), .A2(n21141), .B1(n20740), .B2(n20772), .C1(
        n20905), .C2(n20771), .ZN(P1_U3201) );
  INV_X1 U23691 ( .A(P1_ADDRESS_REG_5__SCAN_IN), .ZN(n20741) );
  OAI222_X1 U23692 ( .A1(n20774), .A2(n21141), .B1(n20741), .B2(n20772), .C1(
        n21008), .C2(n9822), .ZN(P1_U3202) );
  AOI22_X1 U23693 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20808), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20759), .ZN(n20742) );
  OAI21_X1 U23694 ( .B1(n21008), .B2(n20771), .A(n20742), .ZN(P1_U3203) );
  AOI22_X1 U23695 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20808), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20758), .ZN(n20743) );
  OAI21_X1 U23696 ( .B1(n21029), .B2(n9822), .A(n20743), .ZN(P1_U3204) );
  INV_X1 U23697 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21032) );
  INV_X1 U23698 ( .A(P1_ADDRESS_REG_8__SCAN_IN), .ZN(n20744) );
  OAI222_X1 U23699 ( .A1(n9822), .A2(n21032), .B1(n20744), .B2(n20772), .C1(
        n21029), .C2(n20771), .ZN(P1_U3205) );
  INV_X1 U23700 ( .A(P1_ADDRESS_REG_9__SCAN_IN), .ZN(n20745) );
  OAI222_X1 U23701 ( .A1(n9822), .A2(n20987), .B1(n20745), .B2(n20772), .C1(
        n21032), .C2(n20771), .ZN(P1_U3206) );
  INV_X1 U23702 ( .A(P1_ADDRESS_REG_10__SCAN_IN), .ZN(n20746) );
  OAI222_X1 U23703 ( .A1(n9822), .A2(n21154), .B1(n20746), .B2(n20772), .C1(
        n20987), .C2(n20771), .ZN(P1_U3207) );
  INV_X1 U23704 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n20747) );
  OAI222_X1 U23705 ( .A1(n20774), .A2(n21154), .B1(n20747), .B2(n20772), .C1(
        n21138), .C2(n9822), .ZN(P1_U3208) );
  INV_X1 U23706 ( .A(P1_ADDRESS_REG_12__SCAN_IN), .ZN(n20748) );
  INV_X1 U23707 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20917) );
  OAI222_X1 U23708 ( .A1(n20771), .A2(n21138), .B1(n20748), .B2(n20772), .C1(
        n20917), .C2(n9822), .ZN(P1_U3209) );
  INV_X1 U23709 ( .A(P1_ADDRESS_REG_13__SCAN_IN), .ZN(n20749) );
  OAI222_X1 U23710 ( .A1(n20771), .A2(n20917), .B1(n20749), .B2(n20772), .C1(
        n21124), .C2(n9822), .ZN(P1_U3210) );
  INV_X1 U23711 ( .A(P1_ADDRESS_REG_14__SCAN_IN), .ZN(n20750) );
  OAI222_X1 U23712 ( .A1(n9822), .A2(n20752), .B1(n20750), .B2(n20772), .C1(
        n21124), .C2(n20771), .ZN(P1_U3211) );
  INV_X1 U23713 ( .A(P1_ADDRESS_REG_15__SCAN_IN), .ZN(n20751) );
  OAI222_X1 U23714 ( .A1(n20771), .A2(n20752), .B1(n20751), .B2(n20772), .C1(
        n20754), .C2(n9822), .ZN(P1_U3212) );
  INV_X1 U23715 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20753) );
  OAI222_X1 U23716 ( .A1(n20771), .A2(n20754), .B1(n20753), .B2(n20772), .C1(
        n20933), .C2(n9822), .ZN(P1_U3213) );
  INV_X1 U23717 ( .A(P1_ADDRESS_REG_17__SCAN_IN), .ZN(n20755) );
  OAI222_X1 U23718 ( .A1(n20774), .A2(n20933), .B1(n20755), .B2(n20772), .C1(
        n20891), .C2(n9822), .ZN(P1_U3214) );
  INV_X1 U23719 ( .A(P1_ADDRESS_REG_18__SCAN_IN), .ZN(n20756) );
  OAI222_X1 U23720 ( .A1(n9822), .A2(n21026), .B1(n20756), .B2(n20772), .C1(
        n20891), .C2(n20771), .ZN(P1_U3215) );
  AOI222_X1 U23721 ( .A1(n20758), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20808), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20759), .ZN(n20757) );
  INV_X1 U23722 ( .A(n20757), .ZN(P1_U3216) );
  AOI222_X1 U23723 ( .A1(n20759), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20808), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20758), .ZN(n20760) );
  INV_X1 U23724 ( .A(n20760), .ZN(P1_U3217) );
  INV_X1 U23725 ( .A(P1_ADDRESS_REG_21__SCAN_IN), .ZN(n20761) );
  OAI222_X1 U23726 ( .A1(n20774), .A2(n21144), .B1(n20761), .B2(n20772), .C1(
        n20763), .C2(n9822), .ZN(P1_U3218) );
  INV_X1 U23727 ( .A(P1_ADDRESS_REG_22__SCAN_IN), .ZN(n20762) );
  INV_X1 U23728 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21169) );
  OAI222_X1 U23729 ( .A1(n20774), .A2(n20763), .B1(n20762), .B2(n20772), .C1(
        n21169), .C2(n9822), .ZN(P1_U3219) );
  INV_X1 U23730 ( .A(P1_ADDRESS_REG_23__SCAN_IN), .ZN(n20764) );
  OAI222_X1 U23731 ( .A1(n20771), .A2(n21169), .B1(n20764), .B2(n20772), .C1(
        n21140), .C2(n9822), .ZN(P1_U3220) );
  INV_X1 U23732 ( .A(P1_ADDRESS_REG_24__SCAN_IN), .ZN(n20765) );
  OAI222_X1 U23733 ( .A1(n20774), .A2(n21140), .B1(n20765), .B2(n20772), .C1(
        n14344), .C2(n9822), .ZN(P1_U3221) );
  INV_X1 U23734 ( .A(P1_ADDRESS_REG_25__SCAN_IN), .ZN(n20766) );
  OAI222_X1 U23735 ( .A1(n20771), .A2(n14344), .B1(n20766), .B2(n20772), .C1(
        n21027), .C2(n9822), .ZN(P1_U3222) );
  INV_X1 U23736 ( .A(P1_ADDRESS_REG_26__SCAN_IN), .ZN(n20767) );
  OAI222_X1 U23737 ( .A1(n20771), .A2(n21027), .B1(n20767), .B2(n20772), .C1(
        n14523), .C2(n9822), .ZN(P1_U3223) );
  INV_X1 U23738 ( .A(P1_ADDRESS_REG_27__SCAN_IN), .ZN(n20768) );
  INV_X1 U23739 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20770) );
  OAI222_X1 U23740 ( .A1(n20771), .A2(n14523), .B1(n20768), .B2(n20772), .C1(
        n20770), .C2(n9822), .ZN(P1_U3224) );
  INV_X1 U23741 ( .A(P1_ADDRESS_REG_28__SCAN_IN), .ZN(n20769) );
  OAI222_X1 U23742 ( .A1(n20771), .A2(n20770), .B1(n20769), .B2(n20772), .C1(
        n14510), .C2(n9822), .ZN(P1_U3225) );
  INV_X1 U23743 ( .A(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20773) );
  OAI222_X1 U23744 ( .A1(n20774), .A2(n14510), .B1(n20773), .B2(n20772), .C1(
        n20965), .C2(n9822), .ZN(P1_U3226) );
  INV_X1 U23745 ( .A(P1_BE_N_REG_3__SCAN_IN), .ZN(n20775) );
  AOI22_X1 U23746 ( .A1(n20772), .A2(n20913), .B1(n20775), .B2(n20808), .ZN(
        P1_U3458) );
  INV_X1 U23747 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20794) );
  INV_X1 U23748 ( .A(P1_BE_N_REG_2__SCAN_IN), .ZN(n20776) );
  AOI22_X1 U23749 ( .A1(n20772), .A2(n20794), .B1(n20776), .B2(n20808), .ZN(
        P1_U3459) );
  INV_X1 U23750 ( .A(P1_BE_N_REG_1__SCAN_IN), .ZN(n20777) );
  AOI22_X1 U23751 ( .A1(n20772), .A2(n20989), .B1(n20777), .B2(n20808), .ZN(
        P1_U3460) );
  INV_X1 U23752 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21153) );
  INV_X1 U23753 ( .A(P1_BE_N_REG_0__SCAN_IN), .ZN(n20778) );
  AOI22_X1 U23754 ( .A1(n20772), .A2(n21153), .B1(n20778), .B2(n20808), .ZN(
        P1_U3461) );
  INV_X1 U23755 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20781) );
  INV_X1 U23756 ( .A(n20782), .ZN(n20779) );
  AOI21_X1 U23757 ( .B1(n20781), .B2(n20780), .A(n20779), .ZN(P1_U3464) );
  OAI21_X1 U23758 ( .B1(n20784), .B2(n20783), .A(n20782), .ZN(P1_U3465) );
  INV_X1 U23759 ( .A(n20785), .ZN(n20787) );
  OAI22_X1 U23760 ( .A1(n20789), .A2(n20788), .B1(n20787), .B2(n20786), .ZN(
        n20791) );
  MUX2_X1 U23761 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20791), .S(
        n20790), .Z(P1_U3469) );
  AOI21_X1 U23762 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20792) );
  AOI22_X1 U23763 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20792), .B2(n20904), .ZN(n20795) );
  AOI22_X1 U23764 ( .A1(n20797), .A2(n20795), .B1(n20794), .B2(n20793), .ZN(
        P1_U3481) );
  OAI21_X1 U23765 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20797), .ZN(n20796) );
  OAI21_X1 U23766 ( .B1(n20797), .B2(n21153), .A(n20796), .ZN(P1_U3482) );
  AOI22_X1 U23767 ( .A1(n20772), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20968), 
        .B2(n20808), .ZN(P1_U3483) );
  AOI211_X1 U23768 ( .C1(n20801), .C2(n20800), .A(n20799), .B(n20798), .ZN(
        n20807) );
  OAI21_X1 U23769 ( .B1(n10240), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20802) );
  OAI21_X1 U23770 ( .B1(n20803), .B2(n20802), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n20806) );
  NOR2_X1 U23771 ( .A1(n20807), .A2(n20804), .ZN(n20805) );
  AOI22_X1 U23772 ( .A1(n20884), .A2(n20807), .B1(n20806), .B2(n20805), .ZN(
        P1_U3485) );
  INV_X1 U23773 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20809) );
  AOI22_X1 U23774 ( .A1(n20772), .A2(n20809), .B1(n20947), .B2(n20808), .ZN(
        P1_U3486) );
  OAI22_X1 U23775 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput_g126), .B1(
        P1_EBX_REG_2__SCAN_IN), .B2(keyinput_g113), .ZN(n20810) );
  AOI221_X1 U23776 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput_g126), .C1(
        keyinput_g113), .C2(P1_EBX_REG_2__SCAN_IN), .A(n20810), .ZN(n20817) );
  OAI22_X1 U23777 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_g103), .B1(
        DATAI_27_), .B2(keyinput_g5), .ZN(n20811) );
  AOI221_X1 U23778 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_g103), .C1(
        keyinput_g5), .C2(DATAI_27_), .A(n20811), .ZN(n20816) );
  OAI22_X1 U23779 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput_g125), .B1(
        keyinput_g86), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n20812) );
  AOI221_X1 U23780 ( .B1(P1_EAX_REG_22__SCAN_IN), .B2(keyinput_g125), .C1(
        P1_EBX_REG_29__SCAN_IN), .C2(keyinput_g86), .A(n20812), .ZN(n20815) );
  OAI22_X1 U23781 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(keyinput_g102), .B1(
        keyinput_g30), .B2(DATAI_2_), .ZN(n20813) );
  AOI221_X1 U23782 ( .B1(P1_EBX_REG_13__SCAN_IN), .B2(keyinput_g102), .C1(
        DATAI_2_), .C2(keyinput_g30), .A(n20813), .ZN(n20814) );
  NAND4_X1 U23783 ( .A1(n20817), .A2(n20816), .A3(n20815), .A4(n20814), .ZN(
        n20845) );
  OAI22_X1 U23784 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(keyinput_g0), .B2(
        P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n20818) );
  AOI221_X1 U23785 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_g0), .A(n20818), .ZN(n20825)
         );
  OAI22_X1 U23786 ( .A1(P1_EAX_REG_26__SCAN_IN), .A2(keyinput_g121), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .ZN(n20819) );
  AOI221_X1 U23787 ( .B1(P1_EAX_REG_26__SCAN_IN), .B2(keyinput_g121), .C1(
        keyinput_g62), .C2(P1_REIP_REG_21__SCAN_IN), .A(n20819), .ZN(n20824)
         );
  OAI22_X1 U23788 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_g88), .B1(
        keyinput_g104), .B2(P1_EBX_REG_11__SCAN_IN), .ZN(n20820) );
  AOI221_X1 U23789 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_g88), .C1(
        P1_EBX_REG_11__SCAN_IN), .C2(keyinput_g104), .A(n20820), .ZN(n20823)
         );
  OAI22_X1 U23790 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput_g95), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(keyinput_g66), .ZN(n20821) );
  AOI221_X1 U23791 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput_g95), .C1(
        keyinput_g66), .C2(P1_REIP_REG_17__SCAN_IN), .A(n20821), .ZN(n20822)
         );
  NAND4_X1 U23792 ( .A1(n20825), .A2(n20824), .A3(n20823), .A4(n20822), .ZN(
        n20844) );
  OAI22_X1 U23793 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_g44), .B1(
        READY2), .B2(keyinput_g37), .ZN(n20826) );
  AOI221_X1 U23794 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_g44), .C1(
        keyinput_g37), .C2(READY2), .A(n20826), .ZN(n20833) );
  OAI22_X1 U23795 ( .A1(P1_EAX_REG_24__SCAN_IN), .A2(keyinput_g123), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_g108), .ZN(n20827) );
  AOI221_X1 U23796 ( .B1(P1_EAX_REG_24__SCAN_IN), .B2(keyinput_g123), .C1(
        keyinput_g108), .C2(P1_EBX_REG_7__SCAN_IN), .A(n20827), .ZN(n20832) );
  OAI22_X1 U23797 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_g63), .B1(
        keyinput_g2), .B2(DATAI_30_), .ZN(n20828) );
  AOI221_X1 U23798 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_g63), .C1(
        DATAI_30_), .C2(keyinput_g2), .A(n20828), .ZN(n20831) );
  OAI22_X1 U23799 ( .A1(READY1), .A2(keyinput_g36), .B1(keyinput_g112), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n20829) );
  AOI221_X1 U23800 ( .B1(READY1), .B2(keyinput_g36), .C1(P1_EBX_REG_3__SCAN_IN), .C2(keyinput_g112), .A(n20829), .ZN(n20830) );
  NAND4_X1 U23801 ( .A1(n20833), .A2(n20832), .A3(n20831), .A4(n20830), .ZN(
        n20843) );
  OAI22_X1 U23802 ( .A1(DATAI_24_), .A2(keyinput_g8), .B1(keyinput_g12), .B2(
        DATAI_20_), .ZN(n20834) );
  AOI221_X1 U23803 ( .B1(DATAI_24_), .B2(keyinput_g8), .C1(DATAI_20_), .C2(
        keyinput_g12), .A(n20834), .ZN(n20841) );
  OAI22_X1 U23804 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput_g55), .B1(
        keyinput_g31), .B2(DATAI_1_), .ZN(n20835) );
  AOI221_X1 U23805 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .C1(
        DATAI_1_), .C2(keyinput_g31), .A(n20835), .ZN(n20840) );
  OAI22_X1 U23806 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(keyinput_g77), .B1(
        keyinput_g33), .B2(HOLD), .ZN(n20836) );
  AOI221_X1 U23807 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(keyinput_g77), .C1(HOLD), 
        .C2(keyinput_g33), .A(n20836), .ZN(n20839) );
  OAI22_X1 U23808 ( .A1(DATAI_29_), .A2(keyinput_g3), .B1(keyinput_g48), .B2(
        P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20837) );
  AOI221_X1 U23809 ( .B1(DATAI_29_), .B2(keyinput_g3), .C1(
        P1_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput_g48), .A(n20837), .ZN(
        n20838) );
  NAND4_X1 U23810 ( .A1(n20841), .A2(n20840), .A3(n20839), .A4(n20838), .ZN(
        n20842) );
  NOR4_X1 U23811 ( .A1(n20845), .A2(n20844), .A3(n20843), .A4(n20842), .ZN(
        n21197) );
  OAI22_X1 U23812 ( .A1(P1_EBX_REG_31__SCAN_IN), .A2(keyinput_g84), .B1(
        DATAI_25_), .B2(keyinput_g7), .ZN(n20846) );
  AOI221_X1 U23813 ( .B1(P1_EBX_REG_31__SCAN_IN), .B2(keyinput_g84), .C1(
        keyinput_g7), .C2(DATAI_25_), .A(n20846), .ZN(n20853) );
  OAI22_X1 U23814 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_g122), .B1(
        keyinput_g67), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n20847) );
  AOI221_X1 U23815 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_g122), .C1(
        P1_REIP_REG_16__SCAN_IN), .C2(keyinput_g67), .A(n20847), .ZN(n20852)
         );
  OAI22_X1 U23816 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_g116), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n20848) );
  AOI221_X1 U23817 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_g116), .C1(
        keyinput_g60), .C2(P1_REIP_REG_23__SCAN_IN), .A(n20848), .ZN(n20851)
         );
  OAI22_X1 U23818 ( .A1(DATAI_21_), .A2(keyinput_g11), .B1(
        P1_ADS_N_REG_SCAN_IN), .B2(keyinput_g39), .ZN(n20849) );
  AOI221_X1 U23819 ( .B1(DATAI_21_), .B2(keyinput_g11), .C1(keyinput_g39), 
        .C2(P1_ADS_N_REG_SCAN_IN), .A(n20849), .ZN(n20850) );
  NAND4_X1 U23820 ( .A1(n20853), .A2(n20852), .A3(n20851), .A4(n20850), .ZN(
        n20981) );
  OAI22_X1 U23821 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(keyinput_g75), .B1(
        keyinput_g6), .B2(DATAI_26_), .ZN(n20854) );
  AOI221_X1 U23822 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(keyinput_g75), .C1(
        DATAI_26_), .C2(keyinput_g6), .A(n20854), .ZN(n20879) );
  OAI22_X1 U23823 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput_g127), .B1(NA), 
        .B2(keyinput_g34), .ZN(n20855) );
  AOI221_X1 U23824 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput_g127), .C1(
        keyinput_g34), .C2(NA), .A(n20855), .ZN(n20858) );
  OAI22_X1 U23825 ( .A1(P1_EBX_REG_21__SCAN_IN), .A2(keyinput_g94), .B1(
        DATAI_0_), .B2(keyinput_g32), .ZN(n20856) );
  AOI221_X1 U23826 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(keyinput_g94), .C1(
        keyinput_g32), .C2(DATAI_0_), .A(n20856), .ZN(n20857) );
  OAI211_X1 U23827 ( .C1(n21033), .C2(keyinput_g14), .A(n20858), .B(n20857), 
        .ZN(n20859) );
  AOI21_X1 U23828 ( .B1(n21033), .B2(keyinput_g14), .A(n20859), .ZN(n20878) );
  AOI22_X1 U23829 ( .A1(P1_EBX_REG_30__SCAN_IN), .A2(keyinput_g85), .B1(
        P1_EBX_REG_25__SCAN_IN), .B2(keyinput_g90), .ZN(n20860) );
  OAI221_X1 U23830 ( .B1(P1_EBX_REG_30__SCAN_IN), .B2(keyinput_g85), .C1(
        P1_EBX_REG_25__SCAN_IN), .C2(keyinput_g90), .A(n20860), .ZN(n20867) );
  AOI22_X1 U23831 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_g40), .ZN(n20861) );
  OAI221_X1 U23832 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_g40), .A(n20861), .ZN(
        n20866) );
  AOI22_X1 U23833 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_g83), .B1(
        DATAI_15_), .B2(keyinput_g17), .ZN(n20862) );
  OAI221_X1 U23834 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_g83), .C1(
        DATAI_15_), .C2(keyinput_g17), .A(n20862), .ZN(n20865) );
  AOI22_X1 U23835 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_g45), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_g118), .ZN(n20863) );
  OAI221_X1 U23836 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_g118), .A(n20863), .ZN(n20864)
         );
  NOR4_X1 U23837 ( .A1(n20867), .A2(n20866), .A3(n20865), .A4(n20864), .ZN(
        n20877) );
  AOI22_X1 U23838 ( .A1(P1_EBX_REG_6__SCAN_IN), .A2(keyinput_g109), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(keyinput_g119), .ZN(n20868) );
  OAI221_X1 U23839 ( .B1(P1_EBX_REG_6__SCAN_IN), .B2(keyinput_g109), .C1(
        P1_EAX_REG_28__SCAN_IN), .C2(keyinput_g119), .A(n20868), .ZN(n20875)
         );
  AOI22_X1 U23840 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(keyinput_g81), .ZN(n20869) );
  OAI221_X1 U23841 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(
        P1_REIP_REG_2__SCAN_IN), .C2(keyinput_g81), .A(n20869), .ZN(n20874) );
  AOI22_X1 U23842 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(keyinput_g79), .B1(
        P1_REIP_REG_27__SCAN_IN), .B2(keyinput_g56), .ZN(n20870) );
  OAI221_X1 U23843 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(keyinput_g79), .C1(
        P1_REIP_REG_27__SCAN_IN), .C2(keyinput_g56), .A(n20870), .ZN(n20873)
         );
  AOI22_X1 U23844 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(
        P1_EBX_REG_1__SCAN_IN), .B2(keyinput_g114), .ZN(n20871) );
  OAI221_X1 U23845 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(
        P1_EBX_REG_1__SCAN_IN), .C2(keyinput_g114), .A(n20871), .ZN(n20872) );
  NOR4_X1 U23846 ( .A1(n20875), .A2(n20874), .A3(n20873), .A4(n20872), .ZN(
        n20876) );
  NAND4_X1 U23847 ( .A1(n20879), .A2(n20878), .A3(n20877), .A4(n20876), .ZN(
        n20980) );
  AOI22_X1 U23848 ( .A1(DATAI_28_), .A2(keyinput_g4), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n20880) );
  OAI221_X1 U23849 ( .B1(DATAI_28_), .B2(keyinput_g4), .C1(
        P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n20880), .ZN(n20888)
         );
  AOI22_X1 U23850 ( .A1(n21008), .A2(keyinput_g76), .B1(n21144), .B2(
        keyinput_g61), .ZN(n20881) );
  OAI221_X1 U23851 ( .B1(n21008), .B2(keyinput_g76), .C1(n21144), .C2(
        keyinput_g61), .A(n20881), .ZN(n20887) );
  AOI22_X1 U23852 ( .A1(n21140), .A2(keyinput_g58), .B1(n21009), .B2(
        keyinput_g100), .ZN(n20882) );
  OAI221_X1 U23853 ( .B1(n21140), .B2(keyinput_g58), .C1(n21009), .C2(
        keyinput_g100), .A(n20882), .ZN(n20886) );
  AOI22_X1 U23854 ( .A1(n14344), .A2(keyinput_g57), .B1(keyinput_g43), .B2(
        n20884), .ZN(n20883) );
  OAI221_X1 U23855 ( .B1(n14344), .B2(keyinput_g57), .C1(n20884), .C2(
        keyinput_g43), .A(n20883), .ZN(n20885) );
  NOR4_X1 U23856 ( .A1(n20888), .A2(n20887), .A3(n20886), .A4(n20885), .ZN(
        n20927) );
  AOI22_X1 U23857 ( .A1(n20891), .A2(keyinput_g64), .B1(n20890), .B2(
        keyinput_g120), .ZN(n20889) );
  OAI221_X1 U23858 ( .B1(n20891), .B2(keyinput_g64), .C1(n20890), .C2(
        keyinput_g120), .A(n20889), .ZN(n20900) );
  AOI22_X1 U23859 ( .A1(n21135), .A2(keyinput_g16), .B1(n14510), .B2(
        keyinput_g53), .ZN(n20892) );
  OAI221_X1 U23860 ( .B1(n21135), .B2(keyinput_g16), .C1(n14510), .C2(
        keyinput_g53), .A(n20892), .ZN(n20899) );
  AOI22_X1 U23861 ( .A1(n20894), .A2(keyinput_g27), .B1(n20983), .B2(
        keyinput_g26), .ZN(n20893) );
  OAI221_X1 U23862 ( .B1(n20894), .B2(keyinput_g27), .C1(n20983), .C2(
        keyinput_g26), .A(n20893), .ZN(n20898) );
  AOI22_X1 U23863 ( .A1(n20999), .A2(keyinput_g10), .B1(n20896), .B2(
        keyinput_g18), .ZN(n20895) );
  OAI221_X1 U23864 ( .B1(n20999), .B2(keyinput_g10), .C1(n20896), .C2(
        keyinput_g18), .A(n20895), .ZN(n20897) );
  NOR4_X1 U23865 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20926) );
  AOI22_X1 U23866 ( .A1(n21134), .A2(keyinput_g99), .B1(keyinput_g9), .B2(
        n21122), .ZN(n20901) );
  OAI221_X1 U23867 ( .B1(n21134), .B2(keyinput_g99), .C1(n21122), .C2(
        keyinput_g9), .A(n20901), .ZN(n20911) );
  AOI22_X1 U23868 ( .A1(n21138), .A2(keyinput_g70), .B1(n21167), .B2(
        keyinput_g89), .ZN(n20902) );
  OAI221_X1 U23869 ( .B1(n21138), .B2(keyinput_g70), .C1(n21167), .C2(
        keyinput_g89), .A(n20902), .ZN(n20910) );
  AOI22_X1 U23870 ( .A1(n20905), .A2(keyinput_g78), .B1(n20904), .B2(
        keyinput_g82), .ZN(n20903) );
  OAI221_X1 U23871 ( .B1(n20905), .B2(keyinput_g78), .C1(n20904), .C2(
        keyinput_g82), .A(n20903), .ZN(n20909) );
  AOI22_X1 U23872 ( .A1(n20907), .A2(keyinput_g101), .B1(keyinput_g73), .B2(
        n21032), .ZN(n20906) );
  OAI221_X1 U23873 ( .B1(n20907), .B2(keyinput_g101), .C1(n21032), .C2(
        keyinput_g73), .A(n20906), .ZN(n20908) );
  NOR4_X1 U23874 ( .A1(n20911), .A2(n20910), .A3(n20909), .A4(n20908), .ZN(
        n20925) );
  AOI22_X1 U23875 ( .A1(n20913), .A2(keyinput_g51), .B1(n21169), .B2(
        keyinput_g59), .ZN(n20912) );
  OAI221_X1 U23876 ( .B1(n20913), .B2(keyinput_g51), .C1(n21169), .C2(
        keyinput_g59), .A(n20912), .ZN(n20923) );
  INV_X1 U23877 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n20915) );
  AOI22_X1 U23878 ( .A1(n20915), .A2(keyinput_g38), .B1(keyinput_g49), .B2(
        n20989), .ZN(n20914) );
  OAI221_X1 U23879 ( .B1(n20915), .B2(keyinput_g38), .C1(n20989), .C2(
        keyinput_g49), .A(n20914), .ZN(n20922) );
  AOI22_X1 U23880 ( .A1(n21000), .A2(keyinput_g106), .B1(keyinput_g69), .B2(
        n20917), .ZN(n20916) );
  OAI221_X1 U23881 ( .B1(n21000), .B2(keyinput_g106), .C1(n20917), .C2(
        keyinput_g69), .A(n20916), .ZN(n20921) );
  AOI22_X1 U23882 ( .A1(n20919), .A2(keyinput_g21), .B1(n21154), .B2(
        keyinput_g71), .ZN(n20918) );
  OAI221_X1 U23883 ( .B1(n20919), .B2(keyinput_g21), .C1(n21154), .C2(
        keyinput_g71), .A(n20918), .ZN(n20920) );
  NOR4_X1 U23884 ( .A1(n20923), .A2(n20922), .A3(n20921), .A4(n20920), .ZN(
        n20924) );
  NAND4_X1 U23885 ( .A1(n20927), .A2(n20926), .A3(n20925), .A4(n20924), .ZN(
        n20979) );
  AOI22_X1 U23886 ( .A1(n21036), .A2(keyinput_g124), .B1(keyinput_g97), .B2(
        n21059), .ZN(n20928) );
  OAI221_X1 U23887 ( .B1(n21036), .B2(keyinput_g124), .C1(n21059), .C2(
        keyinput_g97), .A(n20928), .ZN(n20940) );
  AOI22_X1 U23888 ( .A1(n20931), .A2(keyinput_g28), .B1(keyinput_g42), .B2(
        n20930), .ZN(n20929) );
  OAI221_X1 U23889 ( .B1(n20931), .B2(keyinput_g28), .C1(n20930), .C2(
        keyinput_g42), .A(n20929), .ZN(n20939) );
  AOI22_X1 U23890 ( .A1(n20934), .A2(keyinput_g80), .B1(n20933), .B2(
        keyinput_g65), .ZN(n20932) );
  OAI221_X1 U23891 ( .B1(n20934), .B2(keyinput_g80), .C1(n20933), .C2(
        keyinput_g65), .A(n20932), .ZN(n20938) );
  AOI22_X1 U23892 ( .A1(n20936), .A2(keyinput_g117), .B1(keyinput_g96), .B2(
        n21125), .ZN(n20935) );
  OAI221_X1 U23893 ( .B1(n20936), .B2(keyinput_g117), .C1(n21125), .C2(
        keyinput_g96), .A(n20935), .ZN(n20937) );
  NOR4_X1 U23894 ( .A1(n20940), .A2(n20939), .A3(n20938), .A4(n20937), .ZN(
        n20977) );
  AOI22_X1 U23895 ( .A1(n13755), .A2(keyinput_g105), .B1(n21157), .B2(
        keyinput_g110), .ZN(n20941) );
  OAI221_X1 U23896 ( .B1(n13755), .B2(keyinput_g105), .C1(n21157), .C2(
        keyinput_g110), .A(n20941), .ZN(n20951) );
  AOI22_X1 U23897 ( .A1(n20943), .A2(keyinput_g35), .B1(n21029), .B2(
        keyinput_g74), .ZN(n20942) );
  OAI221_X1 U23898 ( .B1(n20943), .B2(keyinput_g35), .C1(n21029), .C2(
        keyinput_g74), .A(n20942), .ZN(n20950) );
  AOI22_X1 U23899 ( .A1(n20945), .A2(keyinput_g87), .B1(keyinput_g92), .B2(
        n21020), .ZN(n20944) );
  OAI221_X1 U23900 ( .B1(n20945), .B2(keyinput_g87), .C1(n21020), .C2(
        keyinput_g92), .A(n20944), .ZN(n20949) );
  AOI22_X1 U23901 ( .A1(n20993), .A2(keyinput_g19), .B1(keyinput_g41), .B2(
        n20947), .ZN(n20946) );
  OAI221_X1 U23902 ( .B1(n20993), .B2(keyinput_g19), .C1(n20947), .C2(
        keyinput_g41), .A(n20946), .ZN(n20948) );
  NOR4_X1 U23903 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20976) );
  INV_X1 U23904 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n21150) );
  AOI22_X1 U23905 ( .A1(n21156), .A2(keyinput_g98), .B1(keyinput_g111), .B2(
        n21150), .ZN(n20952) );
  OAI221_X1 U23906 ( .B1(n21156), .B2(keyinput_g98), .C1(n21150), .C2(
        keyinput_g111), .A(n20952), .ZN(n20963) );
  INV_X1 U23907 ( .A(DATAI_8_), .ZN(n20954) );
  INV_X1 U23908 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21019) );
  AOI22_X1 U23909 ( .A1(n20954), .A2(keyinput_g24), .B1(n21019), .B2(
        keyinput_g107), .ZN(n20953) );
  OAI221_X1 U23910 ( .B1(n20954), .B2(keyinput_g24), .C1(n21019), .C2(
        keyinput_g107), .A(n20953), .ZN(n20962) );
  AOI22_X1 U23911 ( .A1(n20957), .A2(keyinput_g1), .B1(keyinput_g25), .B2(
        n20956), .ZN(n20955) );
  OAI221_X1 U23912 ( .B1(n20957), .B2(keyinput_g1), .C1(n20956), .C2(
        keyinput_g25), .A(n20955), .ZN(n20961) );
  AOI22_X1 U23913 ( .A1(n20987), .A2(keyinput_g72), .B1(n20959), .B2(
        keyinput_g93), .ZN(n20958) );
  OAI221_X1 U23914 ( .B1(n20987), .B2(keyinput_g72), .C1(n20959), .C2(
        keyinput_g93), .A(n20958), .ZN(n20960) );
  NOR4_X1 U23915 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n20975) );
  AOI22_X1 U23916 ( .A1(n21124), .A2(keyinput_g68), .B1(n20965), .B2(
        keyinput_g52), .ZN(n20964) );
  OAI221_X1 U23917 ( .B1(n21124), .B2(keyinput_g68), .C1(n20965), .C2(
        keyinput_g52), .A(n20964), .ZN(n20973) );
  INV_X1 U23918 ( .A(DATAI_9_), .ZN(n21006) );
  AOI22_X1 U23919 ( .A1(n21006), .A2(keyinput_g23), .B1(keyinput_g46), .B2(
        n21005), .ZN(n20966) );
  OAI221_X1 U23920 ( .B1(n21006), .B2(keyinput_g23), .C1(n21005), .C2(
        keyinput_g46), .A(n20966), .ZN(n20972) );
  AOI22_X1 U23921 ( .A1(n11648), .A2(keyinput_g115), .B1(keyinput_g47), .B2(
        n20968), .ZN(n20967) );
  OAI221_X1 U23922 ( .B1(n11648), .B2(keyinput_g115), .C1(n20968), .C2(
        keyinput_g47), .A(n20967), .ZN(n20971) );
  AOI22_X1 U23923 ( .A1(n21121), .A2(keyinput_g91), .B1(keyinput_g20), .B2(
        n21016), .ZN(n20969) );
  OAI221_X1 U23924 ( .B1(n21121), .B2(keyinput_g91), .C1(n21016), .C2(
        keyinput_g20), .A(n20969), .ZN(n20970) );
  NOR4_X1 U23925 ( .A1(n20973), .A2(n20972), .A3(n20971), .A4(n20970), .ZN(
        n20974) );
  NAND4_X1 U23926 ( .A1(n20977), .A2(n20976), .A3(n20975), .A4(n20974), .ZN(
        n20978) );
  NOR4_X1 U23927 ( .A1(n20981), .A2(n20980), .A3(n20979), .A4(n20978), .ZN(
        n21196) );
  AOI22_X1 U23928 ( .A1(n20984), .A2(keyinput_f29), .B1(n20983), .B2(
        keyinput_f26), .ZN(n20982) );
  OAI221_X1 U23929 ( .B1(n20984), .B2(keyinput_f29), .C1(n20983), .C2(
        keyinput_f26), .A(n20982), .ZN(n20997) );
  INV_X1 U23930 ( .A(READY2), .ZN(n20986) );
  AOI22_X1 U23931 ( .A1(n20987), .A2(keyinput_f72), .B1(keyinput_f37), .B2(
        n20986), .ZN(n20985) );
  OAI221_X1 U23932 ( .B1(n20987), .B2(keyinput_f72), .C1(n20986), .C2(
        keyinput_f37), .A(n20985), .ZN(n20996) );
  AOI22_X1 U23933 ( .A1(n20990), .A2(keyinput_f86), .B1(keyinput_f49), .B2(
        n20989), .ZN(n20988) );
  OAI221_X1 U23934 ( .B1(n20990), .B2(keyinput_f86), .C1(n20989), .C2(
        keyinput_f49), .A(n20988), .ZN(n20995) );
  AOI22_X1 U23935 ( .A1(n20993), .A2(keyinput_f19), .B1(n20992), .B2(
        keyinput_f90), .ZN(n20991) );
  OAI221_X1 U23936 ( .B1(n20993), .B2(keyinput_f19), .C1(n20992), .C2(
        keyinput_f90), .A(n20991), .ZN(n20994) );
  NOR4_X1 U23937 ( .A1(n20997), .A2(n20996), .A3(n20995), .A4(n20994), .ZN(
        n21190) );
  AOI22_X1 U23938 ( .A1(n21000), .A2(keyinput_f106), .B1(keyinput_f10), .B2(
        n20999), .ZN(n20998) );
  OAI221_X1 U23939 ( .B1(n21000), .B2(keyinput_f106), .C1(n20999), .C2(
        keyinput_f10), .A(n20998), .ZN(n21013) );
  AOI22_X1 U23940 ( .A1(n21003), .A2(keyinput_f12), .B1(n21002), .B2(
        keyinput_f121), .ZN(n21001) );
  OAI221_X1 U23941 ( .B1(n21003), .B2(keyinput_f12), .C1(n21002), .C2(
        keyinput_f121), .A(n21001), .ZN(n21012) );
  AOI22_X1 U23942 ( .A1(n21006), .A2(keyinput_f23), .B1(keyinput_f46), .B2(
        n21005), .ZN(n21004) );
  OAI221_X1 U23943 ( .B1(n21006), .B2(keyinput_f23), .C1(n21005), .C2(
        keyinput_f46), .A(n21004), .ZN(n21011) );
  AOI22_X1 U23944 ( .A1(n21009), .A2(keyinput_f100), .B1(keyinput_f76), .B2(
        n21008), .ZN(n21007) );
  OAI221_X1 U23945 ( .B1(n21009), .B2(keyinput_f100), .C1(n21008), .C2(
        keyinput_f76), .A(n21007), .ZN(n21010) );
  NOR4_X1 U23946 ( .A1(n21013), .A2(n21012), .A3(n21011), .A4(n21010), .ZN(
        n21189) );
  AOI22_X1 U23947 ( .A1(n21016), .A2(keyinput_f20), .B1(keyinput_f8), .B2(
        n21015), .ZN(n21014) );
  OAI221_X1 U23948 ( .B1(n21016), .B2(keyinput_f20), .C1(n21015), .C2(
        keyinput_f8), .A(n21014), .ZN(n21044) );
  AOI22_X1 U23949 ( .A1(n14523), .A2(keyinput_f55), .B1(n14474), .B2(
        keyinput_f125), .ZN(n21017) );
  OAI221_X1 U23950 ( .B1(n14523), .B2(keyinput_f55), .C1(n14474), .C2(
        keyinput_f125), .A(n21017), .ZN(n21043) );
  XOR2_X1 U23951 ( .A(keyinput_f42), .B(P1_D_C_N_REG_SCAN_IN), .Z(n21022) );
  AOI22_X1 U23952 ( .A1(n21020), .A2(keyinput_f92), .B1(keyinput_f107), .B2(
        n21019), .ZN(n21018) );
  OAI221_X1 U23953 ( .B1(n21020), .B2(keyinput_f92), .C1(n21019), .C2(
        keyinput_f107), .A(n21018), .ZN(n21021) );
  AOI211_X1 U23954 ( .C1(n21024), .C2(keyinput_f11), .A(n21022), .B(n21021), 
        .ZN(n21023) );
  OAI21_X1 U23955 ( .B1(n21024), .B2(keyinput_f11), .A(n21023), .ZN(n21042) );
  AOI22_X1 U23956 ( .A1(n21027), .A2(keyinput_f56), .B1(keyinput_f63), .B2(
        n21026), .ZN(n21025) );
  OAI221_X1 U23957 ( .B1(n21027), .B2(keyinput_f56), .C1(n21026), .C2(
        keyinput_f63), .A(n21025), .ZN(n21040) );
  AOI22_X1 U23958 ( .A1(n21030), .A2(keyinput_f113), .B1(keyinput_f74), .B2(
        n21029), .ZN(n21028) );
  OAI221_X1 U23959 ( .B1(n21030), .B2(keyinput_f113), .C1(n21029), .C2(
        keyinput_f74), .A(n21028), .ZN(n21039) );
  AOI22_X1 U23960 ( .A1(n21033), .A2(keyinput_f14), .B1(n21032), .B2(
        keyinput_f73), .ZN(n21031) );
  OAI221_X1 U23961 ( .B1(n21033), .B2(keyinput_f14), .C1(n21032), .C2(
        keyinput_f73), .A(n21031), .ZN(n21038) );
  INV_X1 U23962 ( .A(keyinput_f35), .ZN(n21035) );
  AOI22_X1 U23963 ( .A1(n21036), .A2(keyinput_f124), .B1(BS16), .B2(n21035), 
        .ZN(n21034) );
  OAI221_X1 U23964 ( .B1(n21036), .B2(keyinput_f124), .C1(n21035), .C2(BS16), 
        .A(n21034), .ZN(n21037) );
  OR4_X1 U23965 ( .A1(n21040), .A2(n21039), .A3(n21038), .A4(n21037), .ZN(
        n21041) );
  NOR4_X1 U23966 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21188) );
  OAI22_X1 U23967 ( .A1(P1_EAX_REG_25__SCAN_IN), .A2(keyinput_f122), .B1(
        keyinput_f93), .B2(P1_EBX_REG_22__SCAN_IN), .ZN(n21045) );
  AOI221_X1 U23968 ( .B1(P1_EAX_REG_25__SCAN_IN), .B2(keyinput_f122), .C1(
        P1_EBX_REG_22__SCAN_IN), .C2(keyinput_f93), .A(n21045), .ZN(n21052) );
  OAI22_X1 U23969 ( .A1(P1_EBX_REG_12__SCAN_IN), .A2(keyinput_f103), .B1(
        keyinput_f31), .B2(DATAI_1_), .ZN(n21046) );
  AOI221_X1 U23970 ( .B1(P1_EBX_REG_12__SCAN_IN), .B2(keyinput_f103), .C1(
        DATAI_1_), .C2(keyinput_f31), .A(n21046), .ZN(n21051) );
  OAI22_X1 U23971 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(keyinput_f127), .B1(
        keyinput_f60), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n21047) );
  AOI221_X1 U23972 ( .B1(P1_EAX_REG_20__SCAN_IN), .B2(keyinput_f127), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_f60), .A(n21047), .ZN(n21050)
         );
  OAI22_X1 U23973 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_f45), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_f41), .ZN(n21048) );
  AOI221_X1 U23974 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_f45), .C1(
        keyinput_f41), .C2(P1_M_IO_N_REG_SCAN_IN), .A(n21048), .ZN(n21049) );
  NAND4_X1 U23975 ( .A1(n21052), .A2(n21051), .A3(n21050), .A4(n21049), .ZN(
        n21186) );
  OAI22_X1 U23976 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(keyinput_f53), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(keyinput_f75), .ZN(n21053) );
  AOI221_X1 U23977 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(keyinput_f53), .C1(
        keyinput_f75), .C2(P1_REIP_REG_8__SCAN_IN), .A(n21053), .ZN(n21079) );
  OAI22_X1 U23978 ( .A1(P1_EBX_REG_27__SCAN_IN), .A2(keyinput_f88), .B1(
        keyinput_f47), .B2(P1_W_R_N_REG_SCAN_IN), .ZN(n21054) );
  AOI221_X1 U23979 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(keyinput_f88), .C1(
        P1_W_R_N_REG_SCAN_IN), .C2(keyinput_f47), .A(n21054), .ZN(n21057) );
  OAI22_X1 U23980 ( .A1(DATAI_7_), .A2(keyinput_f25), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .ZN(n21055) );
  AOI221_X1 U23981 ( .B1(DATAI_7_), .B2(keyinput_f25), .C1(keyinput_f38), .C2(
        P1_READREQUEST_REG_SCAN_IN), .A(n21055), .ZN(n21056) );
  OAI211_X1 U23982 ( .C1(n21059), .C2(keyinput_f97), .A(n21057), .B(n21056), 
        .ZN(n21058) );
  AOI21_X1 U23983 ( .B1(n21059), .B2(keyinput_f97), .A(n21058), .ZN(n21078) );
  AOI22_X1 U23984 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(keyinput_f66), .B1(
        P1_EBX_REG_6__SCAN_IN), .B2(keyinput_f109), .ZN(n21060) );
  OAI221_X1 U23985 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(keyinput_f66), .C1(
        P1_EBX_REG_6__SCAN_IN), .C2(keyinput_f109), .A(n21060), .ZN(n21067) );
  AOI22_X1 U23986 ( .A1(DATAI_25_), .A2(keyinput_f7), .B1(
        P1_REIP_REG_5__SCAN_IN), .B2(keyinput_f78), .ZN(n21061) );
  OAI221_X1 U23987 ( .B1(DATAI_25_), .B2(keyinput_f7), .C1(
        P1_REIP_REG_5__SCAN_IN), .C2(keyinput_f78), .A(n21061), .ZN(n21066) );
  AOI22_X1 U23988 ( .A1(READY1), .A2(keyinput_f36), .B1(P1_EAX_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n21062) );
  OAI221_X1 U23989 ( .B1(READY1), .B2(keyinput_f36), .C1(
        P1_EAX_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n21062), .ZN(n21065)
         );
  AOI22_X1 U23990 ( .A1(P1_EBX_REG_11__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_EBX_REG_13__SCAN_IN), .B2(keyinput_f102), .ZN(n21063) );
  OAI221_X1 U23991 ( .B1(P1_EBX_REG_11__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_EBX_REG_13__SCAN_IN), .C2(keyinput_f102), .A(n21063), .ZN(n21064)
         );
  NOR4_X1 U23992 ( .A1(n21067), .A2(n21066), .A3(n21065), .A4(n21064), .ZN(
        n21077) );
  AOI22_X1 U23993 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(keyinput_f83), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(keyinput_f64), .ZN(n21068) );
  OAI221_X1 U23994 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(keyinput_f83), .C1(
        P1_REIP_REG_19__SCAN_IN), .C2(keyinput_f64), .A(n21068), .ZN(n21075)
         );
  AOI22_X1 U23995 ( .A1(DATAI_14_), .A2(keyinput_f18), .B1(
        P1_EBX_REG_1__SCAN_IN), .B2(keyinput_f114), .ZN(n21069) );
  OAI221_X1 U23996 ( .B1(DATAI_14_), .B2(keyinput_f18), .C1(
        P1_EBX_REG_1__SCAN_IN), .C2(keyinput_f114), .A(n21069), .ZN(n21074) );
  AOI22_X1 U23997 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_f0), .B1(
        DATAI_15_), .B2(keyinput_f17), .ZN(n21070) );
  OAI221_X1 U23998 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_f0), .C1(
        DATAI_15_), .C2(keyinput_f17), .A(n21070), .ZN(n21073) );
  AOI22_X1 U23999 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(keyinput_f69), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(keyinput_f84), .ZN(n21071) );
  OAI221_X1 U24000 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(keyinput_f69), .C1(
        P1_EBX_REG_31__SCAN_IN), .C2(keyinput_f84), .A(n21071), .ZN(n21072) );
  NOR4_X1 U24001 ( .A1(n21075), .A2(n21074), .A3(n21073), .A4(n21072), .ZN(
        n21076) );
  NAND4_X1 U24002 ( .A1(n21079), .A2(n21078), .A3(n21077), .A4(n21076), .ZN(
        n21185) );
  AOI22_X1 U24003 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(keyinput_f80), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(keyinput_f108), .ZN(n21080) );
  OAI221_X1 U24004 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(keyinput_f80), .C1(
        P1_EBX_REG_7__SCAN_IN), .C2(keyinput_f108), .A(n21080), .ZN(n21087) );
  AOI22_X1 U24005 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(keyinput_f67), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .ZN(n21081) );
  OAI221_X1 U24006 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(keyinput_f67), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_f62), .A(n21081), .ZN(n21086)
         );
  AOI22_X1 U24007 ( .A1(DATAI_31_), .A2(keyinput_f1), .B1(
        P1_EBX_REG_28__SCAN_IN), .B2(keyinput_f87), .ZN(n21082) );
  OAI221_X1 U24008 ( .B1(DATAI_31_), .B2(keyinput_f1), .C1(
        P1_EBX_REG_28__SCAN_IN), .C2(keyinput_f87), .A(n21082), .ZN(n21085) );
  AOI22_X1 U24009 ( .A1(P1_EBX_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(keyinput_f120), .ZN(n21083) );
  OAI221_X1 U24010 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        P1_EAX_REG_27__SCAN_IN), .C2(keyinput_f120), .A(n21083), .ZN(n21084)
         );
  NOR4_X1 U24011 ( .A1(n21087), .A2(n21086), .A3(n21085), .A4(n21084), .ZN(
        n21116) );
  AOI22_X1 U24012 ( .A1(P1_EAX_REG_31__SCAN_IN), .A2(keyinput_f116), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(keyinput_f119), .ZN(n21088) );
  OAI221_X1 U24013 ( .B1(P1_EAX_REG_31__SCAN_IN), .B2(keyinput_f116), .C1(
        P1_EAX_REG_28__SCAN_IN), .C2(keyinput_f119), .A(n21088), .ZN(n21095)
         );
  AOI22_X1 U24014 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(keyinput_f54), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(keyinput_f118), .ZN(n21089) );
  OAI221_X1 U24015 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_f54), .C1(
        P1_EAX_REG_29__SCAN_IN), .C2(keyinput_f118), .A(n21089), .ZN(n21094)
         );
  AOI22_X1 U24016 ( .A1(P1_EBX_REG_20__SCAN_IN), .A2(keyinput_f95), .B1(
        P1_EBX_REG_21__SCAN_IN), .B2(keyinput_f94), .ZN(n21090) );
  OAI221_X1 U24017 ( .B1(P1_EBX_REG_20__SCAN_IN), .B2(keyinput_f95), .C1(
        P1_EBX_REG_21__SCAN_IN), .C2(keyinput_f94), .A(n21090), .ZN(n21093) );
  AOI22_X1 U24018 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(keyinput_f65), .B1(
        P1_REIP_REG_31__SCAN_IN), .B2(keyinput_f52), .ZN(n21091) );
  OAI221_X1 U24019 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(keyinput_f65), .C1(
        P1_REIP_REG_31__SCAN_IN), .C2(keyinput_f52), .A(n21091), .ZN(n21092)
         );
  NOR4_X1 U24020 ( .A1(n21095), .A2(n21094), .A3(n21093), .A4(n21092), .ZN(
        n21115) );
  AOI22_X1 U24021 ( .A1(DATAI_5_), .A2(keyinput_f27), .B1(
        P1_REIP_REG_1__SCAN_IN), .B2(keyinput_f82), .ZN(n21096) );
  OAI221_X1 U24022 ( .B1(DATAI_5_), .B2(keyinput_f27), .C1(
        P1_REIP_REG_1__SCAN_IN), .C2(keyinput_f82), .A(n21096), .ZN(n21103) );
  AOI22_X1 U24023 ( .A1(keyinput_f51), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        DATAI_19_), .B2(keyinput_f13), .ZN(n21097) );
  OAI221_X1 U24024 ( .B1(keyinput_f51), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), 
        .C1(DATAI_19_), .C2(keyinput_f13), .A(n21097), .ZN(n21102) );
  AOI22_X1 U24025 ( .A1(DATAI_8_), .A2(keyinput_f24), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(keyinput_f126), .ZN(n21098) );
  OAI221_X1 U24026 ( .B1(DATAI_8_), .B2(keyinput_f24), .C1(
        P1_EAX_REG_21__SCAN_IN), .C2(keyinput_f126), .A(n21098), .ZN(n21101)
         );
  AOI22_X1 U24027 ( .A1(keyinput_f39), .A2(P1_ADS_N_REG_SCAN_IN), .B1(
        P1_EBX_REG_0__SCAN_IN), .B2(keyinput_f115), .ZN(n21099) );
  OAI221_X1 U24028 ( .B1(keyinput_f39), .B2(P1_ADS_N_REG_SCAN_IN), .C1(
        P1_EBX_REG_0__SCAN_IN), .C2(keyinput_f115), .A(n21099), .ZN(n21100) );
  NOR4_X1 U24029 ( .A1(n21103), .A2(n21102), .A3(n21101), .A4(n21100), .ZN(
        n21114) );
  AOI22_X1 U24030 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(keyinput_f123), .ZN(n21104) );
  OAI221_X1 U24031 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(
        P1_EAX_REG_24__SCAN_IN), .C2(keyinput_f123), .A(n21104), .ZN(n21112)
         );
  AOI22_X1 U24032 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput_f43), 
        .B1(DATAI_11_), .B2(keyinput_f21), .ZN(n21105) );
  OAI221_X1 U24033 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_f43), 
        .C1(DATAI_11_), .C2(keyinput_f21), .A(n21105), .ZN(n21111) );
  AOI22_X1 U24034 ( .A1(DATAI_4_), .A2(keyinput_f28), .B1(DATAI_30_), .B2(
        keyinput_f2), .ZN(n21106) );
  OAI221_X1 U24035 ( .B1(DATAI_4_), .B2(keyinput_f28), .C1(DATAI_30_), .C2(
        keyinput_f2), .A(n21106), .ZN(n21110) );
  AOI22_X1 U24036 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput_f40), .B1(
        n21108), .B2(keyinput_f32), .ZN(n21107) );
  OAI221_X1 U24037 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_f40), .C1(
        n21108), .C2(keyinput_f32), .A(n21107), .ZN(n21109) );
  NOR4_X1 U24038 ( .A1(n21112), .A2(n21111), .A3(n21110), .A4(n21109), .ZN(
        n21113) );
  NAND4_X1 U24039 ( .A1(n21116), .A2(n21115), .A3(n21114), .A4(n21113), .ZN(
        n21184) );
  AOI22_X1 U24040 ( .A1(n21119), .A2(keyinput_f30), .B1(keyinput_f15), .B2(
        n21118), .ZN(n21117) );
  OAI221_X1 U24041 ( .B1(n21119), .B2(keyinput_f30), .C1(n21118), .C2(
        keyinput_f15), .A(n21117), .ZN(n21132) );
  AOI22_X1 U24042 ( .A1(n21122), .A2(keyinput_f9), .B1(n21121), .B2(
        keyinput_f91), .ZN(n21120) );
  OAI221_X1 U24043 ( .B1(n21122), .B2(keyinput_f9), .C1(n21121), .C2(
        keyinput_f91), .A(n21120), .ZN(n21131) );
  AOI22_X1 U24044 ( .A1(n21125), .A2(keyinput_f96), .B1(keyinput_f68), .B2(
        n21124), .ZN(n21123) );
  OAI221_X1 U24045 ( .B1(n21125), .B2(keyinput_f96), .C1(n21124), .C2(
        keyinput_f68), .A(n21123), .ZN(n21130) );
  AOI22_X1 U24046 ( .A1(n21128), .A2(keyinput_f85), .B1(n21127), .B2(
        keyinput_f44), .ZN(n21126) );
  OAI221_X1 U24047 ( .B1(n21128), .B2(keyinput_f85), .C1(n21127), .C2(
        keyinput_f44), .A(n21126), .ZN(n21129) );
  NOR4_X1 U24048 ( .A1(n21132), .A2(n21131), .A3(n21130), .A4(n21129), .ZN(
        n21182) );
  AOI22_X1 U24049 ( .A1(n21135), .A2(keyinput_f16), .B1(n21134), .B2(
        keyinput_f99), .ZN(n21133) );
  OAI221_X1 U24050 ( .B1(n21135), .B2(keyinput_f16), .C1(n21134), .C2(
        keyinput_f99), .A(n21133), .ZN(n21148) );
  AOI22_X1 U24051 ( .A1(n21138), .A2(keyinput_f70), .B1(keyinput_f5), .B2(
        n21137), .ZN(n21136) );
  OAI221_X1 U24052 ( .B1(n21138), .B2(keyinput_f70), .C1(n21137), .C2(
        keyinput_f5), .A(n21136), .ZN(n21147) );
  AOI22_X1 U24053 ( .A1(n21141), .A2(keyinput_f77), .B1(n21140), .B2(
        keyinput_f58), .ZN(n21139) );
  OAI221_X1 U24054 ( .B1(n21141), .B2(keyinput_f77), .C1(n21140), .C2(
        keyinput_f58), .A(n21139), .ZN(n21146) );
  INV_X1 U24055 ( .A(keyinput_f50), .ZN(n21143) );
  AOI22_X1 U24056 ( .A1(n21144), .A2(keyinput_f61), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n21143), .ZN(n21142) );
  OAI221_X1 U24057 ( .B1(n21144), .B2(keyinput_f61), .C1(n21143), .C2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A(n21142), .ZN(n21145) );
  NOR4_X1 U24058 ( .A1(n21148), .A2(n21147), .A3(n21146), .A4(n21145), .ZN(
        n21181) );
  AOI22_X1 U24059 ( .A1(n21151), .A2(keyinput_f81), .B1(n21150), .B2(
        keyinput_f111), .ZN(n21149) );
  OAI221_X1 U24060 ( .B1(n21151), .B2(keyinput_f81), .C1(n21150), .C2(
        keyinput_f111), .A(n21149), .ZN(n21164) );
  AOI22_X1 U24061 ( .A1(n21154), .A2(keyinput_f71), .B1(keyinput_f48), .B2(
        n21153), .ZN(n21152) );
  OAI221_X1 U24062 ( .B1(n21154), .B2(keyinput_f71), .C1(n21153), .C2(
        keyinput_f48), .A(n21152), .ZN(n21163) );
  AOI22_X1 U24063 ( .A1(n21157), .A2(keyinput_f110), .B1(n21156), .B2(
        keyinput_f98), .ZN(n21155) );
  OAI221_X1 U24064 ( .B1(n21157), .B2(keyinput_f110), .C1(n21156), .C2(
        keyinput_f98), .A(n21155), .ZN(n21162) );
  INV_X1 U24065 ( .A(keyinput_f33), .ZN(n21159) );
  AOI22_X1 U24066 ( .A1(n21160), .A2(keyinput_f3), .B1(HOLD), .B2(n21159), 
        .ZN(n21158) );
  OAI221_X1 U24067 ( .B1(n21160), .B2(keyinput_f3), .C1(n21159), .C2(HOLD), 
        .A(n21158), .ZN(n21161) );
  NOR4_X1 U24068 ( .A1(n21164), .A2(n21163), .A3(n21162), .A4(n21161), .ZN(
        n21180) );
  AOI22_X1 U24069 ( .A1(n21167), .A2(keyinput_f89), .B1(keyinput_f4), .B2(
        n21166), .ZN(n21165) );
  OAI221_X1 U24070 ( .B1(n21167), .B2(keyinput_f89), .C1(n21166), .C2(
        keyinput_f4), .A(n21165), .ZN(n21178) );
  AOI22_X1 U24071 ( .A1(n21170), .A2(keyinput_f79), .B1(n21169), .B2(
        keyinput_f59), .ZN(n21168) );
  OAI221_X1 U24072 ( .B1(n21170), .B2(keyinput_f79), .C1(n21169), .C2(
        keyinput_f59), .A(n21168), .ZN(n21177) );
  AOI22_X1 U24073 ( .A1(n21172), .A2(keyinput_f112), .B1(keyinput_f57), .B2(
        n14344), .ZN(n21171) );
  OAI221_X1 U24074 ( .B1(n21172), .B2(keyinput_f112), .C1(n14344), .C2(
        keyinput_f57), .A(n21171), .ZN(n21176) );
  AOI22_X1 U24075 ( .A1(n13755), .A2(keyinput_f105), .B1(keyinput_f34), .B2(
        n21174), .ZN(n21173) );
  OAI221_X1 U24076 ( .B1(n13755), .B2(keyinput_f105), .C1(n21174), .C2(
        keyinput_f34), .A(n21173), .ZN(n21175) );
  NOR4_X1 U24077 ( .A1(n21178), .A2(n21177), .A3(n21176), .A4(n21175), .ZN(
        n21179) );
  NAND4_X1 U24078 ( .A1(n21182), .A2(n21181), .A3(n21180), .A4(n21179), .ZN(
        n21183) );
  NOR4_X1 U24079 ( .A1(n21186), .A2(n21185), .A3(n21184), .A4(n21183), .ZN(
        n21187) );
  NAND4_X1 U24080 ( .A1(n21190), .A2(n21189), .A3(n21188), .A4(n21187), .ZN(
        n21192) );
  AOI21_X1 U24081 ( .B1(keyinput_f22), .B2(n21192), .A(DATAI_10_), .ZN(n21194)
         );
  INV_X1 U24082 ( .A(keyinput_f22), .ZN(n21191) );
  AOI21_X1 U24083 ( .B1(n21192), .B2(n21191), .A(keyinput_g22), .ZN(n21193) );
  AOI22_X1 U24084 ( .A1(keyinput_g22), .A2(n21194), .B1(DATAI_10_), .B2(n21193), .ZN(n21195) );
  AOI21_X1 U24085 ( .B1(n21197), .B2(n21196), .A(n21195), .ZN(n21199) );
  AOI22_X1 U24086 ( .A1(n16464), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16466), .ZN(n21198) );
  XNOR2_X1 U24087 ( .A(n21199), .B(n21198), .ZN(U355) );
  OR2_X1 U12760 ( .A1(n10338), .A2(n10337), .ZN(n11518) );
  BUF_X1 U11334 ( .A(n13047), .Z(n9819) );
  INV_X4 U11330 ( .A(n21200), .ZN(n9814) );
  CLKBUF_X1 U11293 ( .A(n10680), .Z(n11077) );
  CLKBUF_X1 U11303 ( .A(n10519), .Z(n10561) );
  CLKBUF_X1 U11321 ( .A(n11299), .Z(n17641) );
  CLKBUF_X1 U11333 ( .A(n11659), .Z(n11737) );
  CLKBUF_X1 U12228 ( .A(n12110), .Z(n12125) );
  INV_X2 U12361 ( .A(n10206), .ZN(n12264) );
  CLKBUF_X1 U12429 ( .A(n13029), .Z(n19251) );
  AOI22_X1 U12490 ( .A1(n11325), .A2(n11324), .B1(n11323), .B2(n11322), .ZN(
        n12834) );
  CLKBUF_X1 U12757 ( .A(n16460), .Z(n16454) );
  NAND2_X1 U12761 ( .A1(n14257), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n21200) );
endmodule

