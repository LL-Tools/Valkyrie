

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019;

  NAND2_X1 U3556 ( .A1(n5468), .A2(n5469), .ZN(n5461) );
  AND2_X1 U3557 ( .A1(n6693), .A2(n4392), .ZN(n6095) );
  BUF_X2 U3558 ( .A(n3603), .Z(n5318) );
  CLKBUF_X1 U3559 ( .A(n3688), .Z(n5043) );
  CLKBUF_X2 U3560 ( .A(n3371), .Z(n4145) );
  CLKBUF_X2 U3561 ( .A(n4154), .Z(n4115) );
  CLKBUF_X2 U3562 ( .A(n3299), .Z(n4099) );
  CLKBUF_X2 U3563 ( .A(n3297), .Z(n4152) );
  CLKBUF_X2 U3564 ( .A(n3402), .Z(n4094) );
  CLKBUF_X2 U3565 ( .A(n3298), .Z(n4117) );
  CLKBUF_X2 U3566 ( .A(n3306), .Z(n4143) );
  CLKBUF_X2 U3567 ( .A(n3380), .Z(n4114) );
  CLKBUF_X2 U3568 ( .A(n3270), .Z(n4146) );
  CLKBUF_X2 U3569 ( .A(n3307), .Z(n4142) );
  CLKBUF_X2 U3570 ( .A(n3277), .Z(n4144) );
  AND4_X1 U3571 ( .A1(n3282), .A2(n3281), .A3(n3280), .A4(n3279), .ZN(n3283)
         );
  AND4_X1 U3572 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3268)
         );
  BUF_X2 U3573 ( .A(n3278), .Z(n4154) );
  AND2_X2 U3574 ( .A1(n3192), .A2(n4523), .ZN(n3380) );
  AND2_X1 U3575 ( .A1(n3184), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3189)
         );
  AND2_X1 U3576 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4598) );
  CLKBUF_X2 U3577 ( .A(n3271), .Z(n4116) );
  NOR2_X1 U3578 ( .A1(n3643), .A2(n3317), .ZN(n3665) );
  AND3_X1 U3580 ( .A1(n3319), .A2(n3318), .A3(n3351), .ZN(n3325) );
  NOR2_X1 U3582 ( .A1(n4697), .A2(n6334), .ZN(n3691) );
  CLKBUF_X2 U3583 ( .A(n3272), .Z(n3365) );
  NAND2_X1 U3584 ( .A1(n5412), .A2(n4397), .ZN(n6092) );
  AOI211_X1 U3585 ( .C1(n3117), .C2(n5401), .A(n5402), .B(n5403), .ZN(n4426)
         );
  AND2_X2 U3586 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4523) );
  OAI22_X1 U3587 ( .A1(n5811), .A2(n6044), .B1(n5810), .B2(n6104), .ZN(n5812)
         );
  OAI22_X1 U3588 ( .A1(n5401), .A2(n5698), .B1(n5426), .B2(n5400), .ZN(n5430)
         );
  AND2_X1 U3589 ( .A1(n4547), .A2(n6583), .ZN(n4477) );
  INV_X1 U3590 ( .A(n6096), .ZN(n6108) );
  OAI21_X1 U3591 ( .B1(n3676), .B2(n3433), .A(n3510), .ZN(n3511) );
  AOI21_X1 U3592 ( .B1(n4590), .B2(n6576), .A(n3458), .ZN(n3461) );
  INV_X1 U3593 ( .A(n3355), .ZN(n5092) );
  NAND4_X4 U3594 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3320)
         );
  AND4_X2 U3595 ( .A1(n3213), .A2(n3212), .A3(n3211), .A4(n3210), .ZN(n3229)
         );
  NAND2_X2 U3596 ( .A1(n5529), .A2(n3613), .ZN(n5694) );
  NOR2_X4 U3597 ( .A1(n6095), .A2(n6334), .ZN(n5412) );
  XNOR2_X1 U3598 ( .A(n5423), .B(n4385), .ZN(n5391) );
  CLKBUF_X1 U3599 ( .A(n5555), .Z(n5720) );
  NAND2_X1 U3600 ( .A1(n4975), .A2(n3589), .ZN(n5177) );
  NAND2_X1 U3601 ( .A1(n4977), .A2(n4976), .ZN(n4975) );
  NAND2_X2 U3602 ( .A1(n3141), .A2(n4733), .ZN(n4732) );
  INV_X4 U3603 ( .A(n3602), .ZN(n5554) );
  XNOR2_X1 U3604 ( .A(n3463), .B(n3462), .ZN(n3419) );
  INV_X1 U3605 ( .A(n3342), .ZN(n3421) );
  CLKBUF_X1 U3606 ( .A(n3351), .Z(n4697) );
  NAND2_X2 U3607 ( .A1(n3313), .A2(n3345), .ZN(n4230) );
  AND4_X1 U3608 ( .A1(n3276), .A2(n3275), .A3(n3274), .A4(n3273), .ZN(n3284)
         );
  AND4_X1 U3609 ( .A1(n3263), .A2(n3262), .A3(n3261), .A4(n3260), .ZN(n3269)
         );
  BUF_X2 U3610 ( .A(n3295), .Z(n4153) );
  AOI22_X1 U3611 ( .A1(n3299), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3262) );
  BUF_X2 U3612 ( .A(n3370), .Z(n4147) );
  INV_X2 U3613 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3183) );
  NOR2_X4 U3614 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3191) );
  AOI21_X1 U3615 ( .B1(n5497), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n4383), 
        .ZN(n4384) );
  OR2_X2 U3616 ( .A1(n5424), .A2(n5423), .ZN(n5811) );
  NOR2_X1 U3617 ( .A1(n3165), .A2(n3164), .ZN(n3163) );
  INV_X1 U3618 ( .A(n3165), .ZN(n5423) );
  AOI211_X1 U3619 ( .C1(n6196), .C2(n5834), .A(n5524), .B(n5523), .ZN(n5525)
         );
  CLKBUF_X1 U3620 ( .A(n5440), .Z(n5441) );
  NOR2_X2 U3621 ( .A1(n5461), .A2(n3170), .ZN(n4373) );
  OAI21_X1 U3622 ( .B1(n5340), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5554), 
        .ZN(n3605) );
  OR2_X1 U3623 ( .A1(n5430), .A2(n5429), .ZN(n5810) );
  INV_X1 U3624 ( .A(n5401), .ZN(n4423) );
  INV_X1 U3625 ( .A(n5325), .ZN(n3858) );
  AND2_X2 U3626 ( .A1(n5639), .A2(n5436), .ZN(n3117) );
  XNOR2_X1 U3627 ( .A(n3593), .B(n3581), .ZN(n3732) );
  AND4_X1 U3628 ( .A1(n4623), .A2(n3706), .A3(n4624), .A4(n3172), .ZN(n4629)
         );
  AND2_X1 U3629 ( .A1(n3479), .A2(n3478), .ZN(n4655) );
  NAND2_X1 U3630 ( .A1(n3705), .A2(n4692), .ZN(n4623) );
  XNOR2_X1 U3631 ( .A(n3555), .B(n3556), .ZN(n3718) );
  NAND2_X1 U3632 ( .A1(n3534), .A2(n3533), .ZN(n3555) );
  OR2_X1 U3633 ( .A1(n4461), .A2(n4694), .ZN(n4624) );
  NAND2_X1 U3634 ( .A1(n3683), .A2(n3870), .ZN(n4694) );
  AND2_X1 U3635 ( .A1(n4463), .A2(n4462), .ZN(n4461) );
  CLKBUF_X1 U3636 ( .A(n4643), .Z(n4990) );
  CLKBUF_X1 U3637 ( .A(n4637), .Z(n4993) );
  CLKBUF_X1 U3638 ( .A(n4566), .Z(n6677) );
  AOI21_X2 U3639 ( .B1(n4566), .B2(n6576), .A(n3502), .ZN(n4989) );
  XNOR2_X1 U3640 ( .A(n3419), .B(n3418), .ZN(n4637) );
  XNOR2_X1 U3641 ( .A(n4603), .B(n5131), .ZN(n4566) );
  NAND2_X1 U3642 ( .A1(n3430), .A2(n3119), .ZN(n3465) );
  CLKBUF_X1 U3643 ( .A(n3689), .Z(n3690) );
  NAND2_X1 U3644 ( .A1(n3489), .A2(n3488), .ZN(n5131) );
  CLKBUF_X1 U3645 ( .A(n4212), .Z(n4605) );
  AND2_X1 U3646 ( .A1(n3348), .A2(n3347), .ZN(n4333) );
  INV_X1 U3647 ( .A(n3462), .ZN(n3464) );
  NOR2_X1 U3648 ( .A1(n4232), .A2(n4231), .ZN(n4620) );
  CLKBUF_X1 U3649 ( .A(n4213), .Z(n4537) );
  CLKBUF_X1 U3650 ( .A(n4207), .Z(n4540) );
  AND2_X1 U3651 ( .A1(n3394), .A2(n3393), .ZN(n3462) );
  AND2_X1 U3652 ( .A1(n3350), .A2(n4325), .ZN(n3160) );
  AND2_X1 U3653 ( .A1(n3287), .A2(n4336), .ZN(n3339) );
  OAI21_X1 U3654 ( .B1(n3342), .B2(n3323), .A(n3322), .ZN(n3324) );
  AND3_X1 U3655 ( .A1(n3350), .A2(n3349), .A3(n4325), .ZN(n4207) );
  AND2_X1 U3656 ( .A1(n3421), .A2(n3313), .ZN(n4325) );
  AND2_X1 U3657 ( .A1(n3292), .A2(n3351), .ZN(n3293) );
  CLKBUF_X1 U3658 ( .A(n3315), .Z(n4690) );
  CLKBUF_X1 U3659 ( .A(n3343), .Z(n4445) );
  AND2_X1 U3660 ( .A1(n4335), .A2(n4220), .ZN(n6541) );
  NOR2_X1 U3661 ( .A1(n3342), .A2(n3313), .ZN(n4457) );
  INV_X1 U3662 ( .A(n3469), .ZN(n3420) );
  AND2_X1 U3663 ( .A1(n3317), .A2(n3337), .ZN(n3349) );
  OR2_X1 U3664 ( .A1(n3390), .A2(n3389), .ZN(n3594) );
  NAND2_X1 U3665 ( .A1(n3312), .A2(n3118), .ZN(n3342) );
  NOR2_X2 U3666 ( .A1(n4456), .A2(n6334), .ZN(n3677) );
  NOR2_X1 U3667 ( .A1(n3304), .A2(n3303), .ZN(n3312) );
  AND2_X2 U3668 ( .A1(n3198), .A2(n3197), .ZN(n3317) );
  AND4_X1 U3669 ( .A1(n3251), .A2(n3250), .A3(n3249), .A4(n3248), .ZN(n3257)
         );
  AND4_X1 U3670 ( .A1(n3188), .A2(n3187), .A3(n3186), .A4(n3185), .ZN(n3198)
         );
  NAND2_X1 U3671 ( .A1(n3239), .A2(n3238), .ZN(n3321) );
  NAND2_X2 U3672 ( .A1(n3284), .A2(n3283), .ZN(n3313) );
  AND4_X1 U3673 ( .A1(n3243), .A2(n3242), .A3(n3241), .A4(n3240), .ZN(n3259)
         );
  AND4_X1 U3674 ( .A1(n3247), .A2(n3246), .A3(n3245), .A4(n3244), .ZN(n3258)
         );
  AND4_X1 U3675 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3227)
         );
  AND4_X1 U3676 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3238)
         );
  AND4_X1 U3677 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3226)
         );
  AND4_X1 U3678 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3209)
         );
  AND4_X1 U3679 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3239)
         );
  AND4_X1 U3680 ( .A1(n3196), .A2(n3195), .A3(n3194), .A4(n3193), .ZN(n3197)
         );
  AND4_X1 U3681 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3256)
         );
  AND4_X1 U3682 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3228)
         );
  NOR2_X1 U3683 ( .A1(n6656), .A2(STATE_REG_2__SCAN_IN), .ZN(n6651) );
  BUF_X2 U3684 ( .A(n3305), .Z(n4073) );
  INV_X1 U3686 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6662) );
  AND2_X1 U3687 ( .A1(n3728), .A2(n4682), .ZN(n3109) );
  NOR2_X1 U3688 ( .A1(n5561), .A2(n3167), .ZN(n3110) );
  AND2_X1 U3689 ( .A1(n3111), .A2(n3779), .ZN(n5171) );
  NOR2_X1 U3690 ( .A1(n5173), .A2(n5085), .ZN(n3111) );
  OR2_X1 U3691 ( .A1(n5442), .A2(n5515), .ZN(n3112) );
  NOR2_X1 U3692 ( .A1(n5561), .A2(n3167), .ZN(n5477) );
  NAND2_X1 U3693 ( .A1(n5366), .A2(n5949), .ZN(n5561) );
  NOR2_X1 U3694 ( .A1(n4728), .A2(n4729), .ZN(n4771) );
  NAND2_X1 U3695 ( .A1(n4732), .A2(n3554), .ZN(n3113) );
  CLKBUF_X1 U3696 ( .A(n4811), .Z(n3114) );
  AND2_X2 U3697 ( .A1(n3180), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4531)
         );
  OR2_X4 U3698 ( .A1(n3346), .A2(n3313), .ZN(n4224) );
  NAND2_X2 U3699 ( .A1(n5177), .A2(n5176), .ZN(n5175) );
  NAND2_X1 U3700 ( .A1(n3332), .A2(n3331), .ZN(n3397) );
  NAND2_X2 U3701 ( .A1(n3156), .A2(n3437), .ZN(n6219) );
  NAND2_X2 U3702 ( .A1(n3532), .A2(n3505), .ZN(n3676) );
  NOR2_X2 U3703 ( .A1(n5540), .A2(n4184), .ZN(n5535) );
  NOR2_X2 U3704 ( .A1(n5542), .A2(n5541), .ZN(n5540) );
  INV_X1 U3705 ( .A(n3346), .ZN(n3115) );
  AND2_X2 U3707 ( .A1(n5171), .A2(n5234), .ZN(n5235) );
  AOI22_X2 U3710 ( .A1(n5547), .A2(n5548), .B1(n5582), .B2(n6759), .ZN(n5542)
         );
  AOI22_X2 U3711 ( .A1(n5694), .A2(n5696), .B1(n5554), .B2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5547) );
  NOR3_X4 U3712 ( .A1(n5453), .A2(n5444), .A3(n5640), .ZN(n5639) );
  AOI211_X1 U3713 ( .C1(n5618), .C2(n6107), .A(n4440), .B(n4439), .ZN(n4441)
         );
  NOR2_X2 U3714 ( .A1(n5442), .A2(n5515), .ZN(n5432) );
  AND4_X1 U3715 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3116)
         );
  AND4_X4 U3716 ( .A1(n3259), .A2(n3258), .A3(n3257), .A4(n3256), .ZN(n3346)
         );
  AND2_X2 U3717 ( .A1(n5477), .A2(n3963), .ZN(n5468) );
  NAND2_X1 U3718 ( .A1(n3334), .A2(n3350), .ZN(n3336) );
  INV_X1 U3719 ( .A(n3471), .ZN(n3506) );
  AND2_X2 U3720 ( .A1(n3130), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3192)
         );
  INV_X1 U3721 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3130) );
  NAND2_X1 U3722 ( .A1(n3345), .A2(n3115), .ZN(n4297) );
  INV_X1 U3723 ( .A(n3501), .ZN(n3502) );
  OR2_X1 U3724 ( .A1(n3673), .A2(n3672), .ZN(n4547) );
  AND2_X1 U3725 ( .A1(n4202), .A2(n3671), .ZN(n3672) );
  AOI21_X1 U3726 ( .B1(n3670), .B2(n4202), .A(n3669), .ZN(n3673) );
  OAI22_X1 U3727 ( .A1(n3668), .A2(n3667), .B1(n3666), .B2(n4196), .ZN(n3669)
         );
  INV_X1 U3728 ( .A(n6095), .ZN(n5113) );
  AOI21_X1 U3729 ( .B1(n4643), .B2(n3636), .A(n3474), .ZN(n6221) );
  NAND2_X1 U3730 ( .A1(n4776), .A2(n4775), .ZN(n4984) );
  AND2_X1 U3731 ( .A1(n4349), .A2(n4341), .ZN(n5753) );
  INV_X1 U3732 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U3733 ( .A1(n5033), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3627) );
  NAND2_X1 U3734 ( .A1(n3638), .A2(n3627), .ZN(n3647) );
  AND2_X1 U3735 ( .A1(n3629), .A2(n3628), .ZN(n3646) );
  AOI21_X1 U3736 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6681), .A(n3635), 
        .ZN(n3664) );
  AND2_X1 U3737 ( .A1(n3295), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3203) );
  INV_X1 U3738 ( .A(n3532), .ZN(n3534) );
  NAND2_X1 U3739 ( .A1(n3346), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3490) );
  INV_X1 U3740 ( .A(n5433), .ZN(n4113) );
  NAND2_X1 U3741 ( .A1(n6541), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4133) );
  OR2_X1 U3742 ( .A1(n3457), .A2(n3456), .ZN(n3471) );
  AND2_X1 U3743 ( .A1(n3352), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U3744 ( .A1(n3154), .A2(n3152), .ZN(n3621) );
  NOR2_X1 U3745 ( .A1(n3155), .A2(n3153), .ZN(n3152) );
  INV_X1 U3746 ( .A(n3617), .ZN(n3153) );
  INV_X1 U3747 ( .A(n3125), .ZN(n3155) );
  NAND2_X1 U3748 ( .A1(n3317), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3590) );
  NOR2_X1 U3749 ( .A1(n5241), .A2(n5240), .ZN(n5239) );
  OR2_X1 U3750 ( .A1(n3151), .A2(n3599), .ZN(n3150) );
  INV_X1 U3751 ( .A(n5245), .ZN(n3151) );
  NAND2_X1 U3752 ( .A1(n3411), .A2(n3427), .ZN(n3416) );
  NAND2_X1 U3753 ( .A1(n3441), .A2(n3440), .ZN(n3482) );
  AOI21_X1 U3754 ( .B1(n6578), .B2(n4613), .A(n5386), .ZN(n4709) );
  INV_X1 U3755 ( .A(n5038), .ZN(n5128) );
  AND2_X1 U3756 ( .A1(n4596), .A2(n4595), .ZN(n6550) );
  NOR2_X1 U3757 ( .A1(n6092), .A2(n4401), .ZN(n5270) );
  CLKBUF_X1 U3758 ( .A(n4334), .Z(n4686) );
  NAND2_X1 U3759 ( .A1(n3171), .A2(n4009), .ZN(n3170) );
  INV_X1 U3760 ( .A(n4372), .ZN(n3171) );
  INV_X1 U3761 ( .A(n5461), .ZN(n3169) );
  AND2_X1 U3762 ( .A1(n3762), .A2(n4773), .ZN(n3174) );
  BUF_X4 U3763 ( .A(n4230), .Z(n5683) );
  NAND2_X1 U3764 ( .A1(n3145), .A2(n3143), .ZN(n5580) );
  AOI21_X1 U3765 ( .B1(n3147), .B2(n3144), .A(n3123), .ZN(n3143) );
  OR2_X1 U3766 ( .A1(n5348), .A2(n3148), .ZN(n3145) );
  NAND2_X1 U3767 ( .A1(n5185), .A2(n5184), .ZN(n5241) );
  INV_X1 U3768 ( .A(n4730), .ZN(n3133) );
  NOR2_X1 U3769 ( .A1(n6238), .A2(n6310), .ZN(n5599) );
  NAND2_X1 U3770 ( .A1(n4211), .A2(n4210), .ZN(n4349) );
  INV_X1 U3771 ( .A(n4547), .ZN(n4530) );
  INV_X1 U3772 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4616) );
  AOI22_X1 U3773 ( .A1(n3299), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3279) );
  AND2_X1 U3774 ( .A1(n4990), .A2(n4863), .ZN(n4867) );
  OR3_X1 U3775 ( .A1(n6662), .A2(STATE2_REG_0__SCAN_IN), .A3(n4709), .ZN(n4854) );
  AOI21_X1 U3776 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6372), .A(n5128), .ZN(
        n6414) );
  AND2_X1 U3777 ( .A1(n4616), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3674) );
  INV_X1 U3778 ( .A(n3711), .ZN(n4165) );
  INV_X1 U3779 ( .A(n4438), .ZN(n4439) );
  AND2_X1 U3780 ( .A1(n4434), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4393) );
  INV_X1 U3781 ( .A(n6083), .ZN(n6109) );
  AND2_X1 U3782 ( .A1(n5412), .A2(n4428), .ZN(n6107) );
  AND2_X1 U3783 ( .A1(n5396), .A2(n4698), .ZN(n6134) );
  INV_X1 U3784 ( .A(n5396), .ZN(n6133) );
  INV_X1 U3785 ( .A(n5955), .ZN(n6218) );
  NAND2_X1 U3786 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  OAI21_X1 U3787 ( .B1(n3159), .B2(n3129), .A(n3624), .ZN(n3625) );
  XNOR2_X1 U3788 ( .A(n4188), .B(n4365), .ZN(n4370) );
  NAND2_X1 U3789 ( .A1(n4187), .A2(n4186), .ZN(n4188) );
  INV_X1 U3790 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6372) );
  INV_X1 U3791 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6554) );
  INV_X1 U3792 ( .A(n3670), .ZN(n3658) );
  NOR2_X1 U3793 ( .A1(n3345), .A2(n4195), .ZN(n3357) );
  NOR2_X1 U3794 ( .A1(n4690), .A2(n3317), .ZN(n3333) );
  OR2_X1 U3795 ( .A1(n3346), .A2(n6576), .ZN(n3643) );
  NAND2_X1 U3796 ( .A1(n3630), .A2(n3629), .ZN(n3633) );
  XNOR2_X1 U3797 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3632) );
  INV_X1 U3798 ( .A(n3555), .ZN(n3557) );
  OR2_X1 U3799 ( .A1(n3544), .A2(n3543), .ZN(n3571) );
  OR2_X1 U3800 ( .A1(n3522), .A2(n3521), .ZN(n3547) );
  NAND2_X1 U3801 ( .A1(n3272), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3181)
         );
  OR2_X1 U3802 ( .A1(n3500), .A2(n3499), .ZN(n3525) );
  AOI22_X1 U3803 ( .A1(n3306), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3299), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U3804 ( .A1(n3305), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3236) );
  AOI22_X1 U3805 ( .A1(n3380), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3235) );
  AOI221_X1 U3806 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3664), .C1(
        n6802), .C2(n3664), .A(n3631), .ZN(n4202) );
  INV_X1 U3807 ( .A(n3671), .ZN(n3666) );
  NAND2_X1 U3808 ( .A1(n3590), .A2(n3490), .ZN(n3670) );
  NOR2_X1 U3809 ( .A1(n3116), .A2(n3345), .ZN(n3343) );
  NOR2_X1 U3810 ( .A1(n6883), .A2(n5329), .ZN(n5370) );
  NOR2_X1 U3811 ( .A1(n4420), .A2(n5683), .ZN(n4233) );
  AND2_X1 U3812 ( .A1(n4339), .A2(n6584), .ZN(n3338) );
  NAND2_X1 U3813 ( .A1(n3209), .A2(n3208), .ZN(n3351) );
  INV_X1 U3814 ( .A(n5462), .ZN(n4009) );
  NAND2_X1 U3815 ( .A1(n5694), .A2(n3615), .ZN(n3154) );
  AND2_X1 U3816 ( .A1(n4299), .A2(n5697), .ZN(n5700) );
  NAND2_X1 U3817 ( .A1(n5349), .A2(n5350), .ZN(n3149) );
  INV_X1 U3818 ( .A(n5350), .ZN(n3144) );
  NAND2_X1 U3819 ( .A1(n3142), .A2(n3160), .ZN(n4532) );
  INV_X1 U3820 ( .A(n3675), .ZN(n3142) );
  AND2_X1 U3821 ( .A1(n3337), .A2(n3351), .ZN(n4335) );
  AND2_X2 U3822 ( .A1(n3132), .A2(n3131), .ZN(n4524) );
  INV_X1 U3823 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3132) );
  INV_X1 U3824 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3131) );
  AND2_X2 U3825 ( .A1(n4598), .A2(n4523), .ZN(n3272) );
  INV_X1 U3826 ( .A(n4990), .ZN(n6326) );
  AOI22_X1 U3827 ( .A1(n3307), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3273) );
  INV_X1 U3828 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5033) );
  INV_X1 U3829 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6762) );
  NAND2_X1 U3830 ( .A1(n4477), .A2(n4388), .ZN(n4493) );
  INV_X1 U3831 ( .A(n4537), .ZN(n4388) );
  AND4_X1 U3832 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .A4(n5900), .ZN(n5868) );
  AND2_X1 U3833 ( .A1(n4311), .A2(n4310), .ZN(n5472) );
  INV_X1 U3834 ( .A(n5422), .ZN(n3161) );
  INV_X1 U3835 ( .A(n3346), .ZN(n3135) );
  AOI22_X1 U3836 ( .A1(n4169), .A2(n4168), .B1(n4437), .B2(n4165), .ZN(n4385)
         );
  NAND2_X1 U3837 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4173)
         );
  AND2_X1 U3838 ( .A1(n4087), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4109)
         );
  AOI21_X1 U3839 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n5443) );
  AND2_X1 U3840 ( .A1(n5834), .A2(n4165), .ZN(n4066) );
  OR2_X1 U3841 ( .A1(n4023), .A2(n6822), .ZN(n4046) );
  OR2_X1 U3842 ( .A1(n4046), .A2(n4045), .ZN(n4086) );
  AND2_X1 U3843 ( .A1(n3980), .A2(n3979), .ZN(n5469) );
  NOR2_X1 U3844 ( .A1(n3977), .A2(n6841), .ZN(n4005) );
  AND2_X1 U3845 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3959), .ZN(n3960)
         );
  INV_X1 U3846 ( .A(n3958), .ZN(n3959) );
  NAND2_X1 U3847 ( .A1(n3960), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3977)
         );
  NOR2_X1 U3848 ( .A1(n5559), .A2(n3924), .ZN(n3925) );
  NAND2_X1 U3849 ( .A1(n3925), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3958)
         );
  NAND2_X1 U3850 ( .A1(n3168), .A2(n3909), .ZN(n3167) );
  INV_X1 U3851 ( .A(n5897), .ZN(n3168) );
  INV_X1 U3852 ( .A(n5561), .ZN(n3166) );
  NOR2_X1 U3853 ( .A1(n3889), .A2(n5569), .ZN(n3890) );
  NAND2_X1 U3854 ( .A1(n3890), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3924)
         );
  NAND2_X1 U3855 ( .A1(n3859), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3889)
         );
  CLKBUF_X1 U3856 ( .A(n5366), .Z(n5367) );
  AND2_X1 U3857 ( .A1(n3841), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3859)
         );
  AND2_X1 U3858 ( .A1(n3840), .A2(n5255), .ZN(n3173) );
  NAND2_X1 U3859 ( .A1(n3811), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3825)
         );
  NOR2_X1 U3860 ( .A1(n3796), .A2(n6032), .ZN(n3811) );
  NAND2_X1 U3861 ( .A1(n3780), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3796)
         );
  INV_X1 U3862 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6032) );
  CLKBUF_X1 U3863 ( .A(n5171), .Z(n5172) );
  NOR2_X1 U3864 ( .A1(n3763), .A2(n6051), .ZN(n3780) );
  NOR2_X1 U3865 ( .A1(n6778), .A2(n3729), .ZN(n3747) );
  NOR2_X1 U3866 ( .A1(n3721), .A2(n5098), .ZN(n3722) );
  NAND2_X1 U3867 ( .A1(n3722), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3729)
         );
  NAND2_X1 U3868 ( .A1(n6210), .A2(n3531), .ZN(n3141) );
  INV_X1 U3869 ( .A(n4630), .ZN(n3172) );
  NOR2_X1 U3870 ( .A1(n3699), .A2(n4653), .ZN(n3713) );
  NAND2_X1 U3871 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U3872 ( .A1(n3687), .A2(n3686), .ZN(n4463) );
  NAND2_X1 U3873 ( .A1(n4224), .A2(n5683), .ZN(n5407) );
  AND2_X1 U3874 ( .A1(n3619), .A2(n3158), .ZN(n3157) );
  INV_X1 U3875 ( .A(n5602), .ZN(n3158) );
  NOR2_X1 U3876 ( .A1(n5554), .A2(n5520), .ZN(n3619) );
  AND2_X1 U3877 ( .A1(n3602), .A2(n3175), .ZN(n4185) );
  AND2_X1 U3878 ( .A1(n3602), .A2(n6774), .ZN(n4184) );
  AND2_X1 U3879 ( .A1(n4273), .A2(n4272), .ZN(n5240) );
  NAND2_X1 U3880 ( .A1(n4263), .A2(n4262), .ZN(n5090) );
  NAND2_X1 U3881 ( .A1(n4248), .A2(n3178), .ZN(n4684) );
  AND2_X1 U3882 ( .A1(n4252), .A2(n4251), .ZN(n4780) );
  INV_X1 U3883 ( .A(n3134), .ZN(n4782) );
  NAND2_X1 U3884 ( .A1(n3353), .A2(n3352), .ZN(n4221) );
  CLKBUF_X1 U3885 ( .A(n4632), .Z(n4683) );
  INV_X1 U3886 ( .A(n6219), .ZN(n3477) );
  INV_X1 U3887 ( .A(n6288), .ZN(n6310) );
  AND2_X1 U3888 ( .A1(n4352), .A2(n4351), .ZN(n6239) );
  INV_X1 U3889 ( .A(n5407), .ZN(n4472) );
  INV_X1 U3890 ( .A(n3317), .ZN(n4220) );
  NAND2_X1 U3891 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U3892 ( .A(n3482), .B(n3483), .ZN(n4590) );
  INV_X1 U3893 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4582) );
  NAND2_X1 U3894 ( .A1(n3484), .A2(n3483), .ZN(n4603) );
  AND3_X1 U3895 ( .A1(n4550), .A2(n4549), .A3(n4548), .ZN(n6544) );
  NOR2_X1 U3896 ( .A1(n5191), .A2(n4993), .ZN(n5044) );
  OR2_X1 U3897 ( .A1(n6323), .A2(n4993), .ZN(n4800) );
  AND2_X1 U3898 ( .A1(n4702), .A2(n6677), .ZN(n5283) );
  INV_X1 U3899 ( .A(n5043), .ZN(n4994) );
  INV_X1 U3900 ( .A(n3321), .ZN(n3337) );
  OR2_X1 U3901 ( .A1(n4443), .A2(n6581), .ZN(n5805) );
  INV_X1 U3902 ( .A(n5508), .ZN(n5817) );
  NOR2_X1 U3903 ( .A1(n6637), .A2(n5886), .ZN(n5881) );
  INV_X1 U3904 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6051) );
  INV_X1 U3905 ( .A(n6044), .ZN(n6064) );
  INV_X1 U3906 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5098) );
  AND2_X1 U3907 ( .A1(n5093), .A2(n6044), .ZN(n6116) );
  INV_X1 U3908 ( .A(n5456), .ZN(n6125) );
  INV_X1 U3909 ( .A(n7016), .ZN(n5454) );
  AND2_X1 U3910 ( .A1(n7016), .A2(n5395), .ZN(n6124) );
  AND2_X2 U3911 ( .A1(n4460), .A2(n6583), .ZN(n7016) );
  INV_X1 U3912 ( .A(n6124), .ZN(n7014) );
  INV_X1 U3913 ( .A(n5820), .ZN(n5491) );
  OR2_X1 U3914 ( .A1(n6130), .A2(n6134), .ZN(n5363) );
  NAND2_X1 U3915 ( .A1(n6174), .A2(n4689), .ZN(n5396) );
  OAI21_X1 U3916 ( .B1(n4688), .B2(n4687), .A(n6583), .ZN(n4689) );
  INV_X1 U3917 ( .A(n5363), .ZN(n5088) );
  AND2_X1 U3918 ( .A1(n4480), .A2(n4479), .ZN(n6161) );
  INV_X1 U3919 ( .A(n6161), .ZN(n6166) );
  INV_X1 U3920 ( .A(n6193), .ZN(n6187) );
  XNOR2_X1 U3921 ( .A(n4174), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4434)
         );
  OR2_X1 U3922 ( .A1(n4173), .A2(n4429), .ZN(n4174) );
  INV_X1 U3923 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n6841) );
  INV_X1 U3924 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5559) );
  INV_X1 U3925 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5569) );
  INV_X1 U3926 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U3927 ( .A1(n5955), .A2(n4487), .ZN(n6228) );
  INV_X1 U3928 ( .A(n6228), .ZN(n6196) );
  XNOR2_X1 U3929 ( .A(n5498), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5631)
         );
  NAND2_X1 U3930 ( .A1(n5496), .A2(n3159), .ZN(n5498) );
  AND2_X1 U3931 ( .A1(n5706), .A2(n5526), .ZN(n5663) );
  AND2_X1 U3932 ( .A1(n5668), .A2(n5674), .ZN(n5666) );
  AND2_X1 U3933 ( .A1(n5717), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5706)
         );
  CLKBUF_X1 U3934 ( .A(n5694), .Z(n5695) );
  CLKBUF_X1 U3935 ( .A(n5580), .Z(n5581) );
  NAND2_X1 U3936 ( .A1(n3146), .A2(n5350), .ZN(n5591) );
  OR2_X1 U3937 ( .A1(n5348), .A2(n5349), .ZN(n3146) );
  CLKBUF_X1 U3938 ( .A(n5340), .Z(n5341) );
  NAND2_X1 U3939 ( .A1(n5175), .A2(n3599), .ZN(n5248) );
  CLKBUF_X1 U3940 ( .A(n4657), .Z(n4658) );
  INV_X1 U3941 ( .A(n6292), .ZN(n6317) );
  INV_X1 U3942 ( .A(n6283), .ZN(n6292) );
  CLKBUF_X1 U3943 ( .A(n4647), .Z(n4648) );
  AND2_X1 U3944 ( .A1(n4349), .A2(n6543), .ZN(n5749) );
  CLKBUF_X1 U3945 ( .A(n4518), .Z(n4519) );
  CLKBUF_X1 U3946 ( .A(n4590), .Z(n4591) );
  INV_X1 U3947 ( .A(n6679), .ZN(n6682) );
  INV_X1 U3948 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5388) );
  NOR2_X1 U3949 ( .A1(n6662), .A2(n4530), .ZN(n5386) );
  NAND2_X1 U3950 ( .A1(n6662), .A2(n4616), .ZN(n6670) );
  INV_X1 U3951 ( .A(n4830), .ZN(n5799) );
  INV_X1 U3952 ( .A(n6358), .ZN(n4923) );
  NOR2_X1 U3953 ( .A1(n5191), .A2(n6366), .ZN(n6358) );
  OR2_X1 U3954 ( .A1(n4995), .A2(n5043), .ZN(n6373) );
  INV_X1 U3955 ( .A(n6498), .ZN(n6451) );
  NOR2_X1 U3956 ( .A1(n4800), .A2(n5043), .ZN(n5282) );
  INV_X1 U3957 ( .A(n6419), .ZN(n6502) );
  INV_X1 U3958 ( .A(n6422), .ZN(n6508) );
  INV_X1 U3959 ( .A(n6426), .ZN(n6468) );
  INV_X1 U3960 ( .A(n6429), .ZN(n6514) );
  INV_X1 U3961 ( .A(n6432), .ZN(n6520) );
  INV_X1 U3962 ( .A(n6439), .ZN(n6526) );
  INV_X1 U3963 ( .A(n6445), .ZN(n6535) );
  AND3_X1 U3964 ( .A1(n4870), .A2(n6414), .A3(n4869), .ZN(n4906) );
  NOR2_X1 U3965 ( .A1(n4854), .A2(n3421), .ZN(n6467) );
  NOR2_X1 U3966 ( .A1(n4854), .A2(n4765), .ZN(n6513) );
  NOR2_X1 U3967 ( .A1(n4854), .A2(n3317), .ZN(n6519) );
  NOR2_X1 U3968 ( .A1(n4747), .A2(n4994), .ZN(n4967) );
  NOR2_X1 U3969 ( .A1(n4854), .A2(n5395), .ZN(n6533) );
  INV_X1 U3970 ( .A(n6501), .ZN(n5170) );
  INV_X1 U3971 ( .A(n6507), .ZN(n5158) );
  INV_X1 U3972 ( .A(n6467), .ZN(n5142) );
  INV_X1 U3973 ( .A(n6519), .ZN(n5146) );
  INV_X1 U3974 ( .A(n6481), .ZN(n5154) );
  INV_X1 U3975 ( .A(n6525), .ZN(n5150) );
  INV_X1 U3976 ( .A(n4967), .ZN(n4930) );
  OR2_X1 U3977 ( .A1(n4747), .A2(n5043), .ZN(n5067) );
  INV_X1 U3978 ( .A(n6533), .ZN(n5138) );
  INV_X1 U3979 ( .A(n6701), .ZN(n6578) );
  AND2_X1 U3980 ( .A1(n6566), .A2(n6565), .ZN(n6582) );
  AND2_X1 U3981 ( .A1(n3674), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6583) );
  INV_X1 U3982 ( .A(n6589), .ZN(n6661) );
  INV_X1 U3983 ( .A(n5985), .ZN(n6659) );
  NOR2_X1 U3984 ( .A1(n6838), .A2(STATE_REG_0__SCAN_IN), .ZN(n6706) );
  NOR2_X1 U3985 ( .A1(n4429), .A2(n6109), .ZN(n4440) );
  OAI21_X1 U3986 ( .B1(n5855), .B2(n6211), .A(n4377), .ZN(n4378) );
  AOI21_X1 U3987 ( .B1(n5420), .B2(n5611), .A(n5610), .ZN(n5612) );
  INV_X1 U3988 ( .A(n5609), .ZN(n5610) );
  AOI21_X1 U3989 ( .B1(n5608), .B2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5607), 
        .ZN(n5609) );
  NAND2_X1 U3990 ( .A1(n5235), .A2(n5255), .ZN(n5254) );
  NAND2_X1 U3991 ( .A1(n3166), .A2(n3909), .ZN(n5560) );
  NAND2_X1 U3992 ( .A1(n3169), .A2(n4009), .ZN(n4371) );
  INV_X1 U3993 ( .A(n3159), .ZN(n5497) );
  NAND2_X1 U3994 ( .A1(n3620), .A2(n3157), .ZN(n3159) );
  NAND2_X1 U3995 ( .A1(n3593), .A2(n3592), .ZN(n3602) );
  NAND2_X1 U3996 ( .A1(n4771), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U3997 ( .A1(n5235), .A2(n3173), .ZN(n5325) );
  INV_X1 U3998 ( .A(n4233), .ZN(n4240) );
  NAND2_X1 U3999 ( .A1(n3154), .A2(n3617), .ZN(n5503) );
  AND4_X1 U4000 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3118)
         );
  NAND2_X1 U4001 ( .A1(n3447), .A2(n3446), .ZN(n3483) );
  OR2_X1 U4002 ( .A1(n3590), .A2(n3417), .ZN(n3119) );
  INV_X1 U4003 ( .A(n3345), .ZN(n4752) );
  OR2_X1 U4004 ( .A1(n5391), .A2(n5564), .ZN(n3120) );
  NAND2_X1 U4005 ( .A1(n3620), .A2(n3619), .ZN(n5512) );
  OR2_X1 U4006 ( .A1(n5453), .A2(n5444), .ZN(n3121) );
  XNOR2_X1 U4008 ( .A(n3163), .B(n3162), .ZN(n5419) );
  AND3_X1 U4009 ( .A1(n3340), .A2(n3339), .A3(n3338), .ZN(n3122) );
  AND2_X1 U4010 ( .A1(n5582), .A2(n6949), .ZN(n3123) );
  AND2_X1 U4011 ( .A1(n3150), .A2(n5246), .ZN(n3124) );
  NAND2_X1 U4012 ( .A1(n4381), .A2(n4382), .ZN(n5496) );
  INV_X1 U4013 ( .A(n3148), .ZN(n3147) );
  NAND2_X1 U4014 ( .A1(n5590), .A2(n3149), .ZN(n3148) );
  OAI22_X1 U4015 ( .A1(n5580), .A2(n3607), .B1(n5582), .B2(n3606), .ZN(n5575)
         );
  AND2_X1 U4016 ( .A1(n3345), .A2(n3320), .ZN(n3636) );
  XOR2_X1 U4017 ( .A(n5582), .B(n6788), .Z(n3125) );
  INV_X1 U4018 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6576) );
  AND2_X1 U4019 ( .A1(n4324), .A2(n3135), .ZN(n3126) );
  NAND2_X1 U4020 ( .A1(n5582), .A2(n3610), .ZN(n3127) );
  AND2_X1 U4021 ( .A1(n3161), .A2(n4113), .ZN(n3128) );
  NAND2_X1 U4022 ( .A1(n4349), .A2(n4219), .ZN(n5745) );
  INV_X1 U4023 ( .A(n5745), .ZN(n6315) );
  INV_X1 U4024 ( .A(n5564), .ZN(n6223) );
  NAND2_X1 U4025 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3129) );
  AND2_X2 U4026 ( .A1(n4524), .A2(n3192), .ZN(n3278) );
  AND2_X2 U4027 ( .A1(n3134), .A2(n3133), .ZN(n4776) );
  NOR2_X2 U4028 ( .A1(n4684), .A2(n4780), .ZN(n3134) );
  NOR2_X1 U4029 ( .A1(n4322), .A2(n3135), .ZN(n4193) );
  AOI22_X1 U4030 ( .A1(n5115), .A2(n4322), .B1(n4543), .B2(n3135), .ZN(n3344)
         );
  AOI21_X1 U4031 ( .B1(n6541), .B2(n3320), .A(n3135), .ZN(n3675) );
  NAND2_X1 U4032 ( .A1(n4207), .A2(n3135), .ZN(n4213) );
  OAI22_X1 U4033 ( .A1(n4686), .A2(n4337), .B1(n4336), .B2(n3135), .ZN(n4338)
         );
  NAND2_X1 U4034 ( .A1(n6161), .A2(n3135), .ZN(n4671) );
  NAND3_X1 U4035 ( .A1(n4227), .A2(n3139), .A3(n4226), .ZN(n3136) );
  NAND2_X1 U4036 ( .A1(n3138), .A2(n4471), .ZN(n3137) );
  INV_X1 U4037 ( .A(n4227), .ZN(n3138) );
  INV_X1 U4038 ( .A(n4471), .ZN(n3139) );
  NAND2_X1 U4039 ( .A1(n4226), .A2(n4227), .ZN(n3140) );
  NAND2_X1 U4040 ( .A1(n4466), .A2(n3140), .ZN(n4619) );
  AND2_X2 U4041 ( .A1(n5239), .A2(n4277), .ZN(n5332) );
  NAND2_X2 U4042 ( .A1(n3117), .A2(n5425), .ZN(n5401) );
  OAI21_X1 U4043 ( .B1(n4733), .B2(n3141), .A(n4732), .ZN(n6279) );
  INV_X1 U4044 ( .A(n3603), .ZN(n3601) );
  OAI21_X2 U4045 ( .B1(n5175), .B2(n3151), .A(n3124), .ZN(n3603) );
  NAND2_X1 U4046 ( .A1(n6219), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3475)
         );
  NAND2_X1 U4047 ( .A1(n4647), .A2(n4649), .ZN(n3156) );
  NAND2_X1 U4048 ( .A1(n3425), .A2(n3424), .ZN(n4647) );
  AND3_X2 U4049 ( .A1(n3160), .A2(n3314), .A3(n3339), .ZN(n3327) );
  NAND2_X1 U4050 ( .A1(n5432), .A2(n4113), .ZN(n5435) );
  NAND2_X1 U4051 ( .A1(n5432), .A2(n3128), .ZN(n3165) );
  INV_X1 U4052 ( .A(n4171), .ZN(n3162) );
  INV_X1 U4053 ( .A(n4385), .ZN(n3164) );
  NAND2_X1 U4054 ( .A1(n4629), .A2(n4682), .ZN(n4681) );
  NAND3_X1 U4055 ( .A1(n3706), .A2(n4623), .A3(n4624), .ZN(n4626) );
  NAND2_X1 U4056 ( .A1(n4771), .A2(n3174), .ZN(n4981) );
  INV_X1 U4057 ( .A(n4981), .ZN(n3779) );
  INV_X1 U4058 ( .A(n4404), .ZN(n4442) );
  AND2_X1 U4059 ( .A1(n5435), .A2(n5434), .ZN(n5820) );
  NAND2_X1 U4060 ( .A1(n3359), .A2(n3360), .ZN(n3440) );
  AOI21_X1 U4061 ( .B1(n3442), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3361), 
        .ZN(n3359) );
  NAND2_X1 U4062 ( .A1(n4349), .A2(n4222), .ZN(n6294) );
  AND2_X2 U4063 ( .A1(n4524), .A2(n4598), .ZN(n3295) );
  INV_X1 U4064 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4182) );
  AND2_X1 U4065 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U4066 ( .A1(n6662), .A2(n6334), .ZN(n6694) );
  OR2_X1 U4067 ( .A1(n5407), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3176)
         );
  AOI21_X1 U4068 ( .B1(n4434), .B2(n6196), .A(n4179), .ZN(n4180) );
  INV_X1 U4069 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6778) );
  INV_X1 U4070 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5272) );
  OR2_X1 U4071 ( .A1(n5407), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3177)
         );
  AND2_X1 U4072 ( .A1(n4247), .A2(n4246), .ZN(n3178) );
  INV_X1 U4073 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n3600) );
  INV_X1 U4074 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6802) );
  INV_X1 U4075 ( .A(n3341), .ZN(n3285) );
  OR2_X1 U4076 ( .A1(n3361), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3179)
         );
  NOR2_X1 U4077 ( .A1(n3333), .A2(n4230), .ZN(n3334) );
  NAND2_X1 U4078 ( .A1(n4224), .A2(n4752), .ZN(n3335) );
  NAND2_X1 U4079 ( .A1(n3336), .A2(n3335), .ZN(n3340) );
  NAND2_X1 U4080 ( .A1(n3647), .A2(n3646), .ZN(n3630) );
  NAND2_X1 U4081 ( .A1(n6762), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3629) );
  INV_X1 U4082 ( .A(n4198), .ZN(n3662) );
  INV_X1 U4083 ( .A(n3470), .ZN(n3391) );
  OR2_X1 U4084 ( .A1(n3637), .A2(n3641), .ZN(n3638) );
  INV_X1 U4085 ( .A(n4982), .ZN(n3762) );
  AND2_X1 U4086 ( .A1(n3633), .A2(n3632), .ZN(n3635) );
  OR2_X1 U4087 ( .A1(n3377), .A2(n3376), .ZN(n3470) );
  NAND2_X1 U4088 ( .A1(n3439), .A2(n3438), .ZN(n3441) );
  INV_X1 U4089 ( .A(n3296), .ZN(n3304) );
  AND2_X1 U4090 ( .A1(n3182), .A2(n3181), .ZN(n3188) );
  INV_X1 U4091 ( .A(n5562), .ZN(n3909) );
  INV_X1 U4092 ( .A(n5362), .ZN(n3857) );
  INV_X1 U4093 ( .A(n5326), .ZN(n3840) );
  INV_X1 U4094 ( .A(n5085), .ZN(n3778) );
  OR2_X1 U4095 ( .A1(n3567), .A2(n3566), .ZN(n3583) );
  INV_X1 U4096 ( .A(n4324), .ZN(n3352) );
  AOI21_X1 U4097 ( .B1(n4154), .B2(INSTQUEUE_REG_8__7__SCAN_IN), .A(n3203), 
        .ZN(n3207) );
  INV_X1 U4098 ( .A(n4027), .ZN(n4167) );
  INV_X1 U4099 ( .A(n4779), .ZN(n3728) );
  NOR2_X1 U4100 ( .A1(n4086), .A2(n5522), .ZN(n4087) );
  OR2_X1 U4101 ( .A1(n5867), .A2(n3711), .ZN(n4007) );
  INV_X1 U4102 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3476) );
  AND2_X1 U4103 ( .A1(n3665), .A2(n3636), .ZN(n3671) );
  INV_X1 U4104 ( .A(n5258), .ZN(n4277) );
  OR2_X1 U4105 ( .A1(n3408), .A2(n3407), .ZN(n3469) );
  INV_X1 U4106 ( .A(n3320), .ZN(n3288) );
  INV_X1 U4107 ( .A(n3691), .ZN(n4027) );
  NOR2_X1 U4108 ( .A1(n5406), .A2(n5698), .ZN(n4412) );
  INV_X1 U4109 ( .A(n4985), .ZN(n4262) );
  AND4_X1 U4110 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3208)
         );
  AND2_X1 U4111 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4135)
         );
  AND2_X1 U4112 ( .A1(n4050), .A2(n4049), .ZN(n5448) );
  NOR2_X1 U4113 ( .A1(n3825), .A2(n5272), .ZN(n3841) );
  NAND2_X1 U4114 ( .A1(n3317), .A2(n3320), .ZN(n3341) );
  AND2_X1 U4115 ( .A1(n4296), .A2(n4295), .ZN(n5702) );
  NOR2_X1 U4116 ( .A1(n4344), .A2(n4343), .ZN(n4571) );
  INV_X1 U4117 ( .A(n5769), .ZN(n5797) );
  INV_X1 U4118 ( .A(n6677), .ZN(n6454) );
  OR2_X1 U4119 ( .A1(n4864), .A2(n4591), .ZN(n4824) );
  INV_X1 U4120 ( .A(n5129), .ZN(n5164) );
  AND2_X1 U4121 ( .A1(n3444), .A2(n6328), .ZN(n4935) );
  OR2_X1 U4122 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3711) );
  INV_X1 U4123 ( .A(n3870), .ZN(n4170) );
  AND2_X1 U4124 ( .A1(n4307), .A2(n4306), .ZN(n5481) );
  INV_X1 U4125 ( .A(n6105), .ZN(n5901) );
  NAND2_X1 U4126 ( .A1(n3747), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3763)
         );
  AND3_X1 U4127 ( .A1(n6292), .A2(n4391), .A3(n6587), .ZN(n4392) );
  INV_X2 U4128 ( .A(n4230), .ZN(n5698) );
  AND2_X1 U4129 ( .A1(n4268), .A2(n4267), .ZN(n5089) );
  OR2_X1 U4130 ( .A1(n4135), .A2(n4110), .ZN(n5508) );
  AOI21_X1 U4131 ( .B1(n3727), .B2(n3677), .A(n3726), .ZN(n4779) );
  OR2_X1 U4133 ( .A1(n6670), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6695) );
  OR2_X1 U4134 ( .A1(n5749), .A2(n5753), .ZN(n6238) );
  NAND2_X1 U4135 ( .A1(n3430), .A2(n3429), .ZN(n3688) );
  INV_X1 U4136 ( .A(n3365), .ZN(n4569) );
  OR2_X1 U4137 ( .A1(n6453), .A2(n6677), .ZN(n5767) );
  OR2_X1 U4138 ( .A1(n3682), .A2(n4990), .ZN(n5191) );
  AND2_X1 U4139 ( .A1(n6414), .A2(n4998), .ZN(n5026) );
  OR2_X1 U4140 ( .A1(n4995), .A2(n4994), .ZN(n5230) );
  INV_X1 U4141 ( .A(n5282), .ZN(n5313) );
  INV_X1 U4142 ( .A(n4873), .ZN(n4907) );
  AND2_X1 U4143 ( .A1(n4591), .A2(n4519), .ZN(n6376) );
  INV_X1 U4144 ( .A(n4493), .ZN(n5804) );
  AOI22_X1 U4145 ( .A1(n4167), .A2(EAX_REG_31__SCAN_IN), .B1(n4170), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4171) );
  NOR2_X1 U4146 ( .A1(n5854), .A2(n4402), .ZN(n5830) );
  NAND2_X1 U4147 ( .A1(n4005), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4023)
         );
  NOR2_X1 U4148 ( .A1(n6635), .A2(n5902), .ZN(n5896) );
  INV_X1 U4149 ( .A(n6067), .ZN(n6041) );
  NOR2_X2 U4150 ( .A1(n6095), .A2(n4436), .ZN(n6096) );
  INV_X1 U4151 ( .A(n5916), .ZN(n6131) );
  INV_X1 U4152 ( .A(n4671), .ZN(n6141) );
  INV_X1 U4153 ( .A(n6696), .ZN(n6567) );
  NAND2_X1 U4154 ( .A1(n5804), .A2(n4497), .ZN(n6174) );
  INV_X1 U4155 ( .A(n6174), .ZN(n6190) );
  NAND2_X1 U4156 ( .A1(n3713), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3721)
         );
  INV_X1 U4157 ( .A(n6213), .ZN(n6224) );
  INV_X1 U4158 ( .A(n6294), .ZN(n5611) );
  AND2_X1 U4159 ( .A1(n5663), .A2(n5601), .ZN(n5956) );
  INV_X1 U4160 ( .A(n5736), .ZN(n5967) );
  AND2_X1 U4161 ( .A1(n6310), .A2(n4353), .ZN(n5752) );
  NAND2_X1 U4162 ( .A1(n4813), .A2(n4812), .ZN(n4811) );
  NOR2_X1 U4163 ( .A1(n6695), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6283) );
  AND2_X1 U4164 ( .A1(n4342), .A2(n6238), .ZN(n6318) );
  AND2_X1 U4165 ( .A1(n4192), .A2(n4323), .ZN(n6543) );
  OAI211_X1 U4166 ( .C1(n5041), .C2(n6662), .A(n5040), .B(n6455), .ZN(n5066)
         );
  OAI21_X1 U4167 ( .B1(n4828), .B2(n4827), .A(n6380), .ZN(n4922) );
  INV_X1 U4168 ( .A(n6373), .ZN(n6400) );
  INV_X1 U4169 ( .A(n6404), .ZN(n6440) );
  NOR2_X2 U4170 ( .A1(n4800), .A2(n4994), .ZN(n6494) );
  NOR2_X1 U4171 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4709), .ZN(n5038) );
  NAND2_X1 U4172 ( .A1(n3682), .A2(n6326), .ZN(n6323) );
  INV_X1 U4173 ( .A(n6436), .ZN(n6482) );
  AND2_X1 U4174 ( .A1(n4867), .A2(n4994), .ZN(n4966) );
  NOR2_X1 U4175 ( .A1(n4854), .A2(n3346), .ZN(n6501) );
  NOR2_X1 U4176 ( .A1(n4854), .A2(n4752), .ZN(n6507) );
  NOR2_X1 U4177 ( .A1(n4854), .A2(n3289), .ZN(n6481) );
  INV_X1 U4178 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6593) );
  INV_X1 U4179 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6777) );
  AND2_X1 U4180 ( .A1(n4493), .A2(n5805), .ZN(n6693) );
  INV_X1 U4181 ( .A(n6110), .ZN(n6049) );
  NAND2_X1 U4182 ( .A1(n5113), .A2(n4393), .ZN(n6044) );
  INV_X1 U4183 ( .A(n6107), .ZN(n6104) );
  NAND2_X1 U4184 ( .A1(n7016), .A2(n4697), .ZN(n5456) );
  INV_X1 U4185 ( .A(n5322), .ZN(n6045) );
  NAND2_X1 U4186 ( .A1(n5396), .A2(n4691), .ZN(n5916) );
  INV_X1 U4187 ( .A(n6146), .ZN(n6164) );
  OR2_X1 U4188 ( .A1(n6161), .A2(n6567), .ZN(n6146) );
  INV_X1 U4189 ( .A(n6157), .ZN(n6696) );
  NAND2_X1 U4190 ( .A1(n4477), .A2(n4476), .ZN(n6193) );
  INV_X1 U4191 ( .A(n4378), .ZN(n4379) );
  NAND2_X1 U4192 ( .A1(n6213), .A2(n4176), .ZN(n5955) );
  INV_X1 U4193 ( .A(n6223), .ZN(n6211) );
  OR2_X1 U4194 ( .A1(n6590), .A2(n6694), .ZN(n5564) );
  NAND2_X2 U4195 ( .A1(n4477), .A2(n6557), .ZN(n6213) );
  AND2_X1 U4196 ( .A1(n5666), .A2(n4362), .ZN(n5961) );
  AOI21_X1 U4197 ( .B1(n4354), .B2(n6318), .A(n5752), .ZN(n6236) );
  INV_X1 U4198 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6681) );
  AOI22_X1 U4199 ( .A1(n5772), .A2(n5770), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5768), .ZN(n5803) );
  AOI21_X1 U4200 ( .B1(n6694), .B2(n6335), .A(n6332), .ZN(n6365) );
  OR2_X1 U4201 ( .A1(n6411), .A2(n6366), .ZN(n6404) );
  OR2_X1 U4202 ( .A1(n6411), .A2(n6409), .ZN(n6498) );
  AOI21_X1 U4203 ( .B1(n5286), .B2(n5283), .A(n5280), .ZN(n5317) );
  OR2_X1 U4204 ( .A1(n6323), .A2(n6409), .ZN(n6539) );
  INV_X1 U4205 ( .A(n6513), .ZN(n5162) );
  AND2_X1 U4206 ( .A1(n6573), .A2(n6572), .ZN(n6589) );
  INV_X1 U4207 ( .A(n6659), .ZN(n6592) );
  INV_X1 U4208 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6838) );
  INV_X1 U4209 ( .A(n6651), .ZN(n6648) );
  NAND2_X1 U4210 ( .A1(n4442), .A2(n4441), .ZN(U2797) );
  INV_X1 U4211 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3180) );
  AND2_X4 U4212 ( .A1(n4531), .A2(n3192), .ZN(n3277) );
  NAND2_X1 U4213 ( .A1(n3277), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3182) );
  AND2_X2 U4214 ( .A1(n3183), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3190)
         );
  AND2_X2 U4215 ( .A1(n3190), .A2(n4598), .ZN(n3370) );
  AND2_X2 U4216 ( .A1(n3191), .A2(n4523), .ZN(n3270) );
  AOI22_X1 U4217 ( .A1(n3370), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3187) );
  INV_X1 U4218 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3184) );
  AND2_X2 U4219 ( .A1(n4531), .A2(n3189), .ZN(n3305) );
  AND2_X2 U4220 ( .A1(n3189), .A2(n4523), .ZN(n3306) );
  AOI22_X1 U4221 ( .A1(n3305), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3186) );
  AND2_X2 U4222 ( .A1(n4531), .A2(n4598), .ZN(n3307) );
  AND2_X2 U4223 ( .A1(n3190), .A2(n3191), .ZN(n3402) );
  AOI22_X1 U4224 ( .A1(n3307), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4226 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3299), .B1(n3380), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3196) );
  AND2_X2 U4227 ( .A1(n3190), .A2(n3192), .ZN(n3371) );
  AND2_X2 U4228 ( .A1(n3189), .A2(n4524), .ZN(n3298) );
  AOI22_X1 U4229 ( .A1(n3371), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3195) );
  AND2_X2 U4230 ( .A1(n3190), .A2(n3189), .ZN(n3297) );
  AND2_X2 U4231 ( .A1(n3191), .A2(n4524), .ZN(n3271) );
  AOI22_X1 U4232 ( .A1(n3297), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4233 ( .A1(n3278), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4234 ( .A1(n3307), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3202) );
  AOI22_X1 U4235 ( .A1(n3370), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3201) );
  AOI22_X1 U4236 ( .A1(n3277), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3200) );
  AOI22_X1 U4237 ( .A1(n3305), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4238 ( .A1(n3371), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4239 ( .A1(n3299), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4240 ( .A1(n3297), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4241 ( .A1(n3307), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3213)
         );
  NAND2_X1 U4242 ( .A1(n3370), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3212)
         );
  NAND2_X1 U4243 ( .A1(n3305), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4244 ( .A1(n3380), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3210)
         );
  NAND2_X1 U4245 ( .A1(n3297), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4246 ( .A1(n3371), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3216)
         );
  NAND2_X1 U4247 ( .A1(n3298), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4248 ( .A1(n3295), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3214)
         );
  NAND2_X1 U4249 ( .A1(n3299), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4250 ( .A1(n3278), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U4251 ( .A1(n3272), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3219)
         );
  NAND2_X1 U4252 ( .A1(n3271), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4253 ( .A1(n3402), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4254 ( .A1(n3277), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3224) );
  NAND2_X1 U4255 ( .A1(n3306), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4256 ( .A1(n3270), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4257 ( .A1(n3307), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4258 ( .A1(n3371), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4259 ( .A1(n3370), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3230) );
  AOI22_X1 U4260 ( .A1(n3298), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3237) );
  AOI22_X1 U4261 ( .A1(n3297), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4262 ( .A1(n3288), .A2(n3321), .ZN(n3292) );
  NAND3_X1 U4263 ( .A1(n3317), .A2(n3351), .A3(n3292), .ZN(n4189) );
  NAND2_X1 U4264 ( .A1(n3380), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3243)
         );
  NAND2_X1 U4265 ( .A1(n3277), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4266 ( .A1(n4154), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4267 ( .A1(n3298), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4268 ( .A1(n3402), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3247) );
  NAND2_X1 U4269 ( .A1(n3305), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3246) );
  NAND2_X1 U4270 ( .A1(n3307), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3245)
         );
  NAND2_X1 U4271 ( .A1(n3270), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U4272 ( .A1(n3297), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3251) );
  NAND2_X1 U4273 ( .A1(n3371), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3250)
         );
  NAND2_X1 U4274 ( .A1(n3271), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3249) );
  NAND2_X1 U4275 ( .A1(n3295), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3248)
         );
  NAND2_X1 U4276 ( .A1(n3306), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3255) );
  NAND2_X1 U4277 ( .A1(n3370), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3254)
         );
  NAND2_X1 U4278 ( .A1(n3299), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3253) );
  NAND2_X1 U4279 ( .A1(n3272), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3252)
         );
  AOI22_X1 U4280 ( .A1(n3371), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3263) );
  AOI22_X1 U4281 ( .A1(n3278), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3261) );
  AOI22_X1 U4282 ( .A1(n3297), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4283 ( .A1(n3307), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4284 ( .A1(n3305), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3266) );
  AOI22_X1 U4285 ( .A1(n3277), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3265) );
  AOI22_X1 U4286 ( .A1(n3370), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3264) );
  NAND2_X2 U4287 ( .A1(n3269), .A2(n3268), .ZN(n3345) );
  NAND2_X1 U4288 ( .A1(n4189), .A2(n3343), .ZN(n3287) );
  AOI22_X1 U4289 ( .A1(n3370), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4290 ( .A1(n3297), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4291 ( .A1(n3371), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4292 ( .A1(n3305), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3282) );
  AOI22_X1 U4293 ( .A1(n3402), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3281) );
  AOI22_X1 U4294 ( .A1(n3298), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3278), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3280) );
  INV_X1 U4295 ( .A(n4230), .ZN(n3286) );
  NAND2_X1 U4296 ( .A1(n3286), .A2(n3285), .ZN(n4336) );
  XNOR2_X1 U4297 ( .A(n6593), .B(STATE_REG_1__SCAN_IN), .ZN(n4195) );
  INV_X1 U4298 ( .A(n3357), .ZN(n3290) );
  BUF_X1 U4299 ( .A(n3288), .Z(n3289) );
  NAND2_X1 U4300 ( .A1(n3290), .A2(n3289), .ZN(n3291) );
  NAND2_X1 U4301 ( .A1(n3346), .A2(n4496), .ZN(n4544) );
  AND2_X1 U4302 ( .A1(n3291), .A2(n4544), .ZN(n3314) );
  AND2_X2 U4303 ( .A1(n3337), .A2(n3320), .ZN(n3315) );
  NAND2_X1 U4304 ( .A1(n3315), .A2(n3317), .ZN(n3294) );
  AND2_X2 U4305 ( .A1(n3294), .A2(n3293), .ZN(n3350) );
  AOI22_X1 U4306 ( .A1(n4154), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4307 ( .A1(n3297), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3271), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4308 ( .A1(n3371), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3298), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4309 ( .A1(n3299), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3380), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3300) );
  NAND3_X1 U4310 ( .A1(n3302), .A2(n3301), .A3(n3300), .ZN(n3303) );
  AOI22_X1 U4311 ( .A1(n3370), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4312 ( .A1(n3305), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4313 ( .A1(n3307), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3402), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4314 ( .A1(n3277), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3272), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3308) );
  INV_X1 U4315 ( .A(n3315), .ZN(n3316) );
  NAND2_X1 U4316 ( .A1(n3316), .A2(n3313), .ZN(n3319) );
  INV_X1 U4317 ( .A(n3349), .ZN(n3318) );
  AND2_X1 U4318 ( .A1(n3320), .A2(n4456), .ZN(n3323) );
  NAND2_X1 U4319 ( .A1(n3285), .A2(n3342), .ZN(n3322) );
  NAND2_X2 U4320 ( .A1(n3325), .A2(n3324), .ZN(n3354) );
  OAI21_X1 U4321 ( .B1(n3346), .B2(n3333), .A(n3354), .ZN(n3326) );
  AOI21_X2 U4322 ( .B1(n3327), .B2(n3326), .A(n6576), .ZN(n3442) );
  NAND2_X1 U4323 ( .A1(n3442), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3332) );
  INV_X1 U4324 ( .A(n3674), .ZN(n3329) );
  INV_X1 U4325 ( .A(n6695), .ZN(n3328) );
  MUX2_X1 U4326 ( .A(n3329), .B(n3328), .S(n6372), .Z(n3330) );
  INV_X1 U4327 ( .A(n3330), .ZN(n3331) );
  NAND2_X1 U4328 ( .A1(n6541), .A2(n4457), .ZN(n4339) );
  NOR2_X1 U4329 ( .A1(n6670), .A2(n6576), .ZN(n6584) );
  INV_X1 U4330 ( .A(n4544), .ZN(n5115) );
  NAND2_X1 U4331 ( .A1(n3343), .A2(n4690), .ZN(n4191) );
  AND2_X1 U4332 ( .A1(n3344), .A2(n4191), .ZN(n3348) );
  NAND2_X1 U4333 ( .A1(n4752), .A2(n3346), .ZN(n3355) );
  NAND2_X1 U4334 ( .A1(n3354), .A2(n5092), .ZN(n3347) );
  NAND2_X1 U4335 ( .A1(n3122), .A2(n4333), .ZN(n3395) );
  NAND2_X1 U4336 ( .A1(n3397), .A2(n3395), .ZN(n3439) );
  INV_X1 U4337 ( .A(n3439), .ZN(n3364) );
  XNOR2_X1 U4338 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5279) );
  OAI22_X1 U4339 ( .A1(n6695), .A2(n5279), .B1(n3674), .B2(n5033), .ZN(n3361)
         );
  NAND3_X1 U4340 ( .A1(n5092), .A2(n3289), .A3(n4457), .ZN(n4334) );
  INV_X1 U4341 ( .A(n4334), .ZN(n3353) );
  NAND2_X1 U4342 ( .A1(n4456), .A2(n4697), .ZN(n4324) );
  INV_X1 U4343 ( .A(n3354), .ZN(n4192) );
  NOR2_X1 U4344 ( .A1(n3355), .A2(n4322), .ZN(n3356) );
  NAND2_X1 U4345 ( .A1(n4192), .A2(n3356), .ZN(n4212) );
  OAI211_X1 U4346 ( .C1(n4213), .C2(n3357), .A(n4221), .B(n4212), .ZN(n3358)
         );
  NAND2_X1 U4347 ( .A1(n3358), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3360) );
  INV_X1 U4348 ( .A(n3360), .ZN(n3362) );
  NAND2_X1 U4349 ( .A1(n3362), .A2(n3179), .ZN(n3438) );
  NAND2_X1 U4350 ( .A1(n3440), .A2(n3438), .ZN(n3363) );
  XNOR2_X1 U4351 ( .A(n3364), .B(n3363), .ZN(n4518) );
  NAND2_X1 U4352 ( .A1(n4518), .A2(n6576), .ZN(n3379) );
  AOI22_X1 U4353 ( .A1(n4142), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4354 ( .A1(n4099), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4355 ( .A1(n4114), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4356 ( .A1(n4115), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3366) );
  NAND4_X1 U4357 ( .A1(n3369), .A2(n3368), .A3(n3367), .A4(n3366), .ZN(n3377)
         );
  AOI22_X1 U4358 ( .A1(n3277), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4152), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3375) );
  AOI22_X1 U4359 ( .A1(n4073), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3374) );
  AOI22_X1 U4360 ( .A1(n4147), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3373) );
  AOI22_X1 U4361 ( .A1(n4145), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3372) );
  NAND4_X1 U4362 ( .A1(n3375), .A2(n3374), .A3(n3373), .A4(n3372), .ZN(n3376)
         );
  OR2_X1 U4363 ( .A1(n3590), .A2(n3391), .ZN(n3378) );
  NAND2_X2 U4364 ( .A1(n3379), .A2(n3378), .ZN(n3463) );
  NAND2_X1 U4365 ( .A1(n3665), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4366 ( .A1(n4142), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4367 ( .A1(n4073), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4368 ( .A1(n3371), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4369 ( .A1(n4114), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4370 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  AOI22_X1 U4371 ( .A1(n3277), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4372 ( .A1(n4147), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4373 ( .A1(n4152), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4374 ( .A1(n4154), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4375 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  OAI22_X1 U4376 ( .A1(n3590), .A2(n3594), .B1(n3490), .B2(n3391), .ZN(n3392)
         );
  INV_X1 U4377 ( .A(n3392), .ZN(n3393) );
  INV_X1 U4378 ( .A(n3395), .ZN(n3396) );
  XNOR2_X1 U4379 ( .A(n3397), .B(n3396), .ZN(n3689) );
  NAND2_X1 U4380 ( .A1(n3689), .A2(n6576), .ZN(n3411) );
  INV_X1 U4381 ( .A(n3590), .ZN(n3410) );
  AOI22_X1 U4382 ( .A1(n4073), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3307), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4383 ( .A1(n4152), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4384 ( .A1(n4099), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4385 ( .A1(n4154), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3398) );
  NAND4_X1 U4386 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3408)
         );
  AOI22_X1 U4387 ( .A1(n4094), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4388 ( .A1(n4144), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3405) );
  AOI22_X1 U4389 ( .A1(n4147), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3404) );
  AOI22_X1 U4390 ( .A1(n3371), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3403) );
  NAND4_X1 U4391 ( .A1(n3406), .A2(n3405), .A3(n3404), .A4(n3403), .ZN(n3407)
         );
  XNOR2_X1 U4392 ( .A(n3420), .B(n3594), .ZN(n3409) );
  NAND2_X1 U4393 ( .A1(n3410), .A2(n3409), .ZN(n3427) );
  NAND2_X1 U4394 ( .A1(n3665), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3415) );
  INV_X1 U4395 ( .A(n3594), .ZN(n3417) );
  NAND2_X1 U4396 ( .A1(n3346), .A2(n3469), .ZN(n3412) );
  OAI211_X1 U4397 ( .C1(n3417), .C2(n4220), .A(STATE2_REG_0__SCAN_IN), .B(
        n3412), .ZN(n3413) );
  INV_X1 U4398 ( .A(n3413), .ZN(n3414) );
  NAND2_X1 U4399 ( .A1(n3415), .A2(n3414), .ZN(n3426) );
  NAND2_X1 U4400 ( .A1(n3416), .A2(n3426), .ZN(n3430) );
  INV_X1 U4401 ( .A(n3465), .ZN(n3418) );
  NAND2_X1 U4402 ( .A1(n4637), .A2(n3636), .ZN(n3425) );
  XNOR2_X1 U4403 ( .A(n3420), .B(n3470), .ZN(n3423) );
  NAND2_X1 U4404 ( .A1(n3421), .A2(n3320), .ZN(n3422) );
  AOI21_X1 U4405 ( .B1(n4445), .B2(n3423), .A(n3422), .ZN(n3424) );
  INV_X1 U4406 ( .A(n3426), .ZN(n3428) );
  INV_X1 U4407 ( .A(n3636), .ZN(n3433) );
  INV_X1 U4408 ( .A(n4445), .ZN(n6700) );
  NAND2_X1 U4409 ( .A1(n3346), .A2(n3313), .ZN(n3472) );
  OAI21_X1 U4410 ( .B1(n6700), .B2(n3469), .A(n3472), .ZN(n3431) );
  INV_X1 U4411 ( .A(n3431), .ZN(n3432) );
  OAI21_X2 U4412 ( .B1(n3688), .B2(n3433), .A(n3432), .ZN(n4470) );
  NAND2_X1 U4413 ( .A1(n4470), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3434)
         );
  INV_X1 U4414 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4529) );
  NAND2_X1 U4415 ( .A1(n3434), .A2(n4529), .ZN(n3436) );
  AND2_X1 U4416 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4417 ( .A1(n4470), .A2(n3435), .ZN(n3437) );
  AND2_X1 U4418 ( .A1(n3436), .A2(n3437), .ZN(n4649) );
  NAND2_X1 U4420 ( .A1(n3485), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3447) );
  NAND2_X1 U4421 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3443) );
  NAND2_X1 U4422 ( .A1(n3443), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3444) );
  NOR2_X1 U4423 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n5033), .ZN(n4822)
         );
  NAND2_X1 U4424 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4822), .ZN(n6328) );
  OAI22_X1 U4425 ( .A1(n6695), .A2(n4935), .B1(n3674), .B2(n6762), .ZN(n3445)
         );
  INV_X1 U4426 ( .A(n3445), .ZN(n3446) );
  AOI22_X1 U4427 ( .A1(n4142), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4428 ( .A1(n4073), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4429 ( .A1(n4147), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4430 ( .A1(n4144), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4431 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  AOI22_X1 U4432 ( .A1(n4099), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4433 ( .A1(n4145), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4434 ( .A1(n4152), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4435 ( .A1(n4115), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4436 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  NOR2_X1 U4437 ( .A1(n3590), .A2(n3506), .ZN(n3458) );
  INV_X1 U4438 ( .A(n3665), .ZN(n3580) );
  INV_X1 U4439 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3459) );
  OAI22_X1 U4440 ( .A1(n3580), .A2(n3459), .B1(n3506), .B2(n3490), .ZN(n3460)
         );
  XNOR2_X1 U4441 ( .A(n3461), .B(n3460), .ZN(n3480) );
  OAI21_X1 U4442 ( .B1(n3465), .B2(n3464), .A(n3463), .ZN(n3467) );
  NAND2_X1 U4443 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  NAND2_X1 U4444 ( .A1(n3467), .A2(n3466), .ZN(n3481) );
  INV_X1 U4445 ( .A(n3481), .ZN(n3468) );
  XNOR2_X1 U4446 ( .A(n3480), .B(n3468), .ZN(n4643) );
  NAND2_X1 U4447 ( .A1(n3470), .A2(n3469), .ZN(n3507) );
  XNOR2_X1 U4448 ( .A(n3507), .B(n3471), .ZN(n3473) );
  OAI21_X1 U4449 ( .B1(n3473), .B2(n6700), .A(n3472), .ZN(n3474) );
  NAND2_X1 U4450 ( .A1(n3475), .A2(n6221), .ZN(n3479) );
  NAND2_X1 U4451 ( .A1(n3477), .A2(n3476), .ZN(n3478) );
  NAND2_X1 U4452 ( .A1(n3481), .A2(n3480), .ZN(n3504) );
  INV_X1 U4453 ( .A(n3504), .ZN(n3503) );
  INV_X1 U4454 ( .A(n3482), .ZN(n3484) );
  NAND2_X1 U4455 ( .A1(n3485), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3489) );
  NOR3_X1 U4456 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6762), .A3(n5033), 
        .ZN(n6416) );
  NAND2_X1 U4457 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6416), .ZN(n6406) );
  NAND2_X1 U4458 ( .A1(n6681), .A2(n6406), .ZN(n3486) );
  NOR3_X1 U4459 ( .A1(n6681), .A2(n6762), .A3(n5033), .ZN(n4932) );
  NAND2_X1 U4460 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4932), .ZN(n4862) );
  NAND2_X1 U4461 ( .A1(n3486), .A2(n4862), .ZN(n5037) );
  OAI22_X1 U4462 ( .A1(n6695), .A2(n5037), .B1(n3674), .B2(n6681), .ZN(n3487)
         );
  INV_X1 U4463 ( .A(n3487), .ZN(n3488) );
  AOI22_X1 U4464 ( .A1(n4142), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4465 ( .A1(n4073), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4466 ( .A1(n4147), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3492) );
  INV_X1 U4467 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6890) );
  AOI22_X1 U4468 ( .A1(n4144), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3491) );
  NAND4_X1 U4469 ( .A1(n3494), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3500)
         );
  AOI22_X1 U4470 ( .A1(n4099), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4471 ( .A1(n4145), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4472 ( .A1(n4152), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3496) );
  AOI22_X1 U4473 ( .A1(n4115), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3495) );
  NAND4_X1 U4474 ( .A1(n3498), .A2(n3497), .A3(n3496), .A4(n3495), .ZN(n3499)
         );
  AOI22_X1 U4475 ( .A1(n3665), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3670), 
        .B2(n3525), .ZN(n3501) );
  INV_X1 U4476 ( .A(n4989), .ZN(n4739) );
  NAND2_X2 U4477 ( .A1(n3503), .A2(n4739), .ZN(n3532) );
  NAND2_X1 U4478 ( .A1(n3504), .A2(n4989), .ZN(n3505) );
  NAND2_X1 U4479 ( .A1(n3507), .A2(n3506), .ZN(n3526) );
  INV_X1 U4480 ( .A(n3525), .ZN(n3508) );
  XNOR2_X1 U4481 ( .A(n3526), .B(n3508), .ZN(n3509) );
  NAND2_X1 U4482 ( .A1(n3509), .A2(n4445), .ZN(n3510) );
  INV_X1 U4483 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6808) );
  XNOR2_X1 U4484 ( .A(n3511), .B(n6808), .ZN(n4656) );
  NAND2_X1 U4485 ( .A1(n4655), .A2(n4656), .ZN(n4657) );
  NAND2_X1 U4486 ( .A1(n3511), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3512)
         );
  NAND2_X1 U4487 ( .A1(n4657), .A2(n3512), .ZN(n6208) );
  NAND2_X1 U4488 ( .A1(n3665), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4489 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4094), .B1(n4142), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3516) );
  AOI22_X1 U4490 ( .A1(n4073), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4491 ( .A1(n4147), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4492 ( .A1(n4144), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3513) );
  NAND4_X1 U4493 ( .A1(n3516), .A2(n3515), .A3(n3514), .A4(n3513), .ZN(n3522)
         );
  AOI22_X1 U4494 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n4099), .B1(n4114), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3520) );
  AOI22_X1 U4495 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4145), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3519) );
  AOI22_X1 U4496 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4152), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3518) );
  AOI22_X1 U4497 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4115), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3517) );
  NAND4_X1 U4498 ( .A1(n3520), .A2(n3519), .A3(n3518), .A4(n3517), .ZN(n3521)
         );
  NAND2_X1 U4499 ( .A1(n3670), .A2(n3547), .ZN(n3523) );
  NAND2_X1 U4500 ( .A1(n3524), .A2(n3523), .ZN(n3533) );
  XNOR2_X1 U4501 ( .A(n3532), .B(n3533), .ZN(n3717) );
  NAND2_X1 U4502 ( .A1(n3717), .A2(n3636), .ZN(n3529) );
  NAND2_X1 U4503 ( .A1(n3526), .A2(n3525), .ZN(n3549) );
  XNOR2_X1 U4504 ( .A(n3549), .B(n3547), .ZN(n3527) );
  NAND2_X1 U4505 ( .A1(n3527), .A2(n4445), .ZN(n3528) );
  NAND2_X1 U4506 ( .A1(n3529), .A2(n3528), .ZN(n3530) );
  INV_X1 U4507 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6979) );
  XNOR2_X1 U4508 ( .A(n3530), .B(n6979), .ZN(n6207) );
  NAND2_X1 U4509 ( .A1(n6208), .A2(n6207), .ZN(n6210) );
  NAND2_X1 U4510 ( .A1(n3530), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3531)
         );
  NAND2_X1 U4511 ( .A1(n3665), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3546) );
  AOI22_X1 U4512 ( .A1(n4145), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4513 ( .A1(n4073), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4514 ( .A1(n4094), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3536) );
  AOI22_X1 U4515 ( .A1(n4144), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4516 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AOI22_X1 U4517 ( .A1(n4152), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4518 ( .A1(n4147), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3541) );
  INV_X1 U4519 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6885) );
  AOI22_X1 U4520 ( .A1(n4117), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4521 ( .A1(n4114), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4522 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  NAND2_X1 U4523 ( .A1(n3670), .A2(n3571), .ZN(n3545) );
  NAND2_X1 U4524 ( .A1(n3546), .A2(n3545), .ZN(n3556) );
  NAND2_X1 U4525 ( .A1(n3718), .A2(n3636), .ZN(n3552) );
  INV_X1 U4526 ( .A(n3547), .ZN(n3548) );
  OR2_X1 U4527 ( .A1(n3549), .A2(n3548), .ZN(n3570) );
  XNOR2_X1 U4528 ( .A(n3570), .B(n3571), .ZN(n3550) );
  NAND2_X1 U4529 ( .A1(n3550), .A2(n4445), .ZN(n3551) );
  NAND2_X1 U4530 ( .A1(n3552), .A2(n3551), .ZN(n3553) );
  INV_X1 U4531 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6275) );
  XNOR2_X1 U4532 ( .A(n3553), .B(n6275), .ZN(n4733) );
  NAND2_X1 U4533 ( .A1(n3553), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3554)
         );
  NAND2_X1 U4534 ( .A1(n4732), .A2(n3554), .ZN(n4813) );
  NAND2_X1 U4535 ( .A1(n3557), .A2(n3556), .ZN(n3569) );
  AOI22_X1 U4536 ( .A1(n4142), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4537 ( .A1(n4073), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4538 ( .A1(n4147), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3559) );
  AOI22_X1 U4539 ( .A1(n4144), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3558) );
  NAND4_X1 U4540 ( .A1(n3561), .A2(n3560), .A3(n3559), .A4(n3558), .ZN(n3567)
         );
  AOI22_X1 U4541 ( .A1(n4099), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4542 ( .A1(n4145), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4543 ( .A1(n4152), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4544 ( .A1(n4115), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4545 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3566)
         );
  AOI22_X1 U4546 ( .A1(n3665), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3670), 
        .B2(n3583), .ZN(n3568) );
  OR2_X2 U4547 ( .A1(n3569), .A2(n3568), .ZN(n3593) );
  NAND2_X1 U4548 ( .A1(n3569), .A2(n3568), .ZN(n3727) );
  NAND3_X1 U4549 ( .A1(n3593), .A2(n3727), .A3(n3636), .ZN(n3575) );
  INV_X1 U4550 ( .A(n3570), .ZN(n3572) );
  NAND2_X1 U4551 ( .A1(n3572), .A2(n3571), .ZN(n3582) );
  XNOR2_X1 U4552 ( .A(n3582), .B(n3583), .ZN(n3573) );
  NAND2_X1 U4553 ( .A1(n3573), .A2(n4445), .ZN(n3574) );
  NAND2_X1 U4554 ( .A1(n3575), .A2(n3574), .ZN(n3576) );
  INV_X1 U4555 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4249) );
  XNOR2_X1 U4556 ( .A(n3576), .B(n4249), .ZN(n4812) );
  NAND2_X1 U4557 ( .A1(n3576), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3577)
         );
  NAND2_X1 U4558 ( .A1(n4811), .A2(n3577), .ZN(n4977) );
  INV_X1 U4559 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3579) );
  NAND2_X1 U4560 ( .A1(n3670), .A2(n3594), .ZN(n3578) );
  OAI21_X1 U4561 ( .B1(n3580), .B2(n3579), .A(n3578), .ZN(n3581) );
  NAND2_X1 U4562 ( .A1(n3732), .A2(n3636), .ZN(n3587) );
  INV_X1 U4563 ( .A(n3582), .ZN(n3584) );
  NAND2_X1 U4564 ( .A1(n3584), .A2(n3583), .ZN(n3596) );
  XNOR2_X1 U4565 ( .A(n3596), .B(n3594), .ZN(n3585) );
  NAND2_X1 U4566 ( .A1(n3585), .A2(n4445), .ZN(n3586) );
  NAND2_X1 U4567 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  INV_X1 U4568 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6273) );
  XNOR2_X1 U4569 ( .A(n3588), .B(n6273), .ZN(n4976) );
  NAND2_X1 U4570 ( .A1(n3588), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3589)
         );
  NAND2_X1 U4571 ( .A1(n3636), .A2(n3594), .ZN(n3591) );
  NOR2_X1 U4572 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  NAND2_X1 U4573 ( .A1(n4445), .A2(n3594), .ZN(n3595) );
  OR2_X1 U4574 ( .A1(n3596), .A2(n3595), .ZN(n3597) );
  NAND2_X1 U4575 ( .A1(n3602), .A2(n3597), .ZN(n3598) );
  INV_X1 U4576 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4256) );
  XNOR2_X1 U4577 ( .A(n3598), .B(n4256), .ZN(n5176) );
  NAND2_X1 U4578 ( .A1(n3598), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3599)
         );
  INV_X1 U4579 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U4580 ( .A1(n3602), .A2(n6255), .ZN(n5245) );
  OR2_X1 U4581 ( .A1(n3602), .A2(n6255), .ZN(n5246) );
  NAND2_X1 U4582 ( .A1(n3601), .A2(n3600), .ZN(n5340) );
  NAND3_X1 U4583 ( .A1(n5318), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4584 ( .A1(n3605), .A2(n3604), .ZN(n5348) );
  INV_X1 U4585 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6927) );
  NOR2_X1 U4586 ( .A1(n5582), .A2(n6927), .ZN(n5349) );
  NAND2_X1 U4587 ( .A1(n5582), .A2(n6927), .ZN(n5350) );
  INV_X4 U4588 ( .A(n5554), .ZN(n5582) );
  XNOR2_X1 U4589 ( .A(n5582), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5590)
         );
  INV_X1 U4590 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6949) );
  INV_X1 U4591 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3606) );
  AND2_X1 U4592 ( .A1(n5582), .A2(n3606), .ZN(n3607) );
  INV_X1 U4593 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6993) );
  NOR2_X1 U4594 ( .A1(n5582), .A2(n6993), .ZN(n3609) );
  NAND2_X1 U4595 ( .A1(n5582), .A2(n6993), .ZN(n3608) );
  OAI21_X1 U4596 ( .B1(n5575), .B2(n3609), .A(n3608), .ZN(n5555) );
  INV_X1 U4597 ( .A(n5555), .ZN(n3611) );
  AND2_X1 U4598 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U4599 ( .A1(n4359), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3610) );
  NAND2_X1 U4600 ( .A1(n3611), .A2(n3127), .ZN(n5529) );
  INV_X1 U4601 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5731) );
  INV_X1 U4602 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5966) );
  INV_X1 U4603 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5716) );
  NAND3_X1 U4604 ( .A1(n5731), .A2(n5966), .A3(n5716), .ZN(n3612) );
  NAND2_X1 U4605 ( .A1(n5554), .A2(n3612), .ZN(n3613) );
  AND2_X1 U4606 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5688) );
  AND2_X1 U4607 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3614) );
  NAND2_X1 U4608 ( .A1(n5688), .A2(n3614), .ZN(n4346) );
  NAND2_X1 U4609 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5600) );
  OAI21_X1 U4610 ( .B1(n4346), .B2(n5600), .A(n5582), .ZN(n3615) );
  NOR2_X1 U4611 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4363) );
  NOR2_X1 U4612 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5687) );
  INV_X1 U4613 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n6774) );
  INV_X1 U4614 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4308) );
  NAND4_X1 U4615 ( .A1(n4363), .A2(n5687), .A3(n6774), .A4(n4308), .ZN(n3616)
         );
  NAND2_X1 U4616 ( .A1(n5554), .A2(n3616), .ZN(n3617) );
  INV_X1 U4617 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U4618 ( .A1(n3602), .A2(n6788), .ZN(n3618) );
  NAND2_X1 U4619 ( .A1(n3621), .A2(n3618), .ZN(n4381) );
  INV_X1 U4620 ( .A(n4381), .ZN(n3620) );
  INV_X1 U4621 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U4622 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5602) );
  INV_X1 U4623 ( .A(n3621), .ZN(n3623) );
  INV_X1 U4624 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6843) );
  INV_X1 U4625 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5505) );
  NAND3_X1 U4626 ( .A1(n6843), .A2(n5520), .A3(n5505), .ZN(n3622) );
  NOR2_X1 U4627 ( .A1(n5582), .A2(n3622), .ZN(n4382) );
  INV_X1 U4628 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5614) );
  INV_X1 U4629 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5624) );
  NAND4_X1 U4630 ( .A1(n3623), .A2(n4382), .A3(n5614), .A4(n5624), .ZN(n3624)
         );
  XNOR2_X1 U4631 ( .A(n3625), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5613)
         );
  NAND2_X1 U4632 ( .A1(n3180), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3626) );
  NAND2_X1 U4633 ( .A1(n3627), .A2(n3626), .ZN(n3637) );
  NAND2_X1 U4634 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6372), .ZN(n3641) );
  NAND2_X1 U4635 ( .A1(n5388), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3628) );
  NOR2_X1 U4636 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6554), .ZN(n3631)
         );
  NOR2_X1 U4637 ( .A1(n3633), .A2(n3632), .ZN(n3634) );
  OR2_X1 U4638 ( .A1(n3635), .A2(n3634), .ZN(n4198) );
  OAI21_X1 U4639 ( .B1(n3658), .B2(n4752), .A(n3320), .ZN(n3652) );
  INV_X1 U4640 ( .A(n3637), .ZN(n3640) );
  INV_X1 U4641 ( .A(n3641), .ZN(n3639) );
  OAI21_X1 U4642 ( .B1(n3640), .B2(n3639), .A(n3638), .ZN(n4199) );
  NOR2_X1 U4643 ( .A1(n4199), .A2(n6576), .ZN(n3651) );
  OAI21_X1 U4644 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6372), .A(n3641), 
        .ZN(n3642) );
  INV_X1 U4645 ( .A(n3642), .ZN(n3649) );
  AOI21_X1 U4646 ( .B1(n3649), .B2(n4322), .A(n3643), .ZN(n3644) );
  OAI21_X1 U4647 ( .B1(n3289), .B2(n4496), .A(n3355), .ZN(n3656) );
  OAI22_X1 U4648 ( .A1(n3652), .A2(n3651), .B1(n3644), .B2(n3656), .ZN(n3645)
         );
  INV_X1 U4649 ( .A(n3645), .ZN(n3650) );
  XNOR2_X1 U4650 ( .A(n3647), .B(n3646), .ZN(n4200) );
  INV_X1 U4651 ( .A(n4200), .ZN(n3648) );
  AOI22_X1 U4652 ( .A1(n3650), .A2(n3649), .B1(n3656), .B2(n3648), .ZN(n3655)
         );
  OAI21_X1 U4653 ( .B1(n3650), .B2(n4199), .A(n3671), .ZN(n3654) );
  NAND2_X1 U4654 ( .A1(n3652), .A2(n3651), .ZN(n3653) );
  OAI211_X1 U4655 ( .C1(n3655), .C2(n3658), .A(n3654), .B(n3653), .ZN(n3660)
         );
  AOI21_X1 U4656 ( .B1(n3665), .B2(n4200), .A(n3656), .ZN(n3657) );
  OAI21_X1 U4657 ( .B1(n3658), .B2(n4200), .A(n3657), .ZN(n3659) );
  OAI211_X1 U4658 ( .C1(n3665), .C2(n3662), .A(n3660), .B(n3659), .ZN(n3661)
         );
  OAI21_X1 U4659 ( .B1(n3662), .B2(n3666), .A(n3661), .ZN(n3663) );
  AOI21_X1 U4660 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6576), .A(n3663), 
        .ZN(n3668) );
  NAND3_X1 U4661 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3664), .A3(n6802), .ZN(n4196) );
  NOR2_X1 U4662 ( .A1(n3665), .A2(n4196), .ZN(n3667) );
  NOR2_X1 U4663 ( .A1(n4532), .A2(n4322), .ZN(n6557) );
  INV_X1 U4664 ( .A(n3676), .ZN(n3682) );
  AOI21_X1 U4665 ( .B1(n3699), .B2(n4653), .A(n3713), .ZN(n6088) );
  NAND2_X1 U4666 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4667 ( .A1(n6334), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3870) );
  NOR2_X1 U4668 ( .A1(n3870), .A2(n4653), .ZN(n3678) );
  AOI21_X1 U4669 ( .B1(n4167), .B2(EAX_REG_3__SCAN_IN), .A(n3678), .ZN(n3679)
         );
  OAI211_X1 U4670 ( .C1(n6088), .C2(n3711), .A(n3680), .B(n3679), .ZN(n3681)
         );
  AOI21_X1 U4671 ( .B1(n3682), .B2(n3677), .A(n3681), .ZN(n4625) );
  INV_X1 U4672 ( .A(n4625), .ZN(n3706) );
  NAND2_X1 U4673 ( .A1(n4643), .A2(n3677), .ZN(n3683) );
  NAND2_X1 U4674 ( .A1(n4637), .A2(n3677), .ZN(n3687) );
  AOI22_X1 U4675 ( .A1(n4167), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6334), .ZN(n3685) );
  NAND2_X1 U4676 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3684) );
  AND2_X1 U4677 ( .A1(n3685), .A2(n3684), .ZN(n3686) );
  NAND2_X1 U4678 ( .A1(n5043), .A2(n4335), .ZN(n4481) );
  NAND2_X1 U4679 ( .A1(n3690), .A2(n3677), .ZN(n3695) );
  AOI22_X1 U4680 ( .A1(n3691), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6334), .ZN(n3693) );
  NAND2_X1 U4681 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3692) );
  AND2_X1 U4682 ( .A1(n3693), .A2(n3692), .ZN(n3694) );
  NAND2_X1 U4683 ( .A1(n3695), .A2(n3694), .ZN(n3697) );
  AND2_X1 U4684 ( .A1(n3697), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3696) );
  NAND2_X1 U4685 ( .A1(n4481), .A2(n3696), .ZN(n4484) );
  INV_X1 U4686 ( .A(n3697), .ZN(n4482) );
  NAND2_X1 U4687 ( .A1(n4482), .A2(n4165), .ZN(n3698) );
  NAND2_X1 U4688 ( .A1(n4484), .A2(n3698), .ZN(n4462) );
  NAND2_X1 U4689 ( .A1(n4694), .A2(n4461), .ZN(n3705) );
  NAND2_X1 U4690 ( .A1(n3707), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3704) );
  OAI21_X1 U4691 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3699), .ZN(n6227) );
  NAND2_X1 U4692 ( .A1(n6227), .A2(n4165), .ZN(n3701) );
  NAND2_X1 U4693 ( .A1(n4170), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3700)
         );
  NAND2_X1 U4694 ( .A1(n3701), .A2(n3700), .ZN(n3702) );
  AOI21_X1 U4695 ( .B1(n4167), .B2(EAX_REG_2__SCAN_IN), .A(n3702), .ZN(n3703)
         );
  AND2_X1 U4696 ( .A1(n3704), .A2(n3703), .ZN(n4692) );
  INV_X1 U4697 ( .A(n3707), .ZN(n3710) );
  NAND2_X1 U4698 ( .A1(n6334), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3709)
         );
  NAND2_X1 U4699 ( .A1(n4167), .A2(EAX_REG_4__SCAN_IN), .ZN(n3708) );
  OAI211_X1 U4700 ( .C1(n3710), .C2(n6802), .A(n3709), .B(n3708), .ZN(n3712)
         );
  NAND2_X1 U4701 ( .A1(n3712), .A2(n3711), .ZN(n3715) );
  OAI21_X1 U4702 ( .B1(n3713), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3721), 
        .ZN(n6217) );
  NAND2_X1 U4703 ( .A1(n6217), .A2(n4165), .ZN(n3714) );
  NAND2_X1 U4704 ( .A1(n3715), .A2(n3714), .ZN(n3716) );
  AOI21_X1 U4705 ( .B1(n3717), .B2(n3677), .A(n3716), .ZN(n4630) );
  XOR2_X1 U4706 ( .A(n5098), .B(n3721), .Z(n5095) );
  NAND2_X1 U4707 ( .A1(n3718), .A2(n3677), .ZN(n3720) );
  AOI22_X1 U4708 ( .A1(n3691), .A2(EAX_REG_5__SCAN_IN), .B1(n4170), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3719) );
  OAI211_X1 U4709 ( .C1(n5095), .C2(n3711), .A(n3720), .B(n3719), .ZN(n4682)
         );
  OAI21_X1 U4710 ( .B1(n3722), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3729), 
        .ZN(n6206) );
  INV_X1 U4711 ( .A(n6206), .ZN(n3725) );
  NAND2_X1 U4712 ( .A1(n3691), .A2(EAX_REG_6__SCAN_IN), .ZN(n3724) );
  INV_X1 U4713 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5991) );
  OAI21_X1 U4714 ( .B1(n5991), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6334), 
        .ZN(n3723) );
  AOI22_X1 U4715 ( .A1(n4165), .A2(n3725), .B1(n3724), .B2(n3723), .ZN(n3726)
         );
  NAND2_X1 U4716 ( .A1(n3109), .A2(n4629), .ZN(n4728) );
  AOI21_X1 U4717 ( .B1(n6778), .B2(n3729), .A(n3747), .ZN(n5078) );
  AOI22_X1 U4718 ( .A1(n3691), .A2(EAX_REG_7__SCAN_IN), .B1(n4170), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3730) );
  OAI21_X1 U4719 ( .B1(n5078), .B2(n3711), .A(n3730), .ZN(n3731) );
  AOI21_X1 U4720 ( .B1(n3732), .B2(n3677), .A(n3731), .ZN(n4729) );
  AOI22_X1 U4721 ( .A1(n4147), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4722 ( .A1(n4073), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4723 ( .A1(n4152), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4724 ( .A1(n4145), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3733) );
  NAND4_X1 U4725 ( .A1(n3736), .A2(n3735), .A3(n3734), .A4(n3733), .ZN(n3742)
         );
  AOI22_X1 U4726 ( .A1(n4144), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3740) );
  AOI22_X1 U4727 ( .A1(n4094), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4728 ( .A1(n4115), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4729 ( .A1(n4116), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3737) );
  NAND4_X1 U4730 ( .A1(n3740), .A2(n3739), .A3(n3738), .A4(n3737), .ZN(n3741)
         );
  NOR2_X1 U4731 ( .A1(n3742), .A2(n3741), .ZN(n3746) );
  INV_X1 U4732 ( .A(n3677), .ZN(n3745) );
  XNOR2_X1 U4733 ( .A(n3747), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5179) );
  NAND2_X1 U4734 ( .A1(n5179), .A2(n4165), .ZN(n3744) );
  AOI22_X1 U4735 ( .A1(n3691), .A2(EAX_REG_8__SCAN_IN), .B1(n4170), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3743) );
  OAI211_X1 U4736 ( .C1(n3746), .C2(n3745), .A(n3744), .B(n3743), .ZN(n4773)
         );
  XOR2_X1 U4737 ( .A(n6051), .B(n3763), .Z(n6056) );
  INV_X1 U4738 ( .A(n6056), .ZN(n5250) );
  AOI22_X1 U4739 ( .A1(n4142), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4740 ( .A1(n4073), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4741 ( .A1(n4147), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4742 ( .A1(n4116), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4743 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3757)
         );
  AOI22_X1 U4744 ( .A1(n4144), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4745 ( .A1(n4152), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4746 ( .A1(n4145), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4747 ( .A1(n4099), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3752) );
  NAND4_X1 U4748 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3756)
         );
  OAI21_X1 U4749 ( .B1(n3757), .B2(n3756), .A(n3677), .ZN(n3760) );
  NAND2_X1 U4750 ( .A1(n3691), .A2(EAX_REG_9__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4751 ( .A1(n4170), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3758)
         );
  NAND3_X1 U4752 ( .A1(n3760), .A2(n3759), .A3(n3758), .ZN(n3761) );
  AOI21_X1 U4753 ( .B1(n5250), .B2(n4165), .A(n3761), .ZN(n4982) );
  XNOR2_X1 U4754 ( .A(n3780), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6043)
         );
  AOI22_X1 U4755 ( .A1(n4073), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4756 ( .A1(n4099), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4757 ( .A1(n4117), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4758 ( .A1(n4144), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4759 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3773)
         );
  AOI22_X1 U4760 ( .A1(n4142), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4761 ( .A1(n4152), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3770) );
  AOI22_X1 U4762 ( .A1(n4145), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3769) );
  AOI22_X1 U4763 ( .A1(n4147), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3768) );
  NAND4_X1 U4764 ( .A1(n3771), .A2(n3770), .A3(n3769), .A4(n3768), .ZN(n3772)
         );
  OAI21_X1 U4765 ( .B1(n3773), .B2(n3772), .A(n3677), .ZN(n3776) );
  NAND2_X1 U4766 ( .A1(n3691), .A2(EAX_REG_10__SCAN_IN), .ZN(n3775) );
  NAND2_X1 U4767 ( .A1(n4170), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3774)
         );
  NAND3_X1 U4768 ( .A1(n3776), .A2(n3775), .A3(n3774), .ZN(n3777) );
  AOI21_X1 U4769 ( .B1(n6043), .B2(n4165), .A(n3777), .ZN(n5085) );
  NAND2_X1 U4770 ( .A1(n3779), .A2(n3778), .ZN(n5084) );
  XOR2_X1 U4771 ( .A(n6032), .B(n3796), .Z(n6195) );
  INV_X1 U4772 ( .A(n6195), .ZN(n3795) );
  AOI22_X1 U4773 ( .A1(n4147), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3784) );
  AOI22_X1 U4774 ( .A1(n4073), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3783) );
  AOI22_X1 U4775 ( .A1(n4152), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3782) );
  AOI22_X1 U4776 ( .A1(n4115), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3781) );
  NAND4_X1 U4777 ( .A1(n3784), .A2(n3783), .A3(n3782), .A4(n3781), .ZN(n3790)
         );
  AOI22_X1 U4778 ( .A1(n4145), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3788) );
  AOI22_X1 U4779 ( .A1(n4094), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3787) );
  AOI22_X1 U4780 ( .A1(n4099), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3786) );
  AOI22_X1 U4781 ( .A1(n4144), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3785) );
  NAND4_X1 U4782 ( .A1(n3788), .A2(n3787), .A3(n3786), .A4(n3785), .ZN(n3789)
         );
  OAI21_X1 U4783 ( .B1(n3790), .B2(n3789), .A(n3677), .ZN(n3793) );
  NAND2_X1 U4784 ( .A1(n3691), .A2(EAX_REG_11__SCAN_IN), .ZN(n3792) );
  NAND2_X1 U4785 ( .A1(n4170), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3791)
         );
  NAND3_X1 U4786 ( .A1(n3793), .A2(n3792), .A3(n3791), .ZN(n3794) );
  AOI21_X1 U4787 ( .B1(n3795), .B2(n4165), .A(n3794), .ZN(n5173) );
  XNOR2_X1 U4788 ( .A(n3811), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5355)
         );
  INV_X1 U4789 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5261) );
  AOI21_X1 U4790 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5261), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3798) );
  AND2_X1 U4791 ( .A1(n4167), .A2(EAX_REG_12__SCAN_IN), .ZN(n3797) );
  OAI22_X1 U4792 ( .A1(n5355), .A2(n3711), .B1(n3798), .B2(n3797), .ZN(n3810)
         );
  AOI22_X1 U4793 ( .A1(n4073), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4794 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4099), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4795 ( .A1(n4145), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4796 ( .A1(n4094), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4797 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3808)
         );
  AOI22_X1 U4798 ( .A1(n4147), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4799 ( .A1(n4152), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4800 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4117), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4801 ( .A1(n4144), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4802 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3807)
         );
  OAI21_X1 U4803 ( .B1(n3808), .B2(n3807), .A(n3677), .ZN(n3809) );
  NAND2_X1 U4804 ( .A1(n3810), .A2(n3809), .ZN(n5234) );
  XOR2_X1 U4805 ( .A(n5272), .B(n3825), .Z(n5593) );
  AOI22_X1 U4806 ( .A1(n4147), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3815) );
  AOI22_X1 U4807 ( .A1(n4099), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4808 ( .A1(n4145), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4809 ( .A1(n4143), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3812) );
  NAND4_X1 U4810 ( .A1(n3815), .A2(n3814), .A3(n3813), .A4(n3812), .ZN(n3821)
         );
  AOI22_X1 U4811 ( .A1(n4073), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4812 ( .A1(n4152), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4813 ( .A1(n4142), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4814 ( .A1(n4116), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3816) );
  NAND4_X1 U4815 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3820)
         );
  OR2_X1 U4816 ( .A1(n3821), .A2(n3820), .ZN(n3822) );
  AOI22_X1 U4817 ( .A1(n3677), .A2(n3822), .B1(n4170), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4818 ( .A1(n3691), .A2(EAX_REG_13__SCAN_IN), .ZN(n3823) );
  OAI211_X1 U4819 ( .C1(n5593), .C2(n3711), .A(n3824), .B(n3823), .ZN(n5255)
         );
  XNOR2_X1 U4820 ( .A(n3841), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5585)
         );
  AOI22_X1 U4821 ( .A1(n4147), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4822 ( .A1(n4144), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4823 ( .A1(n4117), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4824 ( .A1(n4152), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4825 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3835)
         );
  AOI22_X1 U4826 ( .A1(n4073), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4827 ( .A1(n4094), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4828 ( .A1(n4099), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4829 ( .A1(n4145), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4830 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  OAI21_X1 U4831 ( .B1(n3835), .B2(n3834), .A(n3677), .ZN(n3838) );
  NAND2_X1 U4832 ( .A1(n3691), .A2(EAX_REG_14__SCAN_IN), .ZN(n3837) );
  NAND2_X1 U4833 ( .A1(n4170), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3836)
         );
  NAND3_X1 U4834 ( .A1(n3838), .A2(n3837), .A3(n3836), .ZN(n3839) );
  AOI21_X1 U4835 ( .B1(n5585), .B2(n4165), .A(n3839), .ZN(n5326) );
  XOR2_X1 U4836 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3859), .Z(n6026) );
  INV_X1 U4837 ( .A(n6026), .ZN(n3856) );
  AOI22_X1 U4838 ( .A1(n4147), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4839 ( .A1(n4073), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4840 ( .A1(n4144), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4841 ( .A1(n4152), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4842 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3851)
         );
  AOI22_X1 U4843 ( .A1(n4143), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4844 ( .A1(n4117), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4845 ( .A1(n4145), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4846 ( .A1(n4099), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4847 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  OAI21_X1 U4848 ( .B1(n3851), .B2(n3850), .A(n3677), .ZN(n3854) );
  NAND2_X1 U4849 ( .A1(n4167), .A2(EAX_REG_15__SCAN_IN), .ZN(n3853) );
  NAND2_X1 U4850 ( .A1(n4170), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3852)
         );
  NAND3_X1 U4851 ( .A1(n3854), .A2(n3853), .A3(n3852), .ZN(n3855) );
  AOI21_X1 U4852 ( .B1(n3856), .B2(n4165), .A(n3855), .ZN(n5362) );
  NAND2_X1 U4853 ( .A1(n3858), .A2(n3857), .ZN(n5360) );
  XNOR2_X1 U4854 ( .A(n3889), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5571)
         );
  INV_X1 U4855 ( .A(n5571), .ZN(n3875) );
  AOI22_X1 U4856 ( .A1(n4073), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4147), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4857 ( .A1(n4099), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4858 ( .A1(n4145), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4859 ( .A1(n4117), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3860) );
  NAND4_X1 U4860 ( .A1(n3863), .A2(n3862), .A3(n3861), .A4(n3860), .ZN(n3869)
         );
  AOI22_X1 U4861 ( .A1(n4142), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4862 ( .A1(n4094), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4863 ( .A1(n4152), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4864 ( .A1(n4144), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3864) );
  NAND4_X1 U4865 ( .A1(n3867), .A2(n3866), .A3(n3865), .A4(n3864), .ZN(n3868)
         );
  NOR2_X1 U4866 ( .A1(n3869), .A2(n3868), .ZN(n3873) );
  NOR2_X1 U4867 ( .A1(n3870), .A2(n5569), .ZN(n3871) );
  AOI21_X1 U4868 ( .B1(n4167), .B2(EAX_REG_16__SCAN_IN), .A(n3871), .ZN(n3872)
         );
  OAI21_X1 U4869 ( .B1(n4133), .B2(n3873), .A(n3872), .ZN(n3874) );
  AOI21_X1 U4870 ( .B1(n3875), .B2(n4165), .A(n3874), .ZN(n5368) );
  NOR2_X2 U4871 ( .A1(n5360), .A2(n5368), .ZN(n5366) );
  AOI22_X1 U4872 ( .A1(n4142), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4873 ( .A1(n4073), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4874 ( .A1(n4099), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4875 ( .A1(n4147), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4876 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  AOI22_X1 U4877 ( .A1(n4152), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4878 ( .A1(n4117), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4879 ( .A1(n4145), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4880 ( .A1(n4094), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4881 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NOR2_X1 U4882 ( .A1(n3885), .A2(n3884), .ZN(n3886) );
  OR2_X1 U4883 ( .A1(n4133), .A2(n3886), .ZN(n3893) );
  NAND2_X1 U4884 ( .A1(n6334), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3887)
         );
  NAND2_X1 U4885 ( .A1(n3711), .A2(n3887), .ZN(n3888) );
  AOI21_X1 U4886 ( .B1(n4167), .B2(EAX_REG_17__SCAN_IN), .A(n3888), .ZN(n3892)
         );
  OAI21_X1 U4887 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3890), .A(n3924), 
        .ZN(n6015) );
  NOR2_X1 U4888 ( .A1(n6015), .A2(n3711), .ZN(n3891) );
  AOI21_X1 U4889 ( .B1(n3893), .B2(n3892), .A(n3891), .ZN(n5949) );
  AOI22_X1 U4890 ( .A1(n4142), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4891 ( .A1(n4145), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3896) );
  AOI22_X1 U4892 ( .A1(n4143), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4893 ( .A1(n4152), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3894) );
  NAND4_X1 U4894 ( .A1(n3897), .A2(n3896), .A3(n3895), .A4(n3894), .ZN(n3903)
         );
  AOI22_X1 U4895 ( .A1(n4073), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4896 ( .A1(n4099), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4897 ( .A1(n4147), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4898 ( .A1(n4117), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3898) );
  NAND4_X1 U4899 ( .A1(n3901), .A2(n3900), .A3(n3899), .A4(n3898), .ZN(n3902)
         );
  NOR2_X1 U4900 ( .A1(n3903), .A2(n3902), .ZN(n3906) );
  OAI21_X1 U4901 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5559), .A(n3711), .ZN(
        n3904) );
  AOI21_X1 U4902 ( .B1(n4167), .B2(EAX_REG_18__SCAN_IN), .A(n3904), .ZN(n3905)
         );
  OAI21_X1 U4903 ( .B1(n4133), .B2(n3906), .A(n3905), .ZN(n3908) );
  XNOR2_X1 U4904 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3924), .ZN(n6007)
         );
  NAND2_X1 U4905 ( .A1(n6007), .A2(n4165), .ZN(n3907) );
  NAND2_X1 U4906 ( .A1(n3908), .A2(n3907), .ZN(n5562) );
  AOI22_X1 U4907 ( .A1(n4147), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4908 ( .A1(n4073), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4909 ( .A1(n4152), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4910 ( .A1(n4099), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4911 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4912 ( .A1(n4094), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4913 ( .A1(n4117), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4914 ( .A1(n4115), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4915 ( .A1(n4143), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4916 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  NOR2_X1 U4917 ( .A1(n3919), .A2(n3918), .ZN(n3923) );
  OAI21_X1 U4918 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5991), .A(n6334), 
        .ZN(n3920) );
  INV_X1 U4919 ( .A(n3920), .ZN(n3921) );
  AOI21_X1 U4920 ( .B1(n4167), .B2(EAX_REG_19__SCAN_IN), .A(n3921), .ZN(n3922)
         );
  OAI21_X1 U4921 ( .B1(n4133), .B2(n3923), .A(n3922), .ZN(n3927) );
  OAI21_X1 U4922 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3925), .A(n3958), 
        .ZN(n5942) );
  OR2_X1 U4923 ( .A1(n3711), .A2(n5942), .ZN(n3926) );
  NAND2_X1 U4924 ( .A1(n3927), .A2(n3926), .ZN(n5897) );
  AOI22_X1 U4925 ( .A1(n4073), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4926 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n4114), .B1(n4099), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4927 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4145), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4928 ( .A1(n4147), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3928) );
  NAND4_X1 U4929 ( .A1(n3931), .A2(n3930), .A3(n3929), .A4(n3928), .ZN(n3937)
         );
  AOI22_X1 U4930 ( .A1(n4142), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4931 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4152), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4932 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4115), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4933 ( .A1(n4144), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3932) );
  NAND4_X1 U4934 ( .A1(n3935), .A2(n3934), .A3(n3933), .A4(n3932), .ZN(n3936)
         );
  NOR2_X1 U4935 ( .A1(n3937), .A2(n3936), .ZN(n3941) );
  NAND2_X1 U4936 ( .A1(n6334), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3938)
         );
  NAND2_X1 U4937 ( .A1(n3711), .A2(n3938), .ZN(n3939) );
  AOI21_X1 U4938 ( .B1(n4167), .B2(EAX_REG_20__SCAN_IN), .A(n3939), .ZN(n3940)
         );
  OAI21_X1 U4939 ( .B1(n4133), .B2(n3941), .A(n3940), .ZN(n3943) );
  XNOR2_X1 U4940 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3958), .ZN(n5889)
         );
  NAND2_X1 U4941 ( .A1(n5889), .A2(n4165), .ZN(n3942) );
  NAND2_X1 U4942 ( .A1(n3943), .A2(n3942), .ZN(n5549) );
  AOI22_X1 U4943 ( .A1(n4073), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4944 ( .A1(n4152), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4145), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4945 ( .A1(n4144), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3945) );
  AOI22_X1 U4946 ( .A1(n4115), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3944) );
  NAND4_X1 U4947 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3953)
         );
  AOI22_X1 U4948 ( .A1(n4094), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4949 ( .A1(n4147), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4950 ( .A1(n4117), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3949) );
  AOI22_X1 U4951 ( .A1(n4099), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3948) );
  NAND4_X1 U4952 ( .A1(n3951), .A2(n3950), .A3(n3949), .A4(n3948), .ZN(n3952)
         );
  NOR2_X1 U4953 ( .A1(n3953), .A2(n3952), .ZN(n3957) );
  NAND2_X1 U4954 ( .A1(n6334), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3954)
         );
  NAND2_X1 U4955 ( .A1(n3711), .A2(n3954), .ZN(n3955) );
  AOI21_X1 U4956 ( .B1(n4167), .B2(EAX_REG_21__SCAN_IN), .A(n3955), .ZN(n3956)
         );
  OAI21_X1 U4957 ( .B1(n4133), .B2(n3957), .A(n3956), .ZN(n3962) );
  OAI21_X1 U4958 ( .B1(n3960), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3977), 
        .ZN(n5879) );
  OR2_X1 U4959 ( .A1(n5879), .A2(n3711), .ZN(n3961) );
  NAND2_X1 U4960 ( .A1(n3962), .A2(n3961), .ZN(n5480) );
  NOR2_X1 U4961 ( .A1(n5549), .A2(n5480), .ZN(n3963) );
  INV_X1 U4962 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U4963 ( .A1(n4142), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4964 ( .A1(n4073), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4965 ( .A1(n4147), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3965) );
  AOI22_X1 U4966 ( .A1(n4144), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3964) );
  NAND4_X1 U4967 ( .A1(n3967), .A2(n3966), .A3(n3965), .A4(n3964), .ZN(n3973)
         );
  AOI22_X1 U4968 ( .A1(n4099), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4969 ( .A1(n4145), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4970 ( .A1(n4152), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U4971 ( .A1(n4115), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3968) );
  NAND4_X1 U4972 ( .A1(n3971), .A2(n3970), .A3(n3969), .A4(n3968), .ZN(n3972)
         );
  NOR2_X1 U4973 ( .A1(n3973), .A2(n3972), .ZN(n3976) );
  AOI21_X1 U4974 ( .B1(n6841), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3974) );
  AOI21_X1 U4975 ( .B1(n4167), .B2(EAX_REG_22__SCAN_IN), .A(n3974), .ZN(n3975)
         );
  OAI21_X1 U4976 ( .B1(n4133), .B2(n3976), .A(n3975), .ZN(n3980) );
  AND2_X1 U4977 ( .A1(n3977), .A2(n6841), .ZN(n3978) );
  NOR2_X1 U4978 ( .A1(n4005), .A2(n3978), .ZN(n5869) );
  NAND2_X1 U4979 ( .A1(n5869), .A2(n4165), .ZN(n3979) );
  AOI22_X1 U4980 ( .A1(n4145), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3984) );
  AOI22_X1 U4981 ( .A1(n4143), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3983) );
  AOI22_X1 U4982 ( .A1(n4099), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4983 ( .A1(n4144), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4984 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n3981), .ZN(n3990)
         );
  AOI22_X1 U4985 ( .A1(n4147), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4986 ( .A1(n4073), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3987) );
  AOI22_X1 U4987 ( .A1(n4152), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3986) );
  AOI22_X1 U4988 ( .A1(n4115), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3985) );
  NAND4_X1 U4989 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n3989)
         );
  NOR2_X1 U4990 ( .A1(n3990), .A2(n3989), .ZN(n4011) );
  AOI22_X1 U4991 ( .A1(n4147), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4992 ( .A1(n4152), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4993 ( .A1(n4073), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4994 ( .A1(n4145), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4995 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n4000)
         );
  AOI22_X1 U4996 ( .A1(n4144), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4997 ( .A1(n4117), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4998 ( .A1(n4094), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4999 ( .A1(n4114), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U5000 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  NOR2_X1 U5001 ( .A1(n4000), .A2(n3999), .ZN(n4010) );
  XNOR2_X1 U5002 ( .A(n4011), .B(n4010), .ZN(n4004) );
  INV_X1 U5003 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4001) );
  AOI21_X1 U5004 ( .B1(n4001), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4002) );
  AOI21_X1 U5005 ( .B1(n4167), .B2(EAX_REG_23__SCAN_IN), .A(n4002), .ZN(n4003)
         );
  OAI21_X1 U5006 ( .B1(n4133), .B2(n4004), .A(n4003), .ZN(n4008) );
  OR2_X1 U5007 ( .A1(n4005), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4006)
         );
  NAND2_X1 U5008 ( .A1(n4023), .A2(n4006), .ZN(n5867) );
  NAND2_X1 U5009 ( .A1(n4008), .A2(n4007), .ZN(n5462) );
  NOR2_X1 U5010 ( .A1(n4011), .A2(n4010), .ZN(n4041) );
  AOI22_X1 U5011 ( .A1(n4142), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U5012 ( .A1(n4073), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U5013 ( .A1(n4147), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U5014 ( .A1(n4144), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U5015 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4021)
         );
  AOI22_X1 U5016 ( .A1(n4099), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U5017 ( .A1(n4145), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4018) );
  AOI22_X1 U5018 ( .A1(n4152), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U5019 ( .A1(n4115), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4016) );
  NAND4_X1 U5020 ( .A1(n4019), .A2(n4018), .A3(n4017), .A4(n4016), .ZN(n4020)
         );
  OR2_X1 U5021 ( .A1(n4021), .A2(n4020), .ZN(n4040) );
  INV_X1 U5022 ( .A(n4040), .ZN(n4022) );
  XNOR2_X1 U5023 ( .A(n4041), .B(n4022), .ZN(n4029) );
  INV_X1 U5024 ( .A(n4133), .ZN(n4163) );
  INV_X1 U5025 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4026) );
  INV_X1 U5026 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6822) );
  NAND2_X1 U5027 ( .A1(n4023), .A2(n6822), .ZN(n4024) );
  NAND2_X1 U5028 ( .A1(n4046), .A2(n4024), .ZN(n5853) );
  AOI22_X1 U5029 ( .A1(n5853), .A2(n4165), .B1(PHYADDRPOINTER_REG_24__SCAN_IN), 
        .B2(n4170), .ZN(n4025) );
  OAI21_X1 U5030 ( .B1(n4027), .B2(n4026), .A(n4025), .ZN(n4028) );
  AOI21_X1 U5031 ( .B1(n4029), .B2(n4163), .A(n4028), .ZN(n4372) );
  AOI22_X1 U5032 ( .A1(n4142), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4033) );
  AOI22_X1 U5033 ( .A1(n4147), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U5034 ( .A1(n4145), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5035 ( .A1(n4115), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4030) );
  NAND4_X1 U5036 ( .A1(n4033), .A2(n4032), .A3(n4031), .A4(n4030), .ZN(n4039)
         );
  AOI22_X1 U5037 ( .A1(n4073), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4037) );
  AOI22_X1 U5038 ( .A1(n4099), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U5039 ( .A1(n4152), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U5040 ( .A1(n4144), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4034) );
  NAND4_X1 U5041 ( .A1(n4037), .A2(n4036), .A3(n4035), .A4(n4034), .ZN(n4038)
         );
  NOR2_X1 U5042 ( .A1(n4039), .A2(n4038), .ZN(n4052) );
  NAND2_X1 U5043 ( .A1(n4041), .A2(n4040), .ZN(n4051) );
  XNOR2_X1 U5044 ( .A(n4052), .B(n4051), .ZN(n4044) );
  INV_X1 U5045 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4045) );
  OAI21_X1 U5046 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4045), .A(n3711), .ZN(
        n4042) );
  AOI21_X1 U5047 ( .B1(n4167), .B2(EAX_REG_25__SCAN_IN), .A(n4042), .ZN(n4043)
         );
  OAI21_X1 U5048 ( .B1(n4044), .B2(n4133), .A(n4043), .ZN(n4050) );
  NAND2_X1 U5049 ( .A1(n4046), .A2(n4045), .ZN(n4047) );
  NAND2_X1 U5050 ( .A1(n4086), .A2(n4047), .ZN(n5940) );
  INV_X1 U5051 ( .A(n5940), .ZN(n4048) );
  NAND2_X1 U5052 ( .A1(n4048), .A2(n4165), .ZN(n4049) );
  NOR2_X1 U5053 ( .A1(n4052), .A2(n4051), .ZN(n4081) );
  AOI22_X1 U5054 ( .A1(n4142), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U5055 ( .A1(n4073), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4055) );
  AOI22_X1 U5056 ( .A1(n4147), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5057 ( .A1(n4144), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4053) );
  NAND4_X1 U5058 ( .A1(n4056), .A2(n4055), .A3(n4054), .A4(n4053), .ZN(n4062)
         );
  AOI22_X1 U5059 ( .A1(n4099), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5060 ( .A1(n4145), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5061 ( .A1(n4152), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5062 ( .A1(n4154), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4057) );
  NAND4_X1 U5063 ( .A1(n4060), .A2(n4059), .A3(n4058), .A4(n4057), .ZN(n4061)
         );
  OR2_X1 U5064 ( .A1(n4062), .A2(n4061), .ZN(n4080) );
  INV_X1 U5065 ( .A(n4080), .ZN(n4063) );
  XNOR2_X1 U5066 ( .A(n4081), .B(n4063), .ZN(n4064) );
  NAND2_X1 U5067 ( .A1(n4064), .A2(n4163), .ZN(n4068) );
  INV_X1 U5068 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5522) );
  OAI21_X1 U5069 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5522), .A(n3711), .ZN(
        n4065) );
  AOI21_X1 U5070 ( .B1(n4167), .B2(EAX_REG_26__SCAN_IN), .A(n4065), .ZN(n4067)
         );
  XNOR2_X1 U5071 ( .A(n4086), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5834)
         );
  AOI22_X1 U5072 ( .A1(n4094), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4072) );
  AOI22_X1 U5073 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n4099), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4071) );
  AOI22_X1 U5074 ( .A1(n4154), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4070) );
  AOI22_X1 U5075 ( .A1(n4114), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4069) );
  NAND4_X1 U5076 ( .A1(n4072), .A2(n4071), .A3(n4070), .A4(n4069), .ZN(n4079)
         );
  AOI22_X1 U5077 ( .A1(n4147), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4142), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4077) );
  AOI22_X1 U5078 ( .A1(n4073), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4076) );
  AOI22_X1 U5079 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4144), .B1(n4152), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4075) );
  AOI22_X1 U5080 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3371), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4074) );
  NAND4_X1 U5081 ( .A1(n4077), .A2(n4076), .A3(n4075), .A4(n4074), .ZN(n4078)
         );
  NOR2_X1 U5082 ( .A1(n4079), .A2(n4078), .ZN(n4093) );
  NAND2_X1 U5083 ( .A1(n4081), .A2(n4080), .ZN(n4092) );
  XNOR2_X1 U5084 ( .A(n4093), .B(n4092), .ZN(n4085) );
  NAND2_X1 U5085 ( .A1(n6334), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4082)
         );
  NAND2_X1 U5086 ( .A1(n3711), .A2(n4082), .ZN(n4083) );
  AOI21_X1 U5087 ( .B1(n4167), .B2(EAX_REG_27__SCAN_IN), .A(n4083), .ZN(n4084)
         );
  OAI21_X1 U5088 ( .B1(n4085), .B2(n4133), .A(n4084), .ZN(n4091) );
  NOR2_X1 U5089 ( .A1(n4087), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4088)
         );
  OR2_X1 U5090 ( .A1(n4109), .A2(n4088), .ZN(n5827) );
  INV_X1 U5091 ( .A(n5827), .ZN(n4089) );
  NAND2_X1 U5092 ( .A1(n4089), .A2(n4165), .ZN(n4090) );
  NAND2_X1 U5093 ( .A1(n4091), .A2(n4090), .ZN(n5515) );
  NOR2_X1 U5094 ( .A1(n4093), .A2(n4092), .ZN(n4129) );
  AOI22_X1 U5095 ( .A1(n4142), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5096 ( .A1(n4073), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4097) );
  AOI22_X1 U5097 ( .A1(n4147), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4096) );
  AOI22_X1 U5098 ( .A1(n4144), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4095) );
  NAND4_X1 U5099 ( .A1(n4098), .A2(n4097), .A3(n4096), .A4(n4095), .ZN(n4105)
         );
  AOI22_X1 U5100 ( .A1(n4099), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5101 ( .A1(n4145), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4117), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4102) );
  AOI22_X1 U5102 ( .A1(n4152), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5103 ( .A1(n4154), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4100) );
  NAND4_X1 U5104 ( .A1(n4103), .A2(n4102), .A3(n4101), .A4(n4100), .ZN(n4104)
         );
  OR2_X1 U5105 ( .A1(n4105), .A2(n4104), .ZN(n4128) );
  XNOR2_X1 U5106 ( .A(n4129), .B(n4128), .ZN(n4108) );
  INV_X1 U5107 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n6998) );
  OAI21_X1 U5108 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6998), .A(n3711), .ZN(
        n4106) );
  AOI21_X1 U5109 ( .B1(n4167), .B2(EAX_REG_28__SCAN_IN), .A(n4106), .ZN(n4107)
         );
  OAI21_X1 U5110 ( .B1(n4108), .B2(n4133), .A(n4107), .ZN(n4112) );
  NOR2_X1 U5111 ( .A1(n4109), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4110)
         );
  NAND2_X1 U5112 ( .A1(n5817), .A2(n4165), .ZN(n4111) );
  NAND2_X1 U5113 ( .A1(n4112), .A2(n4111), .ZN(n5433) );
  AOI22_X1 U5114 ( .A1(n4142), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4121) );
  AOI22_X1 U5115 ( .A1(n4152), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4120) );
  AOI22_X1 U5116 ( .A1(n4145), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4115), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U5117 ( .A1(n4117), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4118) );
  NAND4_X1 U5118 ( .A1(n4121), .A2(n4120), .A3(n4119), .A4(n4118), .ZN(n4127)
         );
  AOI22_X1 U5119 ( .A1(n4073), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4144), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5120 ( .A1(n4094), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5121 ( .A1(n4147), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4123) );
  AOI22_X1 U5122 ( .A1(n4153), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4122) );
  NAND4_X1 U5123 ( .A1(n4125), .A2(n4124), .A3(n4123), .A4(n4122), .ZN(n4126)
         );
  NOR2_X1 U5124 ( .A1(n4127), .A2(n4126), .ZN(n4141) );
  NAND2_X1 U5125 ( .A1(n4129), .A2(n4128), .ZN(n4140) );
  XNOR2_X1 U5126 ( .A(n4141), .B(n4140), .ZN(n4134) );
  NAND2_X1 U5127 ( .A1(n6334), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4130)
         );
  NAND2_X1 U5128 ( .A1(n3711), .A2(n4130), .ZN(n4131) );
  AOI21_X1 U5129 ( .B1(n4167), .B2(EAX_REG_29__SCAN_IN), .A(n4131), .ZN(n4132)
         );
  OAI21_X1 U5130 ( .B1(n4134), .B2(n4133), .A(n4132), .ZN(n4139) );
  OR2_X1 U5131 ( .A1(n4135), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4136)
         );
  NAND2_X1 U5132 ( .A1(n4136), .A2(n4173), .ZN(n5808) );
  INV_X1 U5133 ( .A(n5808), .ZN(n4137) );
  NAND2_X1 U5134 ( .A1(n4137), .A2(n4165), .ZN(n4138) );
  NAND2_X1 U5135 ( .A1(n4139), .A2(n4138), .ZN(n5422) );
  NOR2_X1 U5136 ( .A1(n4141), .A2(n4140), .ZN(n4162) );
  AOI22_X1 U5137 ( .A1(n4142), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4094), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5138 ( .A1(n4144), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4143), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4150) );
  AOI22_X1 U5139 ( .A1(n4145), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4099), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4149) );
  AOI22_X1 U5140 ( .A1(n4147), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4146), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4148) );
  NAND4_X1 U5141 ( .A1(n4151), .A2(n4150), .A3(n4149), .A4(n4148), .ZN(n4160)
         );
  AOI22_X1 U5142 ( .A1(n4152), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4114), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5143 ( .A1(n4117), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4116), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5144 ( .A1(n4154), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4153), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4156) );
  AOI22_X1 U5145 ( .A1(n4073), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3365), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4155) );
  NAND4_X1 U5146 ( .A1(n4158), .A2(n4157), .A3(n4156), .A4(n4155), .ZN(n4159)
         );
  NOR2_X1 U5147 ( .A1(n4160), .A2(n4159), .ZN(n4161) );
  XNOR2_X1 U5148 ( .A(n4162), .B(n4161), .ZN(n4164) );
  NAND2_X1 U5149 ( .A1(n4164), .A2(n4163), .ZN(n4169) );
  INV_X1 U5150 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4429) );
  NOR2_X1 U5151 ( .A1(n4429), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4166) );
  AOI211_X1 U5152 ( .C1(n4167), .C2(EAX_REG_30__SCAN_IN), .A(n4166), .B(n4165), 
        .ZN(n4168) );
  XNOR2_X1 U5153 ( .A(n4173), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4437)
         );
  INV_X1 U5154 ( .A(n5419), .ZN(n4172) );
  AND2_X1 U5155 ( .A1(n6576), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5156 ( .A1(n4390), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6590) );
  NAND2_X1 U5157 ( .A1(n4172), .A2(n6223), .ZN(n4181) );
  NAND2_X1 U5158 ( .A1(n6695), .A2(n6694), .ZN(n4175) );
  NAND2_X1 U5159 ( .A1(n4175), .A2(n6576), .ZN(n4176) );
  NAND2_X1 U5160 ( .A1(n6576), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4178) );
  NAND2_X1 U5161 ( .A1(n5991), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4177) );
  NAND2_X1 U5162 ( .A1(n4178), .A2(n4177), .ZN(n4487) );
  INV_X1 U5163 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6835) );
  NAND2_X1 U5164 ( .A1(n6317), .A2(REIP_REG_31__SCAN_IN), .ZN(n5605) );
  OAI21_X1 U5165 ( .B1(n5955), .B2(n6835), .A(n5605), .ZN(n4179) );
  OAI211_X1 U5166 ( .C1(n5613), .C2(n6213), .A(n4181), .B(n4180), .ZN(U2955)
         );
  XNOR2_X1 U5167 ( .A(n5582), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5696)
         );
  XNOR2_X1 U5168 ( .A(n5582), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5548)
         );
  INV_X1 U5169 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6759) );
  XNOR2_X1 U5170 ( .A(n5582), .B(n6774), .ZN(n5541) );
  NOR2_X1 U5171 ( .A1(n5582), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5534)
         );
  NAND2_X1 U5172 ( .A1(n5540), .A2(n5534), .ZN(n5527) );
  INV_X1 U5173 ( .A(n5527), .ZN(n4183) );
  NAND2_X1 U5174 ( .A1(n4183), .A2(n4182), .ZN(n4187) );
  NAND2_X1 U5175 ( .A1(n5535), .A2(n4185), .ZN(n4186) );
  INV_X1 U5176 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4365) );
  NAND2_X1 U5177 ( .A1(n6541), .A2(n4496), .ZN(n4343) );
  NOR2_X1 U5178 ( .A1(n4690), .A2(n3346), .ZN(n4190) );
  NAND2_X1 U5179 ( .A1(n4190), .A2(n4189), .ZN(n4329) );
  NAND2_X1 U5180 ( .A1(n4329), .A2(n4191), .ZN(n4194) );
  AND2_X1 U5181 ( .A1(n4192), .A2(n4193), .ZN(n4389) );
  INV_X1 U5182 ( .A(n4389), .ZN(n4447) );
  OAI21_X1 U5183 ( .B1(n4532), .B2(n4194), .A(n4447), .ZN(n4542) );
  NAND2_X1 U5184 ( .A1(n4195), .A2(n6777), .ZN(n6598) );
  NAND2_X1 U5185 ( .A1(n4496), .A2(n6598), .ZN(n4204) );
  INV_X1 U5186 ( .A(n4196), .ZN(n4197) );
  NOR4_X1 U5187 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4201)
         );
  NOR2_X1 U5188 ( .A1(n4202), .A2(n4201), .ZN(n4448) );
  INV_X1 U5189 ( .A(n4448), .ZN(n4203) );
  NOR2_X1 U5190 ( .A1(READY_N), .A2(n4203), .ZN(n4533) );
  NAND3_X1 U5191 ( .A1(n4204), .A2(n4533), .A3(n4543), .ZN(n4205) );
  OAI211_X1 U5192 ( .C1(n4547), .C2(n4343), .A(n4542), .B(n4205), .ZN(n4206)
         );
  NAND2_X1 U5193 ( .A1(n4206), .A2(n6583), .ZN(n4211) );
  NAND2_X1 U5194 ( .A1(n4752), .A2(n6598), .ZN(n4395) );
  INV_X1 U5195 ( .A(READY_N), .ZN(n4495) );
  AND2_X1 U5196 ( .A1(n4395), .A2(n4495), .ZN(n4538) );
  NAND2_X1 U5197 ( .A1(n4540), .A2(n4538), .ZN(n4208) );
  AOI21_X1 U5198 ( .B1(n4208), .B2(n3126), .A(n4543), .ZN(n4209) );
  NAND2_X1 U5199 ( .A1(n4477), .A2(n4209), .ZN(n4210) );
  OR2_X1 U5200 ( .A1(n4537), .A2(n4752), .ZN(n4218) );
  INV_X1 U5201 ( .A(n4532), .ZN(n4215) );
  NAND2_X1 U5202 ( .A1(n3355), .A2(n4322), .ZN(n4214) );
  NAND2_X1 U5203 ( .A1(n4215), .A2(n4214), .ZN(n4446) );
  INV_X1 U5204 ( .A(n4221), .ZN(n4216) );
  NAND2_X1 U5205 ( .A1(n4216), .A2(n4220), .ZN(n4217) );
  NAND4_X1 U5206 ( .A1(n4605), .A2(n4218), .A3(n4446), .A4(n4217), .ZN(n4219)
         );
  NAND2_X1 U5207 ( .A1(n4370), .A2(n6315), .ZN(n4369) );
  NAND2_X1 U5208 ( .A1(n4540), .A2(n4445), .ZN(n6571) );
  OAI21_X1 U5209 ( .B1(n4221), .B2(n4220), .A(n6571), .ZN(n4222) );
  BUF_X2 U5210 ( .A(n4297), .Z(n4420) );
  INV_X1 U5211 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4223) );
  NAND2_X1 U5212 ( .A1(n4233), .A2(n4223), .ZN(n4227) );
  NAND2_X1 U5213 ( .A1(n4224), .A2(n4529), .ZN(n4225) );
  OAI211_X1 U5214 ( .C1(n4420), .C2(EBX_REG_1__SCAN_IN), .A(n5683), .B(n4225), 
        .ZN(n4226) );
  NAND2_X1 U5215 ( .A1(n4224), .A2(EBX_REG_0__SCAN_IN), .ZN(n4229) );
  INV_X1 U5216 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U5217 ( .A1(n5683), .A2(n6827), .ZN(n4228) );
  AND2_X1 U5218 ( .A1(n4229), .A2(n4228), .ZN(n4471) );
  OR2_X1 U5219 ( .A1(n4465), .A2(n4420), .ZN(n4466) );
  CLKBUF_X3 U5220 ( .A(n4297), .Z(n5406) );
  MUX2_X1 U5221 ( .A(n4412), .B(n5698), .S(EBX_REG_3__SCAN_IN), .Z(n4232) );
  NOR2_X1 U5222 ( .A1(n5407), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4231)
         );
  INV_X2 U5223 ( .A(n4240), .ZN(n4416) );
  INV_X1 U5224 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4234) );
  NAND2_X1 U5225 ( .A1(n4416), .A2(n4234), .ZN(n4238) );
  NAND2_X1 U5226 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4235)
         );
  NAND2_X1 U5227 ( .A1(n4224), .A2(n4235), .ZN(n4236) );
  OAI21_X1 U5228 ( .B1(n4420), .B2(EBX_REG_2__SCAN_IN), .A(n4236), .ZN(n4237)
         );
  NAND2_X1 U5229 ( .A1(n4238), .A2(n4237), .ZN(n5118) );
  NAND2_X1 U5230 ( .A1(n4620), .A2(n5118), .ZN(n4239) );
  NOR2_X2 U5231 ( .A1(n4619), .A2(n4239), .ZN(n4634) );
  INV_X1 U5232 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U5233 ( .A1(n4416), .A2(n4241), .ZN(n4244) );
  NAND2_X1 U5234 ( .A1(n4224), .A2(n6979), .ZN(n4242) );
  OAI211_X1 U5235 ( .C1(n4420), .C2(EBX_REG_4__SCAN_IN), .A(n5683), .B(n4242), 
        .ZN(n4243) );
  NAND2_X1 U5236 ( .A1(n4244), .A2(n4243), .ZN(n4633) );
  NAND2_X1 U5237 ( .A1(n4634), .A2(n4633), .ZN(n4632) );
  INV_X1 U5238 ( .A(n4632), .ZN(n4248) );
  MUX2_X1 U5239 ( .A(n4412), .B(n5698), .S(EBX_REG_5__SCAN_IN), .Z(n4245) );
  INV_X1 U5240 ( .A(n4245), .ZN(n4247) );
  NAND2_X1 U5241 ( .A1(n4472), .A2(n6275), .ZN(n4246) );
  INV_X1 U5242 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4783) );
  NAND2_X1 U5243 ( .A1(n4416), .A2(n4783), .ZN(n4252) );
  NAND2_X1 U5244 ( .A1(n4224), .A2(n4249), .ZN(n4250) );
  OAI211_X1 U5245 ( .C1(n5406), .C2(EBX_REG_6__SCAN_IN), .A(n5683), .B(n4250), 
        .ZN(n4251) );
  MUX2_X1 U5246 ( .A(n4412), .B(n5698), .S(EBX_REG_7__SCAN_IN), .Z(n4253) );
  INV_X1 U5247 ( .A(n4253), .ZN(n4254) );
  NAND2_X1 U5248 ( .A1(n4254), .A2(n3176), .ZN(n4730) );
  INV_X1 U5249 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U5250 ( .A1(n4416), .A2(n4255), .ZN(n4259) );
  NAND2_X1 U5251 ( .A1(n4224), .A2(n4256), .ZN(n4257) );
  OAI211_X1 U5252 ( .C1(n5406), .C2(EBX_REG_8__SCAN_IN), .A(n5683), .B(n4257), 
        .ZN(n4258) );
  NAND2_X1 U5253 ( .A1(n4259), .A2(n4258), .ZN(n4775) );
  INV_X1 U5254 ( .A(n4984), .ZN(n4263) );
  MUX2_X1 U5255 ( .A(n4412), .B(n5698), .S(EBX_REG_9__SCAN_IN), .Z(n4260) );
  INV_X1 U5256 ( .A(n4260), .ZN(n4261) );
  NAND2_X1 U5257 ( .A1(n4261), .A2(n3177), .ZN(n4985) );
  INV_X1 U5258 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4264) );
  NAND2_X1 U5259 ( .A1(n4416), .A2(n4264), .ZN(n4268) );
  NAND2_X1 U5260 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U5261 ( .A1(n4224), .A2(n4265), .ZN(n4266) );
  OAI21_X1 U5262 ( .B1(n4420), .B2(EBX_REG_10__SCAN_IN), .A(n4266), .ZN(n4267)
         );
  NOR2_X2 U5263 ( .A1(n5090), .A2(n5089), .ZN(n5185) );
  MUX2_X1 U5264 ( .A(n4412), .B(n5698), .S(EBX_REG_11__SCAN_IN), .Z(n4270) );
  NOR2_X1 U5265 ( .A1(n5407), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4269)
         );
  NOR2_X1 U5266 ( .A1(n4270), .A2(n4269), .ZN(n5184) );
  INV_X1 U5267 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6871) );
  NAND2_X1 U5268 ( .A1(n4416), .A2(n6871), .ZN(n4273) );
  NAND2_X1 U5269 ( .A1(n4224), .A2(n6927), .ZN(n4271) );
  OAI211_X1 U5270 ( .C1(n4420), .C2(EBX_REG_12__SCAN_IN), .A(n5683), .B(n4271), 
        .ZN(n4272) );
  MUX2_X1 U5271 ( .A(n4412), .B(n5698), .S(EBX_REG_13__SCAN_IN), .Z(n4274) );
  INV_X1 U5272 ( .A(n4274), .ZN(n4276) );
  NAND2_X1 U5273 ( .A1(n4472), .A2(n6949), .ZN(n4275) );
  NAND2_X1 U5274 ( .A1(n4276), .A2(n4275), .ZN(n5258) );
  INV_X1 U5275 ( .A(EBX_REG_14__SCAN_IN), .ZN(n4278) );
  NAND2_X1 U5276 ( .A1(n4416), .A2(n4278), .ZN(n4282) );
  NAND2_X1 U5277 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U5278 ( .A1(n4224), .A2(n4279), .ZN(n4280) );
  OAI21_X1 U5279 ( .B1(n5406), .B2(EBX_REG_14__SCAN_IN), .A(n4280), .ZN(n4281)
         );
  NAND2_X1 U5280 ( .A1(n4282), .A2(n4281), .ZN(n5331) );
  NAND2_X1 U5281 ( .A1(n5332), .A2(n5331), .ZN(n5739) );
  INV_X1 U5282 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U5283 ( .A1(n4412), .A2(n6122), .ZN(n4285) );
  NAND2_X1 U5284 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4283) );
  OAI211_X1 U5285 ( .C1(n4420), .C2(EBX_REG_15__SCAN_IN), .A(n4224), .B(n4283), 
        .ZN(n4284) );
  NAND2_X1 U5286 ( .A1(n4285), .A2(n4284), .ZN(n5740) );
  OR2_X2 U5287 ( .A1(n5739), .A2(n5740), .ZN(n5737) );
  INV_X1 U5288 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U5289 ( .A1(n4412), .A2(n6918), .ZN(n4288) );
  NAND2_X1 U5290 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4286) );
  OAI211_X1 U5291 ( .C1(n5406), .C2(EBX_REG_17__SCAN_IN), .A(n4224), .B(n4286), 
        .ZN(n4287) );
  AND2_X1 U5292 ( .A1(n4288), .A2(n4287), .ZN(n5725) );
  INV_X1 U5293 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5379) );
  NAND2_X1 U5294 ( .A1(n4416), .A2(n5379), .ZN(n4292) );
  NAND2_X1 U5295 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U5296 ( .A1(n4224), .A2(n4289), .ZN(n4290) );
  OAI21_X1 U5297 ( .B1(n5406), .B2(EBX_REG_16__SCAN_IN), .A(n4290), .ZN(n4291)
         );
  NAND2_X1 U5298 ( .A1(n4292), .A2(n4291), .ZN(n5724) );
  NAND2_X1 U5299 ( .A1(n5725), .A2(n5724), .ZN(n4293) );
  OR2_X2 U5300 ( .A1(n5737), .A2(n4293), .ZN(n5728) );
  INV_X1 U5301 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U5302 ( .A1(n4416), .A2(n5915), .ZN(n4296) );
  INV_X1 U5303 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U5304 ( .A1(n4224), .A2(n5705), .ZN(n4294) );
  OAI211_X1 U5305 ( .C1(n5406), .C2(EBX_REG_19__SCAN_IN), .A(n5683), .B(n4294), 
        .ZN(n4295) );
  NOR2_X2 U5306 ( .A1(n5728), .A2(n5702), .ZN(n5681) );
  INV_X1 U5307 ( .A(EBX_REG_20__SCAN_IN), .ZN(n4302) );
  NAND2_X1 U5308 ( .A1(n4472), .A2(n5716), .ZN(n4299) );
  INV_X1 U5309 ( .A(n4297), .ZN(n4467) );
  INV_X1 U5310 ( .A(EBX_REG_18__SCAN_IN), .ZN(n4298) );
  NAND2_X1 U5311 ( .A1(n4467), .A2(n4298), .ZN(n5697) );
  OAI22_X1 U5312 ( .A1(n5407), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n5406), .B2(EBX_REG_20__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U5313 ( .A1(n5700), .A2(n5684), .ZN(n4301) );
  INV_X1 U5314 ( .A(n5700), .ZN(n5682) );
  NAND2_X1 U5315 ( .A1(n5682), .A2(n5683), .ZN(n4300) );
  OAI211_X1 U5316 ( .C1(n5683), .C2(n4302), .A(n4301), .B(n4300), .ZN(n4303)
         );
  INV_X1 U5317 ( .A(n4303), .ZN(n4304) );
  AND2_X2 U5318 ( .A1(n5681), .A2(n4304), .ZN(n5482) );
  INV_X1 U5319 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U5320 ( .A1(n4412), .A2(n5484), .ZN(n4307) );
  NAND2_X1 U5321 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4305) );
  OAI211_X1 U5322 ( .C1(n4420), .C2(EBX_REG_21__SCAN_IN), .A(n4224), .B(n4305), 
        .ZN(n4306) );
  NAND2_X1 U5323 ( .A1(n5482), .A2(n5481), .ZN(n5471) );
  INV_X1 U5324 ( .A(EBX_REG_22__SCAN_IN), .ZN(n6888) );
  NAND2_X1 U5325 ( .A1(n4416), .A2(n6888), .ZN(n4311) );
  NAND2_X1 U5326 ( .A1(n4224), .A2(n4308), .ZN(n4309) );
  OAI211_X1 U5327 ( .C1(n4420), .C2(EBX_REG_22__SCAN_IN), .A(n5683), .B(n4309), 
        .ZN(n4310) );
  OR2_X2 U5328 ( .A1(n5471), .A2(n5472), .ZN(n5474) );
  INV_X1 U5329 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U5330 ( .A1(n4412), .A2(n5465), .ZN(n4314) );
  NAND2_X1 U5331 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4312) );
  OAI211_X1 U5332 ( .C1(n5406), .C2(EBX_REG_23__SCAN_IN), .A(n4224), .B(n4312), 
        .ZN(n4313) );
  NAND2_X1 U5333 ( .A1(n4314), .A2(n4313), .ZN(n5464) );
  NOR2_X2 U5334 ( .A1(n5474), .A2(n5464), .ZN(n4319) );
  INV_X1 U5335 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U5336 ( .A1(n4416), .A2(n5458), .ZN(n4317) );
  NAND2_X1 U5337 ( .A1(n4224), .A2(n4365), .ZN(n4315) );
  OAI211_X1 U5338 ( .C1(n5406), .C2(EBX_REG_24__SCAN_IN), .A(n5683), .B(n4315), 
        .ZN(n4316) );
  NAND2_X1 U5339 ( .A1(n4317), .A2(n4316), .ZN(n4318) );
  NAND2_X1 U5340 ( .A1(n4319), .A2(n4318), .ZN(n4408) );
  OR2_X1 U5341 ( .A1(n4319), .A2(n4318), .ZN(n4320) );
  NAND2_X1 U5342 ( .A1(n4408), .A2(n4320), .ZN(n5859) );
  INV_X1 U5343 ( .A(n5859), .ZN(n4367) );
  INV_X1 U5344 ( .A(REIP_REG_24__SCAN_IN), .ZN(n4321) );
  NOR2_X1 U5345 ( .A1(n6292), .A2(n4321), .ZN(n4376) );
  NOR2_X1 U5346 ( .A1(n6979), .A2(n6808), .ZN(n6747) );
  NOR2_X1 U5347 ( .A1(n3476), .A2(n4529), .ZN(n6309) );
  AND2_X1 U5348 ( .A1(n6747), .A2(n6309), .ZN(n6278) );
  NAND3_X1 U5349 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n6278), .ZN(n6237) );
  NAND2_X1 U5350 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6260) );
  INV_X1 U5351 ( .A(n6260), .ZN(n6243) );
  NAND3_X1 U5352 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6243), .ZN(n4345) );
  NOR2_X1 U5353 ( .A1(n6237), .A2(n4345), .ZN(n4354) );
  NOR2_X1 U5354 ( .A1(n4322), .A2(n4544), .ZN(n4323) );
  NOR2_X1 U5355 ( .A1(n5749), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4673)
         );
  INV_X1 U5356 ( .A(n4673), .ZN(n4342) );
  AOI22_X1 U5357 ( .A1(n5115), .A2(n4457), .B1(n4543), .B2(n4324), .ZN(n4328)
         );
  INV_X1 U5358 ( .A(n4325), .ZN(n4326) );
  NAND2_X1 U5359 ( .A1(n4326), .A2(n5407), .ZN(n4327) );
  AND2_X1 U5360 ( .A1(n4328), .A2(n4327), .ZN(n4330) );
  OAI211_X1 U5361 ( .C1(n3350), .C2(n5683), .A(n4330), .B(n4329), .ZN(n4331)
         );
  INV_X1 U5362 ( .A(n4331), .ZN(n4332) );
  NAND2_X1 U5363 ( .A1(n4333), .A2(n4332), .ZN(n4344) );
  INV_X1 U5364 ( .A(n4344), .ZN(n4522) );
  INV_X1 U5365 ( .A(n4335), .ZN(n4337) );
  INV_X1 U5366 ( .A(n4338), .ZN(n4340) );
  OR2_X1 U5367 ( .A1(n4339), .A2(n3289), .ZN(n4583) );
  NAND3_X1 U5368 ( .A1(n4522), .A2(n4340), .A3(n4583), .ZN(n4341) );
  NAND2_X1 U5369 ( .A1(n4349), .A2(n4571), .ZN(n6288) );
  INV_X1 U5370 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4528) );
  OAI21_X1 U5371 ( .B1(n4529), .B2(n4528), .A(n3476), .ZN(n6291) );
  NAND2_X1 U5372 ( .A1(n6747), .A2(n6291), .ZN(n6276) );
  NOR2_X1 U5373 ( .A1(n6275), .A2(n6276), .ZN(n4814) );
  NAND2_X1 U5374 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4814), .ZN(n6242)
         );
  NOR2_X1 U5375 ( .A1(n4345), .A2(n6242), .ZN(n4353) );
  INV_X1 U5376 ( .A(n6236), .ZN(n5344) );
  NAND3_X1 U5377 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n5748) );
  NOR2_X1 U5378 ( .A1(n3606), .A2(n5748), .ZN(n4356) );
  NAND2_X1 U5379 ( .A1(n5344), .A2(n4356), .ZN(n5736) );
  NAND3_X1 U5380 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n5967), .ZN(n5732) );
  NOR2_X1 U5381 ( .A1(n5731), .A2(n5732), .ZN(n5717) );
  INV_X1 U5382 ( .A(n4346), .ZN(n5526) );
  INV_X1 U5383 ( .A(n5663), .ZN(n4364) );
  NAND2_X1 U5384 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4347) );
  AND2_X1 U5385 ( .A1(n5688), .A2(n4347), .ZN(n4348) );
  NAND2_X1 U5386 ( .A1(n5706), .A2(n4348), .ZN(n5668) );
  NAND2_X1 U5387 ( .A1(n5753), .A2(n4528), .ZN(n4352) );
  INV_X1 U5388 ( .A(n4349), .ZN(n4350) );
  NAND2_X1 U5389 ( .A1(n4350), .A2(n6292), .ZN(n4351) );
  INV_X1 U5390 ( .A(n6239), .ZN(n6233) );
  INV_X1 U5391 ( .A(n6238), .ZN(n4815) );
  OAI22_X1 U5392 ( .A1(n4815), .A2(n4354), .B1(n4353), .B2(n6288), .ZN(n4355)
         );
  NOR2_X1 U5393 ( .A1(n6233), .A2(n4355), .ZN(n5751) );
  OAI21_X1 U5394 ( .B1(n5599), .B2(n4356), .A(n5751), .ZN(n5964) );
  AND2_X1 U5395 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4357) );
  NOR2_X1 U5396 ( .A1(n5599), .A2(n4357), .ZN(n4358) );
  NOR2_X1 U5397 ( .A1(n5964), .A2(n4358), .ZN(n5730) );
  OR2_X1 U5398 ( .A1(n5599), .A2(n4359), .ZN(n4360) );
  NAND2_X1 U5399 ( .A1(n5730), .A2(n4360), .ZN(n5712) );
  NOR2_X1 U5400 ( .A1(n5599), .A2(n5688), .ZN(n4361) );
  NOR2_X1 U5401 ( .A1(n5712), .A2(n4361), .ZN(n5674) );
  OAI21_X1 U5402 ( .B1(n6318), .B2(n6310), .A(n5600), .ZN(n4362) );
  AOI211_X1 U5403 ( .C1(n4365), .C2(n4364), .A(n4363), .B(n5961), .ZN(n4366)
         );
  AOI211_X1 U5404 ( .C1(n5611), .C2(n4367), .A(n4376), .B(n4366), .ZN(n4368)
         );
  NAND2_X1 U5405 ( .A1(n4369), .A2(n4368), .ZN(U2994) );
  NAND2_X1 U5406 ( .A1(n4370), .A2(n6224), .ZN(n4380) );
  AND2_X1 U5407 ( .A1(n4371), .A2(n4372), .ZN(n4374) );
  OR2_X1 U5408 ( .A1(n4374), .A2(n4373), .ZN(n5855) );
  NOR2_X1 U5409 ( .A1(n6228), .A2(n5853), .ZN(n4375) );
  AOI211_X1 U5410 ( .C1(n6218), .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n4376), 
        .B(n4375), .ZN(n4377) );
  NAND2_X1 U5411 ( .A1(n4380), .A2(n4379), .ZN(U2962) );
  NOR2_X1 U5412 ( .A1(n5496), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4383)
         );
  XNOR2_X1 U5413 ( .A(n4384), .B(n5614), .ZN(n5623) );
  NAND2_X1 U5414 ( .A1(n6317), .A2(REIP_REG_30__SCAN_IN), .ZN(n5615) );
  OAI21_X1 U5415 ( .B1(n5955), .B2(n4429), .A(n5615), .ZN(n4386) );
  AOI21_X1 U5416 ( .B1(n6196), .B2(n4437), .A(n4386), .ZN(n4387) );
  OAI211_X1 U5417 ( .C1(n5623), .C2(n6213), .A(n3120), .B(n4387), .ZN(U2956)
         );
  NAND2_X1 U5418 ( .A1(n4448), .A2(n4389), .ZN(n4443) );
  INV_X1 U5419 ( .A(n6583), .ZN(n6581) );
  NOR2_X1 U5420 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6701) );
  NOR3_X1 U5421 ( .A1(n6576), .A2(n6662), .A3(n6578), .ZN(n6574) );
  INV_X1 U5422 ( .A(n6574), .ZN(n4391) );
  NAND2_X1 U5423 ( .A1(n4390), .A2(n4165), .ZN(n6587) );
  INV_X1 U5424 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6807) );
  INV_X1 U5425 ( .A(REIP_REG_27__SCAN_IN), .ZN(n5829) );
  NOR2_X1 U5426 ( .A1(n6807), .A2(n5829), .ZN(n4398) );
  NAND3_X1 U5427 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4402) );
  NAND3_X1 U5428 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .A3(
        REIP_REG_16__SCAN_IN), .ZN(n4394) );
  INV_X1 U5429 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6897) );
  INV_X1 U5430 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6615) );
  NAND3_X1 U5431 ( .A1(REIP_REG_3__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6072) );
  OR2_X1 U5432 ( .A1(n6615), .A2(n6072), .ZN(n5073) );
  NOR2_X1 U5433 ( .A1(n6897), .A2(n5073), .ZN(n5079) );
  INV_X1 U5434 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U5435 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n5104) );
  NOR2_X1 U5436 ( .A1(n6621), .A2(n5104), .ZN(n6039) );
  AND4_X1 U5437 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n5079), .A4(n6039), .ZN(n6030) );
  NAND2_X1 U5438 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6030), .ZN(n5262) );
  INV_X1 U5439 ( .A(n5262), .ZN(n5260) );
  NAND2_X1 U5440 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5260), .ZN(n4401) );
  NOR2_X1 U5441 ( .A1(n6095), .A2(n4401), .ZN(n5274) );
  NAND3_X1 U5442 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        n5274), .ZN(n5328) );
  NOR2_X1 U5443 ( .A1(n4394), .A2(n5328), .ZN(n5900) );
  NAND4_X1 U5444 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5868), .ZN(n5843) );
  NOR2_X1 U5445 ( .A1(n4402), .A2(n5843), .ZN(n5825) );
  NOR2_X1 U5446 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4431) );
  INV_X1 U5447 ( .A(n4431), .ZN(n4430) );
  NOR2_X1 U5448 ( .A1(n3346), .A2(n4430), .ZN(n4396) );
  AND2_X1 U5449 ( .A1(n4396), .A2(n4395), .ZN(n4397) );
  NAND2_X1 U5450 ( .A1(n6092), .A2(n5113), .ZN(n6105) );
  AOI21_X1 U5451 ( .B1(n4398), .B2(n5825), .A(n5901), .ZN(n5816) );
  INV_X1 U5452 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6650) );
  NAND2_X1 U5453 ( .A1(n6105), .A2(n6650), .ZN(n4399) );
  NAND2_X1 U5454 ( .A1(n4399), .A2(REIP_REG_30__SCAN_IN), .ZN(n4400) );
  NOR2_X1 U5455 ( .A1(n5816), .A2(n4400), .ZN(n5411) );
  INV_X1 U5456 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6637) );
  INV_X1 U5457 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6635) );
  INV_X1 U5458 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U5459 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5270), .ZN(n5329) );
  NAND4_X1 U5460 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5370), .A3(
        REIP_REG_15__SCAN_IN), .A4(REIP_REG_16__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U5461 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5896), .ZN(n5886) );
  NAND4_X1 U5462 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5881), .ZN(n5854) );
  NAND3_X1 U5463 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .A3(
        n5830), .ZN(n5815) );
  NOR2_X1 U5464 ( .A1(n6650), .A2(n5815), .ZN(n5399) );
  NOR2_X1 U5465 ( .A1(REIP_REG_30__SCAN_IN), .A2(n5399), .ZN(n4403) );
  OAI22_X1 U5466 ( .A1(n5391), .A2(n6044), .B1(n5411), .B2(n4403), .ZN(n4404)
         );
  MUX2_X1 U5467 ( .A(n4412), .B(n5698), .S(EBX_REG_25__SCAN_IN), .Z(n4405) );
  INV_X1 U5468 ( .A(n4405), .ZN(n4407) );
  NAND2_X1 U5469 ( .A1(n4472), .A2(n6788), .ZN(n4406) );
  NAND2_X1 U5470 ( .A1(n4407), .A2(n4406), .ZN(n5451) );
  OR2_X2 U5471 ( .A1(n4408), .A2(n5451), .ZN(n5453) );
  INV_X1 U5472 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U5473 ( .A1(n4416), .A2(n5842), .ZN(n4411) );
  NAND2_X1 U5474 ( .A1(n4224), .A2(n5520), .ZN(n4409) );
  OAI211_X1 U5475 ( .C1(n4420), .C2(EBX_REG_26__SCAN_IN), .A(n5683), .B(n4409), 
        .ZN(n4410) );
  AND2_X1 U5476 ( .A1(n4411), .A2(n4410), .ZN(n5444) );
  INV_X1 U5477 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U5478 ( .A1(n4412), .A2(n5909), .ZN(n4415) );
  NAND2_X1 U5479 ( .A1(n5683), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4413) );
  OAI211_X1 U5480 ( .C1(n4420), .C2(EBX_REG_27__SCAN_IN), .A(n4224), .B(n4413), 
        .ZN(n4414) );
  NAND2_X1 U5481 ( .A1(n4415), .A2(n4414), .ZN(n5640) );
  INV_X1 U5482 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U5483 ( .A1(n4416), .A2(n6761), .ZN(n4419) );
  NAND2_X1 U5484 ( .A1(n4224), .A2(n5505), .ZN(n4417) );
  OAI211_X1 U5485 ( .C1(n5406), .C2(EBX_REG_28__SCAN_IN), .A(n5683), .B(n4417), 
        .ZN(n4418) );
  NAND2_X1 U5486 ( .A1(n4419), .A2(n4418), .ZN(n5436) );
  INV_X1 U5487 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5431) );
  AOI22_X1 U5488 ( .A1(n4472), .A2(n5624), .B1(n4467), .B2(n5431), .ZN(n5425)
         );
  NAND2_X1 U5489 ( .A1(n5407), .A2(EBX_REG_30__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5490 ( .A1(n4420), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4421) );
  AND2_X1 U5491 ( .A1(n4422), .A2(n4421), .ZN(n5402) );
  NOR2_X1 U5492 ( .A1(n4423), .A2(n5698), .ZN(n5403) );
  INV_X1 U5493 ( .A(n3117), .ZN(n5400) );
  INV_X1 U5494 ( .A(n5402), .ZN(n4424) );
  AOI211_X1 U5495 ( .C1(n5698), .C2(n5400), .A(n4424), .B(n4423), .ZN(n4425)
         );
  NOR2_X1 U5496 ( .A1(n4426), .A2(n4425), .ZN(n5618) );
  NAND2_X1 U5497 ( .A1(n4430), .A2(EBX_REG_31__SCAN_IN), .ZN(n4427) );
  NOR2_X1 U5498 ( .A1(n5406), .A2(n4427), .ZN(n4428) );
  NOR2_X2 U5499 ( .A1(n6095), .A2(n6662), .ZN(n6083) );
  INV_X1 U5500 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5421) );
  NAND2_X1 U5501 ( .A1(n5421), .A2(n4430), .ZN(n4432) );
  INV_X1 U5502 ( .A(n6598), .ZN(n4479) );
  NAND2_X1 U5503 ( .A1(n4479), .A2(n4431), .ZN(n6570) );
  NAND2_X1 U5504 ( .A1(n4445), .A2(n6570), .ZN(n5413) );
  OAI21_X1 U5505 ( .B1(n3346), .B2(n4432), .A(n5413), .ZN(n4433) );
  AND2_X2 U5506 ( .A1(n5412), .A2(n4433), .ZN(n6110) );
  INV_X1 U5507 ( .A(n4434), .ZN(n4435) );
  NAND2_X1 U5508 ( .A1(n4435), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U5509 ( .A1(EBX_REG_30__SCAN_IN), .A2(n6110), .B1(n4437), .B2(n6096), .ZN(n4438) );
  NAND2_X1 U5510 ( .A1(n4443), .A2(n4537), .ZN(n4444) );
  OAI21_X1 U5511 ( .B1(n4547), .B2(n5092), .A(n4444), .ZN(n5986) );
  OR2_X1 U5512 ( .A1(n4445), .A2(n5115), .ZN(n4455) );
  AOI21_X1 U5513 ( .B1(n4455), .B2(n6598), .A(READY_N), .ZN(n6699) );
  NOR2_X1 U5514 ( .A1(n5986), .A2(n6699), .ZN(n6559) );
  NOR2_X1 U5515 ( .A1(n6559), .A2(n6581), .ZN(n5993) );
  INV_X1 U5516 ( .A(MORE_REG_SCAN_IN), .ZN(n4453) );
  AND2_X1 U5517 ( .A1(n4446), .A2(n4537), .ZN(n4451) );
  OR2_X1 U5518 ( .A1(n4448), .A2(n4447), .ZN(n4450) );
  NAND2_X1 U5519 ( .A1(n4547), .A2(n4571), .ZN(n4449) );
  OAI211_X1 U5520 ( .C1(n4547), .C2(n4451), .A(n4450), .B(n4449), .ZN(n6558)
         );
  NAND2_X1 U5521 ( .A1(n5993), .A2(n6558), .ZN(n4452) );
  OAI21_X1 U5522 ( .B1(n5993), .B2(n4453), .A(n4452), .ZN(U3471) );
  OR2_X1 U5523 ( .A1(n6694), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5988) );
  INV_X1 U5524 ( .A(n5988), .ZN(n5074) );
  OAI21_X1 U5525 ( .B1(n5074), .B2(READREQUEST_REG_SCAN_IN), .A(n6693), .ZN(
        n4454) );
  OAI21_X1 U5526 ( .B1(n6693), .B2(n4455), .A(n4454), .ZN(U3474) );
  NAND2_X1 U5527 ( .A1(n4530), .A2(n4571), .ZN(n4548) );
  INV_X1 U5528 ( .A(n4697), .ZN(n5395) );
  NAND3_X1 U5529 ( .A1(n3317), .A2(n5395), .A3(n4456), .ZN(n4685) );
  INV_X1 U5530 ( .A(n4685), .ZN(n4458) );
  NAND4_X1 U5531 ( .A1(n4467), .A2(n4458), .A3(n3289), .A4(n4457), .ZN(n4459)
         );
  NAND2_X1 U5532 ( .A1(n4548), .A2(n4459), .ZN(n4460) );
  NOR2_X1 U5533 ( .A1(n4463), .A2(n4462), .ZN(n4464) );
  OR2_X1 U5534 ( .A1(n4461), .A2(n4464), .ZN(n6094) );
  INV_X1 U5535 ( .A(n4465), .ZN(n4468) );
  OAI21_X1 U5536 ( .B1(n4468), .B2(n4467), .A(n4466), .ZN(n4678) );
  AOI22_X1 U5537 ( .A1(n6124), .A2(n4678), .B1(n5454), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4469) );
  OAI21_X1 U5538 ( .B1(n5456), .B2(n6094), .A(n4469), .ZN(U2858) );
  XNOR2_X1 U5539 ( .A(n4470), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4492)
         );
  AOI21_X1 U5540 ( .B1(n4472), .B2(n4528), .A(n4471), .ZN(n6106) );
  INV_X1 U5541 ( .A(REIP_REG_0__SCAN_IN), .ZN(n4473) );
  NOR2_X1 U5542 ( .A1(n6292), .A2(n4473), .ZN(n4488) );
  AOI21_X1 U5543 ( .B1(n5611), .B2(n6106), .A(n4488), .ZN(n4475) );
  OAI21_X1 U5544 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6288), .A(n6239), 
        .ZN(n4674) );
  OR2_X1 U5545 ( .A1(n6310), .A2(n5753), .ZN(n5746) );
  OAI22_X1 U5546 ( .A1(n5749), .A2(n4674), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5746), .ZN(n4474) );
  OAI211_X1 U5547 ( .C1(n4492), .C2(n5745), .A(n4475), .B(n4474), .ZN(U3018)
         );
  INV_X1 U5548 ( .A(n6571), .ZN(n4476) );
  NAND2_X1 U5549 ( .A1(n4477), .A2(n6543), .ZN(n4478) );
  NAND2_X1 U5550 ( .A1(n6193), .A2(n4478), .ZN(n4480) );
  NAND2_X1 U5551 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), 
        .ZN(n4613) );
  NOR2_X1 U5552 ( .A1(n4613), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6157) );
  INV_X1 U5553 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n6945) );
  INV_X1 U5554 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6853) );
  INV_X1 U5555 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6858) );
  OAI222_X1 U5556 ( .A1(n6146), .A2(n6945), .B1(n4671), .B2(n6853), .C1(n6858), 
        .C2(n6696), .ZN(U2896) );
  NAND2_X1 U5557 ( .A1(n4481), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4483) );
  NAND2_X1 U5558 ( .A1(n4483), .A2(n4482), .ZN(n4485) );
  NAND2_X1 U5559 ( .A1(n4485), .A2(n4484), .ZN(n6115) );
  INV_X1 U5560 ( .A(n6106), .ZN(n4486) );
  OAI222_X1 U5561 ( .A1(n6115), .A2(n5456), .B1(n6827), .B2(n7016), .C1(n7014), 
        .C2(n4486), .ZN(U2859) );
  OAI21_X1 U5562 ( .B1(n6218), .B2(n4487), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4491) );
  INV_X1 U5563 ( .A(n6115), .ZN(n4489) );
  AOI21_X1 U5564 ( .B1(n4489), .B2(n6223), .A(n4488), .ZN(n4490) );
  OAI211_X1 U5565 ( .C1(n4492), .C2(n6213), .A(n4491), .B(n4490), .ZN(U2986)
         );
  INV_X1 U5566 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4786) );
  NAND2_X1 U5567 ( .A1(n5804), .A2(n4495), .ZN(n4494) );
  AND2_X2 U5568 ( .A1(n4494), .A2(n6193), .ZN(n6191) );
  NAND2_X1 U5569 ( .A1(n6191), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4498) );
  AND2_X1 U5570 ( .A1(n4496), .A2(n4495), .ZN(n4497) );
  NAND2_X1 U5571 ( .A1(n6190), .A2(DATAI_6_), .ZN(n4508) );
  OAI211_X1 U5572 ( .C1(n6193), .C2(n4786), .A(n4498), .B(n4508), .ZN(U2945)
         );
  INV_X1 U5573 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4500) );
  NAND2_X1 U5574 ( .A1(n6191), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4499) );
  NAND2_X1 U5575 ( .A1(n6190), .A2(DATAI_4_), .ZN(n4512) );
  OAI211_X1 U5576 ( .C1(n6193), .C2(n4500), .A(n4499), .B(n4512), .ZN(U2928)
         );
  INV_X1 U5577 ( .A(EAX_REG_1__SCAN_IN), .ZN(n4502) );
  NAND2_X1 U5578 ( .A1(n6191), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4501) );
  INV_X1 U5579 ( .A(DATAI_1_), .ZN(n4701) );
  OR2_X1 U5580 ( .A1(n6174), .A2(n4701), .ZN(n4725) );
  OAI211_X1 U5581 ( .C1(n6193), .C2(n4502), .A(n4501), .B(n4725), .ZN(U2940)
         );
  INV_X1 U5582 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4504) );
  NAND2_X1 U5583 ( .A1(n6191), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4503) );
  INV_X1 U5584 ( .A(DATAI_10_), .ZN(n5087) );
  OR2_X1 U5585 ( .A1(n6174), .A2(n5087), .ZN(n4722) );
  OAI211_X1 U5586 ( .C1(n6193), .C2(n4504), .A(n4503), .B(n4722), .ZN(U2934)
         );
  INV_X1 U5587 ( .A(EAX_REG_19__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U5588 ( .A1(n6191), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4505) );
  INV_X1 U5589 ( .A(DATAI_3_), .ZN(n4715) );
  OR2_X1 U5590 ( .A1(n6174), .A2(n4715), .ZN(n4515) );
  OAI211_X1 U5591 ( .C1(n6193), .C2(n6933), .A(n4505), .B(n4515), .ZN(U2927)
         );
  INV_X1 U5592 ( .A(EAX_REG_0__SCAN_IN), .ZN(n4507) );
  NAND2_X1 U5593 ( .A1(n6191), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5594 ( .A1(n6190), .A2(DATAI_0_), .ZN(n4716) );
  OAI211_X1 U5595 ( .C1(n6193), .C2(n4507), .A(n4506), .B(n4716), .ZN(U2939)
         );
  INV_X1 U5596 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4510) );
  NAND2_X1 U5597 ( .A1(n6191), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4509) );
  OAI211_X1 U5598 ( .C1(n6193), .C2(n4510), .A(n4509), .B(n4508), .ZN(U2930)
         );
  INV_X1 U5599 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U5600 ( .A1(n6191), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4511) );
  NAND2_X1 U5601 ( .A1(n6190), .A2(DATAI_7_), .ZN(n4560) );
  OAI211_X1 U5602 ( .C1(n6193), .C2(n4669), .A(n4511), .B(n4560), .ZN(U2931)
         );
  INV_X1 U5603 ( .A(EAX_REG_4__SCAN_IN), .ZN(n4514) );
  NAND2_X1 U5604 ( .A1(n6191), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4513) );
  OAI211_X1 U5605 ( .C1(n6193), .C2(n4514), .A(n4513), .B(n4512), .ZN(U2943)
         );
  INV_X1 U5606 ( .A(EAX_REG_3__SCAN_IN), .ZN(n4517) );
  NAND2_X1 U5607 ( .A1(n6191), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4516) );
  OAI211_X1 U5608 ( .C1(n6193), .C2(n4517), .A(n4516), .B(n4515), .ZN(U2942)
         );
  INV_X1 U5609 ( .A(n4519), .ZN(n4864) );
  NAND2_X1 U5610 ( .A1(n4686), .A2(n4336), .ZN(n4520) );
  NOR2_X1 U5611 ( .A1(n4540), .A2(n4520), .ZN(n4521) );
  NAND3_X1 U5612 ( .A1(n4522), .A2(n4521), .A3(n4605), .ZN(n6542) );
  INV_X1 U5613 ( .A(n6542), .ZN(n4527) );
  AND2_X1 U5614 ( .A1(n6543), .A2(n3180), .ZN(n4585) );
  INV_X1 U5615 ( .A(n4585), .ZN(n4526) );
  INV_X1 U5616 ( .A(n4523), .ZN(n5387) );
  INV_X1 U5617 ( .A(n4524), .ZN(n4602) );
  NAND3_X1 U5618 ( .A1(n6541), .A2(n5387), .A3(n4602), .ZN(n4525) );
  OAI211_X1 U5619 ( .C1(n4864), .C2(n4527), .A(n4526), .B(n4525), .ZN(n6546)
         );
  INV_X1 U5620 ( .A(n6670), .ZN(n5981) );
  NOR2_X1 U5621 ( .A1(n4616), .A2(n4528), .ZN(n5380) );
  INV_X1 U5622 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5603) );
  AOI22_X1 U5623 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5603), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4529), .ZN(n5381) );
  AOI222_X1 U5624 ( .A1(n6546), .A2(n5981), .B1(n5380), .B2(n5381), .C1(n4531), 
        .C2(n5386), .ZN(n4552) );
  NOR2_X1 U5625 ( .A1(n4532), .A2(n3355), .ZN(n4570) );
  NAND2_X1 U5626 ( .A1(n4547), .A2(n4570), .ZN(n4536) );
  INV_X1 U5627 ( .A(n4533), .ZN(n4534) );
  OR2_X1 U5628 ( .A1(n4605), .A2(n4534), .ZN(n4535) );
  NAND2_X1 U5629 ( .A1(n4536), .A2(n4535), .ZN(n4688) );
  INV_X1 U5630 ( .A(n4688), .ZN(n4550) );
  NAND2_X1 U5631 ( .A1(n4537), .A2(n6598), .ZN(n4539) );
  OAI211_X1 U5632 ( .C1(n4540), .C2(n6543), .A(n4539), .B(n4538), .ZN(n4541)
         );
  INV_X1 U5633 ( .A(n4541), .ZN(n4546) );
  OAI21_X1 U5634 ( .B1(n4544), .B2(n4543), .A(n4542), .ZN(n4545) );
  AOI21_X1 U5635 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(n4549) );
  OR2_X1 U5636 ( .A1(n6576), .A2(n4613), .ZN(n6660) );
  INV_X1 U5637 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5992) );
  OAI22_X1 U5638 ( .A1(n6544), .A2(n6581), .B1(n6660), .B2(n5992), .ZN(n5983)
         );
  AOI21_X1 U5639 ( .B1(n6576), .B2(STATE2_REG_3__SCAN_IN), .A(n5983), .ZN(
        n6664) );
  INV_X1 U5640 ( .A(n5386), .ZN(n6577) );
  NOR2_X1 U5641 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6577), .ZN(n6663)
         );
  OAI21_X1 U5642 ( .B1(n6663), .B2(n6664), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4551) );
  OAI21_X1 U5643 ( .B1(n4552), .B2(n6664), .A(n4551), .ZN(U3460) );
  INV_X1 U5644 ( .A(n6191), .ZN(n6189) );
  INV_X1 U5645 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4555) );
  INV_X1 U5646 ( .A(DATAI_2_), .ZN(n4553) );
  NOR2_X1 U5647 ( .A1(n6174), .A2(n4553), .ZN(n4556) );
  AOI21_X1 U5648 ( .B1(n6187), .B2(EAX_REG_18__SCAN_IN), .A(n4556), .ZN(n4554)
         );
  OAI21_X1 U5649 ( .B1(n6189), .B2(n4555), .A(n4554), .ZN(U2926) );
  INV_X1 U5650 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n4558) );
  AOI21_X1 U5651 ( .B1(n6187), .B2(EAX_REG_2__SCAN_IN), .A(n4556), .ZN(n4557)
         );
  OAI21_X1 U5652 ( .B1(n6189), .B2(n4558), .A(n4557), .ZN(U2941) );
  INV_X1 U5653 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U5654 ( .A1(n6187), .A2(EAX_REG_7__SCAN_IN), .ZN(n4559) );
  OAI211_X1 U5655 ( .C1(n6189), .C2(n4561), .A(n4560), .B(n4559), .ZN(U2946)
         );
  INV_X1 U5656 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4563) );
  AOI22_X1 U5657 ( .A1(n6141), .A2(EAX_REG_19__SCAN_IN), .B1(n6567), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4562) );
  OAI21_X1 U5658 ( .B1(n6146), .B2(n4563), .A(n4562), .ZN(U2904) );
  INV_X1 U5659 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5660 ( .A1(n6141), .A2(EAX_REG_21__SCAN_IN), .B1(n6567), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U5661 ( .B1(n6146), .B2(n4565), .A(n4564), .ZN(U2902) );
  NAND2_X1 U5662 ( .A1(n4523), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5663 ( .A1(n4567), .A2(n4582), .ZN(n4568) );
  NAND2_X1 U5664 ( .A1(n4569), .A2(n4568), .ZN(n5763) );
  OR2_X1 U5665 ( .A1(n4571), .A2(n4570), .ZN(n4584) );
  NOR2_X1 U5666 ( .A1(n4523), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4574)
         );
  AND2_X1 U5667 ( .A1(n4584), .A2(n4574), .ZN(n4592) );
  INV_X1 U5668 ( .A(n4592), .ZN(n4573) );
  NAND2_X1 U5669 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4575) );
  NAND2_X1 U5670 ( .A1(n6543), .A2(n4575), .ZN(n4572) );
  AND2_X1 U5671 ( .A1(n4573), .A2(n4572), .ZN(n4579) );
  INV_X1 U5672 ( .A(n4574), .ZN(n4577) );
  INV_X1 U5673 ( .A(n4575), .ZN(n4576) );
  AOI22_X1 U5674 ( .A1(n4584), .A2(n4577), .B1(n6543), .B2(n4576), .ZN(n4578)
         );
  MUX2_X1 U5675 ( .A(n4579), .B(n4578), .S(n4582), .Z(n4580) );
  OAI21_X1 U5676 ( .B1(n5763), .B2(n4583), .A(n4580), .ZN(n4581) );
  AOI21_X1 U5677 ( .B1(n6677), .B2(n6542), .A(n4581), .ZN(n5764) );
  MUX2_X1 U5678 ( .A(n5764), .B(n4582), .S(n6544), .Z(n6551) );
  INV_X1 U5679 ( .A(n6551), .ZN(n4597) );
  INV_X1 U5680 ( .A(n4583), .ZN(n4587) );
  MUX2_X1 U5681 ( .A(n4584), .B(n4587), .S(n5387), .Z(n4586) );
  NOR2_X1 U5682 ( .A1(n4586), .A2(n4585), .ZN(n4589) );
  AOI22_X1 U5683 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n6543), .B1(n4587), .B2(n4523), .ZN(n4588) );
  MUX2_X1 U5684 ( .A(n4589), .B(n4588), .S(n5388), .Z(n4594) );
  AOI21_X1 U5685 ( .B1(n4591), .B2(n6542), .A(n4592), .ZN(n4593) );
  NAND2_X1 U5686 ( .A1(n4594), .A2(n4593), .ZN(n5385) );
  OR2_X1 U5687 ( .A1(n6544), .A2(n5385), .ZN(n4596) );
  NAND2_X1 U5688 ( .A1(n6544), .A2(n5388), .ZN(n4595) );
  NAND3_X1 U5689 ( .A1(n4597), .A2(n6550), .A3(n4616), .ZN(n4601) );
  NAND2_X1 U5690 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5992), .ZN(n4608) );
  INV_X1 U5691 ( .A(n4608), .ZN(n4599) );
  NAND2_X1 U5692 ( .A1(n4598), .A2(n4599), .ZN(n4600) );
  NAND2_X1 U5693 ( .A1(n4601), .A2(n4600), .ZN(n6564) );
  NAND2_X1 U5694 ( .A1(n6564), .A2(n4602), .ZN(n4615) );
  NAND2_X1 U5695 ( .A1(n6544), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4607) );
  INV_X1 U5696 ( .A(n5131), .ZN(n6375) );
  OR2_X1 U5697 ( .A1(n4603), .A2(n6375), .ZN(n4604) );
  XNOR2_X1 U5698 ( .A(n4604), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6070)
         );
  INV_X1 U5699 ( .A(n4605), .ZN(n5982) );
  NAND2_X1 U5700 ( .A1(n6070), .A2(n5982), .ZN(n4606) );
  NAND2_X1 U5701 ( .A1(n4607), .A2(n4606), .ZN(n4610) );
  NOR2_X1 U5702 ( .A1(n4608), .A2(n6802), .ZN(n4609) );
  AOI21_X1 U5703 ( .B1(n4610), .B2(n4616), .A(n4609), .ZN(n6562) );
  AND2_X1 U5704 ( .A1(n6562), .A2(n5992), .ZN(n4611) );
  AOI21_X1 U5705 ( .B1(n4615), .B2(n4611), .A(n6660), .ZN(n4612) );
  OR2_X1 U5706 ( .A1(n4612), .A2(n5038), .ZN(n6679) );
  INV_X1 U5707 ( .A(n4613), .ZN(n4614) );
  AND3_X1 U5708 ( .A1(n4615), .A2(n6562), .A3(n4614), .ZN(n6575) );
  INV_X1 U5709 ( .A(n3690), .ZN(n6330) );
  NOR2_X1 U5710 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n4616), .ZN(n4639) );
  OAI22_X1 U5711 ( .A1(n5043), .A2(n6694), .B1(n6330), .B2(n4639), .ZN(n4617)
         );
  OAI21_X1 U5712 ( .B1(n6575), .B2(n4617), .A(n6679), .ZN(n4618) );
  OAI21_X1 U5713 ( .B1(n6679), .B2(n6372), .A(n4618), .ZN(U3465) );
  INV_X1 U5714 ( .A(n4619), .ZN(n4621) );
  AOI21_X1 U5715 ( .B1(n4621), .B2(n5118), .A(n4620), .ZN(n4622) );
  OR2_X1 U5716 ( .A1(n4622), .A2(n4634), .ZN(n6082) );
  INV_X1 U5717 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4628) );
  NAND2_X1 U5718 ( .A1(n4623), .A2(n4624), .ZN(n4696) );
  INV_X1 U5719 ( .A(n4696), .ZN(n4627) );
  OAI21_X1 U5720 ( .B1(n4627), .B2(n3706), .A(n4626), .ZN(n6086) );
  OAI222_X1 U5721 ( .A1(n6082), .A2(n7014), .B1(n4628), .B2(n7016), .C1(n6086), 
        .C2(n5456), .ZN(U2856) );
  AND2_X1 U5722 ( .A1(n4626), .A2(n4630), .ZN(n4631) );
  OR2_X1 U5723 ( .A1(n4629), .A2(n4631), .ZN(n6212) );
  OR2_X1 U5724 ( .A1(n4634), .A2(n4633), .ZN(n4635) );
  NAND2_X1 U5725 ( .A1(n4683), .A2(n4635), .ZN(n6293) );
  INV_X1 U5726 ( .A(n6293), .ZN(n6071) );
  AOI22_X1 U5727 ( .A1(n6124), .A2(n6071), .B1(n5454), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4636) );
  OAI21_X1 U5728 ( .B1(n6212), .B2(n5456), .A(n4636), .ZN(U2855) );
  INV_X1 U5729 ( .A(n4993), .ZN(n4638) );
  AOI21_X1 U5730 ( .B1(n4638), .B2(n5991), .A(n6694), .ZN(n4640) );
  NAND2_X1 U5731 ( .A1(n4993), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6410) );
  INV_X1 U5732 ( .A(n4639), .ZN(n6678) );
  AOI22_X1 U5733 ( .A1(n4640), .A2(n6410), .B1(n4519), .B2(n6678), .ZN(n4642)
         );
  NAND2_X1 U5734 ( .A1(n6682), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5735 ( .B1(n6682), .B2(n4642), .A(n4641), .ZN(U3464) );
  XNOR2_X1 U5736 ( .A(n4990), .B(n6410), .ZN(n4644) );
  INV_X1 U5737 ( .A(n6694), .ZN(n6674) );
  AOI22_X1 U5738 ( .A1(n4644), .A2(n6674), .B1(n6678), .B2(n4591), .ZN(n4646)
         );
  NAND2_X1 U5739 ( .A1(n6682), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4645) );
  OAI21_X1 U5740 ( .B1(n6682), .B2(n4646), .A(n4645), .ZN(U3463) );
  XNOR2_X1 U5741 ( .A(n4648), .B(n4649), .ZN(n4680) );
  INV_X1 U5742 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n6099) );
  INV_X1 U5743 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5117) );
  OAI22_X1 U5744 ( .A1(n5955), .A2(n6099), .B1(n6292), .B2(n5117), .ZN(n4651)
         );
  NOR2_X1 U5745 ( .A1(n6094), .A2(n5564), .ZN(n4650) );
  AOI211_X1 U5746 ( .C1(n6196), .C2(n6099), .A(n4651), .B(n4650), .ZN(n4652)
         );
  OAI21_X1 U5747 ( .B1(n4680), .B2(n6213), .A(n4652), .ZN(U2985) );
  NAND2_X1 U5748 ( .A1(n6317), .A2(REIP_REG_3__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U5749 ( .B1(n5955), .B2(n4653), .A(n6301), .ZN(n4654) );
  AOI21_X1 U5750 ( .B1(n6196), .B2(n6088), .A(n4654), .ZN(n4660) );
  OR2_X1 U5751 ( .A1(n4656), .A2(n4655), .ZN(n6302) );
  NAND3_X1 U5752 ( .A1(n6302), .A2(n4658), .A3(n6224), .ZN(n4659) );
  OAI211_X1 U5753 ( .C1(n6086), .C2(n5564), .A(n4660), .B(n4659), .ZN(U2983)
         );
  INV_X1 U5754 ( .A(EAX_REG_30__SCAN_IN), .ZN(n6844) );
  AOI22_X1 U5755 ( .A1(n6567), .A2(UWORD_REG_14__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4661) );
  OAI21_X1 U5756 ( .B1(n6844), .B2(n4671), .A(n4661), .ZN(U2893) );
  INV_X1 U5757 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4663) );
  AOI22_X1 U5758 ( .A1(n6157), .A2(UWORD_REG_12__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4662) );
  OAI21_X1 U5759 ( .B1(n4663), .B2(n4671), .A(n4662), .ZN(U2895) );
  AOI22_X1 U5760 ( .A1(n6157), .A2(UWORD_REG_8__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4664) );
  OAI21_X1 U5761 ( .B1(n4026), .B2(n4671), .A(n4664), .ZN(U2899) );
  INV_X1 U5762 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4666) );
  AOI22_X1 U5763 ( .A1(n6157), .A2(UWORD_REG_13__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4665) );
  OAI21_X1 U5764 ( .B1(n4666), .B2(n4671), .A(n4665), .ZN(U2894) );
  AOI22_X1 U5765 ( .A1(n6157), .A2(UWORD_REG_4__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4667) );
  OAI21_X1 U5766 ( .B1(n4500), .B2(n4671), .A(n4667), .ZN(U2903) );
  AOI22_X1 U5767 ( .A1(n6157), .A2(UWORD_REG_7__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4668) );
  OAI21_X1 U5768 ( .B1(n4669), .B2(n4671), .A(n4668), .ZN(U2900) );
  INV_X1 U5769 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4672) );
  AOI22_X1 U5770 ( .A1(n6567), .A2(UWORD_REG_0__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4670) );
  OAI21_X1 U5771 ( .B1(n4672), .B2(n4671), .A(n4670), .ZN(U2907) );
  NOR2_X1 U5772 ( .A1(n6292), .A2(n5117), .ZN(n4677) );
  NOR2_X1 U5773 ( .A1(n5599), .A2(n4673), .ZN(n4675) );
  MUX2_X1 U5774 ( .A(n4675), .B(n4674), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4676) );
  AOI211_X1 U5775 ( .C1(n5611), .C2(n4678), .A(n4677), .B(n4676), .ZN(n4679)
         );
  OAI21_X1 U5776 ( .B1(n4680), .B2(n5745), .A(n4679), .ZN(U3017) );
  OAI21_X1 U5777 ( .B1(n4629), .B2(n4682), .A(n4681), .ZN(n5102) );
  INV_X1 U5778 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6959) );
  OAI21_X1 U5779 ( .B1(n4248), .B2(n3178), .A(n4684), .ZN(n6280) );
  OAI222_X1 U5780 ( .A1(n5102), .A2(n5456), .B1(n7016), .B2(n6959), .C1(n6280), 
        .C2(n7014), .ZN(U2854) );
  NOR2_X1 U5781 ( .A1(n4686), .A2(n4685), .ZN(n4687) );
  NAND2_X1 U5782 ( .A1(n3316), .A2(n4697), .ZN(n4691) );
  INV_X1 U5783 ( .A(n4692), .ZN(n4693) );
  OR3_X1 U5784 ( .A1(n4461), .A2(n4694), .A3(n4693), .ZN(n4695) );
  NAND2_X1 U5785 ( .A1(n4696), .A2(n4695), .ZN(n6123) );
  AND2_X1 U5786 ( .A1(n5396), .A2(n3352), .ZN(n6130) );
  AND2_X1 U5787 ( .A1(n3289), .A2(n4697), .ZN(n4698) );
  AOI22_X1 U5788 ( .A1(n5363), .A2(DATAI_2_), .B1(EAX_REG_2__SCAN_IN), .B2(
        n6133), .ZN(n4699) );
  OAI21_X1 U5789 ( .B1(n5916), .B2(n6123), .A(n4699), .ZN(U2889) );
  INV_X1 U5790 ( .A(DATAI_5_), .ZN(n6787) );
  INV_X1 U5791 ( .A(EAX_REG_5__SCAN_IN), .ZN(n4700) );
  OAI222_X1 U5792 ( .A1(n5102), .A2(n5916), .B1(n5088), .B2(n6787), .C1(n5396), 
        .C2(n4700), .ZN(U2886) );
  INV_X1 U5793 ( .A(DATAI_4_), .ZN(n6928) );
  OAI222_X1 U5794 ( .A1(n6212), .A2(n5916), .B1(n5088), .B2(n6928), .C1(n5396), 
        .C2(n4514), .ZN(U2887) );
  OAI222_X1 U5795 ( .A1(n6094), .A2(n5916), .B1(n5088), .B2(n4701), .C1(n5396), 
        .C2(n4502), .ZN(U2890) );
  OAI21_X1 U5796 ( .B1(n6323), .B2(n6410), .A(n6674), .ZN(n4708) );
  INV_X1 U5797 ( .A(n4824), .ZN(n4702) );
  NAND2_X1 U5798 ( .A1(n5283), .A2(n3690), .ZN(n4704) );
  INV_X1 U5799 ( .A(n6328), .ZN(n4703) );
  NAND2_X1 U5800 ( .A1(n4703), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5801 ( .A1(n4704), .A2(n4710), .ZN(n4706) );
  NAND2_X1 U5802 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4822), .ZN(n5281) );
  NAND2_X1 U5803 ( .A1(n6694), .A2(n5281), .ZN(n4705) );
  OAI211_X1 U5804 ( .C1(n4708), .C2(n4706), .A(n6414), .B(n4705), .ZN(n6536)
         );
  INV_X1 U5805 ( .A(n6536), .ZN(n4793) );
  INV_X1 U5806 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U5807 ( .A1(DATAI_2_), .A2(n5038), .ZN(n6426) );
  INV_X1 U5808 ( .A(n4706), .ZN(n4707) );
  OAI22_X1 U5809 ( .A1(n4708), .A2(n4707), .B1(n5281), .B2(n6334), .ZN(n6534)
         );
  INV_X1 U5810 ( .A(n4710), .ZN(n6532) );
  AOI22_X1 U5811 ( .A1(n6468), .A2(n6534), .B1(n6467), .B2(n6532), .ZN(n4713)
         );
  INV_X1 U5812 ( .A(DATAI_18_), .ZN(n4711) );
  NOR2_X1 U5813 ( .A1(n6211), .A2(n4711), .ZN(n6469) );
  NAND2_X1 U5814 ( .A1(n4993), .A2(n4994), .ZN(n6409) );
  INV_X1 U5815 ( .A(n6539), .ZN(n4789) );
  NAND2_X1 U5816 ( .A1(n4993), .A2(n5043), .ZN(n6366) );
  NOR2_X2 U5817 ( .A1(n6323), .A2(n6366), .ZN(n6530) );
  NAND2_X1 U5818 ( .A1(n6223), .A2(DATAI_26_), .ZN(n6472) );
  INV_X1 U5819 ( .A(n6472), .ZN(n6423) );
  AOI22_X1 U5820 ( .A1(n6469), .A2(n4789), .B1(n6530), .B2(n6423), .ZN(n4712)
         );
  OAI211_X1 U5821 ( .C1(n4793), .C2(n4714), .A(n4713), .B(n4712), .ZN(U3110)
         );
  OAI222_X1 U5822 ( .A1(n6086), .A2(n5916), .B1(n5088), .B2(n4715), .C1(n5396), 
        .C2(n4517), .ZN(U2888) );
  INV_X1 U5823 ( .A(DATAI_0_), .ZN(n6996) );
  OAI222_X1 U5824 ( .A1(n6115), .A2(n5916), .B1(n5088), .B2(n6996), .C1(n5396), 
        .C2(n4507), .ZN(U2891) );
  NAND2_X1 U5825 ( .A1(n6191), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4717) );
  OAI211_X1 U5826 ( .C1(n6193), .C2(n4672), .A(n4717), .B(n4716), .ZN(U2924)
         );
  NAND2_X1 U5827 ( .A1(n6191), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U5828 ( .A1(n6190), .A2(DATAI_5_), .ZN(n4719) );
  OAI211_X1 U5829 ( .C1(n6193), .C2(n4700), .A(n4718), .B(n4719), .ZN(U2944)
         );
  INV_X1 U5830 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4721) );
  NAND2_X1 U5831 ( .A1(n6191), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4720) );
  OAI211_X1 U5832 ( .C1(n6193), .C2(n4721), .A(n4720), .B(n4719), .ZN(U2929)
         );
  INV_X1 U5833 ( .A(EAX_REG_10__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U5834 ( .A1(n6191), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4723) );
  OAI211_X1 U5835 ( .C1(n6193), .C2(n4724), .A(n4723), .B(n4722), .ZN(U2949)
         );
  INV_X1 U5836 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4727) );
  NAND2_X1 U5837 ( .A1(n6191), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4726) );
  OAI211_X1 U5838 ( .C1(n6193), .C2(n4727), .A(n4726), .B(n4725), .ZN(U2925)
         );
  XNOR2_X1 U5839 ( .A(n4729), .B(n4728), .ZN(n5083) );
  AOI21_X1 U5840 ( .B1(n4730), .B2(n4782), .A(n4776), .ZN(n6267) );
  AOI22_X1 U5841 ( .A1(n6124), .A2(n6267), .B1(n5454), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n4731) );
  OAI21_X1 U5842 ( .B1(n5083), .B2(n5456), .A(n4731), .ZN(U2852) );
  INV_X1 U5843 ( .A(n5102), .ZN(n4737) );
  INV_X1 U5844 ( .A(n5095), .ZN(n4735) );
  AOI22_X1 U5845 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6317), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4734) );
  OAI21_X1 U5846 ( .B1(n6228), .B2(n4735), .A(n4734), .ZN(n4736) );
  AOI21_X1 U5847 ( .B1(n4737), .B2(n6223), .A(n4736), .ZN(n4738) );
  OAI21_X1 U5848 ( .B1(n6213), .B2(n6279), .A(n4738), .ZN(U2981) );
  AND2_X1 U5849 ( .A1(n4993), .A2(n4739), .ZN(n4740) );
  NAND2_X1 U5850 ( .A1(n4990), .A2(n4740), .ZN(n4747) );
  INV_X1 U5851 ( .A(n4747), .ZN(n4741) );
  OR2_X1 U5852 ( .A1(n6694), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6374) );
  OAI21_X1 U5853 ( .B1(n4741), .B2(n5564), .A(n6374), .ZN(n4744) );
  AND2_X1 U5854 ( .A1(n3690), .A2(n6677), .ZN(n4866) );
  NAND2_X1 U5855 ( .A1(n4866), .A2(n6376), .ZN(n4742) );
  NAND2_X1 U5856 ( .A1(n4742), .A2(n4862), .ZN(n4748) );
  INV_X1 U5857 ( .A(n4748), .ZN(n4743) );
  NAND2_X1 U5858 ( .A1(n4744), .A2(n4743), .ZN(n4745) );
  OAI211_X1 U5859 ( .C1(n4932), .C2(n6674), .A(n4745), .B(n6414), .ZN(n4860)
         );
  NAND2_X1 U5860 ( .A1(n6223), .A2(DATAI_31_), .ZN(n6499) );
  INV_X1 U5861 ( .A(DATAI_23_), .ZN(n4746) );
  NOR2_X1 U5862 ( .A1(n5564), .A2(n4746), .ZN(n6493) );
  INV_X1 U5863 ( .A(n6493), .ZN(n6540) );
  OAI22_X1 U5864 ( .A1(n4930), .A2(n6499), .B1(n6540), .B2(n5067), .ZN(n4750)
         );
  NAND2_X1 U5865 ( .A1(DATAI_7_), .A2(n5038), .ZN(n6445) );
  AOI22_X1 U5866 ( .A1(n4748), .A2(n6674), .B1(n4932), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4857) );
  NOR2_X1 U5867 ( .A1(n6445), .A2(n4857), .ZN(n4749) );
  AOI211_X1 U5868 ( .C1(INSTQUEUE_REG_15__7__SCAN_IN), .C2(n4860), .A(n4750), 
        .B(n4749), .ZN(n4751) );
  OAI21_X1 U5869 ( .B1(n4862), .B2(n5138), .A(n4751), .ZN(U3147) );
  INV_X1 U5870 ( .A(DATAI_25_), .ZN(n6951) );
  NOR2_X1 U5871 ( .A1(n6211), .A2(n6951), .ZN(n6506) );
  INV_X1 U5872 ( .A(n6506), .ZN(n6466) );
  INV_X1 U5873 ( .A(DATAI_17_), .ZN(n4753) );
  NOR2_X1 U5874 ( .A1(n6211), .A2(n4753), .ZN(n6463) );
  INV_X1 U5875 ( .A(n6463), .ZN(n6511) );
  OAI22_X1 U5876 ( .A1(n4930), .A2(n6466), .B1(n6511), .B2(n5067), .ZN(n4755)
         );
  NAND2_X1 U5877 ( .A1(DATAI_1_), .A2(n5038), .ZN(n6422) );
  NOR2_X1 U5878 ( .A1(n6422), .A2(n4857), .ZN(n4754) );
  AOI211_X1 U5879 ( .C1(INSTQUEUE_REG_15__1__SCAN_IN), .C2(n4860), .A(n4755), 
        .B(n4754), .ZN(n4756) );
  OAI21_X1 U5880 ( .B1(n4862), .B2(n5158), .A(n4756), .ZN(U3141) );
  INV_X1 U5881 ( .A(DATAI_24_), .ZN(n4757) );
  NOR2_X1 U5882 ( .A1(n6211), .A2(n4757), .ZN(n6500) );
  INV_X1 U5883 ( .A(n6500), .ZN(n6462) );
  INV_X1 U5884 ( .A(DATAI_16_), .ZN(n4758) );
  NOR2_X1 U5885 ( .A1(n6211), .A2(n4758), .ZN(n6459) );
  INV_X1 U5886 ( .A(n6459), .ZN(n6505) );
  OAI22_X1 U5887 ( .A1(n4930), .A2(n6462), .B1(n6505), .B2(n5067), .ZN(n4760)
         );
  NAND2_X1 U5888 ( .A1(DATAI_0_), .A2(n5038), .ZN(n6419) );
  NOR2_X1 U5889 ( .A1(n6419), .A2(n4857), .ZN(n4759) );
  AOI211_X1 U5890 ( .C1(INSTQUEUE_REG_15__0__SCAN_IN), .C2(n4860), .A(n4760), 
        .B(n4759), .ZN(n4761) );
  OAI21_X1 U5891 ( .B1(n4862), .B2(n5170), .A(n4761), .ZN(U3140) );
  INV_X1 U5892 ( .A(n6469), .ZN(n6388) );
  OAI22_X1 U5893 ( .A1(n4930), .A2(n6472), .B1(n6388), .B2(n5067), .ZN(n4763)
         );
  NOR2_X1 U5894 ( .A1(n6426), .A2(n4857), .ZN(n4762) );
  AOI211_X1 U5895 ( .C1(INSTQUEUE_REG_15__2__SCAN_IN), .C2(n4860), .A(n4763), 
        .B(n4762), .ZN(n4764) );
  OAI21_X1 U5896 ( .B1(n4862), .B2(n5142), .A(n4764), .ZN(U3142) );
  INV_X1 U5897 ( .A(n3313), .ZN(n4765) );
  INV_X1 U5898 ( .A(DATAI_27_), .ZN(n4766) );
  NOR2_X1 U5899 ( .A1(n5564), .A2(n4766), .ZN(n6512) );
  INV_X1 U5900 ( .A(n6512), .ZN(n6476) );
  INV_X1 U5901 ( .A(DATAI_19_), .ZN(n4767) );
  NOR2_X1 U5902 ( .A1(n6211), .A2(n4767), .ZN(n6473) );
  INV_X1 U5903 ( .A(n6473), .ZN(n6517) );
  OAI22_X1 U5904 ( .A1(n4930), .A2(n6476), .B1(n6517), .B2(n5067), .ZN(n4769)
         );
  NAND2_X1 U5905 ( .A1(DATAI_3_), .A2(n5038), .ZN(n6429) );
  NOR2_X1 U5906 ( .A1(n6429), .A2(n4857), .ZN(n4768) );
  AOI211_X1 U5907 ( .C1(INSTQUEUE_REG_15__3__SCAN_IN), .C2(n4860), .A(n4769), 
        .B(n4768), .ZN(n4770) );
  OAI21_X1 U5908 ( .B1(n4862), .B2(n5162), .A(n4770), .ZN(U3143) );
  INV_X1 U5909 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6155) );
  INV_X1 U5910 ( .A(DATAI_7_), .ZN(n6975) );
  OAI222_X1 U5911 ( .A1(n5916), .A2(n5083), .B1(n5396), .B2(n6155), .C1(n6975), 
        .C2(n5088), .ZN(U2884) );
  OAI21_X1 U5912 ( .B1(n4771), .B2(n4773), .A(n4772), .ZN(n5183) );
  AOI22_X1 U5913 ( .A1(n5363), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6133), .ZN(n4774) );
  OAI21_X1 U5914 ( .B1(n5183), .B2(n5916), .A(n4774), .ZN(U2883) );
  OAI21_X1 U5915 ( .B1(n4776), .B2(n4775), .A(n4984), .ZN(n5109) );
  INV_X1 U5916 ( .A(n5109), .ZN(n6258) );
  AOI22_X1 U5917 ( .A1(n6124), .A2(n6258), .B1(n5454), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4777) );
  OAI21_X1 U5918 ( .B1(n5183), .B2(n5456), .A(n4777), .ZN(U2851) );
  INV_X1 U5919 ( .A(n4728), .ZN(n4778) );
  AOI21_X1 U5920 ( .B1(n4779), .B2(n4681), .A(n4778), .ZN(n6202) );
  NAND2_X1 U5921 ( .A1(n4684), .A2(n4780), .ZN(n4781) );
  NAND2_X1 U5922 ( .A1(n4782), .A2(n4781), .ZN(n6060) );
  OAI22_X1 U5923 ( .A1(n7014), .A2(n6060), .B1(n4783), .B2(n7016), .ZN(n4784)
         );
  AOI21_X1 U5924 ( .B1(n6202), .B2(n6125), .A(n4784), .ZN(n4785) );
  INV_X1 U5925 ( .A(n4785), .ZN(U2853) );
  INV_X1 U5926 ( .A(n6202), .ZN(n4787) );
  INV_X1 U5927 ( .A(DATAI_6_), .ZN(n6887) );
  OAI222_X1 U5928 ( .A1(n4787), .A2(n5916), .B1(n5088), .B2(n6887), .C1(n4786), 
        .C2(n5396), .ZN(U2885) );
  INV_X1 U5929 ( .A(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4792) );
  NAND2_X1 U5930 ( .A1(DATAI_5_), .A2(n5038), .ZN(n6436) );
  AOI22_X1 U5931 ( .A1(n6482), .A2(n6534), .B1(n6481), .B2(n6532), .ZN(n4791)
         );
  INV_X1 U5932 ( .A(DATAI_21_), .ZN(n4788) );
  NOR2_X1 U5933 ( .A1(n5564), .A2(n4788), .ZN(n6483) );
  NAND2_X1 U5934 ( .A1(n6223), .A2(DATAI_29_), .ZN(n6486) );
  INV_X1 U5935 ( .A(n6486), .ZN(n6433) );
  AOI22_X1 U5936 ( .A1(n6483), .A2(n4789), .B1(n6530), .B2(n6433), .ZN(n4790)
         );
  OAI211_X1 U5937 ( .C1(n4793), .C2(n4792), .A(n4791), .B(n4790), .ZN(U3113)
         );
  NAND3_X1 U5938 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6762), .A3(n5033), .ZN(n6450) );
  NOR2_X1 U5939 ( .A1(n6372), .A2(n6450), .ZN(n4794) );
  INV_X1 U5940 ( .A(n4794), .ZN(n4921) );
  OAI21_X1 U5941 ( .B1(n4800), .B2(n5991), .A(n6674), .ZN(n4798) );
  OR2_X1 U5942 ( .A1(n4591), .A2(n4519), .ZN(n6453) );
  INV_X1 U5943 ( .A(n6453), .ZN(n4795) );
  AOI21_X1 U5944 ( .B1(n4866), .B2(n4795), .A(n4794), .ZN(n4799) );
  INV_X1 U5945 ( .A(n4799), .ZN(n4797) );
  NAND2_X1 U5946 ( .A1(n6694), .A2(n6450), .ZN(n4796) );
  OAI211_X1 U5947 ( .C1(n4798), .C2(n4797), .A(n6414), .B(n4796), .ZN(n4918)
         );
  OAI22_X1 U5948 ( .A1(n4799), .A2(n4798), .B1(n6334), .B2(n6450), .ZN(n4917)
         );
  AOI22_X1 U5949 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4918), .B1(n6535), 
        .B2(n4917), .ZN(n4802) );
  INV_X1 U5950 ( .A(n6499), .ZN(n6531) );
  AOI22_X1 U5951 ( .A1(n6494), .A2(n6531), .B1(n5282), .B2(n6493), .ZN(n4801)
         );
  OAI211_X1 U5952 ( .C1(n4921), .C2(n5138), .A(n4802), .B(n4801), .ZN(U3099)
         );
  AOI22_X1 U5953 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4918), .B1(n6514), 
        .B2(n4917), .ZN(n4804) );
  AOI22_X1 U5954 ( .A1(n6494), .A2(n6512), .B1(n5282), .B2(n6473), .ZN(n4803)
         );
  OAI211_X1 U5955 ( .C1(n4921), .C2(n5162), .A(n4804), .B(n4803), .ZN(U3095)
         );
  AOI22_X1 U5956 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4918), .B1(n6502), 
        .B2(n4917), .ZN(n4806) );
  AOI22_X1 U5957 ( .A1(n6500), .A2(n6494), .B1(n5282), .B2(n6459), .ZN(n4805)
         );
  OAI211_X1 U5958 ( .C1(n4921), .C2(n5170), .A(n4806), .B(n4805), .ZN(U3092)
         );
  AOI22_X1 U5959 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4918), .B1(n6468), 
        .B2(n4917), .ZN(n4808) );
  AOI22_X1 U5960 ( .A1(n6494), .A2(n6423), .B1(n5282), .B2(n6469), .ZN(n4807)
         );
  OAI211_X1 U5961 ( .C1(n4921), .C2(n5142), .A(n4808), .B(n4807), .ZN(U3094)
         );
  AOI22_X1 U5962 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4918), .B1(n6508), 
        .B2(n4917), .ZN(n4810) );
  AOI22_X1 U5963 ( .A1(n6494), .A2(n6506), .B1(n5282), .B2(n6463), .ZN(n4809)
         );
  OAI211_X1 U5964 ( .C1(n4921), .C2(n5158), .A(n4810), .B(n4809), .ZN(U3093)
         );
  OAI21_X1 U5965 ( .B1(n3113), .B2(n4812), .A(n3114), .ZN(n6201) );
  NOR2_X1 U5966 ( .A1(n6294), .A2(n6060), .ZN(n4820) );
  AOI21_X1 U5967 ( .B1(n6309), .B2(n6318), .A(n6310), .ZN(n6289) );
  INV_X1 U5968 ( .A(n4814), .ZN(n4816) );
  NOR2_X1 U5969 ( .A1(n6289), .A2(n4816), .ZN(n4818) );
  INV_X1 U5970 ( .A(n5599), .ZN(n6241) );
  OAI21_X1 U5971 ( .B1(n4815), .B2(n6309), .A(n6239), .ZN(n6316) );
  AOI21_X1 U5972 ( .B1(n6241), .B2(n4816), .A(n6316), .ZN(n6287) );
  INV_X1 U5973 ( .A(n6287), .ZN(n4817) );
  MUX2_X1 U5974 ( .A(n4818), .B(n4817), .S(INSTADDRPOINTER_REG_6__SCAN_IN), 
        .Z(n4819) );
  AOI211_X1 U5975 ( .C1(n6317), .C2(REIP_REG_6__SCAN_IN), .A(n4820), .B(n4819), 
        .ZN(n4821) );
  OAI21_X1 U5976 ( .B1(n5745), .B2(n6201), .A(n4821), .ZN(U3012) );
  NAND2_X1 U5977 ( .A1(n4822), .A2(n6681), .ZN(n6335) );
  NOR2_X1 U5978 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6335), .ZN(n4827)
         );
  INV_X1 U5979 ( .A(n4827), .ZN(n4928) );
  INV_X1 U5980 ( .A(n5044), .ZN(n4823) );
  NOR2_X1 U5981 ( .A1(n4823), .A2(n5043), .ZN(n4830) );
  OAI21_X1 U5982 ( .B1(n4830), .B2(n6358), .A(n6374), .ZN(n4825) );
  OR2_X1 U5983 ( .A1(n4824), .A2(n6677), .ZN(n6331) );
  AOI21_X1 U5984 ( .B1(n4825), .B2(n6331), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4828) );
  AOI21_X1 U5985 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5279), .A(n5128), .ZN(
        n5289) );
  NAND2_X1 U5986 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4826) );
  AND2_X1 U5987 ( .A1(n5289), .A2(n4826), .ZN(n6380) );
  NAND2_X1 U5988 ( .A1(n4922), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4833) );
  NAND2_X1 U5989 ( .A1(n4935), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6448) );
  INV_X1 U5990 ( .A(n6448), .ZN(n5196) );
  INV_X1 U5991 ( .A(n5279), .ZN(n6367) );
  NAND3_X1 U5992 ( .A1(n5196), .A2(n6367), .A3(n6681), .ZN(n4829) );
  OAI21_X1 U5993 ( .B1(n6331), .B2(n6694), .A(n4829), .ZN(n4925) );
  OAI22_X1 U5994 ( .A1(n5799), .A2(n6466), .B1(n6511), .B2(n4923), .ZN(n4831)
         );
  AOI21_X1 U5995 ( .B1(n6508), .B2(n4925), .A(n4831), .ZN(n4832) );
  OAI211_X1 U5996 ( .C1(n4928), .C2(n5158), .A(n4833), .B(n4832), .ZN(U3037)
         );
  NAND2_X1 U5997 ( .A1(n4922), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4836) );
  OAI22_X1 U5998 ( .A1(n5799), .A2(n6476), .B1(n6517), .B2(n4923), .ZN(n4834)
         );
  AOI21_X1 U5999 ( .B1(n6514), .B2(n4925), .A(n4834), .ZN(n4835) );
  OAI211_X1 U6000 ( .C1(n4928), .C2(n5162), .A(n4836), .B(n4835), .ZN(U3039)
         );
  NAND2_X1 U6001 ( .A1(n4922), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4839) );
  OAI22_X1 U6002 ( .A1(n5799), .A2(n6472), .B1(n6388), .B2(n4923), .ZN(n4837)
         );
  AOI21_X1 U6003 ( .B1(n6468), .B2(n4925), .A(n4837), .ZN(n4838) );
  OAI211_X1 U6004 ( .C1(n4928), .C2(n5142), .A(n4839), .B(n4838), .ZN(U3038)
         );
  NAND2_X1 U6005 ( .A1(n4922), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4842) );
  OAI22_X1 U6006 ( .A1(n5799), .A2(n6499), .B1(n6540), .B2(n4923), .ZN(n4840)
         );
  AOI21_X1 U6007 ( .B1(n6535), .B2(n4925), .A(n4840), .ZN(n4841) );
  OAI211_X1 U6008 ( .C1(n4928), .C2(n5138), .A(n4842), .B(n4841), .ZN(U3043)
         );
  NAND2_X1 U6009 ( .A1(n4922), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4845) );
  OAI22_X1 U6010 ( .A1(n5799), .A2(n6462), .B1(n6505), .B2(n4923), .ZN(n4843)
         );
  AOI21_X1 U6011 ( .B1(n6502), .B2(n4925), .A(n4843), .ZN(n4844) );
  OAI211_X1 U6012 ( .C1(n5170), .C2(n4928), .A(n4845), .B(n4844), .ZN(U3036)
         );
  INV_X1 U6013 ( .A(n6483), .ZN(n6395) );
  OAI22_X1 U6014 ( .A1(n4930), .A2(n6486), .B1(n6395), .B2(n5067), .ZN(n4847)
         );
  NOR2_X1 U6015 ( .A1(n6436), .A2(n4857), .ZN(n4846) );
  AOI211_X1 U6016 ( .C1(INSTQUEUE_REG_15__5__SCAN_IN), .C2(n4860), .A(n4847), 
        .B(n4846), .ZN(n4848) );
  OAI21_X1 U6017 ( .B1(n4862), .B2(n5154), .A(n4848), .ZN(U3145) );
  NOR2_X1 U6018 ( .A1(n4854), .A2(n3337), .ZN(n6525) );
  INV_X1 U6019 ( .A(DATAI_30_), .ZN(n4849) );
  NOR2_X1 U6020 ( .A1(n5564), .A2(n4849), .ZN(n6524) );
  INV_X1 U6021 ( .A(n6524), .ZN(n6490) );
  INV_X1 U6022 ( .A(DATAI_22_), .ZN(n4850) );
  NOR2_X1 U6023 ( .A1(n6211), .A2(n4850), .ZN(n6487) );
  INV_X1 U6024 ( .A(n6487), .ZN(n6529) );
  OAI22_X1 U6025 ( .A1(n4930), .A2(n6490), .B1(n6529), .B2(n5067), .ZN(n4852)
         );
  NAND2_X1 U6026 ( .A1(DATAI_6_), .A2(n5038), .ZN(n6439) );
  NOR2_X1 U6027 ( .A1(n6439), .A2(n4857), .ZN(n4851) );
  AOI211_X1 U6028 ( .C1(INSTQUEUE_REG_15__6__SCAN_IN), .C2(n4860), .A(n4852), 
        .B(n4851), .ZN(n4853) );
  OAI21_X1 U6029 ( .B1(n4862), .B2(n5150), .A(n4853), .ZN(U3146) );
  INV_X1 U6030 ( .A(DATAI_28_), .ZN(n4855) );
  NOR2_X1 U6031 ( .A1(n5564), .A2(n4855), .ZN(n6518) );
  INV_X1 U6032 ( .A(n6518), .ZN(n6480) );
  INV_X1 U6033 ( .A(DATAI_20_), .ZN(n4856) );
  NOR2_X1 U6034 ( .A1(n6211), .A2(n4856), .ZN(n6477) );
  INV_X1 U6035 ( .A(n6477), .ZN(n6523) );
  OAI22_X1 U6036 ( .A1(n4930), .A2(n6480), .B1(n6523), .B2(n5067), .ZN(n4859)
         );
  NAND2_X1 U6037 ( .A1(DATAI_4_), .A2(n5038), .ZN(n6432) );
  NOR2_X1 U6038 ( .A1(n6432), .A2(n4857), .ZN(n4858) );
  AOI211_X1 U6039 ( .C1(INSTQUEUE_REG_15__4__SCAN_IN), .C2(n4860), .A(n4859), 
        .B(n4858), .ZN(n4861) );
  OAI21_X1 U6040 ( .B1(n4862), .B2(n5146), .A(n4861), .ZN(U3144) );
  NOR3_X1 U6041 ( .A1(n6762), .A2(n6681), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n5125) );
  INV_X1 U6042 ( .A(n5125), .ZN(n4871) );
  NOR2_X1 U6043 ( .A1(n6372), .A2(n4871), .ZN(n4865) );
  INV_X1 U6044 ( .A(n4865), .ZN(n4911) );
  NOR2_X1 U6045 ( .A1(n4993), .A2(n4989), .ZN(n4863) );
  NAND2_X1 U6046 ( .A1(n4867), .A2(n5043), .ZN(n5129) );
  NAND2_X1 U6047 ( .A1(n4591), .A2(n4864), .ZN(n5190) );
  INV_X1 U6048 ( .A(n5190), .ZN(n5132) );
  AOI21_X1 U6049 ( .B1(n4866), .B2(n5132), .A(n4865), .ZN(n4872) );
  NAND2_X1 U6050 ( .A1(n4867), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6324) );
  NAND2_X1 U6051 ( .A1(n4872), .A2(n6324), .ZN(n4868) );
  OR2_X1 U6052 ( .A1(n6694), .A2(n4868), .ZN(n4870) );
  NAND2_X1 U6053 ( .A1(n6694), .A2(n4871), .ZN(n4869) );
  INV_X1 U6054 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n6818) );
  OAI22_X1 U6055 ( .A1(n5129), .A2(n6499), .B1(n4906), .B2(n6818), .ZN(n4875)
         );
  OAI22_X1 U6056 ( .A1(n4872), .A2(n6694), .B1(n4871), .B2(n6334), .ZN(n4873)
         );
  NOR2_X1 U6057 ( .A1(n6445), .A2(n4907), .ZN(n4874) );
  AOI211_X1 U6058 ( .C1(n4966), .C2(n6493), .A(n4875), .B(n4874), .ZN(n4876)
         );
  OAI21_X1 U6059 ( .B1(n5138), .B2(n4911), .A(n4876), .ZN(U3131) );
  INV_X1 U6060 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4877) );
  OAI22_X1 U6061 ( .A1(n5129), .A2(n6472), .B1(n4906), .B2(n4877), .ZN(n4879)
         );
  NOR2_X1 U6062 ( .A1(n6426), .A2(n4907), .ZN(n4878) );
  AOI211_X1 U6063 ( .C1(n4966), .C2(n6469), .A(n4879), .B(n4878), .ZN(n4880)
         );
  OAI21_X1 U6064 ( .B1(n5142), .B2(n4911), .A(n4880), .ZN(U3126) );
  INV_X1 U6065 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4881) );
  OAI22_X1 U6066 ( .A1(n5129), .A2(n6480), .B1(n4906), .B2(n4881), .ZN(n4883)
         );
  NOR2_X1 U6067 ( .A1(n6432), .A2(n4907), .ZN(n4882) );
  AOI211_X1 U6068 ( .C1(n4966), .C2(n6477), .A(n4883), .B(n4882), .ZN(n4884)
         );
  OAI21_X1 U6069 ( .B1(n5146), .B2(n4911), .A(n4884), .ZN(U3128) );
  INV_X1 U6070 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4885) );
  OAI22_X1 U6071 ( .A1(n5129), .A2(n6490), .B1(n4906), .B2(n4885), .ZN(n4887)
         );
  NOR2_X1 U6072 ( .A1(n6439), .A2(n4907), .ZN(n4886) );
  AOI211_X1 U6073 ( .C1(n4966), .C2(n6487), .A(n4887), .B(n4886), .ZN(n4888)
         );
  OAI21_X1 U6074 ( .B1(n5150), .B2(n4911), .A(n4888), .ZN(U3130) );
  AOI22_X1 U6075 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4918), .B1(n6482), 
        .B2(n4917), .ZN(n4890) );
  AOI22_X1 U6076 ( .A1(n6494), .A2(n6433), .B1(n5282), .B2(n6483), .ZN(n4889)
         );
  OAI211_X1 U6077 ( .C1(n4921), .C2(n5154), .A(n4890), .B(n4889), .ZN(U3097)
         );
  NAND2_X1 U6078 ( .A1(n4922), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4893) );
  OAI22_X1 U6079 ( .A1(n5799), .A2(n6486), .B1(n6395), .B2(n4923), .ZN(n4891)
         );
  AOI21_X1 U6080 ( .B1(n6482), .B2(n4925), .A(n4891), .ZN(n4892) );
  OAI211_X1 U6081 ( .C1(n4928), .C2(n5154), .A(n4893), .B(n4892), .ZN(U3041)
         );
  INV_X1 U6082 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4894) );
  OAI22_X1 U6083 ( .A1(n5129), .A2(n6486), .B1(n4906), .B2(n4894), .ZN(n4896)
         );
  NOR2_X1 U6084 ( .A1(n6436), .A2(n4907), .ZN(n4895) );
  AOI211_X1 U6085 ( .C1(n4966), .C2(n6483), .A(n4896), .B(n4895), .ZN(n4897)
         );
  OAI21_X1 U6086 ( .B1(n5154), .B2(n4911), .A(n4897), .ZN(U3129) );
  INV_X1 U6087 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4898) );
  OAI22_X1 U6088 ( .A1(n5129), .A2(n6476), .B1(n4906), .B2(n4898), .ZN(n4900)
         );
  NOR2_X1 U6089 ( .A1(n6429), .A2(n4907), .ZN(n4899) );
  AOI211_X1 U6090 ( .C1(n4966), .C2(n6473), .A(n4900), .B(n4899), .ZN(n4901)
         );
  OAI21_X1 U6091 ( .B1(n5162), .B2(n4911), .A(n4901), .ZN(U3127) );
  OAI22_X1 U6092 ( .A1(n5129), .A2(n6462), .B1(n4906), .B2(n6824), .ZN(n4903)
         );
  NOR2_X1 U6093 ( .A1(n6419), .A2(n4907), .ZN(n4902) );
  AOI211_X1 U6094 ( .C1(n4966), .C2(n6459), .A(n4903), .B(n4902), .ZN(n4904)
         );
  OAI21_X1 U6095 ( .B1(n5170), .B2(n4911), .A(n4904), .ZN(U3124) );
  INV_X1 U6096 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4905) );
  OAI22_X1 U6097 ( .A1(n5129), .A2(n6466), .B1(n4906), .B2(n4905), .ZN(n4909)
         );
  NOR2_X1 U6098 ( .A1(n6422), .A2(n4907), .ZN(n4908) );
  AOI211_X1 U6099 ( .C1(n4966), .C2(n6463), .A(n4909), .B(n4908), .ZN(n4910)
         );
  OAI21_X1 U6100 ( .B1(n5158), .B2(n4911), .A(n4910), .ZN(U3125) );
  AOI22_X1 U6101 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4918), .B1(n6526), 
        .B2(n4917), .ZN(n4913) );
  AOI22_X1 U6102 ( .A1(n6494), .A2(n6524), .B1(n5282), .B2(n6487), .ZN(n4912)
         );
  OAI211_X1 U6103 ( .C1(n4921), .C2(n5150), .A(n4913), .B(n4912), .ZN(U3098)
         );
  NAND2_X1 U6104 ( .A1(n4922), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4916) );
  OAI22_X1 U6105 ( .A1(n5799), .A2(n6480), .B1(n6523), .B2(n4923), .ZN(n4914)
         );
  AOI21_X1 U6106 ( .B1(n6520), .B2(n4925), .A(n4914), .ZN(n4915) );
  OAI211_X1 U6107 ( .C1(n4928), .C2(n5146), .A(n4916), .B(n4915), .ZN(U3040)
         );
  AOI22_X1 U6108 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4918), .B1(n6520), 
        .B2(n4917), .ZN(n4920) );
  AOI22_X1 U6109 ( .A1(n6494), .A2(n6518), .B1(n5282), .B2(n6477), .ZN(n4919)
         );
  OAI211_X1 U6110 ( .C1(n4921), .C2(n5146), .A(n4920), .B(n4919), .ZN(U3096)
         );
  NAND2_X1 U6111 ( .A1(n4922), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4927) );
  OAI22_X1 U6112 ( .A1(n5799), .A2(n6490), .B1(n6529), .B2(n4923), .ZN(n4924)
         );
  AOI21_X1 U6113 ( .B1(n6526), .B2(n4925), .A(n4924), .ZN(n4926) );
  OAI211_X1 U6114 ( .C1(n4928), .C2(n5150), .A(n4927), .B(n4926), .ZN(U3042)
         );
  INV_X1 U6115 ( .A(n4966), .ZN(n4929) );
  NAND3_X1 U6116 ( .A1(n4930), .A2(n6674), .A3(n4929), .ZN(n4931) );
  AOI22_X1 U6117 ( .A1(n4931), .A2(n6374), .B1(n6376), .B2(n6677), .ZN(n4934)
         );
  AND2_X1 U6118 ( .A1(n6372), .A2(n4932), .ZN(n4971) );
  NAND2_X1 U6119 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6681), .ZN(n5287) );
  OAI211_X1 U6120 ( .C1(n6662), .C2(n4971), .A(n5289), .B(n5287), .ZN(n4933)
         );
  NOR3_X2 U6121 ( .A1(n4934), .A2(n5196), .A3(n4933), .ZN(n4974) );
  INV_X1 U6122 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4941) );
  NOR2_X1 U6123 ( .A1(n6454), .A2(n6694), .ZN(n5126) );
  INV_X1 U6124 ( .A(n4935), .ZN(n4936) );
  NAND2_X1 U6125 ( .A1(n4936), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6455) );
  NOR3_X1 U6126 ( .A1(n6455), .A2(n6681), .A3(n5279), .ZN(n4937) );
  AOI21_X1 U6127 ( .B1(n5126), .B2(n6376), .A(n4937), .ZN(n4969) );
  AOI22_X1 U6128 ( .A1(n6463), .A2(n4967), .B1(n4966), .B2(n6506), .ZN(n4938)
         );
  OAI21_X1 U6129 ( .B1(n6422), .B2(n4969), .A(n4938), .ZN(n4939) );
  AOI21_X1 U6130 ( .B1(n6507), .B2(n4971), .A(n4939), .ZN(n4940) );
  OAI21_X1 U6131 ( .B1(n4974), .B2(n4941), .A(n4940), .ZN(U3133) );
  INV_X1 U6132 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4945) );
  AOI22_X1 U6133 ( .A1(n6469), .A2(n4967), .B1(n4966), .B2(n6423), .ZN(n4942)
         );
  OAI21_X1 U6134 ( .B1(n6426), .B2(n4969), .A(n4942), .ZN(n4943) );
  AOI21_X1 U6135 ( .B1(n6467), .B2(n4971), .A(n4943), .ZN(n4944) );
  OAI21_X1 U6136 ( .B1(n4974), .B2(n4945), .A(n4944), .ZN(U3134) );
  INV_X1 U6137 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4949) );
  AOI22_X1 U6138 ( .A1(n6483), .A2(n4967), .B1(n4966), .B2(n6433), .ZN(n4946)
         );
  OAI21_X1 U6139 ( .B1(n6436), .B2(n4969), .A(n4946), .ZN(n4947) );
  AOI21_X1 U6140 ( .B1(n6481), .B2(n4971), .A(n4947), .ZN(n4948) );
  OAI21_X1 U6141 ( .B1(n4974), .B2(n4949), .A(n4948), .ZN(U3137) );
  INV_X1 U6142 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4953) );
  AOI22_X1 U6143 ( .A1(n6477), .A2(n4967), .B1(n4966), .B2(n6518), .ZN(n4950)
         );
  OAI21_X1 U6144 ( .B1(n6432), .B2(n4969), .A(n4950), .ZN(n4951) );
  AOI21_X1 U6145 ( .B1(n6519), .B2(n4971), .A(n4951), .ZN(n4952) );
  OAI21_X1 U6146 ( .B1(n4974), .B2(n4953), .A(n4952), .ZN(U3136) );
  INV_X1 U6147 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4957) );
  AOI22_X1 U6148 ( .A1(n6459), .A2(n4967), .B1(n4966), .B2(n6500), .ZN(n4954)
         );
  OAI21_X1 U6149 ( .B1(n6419), .B2(n4969), .A(n4954), .ZN(n4955) );
  AOI21_X1 U6150 ( .B1(n6501), .B2(n4971), .A(n4955), .ZN(n4956) );
  OAI21_X1 U6151 ( .B1(n4974), .B2(n4957), .A(n4956), .ZN(U3132) );
  INV_X1 U6152 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U6153 ( .A1(n6487), .A2(n4967), .B1(n4966), .B2(n6524), .ZN(n4958)
         );
  OAI21_X1 U6154 ( .B1(n6439), .B2(n4969), .A(n4958), .ZN(n4959) );
  AOI21_X1 U6155 ( .B1(n6525), .B2(n4971), .A(n4959), .ZN(n4960) );
  OAI21_X1 U6156 ( .B1(n4974), .B2(n4961), .A(n4960), .ZN(U3138) );
  INV_X1 U6157 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U6158 ( .A1(n6473), .A2(n4967), .B1(n4966), .B2(n6512), .ZN(n4962)
         );
  OAI21_X1 U6159 ( .B1(n6429), .B2(n4969), .A(n4962), .ZN(n4963) );
  AOI21_X1 U6160 ( .B1(n6513), .B2(n4971), .A(n4963), .ZN(n4964) );
  OAI21_X1 U6161 ( .B1(n4974), .B2(n4965), .A(n4964), .ZN(U3135) );
  INV_X1 U6162 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U6163 ( .A1(n6493), .A2(n4967), .B1(n4966), .B2(n6531), .ZN(n4968)
         );
  OAI21_X1 U6164 ( .B1(n6445), .B2(n4969), .A(n4968), .ZN(n4970) );
  AOI21_X1 U6165 ( .B1(n6533), .B2(n4971), .A(n4970), .ZN(n4972) );
  OAI21_X1 U6166 ( .B1(n4974), .B2(n4973), .A(n4972), .ZN(U3139) );
  OAI21_X1 U6167 ( .B1(n4977), .B2(n4976), .A(n4975), .ZN(n6268) );
  NAND2_X1 U6168 ( .A1(n6317), .A2(REIP_REG_7__SCAN_IN), .ZN(n6265) );
  OAI21_X1 U6169 ( .B1(n5955), .B2(n6778), .A(n6265), .ZN(n4979) );
  NOR2_X1 U6170 ( .A1(n5083), .A2(n5564), .ZN(n4978) );
  AOI211_X1 U6171 ( .C1(n6196), .C2(n5078), .A(n4979), .B(n4978), .ZN(n4980)
         );
  OAI21_X1 U6172 ( .B1(n6213), .B2(n6268), .A(n4980), .ZN(U2979) );
  AOI21_X1 U6173 ( .B1(n4982), .B2(n4772), .A(n3779), .ZN(n6054) );
  INV_X1 U6174 ( .A(n6054), .ZN(n4988) );
  INV_X1 U6175 ( .A(n5090), .ZN(n4983) );
  AOI21_X1 U6176 ( .B1(n4985), .B2(n4984), .A(n4983), .ZN(n6249) );
  AOI22_X1 U6177 ( .A1(n6124), .A2(n6249), .B1(n5454), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n4986) );
  OAI21_X1 U6178 ( .B1(n4988), .B2(n5456), .A(n4986), .ZN(U2850) );
  AOI22_X1 U6179 ( .A1(n5363), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6133), .ZN(n4987) );
  OAI21_X1 U6180 ( .B1(n4988), .B2(n5916), .A(n4987), .ZN(U2882) );
  NAND3_X1 U6181 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6681), .A3(n5033), .ZN(n5188) );
  NOR2_X1 U6182 ( .A1(n6372), .A2(n5188), .ZN(n4992) );
  INV_X1 U6183 ( .A(n4992), .ZN(n5032) );
  NAND2_X1 U6184 ( .A1(n4990), .A2(n4989), .ZN(n6411) );
  OR3_X1 U6185 ( .A1(n6411), .A2(n4993), .A3(n5991), .ZN(n4991) );
  NAND2_X1 U6186 ( .A1(n4991), .A2(n6674), .ZN(n5192) );
  NOR2_X1 U6187 ( .A1(n5190), .A2(n5131), .ZN(n5193) );
  AOI21_X1 U6188 ( .B1(n5193), .B2(n3690), .A(n4992), .ZN(n4997) );
  OAI22_X1 U6189 ( .A1(n5192), .A2(n4997), .B1(n5188), .B2(n6334), .ZN(n5030)
         );
  OR2_X1 U6190 ( .A1(n6411), .A2(n4993), .ZN(n4995) );
  NOR2_X1 U6191 ( .A1(n5230), .A2(n6486), .ZN(n5001) );
  INV_X1 U6192 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4999) );
  INV_X1 U6193 ( .A(n5192), .ZN(n4996) );
  AOI22_X1 U6194 ( .A1(n4997), .A2(n4996), .B1(n5188), .B2(n6694), .ZN(n4998)
         );
  OAI22_X1 U6195 ( .A1(n6373), .A2(n6395), .B1(n4999), .B2(n5026), .ZN(n5000)
         );
  AOI211_X1 U6196 ( .C1(n6482), .C2(n5030), .A(n5001), .B(n5000), .ZN(n5002)
         );
  OAI21_X1 U6197 ( .B1(n5154), .B2(n5032), .A(n5002), .ZN(U3065) );
  NOR2_X1 U6198 ( .A1(n5230), .A2(n6472), .ZN(n5005) );
  INV_X1 U6199 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n5003) );
  OAI22_X1 U6200 ( .A1(n6373), .A2(n6388), .B1(n5003), .B2(n5026), .ZN(n5004)
         );
  AOI211_X1 U6201 ( .C1(n6468), .C2(n5030), .A(n5005), .B(n5004), .ZN(n5006)
         );
  OAI21_X1 U6202 ( .B1(n5142), .B2(n5032), .A(n5006), .ZN(U3062) );
  NOR2_X1 U6203 ( .A1(n5230), .A2(n6490), .ZN(n5009) );
  INV_X1 U6204 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5007) );
  OAI22_X1 U6205 ( .A1(n6373), .A2(n6529), .B1(n5007), .B2(n5026), .ZN(n5008)
         );
  AOI211_X1 U6206 ( .C1(n6526), .C2(n5030), .A(n5009), .B(n5008), .ZN(n5010)
         );
  OAI21_X1 U6207 ( .B1(n5150), .B2(n5032), .A(n5010), .ZN(U3066) );
  NOR2_X1 U6208 ( .A1(n5230), .A2(n6480), .ZN(n5013) );
  INV_X1 U6209 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5011) );
  OAI22_X1 U6210 ( .A1(n6373), .A2(n6523), .B1(n5011), .B2(n5026), .ZN(n5012)
         );
  AOI211_X1 U6211 ( .C1(n6520), .C2(n5030), .A(n5013), .B(n5012), .ZN(n5014)
         );
  OAI21_X1 U6212 ( .B1(n5146), .B2(n5032), .A(n5014), .ZN(U3064) );
  NOR2_X1 U6213 ( .A1(n5230), .A2(n6462), .ZN(n5017) );
  INV_X1 U6214 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n5015) );
  OAI22_X1 U6215 ( .A1(n6373), .A2(n6505), .B1(n5015), .B2(n5026), .ZN(n5016)
         );
  AOI211_X1 U6216 ( .C1(n6502), .C2(n5030), .A(n5017), .B(n5016), .ZN(n5018)
         );
  OAI21_X1 U6217 ( .B1(n5170), .B2(n5032), .A(n5018), .ZN(U3060) );
  NOR2_X1 U6218 ( .A1(n5230), .A2(n6466), .ZN(n5020) );
  INV_X1 U6219 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6914) );
  OAI22_X1 U6220 ( .A1(n6373), .A2(n6511), .B1(n6914), .B2(n5026), .ZN(n5019)
         );
  AOI211_X1 U6221 ( .C1(n6508), .C2(n5030), .A(n5020), .B(n5019), .ZN(n5021)
         );
  OAI21_X1 U6222 ( .B1(n5158), .B2(n5032), .A(n5021), .ZN(U3061) );
  NOR2_X1 U6223 ( .A1(n5230), .A2(n6499), .ZN(n5024) );
  INV_X1 U6224 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5022) );
  OAI22_X1 U6225 ( .A1(n6373), .A2(n6540), .B1(n5022), .B2(n5026), .ZN(n5023)
         );
  AOI211_X1 U6226 ( .C1(n6535), .C2(n5030), .A(n5024), .B(n5023), .ZN(n5025)
         );
  OAI21_X1 U6227 ( .B1(n5138), .B2(n5032), .A(n5025), .ZN(U3067) );
  NOR2_X1 U6228 ( .A1(n5230), .A2(n6476), .ZN(n5029) );
  INV_X1 U6229 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5027) );
  OAI22_X1 U6230 ( .A1(n6373), .A2(n6517), .B1(n5027), .B2(n5026), .ZN(n5028)
         );
  AOI211_X1 U6231 ( .C1(n6514), .C2(n5030), .A(n5029), .B(n5028), .ZN(n5031)
         );
  OAI21_X1 U6232 ( .B1(n5162), .B2(n5032), .A(n5031), .ZN(U3063) );
  NAND3_X1 U6233 ( .A1(n6681), .A2(n6762), .A3(n5033), .ZN(n5771) );
  NOR2_X1 U6234 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5771), .ZN(n5041)
         );
  INV_X1 U6235 ( .A(n5041), .ZN(n5072) );
  INV_X1 U6236 ( .A(n5067), .ZN(n5036) );
  INV_X1 U6237 ( .A(n5767), .ZN(n5035) );
  OAI21_X1 U6238 ( .B1(n5044), .B2(n6694), .A(n6374), .ZN(n5772) );
  INV_X1 U6239 ( .A(n5772), .ZN(n5034) );
  AOI211_X1 U6240 ( .C1(n5036), .C2(n6374), .A(n5035), .B(n5034), .ZN(n5039)
         );
  INV_X1 U6241 ( .A(n5037), .ZN(n5127) );
  NOR2_X1 U6242 ( .A1(n6367), .A2(n5127), .ZN(n5042) );
  OAI21_X1 U6243 ( .B1(n5042), .B2(n6334), .A(n5038), .ZN(n5195) );
  NOR2_X1 U6244 ( .A1(n5039), .A2(n5195), .ZN(n5040) );
  NAND2_X1 U6245 ( .A1(n5066), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5047) );
  INV_X1 U6246 ( .A(n5042), .ZN(n5189) );
  OAI22_X1 U6247 ( .A1(n5767), .A2(n6694), .B1(n6448), .B2(n5189), .ZN(n5069)
         );
  NAND2_X1 U6248 ( .A1(n5044), .A2(n5043), .ZN(n5769) );
  OAI22_X1 U6249 ( .A1(n5769), .A2(n6523), .B1(n6480), .B2(n5067), .ZN(n5045)
         );
  AOI21_X1 U6250 ( .B1(n6520), .B2(n5069), .A(n5045), .ZN(n5046) );
  OAI211_X1 U6251 ( .C1(n5072), .C2(n5146), .A(n5047), .B(n5046), .ZN(U3024)
         );
  NAND2_X1 U6252 ( .A1(n5066), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5050) );
  OAI22_X1 U6253 ( .A1(n5769), .A2(n6529), .B1(n6490), .B2(n5067), .ZN(n5048)
         );
  AOI21_X1 U6254 ( .B1(n6526), .B2(n5069), .A(n5048), .ZN(n5049) );
  OAI211_X1 U6255 ( .C1(n5072), .C2(n5150), .A(n5050), .B(n5049), .ZN(U3026)
         );
  NAND2_X1 U6256 ( .A1(n5066), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n5053) );
  OAI22_X1 U6257 ( .A1(n5769), .A2(n6395), .B1(n6486), .B2(n5067), .ZN(n5051)
         );
  AOI21_X1 U6258 ( .B1(n6482), .B2(n5069), .A(n5051), .ZN(n5052) );
  OAI211_X1 U6259 ( .C1(n5072), .C2(n5154), .A(n5053), .B(n5052), .ZN(U3025)
         );
  NAND2_X1 U6260 ( .A1(n5066), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n5056) );
  OAI22_X1 U6261 ( .A1(n5769), .A2(n6511), .B1(n6466), .B2(n5067), .ZN(n5054)
         );
  AOI21_X1 U6262 ( .B1(n6508), .B2(n5069), .A(n5054), .ZN(n5055) );
  OAI211_X1 U6263 ( .C1(n5072), .C2(n5158), .A(n5056), .B(n5055), .ZN(U3021)
         );
  NAND2_X1 U6264 ( .A1(n5066), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n5059) );
  OAI22_X1 U6265 ( .A1(n5769), .A2(n6505), .B1(n6462), .B2(n5067), .ZN(n5057)
         );
  AOI21_X1 U6266 ( .B1(n6502), .B2(n5069), .A(n5057), .ZN(n5058) );
  OAI211_X1 U6267 ( .C1(n5170), .C2(n5072), .A(n5059), .B(n5058), .ZN(U3020)
         );
  NAND2_X1 U6268 ( .A1(n5066), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5062) );
  OAI22_X1 U6269 ( .A1(n5769), .A2(n6388), .B1(n6472), .B2(n5067), .ZN(n5060)
         );
  AOI21_X1 U6270 ( .B1(n6468), .B2(n5069), .A(n5060), .ZN(n5061) );
  OAI211_X1 U6271 ( .C1(n5072), .C2(n5142), .A(n5062), .B(n5061), .ZN(U3022)
         );
  NAND2_X1 U6272 ( .A1(n5066), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n5065) );
  OAI22_X1 U6273 ( .A1(n5769), .A2(n6517), .B1(n6476), .B2(n5067), .ZN(n5063)
         );
  AOI21_X1 U6274 ( .B1(n6514), .B2(n5069), .A(n5063), .ZN(n5064) );
  OAI211_X1 U6275 ( .C1(n5072), .C2(n5162), .A(n5065), .B(n5064), .ZN(U3023)
         );
  NAND2_X1 U6276 ( .A1(n5066), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n5071) );
  OAI22_X1 U6277 ( .A1(n5769), .A2(n6540), .B1(n6499), .B2(n5067), .ZN(n5068)
         );
  AOI21_X1 U6278 ( .B1(n6535), .B2(n5069), .A(n5068), .ZN(n5070) );
  OAI211_X1 U6279 ( .C1(n5072), .C2(n5138), .A(n5071), .B(n5070), .ZN(U3027)
         );
  INV_X1 U6280 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6619) );
  NOR2_X1 U6281 ( .A1(n6092), .A2(n5073), .ZN(n5094) );
  AND2_X1 U6282 ( .A1(n5094), .A2(REIP_REG_5__SCAN_IN), .ZN(n6038) );
  INV_X1 U6283 ( .A(n6038), .ZN(n5103) );
  NOR3_X1 U6284 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6619), .A3(n5103), .ZN(n5077)
         );
  AOI22_X1 U6285 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6110), .B1(n6107), .B2(n6267), 
        .ZN(n5075) );
  NAND2_X1 U6286 ( .A1(n5113), .A2(n5074), .ZN(n6067) );
  OAI211_X1 U6287 ( .C1(n6109), .C2(n6778), .A(n5075), .B(n6067), .ZN(n5076)
         );
  AOI211_X1 U6288 ( .C1(n6096), .C2(n5078), .A(n5077), .B(n5076), .ZN(n5082)
         );
  OR2_X1 U6289 ( .A1(n6092), .A2(n5079), .ZN(n5080) );
  NAND2_X1 U6290 ( .A1(n5080), .A2(n5113), .ZN(n6063) );
  NOR2_X1 U6291 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5103), .ZN(n6062) );
  OAI21_X1 U6292 ( .B1(n6063), .B2(n6062), .A(REIP_REG_7__SCAN_IN), .ZN(n5081)
         );
  OAI211_X1 U6293 ( .C1(n5083), .C2(n6044), .A(n5082), .B(n5081), .ZN(U2820)
         );
  NAND2_X1 U6294 ( .A1(n4981), .A2(n5085), .ZN(n5086) );
  AND2_X1 U6295 ( .A1(n5084), .A2(n5086), .ZN(n5322) );
  OAI222_X1 U6296 ( .A1(n6045), .A2(n5916), .B1(n5088), .B2(n5087), .C1(n5396), 
        .C2(n4724), .ZN(U2881) );
  AND2_X1 U6297 ( .A1(n5090), .A2(n5089), .ZN(n5091) );
  OR2_X1 U6298 ( .A1(n5091), .A2(n5185), .ZN(n6244) );
  OAI222_X1 U6299 ( .A1(n6045), .A2(n5456), .B1(n7016), .B2(n4264), .C1(n6244), 
        .C2(n7014), .ZN(U2849) );
  NAND2_X1 U6300 ( .A1(n5412), .A2(n5092), .ZN(n5093) );
  OAI21_X1 U6301 ( .B1(n5094), .B2(REIP_REG_5__SCAN_IN), .A(n6063), .ZN(n5097)
         );
  AOI21_X1 U6302 ( .B1(n6096), .B2(n5095), .A(n6041), .ZN(n5096) );
  OAI211_X1 U6303 ( .C1(n6280), .C2(n6104), .A(n5097), .B(n5096), .ZN(n5100)
         );
  OAI22_X1 U6304 ( .A1(n6959), .A2(n6049), .B1(n5098), .B2(n6109), .ZN(n5099)
         );
  NOR2_X1 U6305 ( .A1(n5100), .A2(n5099), .ZN(n5101) );
  OAI21_X1 U6306 ( .B1(n6116), .B2(n5102), .A(n5101), .ZN(U2822) );
  OAI21_X1 U6307 ( .B1(n5104), .B2(n5103), .A(n6621), .ZN(n5111) );
  INV_X1 U6308 ( .A(n6063), .ZN(n5105) );
  OAI21_X1 U6309 ( .B1(n6039), .B2(n6092), .A(n5105), .ZN(n6055) );
  AOI22_X1 U6310 ( .A1(EBX_REG_8__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n6083), .ZN(n5108) );
  INV_X1 U6311 ( .A(n5179), .ZN(n5106) );
  AOI21_X1 U6312 ( .B1(n6096), .B2(n5106), .A(n6041), .ZN(n5107) );
  OAI211_X1 U6313 ( .C1(n6104), .C2(n5109), .A(n5108), .B(n5107), .ZN(n5110)
         );
  AOI21_X1 U6314 ( .B1(n5111), .B2(n6055), .A(n5110), .ZN(n5112) );
  OAI21_X1 U6315 ( .B1(n6044), .B2(n5183), .A(n5112), .ZN(U2819) );
  OR2_X1 U6316 ( .A1(n6092), .A2(REIP_REG_1__SCAN_IN), .ZN(n5114) );
  NAND2_X1 U6317 ( .A1(n5114), .A2(n5113), .ZN(n6080) );
  AND2_X1 U6318 ( .A1(n5412), .A2(n5115), .ZN(n6111) );
  AOI22_X1 U6319 ( .A1(n6110), .A2(EBX_REG_2__SCAN_IN), .B1(n6111), .B2(n4591), 
        .ZN(n5122) );
  INV_X1 U6320 ( .A(n6227), .ZN(n5116) );
  AOI22_X1 U6321 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n6083), .B1(n6096), 
        .B2(n5116), .ZN(n5121) );
  OR3_X1 U6322 ( .A1(n6092), .A2(REIP_REG_2__SCAN_IN), .A3(n5117), .ZN(n5120)
         );
  XNOR2_X1 U6323 ( .A(n4619), .B(n5118), .ZN(n6313) );
  NAND2_X1 U6324 ( .A1(n6107), .A2(n6313), .ZN(n5119) );
  NAND4_X1 U6325 ( .A1(n5122), .A2(n5121), .A3(n5120), .A4(n5119), .ZN(n5123)
         );
  AOI21_X1 U6326 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6080), .A(n5123), .ZN(n5124)
         );
  OAI21_X1 U6327 ( .B1(n6116), .B2(n6123), .A(n5124), .ZN(U2825) );
  NAND2_X1 U6328 ( .A1(n6372), .A2(n5125), .ZN(n5169) );
  INV_X1 U6329 ( .A(n5126), .ZN(n6449) );
  NAND2_X1 U6330 ( .A1(n5127), .A2(n5279), .ZN(n6447) );
  OAI22_X1 U6331 ( .A1(n6449), .A2(n5190), .B1(n6455), .B2(n6447), .ZN(n5167)
         );
  AOI21_X1 U6332 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6447), .A(n5128), .ZN(
        n6456) );
  AOI21_X1 U6333 ( .B1(n6539), .B2(n5129), .A(n5991), .ZN(n5130) );
  AOI211_X1 U6334 ( .C1(n5132), .C2(n5131), .A(n5130), .B(n6694), .ZN(n5133)
         );
  AOI211_X1 U6335 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5169), .A(n5133), .B(
        n5196), .ZN(n5134) );
  NAND2_X1 U6336 ( .A1(n6456), .A2(n5134), .ZN(n5163) );
  AOI22_X1 U6337 ( .A1(n5164), .A2(n6493), .B1(INSTQUEUE_REG_12__7__SCAN_IN), 
        .B2(n5163), .ZN(n5135) );
  OAI21_X1 U6338 ( .B1(n6499), .B2(n6539), .A(n5135), .ZN(n5136) );
  AOI21_X1 U6339 ( .B1(n6535), .B2(n5167), .A(n5136), .ZN(n5137) );
  OAI21_X1 U6340 ( .B1(n5138), .B2(n5169), .A(n5137), .ZN(U3123) );
  AOI22_X1 U6341 ( .A1(n5164), .A2(n6469), .B1(INSTQUEUE_REG_12__2__SCAN_IN), 
        .B2(n5163), .ZN(n5139) );
  OAI21_X1 U6342 ( .B1(n6472), .B2(n6539), .A(n5139), .ZN(n5140) );
  AOI21_X1 U6343 ( .B1(n6468), .B2(n5167), .A(n5140), .ZN(n5141) );
  OAI21_X1 U6344 ( .B1(n5142), .B2(n5169), .A(n5141), .ZN(U3118) );
  AOI22_X1 U6345 ( .A1(n5164), .A2(n6477), .B1(INSTQUEUE_REG_12__4__SCAN_IN), 
        .B2(n5163), .ZN(n5143) );
  OAI21_X1 U6346 ( .B1(n6480), .B2(n6539), .A(n5143), .ZN(n5144) );
  AOI21_X1 U6347 ( .B1(n6520), .B2(n5167), .A(n5144), .ZN(n5145) );
  OAI21_X1 U6348 ( .B1(n5146), .B2(n5169), .A(n5145), .ZN(U3120) );
  AOI22_X1 U6349 ( .A1(n5164), .A2(n6487), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n5163), .ZN(n5147) );
  OAI21_X1 U6350 ( .B1(n6490), .B2(n6539), .A(n5147), .ZN(n5148) );
  AOI21_X1 U6351 ( .B1(n6526), .B2(n5167), .A(n5148), .ZN(n5149) );
  OAI21_X1 U6352 ( .B1(n5150), .B2(n5169), .A(n5149), .ZN(U3122) );
  AOI22_X1 U6353 ( .A1(n5164), .A2(n6483), .B1(INSTQUEUE_REG_12__5__SCAN_IN), 
        .B2(n5163), .ZN(n5151) );
  OAI21_X1 U6354 ( .B1(n6486), .B2(n6539), .A(n5151), .ZN(n5152) );
  AOI21_X1 U6355 ( .B1(n6482), .B2(n5167), .A(n5152), .ZN(n5153) );
  OAI21_X1 U6356 ( .B1(n5154), .B2(n5169), .A(n5153), .ZN(U3121) );
  AOI22_X1 U6357 ( .A1(n5164), .A2(n6463), .B1(INSTQUEUE_REG_12__1__SCAN_IN), 
        .B2(n5163), .ZN(n5155) );
  OAI21_X1 U6358 ( .B1(n6466), .B2(n6539), .A(n5155), .ZN(n5156) );
  AOI21_X1 U6359 ( .B1(n6508), .B2(n5167), .A(n5156), .ZN(n5157) );
  OAI21_X1 U6360 ( .B1(n5158), .B2(n5169), .A(n5157), .ZN(U3117) );
  AOI22_X1 U6361 ( .A1(n5164), .A2(n6473), .B1(INSTQUEUE_REG_12__3__SCAN_IN), 
        .B2(n5163), .ZN(n5159) );
  OAI21_X1 U6362 ( .B1(n6476), .B2(n6539), .A(n5159), .ZN(n5160) );
  AOI21_X1 U6363 ( .B1(n6514), .B2(n5167), .A(n5160), .ZN(n5161) );
  OAI21_X1 U6364 ( .B1(n5162), .B2(n5169), .A(n5161), .ZN(U3119) );
  AOI22_X1 U6365 ( .A1(n5164), .A2(n6459), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n5163), .ZN(n5165) );
  OAI21_X1 U6366 ( .B1(n6462), .B2(n6539), .A(n5165), .ZN(n5166) );
  AOI21_X1 U6367 ( .B1(n6502), .B2(n5167), .A(n5166), .ZN(n5168) );
  OAI21_X1 U6368 ( .B1(n5170), .B2(n5169), .A(n5168), .ZN(U3116) );
  AOI21_X1 U6369 ( .B1(n5173), .B2(n5084), .A(n5172), .ZN(n6197) );
  INV_X1 U6370 ( .A(n6197), .ZN(n5187) );
  AOI22_X1 U6371 ( .A1(n5363), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6133), .ZN(n5174) );
  OAI21_X1 U6372 ( .B1(n5187), .B2(n5916), .A(n5174), .ZN(U2880) );
  OAI21_X1 U6373 ( .B1(n5177), .B2(n5176), .A(n5175), .ZN(n5178) );
  INV_X1 U6374 ( .A(n5178), .ZN(n6259) );
  NAND2_X1 U6375 ( .A1(n6259), .A2(n6224), .ZN(n5182) );
  AND2_X1 U6376 ( .A1(n6317), .A2(REIP_REG_8__SCAN_IN), .ZN(n6257) );
  NOR2_X1 U6377 ( .A1(n6228), .A2(n5179), .ZN(n5180) );
  AOI211_X1 U6378 ( .C1(n6218), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6257), 
        .B(n5180), .ZN(n5181) );
  OAI211_X1 U6379 ( .C1(n6211), .C2(n5183), .A(n5182), .B(n5181), .ZN(U2978)
         );
  INV_X1 U6380 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5186) );
  OAI21_X1 U6381 ( .B1(n5185), .B2(n5184), .A(n5241), .ZN(n5345) );
  OAI222_X1 U6382 ( .A1(n5187), .A2(n5456), .B1(n5186), .B2(n7016), .C1(n7014), 
        .C2(n5345), .ZN(U2848) );
  NOR2_X1 U6383 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5188), .ZN(n5232)
         );
  NAND2_X1 U6384 ( .A1(n6454), .A2(n6674), .ZN(n6371) );
  OAI22_X1 U6385 ( .A1(n6371), .A2(n5190), .B1(n5189), .B2(n6455), .ZN(n5226)
         );
  NAND2_X1 U6386 ( .A1(n6520), .A2(n5226), .ZN(n5199) );
  NOR2_X2 U6387 ( .A1(n5191), .A2(n6409), .ZN(n6361) );
  AOI211_X1 U6388 ( .C1(n6361), .C2(n6374), .A(n5193), .B(n5192), .ZN(n5194)
         );
  NOR3_X1 U6389 ( .A1(n5196), .A2(n5195), .A3(n5194), .ZN(n5197) );
  OAI21_X1 U6390 ( .B1(n5232), .B2(n6662), .A(n5197), .ZN(n5227) );
  AOI22_X1 U6391 ( .A1(n6361), .A2(n6518), .B1(INSTQUEUE_REG_4__4__SCAN_IN), 
        .B2(n5227), .ZN(n5198) );
  OAI211_X1 U6392 ( .C1(n5230), .C2(n6523), .A(n5199), .B(n5198), .ZN(n5200)
         );
  AOI21_X1 U6393 ( .B1(n6519), .B2(n5232), .A(n5200), .ZN(n5201) );
  INV_X1 U6394 ( .A(n5201), .ZN(U3056) );
  NAND2_X1 U6395 ( .A1(n6508), .A2(n5226), .ZN(n5203) );
  AOI22_X1 U6396 ( .A1(n6361), .A2(n6506), .B1(INSTQUEUE_REG_4__1__SCAN_IN), 
        .B2(n5227), .ZN(n5202) );
  OAI211_X1 U6397 ( .C1(n5230), .C2(n6511), .A(n5203), .B(n5202), .ZN(n5204)
         );
  AOI21_X1 U6398 ( .B1(n6507), .B2(n5232), .A(n5204), .ZN(n5205) );
  INV_X1 U6399 ( .A(n5205), .ZN(U3053) );
  NAND2_X1 U6400 ( .A1(n6535), .A2(n5226), .ZN(n5207) );
  AOI22_X1 U6401 ( .A1(n6361), .A2(n6531), .B1(INSTQUEUE_REG_4__7__SCAN_IN), 
        .B2(n5227), .ZN(n5206) );
  OAI211_X1 U6402 ( .C1(n5230), .C2(n6540), .A(n5207), .B(n5206), .ZN(n5208)
         );
  AOI21_X1 U6403 ( .B1(n6533), .B2(n5232), .A(n5208), .ZN(n5209) );
  INV_X1 U6404 ( .A(n5209), .ZN(U3059) );
  NAND2_X1 U6405 ( .A1(n6468), .A2(n5226), .ZN(n5211) );
  AOI22_X1 U6406 ( .A1(n6361), .A2(n6423), .B1(INSTQUEUE_REG_4__2__SCAN_IN), 
        .B2(n5227), .ZN(n5210) );
  OAI211_X1 U6407 ( .C1(n5230), .C2(n6388), .A(n5211), .B(n5210), .ZN(n5212)
         );
  AOI21_X1 U6408 ( .B1(n6467), .B2(n5232), .A(n5212), .ZN(n5213) );
  INV_X1 U6409 ( .A(n5213), .ZN(U3054) );
  NAND2_X1 U6410 ( .A1(n6526), .A2(n5226), .ZN(n5215) );
  AOI22_X1 U6411 ( .A1(n6361), .A2(n6524), .B1(INSTQUEUE_REG_4__6__SCAN_IN), 
        .B2(n5227), .ZN(n5214) );
  OAI211_X1 U6412 ( .C1(n5230), .C2(n6529), .A(n5215), .B(n5214), .ZN(n5216)
         );
  AOI21_X1 U6413 ( .B1(n6525), .B2(n5232), .A(n5216), .ZN(n5217) );
  INV_X1 U6414 ( .A(n5217), .ZN(U3058) );
  NAND2_X1 U6415 ( .A1(n6514), .A2(n5226), .ZN(n5219) );
  AOI22_X1 U6416 ( .A1(n6361), .A2(n6512), .B1(INSTQUEUE_REG_4__3__SCAN_IN), 
        .B2(n5227), .ZN(n5218) );
  OAI211_X1 U6417 ( .C1(n5230), .C2(n6517), .A(n5219), .B(n5218), .ZN(n5220)
         );
  AOI21_X1 U6418 ( .B1(n6513), .B2(n5232), .A(n5220), .ZN(n5221) );
  INV_X1 U6419 ( .A(n5221), .ZN(U3055) );
  NAND2_X1 U6420 ( .A1(n6502), .A2(n5226), .ZN(n5223) );
  AOI22_X1 U6421 ( .A1(n6361), .A2(n6500), .B1(INSTQUEUE_REG_4__0__SCAN_IN), 
        .B2(n5227), .ZN(n5222) );
  OAI211_X1 U6422 ( .C1(n5230), .C2(n6505), .A(n5223), .B(n5222), .ZN(n5224)
         );
  AOI21_X1 U6423 ( .B1(n6501), .B2(n5232), .A(n5224), .ZN(n5225) );
  INV_X1 U6424 ( .A(n5225), .ZN(U3052) );
  NAND2_X1 U6425 ( .A1(n6482), .A2(n5226), .ZN(n5229) );
  AOI22_X1 U6426 ( .A1(n6361), .A2(n6433), .B1(INSTQUEUE_REG_4__5__SCAN_IN), 
        .B2(n5227), .ZN(n5228) );
  OAI211_X1 U6427 ( .C1(n5230), .C2(n6395), .A(n5229), .B(n5228), .ZN(n5231)
         );
  AOI21_X1 U6428 ( .B1(n6481), .B2(n5232), .A(n5231), .ZN(n5233) );
  INV_X1 U6429 ( .A(n5233), .ZN(U3057) );
  INV_X1 U6430 ( .A(n5234), .ZN(n5237) );
  INV_X1 U6431 ( .A(n5172), .ZN(n5236) );
  AOI21_X1 U6432 ( .B1(n5237), .B2(n5236), .A(n5235), .ZN(n5357) );
  INV_X1 U6433 ( .A(n5357), .ZN(n5269) );
  AOI22_X1 U6434 ( .A1(n5363), .A2(DATAI_12_), .B1(EAX_REG_12__SCAN_IN), .B2(
        n6133), .ZN(n5238) );
  OAI21_X1 U6435 ( .B1(n5269), .B2(n5916), .A(n5238), .ZN(U2879) );
  INV_X1 U6436 ( .A(n5239), .ZN(n5257) );
  NAND2_X1 U6437 ( .A1(n5241), .A2(n5240), .ZN(n5242) );
  NAND2_X1 U6438 ( .A1(n5257), .A2(n5242), .ZN(n6229) );
  INV_X1 U6439 ( .A(n6229), .ZN(n5243) );
  AOI22_X1 U6440 ( .A1(n6124), .A2(n5243), .B1(n5454), .B2(EBX_REG_12__SCAN_IN), .ZN(n5244) );
  OAI21_X1 U6441 ( .B1(n5269), .B2(n5456), .A(n5244), .ZN(U2847) );
  NAND2_X1 U6442 ( .A1(n5246), .A2(n5245), .ZN(n5247) );
  XNOR2_X1 U6443 ( .A(n5248), .B(n5247), .ZN(n6253) );
  INV_X1 U6444 ( .A(n6253), .ZN(n5253) );
  AOI22_X1 U6445 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6317), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5249) );
  OAI21_X1 U6446 ( .B1(n5250), .B2(n6228), .A(n5249), .ZN(n5251) );
  AOI21_X1 U6447 ( .B1(n6054), .B2(n6223), .A(n5251), .ZN(n5252) );
  OAI21_X1 U6448 ( .B1(n5253), .B2(n6213), .A(n5252), .ZN(U2977) );
  OAI21_X1 U6449 ( .B1(n5235), .B2(n5255), .A(n5254), .ZN(n5596) );
  AOI22_X1 U6450 ( .A1(n5363), .A2(DATAI_13_), .B1(EAX_REG_13__SCAN_IN), .B2(
        n6133), .ZN(n5256) );
  OAI21_X1 U6451 ( .B1(n5596), .B2(n5916), .A(n5256), .ZN(U2878) );
  AOI21_X1 U6452 ( .B1(n5258), .B2(n5257), .A(n5332), .ZN(n5975) );
  AOI22_X1 U6453 ( .A1(n5975), .A2(n6124), .B1(EBX_REG_13__SCAN_IN), .B2(n5454), .ZN(n5259) );
  OAI21_X1 U6454 ( .B1(n5596), .B2(n5456), .A(n5259), .ZN(U2846) );
  NOR2_X1 U6455 ( .A1(n6092), .A2(n5260), .ZN(n6029) );
  NOR2_X1 U6456 ( .A1(n6029), .A2(n6095), .ZN(n6033) );
  INV_X1 U6457 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6628) );
  NOR2_X1 U6458 ( .A1(n6033), .A2(n6628), .ZN(n5267) );
  OAI22_X1 U6459 ( .A1(n5261), .A2(n6109), .B1(n6104), .B2(n6229), .ZN(n5266)
         );
  AND2_X1 U6460 ( .A1(n6110), .A2(EBX_REG_12__SCAN_IN), .ZN(n5265) );
  OR3_X1 U6461 ( .A1(n6092), .A2(REIP_REG_12__SCAN_IN), .A3(n5262), .ZN(n5263)
         );
  OAI211_X1 U6462 ( .C1(n6108), .C2(n5355), .A(n5263), .B(n6067), .ZN(n5264)
         );
  NOR4_X1 U6463 ( .A1(n5267), .A2(n5266), .A3(n5265), .A4(n5264), .ZN(n5268)
         );
  OAI21_X1 U6464 ( .B1(n5269), .B2(n6044), .A(n5268), .ZN(U2815) );
  INV_X1 U6465 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6629) );
  AOI22_X1 U6466 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6110), .B1(n5270), .B2(n6629), .ZN(n5271) );
  OAI211_X1 U6467 ( .C1(n6109), .C2(n5272), .A(n5271), .B(n6067), .ZN(n5273)
         );
  AOI21_X1 U6468 ( .B1(n5593), .B2(n6096), .A(n5273), .ZN(n5277) );
  NOR2_X1 U6469 ( .A1(n5901), .A2(n5274), .ZN(n5275) );
  AOI22_X1 U6470 ( .A1(n5275), .A2(REIP_REG_13__SCAN_IN), .B1(n6107), .B2(
        n5975), .ZN(n5276) );
  OAI211_X1 U6471 ( .C1(n5596), .C2(n6044), .A(n5277), .B(n5276), .ZN(U2814)
         );
  OR2_X1 U6472 ( .A1(n5282), .A2(n6530), .ZN(n5278) );
  AOI21_X1 U6473 ( .B1(n5278), .B2(STATEBS16_REG_SCAN_IN), .A(n6694), .ZN(
        n5286) );
  NOR3_X1 U6474 ( .A1(n6448), .A2(n6681), .A3(n5279), .ZN(n5280) );
  NOR2_X1 U6475 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5281), .ZN(n5315)
         );
  INV_X1 U6476 ( .A(n5283), .ZN(n5285) );
  INV_X1 U6477 ( .A(n5315), .ZN(n5284) );
  AOI22_X1 U6478 ( .A1(n5286), .A2(n5285), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5284), .ZN(n5288) );
  NAND4_X1 U6479 ( .A1(n5289), .A2(n5288), .A3(n5287), .A4(n6455), .ZN(n5311)
         );
  AOI22_X1 U6480 ( .A1(n6530), .A2(n6469), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5311), .ZN(n5290) );
  OAI21_X1 U6481 ( .B1(n5313), .B2(n6472), .A(n5290), .ZN(n5291) );
  AOI21_X1 U6482 ( .B1(n6467), .B2(n5315), .A(n5291), .ZN(n5292) );
  OAI21_X1 U6483 ( .B1(n5317), .B2(n6426), .A(n5292), .ZN(U3102) );
  AOI22_X1 U6484 ( .A1(n6530), .A2(n6493), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5311), .ZN(n5293) );
  OAI21_X1 U6485 ( .B1(n5313), .B2(n6499), .A(n5293), .ZN(n5294) );
  AOI21_X1 U6486 ( .B1(n6533), .B2(n5315), .A(n5294), .ZN(n5295) );
  OAI21_X1 U6487 ( .B1(n5317), .B2(n6445), .A(n5295), .ZN(U3107) );
  AOI22_X1 U6488 ( .A1(n6530), .A2(n6487), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5311), .ZN(n5296) );
  OAI21_X1 U6489 ( .B1(n5313), .B2(n6490), .A(n5296), .ZN(n5297) );
  AOI21_X1 U6490 ( .B1(n6525), .B2(n5315), .A(n5297), .ZN(n5298) );
  OAI21_X1 U6491 ( .B1(n5317), .B2(n6439), .A(n5298), .ZN(U3106) );
  AOI22_X1 U6492 ( .A1(n6530), .A2(n6477), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5311), .ZN(n5299) );
  OAI21_X1 U6493 ( .B1(n5313), .B2(n6480), .A(n5299), .ZN(n5300) );
  AOI21_X1 U6494 ( .B1(n6519), .B2(n5315), .A(n5300), .ZN(n5301) );
  OAI21_X1 U6495 ( .B1(n5317), .B2(n6432), .A(n5301), .ZN(U3104) );
  AOI22_X1 U6496 ( .A1(n6530), .A2(n6483), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5311), .ZN(n5302) );
  OAI21_X1 U6497 ( .B1(n5313), .B2(n6486), .A(n5302), .ZN(n5303) );
  AOI21_X1 U6498 ( .B1(n6481), .B2(n5315), .A(n5303), .ZN(n5304) );
  OAI21_X1 U6499 ( .B1(n5317), .B2(n6436), .A(n5304), .ZN(U3105) );
  AOI22_X1 U6500 ( .A1(n6530), .A2(n6473), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5311), .ZN(n5305) );
  OAI21_X1 U6501 ( .B1(n5313), .B2(n6476), .A(n5305), .ZN(n5306) );
  AOI21_X1 U6502 ( .B1(n6513), .B2(n5315), .A(n5306), .ZN(n5307) );
  OAI21_X1 U6503 ( .B1(n5317), .B2(n6429), .A(n5307), .ZN(U3103) );
  AOI22_X1 U6504 ( .A1(n6530), .A2(n6459), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5311), .ZN(n5308) );
  OAI21_X1 U6505 ( .B1(n5313), .B2(n6462), .A(n5308), .ZN(n5309) );
  AOI21_X1 U6506 ( .B1(n6501), .B2(n5315), .A(n5309), .ZN(n5310) );
  OAI21_X1 U6507 ( .B1(n5317), .B2(n6419), .A(n5310), .ZN(U3100) );
  AOI22_X1 U6508 ( .A1(n6530), .A2(n6463), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5311), .ZN(n5312) );
  OAI21_X1 U6509 ( .B1(n5313), .B2(n6466), .A(n5312), .ZN(n5314) );
  AOI21_X1 U6510 ( .B1(n6507), .B2(n5315), .A(n5314), .ZN(n5316) );
  OAI21_X1 U6511 ( .B1(n5317), .B2(n6422), .A(n5316), .ZN(U3101) );
  XNOR2_X1 U6512 ( .A(n5554), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5319)
         );
  XNOR2_X1 U6513 ( .A(n5318), .B(n5319), .ZN(n6247) );
  INV_X1 U6514 ( .A(n6247), .ZN(n5324) );
  AOI22_X1 U6515 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6317), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5320) );
  OAI21_X1 U6516 ( .B1(n6043), .B2(n6228), .A(n5320), .ZN(n5321) );
  AOI21_X1 U6517 ( .B1(n5322), .B2(n6223), .A(n5321), .ZN(n5323) );
  OAI21_X1 U6518 ( .B1(n5324), .B2(n6213), .A(n5323), .ZN(U2976) );
  AOI21_X1 U6519 ( .B1(n5326), .B2(n5254), .A(n3858), .ZN(n5587) );
  INV_X1 U6520 ( .A(n5587), .ZN(n5339) );
  AOI22_X1 U6521 ( .A1(n5363), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6133), .ZN(n5327) );
  OAI21_X1 U6522 ( .B1(n5339), .B2(n5916), .A(n5327), .ZN(U2877) );
  AND2_X1 U6523 ( .A1(n6105), .A2(n5328), .ZN(n6022) );
  NAND2_X1 U6524 ( .A1(n6883), .A2(n5329), .ZN(n5337) );
  NAND2_X1 U6525 ( .A1(n6110), .A2(EBX_REG_14__SCAN_IN), .ZN(n5330) );
  OAI211_X1 U6526 ( .C1(n6108), .C2(n5585), .A(n5330), .B(n6067), .ZN(n5336)
         );
  INV_X1 U6527 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5334) );
  OR2_X1 U6528 ( .A1(n5332), .A2(n5331), .ZN(n5333) );
  NAND2_X1 U6529 ( .A1(n5739), .A2(n5333), .ZN(n5758) );
  OAI22_X1 U6530 ( .A1(n5334), .A2(n6109), .B1(n6104), .B2(n5758), .ZN(n5335)
         );
  AOI211_X1 U6531 ( .C1(n6022), .C2(n5337), .A(n5336), .B(n5335), .ZN(n5338)
         );
  OAI21_X1 U6532 ( .B1(n5339), .B2(n6044), .A(n5338), .ZN(U2813) );
  OAI222_X1 U6533 ( .A1(n5339), .A2(n5456), .B1(n7016), .B2(n4278), .C1(n5758), 
        .C2(n7014), .ZN(U2845) );
  AOI22_X1 U6534 ( .A1(n5341), .A2(n5554), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5318), .ZN(n5343) );
  XNOR2_X1 U6535 ( .A(n5554), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5342)
         );
  XNOR2_X1 U6536 ( .A(n5343), .B(n5342), .ZN(n6200) );
  NAND2_X1 U6537 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n5751), .ZN(n6232) );
  OAI21_X1 U6538 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5344), .A(n6232), 
        .ZN(n5347) );
  INV_X1 U6539 ( .A(n5345), .ZN(n6031) );
  AOI22_X1 U6540 ( .A1(n5611), .A2(n6031), .B1(n6317), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5346) );
  OAI211_X1 U6541 ( .C1(n6200), .C2(n5745), .A(n5347), .B(n5346), .ZN(U3007)
         );
  CLKBUF_X1 U6542 ( .A(n5348), .Z(n5353) );
  INV_X1 U6543 ( .A(n5349), .ZN(n5351) );
  NAND2_X1 U6544 ( .A1(n5351), .A2(n5350), .ZN(n5352) );
  XNOR2_X1 U6545 ( .A(n5353), .B(n5352), .ZN(n6231) );
  INV_X1 U6546 ( .A(n6231), .ZN(n5359) );
  AOI22_X1 U6547 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .B1(n6317), 
        .B2(REIP_REG_12__SCAN_IN), .ZN(n5354) );
  OAI21_X1 U6548 ( .B1(n5355), .B2(n6228), .A(n5354), .ZN(n5356) );
  AOI21_X1 U6549 ( .B1(n5357), .B2(n6223), .A(n5356), .ZN(n5358) );
  OAI21_X1 U6550 ( .B1(n5359), .B2(n6213), .A(n5358), .ZN(U2974) );
  INV_X1 U6551 ( .A(n5360), .ZN(n5361) );
  AOI21_X1 U6552 ( .B1(n5362), .B2(n5325), .A(n5361), .ZN(n6120) );
  INV_X1 U6553 ( .A(n6120), .ZN(n5365) );
  AOI22_X1 U6554 ( .A1(n5363), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6133), .ZN(n5364) );
  OAI21_X1 U6555 ( .B1(n5365), .B2(n5916), .A(n5364), .ZN(U2876) );
  AOI21_X1 U6556 ( .B1(n5368), .B2(n5360), .A(n5367), .ZN(n5369) );
  INV_X1 U6557 ( .A(n5369), .ZN(n5574) );
  INV_X1 U6558 ( .A(n5370), .ZN(n5373) );
  NOR2_X1 U6559 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5373), .ZN(n6025) );
  AOI22_X1 U6560 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6110), .B1(n5571), .B2(n6096), .ZN(n5371) );
  OAI211_X1 U6561 ( .C1(n6109), .C2(n5569), .A(n5371), .B(n6067), .ZN(n5372)
         );
  AOI221_X1 U6562 ( .B1(n6022), .B2(REIP_REG_16__SCAN_IN), .C1(n6025), .C2(
        REIP_REG_16__SCAN_IN), .A(n5372), .ZN(n5375) );
  INV_X1 U6563 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6977) );
  NOR2_X1 U6564 ( .A1(n5373), .A2(n6977), .ZN(n6013) );
  INV_X1 U6565 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6633) );
  XNOR2_X1 U6566 ( .A(n5737), .B(n5724), .ZN(n5962) );
  AOI22_X1 U6567 ( .A1(n6013), .A2(n6633), .B1(n6107), .B2(n5962), .ZN(n5374)
         );
  OAI211_X1 U6568 ( .C1(n5574), .C2(n6044), .A(n5375), .B(n5374), .ZN(U2811)
         );
  AOI22_X1 U6569 ( .A1(n6130), .A2(DATAI_16_), .B1(n6133), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6570 ( .A1(n6134), .A2(DATAI_0_), .ZN(n5376) );
  OAI211_X1 U6571 ( .C1(n5574), .C2(n5916), .A(n5377), .B(n5376), .ZN(U2875)
         );
  INV_X1 U6572 ( .A(n5962), .ZN(n5378) );
  OAI222_X1 U6573 ( .A1(n5574), .A2(n5456), .B1(n5379), .B2(n7016), .C1(n7014), 
        .C2(n5378), .ZN(U2843) );
  INV_X1 U6574 ( .A(n5380), .ZN(n5382) );
  NOR2_X1 U6575 ( .A1(n5382), .A2(n5381), .ZN(n5384) );
  NOR3_X1 U6576 ( .A1(n5387), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n6577), 
        .ZN(n5383) );
  AOI211_X1 U6577 ( .C1(n5385), .C2(n5981), .A(n5384), .B(n5383), .ZN(n5390)
         );
  AOI21_X1 U6578 ( .B1(n5387), .B2(n5386), .A(n6664), .ZN(n5389) );
  OAI22_X1 U6579 ( .A1(n5390), .A2(n6664), .B1(n5389), .B2(n5388), .ZN(U3459)
         );
  AOI22_X1 U6580 ( .A1(n5618), .A2(n6124), .B1(EBX_REG_30__SCAN_IN), .B2(n5454), .ZN(n5392) );
  OAI21_X1 U6581 ( .B1(n5391), .B2(n5456), .A(n5392), .ZN(U2829) );
  AOI22_X1 U6582 ( .A1(n6134), .A2(DATAI_14_), .B1(n6133), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5394) );
  NAND2_X1 U6583 ( .A1(n6130), .A2(DATAI_30_), .ZN(n5393) );
  OAI211_X1 U6584 ( .C1(n5391), .C2(n5916), .A(n5394), .B(n5393), .ZN(U2861)
         );
  NAND2_X1 U6585 ( .A1(n5396), .A2(n5395), .ZN(n5398) );
  AOI22_X1 U6586 ( .A1(n6130), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6133), .ZN(n5397) );
  OAI21_X1 U6587 ( .B1(n5419), .B2(n5398), .A(n5397), .ZN(U2860) );
  INV_X1 U6588 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6768) );
  NAND3_X1 U6589 ( .A1(REIP_REG_30__SCAN_IN), .A2(n5399), .A3(n6768), .ZN(
        n5418) );
  NAND2_X1 U6590 ( .A1(n4416), .A2(n5431), .ZN(n5426) );
  NAND2_X1 U6591 ( .A1(n5430), .A2(n5402), .ZN(n5405) );
  INV_X1 U6592 ( .A(n5403), .ZN(n5404) );
  NAND2_X1 U6593 ( .A1(n5405), .A2(n5404), .ZN(n5410) );
  OAI22_X1 U6594 ( .A1(n5407), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5406), .B2(EBX_REG_31__SCAN_IN), .ZN(n5408) );
  INV_X1 U6595 ( .A(n5408), .ZN(n5409) );
  XNOR2_X1 U6596 ( .A(n5410), .B(n5409), .ZN(n5420) );
  NOR3_X1 U6597 ( .A1(n5411), .A2(n5901), .A3(n6768), .ZN(n5416) );
  NAND2_X1 U6598 ( .A1(EBX_REG_31__SCAN_IN), .A2(n5412), .ZN(n5414) );
  OAI22_X1 U6599 ( .A1(n6109), .A2(n6835), .B1(n5414), .B2(n5413), .ZN(n5415)
         );
  AOI211_X1 U6600 ( .C1(n5420), .C2(n6107), .A(n5416), .B(n5415), .ZN(n5417)
         );
  OAI211_X1 U6601 ( .C1(n5419), .C2(n6044), .A(n5418), .B(n5417), .ZN(U2796)
         );
  INV_X1 U6602 ( .A(n5420), .ZN(n5597) );
  OAI22_X1 U6603 ( .A1(n5597), .A2(n7014), .B1(n5421), .B2(n7016), .ZN(U2828)
         );
  AND2_X1 U6604 ( .A1(n5435), .A2(n5422), .ZN(n5424) );
  NAND2_X1 U6605 ( .A1(n5425), .A2(n5683), .ZN(n5427) );
  NAND2_X1 U6606 ( .A1(n5427), .A2(n5426), .ZN(n5428) );
  NOR2_X1 U6607 ( .A1(n3117), .A2(n5428), .ZN(n5429) );
  OAI222_X1 U6608 ( .A1(n5456), .A2(n5811), .B1(n5431), .B2(n7016), .C1(n5810), 
        .C2(n7014), .ZN(U2830) );
  NAND2_X1 U6609 ( .A1(n3112), .A2(n5433), .ZN(n5434) );
  NOR2_X1 U6610 ( .A1(n5639), .A2(n5436), .ZN(n5437) );
  OR2_X1 U6611 ( .A1(n3117), .A2(n5437), .ZN(n5818) );
  OAI22_X1 U6612 ( .A1(n5818), .A2(n7014), .B1(n6761), .B2(n7016), .ZN(n5438)
         );
  INV_X1 U6613 ( .A(n5438), .ZN(n5439) );
  OAI21_X1 U6614 ( .B1(n5491), .B2(n5456), .A(n5439), .ZN(U2831) );
  OAI21_X1 U6615 ( .B1(n5441), .B2(n5443), .A(n5442), .ZN(n5836) );
  NAND2_X1 U6616 ( .A1(n5453), .A2(n5444), .ZN(n5445) );
  NAND2_X1 U6617 ( .A1(n3121), .A2(n5445), .ZN(n5835) );
  INV_X1 U6618 ( .A(n5835), .ZN(n5446) );
  AOI22_X1 U6619 ( .A1(n5446), .A2(n6124), .B1(EBX_REG_26__SCAN_IN), .B2(n5454), .ZN(n5447) );
  OAI21_X1 U6620 ( .B1(n5836), .B2(n5456), .A(n5447), .ZN(U2833) );
  INV_X1 U6621 ( .A(n5448), .ZN(n5450) );
  INV_X1 U6622 ( .A(n4373), .ZN(n5449) );
  AOI21_X1 U6623 ( .B1(n5450), .B2(n5449), .A(n5441), .ZN(n5937) );
  INV_X1 U6624 ( .A(n5937), .ZN(n5457) );
  NAND2_X1 U6625 ( .A1(n4408), .A2(n5451), .ZN(n5452) );
  AND2_X1 U6626 ( .A1(n5453), .A2(n5452), .ZN(n5957) );
  AOI22_X1 U6627 ( .A1(n5957), .A2(n6124), .B1(EBX_REG_25__SCAN_IN), .B2(n5454), .ZN(n5455) );
  OAI21_X1 U6628 ( .B1(n5457), .B2(n5456), .A(n5455), .ZN(U2834) );
  OAI22_X1 U6629 ( .A1(n5859), .A2(n7014), .B1(n5458), .B2(n7016), .ZN(n5459)
         );
  INV_X1 U6630 ( .A(n5459), .ZN(n5460) );
  OAI21_X1 U6631 ( .B1(n5855), .B2(n5456), .A(n5460), .ZN(U2835) );
  NAND2_X1 U6632 ( .A1(n5461), .A2(n5462), .ZN(n5463) );
  AND2_X1 U6633 ( .A1(n4371), .A2(n5463), .ZN(n5922) );
  XNOR2_X1 U6634 ( .A(n5474), .B(n5464), .ZN(n5861) );
  OAI22_X1 U6635 ( .A1(n5861), .A2(n7014), .B1(n5465), .B2(n7016), .ZN(n5466)
         );
  AOI21_X1 U6636 ( .B1(n5922), .B2(n6125), .A(n5466), .ZN(n5467) );
  INV_X1 U6637 ( .A(n5467), .ZN(U2836) );
  OR2_X1 U6638 ( .A1(n5468), .A2(n5469), .ZN(n5470) );
  NAND2_X1 U6639 ( .A1(n5461), .A2(n5470), .ZN(n5871) );
  INV_X1 U6640 ( .A(n5871), .ZN(n5925) );
  NAND2_X1 U6641 ( .A1(n5471), .A2(n5472), .ZN(n5473) );
  NAND2_X1 U6642 ( .A1(n5474), .A2(n5473), .ZN(n5870) );
  OAI22_X1 U6643 ( .A1(n5870), .A2(n7014), .B1(n6888), .B2(n7016), .ZN(n5475)
         );
  AOI21_X1 U6644 ( .B1(n5925), .B2(n6125), .A(n5475), .ZN(n5476) );
  INV_X1 U6645 ( .A(n5476), .ZN(U2837) );
  INV_X1 U6646 ( .A(n5549), .ZN(n5478) );
  NAND2_X1 U6647 ( .A1(n3110), .A2(n5478), .ZN(n5479) );
  AOI21_X1 U6648 ( .B1(n5480), .B2(n5479), .A(n5468), .ZN(n5928) );
  OR2_X1 U6649 ( .A1(n5482), .A2(n5481), .ZN(n5483) );
  NAND2_X1 U6650 ( .A1(n5471), .A2(n5483), .ZN(n5884) );
  OAI22_X1 U6651 ( .A1(n5884), .A2(n7014), .B1(n5484), .B2(n7016), .ZN(n5485)
         );
  AOI21_X1 U6652 ( .B1(n5928), .B2(n6125), .A(n5485), .ZN(n5486) );
  INV_X1 U6653 ( .A(n5486), .ZN(U2838) );
  AOI22_X1 U6654 ( .A1(n6134), .A2(DATAI_13_), .B1(n6133), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5488) );
  NAND2_X1 U6655 ( .A1(n6130), .A2(DATAI_29_), .ZN(n5487) );
  OAI211_X1 U6656 ( .C1(n5811), .C2(n5916), .A(n5488), .B(n5487), .ZN(U2862)
         );
  AOI22_X1 U6657 ( .A1(n6134), .A2(DATAI_12_), .B1(n6133), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6658 ( .A1(n6130), .A2(DATAI_28_), .ZN(n5489) );
  OAI211_X1 U6659 ( .C1(n5491), .C2(n5916), .A(n5490), .B(n5489), .ZN(U2863)
         );
  AOI22_X1 U6660 ( .A1(n6134), .A2(DATAI_10_), .B1(n6133), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6661 ( .A1(n6130), .A2(DATAI_26_), .ZN(n5492) );
  OAI211_X1 U6662 ( .C1(n5836), .C2(n5916), .A(n5493), .B(n5492), .ZN(U2865)
         );
  AOI22_X1 U6663 ( .A1(n6134), .A2(DATAI_8_), .B1(n6133), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U6664 ( .A1(n6130), .A2(DATAI_24_), .ZN(n5494) );
  OAI211_X1 U6665 ( .C1(n5855), .C2(n5916), .A(n5495), .B(n5494), .ZN(U2867)
         );
  INV_X1 U6666 ( .A(n5811), .ZN(n5501) );
  NAND2_X1 U6667 ( .A1(n6317), .A2(REIP_REG_29__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6668 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5499)
         );
  OAI211_X1 U6669 ( .C1(n6228), .C2(n5808), .A(n5627), .B(n5499), .ZN(n5500)
         );
  AOI21_X1 U6670 ( .B1(n5501), .B2(n6223), .A(n5500), .ZN(n5502) );
  OAI21_X1 U6671 ( .B1(n5631), .B2(n6213), .A(n5502), .ZN(U2957) );
  NOR3_X1 U6672 ( .A1(n4381), .A2(n5554), .A3(n6843), .ZN(n5504) );
  NAND2_X1 U6673 ( .A1(n6788), .A2(n5520), .ZN(n5651) );
  NOR3_X1 U6674 ( .A1(n5503), .A2(n5582), .A3(n5651), .ZN(n5511) );
  OAI22_X1 U6675 ( .A1(n5504), .A2(n5511), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n6843), .ZN(n5506) );
  XNOR2_X1 U6676 ( .A(n5506), .B(n5505), .ZN(n5638) );
  NOR2_X1 U6677 ( .A1(n6292), .A2(n6807), .ZN(n5632) );
  AOI21_X1 U6678 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5632), 
        .ZN(n5507) );
  OAI21_X1 U6679 ( .B1(n5508), .B2(n6228), .A(n5507), .ZN(n5509) );
  AOI21_X1 U6680 ( .B1(n5820), .B2(n6223), .A(n5509), .ZN(n5510) );
  OAI21_X1 U6681 ( .B1(n5638), .B2(n6213), .A(n5510), .ZN(U2958) );
  INV_X1 U6682 ( .A(n5511), .ZN(n5513) );
  NAND2_X1 U6683 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  XNOR2_X1 U6684 ( .A(n5514), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5649)
         );
  NAND2_X1 U6685 ( .A1(n5442), .A2(n5515), .ZN(n5516) );
  AND2_X1 U6686 ( .A1(n3112), .A2(n5516), .ZN(n5917) );
  NAND2_X1 U6687 ( .A1(n6317), .A2(REIP_REG_27__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U6688 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5517)
         );
  OAI211_X1 U6689 ( .C1(n6228), .C2(n5827), .A(n5643), .B(n5517), .ZN(n5518)
         );
  AOI21_X1 U6690 ( .B1(n5917), .B2(n6223), .A(n5518), .ZN(n5519) );
  OAI21_X1 U6691 ( .B1(n5649), .B2(n6213), .A(n5519), .ZN(U2959) );
  XNOR2_X1 U6692 ( .A(n5582), .B(n5520), .ZN(n5521) );
  XNOR2_X1 U6693 ( .A(n4381), .B(n5521), .ZN(n5655) );
  NAND2_X1 U6694 ( .A1(n6317), .A2(REIP_REG_26__SCAN_IN), .ZN(n5653) );
  OAI21_X1 U6695 ( .B1(n5955), .B2(n5522), .A(n5653), .ZN(n5524) );
  NOR2_X1 U6696 ( .A1(n5836), .A2(n5564), .ZN(n5523) );
  OAI21_X1 U6697 ( .B1(n6213), .B2(n5655), .A(n5525), .ZN(U2960) );
  NAND2_X1 U6698 ( .A1(n3602), .A2(n5526), .ZN(n5528) );
  OAI21_X1 U6699 ( .B1(n5529), .B2(n5528), .A(n5527), .ZN(n5530) );
  XNOR2_X1 U6700 ( .A(n5530), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5665)
         );
  NAND2_X1 U6701 ( .A1(n6317), .A2(REIP_REG_23__SCAN_IN), .ZN(n5660) );
  NAND2_X1 U6702 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5531)
         );
  OAI211_X1 U6703 ( .C1(n6228), .C2(n5867), .A(n5660), .B(n5531), .ZN(n5532)
         );
  AOI21_X1 U6704 ( .B1(n5922), .B2(n6223), .A(n5532), .ZN(n5533) );
  OAI21_X1 U6705 ( .B1(n5665), .B2(n6213), .A(n5533), .ZN(U2963) );
  AOI21_X1 U6706 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5582), .A(n5534), 
        .ZN(n5536) );
  XOR2_X1 U6707 ( .A(n5536), .B(n5535), .Z(n5673) );
  NAND2_X1 U6708 ( .A1(n6317), .A2(REIP_REG_22__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U6709 ( .B1(n5955), .B2(n6841), .A(n5667), .ZN(n5538) );
  NOR2_X1 U6710 ( .A1(n5871), .A2(n5564), .ZN(n5537) );
  AOI211_X1 U6711 ( .C1(n6196), .C2(n5869), .A(n5538), .B(n5537), .ZN(n5539)
         );
  OAI21_X1 U6712 ( .B1(n5673), .B2(n6213), .A(n5539), .ZN(U2964) );
  AOI21_X1 U6713 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5680) );
  INV_X1 U6714 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5543) );
  NOR2_X1 U6715 ( .A1(n6292), .A2(n5543), .ZN(n5676) );
  AOI21_X1 U6716 ( .B1(n6218), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5676), 
        .ZN(n5544) );
  OAI21_X1 U6717 ( .B1(n5879), .B2(n6228), .A(n5544), .ZN(n5545) );
  AOI21_X1 U6718 ( .B1(n5928), .B2(n6223), .A(n5545), .ZN(n5546) );
  OAI21_X1 U6719 ( .B1(n5680), .B2(n6213), .A(n5546), .ZN(U2965) );
  XOR2_X1 U6720 ( .A(n5548), .B(n5547), .Z(n5693) );
  XNOR2_X1 U6721 ( .A(n3110), .B(n5549), .ZN(n5931) );
  INV_X1 U6722 ( .A(n5889), .ZN(n5551) );
  NAND2_X1 U6723 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5550)
         );
  NAND2_X1 U6724 ( .A1(n6317), .A2(REIP_REG_20__SCAN_IN), .ZN(n5686) );
  OAI211_X1 U6725 ( .C1(n6228), .C2(n5551), .A(n5550), .B(n5686), .ZN(n5552)
         );
  AOI21_X1 U6726 ( .B1(n5931), .B2(n6223), .A(n5552), .ZN(n5553) );
  OAI21_X1 U6727 ( .B1(n5693), .B2(n6213), .A(n5553), .ZN(U2966) );
  NAND2_X1 U6728 ( .A1(n5554), .A2(n5966), .ZN(n5721) );
  NOR2_X1 U6729 ( .A1(n5721), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5557)
         );
  NAND2_X1 U6730 ( .A1(n5582), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5722) );
  NOR3_X1 U6731 ( .A1(n5720), .A2(n5731), .A3(n5722), .ZN(n5556) );
  AOI21_X1 U6732 ( .B1(n5557), .B2(n5720), .A(n5556), .ZN(n5558) );
  XNOR2_X1 U6733 ( .A(n5558), .B(n5716), .ZN(n5719) );
  NAND2_X1 U6734 ( .A1(n6317), .A2(REIP_REG_18__SCAN_IN), .ZN(n5713) );
  OAI21_X1 U6735 ( .B1(n5955), .B2(n5559), .A(n5713), .ZN(n5566) );
  NAND2_X1 U6736 ( .A1(n5561), .A2(n5562), .ZN(n5563) );
  NAND2_X1 U6737 ( .A1(n5560), .A2(n5563), .ZN(n7017) );
  NOR2_X1 U6738 ( .A1(n7017), .A2(n5564), .ZN(n5565) );
  AOI211_X1 U6739 ( .C1(n6196), .C2(n6007), .A(n5566), .B(n5565), .ZN(n5567)
         );
  OAI21_X1 U6740 ( .B1(n5719), .B2(n6213), .A(n5567), .ZN(U2968) );
  NAND2_X1 U6741 ( .A1(n5721), .A2(n5722), .ZN(n5568) );
  XNOR2_X1 U6742 ( .A(n5720), .B(n5568), .ZN(n5963) );
  NAND2_X1 U6743 ( .A1(n5963), .A2(n6224), .ZN(n5573) );
  OAI22_X1 U6744 ( .A1(n5955), .A2(n5569), .B1(n6292), .B2(n6633), .ZN(n5570)
         );
  AOI21_X1 U6745 ( .B1(n6196), .B2(n5571), .A(n5570), .ZN(n5572) );
  OAI211_X1 U6746 ( .C1(n6211), .C2(n5574), .A(n5573), .B(n5572), .ZN(U2970)
         );
  XNOR2_X1 U6747 ( .A(n5582), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5576)
         );
  XNOR2_X1 U6748 ( .A(n5575), .B(n5576), .ZN(n5744) );
  AND2_X1 U6749 ( .A1(n6317), .A2(REIP_REG_15__SCAN_IN), .ZN(n5741) );
  AND2_X1 U6750 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5577)
         );
  AOI211_X1 U6751 ( .C1(n6196), .C2(n6026), .A(n5741), .B(n5577), .ZN(n5579)
         );
  NAND2_X1 U6752 ( .A1(n6120), .A2(n6223), .ZN(n5578) );
  OAI211_X1 U6753 ( .C1(n5744), .C2(n6213), .A(n5579), .B(n5578), .ZN(U2971)
         );
  XNOR2_X1 U6754 ( .A(n5582), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5583)
         );
  XNOR2_X1 U6755 ( .A(n5581), .B(n5583), .ZN(n5761) );
  INV_X1 U6756 ( .A(n5761), .ZN(n5589) );
  NAND2_X1 U6757 ( .A1(n6317), .A2(REIP_REG_14__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U6758 ( .A1(n6218), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5584)
         );
  OAI211_X1 U6759 ( .C1(n6228), .C2(n5585), .A(n5757), .B(n5584), .ZN(n5586)
         );
  AOI21_X1 U6760 ( .B1(n5587), .B2(n6223), .A(n5586), .ZN(n5588) );
  OAI21_X1 U6761 ( .B1(n5589), .B2(n6213), .A(n5588), .ZN(U2972) );
  XNOR2_X1 U6762 ( .A(n5591), .B(n5590), .ZN(n5977) );
  NAND2_X1 U6763 ( .A1(n5977), .A2(n6224), .ZN(n5595) );
  NAND2_X1 U6764 ( .A1(n6317), .A2(REIP_REG_13__SCAN_IN), .ZN(n5973) );
  OAI21_X1 U6765 ( .B1(n5955), .B2(n5272), .A(n5973), .ZN(n5592) );
  AOI21_X1 U6766 ( .B1(n6196), .B2(n5593), .A(n5592), .ZN(n5594) );
  OAI211_X1 U6767 ( .C1(n6211), .C2(n5596), .A(n5595), .B(n5594), .ZN(U2973)
         );
  AND2_X1 U6768 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5604) );
  NAND2_X1 U6769 ( .A1(n5961), .A2(n5599), .ZN(n5620) );
  AND2_X1 U6770 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5650) );
  OR2_X1 U6771 ( .A1(n5599), .A2(n5650), .ZN(n5598) );
  NAND2_X1 U6772 ( .A1(n5961), .A2(n5598), .ZN(n5647) );
  AOI21_X1 U6773 ( .B1(n5602), .B2(n5620), .A(n5647), .ZN(n5619) );
  OAI21_X1 U6774 ( .B1(n5599), .B2(n5604), .A(n5619), .ZN(n5608) );
  INV_X1 U6775 ( .A(n5600), .ZN(n5601) );
  NAND2_X1 U6776 ( .A1(n5956), .A2(n5650), .ZN(n5644) );
  NOR2_X1 U6777 ( .A1(n5644), .A2(n5602), .ZN(n5625) );
  NAND3_X1 U6778 ( .A1(n5625), .A2(n5604), .A3(n5603), .ZN(n5606) );
  OAI21_X1 U6779 ( .B1(n5613), .B2(n5745), .A(n5612), .ZN(U2987) );
  AND3_X1 U6780 ( .A1(n5625), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5614), 
        .ZN(n5617) );
  INV_X1 U6781 ( .A(n5615), .ZN(n5616) );
  AOI211_X2 U6782 ( .C1(n5618), .C2(n5611), .A(n5617), .B(n5616), .ZN(n5622)
         );
  INV_X1 U6783 ( .A(n5619), .ZN(n5629) );
  OAI211_X1 U6784 ( .C1(n5629), .C2(n5624), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5620), .ZN(n5621) );
  OAI211_X1 U6785 ( .C1(n5623), .C2(n5745), .A(n5622), .B(n5621), .ZN(U2988)
         );
  NAND2_X1 U6786 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  OAI211_X1 U6787 ( .C1(n5810), .C2(n6294), .A(n5627), .B(n5626), .ZN(n5628)
         );
  AOI21_X1 U6788 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5629), .A(n5628), 
        .ZN(n5630) );
  OAI21_X1 U6789 ( .B1(n5631), .B2(n5745), .A(n5630), .ZN(U2989) );
  XNOR2_X1 U6790 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5635) );
  INV_X1 U6791 ( .A(n5818), .ZN(n5633) );
  AOI21_X1 U6792 ( .B1(n5633), .B2(n5611), .A(n5632), .ZN(n5634) );
  OAI21_X1 U6793 ( .B1(n5644), .B2(n5635), .A(n5634), .ZN(n5636) );
  AOI21_X1 U6794 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5647), .A(n5636), 
        .ZN(n5637) );
  OAI21_X1 U6795 ( .B1(n5638), .B2(n5745), .A(n5637), .ZN(U2990) );
  INV_X1 U6796 ( .A(n5639), .ZN(n5642) );
  NAND2_X1 U6797 ( .A1(n3121), .A2(n5640), .ZN(n5641) );
  NAND2_X1 U6798 ( .A1(n5642), .A2(n5641), .ZN(n5906) );
  OAI21_X1 U6799 ( .B1(n5906), .B2(n6294), .A(n5643), .ZN(n5646) );
  NOR2_X1 U6800 ( .A1(n5644), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5645)
         );
  AOI211_X1 U6801 ( .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n5647), .A(n5646), .B(n5645), .ZN(n5648) );
  OAI21_X1 U6802 ( .B1(n5649), .B2(n5745), .A(n5648), .ZN(U2991) );
  INV_X1 U6803 ( .A(n5961), .ZN(n5658) );
  INV_X1 U6804 ( .A(n5650), .ZN(n5652) );
  NAND3_X1 U6805 ( .A1(n5956), .A2(n5652), .A3(n5651), .ZN(n5654) );
  OAI211_X1 U6806 ( .C1(n6294), .C2(n5835), .A(n5654), .B(n5653), .ZN(n5657)
         );
  NOR2_X1 U6807 ( .A1(n5655), .A2(n5745), .ZN(n5656) );
  AOI211_X1 U6808 ( .C1(INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n5658), .A(n5657), .B(n5656), .ZN(n5659) );
  INV_X1 U6809 ( .A(n5659), .ZN(U2992) );
  OAI21_X1 U6810 ( .B1(n5861), .B2(n6294), .A(n5660), .ZN(n5662) );
  NOR2_X1 U6811 ( .A1(n5666), .A2(n4182), .ZN(n5661) );
  AOI211_X1 U6812 ( .C1(n5663), .C2(n4182), .A(n5662), .B(n5661), .ZN(n5664)
         );
  OAI21_X1 U6813 ( .B1(n5665), .B2(n5745), .A(n5664), .ZN(U2995) );
  INV_X1 U6814 ( .A(n5666), .ZN(n5671) );
  OAI21_X1 U6815 ( .B1(n5870), .B2(n6294), .A(n5667), .ZN(n5670) );
  NOR2_X1 U6816 ( .A1(n5668), .A2(n6774), .ZN(n5669) );
  AOI211_X1 U6817 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5671), .A(n5670), .B(n5669), .ZN(n5672) );
  OAI21_X1 U6818 ( .B1(n5673), .B2(n5745), .A(n5672), .ZN(U2996) );
  INV_X1 U6819 ( .A(n5884), .ZN(n5677) );
  NOR2_X1 U6820 ( .A1(n5674), .A2(n6774), .ZN(n5675) );
  AOI211_X1 U6821 ( .C1(n5611), .C2(n5677), .A(n5676), .B(n5675), .ZN(n5679)
         );
  NAND3_X1 U6822 ( .A1(n5706), .A2(n5688), .A3(n6774), .ZN(n5678) );
  OAI211_X1 U6823 ( .C1(n5680), .C2(n5745), .A(n5679), .B(n5678), .ZN(U2997)
         );
  MUX2_X1 U6824 ( .A(n5683), .B(n5682), .S(n5681), .Z(n5685) );
  XNOR2_X1 U6825 ( .A(n5685), .B(n5684), .ZN(n5885) );
  OAI21_X1 U6826 ( .B1(n5885), .B2(n6294), .A(n5686), .ZN(n5691) );
  INV_X1 U6827 ( .A(n5706), .ZN(n5689) );
  NOR3_X1 U6828 ( .A1(n5689), .A2(n5688), .A3(n5687), .ZN(n5690) );
  AOI211_X1 U6829 ( .C1(INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n5712), .A(n5691), .B(n5690), .ZN(n5692) );
  OAI21_X1 U6830 ( .B1(n5693), .B2(n5745), .A(n5692), .ZN(U2998) );
  XNOR2_X1 U6831 ( .A(n5695), .B(n5696), .ZN(n5941) );
  INV_X1 U6832 ( .A(n5728), .ZN(n5701) );
  INV_X1 U6833 ( .A(n5697), .ZN(n5699) );
  MUX2_X1 U6834 ( .A(n5700), .B(n5699), .S(n5698), .Z(n5708) );
  NAND2_X1 U6835 ( .A1(n5701), .A2(n5708), .ZN(n5711) );
  XNOR2_X1 U6836 ( .A(n5711), .B(n5702), .ZN(n5912) );
  NAND2_X1 U6837 ( .A1(n5712), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U6838 ( .A1(n6317), .A2(REIP_REG_19__SCAN_IN), .ZN(n5946) );
  OAI211_X1 U6839 ( .C1(n5912), .C2(n6294), .A(n5703), .B(n5946), .ZN(n5704)
         );
  AOI21_X1 U6840 ( .B1(n5706), .B2(n5705), .A(n5704), .ZN(n5707) );
  OAI21_X1 U6841 ( .B1(n5941), .B2(n5745), .A(n5707), .ZN(U2999) );
  INV_X1 U6842 ( .A(n5708), .ZN(n5709) );
  NAND2_X1 U6843 ( .A1(n5728), .A2(n5709), .ZN(n5710) );
  NAND2_X1 U6844 ( .A1(n5711), .A2(n5710), .ZN(n7015) );
  NAND2_X1 U6845 ( .A1(n5712), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5714) );
  OAI211_X1 U6846 ( .C1(n6294), .C2(n7015), .A(n5714), .B(n5713), .ZN(n5715)
         );
  AOI21_X1 U6847 ( .B1(n5717), .B2(n5716), .A(n5715), .ZN(n5718) );
  OAI21_X1 U6848 ( .B1(n5719), .B2(n5745), .A(n5718), .ZN(U3000) );
  MUX2_X1 U6849 ( .A(n5722), .B(n5721), .S(n5720), .Z(n5723) );
  XNOR2_X1 U6850 ( .A(n5723), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5952)
         );
  INV_X1 U6851 ( .A(n5952), .ZN(n5735) );
  INV_X1 U6852 ( .A(n5724), .ZN(n5727) );
  INV_X1 U6853 ( .A(n5725), .ZN(n5726) );
  OAI21_X1 U6854 ( .B1(n5737), .B2(n5727), .A(n5726), .ZN(n5729) );
  AND2_X1 U6855 ( .A1(n5729), .A2(n5728), .ZN(n6117) );
  NAND2_X1 U6856 ( .A1(n6317), .A2(REIP_REG_17__SCAN_IN), .ZN(n5953) );
  OAI221_X1 U6857 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5732), .C1(
        n5731), .C2(n5730), .A(n5953), .ZN(n5733) );
  AOI21_X1 U6858 ( .B1(n6117), .B2(n5611), .A(n5733), .ZN(n5734) );
  OAI21_X1 U6859 ( .B1(n5735), .B2(n5745), .A(n5734), .ZN(U3001) );
  NOR2_X1 U6860 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5736), .ZN(n5965)
         );
  AOI21_X1 U6861 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n5964), .A(n5965), 
        .ZN(n5743) );
  INV_X1 U6862 ( .A(n5737), .ZN(n5738) );
  AOI21_X1 U6863 ( .B1(n5740), .B2(n5739), .A(n5738), .ZN(n6119) );
  AOI21_X1 U6864 ( .B1(n6119), .B2(n5611), .A(n5741), .ZN(n5742) );
  OAI211_X1 U6865 ( .C1(n5744), .C2(n5745), .A(n5743), .B(n5742), .ZN(U3003)
         );
  NOR2_X1 U6866 ( .A1(n6236), .A2(n5748), .ZN(n5756) );
  NAND2_X1 U6867 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5747) );
  NOR2_X1 U6868 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5747), .ZN(n5972)
         );
  AOI22_X1 U6869 ( .A1(n5749), .A2(n5748), .B1(n5747), .B2(n5746), .ZN(n5750)
         );
  NAND2_X1 U6870 ( .A1(n5751), .A2(n5750), .ZN(n5976) );
  AOI221_X1 U6871 ( .B1(n5753), .B2(n5972), .C1(n5752), .C2(n5972), .A(n5976), 
        .ZN(n5754) );
  INV_X1 U6872 ( .A(n5754), .ZN(n5755) );
  MUX2_X1 U6873 ( .A(n5756), .B(n5755), .S(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .Z(n5760) );
  OAI21_X1 U6874 ( .B1(n5758), .B2(n6294), .A(n5757), .ZN(n5759) );
  AOI211_X1 U6875 ( .C1(n5761), .C2(n6315), .A(n5760), .B(n5759), .ZN(n5762)
         );
  INV_X1 U6876 ( .A(n5762), .ZN(U3004) );
  OAI22_X1 U6877 ( .A1(n5764), .A2(n6670), .B1(n5763), .B2(n6577), .ZN(n5765)
         );
  INV_X1 U6878 ( .A(n6664), .ZN(n6668) );
  MUX2_X1 U6879 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5765), .S(n6668), 
        .Z(U3456) );
  NOR2_X1 U6880 ( .A1(n6372), .A2(n5771), .ZN(n5801) );
  INV_X1 U6881 ( .A(n5801), .ZN(n5766) );
  OAI21_X1 U6882 ( .B1(n5767), .B2(n6330), .A(n5766), .ZN(n5770) );
  INV_X1 U6883 ( .A(n5771), .ZN(n5768) );
  INV_X1 U6884 ( .A(n5770), .ZN(n5773) );
  AOI22_X1 U6885 ( .A1(n5773), .A2(n5772), .B1(n5771), .B2(n6694), .ZN(n5774)
         );
  NAND2_X1 U6886 ( .A1(n6414), .A2(n5774), .ZN(n5796) );
  AOI22_X1 U6887 ( .A1(n5797), .A2(n6500), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n5796), .ZN(n5775) );
  OAI21_X1 U6888 ( .B1(n5799), .B2(n6505), .A(n5775), .ZN(n5776) );
  AOI21_X1 U6889 ( .B1(n6501), .B2(n5801), .A(n5776), .ZN(n5777) );
  OAI21_X1 U6890 ( .B1(n5803), .B2(n6419), .A(n5777), .ZN(U3028) );
  AOI22_X1 U6891 ( .A1(n5797), .A2(n6506), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n5796), .ZN(n5778) );
  OAI21_X1 U6892 ( .B1(n5799), .B2(n6511), .A(n5778), .ZN(n5779) );
  AOI21_X1 U6893 ( .B1(n6507), .B2(n5801), .A(n5779), .ZN(n5780) );
  OAI21_X1 U6894 ( .B1(n5803), .B2(n6422), .A(n5780), .ZN(U3029) );
  AOI22_X1 U6895 ( .A1(n5797), .A2(n6423), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n5796), .ZN(n5781) );
  OAI21_X1 U6896 ( .B1(n5799), .B2(n6388), .A(n5781), .ZN(n5782) );
  AOI21_X1 U6897 ( .B1(n6467), .B2(n5801), .A(n5782), .ZN(n5783) );
  OAI21_X1 U6898 ( .B1(n5803), .B2(n6426), .A(n5783), .ZN(U3030) );
  AOI22_X1 U6899 ( .A1(n5797), .A2(n6512), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n5796), .ZN(n5784) );
  OAI21_X1 U6900 ( .B1(n5799), .B2(n6517), .A(n5784), .ZN(n5785) );
  AOI21_X1 U6901 ( .B1(n6513), .B2(n5801), .A(n5785), .ZN(n5786) );
  OAI21_X1 U6902 ( .B1(n5803), .B2(n6429), .A(n5786), .ZN(U3031) );
  AOI22_X1 U6903 ( .A1(n5797), .A2(n6518), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n5796), .ZN(n5787) );
  OAI21_X1 U6904 ( .B1(n5799), .B2(n6523), .A(n5787), .ZN(n5788) );
  AOI21_X1 U6905 ( .B1(n6519), .B2(n5801), .A(n5788), .ZN(n5789) );
  OAI21_X1 U6906 ( .B1(n5803), .B2(n6432), .A(n5789), .ZN(U3032) );
  AOI22_X1 U6907 ( .A1(n5797), .A2(n6433), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n5796), .ZN(n5790) );
  OAI21_X1 U6908 ( .B1(n5799), .B2(n6395), .A(n5790), .ZN(n5791) );
  AOI21_X1 U6909 ( .B1(n6481), .B2(n5801), .A(n5791), .ZN(n5792) );
  OAI21_X1 U6910 ( .B1(n5803), .B2(n6436), .A(n5792), .ZN(U3033) );
  AOI22_X1 U6911 ( .A1(n5797), .A2(n6524), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n5796), .ZN(n5793) );
  OAI21_X1 U6912 ( .B1(n5799), .B2(n6529), .A(n5793), .ZN(n5794) );
  AOI21_X1 U6913 ( .B1(n6525), .B2(n5801), .A(n5794), .ZN(n5795) );
  OAI21_X1 U6914 ( .B1(n5803), .B2(n6439), .A(n5795), .ZN(U3034) );
  AOI22_X1 U6915 ( .A1(n5797), .A2(n6531), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n5796), .ZN(n5798) );
  OAI21_X1 U6916 ( .B1(n5799), .B2(n6540), .A(n5798), .ZN(n5800) );
  AOI21_X1 U6917 ( .B1(n6533), .B2(n5801), .A(n5800), .ZN(n5802) );
  OAI21_X1 U6918 ( .B1(n5803), .B2(n6445), .A(n5802), .ZN(U3035) );
  AND2_X1 U6919 ( .A1(n6164), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6920 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5805), .A(n5804), .ZN(
        n5806) );
  NAND2_X1 U6921 ( .A1(n5988), .A2(n5806), .ZN(U2788) );
  AOI22_X1 U6922 ( .A1(EBX_REG_29__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6083), .ZN(n5807) );
  OAI21_X1 U6923 ( .B1(n5808), .B2(n6108), .A(n5807), .ZN(n5809) );
  AOI21_X1 U6924 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5816), .A(n5809), .ZN(n5814) );
  INV_X1 U6925 ( .A(n5812), .ZN(n5813) );
  OAI211_X1 U6926 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5815), .A(n5814), .B(n5813), .ZN(U2798) );
  AOI22_X1 U6927 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6083), .ZN(n5824) );
  AOI22_X1 U6928 ( .A1(n5817), .A2(n6096), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5816), .ZN(n5823) );
  NOR2_X1 U6929 ( .A1(n5818), .A2(n6104), .ZN(n5819) );
  AOI21_X1 U6930 ( .B1(n5820), .B2(n6064), .A(n5819), .ZN(n5822) );
  NAND3_X1 U6931 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5830), .A3(n6807), .ZN(
        n5821) );
  NAND4_X1 U6932 ( .A1(n5824), .A2(n5823), .A3(n5822), .A4(n5821), .ZN(U2799)
         );
  NOR2_X1 U6933 ( .A1(n5901), .A2(n5825), .ZN(n5839) );
  AOI22_X1 U6934 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6083), .ZN(n5826) );
  OAI21_X1 U6935 ( .B1(n5827), .B2(n6108), .A(n5826), .ZN(n5828) );
  AOI221_X1 U6936 ( .B1(n5839), .B2(REIP_REG_27__SCAN_IN), .C1(n5830), .C2(
        n5829), .A(n5828), .ZN(n5833) );
  NOR2_X1 U6937 ( .A1(n5906), .A2(n6104), .ZN(n5831) );
  AOI21_X1 U6938 ( .B1(n5917), .B2(n6064), .A(n5831), .ZN(n5832) );
  NAND2_X1 U6939 ( .A1(n5833), .A2(n5832), .ZN(U2800) );
  AOI22_X1 U6940 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6083), .B1(n5834), 
        .B2(n6096), .ZN(n5841) );
  NAND2_X1 U6941 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5845) );
  INV_X1 U6942 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6805) );
  OAI21_X1 U6943 ( .B1(n5854), .B2(n5845), .A(n6805), .ZN(n5838) );
  OAI22_X1 U6944 ( .A1(n5836), .A2(n6044), .B1(n5835), .B2(n6104), .ZN(n5837)
         );
  AOI21_X1 U6945 ( .B1(n5839), .B2(n5838), .A(n5837), .ZN(n5840) );
  OAI211_X1 U6946 ( .C1(n5842), .C2(n6049), .A(n5841), .B(n5840), .ZN(U2801)
         );
  AOI22_X1 U6947 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6083), .ZN(n5850) );
  INV_X1 U6948 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U6949 ( .A1(n6105), .A2(n5843), .ZN(n5862) );
  OAI22_X1 U6950 ( .A1(n5940), .A2(n6108), .B1(n6643), .B2(n5862), .ZN(n5844)
         );
  INV_X1 U6951 ( .A(n5844), .ZN(n5849) );
  AOI22_X1 U6952 ( .A1(n5937), .A2(n6064), .B1(n6107), .B2(n5957), .ZN(n5848)
         );
  INV_X1 U6953 ( .A(n5854), .ZN(n5846) );
  OAI211_X1 U6954 ( .C1(REIP_REG_24__SCAN_IN), .C2(REIP_REG_25__SCAN_IN), .A(
        n5846), .B(n5845), .ZN(n5847) );
  NAND4_X1 U6955 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(U2802)
         );
  INV_X1 U6956 ( .A(n5862), .ZN(n5851) );
  AOI22_X1 U6957 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5851), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n6083), .ZN(n5852) );
  OAI21_X1 U6958 ( .B1(n5853), .B2(n6108), .A(n5852), .ZN(n5857) );
  OAI22_X1 U6959 ( .A1(n5855), .A2(n6044), .B1(REIP_REG_24__SCAN_IN), .B2(
        n5854), .ZN(n5856) );
  AOI211_X1 U6960 ( .C1(EBX_REG_24__SCAN_IN), .C2(n6110), .A(n5857), .B(n5856), 
        .ZN(n5858) );
  OAI21_X1 U6961 ( .B1(n5859), .B2(n6104), .A(n5858), .ZN(U2803) );
  AOI22_X1 U6962 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6083), .ZN(n5866) );
  NAND2_X1 U6963 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5873) );
  INV_X1 U6964 ( .A(n5873), .ZN(n5860) );
  AOI21_X1 U6965 ( .B1(n5881), .B2(n5860), .A(REIP_REG_23__SCAN_IN), .ZN(n5863) );
  OAI22_X1 U6966 ( .A1(n5863), .A2(n5862), .B1(n5861), .B2(n6104), .ZN(n5864)
         );
  AOI21_X1 U6967 ( .B1(n5922), .B2(n6064), .A(n5864), .ZN(n5865) );
  OAI211_X1 U6968 ( .C1(n5867), .C2(n6108), .A(n5866), .B(n5865), .ZN(U2804)
         );
  AOI22_X1 U6969 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6083), .ZN(n5877) );
  NOR2_X1 U6970 ( .A1(n5901), .A2(n5868), .ZN(n5887) );
  AOI22_X1 U6971 ( .A1(n5869), .A2(n6096), .B1(REIP_REG_22__SCAN_IN), .B2(
        n5887), .ZN(n5876) );
  OAI22_X1 U6972 ( .A1(n5871), .A2(n6044), .B1(n5870), .B2(n6104), .ZN(n5872)
         );
  INV_X1 U6973 ( .A(n5872), .ZN(n5875) );
  OAI211_X1 U6974 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5881), .B(n5873), .ZN(n5874) );
  NAND4_X1 U6975 ( .A1(n5877), .A2(n5876), .A3(n5875), .A4(n5874), .ZN(U2805)
         );
  AOI22_X1 U6976 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6083), .ZN(n5878) );
  OAI21_X1 U6977 ( .B1(n5879), .B2(n6108), .A(n5878), .ZN(n5880) );
  AOI221_X1 U6978 ( .B1(n5887), .B2(REIP_REG_21__SCAN_IN), .C1(n5881), .C2(
        n5543), .A(n5880), .ZN(n5883) );
  NAND2_X1 U6979 ( .A1(n5928), .A2(n6064), .ZN(n5882) );
  OAI211_X1 U6980 ( .C1(n6104), .C2(n5884), .A(n5883), .B(n5882), .ZN(U2806)
         );
  AOI22_X1 U6981 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6083), .ZN(n5893) );
  INV_X1 U6982 ( .A(n5885), .ZN(n5910) );
  AOI22_X1 U6983 ( .A1(n5931), .A2(n6064), .B1(n5910), .B2(n6107), .ZN(n5892)
         );
  INV_X1 U6984 ( .A(n5886), .ZN(n5888) );
  OAI21_X1 U6985 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5888), .A(n5887), .ZN(n5891) );
  NAND2_X1 U6986 ( .A1(n5889), .A2(n6096), .ZN(n5890) );
  NAND4_X1 U6987 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(U2807)
         );
  INV_X1 U6988 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6636) );
  INV_X1 U6989 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5948) );
  OAI21_X1 U6990 ( .B1(n6109), .B2(n5948), .A(n6067), .ZN(n5895) );
  OAI22_X1 U6991 ( .A1(n5915), .A2(n6049), .B1(n5942), .B2(n6108), .ZN(n5894)
         );
  AOI211_X1 U6992 ( .C1(n5896), .C2(n6636), .A(n5895), .B(n5894), .ZN(n5905)
         );
  AND2_X1 U6993 ( .A1(n5560), .A2(n5897), .ZN(n5898) );
  NOR2_X1 U6994 ( .A1(n3110), .A2(n5898), .ZN(n5943) );
  NOR2_X1 U6995 ( .A1(n5912), .A2(n6104), .ZN(n5899) );
  AOI21_X1 U6996 ( .B1(n5943), .B2(n6064), .A(n5899), .ZN(n5904) );
  NOR2_X1 U6997 ( .A1(n5901), .A2(n5900), .ZN(n6014) );
  NOR2_X1 U6998 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5902), .ZN(n6011) );
  OAI21_X1 U6999 ( .B1(n6014), .B2(n6011), .A(REIP_REG_19__SCAN_IN), .ZN(n5903) );
  NAND3_X1 U7000 ( .A1(n5905), .A2(n5904), .A3(n5903), .ZN(U2808) );
  NOR2_X1 U7001 ( .A1(n5906), .A2(n7014), .ZN(n5907) );
  AOI21_X1 U7002 ( .B1(n5917), .B2(n6125), .A(n5907), .ZN(n5908) );
  OAI21_X1 U7003 ( .B1(n7016), .B2(n5909), .A(n5908), .ZN(U2832) );
  AOI22_X1 U7004 ( .A1(n5931), .A2(n6125), .B1(n5910), .B2(n6124), .ZN(n5911)
         );
  OAI21_X1 U7005 ( .B1(n7016), .B2(n4302), .A(n5911), .ZN(U2839) );
  NOR2_X1 U7006 ( .A1(n5912), .A2(n7014), .ZN(n5913) );
  AOI21_X1 U7007 ( .B1(n5943), .B2(n6125), .A(n5913), .ZN(n5914) );
  OAI21_X1 U7008 ( .B1(n7016), .B2(n5915), .A(n5914), .ZN(U2840) );
  AOI22_X1 U7009 ( .A1(n5917), .A2(n6131), .B1(n6130), .B2(DATAI_27_), .ZN(
        n5919) );
  AOI22_X1 U7010 ( .A1(n6134), .A2(DATAI_11_), .B1(n6133), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5918) );
  NAND2_X1 U7011 ( .A1(n5919), .A2(n5918), .ZN(U2864) );
  AOI22_X1 U7012 ( .A1(n5937), .A2(n6131), .B1(n6130), .B2(DATAI_25_), .ZN(
        n5921) );
  AOI22_X1 U7013 ( .A1(n6134), .A2(DATAI_9_), .B1(n6133), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5920) );
  NAND2_X1 U7014 ( .A1(n5921), .A2(n5920), .ZN(U2866) );
  AOI22_X1 U7015 ( .A1(n5922), .A2(n6131), .B1(n6130), .B2(DATAI_23_), .ZN(
        n5924) );
  AOI22_X1 U7016 ( .A1(n6134), .A2(DATAI_7_), .B1(n6133), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7017 ( .A1(n5924), .A2(n5923), .ZN(U2868) );
  AOI22_X1 U7018 ( .A1(n5925), .A2(n6131), .B1(n6130), .B2(DATAI_22_), .ZN(
        n5927) );
  AOI22_X1 U7019 ( .A1(n6134), .A2(DATAI_6_), .B1(n6133), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7020 ( .A1(n5927), .A2(n5926), .ZN(U2869) );
  AOI22_X1 U7021 ( .A1(n5928), .A2(n6131), .B1(n6130), .B2(DATAI_21_), .ZN(
        n5930) );
  AOI22_X1 U7022 ( .A1(n6134), .A2(DATAI_5_), .B1(n6133), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5929) );
  NAND2_X1 U7023 ( .A1(n5930), .A2(n5929), .ZN(U2870) );
  AOI22_X1 U7024 ( .A1(n5931), .A2(n6131), .B1(n6130), .B2(DATAI_20_), .ZN(
        n5933) );
  AOI22_X1 U7025 ( .A1(n6134), .A2(DATAI_4_), .B1(n6133), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5932) );
  NAND2_X1 U7026 ( .A1(n5933), .A2(n5932), .ZN(U2871) );
  AOI22_X1 U7027 ( .A1(n5943), .A2(n6131), .B1(n6130), .B2(DATAI_19_), .ZN(
        n5935) );
  AOI22_X1 U7028 ( .A1(n6134), .A2(DATAI_3_), .B1(n6133), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7029 ( .A1(n5935), .A2(n5934), .ZN(U2872) );
  AOI22_X1 U7030 ( .A1(n6283), .A2(REIP_REG_25__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5939) );
  INV_X1 U7031 ( .A(n5503), .ZN(n5936) );
  OAI21_X1 U7032 ( .B1(n5936), .B2(n3125), .A(n3621), .ZN(n5958) );
  AOI22_X1 U7033 ( .A1(n5937), .A2(n6223), .B1(n6224), .B2(n5958), .ZN(n5938)
         );
  OAI211_X1 U7034 ( .C1(n6228), .C2(n5940), .A(n5939), .B(n5938), .ZN(U2961)
         );
  INV_X1 U7035 ( .A(n5941), .ZN(n5945) );
  INV_X1 U7036 ( .A(n5942), .ZN(n5944) );
  AOI222_X1 U7037 ( .A1(n5945), .A2(n6224), .B1(n5944), .B2(n6196), .C1(n6223), 
        .C2(n5943), .ZN(n5947) );
  OAI211_X1 U7038 ( .C1(n5948), .C2(n5955), .A(n5947), .B(n5946), .ZN(U2967)
         );
  INV_X1 U7039 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6016) );
  OR2_X1 U7040 ( .A1(n5367), .A2(n5949), .ZN(n5950) );
  AND2_X1 U7041 ( .A1(n5950), .A2(n5561), .ZN(n6132) );
  INV_X1 U7042 ( .A(n6015), .ZN(n5951) );
  AOI222_X1 U7043 ( .A1(n5952), .A2(n6224), .B1(n6223), .B2(n6132), .C1(n5951), 
        .C2(n6196), .ZN(n5954) );
  OAI211_X1 U7044 ( .C1(n6016), .C2(n5955), .A(n5954), .B(n5953), .ZN(U2969)
         );
  AOI22_X1 U7045 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6283), .B1(n5956), .B2(
        n6788), .ZN(n5960) );
  AOI22_X1 U7046 ( .A1(n5958), .A2(n6315), .B1(n5611), .B2(n5957), .ZN(n5959)
         );
  OAI211_X1 U7047 ( .C1(n5961), .C2(n6788), .A(n5960), .B(n5959), .ZN(U2993)
         );
  AOI22_X1 U7048 ( .A1(n5963), .A2(n6315), .B1(n5611), .B2(n5962), .ZN(n5971)
         );
  NAND2_X1 U7049 ( .A1(n6283), .A2(REIP_REG_16__SCAN_IN), .ZN(n5970) );
  OAI21_X1 U7050 ( .B1(n5965), .B2(n5964), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5969) );
  NAND3_X1 U7051 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5967), .A3(n5966), .ZN(n5968) );
  NAND4_X1 U7052 ( .A1(n5971), .A2(n5970), .A3(n5969), .A4(n5968), .ZN(U3002)
         );
  INV_X1 U7053 ( .A(n5972), .ZN(n5980) );
  INV_X1 U7054 ( .A(n5973), .ZN(n5974) );
  AOI21_X1 U7055 ( .B1(n5975), .B2(n5611), .A(n5974), .ZN(n5979) );
  AOI22_X1 U7056 ( .A1(n5977), .A2(n6315), .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5976), .ZN(n5978) );
  OAI211_X1 U7057 ( .C1(n6236), .C2(n5980), .A(n5979), .B(n5978), .ZN(U3005)
         );
  NAND4_X1 U7058 ( .A1(n5983), .A2(n5982), .A3(n5981), .A4(n6070), .ZN(n5984)
         );
  OAI21_X1 U7059 ( .B1(n6668), .B2(n6802), .A(n5984), .ZN(U3455) );
  INV_X1 U7060 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6794) );
  INV_X2 U7061 ( .A(n6706), .ZN(n6656) );
  OAI221_X1 U7062 ( .B1(n6593), .B2(n6777), .C1(STATE_REG_1__SCAN_IN), .C2(
        n6777), .A(n6656), .ZN(n5985) );
  OAI21_X1 U7063 ( .B1(n6706), .B2(n6794), .A(n6592), .ZN(U2789) );
  OAI21_X1 U7064 ( .B1(n5986), .B2(n6581), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5987) );
  OAI21_X1 U7065 ( .B1(n5988), .B2(n6576), .A(n5987), .ZN(U2790) );
  NOR2_X1 U7066 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5990) );
  OAI21_X1 U7067 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5990), .A(n6656), .ZN(n5989)
         );
  OAI21_X1 U7068 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6656), .A(n5989), .ZN(
        U2791) );
  OAI21_X1 U7069 ( .B1(n5990), .B2(BS16_N), .A(n6659), .ZN(n6658) );
  OAI21_X1 U7070 ( .B1(n6659), .B2(n5991), .A(n6658), .ZN(U2792) );
  OAI21_X1 U7071 ( .B1(n5993), .B2(n5992), .A(n6213), .ZN(U2793) );
  NOR4_X1 U7072 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5997) );
  NOR4_X1 U7073 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5996) );
  NOR4_X1 U7074 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n5995) );
  NOR4_X1 U7075 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5994) );
  NAND4_X1 U7076 ( .A1(n5997), .A2(n5996), .A3(n5995), .A4(n5994), .ZN(n6003)
         );
  NOR4_X1 U7077 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6001) );
  AOI211_X1 U7078 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_12__SCAN_IN), .B(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6000) );
  NOR4_X1 U7079 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n5999)
         );
  NOR4_X1 U7080 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5998) );
  NAND4_X1 U7081 ( .A1(n6001), .A2(n6000), .A3(n5999), .A4(n5998), .ZN(n6002)
         );
  NOR2_X1 U7082 ( .A1(n6003), .A2(n6002), .ZN(n6686) );
  INV_X1 U7083 ( .A(n6686), .ZN(n6690) );
  NAND2_X1 U7084 ( .A1(n6686), .A2(n4473), .ZN(n6685) );
  NOR3_X1 U7085 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6685), .ZN(n6005) );
  AOI21_X1 U7086 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6690), .A(n6005), .ZN(
        n6004) );
  OAI21_X1 U7087 ( .B1(n5117), .B2(n6690), .A(n6004), .ZN(U2794) );
  NOR2_X1 U7088 ( .A1(n6690), .A2(REIP_REG_1__SCAN_IN), .ZN(n6691) );
  INV_X1 U7089 ( .A(n6691), .ZN(n6683) );
  AOI21_X1 U7090 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n6690), .A(n6005), .ZN(
        n6006) );
  OAI21_X1 U7091 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6683), .A(n6006), .ZN(
        U2795) );
  INV_X1 U7092 ( .A(n7017), .ZN(n6127) );
  AOI22_X1 U7093 ( .A1(n6007), .A2(n6096), .B1(REIP_REG_18__SCAN_IN), .B2(
        n6014), .ZN(n6009) );
  AOI21_X1 U7094 ( .B1(n6083), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n6041), 
        .ZN(n6008) );
  OAI211_X1 U7095 ( .C1(n4298), .C2(n6049), .A(n6009), .B(n6008), .ZN(n6010)
         );
  AOI211_X1 U7096 ( .C1(n6127), .C2(n6064), .A(n6011), .B(n6010), .ZN(n6012)
         );
  OAI21_X1 U7097 ( .B1(n6104), .B2(n7015), .A(n6012), .ZN(U2809) );
  AOI21_X1 U7098 ( .B1(REIP_REG_16__SCAN_IN), .B2(n6013), .A(
        REIP_REG_17__SCAN_IN), .ZN(n6021) );
  INV_X1 U7099 ( .A(n6014), .ZN(n6020) );
  OAI22_X1 U7100 ( .A1(n6016), .A2(n6109), .B1(n6015), .B2(n6108), .ZN(n6017)
         );
  AOI211_X1 U7101 ( .C1(n6110), .C2(EBX_REG_17__SCAN_IN), .A(n6041), .B(n6017), 
        .ZN(n6019) );
  AOI22_X1 U7102 ( .A1(n6132), .A2(n6064), .B1(n6117), .B2(n6107), .ZN(n6018)
         );
  OAI211_X1 U7103 ( .C1(n6021), .C2(n6020), .A(n6019), .B(n6018), .ZN(U2810)
         );
  AOI22_X1 U7104 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6083), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6022), .ZN(n6023) );
  OAI211_X1 U7105 ( .C1(n6049), .C2(n6122), .A(n6023), .B(n6067), .ZN(n6024)
         );
  AOI211_X1 U7106 ( .C1(n6119), .C2(n6107), .A(n6025), .B(n6024), .ZN(n6028)
         );
  AOI22_X1 U7107 ( .A1(n6120), .A2(n6064), .B1(n6026), .B2(n6096), .ZN(n6027)
         );
  NAND2_X1 U7108 ( .A1(n6028), .A2(n6027), .ZN(U2812) );
  AOI22_X1 U7109 ( .A1(n6107), .A2(n6031), .B1(n6030), .B2(n6029), .ZN(n6037)
         );
  INV_X1 U7110 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6625) );
  OAI22_X1 U7111 ( .A1(n6033), .A2(n6625), .B1(n6032), .B2(n6109), .ZN(n6034)
         );
  AOI211_X1 U7112 ( .C1(n6110), .C2(EBX_REG_11__SCAN_IN), .A(n6041), .B(n6034), 
        .ZN(n6036) );
  AOI22_X1 U7113 ( .A1(n6197), .A2(n6064), .B1(n6096), .B2(n6195), .ZN(n6035)
         );
  NAND3_X1 U7114 ( .A1(n6037), .A2(n6036), .A3(n6035), .ZN(U2816) );
  INV_X1 U7115 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6902) );
  NAND2_X1 U7116 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6902), .ZN(n6726) );
  NAND2_X1 U7117 ( .A1(n6039), .A2(n6038), .ZN(n6042) );
  OAI22_X1 U7118 ( .A1(n6104), .A2(n6244), .B1(n6726), .B2(n6042), .ZN(n6040)
         );
  AOI211_X1 U7119 ( .C1(n6083), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6041), 
        .B(n6040), .ZN(n6048) );
  NOR2_X1 U7120 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6042), .ZN(n6052) );
  OAI22_X1 U7121 ( .A1(n6045), .A2(n6044), .B1(n6043), .B2(n6108), .ZN(n6046)
         );
  AOI221_X1 U7122 ( .B1(n6052), .B2(REIP_REG_10__SCAN_IN), .C1(n6055), .C2(
        REIP_REG_10__SCAN_IN), .A(n6046), .ZN(n6047) );
  OAI211_X1 U7123 ( .C1(n4264), .C2(n6049), .A(n6048), .B(n6047), .ZN(U2817)
         );
  AOI22_X1 U7124 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6110), .B1(n6107), .B2(n6249), 
        .ZN(n6050) );
  OAI211_X1 U7125 ( .C1(n6109), .C2(n6051), .A(n6050), .B(n6067), .ZN(n6053)
         );
  AOI211_X1 U7126 ( .C1(n6054), .C2(n6064), .A(n6053), .B(n6052), .ZN(n6058)
         );
  AOI22_X1 U7127 ( .A1(n6056), .A2(n6096), .B1(REIP_REG_9__SCAN_IN), .B2(n6055), .ZN(n6057) );
  NAND2_X1 U7128 ( .A1(n6058), .A2(n6057), .ZN(U2818) );
  AOI22_X1 U7129 ( .A1(EBX_REG_6__SCAN_IN), .A2(n6110), .B1(
        PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6083), .ZN(n6059) );
  OAI211_X1 U7130 ( .C1(n6104), .C2(n6060), .A(n6059), .B(n6067), .ZN(n6061)
         );
  AOI211_X1 U7131 ( .C1(REIP_REG_6__SCAN_IN), .C2(n6063), .A(n6062), .B(n6061), 
        .ZN(n6066) );
  NAND2_X1 U7132 ( .A1(n6202), .A2(n6064), .ZN(n6065) );
  OAI211_X1 U7133 ( .C1(n6108), .C2(n6206), .A(n6066), .B(n6065), .ZN(U2821)
         );
  INV_X1 U7134 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6958) );
  OAI21_X1 U7135 ( .B1(n6109), .B2(n6958), .A(n6067), .ZN(n6069) );
  OAI21_X1 U7136 ( .B1(n6095), .B2(n6072), .A(n6105), .ZN(n6091) );
  NOR2_X1 U7137 ( .A1(n6091), .A2(n6615), .ZN(n6068) );
  AOI211_X1 U7138 ( .C1(n6111), .C2(n6070), .A(n6069), .B(n6068), .ZN(n6079)
         );
  NOR2_X1 U7139 ( .A1(n6116), .A2(n6212), .ZN(n6077) );
  NAND2_X1 U7140 ( .A1(n6107), .A2(n6071), .ZN(n6075) );
  NAND2_X1 U7141 ( .A1(n6110), .A2(EBX_REG_4__SCAN_IN), .ZN(n6074) );
  OR3_X1 U7142 ( .A1(n6092), .A2(REIP_REG_4__SCAN_IN), .A3(n6072), .ZN(n6073)
         );
  NAND3_X1 U7143 ( .A1(n6075), .A2(n6074), .A3(n6073), .ZN(n6076) );
  NOR2_X1 U7144 ( .A1(n6077), .A2(n6076), .ZN(n6078) );
  OAI211_X1 U7145 ( .C1(n6217), .C2(n6108), .A(n6079), .B(n6078), .ZN(U2823)
         );
  INV_X1 U7146 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6753) );
  INV_X1 U7147 ( .A(n6080), .ZN(n6081) );
  NAND2_X1 U7148 ( .A1(n6081), .A2(REIP_REG_2__SCAN_IN), .ZN(n6090) );
  INV_X1 U7149 ( .A(n6082), .ZN(n6305) );
  AOI22_X1 U7150 ( .A1(n6107), .A2(n6305), .B1(n6110), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n6085) );
  AOI22_X1 U7151 ( .A1(n6111), .A2(n6677), .B1(n6083), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6084) );
  OAI211_X1 U7152 ( .C1(n6116), .C2(n6086), .A(n6085), .B(n6084), .ZN(n6087)
         );
  AOI21_X1 U7153 ( .B1(n6088), .B2(n6096), .A(n6087), .ZN(n6089) );
  OAI221_X1 U7154 ( .B1(n6091), .B2(n6753), .C1(n6091), .C2(n6090), .A(n6089), 
        .ZN(U2824) );
  INV_X1 U7155 ( .A(n6092), .ZN(n6093) );
  AOI22_X1 U7156 ( .A1(n6093), .A2(n5117), .B1(n6110), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n6103) );
  NOR2_X1 U7157 ( .A1(n6116), .A2(n6094), .ZN(n6101) );
  NAND2_X1 U7158 ( .A1(n6111), .A2(n4519), .ZN(n6098) );
  AOI22_X1 U7159 ( .A1(n6096), .A2(n6099), .B1(REIP_REG_1__SCAN_IN), .B2(n6095), .ZN(n6097) );
  OAI211_X1 U7160 ( .C1(n6099), .C2(n6109), .A(n6098), .B(n6097), .ZN(n6100)
         );
  NOR2_X1 U7161 ( .A1(n6101), .A2(n6100), .ZN(n6102) );
  OAI211_X1 U7162 ( .C1(n4465), .C2(n6104), .A(n6103), .B(n6102), .ZN(U2826)
         );
  AOI22_X1 U7163 ( .A1(n6107), .A2(n6106), .B1(REIP_REG_0__SCAN_IN), .B2(n6105), .ZN(n6114) );
  NAND2_X1 U7164 ( .A1(n6109), .A2(n6108), .ZN(n6112) );
  AOI222_X1 U7165 ( .A1(n6112), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n6111), 
        .B2(n3690), .C1(EBX_REG_0__SCAN_IN), .C2(n6110), .ZN(n6113) );
  OAI211_X1 U7166 ( .C1(n6116), .C2(n6115), .A(n6114), .B(n6113), .ZN(U2827)
         );
  AOI22_X1 U7167 ( .A1(n6132), .A2(n6125), .B1(n6117), .B2(n6124), .ZN(n6118)
         );
  OAI21_X1 U7168 ( .B1(n7016), .B2(n6918), .A(n6118), .ZN(U2842) );
  AOI22_X1 U7169 ( .A1(n6120), .A2(n6125), .B1(n6124), .B2(n6119), .ZN(n6121)
         );
  OAI21_X1 U7170 ( .B1(n7016), .B2(n6122), .A(n6121), .ZN(U2844) );
  INV_X1 U7171 ( .A(n6123), .ZN(n6222) );
  AOI22_X1 U7172 ( .A1(n6222), .A2(n6125), .B1(n6124), .B2(n6313), .ZN(n6126)
         );
  OAI21_X1 U7173 ( .B1(n7016), .B2(n4234), .A(n6126), .ZN(U2857) );
  AOI22_X1 U7174 ( .A1(n6127), .A2(n6131), .B1(n6130), .B2(DATAI_18_), .ZN(
        n6129) );
  AOI22_X1 U7175 ( .A1(n6134), .A2(DATAI_2_), .B1(n6133), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6128) );
  NAND2_X1 U7176 ( .A1(n6129), .A2(n6128), .ZN(U2873) );
  AOI22_X1 U7177 ( .A1(n6132), .A2(n6131), .B1(n6130), .B2(DATAI_17_), .ZN(
        n6136) );
  AOI22_X1 U7178 ( .A1(n6134), .A2(DATAI_1_), .B1(n6133), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7179 ( .A1(n6136), .A2(n6135), .ZN(U2874) );
  INV_X1 U7180 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n6904) );
  AOI22_X1 U7181 ( .A1(n6141), .A2(EAX_REG_26__SCAN_IN), .B1(n6567), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6137) );
  OAI21_X1 U7182 ( .B1(n6904), .B2(n6146), .A(n6137), .ZN(U2897) );
  INV_X1 U7183 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6982) );
  AOI22_X1 U7184 ( .A1(n6141), .A2(EAX_REG_25__SCAN_IN), .B1(n6567), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7185 ( .B1(n6982), .B2(n6146), .A(n6138), .ZN(U2898) );
  INV_X1 U7186 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6756) );
  AOI22_X1 U7187 ( .A1(n6141), .A2(EAX_REG_22__SCAN_IN), .B1(n6567), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6139) );
  OAI21_X1 U7188 ( .B1(n6756), .B2(n6146), .A(n6139), .ZN(U2901) );
  AOI22_X1 U7189 ( .A1(n6164), .A2(DATAO_REG_18__SCAN_IN), .B1(n6141), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7190 ( .B1(n4555), .B2(n6696), .A(n6140), .ZN(U2905) );
  INV_X1 U7191 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U7192 ( .A1(n6141), .A2(EAX_REG_17__SCAN_IN), .B1(n6567), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n6142) );
  OAI21_X1 U7193 ( .B1(n6772), .B2(n6146), .A(n6142), .ZN(U2906) );
  INV_X1 U7194 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6194) );
  AOI22_X1 U7195 ( .A1(n6567), .A2(LWORD_REG_15__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6143) );
  OAI21_X1 U7196 ( .B1(n6194), .B2(n6166), .A(n6143), .ZN(U2908) );
  INV_X1 U7197 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6968) );
  AOI22_X1 U7198 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6161), .B1(n6164), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6144) );
  OAI21_X1 U7199 ( .B1(n6968), .B2(n6696), .A(n6144), .ZN(U2909) );
  INV_X1 U7200 ( .A(DATAO_REG_13__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U7201 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6161), .B1(n6157), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6145) );
  OAI21_X1 U7202 ( .B1(n6803), .B2(n6146), .A(n6145), .ZN(U2910) );
  INV_X1 U7203 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6148) );
  AOI22_X1 U7204 ( .A1(n6567), .A2(LWORD_REG_12__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6147) );
  OAI21_X1 U7205 ( .B1(n6148), .B2(n6166), .A(n6147), .ZN(U2911) );
  AOI222_X1 U7206 ( .A1(n6157), .A2(LWORD_REG_11__SCAN_IN), .B1(n6161), .B2(
        EAX_REG_11__SCAN_IN), .C1(DATAO_REG_11__SCAN_IN), .C2(n6164), .ZN(
        n6149) );
  INV_X1 U7207 ( .A(n6149), .ZN(U2912) );
  AOI222_X1 U7208 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6157), .B1(n6161), .B2(
        EAX_REG_10__SCAN_IN), .C1(DATAO_REG_10__SCAN_IN), .C2(n6164), .ZN(
        n6150) );
  INV_X1 U7209 ( .A(n6150), .ZN(U2913) );
  INV_X1 U7210 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6152) );
  AOI22_X1 U7211 ( .A1(n6567), .A2(LWORD_REG_9__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6151) );
  OAI21_X1 U7212 ( .B1(n6152), .B2(n6166), .A(n6151), .ZN(U2914) );
  AOI222_X1 U7213 ( .A1(n6164), .A2(DATAO_REG_8__SCAN_IN), .B1(n6161), .B2(
        EAX_REG_8__SCAN_IN), .C1(LWORD_REG_8__SCAN_IN), .C2(n6567), .ZN(n6153)
         );
  INV_X1 U7214 ( .A(n6153), .ZN(U2915) );
  AOI22_X1 U7215 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6567), .B1(n6164), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7216 ( .B1(n6155), .B2(n6166), .A(n6154), .ZN(U2916) );
  INV_X1 U7217 ( .A(LWORD_REG_6__SCAN_IN), .ZN(n6837) );
  AOI22_X1 U7218 ( .A1(EAX_REG_6__SCAN_IN), .A2(n6161), .B1(n6164), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6156) );
  OAI21_X1 U7219 ( .B1(n6837), .B2(n6696), .A(n6156), .ZN(U2917) );
  AOI222_X1 U7220 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6157), .B1(n6161), .B2(
        EAX_REG_5__SCAN_IN), .C1(DATAO_REG_5__SCAN_IN), .C2(n6164), .ZN(n6158)
         );
  INV_X1 U7221 ( .A(n6158), .ZN(U2918) );
  AOI22_X1 U7222 ( .A1(n6567), .A2(LWORD_REG_4__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6159) );
  OAI21_X1 U7223 ( .B1(n4514), .B2(n6166), .A(n6159), .ZN(U2919) );
  AOI222_X1 U7224 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6567), .B1(n6161), .B2(
        EAX_REG_3__SCAN_IN), .C1(DATAO_REG_3__SCAN_IN), .C2(n6164), .ZN(n6160)
         );
  INV_X1 U7225 ( .A(n6160), .ZN(U2920) );
  AOI222_X1 U7226 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6567), .B1(n6161), .B2(
        EAX_REG_2__SCAN_IN), .C1(DATAO_REG_2__SCAN_IN), .C2(n6164), .ZN(n6162)
         );
  INV_X1 U7227 ( .A(n6162), .ZN(U2921) );
  AOI22_X1 U7228 ( .A1(n6567), .A2(LWORD_REG_1__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6163) );
  OAI21_X1 U7229 ( .B1(n4502), .B2(n6166), .A(n6163), .ZN(U2922) );
  AOI22_X1 U7230 ( .A1(n6567), .A2(LWORD_REG_0__SCAN_IN), .B1(n6164), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6165) );
  OAI21_X1 U7231 ( .B1(n4507), .B2(n6166), .A(n6165), .ZN(U2923) );
  AOI22_X1 U7232 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7233 ( .A1(n6190), .A2(DATAI_8_), .ZN(n6176) );
  NAND2_X1 U7234 ( .A1(n6167), .A2(n6176), .ZN(U2932) );
  AOI22_X1 U7235 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6168) );
  NAND2_X1 U7236 ( .A1(n6190), .A2(DATAI_9_), .ZN(n6178) );
  NAND2_X1 U7237 ( .A1(n6168), .A2(n6178), .ZN(U2933) );
  INV_X1 U7238 ( .A(DATAI_11_), .ZN(n6169) );
  NOR2_X1 U7239 ( .A1(n6174), .A2(n6169), .ZN(n6180) );
  AOI21_X1 U7240 ( .B1(n6191), .B2(UWORD_REG_11__SCAN_IN), .A(n6180), .ZN(
        n6170) );
  OAI21_X1 U7241 ( .B1(n6853), .B2(n6193), .A(n6170), .ZN(U2935) );
  AOI22_X1 U7242 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7243 ( .A1(n6190), .A2(DATAI_12_), .ZN(n6182) );
  NAND2_X1 U7244 ( .A1(n6171), .A2(n6182), .ZN(U2936) );
  AOI22_X1 U7245 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7246 ( .A1(n6190), .A2(DATAI_13_), .ZN(n6184) );
  NAND2_X1 U7247 ( .A1(n6172), .A2(n6184), .ZN(U2937) );
  INV_X1 U7248 ( .A(DATAI_14_), .ZN(n6173) );
  NOR2_X1 U7249 ( .A1(n6174), .A2(n6173), .ZN(n6186) );
  AOI21_X1 U7250 ( .B1(n6191), .B2(UWORD_REG_14__SCAN_IN), .A(n6186), .ZN(
        n6175) );
  OAI21_X1 U7251 ( .B1(n6844), .B2(n6193), .A(n6175), .ZN(U2938) );
  AOI22_X1 U7252 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6187), .B1(
        LWORD_REG_8__SCAN_IN), .B2(n6191), .ZN(n6177) );
  NAND2_X1 U7253 ( .A1(n6177), .A2(n6176), .ZN(U2947) );
  AOI22_X1 U7254 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7255 ( .A1(n6179), .A2(n6178), .ZN(U2948) );
  INV_X1 U7256 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6866) );
  AOI21_X1 U7257 ( .B1(n6187), .B2(EAX_REG_11__SCAN_IN), .A(n6180), .ZN(n6181)
         );
  OAI21_X1 U7258 ( .B1(n6866), .B2(n6189), .A(n6181), .ZN(U2950) );
  AOI22_X1 U7259 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7260 ( .A1(n6183), .A2(n6182), .ZN(U2951) );
  AOI22_X1 U7261 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6187), .B1(n6191), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6185) );
  NAND2_X1 U7262 ( .A1(n6185), .A2(n6184), .ZN(U2952) );
  AOI21_X1 U7263 ( .B1(n6187), .B2(EAX_REG_14__SCAN_IN), .A(n6186), .ZN(n6188)
         );
  OAI21_X1 U7264 ( .B1(n6968), .B2(n6189), .A(n6188), .ZN(U2953) );
  AOI22_X1 U7265 ( .A1(n6191), .A2(LWORD_REG_15__SCAN_IN), .B1(n6190), .B2(
        DATAI_15_), .ZN(n6192) );
  OAI21_X1 U7266 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(U2954) );
  AOI22_X1 U7267 ( .A1(n6283), .A2(REIP_REG_11__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6199) );
  AOI22_X1 U7268 ( .A1(n6197), .A2(n6223), .B1(n6196), .B2(n6195), .ZN(n6198)
         );
  OAI211_X1 U7269 ( .C1(n6200), .C2(n6213), .A(n6199), .B(n6198), .ZN(U2975)
         );
  AOI22_X1 U7270 ( .A1(n6283), .A2(REIP_REG_6__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6205) );
  INV_X1 U7271 ( .A(n6201), .ZN(n6203) );
  AOI22_X1 U7272 ( .A1(n6224), .A2(n6203), .B1(n6202), .B2(n6223), .ZN(n6204)
         );
  OAI211_X1 U7273 ( .C1(n6228), .C2(n6206), .A(n6205), .B(n6204), .ZN(U2980)
         );
  AOI22_X1 U7274 ( .A1(n6283), .A2(REIP_REG_4__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6216) );
  OR2_X1 U7275 ( .A1(n6208), .A2(n6207), .ZN(n6209) );
  NAND2_X1 U7276 ( .A1(n6210), .A2(n6209), .ZN(n6297) );
  OAI22_X1 U7277 ( .A1(n6213), .A2(n6297), .B1(n6212), .B2(n6211), .ZN(n6214)
         );
  INV_X1 U7278 ( .A(n6214), .ZN(n6215) );
  OAI211_X1 U7279 ( .C1(n6228), .C2(n6217), .A(n6216), .B(n6215), .ZN(U2982)
         );
  AOI22_X1 U7280 ( .A1(n6283), .A2(REIP_REG_2__SCAN_IN), .B1(n6218), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6226) );
  XOR2_X1 U7281 ( .A(n6219), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n6220) );
  XNOR2_X1 U7282 ( .A(n6221), .B(n6220), .ZN(n6314) );
  AOI22_X1 U7283 ( .A1(n6314), .A2(n6224), .B1(n6223), .B2(n6222), .ZN(n6225)
         );
  OAI211_X1 U7284 ( .C1(n6228), .C2(n6227), .A(n6226), .B(n6225), .ZN(U2984)
         );
  NAND2_X1 U7285 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6927), .ZN(n6709) );
  OAI22_X1 U7286 ( .A1(n6294), .A2(n6229), .B1(n6628), .B2(n6292), .ZN(n6230)
         );
  AOI21_X1 U7287 ( .B1(n6231), .B2(n6315), .A(n6230), .ZN(n6235) );
  OAI211_X1 U7288 ( .C1(n6241), .C2(n6233), .A(INSTADDRPOINTER_REG_12__SCAN_IN), .B(n6232), .ZN(n6234) );
  OAI211_X1 U7289 ( .C1(n6236), .C2(n6709), .A(n6235), .B(n6234), .ZN(U3006)
         );
  AOI22_X1 U7290 ( .A1(n6310), .A2(n6242), .B1(n6238), .B2(n6237), .ZN(n6240)
         );
  NAND2_X1 U7291 ( .A1(n6240), .A2(n6239), .ZN(n6264) );
  AOI21_X1 U7292 ( .B1(n6241), .B2(n6260), .A(n6264), .ZN(n6256) );
  NOR2_X1 U7293 ( .A1(n6289), .A2(n6242), .ZN(n6269) );
  NAND2_X1 U7294 ( .A1(n6243), .A2(n6269), .ZN(n6251) );
  AOI221_X1 U7295 ( .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n3600), .C2(n6255), .A(n6251), 
        .ZN(n6246) );
  OAI22_X1 U7296 ( .A1(n6294), .A2(n6244), .B1(n6902), .B2(n6292), .ZN(n6245)
         );
  AOI211_X1 U7297 ( .C1(n6247), .C2(n6315), .A(n6246), .B(n6245), .ZN(n6248)
         );
  OAI21_X1 U7298 ( .B1(n6256), .B2(n3600), .A(n6248), .ZN(U3008) );
  AOI22_X1 U7299 ( .A1(n5611), .A2(n6249), .B1(n6317), .B2(REIP_REG_9__SCAN_IN), .ZN(n6250) );
  OAI21_X1 U7300 ( .B1(n6251), .B2(INSTADDRPOINTER_REG_9__SCAN_IN), .A(n6250), 
        .ZN(n6252) );
  AOI21_X1 U7301 ( .B1(n6253), .B2(n6315), .A(n6252), .ZN(n6254) );
  OAI21_X1 U7302 ( .B1(n6256), .B2(n6255), .A(n6254), .ZN(U3009) );
  AOI21_X1 U7303 ( .B1(n5611), .B2(n6258), .A(n6257), .ZN(n6263) );
  AOI22_X1 U7304 ( .A1(n6259), .A2(n6315), .B1(INSTADDRPOINTER_REG_8__SCAN_IN), 
        .B2(n6264), .ZN(n6262) );
  OAI211_X1 U7305 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6269), .B(n6260), .ZN(n6261) );
  NAND3_X1 U7306 ( .A1(n6263), .A2(n6262), .A3(n6261), .ZN(U3010) );
  INV_X1 U7307 ( .A(n6264), .ZN(n6274) );
  INV_X1 U7308 ( .A(n6265), .ZN(n6266) );
  AOI21_X1 U7309 ( .B1(n5611), .B2(n6267), .A(n6266), .ZN(n6272) );
  INV_X1 U7310 ( .A(n6268), .ZN(n6270) );
  AOI22_X1 U7311 ( .A1(n6270), .A2(n6315), .B1(n6269), .B2(n6273), .ZN(n6271)
         );
  OAI211_X1 U7312 ( .C1(n6274), .C2(n6273), .A(n6272), .B(n6271), .ZN(U3011)
         );
  OAI21_X1 U7313 ( .B1(n6288), .B2(n6276), .A(n6275), .ZN(n6277) );
  AOI21_X1 U7314 ( .B1(n6278), .B2(n6318), .A(n6277), .ZN(n6286) );
  INV_X1 U7315 ( .A(n6279), .ZN(n6282) );
  INV_X1 U7316 ( .A(n6280), .ZN(n6281) );
  AOI22_X1 U7317 ( .A1(n6282), .A2(n6315), .B1(n5611), .B2(n6281), .ZN(n6285)
         );
  NAND2_X1 U7318 ( .A1(n6283), .A2(REIP_REG_5__SCAN_IN), .ZN(n6284) );
  OAI211_X1 U7319 ( .C1(n6287), .C2(n6286), .A(n6285), .B(n6284), .ZN(U3013)
         );
  NOR2_X1 U7320 ( .A1(n6288), .A2(n6291), .ZN(n6312) );
  NOR2_X1 U7321 ( .A1(n6312), .A2(n6316), .ZN(n6307) );
  INV_X1 U7322 ( .A(n6289), .ZN(n6290) );
  NAND2_X1 U7323 ( .A1(n6291), .A2(n6290), .ZN(n6308) );
  AOI211_X1 U7324 ( .C1(n6979), .C2(n6808), .A(n6747), .B(n6308), .ZN(n6299)
         );
  OAI22_X1 U7325 ( .A1(n6294), .A2(n6293), .B1(n6615), .B2(n6292), .ZN(n6295)
         );
  INV_X1 U7326 ( .A(n6295), .ZN(n6296) );
  OAI21_X1 U7327 ( .B1(n6297), .B2(n5745), .A(n6296), .ZN(n6298) );
  NOR2_X1 U7328 ( .A1(n6299), .A2(n6298), .ZN(n6300) );
  OAI21_X1 U7329 ( .B1(n6307), .B2(n6979), .A(n6300), .ZN(U3014) );
  INV_X1 U7330 ( .A(n6301), .ZN(n6304) );
  AND3_X1 U7331 ( .A1(n4658), .A2(n6315), .A3(n6302), .ZN(n6303) );
  AOI211_X1 U7332 ( .C1(n5611), .C2(n6305), .A(n6304), .B(n6303), .ZN(n6306)
         );
  OAI221_X1 U7333 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n6308), .C1(n6808), .C2(n6307), .A(n6306), .ZN(U3015) );
  AND3_X1 U7334 ( .A1(n6310), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(n6309), 
        .ZN(n6311) );
  AOI211_X1 U7335 ( .C1(n5611), .C2(n6313), .A(n6312), .B(n6311), .ZN(n6322)
         );
  AOI22_X1 U7336 ( .A1(n6316), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6315), 
        .B2(n6314), .ZN(n6321) );
  NAND2_X1 U7337 ( .A1(n6317), .A2(REIP_REG_2__SCAN_IN), .ZN(n6320) );
  NAND3_X1 U7338 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6318), .A3(n3476), 
        .ZN(n6319) );
  NAND4_X1 U7339 ( .A1(n6322), .A2(n6321), .A3(n6320), .A4(n6319), .ZN(U3016)
         );
  NOR2_X1 U7340 ( .A1(n6554), .A2(n6679), .ZN(U3019) );
  NAND2_X1 U7341 ( .A1(n6324), .A2(n6323), .ZN(n6673) );
  INV_X1 U7342 ( .A(n6410), .ZN(n6325) );
  NAND2_X1 U7343 ( .A1(n6326), .A2(n6325), .ZN(n6327) );
  OAI21_X1 U7344 ( .B1(n6673), .B2(n6327), .A(n6674), .ZN(n6337) );
  NOR2_X1 U7345 ( .A1(n6328), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6359)
         );
  INV_X1 U7346 ( .A(n6359), .ZN(n6329) );
  OAI21_X1 U7347 ( .B1(n6331), .B2(n6330), .A(n6329), .ZN(n6333) );
  OAI21_X1 U7348 ( .B1(n6337), .B2(n6333), .A(n6414), .ZN(n6332) );
  INV_X1 U7349 ( .A(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n6911) );
  AOI22_X1 U7350 ( .A1(n6501), .A2(n6359), .B1(n6500), .B2(n6358), .ZN(n6339)
         );
  INV_X1 U7351 ( .A(n6333), .ZN(n6336) );
  OAI22_X1 U7352 ( .A1(n6337), .A2(n6336), .B1(n6335), .B2(n6334), .ZN(n6360)
         );
  AOI22_X1 U7353 ( .A1(n6459), .A2(n6361), .B1(n6502), .B2(n6360), .ZN(n6338)
         );
  OAI211_X1 U7354 ( .C1(n6365), .C2(n6911), .A(n6339), .B(n6338), .ZN(U3044)
         );
  INV_X1 U7355 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6342) );
  AOI22_X1 U7356 ( .A1(n6507), .A2(n6359), .B1(n6506), .B2(n6358), .ZN(n6341)
         );
  AOI22_X1 U7357 ( .A1(n6463), .A2(n6361), .B1(n6508), .B2(n6360), .ZN(n6340)
         );
  OAI211_X1 U7358 ( .C1(n6365), .C2(n6342), .A(n6341), .B(n6340), .ZN(U3045)
         );
  INV_X1 U7359 ( .A(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n6345) );
  AOI22_X1 U7360 ( .A1(n6467), .A2(n6359), .B1(n6423), .B2(n6358), .ZN(n6344)
         );
  AOI22_X1 U7361 ( .A1(n6469), .A2(n6361), .B1(n6468), .B2(n6360), .ZN(n6343)
         );
  OAI211_X1 U7362 ( .C1(n6365), .C2(n6345), .A(n6344), .B(n6343), .ZN(U3046)
         );
  INV_X1 U7363 ( .A(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n6348) );
  AOI22_X1 U7364 ( .A1(n6513), .A2(n6359), .B1(n6512), .B2(n6358), .ZN(n6347)
         );
  AOI22_X1 U7365 ( .A1(n6473), .A2(n6361), .B1(n6514), .B2(n6360), .ZN(n6346)
         );
  OAI211_X1 U7366 ( .C1(n6365), .C2(n6348), .A(n6347), .B(n6346), .ZN(U3047)
         );
  INV_X1 U7367 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n6351) );
  AOI22_X1 U7368 ( .A1(n6519), .A2(n6359), .B1(n6518), .B2(n6358), .ZN(n6350)
         );
  AOI22_X1 U7369 ( .A1(n6477), .A2(n6361), .B1(n6520), .B2(n6360), .ZN(n6349)
         );
  OAI211_X1 U7370 ( .C1(n6365), .C2(n6351), .A(n6350), .B(n6349), .ZN(U3048)
         );
  INV_X1 U7371 ( .A(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n6354) );
  AOI22_X1 U7372 ( .A1(n6481), .A2(n6359), .B1(n6433), .B2(n6358), .ZN(n6353)
         );
  AOI22_X1 U7373 ( .A1(n6483), .A2(n6361), .B1(n6482), .B2(n6360), .ZN(n6352)
         );
  OAI211_X1 U7374 ( .C1(n6365), .C2(n6354), .A(n6353), .B(n6352), .ZN(U3049)
         );
  INV_X1 U7375 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6357) );
  AOI22_X1 U7376 ( .A1(n6525), .A2(n6359), .B1(n6524), .B2(n6358), .ZN(n6356)
         );
  AOI22_X1 U7377 ( .A1(n6487), .A2(n6361), .B1(n6526), .B2(n6360), .ZN(n6355)
         );
  OAI211_X1 U7378 ( .C1(n6365), .C2(n6357), .A(n6356), .B(n6355), .ZN(U3050)
         );
  INV_X1 U7379 ( .A(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n6364) );
  AOI22_X1 U7380 ( .A1(n6533), .A2(n6359), .B1(n6531), .B2(n6358), .ZN(n6363)
         );
  AOI22_X1 U7381 ( .A1(n6493), .A2(n6361), .B1(n6535), .B2(n6360), .ZN(n6362)
         );
  OAI211_X1 U7382 ( .C1(n6365), .C2(n6364), .A(n6363), .B(n6362), .ZN(U3051)
         );
  INV_X1 U7383 ( .A(n6376), .ZN(n6370) );
  INV_X1 U7384 ( .A(n6455), .ZN(n6368) );
  NAND3_X1 U7385 ( .A1(n6368), .A2(n6367), .A3(n6681), .ZN(n6369) );
  OAI21_X1 U7386 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6399) );
  NAND2_X1 U7387 ( .A1(n6372), .A2(n6416), .ZN(n6378) );
  INV_X1 U7388 ( .A(n6378), .ZN(n6398) );
  AOI22_X1 U7389 ( .A1(n6502), .A2(n6399), .B1(n6501), .B2(n6398), .ZN(n6383)
         );
  NOR3_X1 U7390 ( .A1(n6400), .A2(n6440), .A3(n6694), .ZN(n6377) );
  INV_X1 U7391 ( .A(n6374), .ZN(n6676) );
  NAND2_X1 U7392 ( .A1(n6376), .A2(n6375), .ZN(n6405) );
  OAI21_X1 U7393 ( .B1(n6377), .B2(n6676), .A(n6405), .ZN(n6381) );
  NAND2_X1 U7394 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6378), .ZN(n6379) );
  NAND4_X1 U7395 ( .A1(n6381), .A2(n6380), .A3(n6448), .A4(n6379), .ZN(n6401)
         );
  AOI22_X1 U7396 ( .A1(n6401), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6500), 
        .B2(n6400), .ZN(n6382) );
  OAI211_X1 U7397 ( .C1(n6505), .C2(n6404), .A(n6383), .B(n6382), .ZN(U3068)
         );
  AOI22_X1 U7398 ( .A1(n6508), .A2(n6399), .B1(n6507), .B2(n6398), .ZN(n6385)
         );
  AOI22_X1 U7399 ( .A1(n6401), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6506), 
        .B2(n6400), .ZN(n6384) );
  OAI211_X1 U7400 ( .C1(n6511), .C2(n6404), .A(n6385), .B(n6384), .ZN(U3069)
         );
  AOI22_X1 U7401 ( .A1(n6468), .A2(n6399), .B1(n6467), .B2(n6398), .ZN(n6387)
         );
  AOI22_X1 U7402 ( .A1(n6401), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6423), 
        .B2(n6400), .ZN(n6386) );
  OAI211_X1 U7403 ( .C1(n6388), .C2(n6404), .A(n6387), .B(n6386), .ZN(U3070)
         );
  AOI22_X1 U7404 ( .A1(n6514), .A2(n6399), .B1(n6513), .B2(n6398), .ZN(n6390)
         );
  AOI22_X1 U7405 ( .A1(n6401), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6512), 
        .B2(n6400), .ZN(n6389) );
  OAI211_X1 U7406 ( .C1(n6517), .C2(n6404), .A(n6390), .B(n6389), .ZN(U3071)
         );
  AOI22_X1 U7407 ( .A1(n6520), .A2(n6399), .B1(n6519), .B2(n6398), .ZN(n6392)
         );
  AOI22_X1 U7408 ( .A1(n6401), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6518), 
        .B2(n6400), .ZN(n6391) );
  OAI211_X1 U7409 ( .C1(n6523), .C2(n6404), .A(n6392), .B(n6391), .ZN(U3072)
         );
  AOI22_X1 U7410 ( .A1(n6482), .A2(n6399), .B1(n6481), .B2(n6398), .ZN(n6394)
         );
  AOI22_X1 U7411 ( .A1(n6401), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6433), 
        .B2(n6400), .ZN(n6393) );
  OAI211_X1 U7412 ( .C1(n6395), .C2(n6404), .A(n6394), .B(n6393), .ZN(U3073)
         );
  AOI22_X1 U7413 ( .A1(n6526), .A2(n6399), .B1(n6525), .B2(n6398), .ZN(n6397)
         );
  AOI22_X1 U7414 ( .A1(n6401), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6524), 
        .B2(n6400), .ZN(n6396) );
  OAI211_X1 U7415 ( .C1(n6529), .C2(n6404), .A(n6397), .B(n6396), .ZN(U3074)
         );
  AOI22_X1 U7416 ( .A1(n6535), .A2(n6399), .B1(n6533), .B2(n6398), .ZN(n6403)
         );
  AOI22_X1 U7417 ( .A1(n6401), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6531), 
        .B2(n6400), .ZN(n6402) );
  OAI211_X1 U7418 ( .C1(n6540), .C2(n6404), .A(n6403), .B(n6402), .ZN(U3075)
         );
  INV_X1 U7419 ( .A(n6405), .ZN(n6407) );
  INV_X1 U7420 ( .A(n6406), .ZN(n6441) );
  AOI21_X1 U7421 ( .B1(n6407), .B2(n3690), .A(n6441), .ZN(n6412) );
  NOR2_X1 U7422 ( .A1(n6412), .A2(n6694), .ZN(n6408) );
  AOI21_X1 U7423 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6416), .A(n6408), .ZN(
        n6446) );
  AOI22_X1 U7424 ( .A1(n6501), .A2(n6441), .B1(n6459), .B2(n6451), .ZN(n6418)
         );
  NOR2_X1 U7425 ( .A1(n6411), .A2(n6410), .ZN(n6672) );
  INV_X1 U7426 ( .A(n6672), .ZN(n6413) );
  NAND3_X1 U7427 ( .A1(n6413), .A2(n6674), .A3(n6412), .ZN(n6415) );
  OAI211_X1 U7428 ( .C1(n6416), .C2(n6674), .A(n6415), .B(n6414), .ZN(n6442)
         );
  AOI22_X1 U7429 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6442), .B1(n6500), 
        .B2(n6440), .ZN(n6417) );
  OAI211_X1 U7430 ( .C1(n6446), .C2(n6419), .A(n6418), .B(n6417), .ZN(U3076)
         );
  AOI22_X1 U7431 ( .A1(n6507), .A2(n6441), .B1(n6463), .B2(n6451), .ZN(n6421)
         );
  AOI22_X1 U7432 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6442), .B1(n6506), 
        .B2(n6440), .ZN(n6420) );
  OAI211_X1 U7433 ( .C1(n6446), .C2(n6422), .A(n6421), .B(n6420), .ZN(U3077)
         );
  AOI22_X1 U7434 ( .A1(n6467), .A2(n6441), .B1(n6423), .B2(n6440), .ZN(n6425)
         );
  AOI22_X1 U7435 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6442), .B1(n6469), 
        .B2(n6451), .ZN(n6424) );
  OAI211_X1 U7436 ( .C1(n6446), .C2(n6426), .A(n6425), .B(n6424), .ZN(U3078)
         );
  AOI22_X1 U7437 ( .A1(n6513), .A2(n6441), .B1(n6473), .B2(n6451), .ZN(n6428)
         );
  AOI22_X1 U7438 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6442), .B1(n6512), 
        .B2(n6440), .ZN(n6427) );
  OAI211_X1 U7439 ( .C1(n6446), .C2(n6429), .A(n6428), .B(n6427), .ZN(U3079)
         );
  AOI22_X1 U7440 ( .A1(n6519), .A2(n6441), .B1(n6477), .B2(n6451), .ZN(n6431)
         );
  AOI22_X1 U7441 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6442), .B1(n6518), 
        .B2(n6440), .ZN(n6430) );
  OAI211_X1 U7442 ( .C1(n6446), .C2(n6432), .A(n6431), .B(n6430), .ZN(U3080)
         );
  AOI22_X1 U7443 ( .A1(n6481), .A2(n6441), .B1(n6433), .B2(n6440), .ZN(n6435)
         );
  AOI22_X1 U7444 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6442), .B1(n6483), 
        .B2(n6451), .ZN(n6434) );
  OAI211_X1 U7445 ( .C1(n6446), .C2(n6436), .A(n6435), .B(n6434), .ZN(U3081)
         );
  AOI22_X1 U7446 ( .A1(n6525), .A2(n6441), .B1(n6487), .B2(n6451), .ZN(n6438)
         );
  AOI22_X1 U7447 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6442), .B1(n6524), 
        .B2(n6440), .ZN(n6437) );
  OAI211_X1 U7448 ( .C1(n6446), .C2(n6439), .A(n6438), .B(n6437), .ZN(U3082)
         );
  AOI22_X1 U7449 ( .A1(n6533), .A2(n6441), .B1(n6531), .B2(n6440), .ZN(n6444)
         );
  AOI22_X1 U7450 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6442), .B1(n6493), 
        .B2(n6451), .ZN(n6443) );
  OAI211_X1 U7451 ( .C1(n6446), .C2(n6445), .A(n6444), .B(n6443), .ZN(U3083)
         );
  OAI22_X1 U7452 ( .A1(n6449), .A2(n6453), .B1(n6448), .B2(n6447), .ZN(n6492)
         );
  NOR2_X1 U7453 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6450), .ZN(n6491)
         );
  AOI22_X1 U7454 ( .A1(n6502), .A2(n6492), .B1(n6501), .B2(n6491), .ZN(n6461)
         );
  OAI21_X1 U7455 ( .B1(n6494), .B2(n6451), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6452) );
  OAI211_X1 U7456 ( .C1(n6454), .C2(n6453), .A(n6452), .B(n6674), .ZN(n6458)
         );
  OR2_X1 U7457 ( .A1(n6662), .A2(n6491), .ZN(n6457) );
  NAND4_X1 U7458 ( .A1(n6458), .A2(n6457), .A3(n6456), .A4(n6455), .ZN(n6495)
         );
  AOI22_X1 U7459 ( .A1(n6495), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n6494), 
        .B2(n6459), .ZN(n6460) );
  OAI211_X1 U7460 ( .C1(n6462), .C2(n6498), .A(n6461), .B(n6460), .ZN(U3084)
         );
  AOI22_X1 U7461 ( .A1(n6508), .A2(n6492), .B1(n6507), .B2(n6491), .ZN(n6465)
         );
  AOI22_X1 U7462 ( .A1(n6495), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6494), 
        .B2(n6463), .ZN(n6464) );
  OAI211_X1 U7463 ( .C1(n6466), .C2(n6498), .A(n6465), .B(n6464), .ZN(U3085)
         );
  AOI22_X1 U7464 ( .A1(n6468), .A2(n6492), .B1(n6467), .B2(n6491), .ZN(n6471)
         );
  AOI22_X1 U7465 ( .A1(n6495), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n6494), 
        .B2(n6469), .ZN(n6470) );
  OAI211_X1 U7466 ( .C1(n6472), .C2(n6498), .A(n6471), .B(n6470), .ZN(U3086)
         );
  AOI22_X1 U7467 ( .A1(n6514), .A2(n6492), .B1(n6513), .B2(n6491), .ZN(n6475)
         );
  AOI22_X1 U7468 ( .A1(n6495), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6494), 
        .B2(n6473), .ZN(n6474) );
  OAI211_X1 U7469 ( .C1(n6476), .C2(n6498), .A(n6475), .B(n6474), .ZN(U3087)
         );
  AOI22_X1 U7470 ( .A1(n6520), .A2(n6492), .B1(n6519), .B2(n6491), .ZN(n6479)
         );
  AOI22_X1 U7471 ( .A1(n6495), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n6494), 
        .B2(n6477), .ZN(n6478) );
  OAI211_X1 U7472 ( .C1(n6480), .C2(n6498), .A(n6479), .B(n6478), .ZN(U3088)
         );
  AOI22_X1 U7473 ( .A1(n6482), .A2(n6492), .B1(n6481), .B2(n6491), .ZN(n6485)
         );
  AOI22_X1 U7474 ( .A1(n6495), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n6494), 
        .B2(n6483), .ZN(n6484) );
  OAI211_X1 U7475 ( .C1(n6486), .C2(n6498), .A(n6485), .B(n6484), .ZN(U3089)
         );
  AOI22_X1 U7476 ( .A1(n6526), .A2(n6492), .B1(n6525), .B2(n6491), .ZN(n6489)
         );
  AOI22_X1 U7477 ( .A1(n6495), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n6494), 
        .B2(n6487), .ZN(n6488) );
  OAI211_X1 U7478 ( .C1(n6490), .C2(n6498), .A(n6489), .B(n6488), .ZN(U3090)
         );
  AOI22_X1 U7479 ( .A1(n6535), .A2(n6492), .B1(n6533), .B2(n6491), .ZN(n6497)
         );
  AOI22_X1 U7480 ( .A1(n6495), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n6494), 
        .B2(n6493), .ZN(n6496) );
  OAI211_X1 U7481 ( .C1(n6499), .C2(n6498), .A(n6497), .B(n6496), .ZN(U3091)
         );
  AOI22_X1 U7482 ( .A1(n6501), .A2(n6532), .B1(n6500), .B2(n6530), .ZN(n6504)
         );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6536), .B1(n6502), 
        .B2(n6534), .ZN(n6503) );
  OAI211_X1 U7484 ( .C1(n6505), .C2(n6539), .A(n6504), .B(n6503), .ZN(U3108)
         );
  AOI22_X1 U7485 ( .A1(n6507), .A2(n6532), .B1(n6506), .B2(n6530), .ZN(n6510)
         );
  AOI22_X1 U7486 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6536), .B1(n6508), 
        .B2(n6534), .ZN(n6509) );
  OAI211_X1 U7487 ( .C1(n6511), .C2(n6539), .A(n6510), .B(n6509), .ZN(U3109)
         );
  AOI22_X1 U7488 ( .A1(n6513), .A2(n6532), .B1(n6512), .B2(n6530), .ZN(n6516)
         );
  AOI22_X1 U7489 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6536), .B1(n6514), 
        .B2(n6534), .ZN(n6515) );
  OAI211_X1 U7490 ( .C1(n6517), .C2(n6539), .A(n6516), .B(n6515), .ZN(U3111)
         );
  AOI22_X1 U7491 ( .A1(n6519), .A2(n6532), .B1(n6518), .B2(n6530), .ZN(n6522)
         );
  AOI22_X1 U7492 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6536), .B1(n6520), 
        .B2(n6534), .ZN(n6521) );
  OAI211_X1 U7493 ( .C1(n6523), .C2(n6539), .A(n6522), .B(n6521), .ZN(U3112)
         );
  AOI22_X1 U7494 ( .A1(n6525), .A2(n6532), .B1(n6524), .B2(n6530), .ZN(n6528)
         );
  AOI22_X1 U7495 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6536), .B1(n6526), 
        .B2(n6534), .ZN(n6527) );
  OAI211_X1 U7496 ( .C1(n6529), .C2(n6539), .A(n6528), .B(n6527), .ZN(U3114)
         );
  AOI22_X1 U7497 ( .A1(n6533), .A2(n6532), .B1(n6531), .B2(n6530), .ZN(n6538)
         );
  AOI22_X1 U7498 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6536), .B1(n6535), 
        .B2(n6534), .ZN(n6537) );
  OAI211_X1 U7499 ( .C1(n6540), .C2(n6539), .A(n6538), .B(n6537), .ZN(U3115)
         );
  AOI22_X1 U7500 ( .A1(n3690), .A2(n6542), .B1(n6541), .B2(n3183), .ZN(n6666)
         );
  NAND2_X1 U7501 ( .A1(n6543), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6671) );
  AND3_X1 U7502 ( .A1(n6666), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6671), 
        .ZN(n6548) );
  AOI21_X1 U7503 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6548), .A(n6544), 
        .ZN(n6545) );
  NAND2_X1 U7504 ( .A1(n6546), .A2(n6545), .ZN(n6547) );
  OAI21_X1 U7505 ( .B1(n6548), .B2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n6547), 
        .ZN(n6549) );
  AOI222_X1 U7506 ( .A1(n6762), .A2(n6550), .B1(n6762), .B2(n6549), .C1(n6550), 
        .C2(n6549), .ZN(n6553) );
  OR2_X1 U7507 ( .A1(n6553), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6552)
         );
  NAND2_X1 U7508 ( .A1(n6552), .A2(n6551), .ZN(n6556) );
  NAND2_X1 U7509 ( .A1(n6553), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6555) );
  NAND3_X1 U7510 ( .A1(n6556), .A2(n6555), .A3(n6554), .ZN(n6566) );
  NOR2_X1 U7511 ( .A1(n6558), .A2(n6557), .ZN(n6561) );
  OAI21_X1 U7512 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6559), 
        .ZN(n6560) );
  NAND3_X1 U7513 ( .A1(n6562), .A2(n6561), .A3(n6560), .ZN(n6563) );
  NOR2_X1 U7514 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  NAND2_X1 U7515 ( .A1(n6582), .A2(n6583), .ZN(n6569) );
  NAND2_X1 U7516 ( .A1(READY_N), .A2(n6567), .ZN(n6568) );
  NAND2_X1 U7517 ( .A1(n6569), .A2(n6568), .ZN(n6573) );
  OR2_X1 U7518 ( .A1(n6571), .A2(n6570), .ZN(n6572) );
  OAI21_X1 U7519 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4495), .A(n6661), .ZN(
        n6585) );
  AOI221_X1 U7520 ( .B1(n6575), .B2(STATE2_REG_0__SCAN_IN), .C1(n6585), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6574), .ZN(n6580) );
  OAI211_X1 U7521 ( .C1(n6578), .C2(n6577), .A(n6576), .B(n6661), .ZN(n6579)
         );
  OAI211_X1 U7522 ( .C1(n6582), .C2(n6581), .A(n6580), .B(n6579), .ZN(U3148)
         );
  AOI21_X1 U7523 ( .B1(n6584), .B2(n4495), .A(n6583), .ZN(n6588) );
  OAI211_X1 U7524 ( .C1(STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_2__SCAN_IN), 
        .A(STATE2_REG_1__SCAN_IN), .B(n6585), .ZN(n6586) );
  OAI211_X1 U7525 ( .C1(n6589), .C2(n6588), .A(n6587), .B(n6586), .ZN(U3149)
         );
  OAI221_X1 U7526 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(n4495), .A(n6660), .ZN(n6591) );
  OAI21_X1 U7527 ( .B1(n6701), .B2(n6591), .A(n6590), .ZN(U3150) );
  INV_X1 U7528 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6828) );
  NOR2_X1 U7529 ( .A1(n6659), .A2(n6828), .ZN(U3151) );
  AND2_X1 U7530 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6592), .ZN(U3152) );
  AND2_X1 U7531 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6592), .ZN(U3153) );
  AND2_X1 U7532 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6592), .ZN(U3154) );
  AND2_X1 U7533 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6592), .ZN(U3155) );
  INV_X1 U7534 ( .A(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6974) );
  NOR2_X1 U7535 ( .A1(n6659), .A2(n6974), .ZN(U3156) );
  AND2_X1 U7536 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6592), .ZN(U3157) );
  AND2_X1 U7537 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6592), .ZN(U3158) );
  AND2_X1 U7538 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6592), .ZN(U3159) );
  AND2_X1 U7539 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6592), .ZN(U3160) );
  AND2_X1 U7540 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6592), .ZN(U3161) );
  AND2_X1 U7541 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6592), .ZN(U3162) );
  AND2_X1 U7542 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6592), .ZN(U3163) );
  AND2_X1 U7543 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6592), .ZN(U3164) );
  AND2_X1 U7544 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6592), .ZN(U3165) );
  AND2_X1 U7545 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6592), .ZN(U3166) );
  AND2_X1 U7546 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6592), .ZN(U3167) );
  AND2_X1 U7547 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6592), .ZN(U3168) );
  AND2_X1 U7548 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6592), .ZN(U3169) );
  INV_X1 U7549 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U7550 ( .A1(n6659), .A2(n6925), .ZN(U3170) );
  AND2_X1 U7551 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6592), .ZN(U3171) );
  AND2_X1 U7552 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6592), .ZN(U3172) );
  AND2_X1 U7553 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6592), .ZN(U3173) );
  INV_X1 U7554 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6819) );
  NOR2_X1 U7555 ( .A1(n6659), .A2(n6819), .ZN(U3174) );
  AND2_X1 U7556 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6592), .ZN(U3175) );
  AND2_X1 U7557 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6592), .ZN(U3176) );
  AND2_X1 U7558 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6592), .ZN(U3177) );
  AND2_X1 U7559 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6592), .ZN(U3178) );
  AND2_X1 U7560 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6592), .ZN(U3179) );
  AND2_X1 U7561 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6592), .ZN(U3180) );
  NOR2_X1 U7562 ( .A1(n6838), .A2(n6593), .ZN(n6599) );
  AOI22_X1 U7563 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6610) );
  OAI221_X1 U7564 ( .B1(n6593), .B2(NA_N), .C1(n6593), .C2(n6838), .A(n6777), 
        .ZN(n6607) );
  AND2_X1 U7565 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6596) );
  INV_X1 U7566 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6595) );
  OAI21_X1 U7567 ( .B1(n6596), .B2(n6595), .A(n6656), .ZN(n6594) );
  OAI211_X1 U7568 ( .C1(n6599), .C2(n6610), .A(n6607), .B(n6594), .ZN(U3181)
         );
  NOR2_X1 U7569 ( .A1(n6777), .A2(n6595), .ZN(n6603) );
  NAND2_X1 U7570 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6601) );
  OAI21_X1 U7571 ( .B1(n6603), .B2(n6596), .A(n6601), .ZN(n6597) );
  OAI211_X1 U7572 ( .C1(n6838), .C2(n4495), .A(n6598), .B(n6597), .ZN(U3182)
         );
  INV_X1 U7573 ( .A(n6599), .ZN(n6609) );
  NOR2_X1 U7574 ( .A1(NA_N), .A2(n4495), .ZN(n6600) );
  OAI21_X1 U7575 ( .B1(n6600), .B2(n6838), .A(HOLD), .ZN(n6602) );
  OAI211_X1 U7576 ( .C1(REQUESTPENDING_REG_SCAN_IN), .C2(n6602), .A(
        STATE_REG_0__SCAN_IN), .B(n6601), .ZN(n6606) );
  INV_X1 U7577 ( .A(n6603), .ZN(n6604) );
  NOR4_X1 U7578 ( .A1(NA_N), .A2(n6838), .A3(n4495), .A4(n6604), .ZN(n6605) );
  AOI21_X1 U7579 ( .B1(n6607), .B2(n6606), .A(n6605), .ZN(n6608) );
  OAI21_X1 U7580 ( .B1(n6610), .B2(n6609), .A(n6608), .ZN(U3183) );
  INV_X1 U7581 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U7582 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6706), .ZN(n6653) );
  INV_X1 U7583 ( .A(n6653), .ZN(n6646) );
  AOI22_X1 U7584 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6656), .ZN(n6611) );
  OAI21_X1 U7585 ( .B1(n6612), .B2(n6648), .A(n6611), .ZN(U3184) );
  AOI22_X1 U7586 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6656), .ZN(n6613) );
  OAI21_X1 U7587 ( .B1(n6753), .B2(n6648), .A(n6613), .ZN(U3185) );
  AOI22_X1 U7588 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6656), .ZN(n6614) );
  OAI21_X1 U7589 ( .B1(n6615), .B2(n6648), .A(n6614), .ZN(U3186) );
  AOI22_X1 U7590 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6656), .ZN(n6616) );
  OAI21_X1 U7591 ( .B1(n6897), .B2(n6648), .A(n6616), .ZN(U3187) );
  AOI22_X1 U7592 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6656), .ZN(n6617) );
  OAI21_X1 U7593 ( .B1(n6619), .B2(n6648), .A(n6617), .ZN(U3188) );
  AOI22_X1 U7594 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6656), .ZN(n6618) );
  OAI21_X1 U7595 ( .B1(n6619), .B2(n6653), .A(n6618), .ZN(U3189) );
  AOI22_X1 U7596 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6656), .ZN(n6620) );
  OAI21_X1 U7597 ( .B1(n6621), .B2(n6648), .A(n6620), .ZN(U3190) );
  INV_X1 U7598 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6821) );
  AOI22_X1 U7599 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6656), .ZN(n6622) );
  OAI21_X1 U7600 ( .B1(n6821), .B2(n6648), .A(n6622), .ZN(U3191) );
  AOI22_X1 U7601 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6656), .ZN(n6623) );
  OAI21_X1 U7602 ( .B1(n6821), .B2(n6653), .A(n6623), .ZN(U3192) );
  AOI22_X1 U7603 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6656), .ZN(n6624) );
  OAI21_X1 U7604 ( .B1(n6625), .B2(n6648), .A(n6624), .ZN(U3193) );
  AOI22_X1 U7605 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6656), .ZN(n6626) );
  OAI21_X1 U7606 ( .B1(n6628), .B2(n6648), .A(n6626), .ZN(U3194) );
  AOI22_X1 U7607 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6656), .ZN(n6627) );
  OAI21_X1 U7608 ( .B1(n6628), .B2(n6653), .A(n6627), .ZN(U3195) );
  INV_X1 U7609 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n6948) );
  OAI222_X1 U7610 ( .A1(n6653), .A2(n6629), .B1(n6948), .B2(n6706), .C1(n6883), 
        .C2(n6648), .ZN(U3196) );
  AOI22_X1 U7611 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6656), .ZN(n6630) );
  OAI21_X1 U7612 ( .B1(n6883), .B2(n6653), .A(n6630), .ZN(U3197) );
  AOI22_X1 U7613 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6656), .ZN(n6631) );
  OAI21_X1 U7614 ( .B1(n6633), .B2(n6648), .A(n6631), .ZN(U3198) );
  AOI22_X1 U7615 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6656), .ZN(n6632) );
  OAI21_X1 U7616 ( .B1(n6633), .B2(n6653), .A(n6632), .ZN(U3199) );
  AOI222_X1 U7617 ( .A1(n6651), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6656), .C1(REIP_REG_17__SCAN_IN), .C2(
        n6646), .ZN(n6634) );
  INV_X1 U7618 ( .A(n6634), .ZN(U3200) );
  INV_X1 U7619 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6946) );
  OAI222_X1 U7620 ( .A1(n6653), .A2(n6635), .B1(n6946), .B2(n6706), .C1(n6636), 
        .C2(n6648), .ZN(U3201) );
  INV_X1 U7621 ( .A(ADDRESS_REG_18__SCAN_IN), .ZN(n6771) );
  OAI222_X1 U7622 ( .A1(n6653), .A2(n6636), .B1(n6771), .B2(n6706), .C1(n6637), 
        .C2(n6648), .ZN(U3202) );
  INV_X1 U7623 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6825) );
  OAI222_X1 U7624 ( .A1(n6653), .A2(n6637), .B1(n6825), .B2(n6706), .C1(n5543), 
        .C2(n6648), .ZN(U3203) );
  INV_X1 U7625 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6640) );
  AOI22_X1 U7626 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6656), .ZN(n6638) );
  OAI21_X1 U7627 ( .B1(n6640), .B2(n6648), .A(n6638), .ZN(U3204) );
  AOI22_X1 U7628 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6656), .ZN(n6639) );
  OAI21_X1 U7629 ( .B1(n6640), .B2(n6653), .A(n6639), .ZN(U3205) );
  AOI22_X1 U7630 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6656), .ZN(n6641) );
  OAI21_X1 U7631 ( .B1(n4321), .B2(n6648), .A(n6641), .ZN(U3206) );
  INV_X1 U7632 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6919) );
  OAI222_X1 U7633 ( .A1(n6648), .A2(n6643), .B1(n6919), .B2(n6706), .C1(n4321), 
        .C2(n6653), .ZN(U3207) );
  AOI22_X1 U7634 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6656), .ZN(n6642) );
  OAI21_X1 U7635 ( .B1(n6643), .B2(n6653), .A(n6642), .ZN(U3208) );
  AOI22_X1 U7636 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6656), .ZN(n6644) );
  OAI21_X1 U7637 ( .B1(n6805), .B2(n6653), .A(n6644), .ZN(U3209) );
  AOI22_X1 U7638 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6656), .ZN(n6645) );
  OAI21_X1 U7639 ( .B1(n6807), .B2(n6648), .A(n6645), .ZN(U3210) );
  AOI22_X1 U7640 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6646), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6656), .ZN(n6647) );
  OAI21_X1 U7641 ( .B1(n6650), .B2(n6648), .A(n6647), .ZN(U3211) );
  AOI22_X1 U7642 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6656), .ZN(n6649) );
  OAI21_X1 U7643 ( .B1(n6650), .B2(n6653), .A(n6649), .ZN(U3212) );
  INV_X1 U7644 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6654) );
  AOI22_X1 U7645 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6651), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6656), .ZN(n6652) );
  OAI21_X1 U7646 ( .B1(n6654), .B2(n6653), .A(n6652), .ZN(U3213) );
  OAI22_X1 U7647 ( .A1(n6656), .A2(BYTEENABLE_REG_3__SCAN_IN), .B1(
        BE_N_REG_3__SCAN_IN), .B2(n6706), .ZN(n6655) );
  INV_X1 U7648 ( .A(n6655), .ZN(U3445) );
  MUX2_X1 U7649 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6656), .Z(U3446) );
  MUX2_X1 U7650 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6656), .Z(U3447) );
  INV_X1 U7651 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6689) );
  INV_X1 U7652 ( .A(BE_N_REG_0__SCAN_IN), .ZN(n6967) );
  AOI22_X1 U7653 ( .A1(n6706), .A2(n6689), .B1(n6967), .B2(n6656), .ZN(U3448)
         );
  OAI21_X1 U7654 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6659), .A(n6658), .ZN(
        n6657) );
  INV_X1 U7655 ( .A(n6657), .ZN(U3451) );
  INV_X1 U7656 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6684) );
  OAI21_X1 U7657 ( .B1(n6659), .B2(n6684), .A(n6658), .ZN(U3452) );
  OAI221_X1 U7658 ( .B1(n6662), .B2(STATE2_REG_0__SCAN_IN), .C1(n6662), .C2(
        n6661), .A(n6660), .ZN(U3453) );
  AOI211_X1 U7659 ( .C1(STATE2_REG_1__SCAN_IN), .C2(n4528), .A(n6664), .B(
        n6663), .ZN(n6665) );
  OAI21_X1 U7660 ( .B1(n6666), .B2(n6670), .A(n6665), .ZN(n6667) );
  OAI21_X1 U7661 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6668), .A(n6667), 
        .ZN(n6669) );
  OAI21_X1 U7662 ( .B1(n6671), .B2(n6670), .A(n6669), .ZN(U3461) );
  OR2_X1 U7663 ( .A1(n6673), .A2(n6672), .ZN(n6675) );
  AOI222_X1 U7664 ( .A1(n6678), .A2(n6677), .B1(n3682), .B2(n6676), .C1(n6675), 
        .C2(n6674), .ZN(n6680) );
  AOI22_X1 U7665 ( .A1(n6682), .A2(n6681), .B1(n6680), .B2(n6679), .ZN(U3462)
         );
  INV_X1 U7666 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6855) );
  AOI221_X1 U7667 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n4473), .C1(n6855), 
        .C2(n6684), .A(n6683), .ZN(n6688) );
  OAI22_X1 U7668 ( .A1(n6686), .A2(BYTEENABLE_REG_2__SCAN_IN), .B1(n5117), 
        .B2(n6685), .ZN(n6687) );
  NOR2_X1 U7669 ( .A1(n6688), .A2(n6687), .ZN(U3468) );
  AOI22_X1 U7670 ( .A1(n6691), .A2(n4473), .B1(n6690), .B2(n6689), .ZN(U3469)
         );
  NAND2_X1 U7671 ( .A1(n6656), .A2(W_R_N_REG_SCAN_IN), .ZN(n6692) );
  OAI21_X1 U7672 ( .B1(n6656), .B2(READREQUEST_REG_SCAN_IN), .A(n6692), .ZN(
        U3470) );
  INV_X1 U7673 ( .A(n6693), .ZN(n6698) );
  OAI211_X1 U7674 ( .C1(n6696), .C2(READY_N), .A(n6695), .B(n6694), .ZN(n6697)
         );
  NOR2_X1 U7675 ( .A1(n6698), .A2(n6697), .ZN(n6705) );
  OAI211_X1 U7676 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6700), .A(n6699), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6702) );
  AOI21_X1 U7677 ( .B1(n6702), .B2(STATE2_REG_0__SCAN_IN), .A(n6701), .ZN(
        n6704) );
  NAND2_X1 U7678 ( .A1(n6705), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6703) );
  OAI21_X1 U7679 ( .B1(n6705), .B2(n6704), .A(n6703), .ZN(U3472) );
  OAI22_X1 U7680 ( .A1(n6656), .A2(MEMORYFETCH_REG_SCAN_IN), .B1(
        M_IO_N_REG_SCAN_IN), .B2(n6706), .ZN(n6707) );
  INV_X1 U7681 ( .A(n6707), .ZN(U3473) );
  INV_X1 U7682 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6898) );
  NOR4_X1 U7683 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(
        INSTQUEUE_REG_11__5__SCAN_IN), .A3(n6885), .A4(n6898), .ZN(n6717) );
  NOR4_X1 U7684 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(
        INSTQUEUE_REG_3__0__SCAN_IN), .A3(INSTQUEUE_REG_6__0__SCAN_IN), .A4(
        n5015), .ZN(n6716) );
  NAND4_X1 U7685 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6918), .A3(n6949), .A4(n6871), .ZN(n6708) );
  NOR4_X1 U7686 ( .A1(EBX_REG_5__SCAN_IN), .A2(EBX_REG_2__SCAN_IN), .A3(n6709), 
        .A4(n6708), .ZN(n6715) );
  NAND4_X1 U7687 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(
        EAX_REG_10__SCAN_IN), .A3(PHYADDRPOINTER_REG_0__SCAN_IN), .A4(n6762), 
        .ZN(n6713) );
  INV_X1 U7688 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6900) );
  NAND4_X1 U7689 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(
        INSTQUEUE_REG_14__5__SCAN_IN), .A3(n4898), .A4(n6900), .ZN(n6712) );
  NAND4_X1 U7690 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .A3(PHYADDRPOINTER_REG_22__SCAN_IN), 
        .A4(REIP_REG_14__SCAN_IN), .ZN(n6711) );
  NAND4_X1 U7691 ( .A1(EBX_REG_28__SCAN_IN), .A2(EBX_REG_0__SCAN_IN), .A3(
        CODEFETCH_REG_SCAN_IN), .A4(D_C_N_REG_SCAN_IN), .ZN(n6710) );
  NOR4_X1 U7692 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6714)
         );
  NAND4_X1 U7693 ( .A1(n6717), .A2(n6716), .A3(n6715), .A4(n6714), .ZN(n6751)
         );
  NOR4_X1 U7694 ( .A1(EBX_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .A3(REIP_REG_3__SCAN_IN), .A4(
        DATAWIDTH_REG_0__SCAN_IN), .ZN(n6721) );
  NOR4_X1 U7695 ( .A1(DATAO_REG_10__SCAN_IN), .A2(DATAO_REG_19__SCAN_IN), .A3(
        UWORD_REG_5__SCAN_IN), .A4(DATAO_REG_21__SCAN_IN), .ZN(n6720) );
  NOR4_X1 U7696 ( .A1(EAX_REG_30__SCAN_IN), .A2(EAX_REG_27__SCAN_IN), .A3(
        DATAI_25_), .A4(DATAI_6_), .ZN(n6719) );
  NOR4_X1 U7697 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .A3(EAX_REG_19__SCAN_IN), .A4(
        DATAI_5_), .ZN(n6718) );
  NAND4_X1 U7698 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6750)
         );
  NOR4_X1 U7699 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(ADDRESS_REG_18__SCAN_IN), 
        .A3(DATAO_REG_26__SCAN_IN), .A4(DATAO_REG_27__SCAN_IN), .ZN(n6725) );
  NOR4_X1 U7700 ( .A1(DATAO_REG_22__SCAN_IN), .A2(DATAO_REG_25__SCAN_IN), .A3(
        ADDRESS_REG_17__SCAN_IN), .A4(ADDRESS_REG_16__SCAN_IN), .ZN(n6724) );
  NOR4_X1 U7701 ( .A1(LWORD_REG_11__SCAN_IN), .A2(LWORD_REG_7__SCAN_IN), .A3(
        UWORD_REG_2__SCAN_IN), .A4(DATAO_REG_5__SCAN_IN), .ZN(n6723) );
  NOR4_X1 U7702 ( .A1(READY_N), .A2(DATAWIDTH_REG_12__SCAN_IN), .A3(
        DATAWIDTH_REG_31__SCAN_IN), .A4(M_IO_N_REG_SCAN_IN), .ZN(n6722) );
  NAND4_X1 U7703 ( .A1(n6725), .A2(n6724), .A3(n6723), .A4(n6722), .ZN(n6749)
         );
  INV_X1 U7704 ( .A(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n6931) );
  NOR4_X1 U7705 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6931), .A3(n6656), 
        .A4(n6726), .ZN(n6746) );
  INV_X1 U7706 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6791) );
  INV_X1 U7707 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6757) );
  NOR4_X1 U7708 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(
        INSTQUEUE_REG_8__6__SCAN_IN), .A3(n6757), .A4(n6840), .ZN(n6727) );
  NAND3_X1 U7709 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(
        INSTQUEUE_REG_2__6__SCAN_IN), .A3(n6727), .ZN(n6733) );
  INV_X1 U7710 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6800) );
  NOR4_X1 U7711 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(
        INSTQUEUE_REG_12__7__SCAN_IN), .A3(n6818), .A4(n6800), .ZN(n6731) );
  INV_X1 U7712 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6775) );
  NOR4_X1 U7713 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(
        INSTQUEUE_REG_9__4__SCAN_IN), .A3(INSTQUEUE_REG_15__4__SCAN_IN), .A4(
        n6775), .ZN(n6730) );
  INV_X1 U7714 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n6873) );
  NOR4_X1 U7715 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(
        INSTQUEUE_REG_2__1__SCAN_IN), .A3(n4905), .A4(n6873), .ZN(n6729) );
  NOR4_X1 U7716 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(
        INSTQUEUE_REG_4__1__SCAN_IN), .A3(PHYADDRPOINTER_REG_4__SCAN_IN), .A4(
        n6778), .ZN(n6728) );
  NAND4_X1 U7717 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6732)
         );
  NOR4_X1 U7718 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6791), .A3(n6733), 
        .A4(n6732), .ZN(n6745) );
  NOR4_X1 U7719 ( .A1(LWORD_REG_14__SCAN_IN), .A2(ADS_N_REG_SCAN_IN), .A3(
        DATAO_REG_8__SCAN_IN), .A4(n6996), .ZN(n6734) );
  NAND3_X1 U7720 ( .A1(DATAO_REG_2__SCAN_IN), .A2(DATAO_REG_13__SCAN_IN), .A3(
        n6734), .ZN(n6743) );
  NAND4_X1 U7721 ( .A1(BE_N_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), 
        .A3(DATAO_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_26__SCAN_IN), .ZN(n6735)
         );
  NOR3_X1 U7722 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(DATAI_31_), .A3(
        n6735), .ZN(n6741) );
  NAND4_X1 U7723 ( .A1(EBX_REG_20__SCAN_IN), .A2(DATAI_4_), .A3(n6805), .A4(
        n4045), .ZN(n6739) );
  NAND4_X1 U7724 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(
        REIP_REG_31__SCAN_IN), .A3(REIP_REG_28__SCAN_IN), .A4(DATAI_7_), .ZN(
        n6738) );
  NAND4_X1 U7725 ( .A1(BE_N_REG_3__SCAN_IN), .A2(LWORD_REG_6__SCAN_IN), .A3(
        LWORD_REG_8__SCAN_IN), .A4(DATAO_REG_3__SCAN_IN), .ZN(n6737) );
  NAND4_X1 U7726 ( .A1(ADDRESS_REG_12__SCAN_IN), .A2(DATAO_REG_17__SCAN_IN), 
        .A3(ADDRESS_REG_23__SCAN_IN), .A4(UWORD_REG_11__SCAN_IN), .ZN(n6736)
         );
  NOR4_X1 U7727 ( .A1(n6739), .A2(n6738), .A3(n6737), .A4(n6736), .ZN(n6740)
         );
  INV_X1 U7728 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n6793) );
  NAND4_X1 U7729 ( .A1(n6741), .A2(n6740), .A3(n6793), .A4(n6977), .ZN(n6742)
         );
  NOR4_X1 U7730 ( .A1(n6888), .A2(n6897), .A3(n6743), .A4(n6742), .ZN(n6744)
         );
  NAND4_X1 U7731 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6748)
         );
  NOR4_X1 U7732 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n7013)
         );
  INV_X1 U7733 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6754) );
  AOI22_X1 U7734 ( .A1(n6754), .A2(keyinput63), .B1(keyinput42), .B2(n6753), 
        .ZN(n6752) );
  OAI221_X1 U7735 ( .B1(n6754), .B2(keyinput63), .C1(n6753), .C2(keyinput42), 
        .A(n6752), .ZN(n6766) );
  AOI22_X1 U7736 ( .A1(n6757), .A2(keyinput127), .B1(keyinput65), .B2(n6756), 
        .ZN(n6755) );
  OAI221_X1 U7737 ( .B1(n6757), .B2(keyinput127), .C1(n6756), .C2(keyinput65), 
        .A(n6755), .ZN(n6765) );
  AOI22_X1 U7738 ( .A1(n4045), .A2(keyinput37), .B1(n6759), .B2(keyinput78), 
        .ZN(n6758) );
  OAI221_X1 U7739 ( .B1(n4045), .B2(keyinput37), .C1(n6759), .C2(keyinput78), 
        .A(n6758), .ZN(n6764) );
  AOI22_X1 U7740 ( .A1(n6762), .A2(keyinput38), .B1(keyinput24), .B2(n6761), 
        .ZN(n6760) );
  OAI221_X1 U7741 ( .B1(n6762), .B2(keyinput38), .C1(n6761), .C2(keyinput24), 
        .A(n6760), .ZN(n6763) );
  NOR4_X1 U7742 ( .A1(n6766), .A2(n6765), .A3(n6764), .A4(n6763), .ZN(n6816)
         );
  INV_X1 U7743 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6769) );
  AOI22_X1 U7744 ( .A1(n6769), .A2(keyinput83), .B1(n6768), .B2(keyinput69), 
        .ZN(n6767) );
  OAI221_X1 U7745 ( .B1(n6769), .B2(keyinput83), .C1(n6768), .C2(keyinput69), 
        .A(n6767), .ZN(n6782) );
  AOI22_X1 U7746 ( .A1(n6772), .A2(keyinput0), .B1(keyinput124), .B2(n6771), 
        .ZN(n6770) );
  OAI221_X1 U7747 ( .B1(n6772), .B2(keyinput0), .C1(n6771), .C2(keyinput124), 
        .A(n6770), .ZN(n6781) );
  AOI22_X1 U7748 ( .A1(n6775), .A2(keyinput72), .B1(keyinput74), .B2(n6774), 
        .ZN(n6773) );
  OAI221_X1 U7749 ( .B1(n6775), .B2(keyinput72), .C1(n6774), .C2(keyinput74), 
        .A(n6773), .ZN(n6780) );
  AOI22_X1 U7750 ( .A1(n6778), .A2(keyinput87), .B1(n6777), .B2(keyinput55), 
        .ZN(n6776) );
  OAI221_X1 U7751 ( .B1(n6778), .B2(keyinput87), .C1(n6777), .C2(keyinput55), 
        .A(n6776), .ZN(n6779) );
  NOR4_X1 U7752 ( .A1(n6782), .A2(n6781), .A3(n6780), .A4(n6779), .ZN(n6815)
         );
  INV_X1 U7753 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6785) );
  INV_X1 U7754 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6784) );
  AOI22_X1 U7755 ( .A1(n6785), .A2(keyinput68), .B1(n6784), .B2(keyinput20), 
        .ZN(n6783) );
  OAI221_X1 U7756 ( .B1(n6785), .B2(keyinput68), .C1(n6784), .C2(keyinput20), 
        .A(n6783), .ZN(n6798) );
  AOI22_X1 U7757 ( .A1(n6788), .A2(keyinput56), .B1(keyinput101), .B2(n6787), 
        .ZN(n6786) );
  OAI221_X1 U7758 ( .B1(n6788), .B2(keyinput56), .C1(n6787), .C2(keyinput101), 
        .A(n6786), .ZN(n6797) );
  INV_X1 U7759 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6790) );
  AOI22_X1 U7760 ( .A1(n6791), .A2(keyinput67), .B1(keyinput99), .B2(n6790), 
        .ZN(n6789) );
  OAI221_X1 U7761 ( .B1(n6791), .B2(keyinput67), .C1(n6790), .C2(keyinput99), 
        .A(n6789), .ZN(n6796) );
  AOI22_X1 U7762 ( .A1(n6794), .A2(keyinput45), .B1(n6793), .B2(keyinput53), 
        .ZN(n6792) );
  OAI221_X1 U7763 ( .B1(n6794), .B2(keyinput45), .C1(n6793), .C2(keyinput53), 
        .A(n6792), .ZN(n6795) );
  NOR4_X1 U7764 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n6814)
         );
  AOI22_X1 U7765 ( .A1(n5022), .A2(keyinput116), .B1(n6800), .B2(keyinput35), 
        .ZN(n6799) );
  OAI221_X1 U7766 ( .B1(n5022), .B2(keyinput116), .C1(n6800), .C2(keyinput35), 
        .A(n6799), .ZN(n6812) );
  AOI22_X1 U7767 ( .A1(n6803), .A2(keyinput44), .B1(n6802), .B2(keyinput32), 
        .ZN(n6801) );
  OAI221_X1 U7768 ( .B1(n6803), .B2(keyinput44), .C1(n6802), .C2(keyinput32), 
        .A(n6801), .ZN(n6811) );
  AOI22_X1 U7769 ( .A1(n6805), .A2(keyinput57), .B1(n4905), .B2(keyinput84), 
        .ZN(n6804) );
  OAI221_X1 U7770 ( .B1(n6805), .B2(keyinput57), .C1(n4905), .C2(keyinput84), 
        .A(n6804), .ZN(n6810) );
  AOI22_X1 U7771 ( .A1(n6808), .A2(keyinput5), .B1(keyinput50), .B2(n6807), 
        .ZN(n6806) );
  OAI221_X1 U7772 ( .B1(n6808), .B2(keyinput5), .C1(n6807), .C2(keyinput50), 
        .A(n6806), .ZN(n6809) );
  NOR4_X1 U7773 ( .A1(n6812), .A2(n6811), .A3(n6810), .A4(n6809), .ZN(n6813)
         );
  NAND4_X1 U7774 ( .A1(n6816), .A2(n6815), .A3(n6814), .A4(n6813), .ZN(n7011)
         );
  AOI22_X1 U7775 ( .A1(n6819), .A2(keyinput31), .B1(n6818), .B2(keyinput1), 
        .ZN(n6817) );
  OAI221_X1 U7776 ( .B1(n6819), .B2(keyinput31), .C1(n6818), .C2(keyinput1), 
        .A(n6817), .ZN(n6832) );
  AOI22_X1 U7777 ( .A1(n6822), .A2(keyinput100), .B1(keyinput61), .B2(n6821), 
        .ZN(n6820) );
  OAI221_X1 U7778 ( .B1(n6822), .B2(keyinput100), .C1(n6821), .C2(keyinput61), 
        .A(n6820), .ZN(n6831) );
  INV_X1 U7779 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6824) );
  AOI22_X1 U7780 ( .A1(n6825), .A2(keyinput125), .B1(n6824), .B2(keyinput19), 
        .ZN(n6823) );
  OAI221_X1 U7781 ( .B1(n6825), .B2(keyinput125), .C1(n6824), .C2(keyinput19), 
        .A(n6823), .ZN(n6830) );
  AOI22_X1 U7782 ( .A1(n6828), .A2(keyinput12), .B1(n6827), .B2(keyinput59), 
        .ZN(n6826) );
  OAI221_X1 U7783 ( .B1(n6828), .B2(keyinput12), .C1(n6827), .C2(keyinput59), 
        .A(n6826), .ZN(n6829) );
  NOR4_X1 U7784 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n6881)
         );
  INV_X1 U7785 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6834) );
  AOI22_X1 U7786 ( .A1(n6835), .A2(keyinput123), .B1(keyinput10), .B2(n6834), 
        .ZN(n6833) );
  OAI221_X1 U7787 ( .B1(n6835), .B2(keyinput123), .C1(n6834), .C2(keyinput10), 
        .A(n6833), .ZN(n6848) );
  AOI22_X1 U7788 ( .A1(n6838), .A2(keyinput105), .B1(keyinput110), .B2(n6837), 
        .ZN(n6836) );
  OAI221_X1 U7789 ( .B1(n6838), .B2(keyinput105), .C1(n6837), .C2(keyinput110), 
        .A(n6836), .ZN(n6847) );
  AOI22_X1 U7790 ( .A1(n6841), .A2(keyinput111), .B1(n6840), .B2(keyinput108), 
        .ZN(n6839) );
  OAI221_X1 U7791 ( .B1(n6841), .B2(keyinput111), .C1(n6840), .C2(keyinput108), 
        .A(n6839), .ZN(n6846) );
  AOI22_X1 U7792 ( .A1(n6844), .A2(keyinput58), .B1(n6843), .B2(keyinput104), 
        .ZN(n6842) );
  OAI221_X1 U7793 ( .B1(n6844), .B2(keyinput58), .C1(n6843), .C2(keyinput104), 
        .A(n6842), .ZN(n6845) );
  NOR4_X1 U7794 ( .A1(n6848), .A2(n6847), .A3(n6846), .A4(n6845), .ZN(n6880)
         );
  INV_X1 U7795 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6850) );
  AOI22_X1 U7796 ( .A1(n4563), .A2(keyinput26), .B1(n6850), .B2(keyinput66), 
        .ZN(n6849) );
  OAI221_X1 U7797 ( .B1(n4563), .B2(keyinput26), .C1(n6850), .C2(keyinput66), 
        .A(n6849), .ZN(n6862) );
  INV_X1 U7798 ( .A(ADDRESS_REG_16__SCAN_IN), .ZN(n6852) );
  AOI22_X1 U7799 ( .A1(n6853), .A2(keyinput86), .B1(keyinput107), .B2(n6852), 
        .ZN(n6851) );
  OAI221_X1 U7800 ( .B1(n6853), .B2(keyinput86), .C1(n6852), .C2(keyinput107), 
        .A(n6851), .ZN(n6861) );
  INV_X1 U7801 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6856) );
  AOI22_X1 U7802 ( .A1(n6856), .A2(keyinput36), .B1(keyinput16), .B2(n6855), 
        .ZN(n6854) );
  OAI221_X1 U7803 ( .B1(n6856), .B2(keyinput36), .C1(n6855), .C2(keyinput16), 
        .A(n6854), .ZN(n6860) );
  AOI22_X1 U7804 ( .A1(n4792), .A2(keyinput115), .B1(keyinput15), .B2(n6858), 
        .ZN(n6857) );
  OAI221_X1 U7805 ( .B1(n4792), .B2(keyinput115), .C1(n6858), .C2(keyinput15), 
        .A(n6857), .ZN(n6859) );
  NOR4_X1 U7806 ( .A1(n6862), .A2(n6861), .A3(n6860), .A4(n6859), .ZN(n6879)
         );
  INV_X1 U7807 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6865) );
  INV_X1 U7808 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6864) );
  AOI22_X1 U7809 ( .A1(n6865), .A2(keyinput90), .B1(n6864), .B2(keyinput54), 
        .ZN(n6863) );
  OAI221_X1 U7810 ( .B1(n6865), .B2(keyinput90), .C1(n6864), .C2(keyinput54), 
        .A(n6863), .ZN(n6869) );
  XNOR2_X1 U7811 ( .A(n3183), .B(keyinput117), .ZN(n6868) );
  XNOR2_X1 U7812 ( .A(n6866), .B(keyinput81), .ZN(n6867) );
  OR3_X1 U7813 ( .A1(n6869), .A2(n6868), .A3(n6867), .ZN(n6877) );
  AOI22_X1 U7814 ( .A1(n4898), .A2(keyinput93), .B1(keyinput43), .B2(n6871), 
        .ZN(n6870) );
  OAI221_X1 U7815 ( .B1(n4898), .B2(keyinput93), .C1(n6871), .C2(keyinput43), 
        .A(n6870), .ZN(n6876) );
  INV_X1 U7816 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6874) );
  AOI22_X1 U7817 ( .A1(n6874), .A2(keyinput9), .B1(keyinput118), .B2(n6873), 
        .ZN(n6872) );
  OAI221_X1 U7818 ( .B1(n6874), .B2(keyinput9), .C1(n6873), .C2(keyinput118), 
        .A(n6872), .ZN(n6875) );
  NOR3_X1 U7819 ( .A1(n6877), .A2(n6876), .A3(n6875), .ZN(n6878) );
  NAND4_X1 U7820 ( .A1(n6881), .A2(n6880), .A3(n6879), .A4(n6878), .ZN(n7010)
         );
  AOI22_X1 U7821 ( .A1(n6883), .A2(keyinput52), .B1(n5015), .B2(keyinput2), 
        .ZN(n6882) );
  OAI221_X1 U7822 ( .B1(n6883), .B2(keyinput52), .C1(n5015), .C2(keyinput2), 
        .A(n6882), .ZN(n6895) );
  AOI22_X1 U7823 ( .A1(n6885), .A2(keyinput17), .B1(keyinput121), .B2(n4724), 
        .ZN(n6884) );
  OAI221_X1 U7824 ( .B1(n6885), .B2(keyinput17), .C1(n4724), .C2(keyinput121), 
        .A(n6884), .ZN(n6894) );
  AOI22_X1 U7825 ( .A1(n6888), .A2(keyinput41), .B1(keyinput3), .B2(n6887), 
        .ZN(n6886) );
  OAI221_X1 U7826 ( .B1(n6888), .B2(keyinput41), .C1(n6887), .C2(keyinput3), 
        .A(n6886), .ZN(n6893) );
  INV_X1 U7827 ( .A(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U7828 ( .A1(n6891), .A2(keyinput49), .B1(keyinput46), .B2(n6890), 
        .ZN(n6889) );
  OAI221_X1 U7829 ( .B1(n6891), .B2(keyinput49), .C1(n6890), .C2(keyinput46), 
        .A(n6889), .ZN(n6892) );
  NOR4_X1 U7830 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n6941)
         );
  AOI22_X1 U7831 ( .A1(n6898), .A2(keyinput13), .B1(keyinput47), .B2(n6897), 
        .ZN(n6896) );
  OAI221_X1 U7832 ( .B1(n6898), .B2(keyinput13), .C1(n6897), .C2(keyinput47), 
        .A(n6896), .ZN(n6908) );
  AOI22_X1 U7833 ( .A1(n6900), .A2(keyinput39), .B1(keyinput95), .B2(n4565), 
        .ZN(n6899) );
  OAI221_X1 U7834 ( .B1(n6900), .B2(keyinput39), .C1(n4565), .C2(keyinput95), 
        .A(n6899), .ZN(n6907) );
  AOI22_X1 U7835 ( .A1(n6902), .A2(keyinput82), .B1(keyinput106), .B2(n4555), 
        .ZN(n6901) );
  OAI221_X1 U7836 ( .B1(n6902), .B2(keyinput82), .C1(n4555), .C2(keyinput106), 
        .A(n6901), .ZN(n6906) );
  AOI22_X1 U7837 ( .A1(n4302), .A2(keyinput91), .B1(keyinput88), .B2(n6904), 
        .ZN(n6903) );
  OAI221_X1 U7838 ( .B1(n4302), .B2(keyinput91), .C1(n6904), .C2(keyinput88), 
        .A(n6903), .ZN(n6905) );
  NOR4_X1 U7839 ( .A1(n6908), .A2(n6907), .A3(n6906), .A4(n6905), .ZN(n6940)
         );
  INV_X1 U7840 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6910) );
  AOI22_X1 U7841 ( .A1(n6911), .A2(keyinput114), .B1(keyinput28), .B2(n6910), 
        .ZN(n6909) );
  OAI221_X1 U7842 ( .B1(n6911), .B2(keyinput114), .C1(n6910), .C2(keyinput28), 
        .A(n6909), .ZN(n6923) );
  INV_X1 U7843 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6913) );
  AOI22_X1 U7844 ( .A1(n6914), .A2(keyinput29), .B1(keyinput51), .B2(n6913), 
        .ZN(n6912) );
  OAI221_X1 U7845 ( .B1(n6914), .B2(keyinput29), .C1(n6913), .C2(keyinput51), 
        .A(n6912), .ZN(n6922) );
  INV_X1 U7846 ( .A(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6916) );
  AOI22_X1 U7847 ( .A1(n4561), .A2(keyinput113), .B1(n6916), .B2(keyinput103), 
        .ZN(n6915) );
  OAI221_X1 U7848 ( .B1(n4561), .B2(keyinput113), .C1(n6916), .C2(keyinput103), 
        .A(n6915), .ZN(n6921) );
  AOI22_X1 U7849 ( .A1(n6919), .A2(keyinput4), .B1(n6918), .B2(keyinput94), 
        .ZN(n6917) );
  OAI221_X1 U7850 ( .B1(n6919), .B2(keyinput4), .C1(n6918), .C2(keyinput94), 
        .A(n6917), .ZN(n6920) );
  NOR4_X1 U7851 ( .A1(n6923), .A2(n6922), .A3(n6921), .A4(n6920), .ZN(n6939)
         );
  AOI22_X1 U7852 ( .A1(n6925), .A2(keyinput11), .B1(n4234), .B2(keyinput73), 
        .ZN(n6924) );
  OAI221_X1 U7853 ( .B1(n6925), .B2(keyinput11), .C1(n4234), .C2(keyinput73), 
        .A(n6924), .ZN(n6937) );
  AOI22_X1 U7854 ( .A1(n6928), .A2(keyinput25), .B1(n6927), .B2(keyinput22), 
        .ZN(n6926) );
  OAI221_X1 U7855 ( .B1(n6928), .B2(keyinput25), .C1(n6927), .C2(keyinput22), 
        .A(n6926), .ZN(n6936) );
  INV_X1 U7856 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U7857 ( .A1(n6931), .A2(keyinput8), .B1(keyinput18), .B2(n6930), 
        .ZN(n6929) );
  OAI221_X1 U7858 ( .B1(n6931), .B2(keyinput8), .C1(n6930), .C2(keyinput18), 
        .A(n6929), .ZN(n6935) );
  AOI22_X1 U7859 ( .A1(n4495), .A2(keyinput102), .B1(keyinput122), .B2(n6933), 
        .ZN(n6932) );
  OAI221_X1 U7860 ( .B1(n4495), .B2(keyinput102), .C1(n6933), .C2(keyinput122), 
        .A(n6932), .ZN(n6934) );
  NOR4_X1 U7861 ( .A1(n6937), .A2(n6936), .A3(n6935), .A4(n6934), .ZN(n6938)
         );
  NAND4_X1 U7862 ( .A1(n6941), .A2(n6940), .A3(n6939), .A4(n6938), .ZN(n7009)
         );
  INV_X1 U7863 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6943) );
  AOI22_X1 U7864 ( .A1(n6943), .A2(keyinput21), .B1(n4949), .B2(keyinput70), 
        .ZN(n6942) );
  OAI221_X1 U7865 ( .B1(n6943), .B2(keyinput21), .C1(n4949), .C2(keyinput70), 
        .A(n6942), .ZN(n6956) );
  AOI22_X1 U7866 ( .A1(n6946), .A2(keyinput126), .B1(keyinput119), .B2(n6945), 
        .ZN(n6944) );
  OAI221_X1 U7867 ( .B1(n6946), .B2(keyinput126), .C1(n6945), .C2(keyinput119), 
        .A(n6944), .ZN(n6955) );
  AOI22_X1 U7868 ( .A1(n6949), .A2(keyinput92), .B1(keyinput75), .B2(n6948), 
        .ZN(n6947) );
  OAI221_X1 U7869 ( .B1(n6949), .B2(keyinput92), .C1(n6948), .C2(keyinput75), 
        .A(n6947), .ZN(n6954) );
  INV_X1 U7870 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6952) );
  AOI22_X1 U7871 ( .A1(n6952), .A2(keyinput23), .B1(n6951), .B2(keyinput30), 
        .ZN(n6950) );
  OAI221_X1 U7872 ( .B1(n6952), .B2(keyinput23), .C1(n6951), .C2(keyinput30), 
        .A(n6950), .ZN(n6953) );
  NOR4_X1 U7873 ( .A1(n6956), .A2(n6955), .A3(n6954), .A4(n6953), .ZN(n7007)
         );
  AOI22_X1 U7874 ( .A1(n6959), .A2(keyinput48), .B1(keyinput85), .B2(n6958), 
        .ZN(n6957) );
  OAI221_X1 U7875 ( .B1(n6959), .B2(keyinput48), .C1(n6958), .C2(keyinput85), 
        .A(n6957), .ZN(n6972) );
  INV_X1 U7876 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6962) );
  INV_X1 U7877 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6961) );
  AOI22_X1 U7878 ( .A1(n6962), .A2(keyinput60), .B1(keyinput64), .B2(n6961), 
        .ZN(n6960) );
  OAI221_X1 U7879 ( .B1(n6962), .B2(keyinput60), .C1(n6961), .C2(keyinput64), 
        .A(n6960), .ZN(n6971) );
  INV_X1 U7880 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6965) );
  INV_X1 U7881 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6964) );
  AOI22_X1 U7882 ( .A1(n6965), .A2(keyinput96), .B1(keyinput80), .B2(n6964), 
        .ZN(n6963) );
  OAI221_X1 U7883 ( .B1(n6965), .B2(keyinput96), .C1(n6964), .C2(keyinput80), 
        .A(n6963), .ZN(n6970) );
  AOI22_X1 U7884 ( .A1(n6968), .A2(keyinput6), .B1(n6967), .B2(keyinput109), 
        .ZN(n6966) );
  OAI221_X1 U7885 ( .B1(n6968), .B2(keyinput6), .C1(n6967), .C2(keyinput109), 
        .A(n6966), .ZN(n6969) );
  NOR4_X1 U7886 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n7006)
         );
  AOI22_X1 U7887 ( .A1(n6975), .A2(keyinput62), .B1(keyinput71), .B2(n6974), 
        .ZN(n6973) );
  OAI221_X1 U7888 ( .B1(n6975), .B2(keyinput62), .C1(n6974), .C2(keyinput71), 
        .A(n6973), .ZN(n6987) );
  AOI22_X1 U7889 ( .A1(n6977), .A2(keyinput76), .B1(n4961), .B2(keyinput33), 
        .ZN(n6976) );
  OAI221_X1 U7890 ( .B1(n6977), .B2(keyinput76), .C1(n4961), .C2(keyinput33), 
        .A(n6976), .ZN(n6986) );
  INV_X1 U7891 ( .A(DATAI_31_), .ZN(n6980) );
  AOI22_X1 U7892 ( .A1(n6980), .A2(keyinput79), .B1(n6979), .B2(keyinput7), 
        .ZN(n6978) );
  OAI221_X1 U7893 ( .B1(n6980), .B2(keyinput79), .C1(n6979), .C2(keyinput7), 
        .A(n6978), .ZN(n6985) );
  INV_X1 U7894 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U7895 ( .A1(n6983), .A2(keyinput112), .B1(keyinput40), .B2(n6982), 
        .ZN(n6981) );
  OAI221_X1 U7896 ( .B1(n6983), .B2(keyinput112), .C1(n6982), .C2(keyinput40), 
        .A(n6981), .ZN(n6984) );
  NOR4_X1 U7897 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n7005)
         );
  INV_X1 U7898 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6990) );
  INV_X1 U7899 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6989) );
  AOI22_X1 U7900 ( .A1(n6990), .A2(keyinput34), .B1(keyinput120), .B2(n6989), 
        .ZN(n6988) );
  OAI221_X1 U7901 ( .B1(n6990), .B2(keyinput34), .C1(n6989), .C2(keyinput120), 
        .A(n6988), .ZN(n7003) );
  INV_X1 U7902 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6992) );
  AOI22_X1 U7903 ( .A1(n6993), .A2(keyinput97), .B1(n6992), .B2(keyinput14), 
        .ZN(n6991) );
  OAI221_X1 U7904 ( .B1(n6993), .B2(keyinput97), .C1(n6992), .C2(keyinput14), 
        .A(n6991), .ZN(n7002) );
  INV_X1 U7905 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6995) );
  AOI22_X1 U7906 ( .A1(n6996), .A2(keyinput89), .B1(n6995), .B2(keyinput27), 
        .ZN(n6994) );
  OAI221_X1 U7907 ( .B1(n6996), .B2(keyinput89), .C1(n6995), .C2(keyinput27), 
        .A(n6994), .ZN(n7001) );
  INV_X1 U7908 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n6999) );
  AOI22_X1 U7909 ( .A1(n6999), .A2(keyinput98), .B1(keyinput77), .B2(n6998), 
        .ZN(n6997) );
  OAI221_X1 U7910 ( .B1(n6999), .B2(keyinput98), .C1(n6998), .C2(keyinput77), 
        .A(n6997), .ZN(n7000) );
  NOR4_X1 U7911 ( .A1(n7003), .A2(n7002), .A3(n7001), .A4(n7000), .ZN(n7004)
         );
  NAND4_X1 U7912 ( .A1(n7007), .A2(n7006), .A3(n7005), .A4(n7004), .ZN(n7008)
         );
  NOR4_X1 U7913 ( .A1(n7011), .A2(n7010), .A3(n7009), .A4(n7008), .ZN(n7012)
         );
  XNOR2_X1 U7914 ( .A(n7013), .B(n7012), .ZN(n7019) );
  OAI222_X1 U7915 ( .A1(n5456), .A2(n7017), .B1(n7016), .B2(n4298), .C1(n7015), 
        .C2(n7014), .ZN(n7018) );
  XNOR2_X1 U7916 ( .A(n7019), .B(n7018), .ZN(U2841) );
  AND2_X2 U4225 ( .A1(n4531), .A2(n3191), .ZN(n3299) );
  AND2_X1 U3709 ( .A1(n4373), .A2(n5448), .ZN(n5440) );
  OAI211_X1 U3706 ( .C1(n4226), .C2(n3139), .A(n3137), .B(n3136), .ZN(n4465)
         );
  CLKBUF_X1 U3579 ( .A(n3442), .Z(n3485) );
  CLKBUF_X1 U3581 ( .A(n3342), .Z(n4543) );
  CLKBUF_X1 U3685 ( .A(n3321), .Z(n4456) );
  CLKBUF_X1 U3708 ( .A(n3345), .Z(n4496) );
  CLKBUF_X1 U4007 ( .A(n3341), .Z(n4322) );
  NAND2_X1 U4132 ( .A1(n5440), .A2(n5443), .ZN(n5442) );
endmodule

