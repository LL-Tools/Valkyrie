

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, 
        REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, 
        REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, 
        REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, 
        REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, 
        REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, 
        REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, 
        REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, 
        REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, 
        IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, 
        IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, 
        IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, 
        IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, 
        IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, 
        IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, 
        IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, 
        IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, 
        IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, 
        IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, 
        D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, 
        D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, 
        D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, 
        D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, 
        D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, 
        D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, 
        D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, 
        D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, 
        D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, 
        D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, 
        REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, 
        REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, 
        REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, 
        REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, 
        REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, 
        REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, 
        REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, 
        REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, 
        REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, 
        REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, 
        REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, 
        REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, 
        REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, 
        REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, 
        REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, 
        REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, 
        REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, 
        REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, 
        REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, 
        REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, 
        REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, 
        REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, 
        REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, 
        REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, 
        REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, 
        REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, 
        REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, 
        REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, 
        REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, 
        REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, 
        REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, 
        REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, 
        ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, 
        ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, 
        ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, 
        ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, 
        ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, 
        ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, 
        ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, 
        DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, 
        DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, 
        DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, 
        DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, 
        DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, 
        DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, 
        DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, 
        DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, 
        DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, 
        DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, 
        DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, 
        REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, 
        REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, 
        U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343, U3342, 
        U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333, U3332, 
        U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323, U3322, 
        U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315, U3314, 
        U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305, U3304, 
        U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295, U3294, 
        U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477, U3479, 
        U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497, U3499, 
        U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511, U3512, 
        U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521, U3522, 
        U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531, U3532, 
        U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541, U3542, 
        U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289, U3288, 
        U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279, U3278, 
        U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269, U3268, 
        U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260, U3259, 
        U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250, U3249, 
        U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240, U3550, 
        U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559, U3560, 
        U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569, U3570, 
        U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579, U3580, 
        U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232, U3231, 
        U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222, U3221, 
        U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212, U3211, 
        U3210, U3149, U3148, U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, DATAI_31_, DATAI_30_, DATAI_29_,
         DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
         DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
         DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
         DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
         DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN,
         REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
         REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
         REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
         REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
         REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
         REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
         REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
         REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
         IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
         IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
         IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
         IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
         IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
         IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
         IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
         IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
         IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
         IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
         D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN,
         D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, D_REG_5__SCAN_IN,
         D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN,
         D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN,
         D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN,
         D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN,
         D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN,
         D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN,
         D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN,
         D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN,
         D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN,
         REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN,
         REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN,
         REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN,
         REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN,
         REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN,
         REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN,
         REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN,
         REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN,
         REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN,
         REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN,
         REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN,
         REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN,
         REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN,
         REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN,
         REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN,
         REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN,
         REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN,
         REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN,
         REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN,
         REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN,
         REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN,
         REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN,
         REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN,
         REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN,
         REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN,
         REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN,
         REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN,
         REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN,
         REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN,
         REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN,
         REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN,
         REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN,
         ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN,
         ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN,
         ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN,
         ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN,
         ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN,
         ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN,
         ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN,
         REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN,
         REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062;

  INV_X2 U2295 ( .A(IR_REG_31__SCAN_IN), .ZN(n3190) );
  INV_X1 U2296 ( .A(n3596), .ZN(n3566) );
  OAI211_X1 U2297 ( .C1(n4238), .C2(n4232), .A(n4233), .B(n4231), .ZN(n4230)
         );
  OAI21_X1 U2298 ( .B1(n3326), .B2(n2525), .A(n2521), .ZN(n3719) );
  NOR3_X1 U2299 ( .A1(n4335), .A2(n2326), .A3(n5049), .ZN(n2328) );
  NOR2_X2 U2300 ( .A1(n3153), .A2(IR_REG_9__SCAN_IN), .ZN(n3189) );
  OR2_X2 U2301 ( .A1(n2827), .A2(n2286), .ZN(n2479) );
  NOR2_X1 U2302 ( .A1(n2671), .A2(n2672), .ZN(n3961) );
  INV_X2 U2303 ( .A(n5058), .ZN(n2260) );
  INV_X1 U2304 ( .A(n2713), .ZN(n2719) );
  NAND4_X1 U2305 ( .A1(n2778), .A2(n2777), .A3(n2776), .A4(n2775), .ZN(n3931)
         );
  AOI21_X1 U2306 ( .B1(n2650), .B2(REG1_REG_3__SCAN_IN), .A(n2477), .ZN(n2654)
         );
  NOR2_X1 U2307 ( .A1(n2276), .A2(n2330), .ZN(n2329) );
  NAND2_X1 U2308 ( .A1(n2456), .A2(n4068), .ZN(n4108) );
  OAI21_X1 U2309 ( .B1(n2519), .B2(n2517), .A(n2516), .ZN(n3374) );
  OAI21_X1 U2310 ( .B1(n4253), .B2(n2470), .A(n2469), .ZN(n2468) );
  NAND2_X1 U2311 ( .A1(n2472), .A2(n2471), .ZN(n4253) );
  NOR3_X2 U2312 ( .A1(n4172), .A2(n2324), .A3(n4156), .ZN(n4117) );
  NAND2_X1 U2313 ( .A1(n4189), .A2(n4173), .ZN(n4172) );
  NAND2_X1 U2314 ( .A1(n3057), .A2(n3056), .ZN(n3082) );
  AND2_X2 U2315 ( .A1(n2927), .A2(n4950), .ZN(n5058) );
  NOR2_X2 U2316 ( .A1(n2630), .A2(n2629), .ZN(n4869) );
  NAND2_X1 U2317 ( .A1(n2719), .A2(n4876), .ZN(n5007) );
  INV_X1 U2318 ( .A(n2928), .ZN(n2757) );
  NAND2_X1 U2319 ( .A1(n2805), .A2(n2804), .ZN(n2843) );
  NAND2_X2 U2320 ( .A1(n2719), .A2(n3797), .ZN(n2928) );
  INV_X1 U2321 ( .A(n2748), .ZN(n4034) );
  NAND4_X1 U2322 ( .A1(n2852), .A2(n2851), .A3(n2850), .A4(n2849), .ZN(n3930)
         );
  CLKBUF_X1 U2323 ( .A(n2713), .Z(n2262) );
  INV_X1 U2324 ( .A(n3795), .ZN(n2314) );
  OAI21_X1 U2325 ( .B1(n2596), .B2(n2378), .A(IR_REG_31__SCAN_IN), .ZN(n2380)
         );
  XNOR2_X1 U2326 ( .A(n2567), .B(IR_REG_24__SCAN_IN), .ZN(n2726) );
  NAND2_X1 U2327 ( .A1(n2584), .A2(n2297), .ZN(n2596) );
  AND2_X2 U2328 ( .A1(n2706), .A2(n2708), .ZN(n3774) );
  INV_X1 U2329 ( .A(n2708), .ZN(n2707) );
  NAND2_X1 U2330 ( .A1(n2602), .A2(n3353), .ZN(n2708) );
  XNOR2_X1 U2331 ( .A(n2705), .B(n3350), .ZN(n2706) );
  MUX2_X1 U2332 ( .A(IR_REG_31__SCAN_IN), .B(n2600), .S(IR_REG_29__SCAN_IN), 
        .Z(n2602) );
  OR2_X1 U2333 ( .A1(n2704), .A2(n3190), .ZN(n2705) );
  NAND2_X1 U2334 ( .A1(n3359), .A2(IR_REG_31__SCAN_IN), .ZN(n3368) );
  AND2_X1 U2335 ( .A1(n2475), .A2(n2543), .ZN(n2474) );
  NOR2_X1 U2336 ( .A1(n3357), .A2(IR_REG_26__SCAN_IN), .ZN(n2318) );
  AND2_X1 U2337 ( .A1(n2277), .A2(n2562), .ZN(n2543) );
  NAND2_X1 U2338 ( .A1(n2512), .A2(n2513), .ZN(n4766) );
  NOR2_X1 U2339 ( .A1(n2548), .A2(n2569), .ZN(n2547) );
  NAND2_X1 U2340 ( .A1(n2597), .A2(n2379), .ZN(n2378) );
  AND3_X1 U2341 ( .A1(n2617), .A2(n4594), .A3(n4721), .ZN(n2560) );
  NOR2_X1 U2342 ( .A1(n2595), .A2(IR_REG_19__SCAN_IN), .ZN(n2379) );
  NOR2_X2 U2343 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2615)
         );
  NOR2_X1 U2344 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2559)
         );
  INV_X1 U2345 ( .A(IR_REG_23__SCAN_IN), .ZN(n2576) );
  INV_X1 U2346 ( .A(IR_REG_15__SCAN_IN), .ZN(n3393) );
  NOR2_X1 U2347 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2558)
         );
  BUF_X4 U2348 ( .A(n3778), .Z(n2261) );
  NAND2_X1 U2349 ( .A1(n2624), .A2(n2623), .ZN(n3778) );
  NAND4_X2 U2350 ( .A1(n2762), .A2(n2761), .A3(n2760), .A4(n2759), .ZN(n2906)
         );
  INV_X4 U2351 ( .A(n3595), .ZN(n3548) );
  INV_X1 U2352 ( .A(IR_REG_13__SCAN_IN), .ZN(n2562) );
  AND2_X1 U2353 ( .A1(n2289), .A2(n2263), .ZN(n2448) );
  INV_X1 U2354 ( .A(n2797), .ZN(n3603) );
  AND2_X1 U2355 ( .A1(n3851), .A2(n4085), .ZN(n2402) );
  INV_X1 U2356 ( .A(n4087), .ZN(n2401) );
  AOI21_X1 U2357 ( .B1(n2525), .B2(n2518), .A(n3635), .ZN(n2516) );
  AND2_X1 U2358 ( .A1(n2438), .A2(n2278), .ZN(n2437) );
  NOR2_X1 U2359 ( .A1(n2442), .A2(n4333), .ZN(n2441) );
  INV_X1 U2360 ( .A(n2444), .ZN(n2442) );
  AOI21_X1 U2361 ( .B1(n2463), .B2(n3081), .A(n2285), .ZN(n2461) );
  AND2_X1 U2362 ( .A1(n2543), .A2(n2476), .ZN(n2473) );
  AND2_X1 U2363 ( .A1(n2547), .A2(n2476), .ZN(n2475) );
  INV_X1 U2364 ( .A(n3647), .ZN(n3517) );
  INV_X1 U2365 ( .A(n2802), .ZN(n3604) );
  NAND2_X1 U2366 ( .A1(n2691), .A2(n2662), .ZN(n2663) );
  NOR2_X1 U2367 ( .A1(n2687), .A2(n2515), .ZN(n2680) );
  AND2_X1 U2368 ( .A1(n4762), .A2(REG2_REG_5__SCAN_IN), .ZN(n2515) );
  OR2_X1 U2369 ( .A1(n4802), .A2(n4803), .ZN(n2514) );
  NOR2_X1 U2370 ( .A1(n3961), .A2(n3962), .ZN(n4813) );
  OAI22_X1 U2371 ( .A1(n4832), .A2(n4830), .B1(n3965), .B2(
        REG1_REG_11__SCAN_IN), .ZN(n3966) );
  AOI21_X1 U2372 ( .B1(n2460), .B2(n2459), .A(n2458), .ZN(n4125) );
  NAND2_X1 U2373 ( .A1(n4065), .A2(n4156), .ZN(n2459) );
  AND2_X1 U2374 ( .A1(n4169), .A2(n4066), .ZN(n2458) );
  INV_X1 U2375 ( .A(n4144), .ZN(n2460) );
  OR2_X1 U2376 ( .A1(n3556), .A2(n3747), .ZN(n3572) );
  OR2_X1 U2377 ( .A1(n4061), .A2(n4213), .ZN(n4062) );
  NAND2_X1 U2378 ( .A1(n2451), .A2(n2552), .ZN(n2450) );
  OR2_X1 U2379 ( .A1(n3509), .A2(n4514), .ZN(n3536) );
  INV_X1 U2380 ( .A(n2468), .ZN(n4238) );
  AND2_X1 U2381 ( .A1(n4279), .A2(n5049), .ZN(n2470) );
  NAND2_X1 U2382 ( .A1(n5031), .A2(n4057), .ZN(n2469) );
  NAND2_X1 U2383 ( .A1(n3796), .A2(n2912), .ZN(n3882) );
  OAI22_X1 U2384 ( .A1(n2740), .A2(D_REG_0__SCAN_IN), .B1(n2737), .B2(n2726), 
        .ZN(n3002) );
  NOR2_X1 U2385 ( .A1(n2573), .A2(n2738), .ZN(n2575) );
  INV_X1 U2386 ( .A(n3466), .ZN(n2541) );
  NOR2_X1 U2387 ( .A1(n3715), .A2(n2522), .ZN(n2518) );
  NAND2_X1 U2388 ( .A1(n2549), .A2(n2589), .ZN(n2548) );
  INV_X1 U2389 ( .A(IR_REG_25__SCAN_IN), .ZN(n2549) );
  NOR2_X1 U2390 ( .A1(n2539), .A2(n3725), .ZN(n2362) );
  INV_X1 U2391 ( .A(n3725), .ZN(n2364) );
  NOR2_X1 U2392 ( .A1(n3190), .A2(n2316), .ZN(n2315) );
  AND2_X1 U2393 ( .A1(n3868), .A2(n4181), .ZN(n4084) );
  NAND2_X1 U2394 ( .A1(n2496), .A2(n2495), .ZN(n2494) );
  NOR2_X1 U2395 ( .A1(n2493), .A2(n2766), .ZN(n2492) );
  INV_X1 U2396 ( .A(n2664), .ZN(n2493) );
  AND2_X1 U2397 ( .A1(n2491), .A2(n2489), .ZN(n3962) );
  NOR2_X1 U2398 ( .A1(n2668), .A2(n2490), .ZN(n2489) );
  INV_X1 U2399 ( .A(n2494), .ZN(n2490) );
  INV_X1 U2400 ( .A(n4818), .ZN(n2344) );
  NOR2_X1 U2401 ( .A1(n2344), .A2(n3106), .ZN(n2341) );
  NAND2_X1 U2402 ( .A1(n2287), .A2(n3782), .ZN(n2395) );
  NAND2_X1 U2403 ( .A1(n2399), .A2(n2400), .ZN(n2398) );
  INV_X1 U2404 ( .A(n2402), .ZN(n2399) );
  INV_X1 U2405 ( .A(n4333), .ZN(n2415) );
  AND2_X1 U2406 ( .A1(n2419), .A2(n4078), .ZN(n2418) );
  INV_X1 U2407 ( .A(n4079), .ZN(n2419) );
  AND2_X1 U2408 ( .A1(n2440), .A2(n2278), .ZN(n2435) );
  INV_X1 U2409 ( .A(n3844), .ZN(n4078) );
  NAND2_X1 U2410 ( .A1(n4075), .A2(n4074), .ZN(n2383) );
  AND2_X1 U2411 ( .A1(n4386), .A2(n3755), .ZN(n3833) );
  AOI21_X1 U2412 ( .B1(n3820), .B2(n3815), .A(n2389), .ZN(n2388) );
  INV_X1 U2413 ( .A(n3817), .ZN(n2389) );
  INV_X1 U2414 ( .A(n3815), .ZN(n2390) );
  OR2_X1 U2415 ( .A1(n3207), .A2(n3206), .ZN(n3252) );
  AND2_X1 U2416 ( .A1(n3083), .A2(n2464), .ZN(n2463) );
  INV_X1 U2417 ( .A(n3824), .ZN(n2405) );
  NOR2_X1 U2418 ( .A1(n3058), .A2(n2412), .ZN(n2411) );
  NAND2_X1 U2419 ( .A1(n2403), .A2(n3824), .ZN(n2408) );
  NAND2_X1 U2420 ( .A1(n2411), .A2(n2972), .ZN(n2403) );
  INV_X1 U2421 ( .A(n2843), .ZN(n2963) );
  NAND2_X1 U2422 ( .A1(n2920), .A2(n2995), .ZN(n3799) );
  NAND2_X1 U2423 ( .A1(n3799), .A2(n3802), .ZN(n2914) );
  AND2_X1 U2424 ( .A1(n2547), .A2(n2599), .ZN(n2545) );
  NOR2_X1 U2425 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2599)
         );
  NOR2_X1 U2426 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2565)
         );
  NAND2_X1 U2427 ( .A1(n3393), .A2(n2563), .ZN(n3409) );
  INV_X1 U2428 ( .A(IR_REG_16__SCAN_IN), .ZN(n2563) );
  INV_X1 U2429 ( .A(IR_REG_5__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U2430 ( .A1(n2376), .A2(n2306), .ZN(n2375) );
  INV_X1 U2431 ( .A(n3121), .ZN(n2376) );
  INV_X1 U2432 ( .A(n3745), .ZN(n2532) );
  NAND2_X1 U2433 ( .A1(n3719), .A2(n3715), .ZN(n3377) );
  AND2_X1 U2434 ( .A1(n2717), .A2(n2716), .ZN(n2782) );
  INV_X1 U2435 ( .A(n3675), .ZN(n3677) );
  NAND2_X1 U2436 ( .A1(n3675), .A2(n3674), .ZN(n3706) );
  INV_X1 U2437 ( .A(n5050), .ZN(n3748) );
  OR2_X1 U2438 ( .A1(n3237), .A2(n4699), .ZN(n3385) );
  NAND2_X1 U2439 ( .A1(n3939), .A2(n3938), .ZN(n3937) );
  AOI22_X1 U2440 ( .A1(n2683), .A2(REG2_REG_7__SCAN_IN), .B1(n2682), .B2(n4761), .ZN(n3947) );
  NOR2_X1 U2441 ( .A1(REG2_REG_7__SCAN_IN), .A2(n2357), .ZN(n2356) );
  INV_X1 U2442 ( .A(n2275), .ZN(n2357) );
  NOR3_X1 U2443 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .A3(
        IR_REG_11__SCAN_IN), .ZN(n2561) );
  INV_X1 U2444 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U2445 ( .A1(n2310), .A2(n3969), .ZN(n3979) );
  NAND2_X1 U2446 ( .A1(n4853), .A2(n4851), .ZN(n2310) );
  OR2_X1 U2447 ( .A1(n4856), .A2(n2333), .ZN(n2331) );
  OR2_X1 U2448 ( .A1(n4855), .A2(n4759), .ZN(n2333) );
  OR2_X1 U2449 ( .A1(n4759), .A2(n2338), .ZN(n2332) );
  NOR2_X1 U2450 ( .A1(n2337), .A2(n3957), .ZN(n2336) );
  OR2_X1 U2451 ( .A1(n4856), .A2(n4855), .ZN(n2339) );
  INV_X1 U2452 ( .A(n2338), .ZN(n2337) );
  NAND2_X1 U2453 ( .A1(n2505), .A2(n2504), .ZN(n4002) );
  INV_X1 U2454 ( .A(n3976), .ZN(n2504) );
  INV_X1 U2455 ( .A(n3984), .ZN(n2482) );
  NOR2_X1 U2456 ( .A1(n2487), .A2(n4003), .ZN(n2484) );
  OR2_X1 U2457 ( .A1(n4871), .A2(REG1_REG_16__SCAN_IN), .ZN(n2309) );
  AND2_X1 U2458 ( .A1(n4002), .A2(n4001), .ZN(n4004) );
  NAND2_X1 U2459 ( .A1(n2349), .A2(n2355), .ZN(n2346) );
  NAND2_X1 U2460 ( .A1(n4117), .A2(n4101), .ZN(n4415) );
  OAI21_X1 U2461 ( .B1(n4164), .B2(n2396), .A(n2395), .ZN(n4109) );
  OR2_X1 U2462 ( .A1(n3628), .A2(n3603), .ZN(n3579) );
  NAND2_X1 U2463 ( .A1(n2447), .A2(n2446), .ZN(n4161) );
  AOI21_X1 U2464 ( .B1(n2448), .B2(n2452), .A(n2284), .ZN(n2446) );
  NAND2_X1 U2465 ( .A1(n3522), .A2(REG3_REG_24__SCAN_IN), .ZN(n3538) );
  INV_X1 U2466 ( .A(n3536), .ZN(n3522) );
  INV_X1 U2467 ( .A(n2552), .ZN(n2452) );
  NAND2_X1 U2468 ( .A1(n4242), .A2(n4058), .ZN(n4059) );
  OR2_X1 U2469 ( .A1(n4259), .A2(n4284), .ZN(n2471) );
  NAND2_X1 U2470 ( .A1(n4282), .A2(n2295), .ZN(n2472) );
  INV_X1 U2471 ( .A(n2441), .ZN(n2440) );
  AOI21_X1 U2472 ( .B1(n2441), .B2(n2439), .A(n2294), .ZN(n2438) );
  INV_X1 U2473 ( .A(n4054), .ZN(n2439) );
  AOI21_X1 U2474 ( .B1(n4054), .B2(n4359), .A(n2445), .ZN(n2444) );
  INV_X1 U2475 ( .A(n4056), .ZN(n2445) );
  AND2_X1 U2476 ( .A1(n4078), .A2(n3869), .ZN(n4333) );
  NAND2_X1 U2477 ( .A1(n3226), .A2(n3831), .ZN(n4388) );
  OAI21_X1 U2478 ( .B1(n4938), .B2(n2426), .A(n2423), .ZN(n3187) );
  AOI21_X1 U2479 ( .B1(n2427), .B2(n2425), .A(n2424), .ZN(n2423) );
  INV_X1 U2480 ( .A(n2427), .ZN(n2426) );
  INV_X1 U2481 ( .A(n3826), .ZN(n2424) );
  OAI21_X1 U2482 ( .B1(n4938), .B2(n3092), .A(n3823), .ZN(n3156) );
  NAND2_X1 U2483 ( .A1(n2466), .A2(n2465), .ZN(n2464) );
  AND2_X1 U2484 ( .A1(n3811), .A2(n3823), .ZN(n4937) );
  NAND2_X1 U2485 ( .A1(n2715), .A2(n2606), .ZN(n2756) );
  INV_X1 U2486 ( .A(n3931), .ZN(n2920) );
  INV_X1 U2487 ( .A(n2914), .ZN(n3884) );
  NAND2_X1 U2488 ( .A1(n3882), .A2(n2946), .ZN(n2945) );
  INV_X1 U2489 ( .A(n4880), .ZN(n4944) );
  AND2_X1 U2490 ( .A1(n2720), .A2(n3908), .ZN(n4876) );
  AOI21_X1 U2491 ( .B1(n4097), .B2(n4878), .A(n4096), .ZN(n4422) );
  OR2_X1 U2492 ( .A1(n4885), .A2(n3920), .ZN(n4983) );
  NAND2_X1 U2493 ( .A1(n2605), .A2(n2737), .ZN(n2740) );
  INV_X1 U2494 ( .A(n2597), .ZN(n2377) );
  AND2_X1 U2495 ( .A1(n3234), .A2(n3225), .ZN(n3965) );
  AND2_X1 U2496 ( .A1(n2643), .A2(n2642), .ZN(n2656) );
  AOI21_X1 U2497 ( .B1(n2373), .B2(n3122), .A(n2280), .ZN(n2372) );
  NAND2_X1 U2498 ( .A1(n2313), .A2(n4766), .ZN(n2312) );
  INV_X1 U2499 ( .A(n2261), .ZN(n2313) );
  AND2_X1 U2500 ( .A1(n2858), .A2(n2857), .ZN(n5054) );
  AND2_X1 U2501 ( .A1(n2758), .A2(n2751), .ZN(n5048) );
  NAND2_X1 U2502 ( .A1(n3563), .A2(n3562), .ZN(n4065) );
  NAND2_X1 U2503 ( .A1(n3529), .A2(n3528), .ZN(n4150) );
  OR2_X1 U2504 ( .A1(n3684), .A2(n3603), .ZN(n3529) );
  OAI211_X1 U2505 ( .C1(n4215), .C2(n3603), .A(n3512), .B(n3511), .ZN(n4224)
         );
  NAND2_X1 U2506 ( .A1(n2797), .A2(REG3_REG_1__SCAN_IN), .ZN(n2760) );
  AND2_X1 U2507 ( .A1(n3936), .A2(n2613), .ZN(n2829) );
  NAND2_X1 U2508 ( .A1(n2514), .A2(n2275), .ZN(n2683) );
  NAND2_X1 U2509 ( .A1(n4806), .A2(n2664), .ZN(n2769) );
  NAND2_X1 U2510 ( .A1(n3949), .A2(n3950), .ZN(n4817) );
  NAND2_X1 U2511 ( .A1(n4822), .A2(n3964), .ZN(n4832) );
  XNOR2_X1 U2512 ( .A(n3966), .B(n4980), .ZN(n4842) );
  NOR2_X1 U2513 ( .A1(n4842), .A2(n4843), .ZN(n4841) );
  XNOR2_X1 U2514 ( .A(n4004), .B(n4003), .ZN(n4866) );
  NAND2_X1 U2515 ( .A1(n4866), .A2(n4340), .ZN(n4865) );
  NAND2_X1 U2516 ( .A1(n4415), .A2(n4102), .ZN(n4423) );
  OR2_X1 U2517 ( .A1(n4117), .A2(n4101), .ZN(n4102) );
  INV_X1 U2518 ( .A(n4810), .ZN(n4959) );
  XNOR2_X1 U2519 ( .A(n2609), .B(IR_REG_2__SCAN_IN), .ZN(n4765) );
  NAND2_X1 U2520 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2609) );
  INV_X1 U2521 ( .A(n2615), .ZN(n2360) );
  INV_X1 U2522 ( .A(n2518), .ZN(n2517) );
  NAND2_X1 U2523 ( .A1(n3645), .A2(n3521), .ZN(n3675) );
  OR2_X1 U2524 ( .A1(n5030), .A2(n2541), .ZN(n2540) );
  NAND2_X1 U2525 ( .A1(n4982), .A2(n4402), .ZN(n2338) );
  NAND2_X1 U2526 ( .A1(n3990), .A2(n2486), .ZN(n3992) );
  INV_X1 U2527 ( .A(n3997), .ZN(n2499) );
  NOR2_X1 U2528 ( .A1(n2551), .A2(n2354), .ZN(n2347) );
  OR2_X1 U2529 ( .A1(n4088), .A2(n3853), .ZN(n3900) );
  INV_X1 U2530 ( .A(n4059), .ZN(n2451) );
  INV_X1 U2531 ( .A(n4378), .ZN(n4370) );
  AOI21_X1 U2532 ( .B1(n3092), .B2(n3823), .A(n2428), .ZN(n2427) );
  INV_X1 U2533 ( .A(n3814), .ZN(n2428) );
  NAND2_X1 U2534 ( .A1(n2906), .A2(n2947), .ZN(n3796) );
  AND2_X1 U2535 ( .A1(n3920), .A2(n3797), .ZN(n2917) );
  AOI21_X1 U2536 ( .B1(n2394), .B2(n2396), .A(n2393), .ZN(n2392) );
  INV_X1 U2537 ( .A(n4090), .ZN(n2393) );
  NAND2_X1 U2538 ( .A1(n2397), .A2(n2400), .ZN(n4127) );
  AND2_X1 U2539 ( .A1(n4227), .A2(n4213), .ZN(n4190) );
  NAND2_X1 U2540 ( .A1(n2327), .A2(n4284), .ZN(n2326) );
  NOR2_X1 U2541 ( .A1(n3761), .A2(n4317), .ZN(n2327) );
  INV_X1 U2542 ( .A(n3307), .ZN(n3271) );
  AND2_X1 U2543 ( .A1(n2322), .A2(n3170), .ZN(n2321) );
  AND2_X1 U2544 ( .A1(n4940), .A2(n3151), .ZN(n2322) );
  INV_X1 U2545 ( .A(IR_REG_24__SCAN_IN), .ZN(n2568) );
  INV_X1 U2546 ( .A(IR_REG_19__SCAN_IN), .ZN(n2744) );
  OR2_X1 U2547 ( .A1(n2658), .A2(IR_REG_6__SCAN_IN), .ZN(n2648) );
  NAND2_X1 U2548 ( .A1(n2366), .A2(n2364), .ZN(n2363) );
  AOI21_X1 U2549 ( .B1(n2366), .B2(n2362), .A(n2296), .ZN(n2361) );
  NAND2_X1 U2550 ( .A1(n3287), .A2(n3286), .ZN(n2542) );
  AND2_X1 U2551 ( .A1(n3157), .A2(REG3_REG_10__SCAN_IN), .ZN(n3192) );
  INV_X1 U2552 ( .A(n3619), .ZN(n2374) );
  INV_X1 U2553 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4507) );
  AND2_X1 U2554 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2883) );
  XNOR2_X1 U2555 ( .A(n2842), .B(n3596), .ZN(n2866) );
  NAND2_X1 U2556 ( .A1(n2875), .A2(n2874), .ZN(n2935) );
  OR2_X1 U2557 ( .A1(n3084), .A2(n4573), .ZN(n3094) );
  NOR2_X1 U2558 ( .A1(n3094), .A2(n3093), .ZN(n3157) );
  NAND2_X1 U2559 ( .A1(n2725), .A2(n2724), .ZN(n2784) );
  NAND2_X1 U2560 ( .A1(n5029), .A2(n5030), .ZN(n5028) );
  NAND2_X1 U2561 ( .A1(n3480), .A2(n3481), .ZN(n5042) );
  NAND2_X1 U2562 ( .A1(n2524), .A2(n3331), .ZN(n2523) );
  INV_X1 U2563 ( .A(n3325), .ZN(n2524) );
  INV_X1 U2564 ( .A(n3331), .ZN(n2526) );
  INV_X1 U2565 ( .A(n2367), .ZN(n2366) );
  OAI21_X1 U2566 ( .B1(n2368), .B2(n2267), .A(n3661), .ZN(n2367) );
  AOI22_X1 U2567 ( .A1(n2906), .A2(n3548), .B1(n3477), .B2(n3656), .ZN(n2791)
         );
  NAND2_X1 U2568 ( .A1(n2786), .A2(n3656), .ZN(n2787) );
  OR2_X1 U2569 ( .A1(n2795), .A2(n2796), .ZN(n2847) );
  NAND2_X1 U2570 ( .A1(n3689), .A2(n3690), .ZN(n2538) );
  AOI22_X1 U2571 ( .A1(n4329), .A2(n3548), .B1(n3477), .B2(n4996), .ZN(n5000)
         );
  OAI21_X1 U2572 ( .B1(n2627), .B2(IR_REG_28__SCAN_IN), .A(n2621), .ZN(n2624)
         );
  NAND2_X1 U2573 ( .A1(n4034), .A2(n3920), .ZN(n2806) );
  AND2_X1 U2574 ( .A1(n3594), .A2(n3593), .ZN(n4128) );
  OR2_X1 U2575 ( .A1(n2802), .A2(n2954), .ZN(n2759) );
  OAI211_X1 U2576 ( .C1(n2512), .C2(REG2_REG_1__SCAN_IN), .A(n2510), .B(n2509), 
        .ZN(n3939) );
  NAND2_X1 U2577 ( .A1(n2511), .A2(n2954), .ZN(n2510) );
  NAND2_X1 U2578 ( .A1(n2512), .A2(n2281), .ZN(n2509) );
  INV_X1 U2579 ( .A(n2513), .ZN(n2511) );
  NOR2_X1 U2580 ( .A1(n2819), .A2(n2679), .ZN(n2689) );
  AND2_X1 U2581 ( .A1(n2479), .A2(n4764), .ZN(n2477) );
  INV_X1 U2582 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3045) );
  NAND2_X1 U2583 ( .A1(n2670), .A2(n2311), .ZN(n2671) );
  NAND2_X1 U2584 ( .A1(n2669), .A2(n2668), .ZN(n2311) );
  NAND2_X1 U2585 ( .A1(n2342), .A2(n2340), .ZN(n3952) );
  INV_X1 U2586 ( .A(n2343), .ZN(n2342) );
  OAI21_X1 U2587 ( .B1(n3950), .B2(n2344), .A(n2304), .ZN(n2343) );
  NAND2_X1 U2588 ( .A1(n2488), .A2(REG1_REG_10__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U2589 ( .A1(n3954), .A2(n4836), .ZN(n3955) );
  NAND2_X1 U2590 ( .A1(n2544), .A2(n2562), .ZN(n3359) );
  NAND2_X1 U2591 ( .A1(n2506), .A2(n2335), .ZN(n2505) );
  NOR2_X1 U2592 ( .A1(n2301), .A2(n3983), .ZN(n3984) );
  INV_X1 U2593 ( .A(n2352), .ZN(n2350) );
  NAND2_X1 U2594 ( .A1(n4012), .A2(n4321), .ZN(n2352) );
  INV_X1 U2595 ( .A(n4013), .ZN(n2500) );
  NAND2_X1 U2596 ( .A1(n2501), .A2(n3997), .ZN(n4014) );
  XNOR2_X1 U2597 ( .A(n4030), .B(n4029), .ZN(n4033) );
  NAND2_X1 U2598 ( .A1(n2308), .A2(n2498), .ZN(n4030) );
  AOI21_X1 U2599 ( .B1(n2272), .B2(n2499), .A(n2307), .ZN(n2498) );
  NAND2_X1 U2600 ( .A1(n3996), .A2(n2272), .ZN(n2308) );
  NOR2_X1 U2601 ( .A1(n4415), .A2(n4418), .ZN(n4414) );
  OR2_X1 U2602 ( .A1(n4134), .A2(n4069), .ZN(n2324) );
  NAND2_X1 U2603 ( .A1(n4125), .A2(n2457), .ZN(n2456) );
  NAND2_X1 U2604 ( .A1(n4152), .A2(n4129), .ZN(n2457) );
  NOR2_X1 U2605 ( .A1(n2274), .A2(n4134), .ZN(n4133) );
  INV_X1 U2606 ( .A(n3900), .ZN(n4126) );
  INV_X1 U2607 ( .A(n4066), .ZN(n4156) );
  NAND2_X1 U2608 ( .A1(n4164), .A2(n4085), .ZN(n4147) );
  NOR2_X1 U2609 ( .A1(n4150), .A2(n4167), .ZN(n4064) );
  AND2_X1 U2610 ( .A1(n4190), .A2(n4100), .ZN(n4189) );
  INV_X1 U2611 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4514) );
  INV_X1 U2612 ( .A(n3499), .ZN(n3498) );
  INV_X1 U2613 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4686) );
  INV_X1 U2614 ( .A(n2417), .ZN(n2416) );
  AOI21_X1 U2615 ( .B1(n2417), .B2(n2415), .A(n2414), .ZN(n2413) );
  AND2_X1 U2616 ( .A1(n2418), .A2(n3888), .ZN(n2417) );
  OR2_X1 U2617 ( .A1(n3453), .A2(n3452), .ZN(n3468) );
  NAND2_X1 U2618 ( .A1(n3467), .A2(REG3_REG_20__SCAN_IN), .ZN(n3484) );
  INV_X1 U2619 ( .A(n3468), .ZN(n3467) );
  NAND2_X1 U2620 ( .A1(n4326), .A2(n2418), .ZN(n4255) );
  NAND2_X1 U2621 ( .A1(n3436), .A2(REG3_REG_18__SCAN_IN), .ZN(n3453) );
  NAND2_X1 U2622 ( .A1(n2436), .A2(n2433), .ZN(n4299) );
  AOI21_X1 U2623 ( .B1(n2435), .B2(n2438), .A(n2434), .ZN(n2433) );
  NOR2_X1 U2624 ( .A1(n4293), .A2(n4317), .ZN(n2434) );
  NAND2_X1 U2625 ( .A1(n4326), .A2(n4078), .ZN(n4310) );
  NOR2_X1 U2626 ( .A1(n4335), .A2(n4317), .ZN(n4319) );
  NOR2_X1 U2627 ( .A1(n3385), .A2(n3384), .ZN(n3402) );
  NAND2_X1 U2628 ( .A1(n4327), .A2(n4333), .ZN(n4326) );
  NOR2_X1 U2629 ( .A1(n4364), .A2(n2382), .ZN(n2381) );
  INV_X1 U2630 ( .A(n4076), .ZN(n2382) );
  NAND2_X1 U2631 ( .A1(n2383), .A2(n4076), .ZN(n4347) );
  INV_X1 U2632 ( .A(n4996), .ZN(n4351) );
  AND2_X1 U2633 ( .A1(n4398), .A2(n4370), .ZN(n4377) );
  NAND2_X1 U2634 ( .A1(n3758), .A2(n3836), .ZN(n4075) );
  NOR2_X1 U2635 ( .A1(n2273), .A2(n4399), .ZN(n4398) );
  NAND2_X1 U2636 ( .A1(n3192), .A2(REG3_REG_11__SCAN_IN), .ZN(n3227) );
  AND2_X1 U2637 ( .A1(n3831), .A2(n3818), .ZN(n4041) );
  AOI21_X1 U2638 ( .B1(n2388), .B2(n2390), .A(n2386), .ZN(n2385) );
  INV_X1 U2639 ( .A(n3829), .ZN(n2386) );
  NAND2_X1 U2640 ( .A1(n2387), .A2(n3815), .ZN(n3220) );
  NAND2_X1 U2641 ( .A1(n3188), .A2(n3827), .ZN(n2387) );
  NAND2_X1 U2642 ( .A1(n2462), .A2(n2461), .ZN(n3213) );
  NOR2_X1 U2643 ( .A1(n2895), .A2(n3045), .ZN(n3039) );
  OAI21_X1 U2644 ( .B1(n3008), .B2(n2408), .A(n2407), .ZN(n3091) );
  AND2_X1 U2645 ( .A1(n2404), .A2(n3825), .ZN(n2407) );
  OR2_X1 U2646 ( .A1(n2411), .A2(n2405), .ZN(n2404) );
  NAND2_X1 U2647 ( .A1(n2406), .A2(n2410), .ZN(n3090) );
  NAND2_X1 U2648 ( .A1(n3008), .A2(n2411), .ZN(n2406) );
  NAND2_X1 U2649 ( .A1(n2409), .A2(n3808), .ZN(n3059) );
  OR2_X1 U2650 ( .A1(n3008), .A2(n2972), .ZN(n2409) );
  OR2_X1 U2651 ( .A1(n3018), .A2(n3019), .ZN(n3016) );
  NAND2_X1 U2652 ( .A1(n2455), .A2(n2453), .ZN(n3011) );
  NOR2_X1 U2653 ( .A1(n2268), .A2(n2454), .ZN(n2453) );
  NAND2_X1 U2654 ( .A1(n2971), .A2(n3804), .ZN(n3008) );
  AND2_X1 U2655 ( .A1(n3804), .A2(n3801), .ZN(n3892) );
  NAND2_X1 U2656 ( .A1(n2913), .A2(n2912), .ZN(n2989) );
  OR2_X1 U2657 ( .A1(n3882), .A2(n3867), .ZN(n2913) );
  NAND2_X1 U2658 ( .A1(n2911), .A2(n4034), .ZN(n4397) );
  NAND2_X1 U2659 ( .A1(n2918), .A2(n2917), .ZN(n4880) );
  INV_X1 U2660 ( .A(n4939), .ZN(n4417) );
  INV_X1 U2661 ( .A(n4407), .ZN(n4418) );
  NOR2_X1 U2662 ( .A1(n4245), .A2(n4058), .ZN(n4227) );
  INV_X1 U2663 ( .A(IR_REG_7__SCAN_IN), .ZN(n4717) );
  OR2_X1 U2664 ( .A1(n4264), .A2(n4099), .ZN(n4245) );
  INV_X1 U2665 ( .A(n5026), .ZN(n4284) );
  NOR2_X1 U2666 ( .A1(n4335), .A2(n2325), .ZN(n4301) );
  INV_X1 U2667 ( .A(n2327), .ZN(n2325) );
  NAND2_X1 U2668 ( .A1(n4377), .A2(n4351), .ZN(n4353) );
  OR2_X1 U2669 ( .A1(n4353), .A2(n4328), .ZN(n4335) );
  AND2_X1 U2670 ( .A1(n4929), .A2(n2319), .ZN(n3272) );
  AND2_X1 U2671 ( .A1(n2321), .A2(n2320), .ZN(n2319) );
  NAND2_X1 U2672 ( .A1(n4929), .A2(n4940), .ZN(n4928) );
  NOR2_X1 U2673 ( .A1(n3016), .A2(n3055), .ZN(n3063) );
  AND2_X1 U2674 ( .A1(n3063), .A2(n2465), .ZN(n4929) );
  NAND2_X1 U2675 ( .A1(n2314), .A2(n2947), .ZN(n2996) );
  NOR2_X1 U2676 ( .A1(n2996), .A2(n2995), .ZN(n2998) );
  INV_X1 U2677 ( .A(n5010), .ZN(n5015) );
  AND3_X1 U2678 ( .A1(n2983), .A2(n2982), .A3(n2981), .ZN(n3003) );
  AND2_X1 U2679 ( .A1(n2545), .A2(n2430), .ZN(n2429) );
  AND2_X1 U2680 ( .A1(n2622), .A2(n2431), .ZN(n2430) );
  INV_X1 U2681 ( .A(IR_REG_29__SCAN_IN), .ZN(n2431) );
  AND2_X1 U2682 ( .A1(n2317), .A2(IR_REG_31__SCAN_IN), .ZN(n2627) );
  NOR2_X1 U2683 ( .A1(n2569), .A2(IR_REG_22__SCAN_IN), .ZN(n2546) );
  AND2_X1 U2684 ( .A1(n2579), .A2(n2578), .ZN(n2620) );
  XNOR2_X1 U2685 ( .A(n2581), .B(n2476), .ZN(n3908) );
  AND2_X1 U2686 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2595)
         );
  INV_X1 U2687 ( .A(n3392), .ZN(n2584) );
  NAND2_X1 U2688 ( .A1(n3190), .A2(IR_REG_1__SCAN_IN), .ZN(n2513) );
  OAI21_X1 U2689 ( .B1(IR_REG_0__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(n2497), 
        .ZN(n2512) );
  NAND2_X1 U2690 ( .A1(n2507), .A2(IR_REG_0__SCAN_IN), .ZN(n2497) );
  NAND2_X1 U2691 ( .A1(n2508), .A2(IR_REG_31__SCAN_IN), .ZN(n2507) );
  INV_X1 U2692 ( .A(IR_REG_1__SCAN_IN), .ZN(n2508) );
  AND2_X1 U2693 ( .A1(n2375), .A2(n3123), .ZN(n3617) );
  NAND2_X1 U2694 ( .A1(n2375), .A2(n2373), .ZN(n3618) );
  INV_X1 U2695 ( .A(n2535), .ZN(n2534) );
  OAI21_X1 U2696 ( .B1(n2536), .B2(n3745), .A(n3743), .ZN(n2535) );
  NAND2_X1 U2697 ( .A1(n2542), .A2(n3291), .ZN(n3316) );
  XNOR2_X1 U2698 ( .A(n2790), .B(n2791), .ZN(n3654) );
  NAND2_X1 U2699 ( .A1(n2520), .A2(n3331), .ZN(n3356) );
  NAND2_X1 U2700 ( .A1(n3326), .A2(n3325), .ZN(n2520) );
  NAND2_X1 U2701 ( .A1(n2537), .A2(n2536), .ZN(n2533) );
  NAND2_X1 U2702 ( .A1(n2261), .A2(DATAI_0_), .ZN(n2714) );
  INV_X1 U2703 ( .A(n4057), .ZN(n5049) );
  NAND2_X1 U2704 ( .A1(n5028), .A2(n3466), .ZN(n5043) );
  NAND2_X1 U2705 ( .A1(n2279), .A2(n2528), .ZN(n2527) );
  NAND2_X1 U2706 ( .A1(n2530), .A2(n2880), .ZN(n2528) );
  NAND2_X1 U2707 ( .A1(n2750), .A2(n4950), .ZN(n5050) );
  INV_X1 U2708 ( .A(n4128), .ZN(n4070) );
  OR2_X1 U2709 ( .A1(n4193), .A2(n3603), .ZN(n3544) );
  OAI211_X1 U2710 ( .C1(n4247), .C2(n3603), .A(n3489), .B(n3488), .ZN(n5039)
         );
  NAND4_X1 U2711 ( .A1(n3459), .A2(n3458), .A3(n3457), .A4(n3456), .ZN(n5046)
         );
  OR2_X1 U2712 ( .A1(n2802), .A2(n2774), .ZN(n2775) );
  OR2_X1 U2713 ( .A1(n2802), .A2(n4889), .ZN(n2709) );
  INV_X2 U2714 ( .A(U4043), .ZN(n3932) );
  NAND2_X1 U2715 ( .A1(n2503), .A2(n2636), .ZN(n2502) );
  NAND2_X1 U2716 ( .A1(n2833), .A2(n2832), .ZN(n2503) );
  XNOR2_X1 U2717 ( .A(n2479), .B(n2478), .ZN(n2650) );
  XNOR2_X1 U2718 ( .A(n2663), .B(n4927), .ZN(n4807) );
  NAND2_X1 U2719 ( .A1(n4807), .A2(REG1_REG_6__SCAN_IN), .ZN(n4806) );
  XNOR2_X1 U2720 ( .A(n2680), .B(n4927), .ZN(n4802) );
  INV_X1 U2721 ( .A(n2514), .ZN(n4801) );
  INV_X1 U2722 ( .A(n2765), .ZN(n2359) );
  NAND2_X1 U2723 ( .A1(n2684), .A2(REG2_REG_8__SCAN_IN), .ZN(n3949) );
  XNOR2_X1 U2724 ( .A(n3952), .B(n3951), .ZN(n4825) );
  NOR2_X1 U2725 ( .A1(n4841), .A2(n3968), .ZN(n4853) );
  XNOR2_X1 U2726 ( .A(n3979), .B(n4759), .ZN(n3970) );
  NAND2_X1 U2727 ( .A1(n2335), .A2(n2334), .ZN(n3958) );
  AND2_X1 U2728 ( .A1(n2331), .A2(n2332), .ZN(n2334) );
  NAND2_X1 U2729 ( .A1(n3985), .A2(n3984), .ZN(n3990) );
  INV_X1 U2730 ( .A(n2484), .ZN(n2483) );
  AOI21_X1 U2731 ( .B1(n2484), .B2(n2482), .A(n2269), .ZN(n2481) );
  INV_X1 U2732 ( .A(n2309), .ZN(n4872) );
  NAND2_X1 U2733 ( .A1(n4865), .A2(n4005), .ZN(n4019) );
  NAND2_X1 U2734 ( .A1(n2351), .A2(n2352), .ZN(n4021) );
  NAND2_X1 U2735 ( .A1(n4014), .A2(n2272), .ZN(n4028) );
  OAI21_X1 U2736 ( .B1(n4115), .B2(n4946), .A(n4114), .ZN(n4116) );
  NOR2_X1 U2737 ( .A1(n4113), .A2(n4112), .ZN(n4114) );
  AND2_X1 U2738 ( .A1(n4111), .A2(n4944), .ZN(n4112) );
  AND2_X1 U2739 ( .A1(n3572), .A2(n3557), .ZN(n4155) );
  NAND2_X1 U2740 ( .A1(n2449), .A2(n2263), .ZN(n4180) );
  OR2_X1 U2741 ( .A1(n4230), .A2(n2452), .ZN(n2449) );
  NAND2_X1 U2742 ( .A1(n4230), .A2(n4059), .ZN(n4198) );
  OR2_X1 U2743 ( .A1(n4357), .A2(n2440), .ZN(n2432) );
  NAND2_X1 U2744 ( .A1(n2443), .A2(n2444), .ZN(n4334) );
  NAND2_X1 U2745 ( .A1(n4357), .A2(n4054), .ZN(n2443) );
  NAND2_X1 U2746 ( .A1(n2467), .A2(n2464), .ZN(n4932) );
  NAND2_X1 U2747 ( .A1(n2945), .A2(n2908), .ZN(n2987) );
  INV_X1 U2748 ( .A(n4338), .ZN(n5059) );
  AND2_X1 U2749 ( .A1(n4406), .A2(n2944), .ZN(n4325) );
  OR2_X1 U2750 ( .A1(n2262), .A2(n4034), .ZN(n4885) );
  INV_X1 U2751 ( .A(n4950), .ZN(n4897) );
  AND2_X2 U2752 ( .A1(n3003), .A2(n2984), .ZN(n5022) );
  OAI21_X1 U2753 ( .B1(n4423), .B2(n5007), .A(n2329), .ZN(n4494) );
  INV_X1 U2754 ( .A(n4422), .ZN(n2330) );
  NAND2_X1 U2755 ( .A1(n2740), .A2(n2742), .ZN(n4769) );
  XNOR2_X1 U2756 ( .A(n2574), .B(IR_REG_26__SCAN_IN), .ZN(n2737) );
  INV_X1 U2757 ( .A(n3908), .ZN(n3797) );
  CLKBUF_X1 U2758 ( .A(n2748), .Z(n4936) );
  NOR2_X1 U2759 ( .A1(n2660), .A2(n2659), .ZN(n4762) );
  AOI21_X1 U2760 ( .B1(n3713), .B2(n5048), .A(n3712), .ZN(n3714) );
  NOR2_X1 U2761 ( .A1(n4864), .A2(n2502), .ZN(n2837) );
  NOR2_X1 U2762 ( .A1(n2358), .A2(n4864), .ZN(n2773) );
  NAND2_X1 U2763 ( .A1(n4817), .A2(n4818), .ZN(n4816) );
  NAND2_X1 U2764 ( .A1(n2422), .A2(n2420), .ZN(U3547) );
  OR2_X1 U2765 ( .A1(n5022), .A2(n2421), .ZN(n2420) );
  NAND2_X1 U2766 ( .A1(n4494), .A2(n5022), .ZN(n2422) );
  INV_X1 U2767 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2421) );
  AND3_X1 U2768 ( .A1(n2429), .A2(n2473), .A3(n2544), .ZN(n2704) );
  AND2_X1 U2769 ( .A1(n2450), .A2(n4062), .ZN(n2263) );
  NAND2_X1 U2770 ( .A1(n2785), .A2(n2312), .ZN(n3656) );
  NAND2_X1 U2771 ( .A1(n2544), .A2(n2543), .ZN(n2580) );
  NAND2_X1 U2772 ( .A1(n2474), .A2(n2544), .ZN(n2264) );
  AND2_X1 U2773 ( .A1(n2279), .A2(n2874), .ZN(n2265) );
  AND2_X1 U2774 ( .A1(n2473), .A2(n2544), .ZN(n2587) );
  AND2_X1 U2775 ( .A1(n2288), .A2(n2309), .ZN(n3996) );
  INV_X1 U2776 ( .A(n3996), .ZN(n2501) );
  OR2_X1 U2777 ( .A1(n3355), .A2(n2526), .ZN(n2525) );
  AND2_X1 U2778 ( .A1(n3295), .A2(n3291), .ZN(n2266) );
  INV_X1 U2779 ( .A(n3080), .ZN(n2465) );
  AND2_X1 U2780 ( .A1(n2540), .A2(n5042), .ZN(n2267) );
  INV_X1 U2781 ( .A(n3319), .ZN(n2320) );
  AND2_X1 U2782 ( .A1(n3805), .A2(n3808), .ZN(n2268) );
  NAND2_X1 U2783 ( .A1(n4929), .A2(n2322), .ZN(n2323) );
  NOR2_X1 U2784 ( .A1(n2486), .A2(n2485), .ZN(n2269) );
  AND2_X1 U2785 ( .A1(n3984), .A2(n4003), .ZN(n2270) );
  AND2_X1 U2786 ( .A1(n2332), .A2(REG2_REG_14__SCAN_IN), .ZN(n2271) );
  NOR2_X1 U2787 ( .A1(n4015), .A2(n2500), .ZN(n2272) );
  INV_X1 U2788 ( .A(n2551), .ZN(n2355) );
  OR2_X1 U2789 ( .A1(n3270), .A2(n4040), .ZN(n2273) );
  OR2_X1 U2790 ( .A1(n4172), .A2(n4156), .ZN(n2274) );
  OR2_X1 U2791 ( .A1(n2680), .A2(n4927), .ZN(n2275) );
  NAND2_X1 U2792 ( .A1(n2339), .A2(n2336), .ZN(n2335) );
  NAND2_X1 U2793 ( .A1(n2575), .A2(n2737), .ZN(n2715) );
  NAND4_X1 U2794 ( .A1(n2712), .A2(n2711), .A3(n2710), .A4(n2709), .ZN(n2907)
         );
  OAI21_X1 U2795 ( .B1(n5029), .B2(n2368), .A(n2366), .ZN(n3724) );
  NAND2_X1 U2796 ( .A1(n2531), .A2(n2534), .ZN(n3626) );
  INV_X1 U2797 ( .A(n2533), .ZN(n3670) );
  AND2_X1 U2798 ( .A1(n2619), .A2(n2651), .ZN(n4764) );
  INV_X1 U2799 ( .A(n4764), .ZN(n2478) );
  AND2_X1 U2800 ( .A1(n4421), .A2(n5010), .ZN(n2276) );
  AND4_X1 U2801 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2744), .ZN(n2277)
         );
  NAND2_X1 U2802 ( .A1(n4293), .A2(n4317), .ZN(n2278) );
  XNOR2_X1 U2803 ( .A(n2789), .B(n3596), .ZN(n2790) );
  INV_X1 U2804 ( .A(IR_REG_3__SCAN_IN), .ZN(n2617) );
  OR2_X1 U2805 ( .A1(n3024), .A2(n3025), .ZN(n2279) );
  AND2_X1 U2806 ( .A1(n3131), .A2(n3130), .ZN(n2280) );
  NAND2_X1 U2807 ( .A1(n3518), .A2(n3517), .ZN(n3645) );
  AND2_X1 U2808 ( .A1(REG2_REG_1__SCAN_IN), .A2(n2513), .ZN(n2281) );
  AND2_X1 U2809 ( .A1(n2351), .A2(n2348), .ZN(n2282) );
  INV_X1 U2810 ( .A(n2522), .ZN(n2521) );
  OAI21_X1 U2811 ( .B1(n2523), .B2(n3355), .A(n3354), .ZN(n2522) );
  AND2_X1 U2812 ( .A1(n4014), .A2(n4013), .ZN(n2283) );
  AND2_X1 U2813 ( .A1(n4063), .A2(n4100), .ZN(n2284) );
  NAND2_X1 U2814 ( .A1(n3208), .A2(n3252), .ZN(n2285) );
  NAND2_X1 U2815 ( .A1(n2400), .A2(n3782), .ZN(n2396) );
  NAND2_X1 U2816 ( .A1(n2401), .A2(n3851), .ZN(n2400) );
  AND2_X1 U2817 ( .A1(n4765), .A2(REG1_REG_2__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U2818 ( .A1(n4126), .A2(n2398), .ZN(n2287) );
  OR2_X1 U2819 ( .A1(n4003), .A2(n3992), .ZN(n2288) );
  NOR2_X1 U2820 ( .A1(n3124), .A2(n2374), .ZN(n2373) );
  NAND2_X1 U2821 ( .A1(n4209), .A2(n4191), .ZN(n2289) );
  NAND2_X1 U2822 ( .A1(n2587), .A2(n2546), .ZN(n2290) );
  AND2_X1 U2823 ( .A1(n2395), .A2(n4089), .ZN(n2394) );
  INV_X1 U2824 ( .A(n3477), .ZN(n3533) );
  INV_X1 U2825 ( .A(n3928), .ZN(n2466) );
  NAND2_X1 U2826 ( .A1(n4930), .A2(n3208), .ZN(n3251) );
  INV_X1 U2827 ( .A(n3823), .ZN(n2425) );
  NAND2_X1 U2828 ( .A1(n3699), .A2(n3432), .ZN(n2291) );
  NAND2_X1 U2829 ( .A1(n2432), .A2(n2438), .ZN(n4308) );
  NAND2_X1 U2830 ( .A1(n3314), .A2(n3300), .ZN(n3326) );
  NAND2_X1 U2831 ( .A1(n2538), .A2(n3418), .ZN(n3697) );
  AND2_X1 U2832 ( .A1(n3555), .A2(n3521), .ZN(n2292) );
  OR2_X1 U2833 ( .A1(n2596), .A2(n2595), .ZN(n2293) );
  INV_X1 U2834 ( .A(IR_REG_21__SCAN_IN), .ZN(n2476) );
  INV_X1 U2835 ( .A(IR_REG_30__SCAN_IN), .ZN(n3350) );
  AND2_X1 U2836 ( .A1(n4314), .A2(n4328), .ZN(n2294) );
  NAND4_X1 U2837 ( .A1(n2560), .A2(n2615), .A3(n2559), .A4(n2558), .ZN(n3153)
         );
  OR2_X1 U2838 ( .A1(n5046), .A2(n5026), .ZN(n2295) );
  AND2_X1 U2839 ( .A1(n3508), .A2(n3507), .ZN(n2296) );
  AOI21_X1 U2840 ( .B1(n2267), .B2(n2541), .A(n2298), .ZN(n2539) );
  INV_X1 U2841 ( .A(n4080), .ZN(n2414) );
  AND2_X1 U2842 ( .A1(n3579), .A2(n3578), .ZN(n4152) );
  INV_X1 U2843 ( .A(n4152), .ZN(n4067) );
  NAND2_X1 U2844 ( .A1(n3409), .A2(IR_REG_31__SCAN_IN), .ZN(n2297) );
  INV_X1 U2845 ( .A(IR_REG_28__SCAN_IN), .ZN(n2622) );
  NAND2_X1 U2846 ( .A1(n5041), .A2(n3660), .ZN(n2298) );
  AND2_X1 U2847 ( .A1(n2291), .A2(n3418), .ZN(n2299) );
  AND2_X1 U2848 ( .A1(n2292), .A2(n2532), .ZN(n2300) );
  OAI21_X1 U2849 ( .B1(n2261), .B2(n3934), .A(n2714), .ZN(n3795) );
  AND2_X1 U2850 ( .A1(n4758), .A2(REG1_REG_15__SCAN_IN), .ZN(n2301) );
  OAI21_X1 U2851 ( .B1(n3178), .B2(n3177), .A(n3176), .ZN(n3287) );
  NAND2_X1 U2852 ( .A1(n2935), .A2(n2880), .ZN(n3026) );
  INV_X1 U2853 ( .A(n2408), .ZN(n2410) );
  NAND2_X1 U2854 ( .A1(n2455), .A2(n2964), .ZN(n3009) );
  INV_X1 U2855 ( .A(n2487), .ZN(n2486) );
  OR2_X1 U2856 ( .A1(n4335), .A2(n2326), .ZN(n2302) );
  NAND3_X1 U2857 ( .A1(n2473), .A2(n2544), .A3(n2545), .ZN(n2303) );
  OR2_X1 U2858 ( .A1(n4959), .A2(n3096), .ZN(n2304) );
  NAND2_X1 U2859 ( .A1(n2529), .A2(n2527), .ZN(n3121) );
  NAND2_X1 U2860 ( .A1(n2847), .A2(n2846), .ZN(n2865) );
  AND2_X1 U2861 ( .A1(n4929), .A2(n2321), .ZN(n2305) );
  INV_X1 U2862 ( .A(IR_REG_27__SCAN_IN), .ZN(n2316) );
  INV_X1 U2863 ( .A(n4129), .ZN(n4134) );
  INV_X1 U2864 ( .A(n4003), .ZN(n2485) );
  NAND2_X1 U2865 ( .A1(n3033), .A2(n3034), .ZN(n2306) );
  NOR2_X1 U2866 ( .A1(n4027), .A2(n4471), .ZN(n2307) );
  INV_X1 U2867 ( .A(n2354), .ZN(n2353) );
  NOR2_X1 U2868 ( .A1(n4012), .A2(n4321), .ZN(n2354) );
  INV_X1 U2869 ( .A(n2349), .ZN(n2348) );
  OR2_X1 U2870 ( .A1(n4022), .A2(n2350), .ZN(n2349) );
  AND2_X1 U2871 ( .A1(n2667), .A2(n2666), .ZN(n4761) );
  INV_X1 U2872 ( .A(n4761), .ZN(n2496) );
  INV_X1 U2873 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2495) );
  INV_X1 U2874 ( .A(IR_REG_8__SCAN_IN), .ZN(n4721) );
  INV_X1 U2875 ( .A(IR_REG_4__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U2876 ( .A1(n2692), .A2(n2693), .ZN(n2691) );
  XNOR2_X1 U2877 ( .A(n3963), .B(n3951), .ZN(n2488) );
  NOR2_X1 U2878 ( .A1(n2829), .A2(n2828), .ZN(n2827) );
  NAND2_X1 U2879 ( .A1(n2317), .A2(n2315), .ZN(n2621) );
  NAND2_X1 U2880 ( .A1(n2474), .A2(n2318), .ZN(n2317) );
  INV_X2 U2881 ( .A(n3357), .ZN(n2544) );
  INV_X1 U2882 ( .A(n2323), .ZN(n3171) );
  INV_X1 U2883 ( .A(n2328), .ZN(n4264) );
  NAND3_X1 U2884 ( .A1(n2335), .A2(n2331), .A3(n2271), .ZN(n2506) );
  NAND2_X1 U2885 ( .A1(n2684), .A2(n2341), .ZN(n2340) );
  NAND2_X1 U2886 ( .A1(n4019), .A2(n2347), .ZN(n2345) );
  NAND2_X1 U2887 ( .A1(n2345), .A2(n2346), .ZN(n4031) );
  NAND2_X1 U2888 ( .A1(n4019), .A2(n2353), .ZN(n2351) );
  NAND2_X1 U2889 ( .A1(n2514), .A2(n2356), .ZN(n2682) );
  XNOR2_X1 U2890 ( .A(n2683), .B(n2359), .ZN(n2358) );
  INV_X1 U2891 ( .A(n5029), .ZN(n2365) );
  OAI21_X2 U2892 ( .B1(n2365), .B2(n2363), .A(n2361), .ZN(n3644) );
  INV_X1 U2893 ( .A(n2539), .ZN(n2368) );
  NAND2_X1 U2894 ( .A1(n2795), .A2(n2846), .ZN(n2370) );
  NAND2_X1 U2895 ( .A1(n2796), .A2(n2846), .ZN(n2369) );
  NAND3_X1 U2896 ( .A1(n2370), .A2(n2864), .A3(n2369), .ZN(n2870) );
  NAND2_X1 U2897 ( .A1(n3121), .A2(n2373), .ZN(n2371) );
  NAND2_X1 U2898 ( .A1(n2371), .A2(n2372), .ZN(n3178) );
  OR3_X1 U2899 ( .A1(n2596), .A2(n2377), .A3(n2595), .ZN(n2745) );
  XNOR2_X1 U2900 ( .A(n2380), .B(IR_REG_20__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U2901 ( .A1(n2383), .A2(n2381), .ZN(n4345) );
  NAND2_X1 U2902 ( .A1(n3188), .A2(n2388), .ZN(n2384) );
  NAND2_X1 U2903 ( .A1(n2384), .A2(n2385), .ZN(n3262) );
  NAND2_X1 U2904 ( .A1(n4164), .A2(n2394), .ZN(n2391) );
  NAND2_X1 U2905 ( .A1(n2391), .A2(n2392), .ZN(n4091) );
  NAND2_X1 U2906 ( .A1(n4164), .A2(n2402), .ZN(n2397) );
  INV_X1 U2907 ( .A(n3808), .ZN(n2412) );
  OAI21_X1 U2908 ( .B1(n4327), .B2(n2416), .A(n2413), .ZN(n4240) );
  NAND4_X1 U2909 ( .A1(n2473), .A2(n2544), .A3(n2545), .A4(n2622), .ZN(n2601)
         );
  OAI21_X1 U2910 ( .B1(n4240), .B2(n4083), .A(n4082), .ZN(n4182) );
  NAND2_X1 U2911 ( .A1(n3091), .A2(n3810), .ZN(n4938) );
  NAND2_X1 U2912 ( .A1(n4182), .A2(n4084), .ZN(n4164) );
  NAND2_X1 U2913 ( .A1(n4388), .A2(n3833), .ZN(n3758) );
  OAI21_X1 U2914 ( .B1(n4037), .B2(n2557), .A(n4036), .ZN(n4039) );
  NAND2_X1 U2915 ( .A1(n2830), .A2(n2831), .ZN(n2636) );
  NAND2_X1 U2916 ( .A1(n4357), .A2(n2437), .ZN(n2436) );
  NAND2_X1 U2917 ( .A1(n4230), .A2(n2448), .ZN(n2447) );
  INV_X1 U2918 ( .A(n2964), .ZN(n2454) );
  NAND2_X1 U2919 ( .A1(n2961), .A2(n2960), .ZN(n2455) );
  NAND2_X1 U2920 ( .A1(n3082), .A2(n2463), .ZN(n2462) );
  NAND2_X1 U2921 ( .A1(n2467), .A2(n2463), .ZN(n4930) );
  OR2_X1 U2922 ( .A1(n3082), .A2(n3081), .ZN(n2467) );
  NAND3_X1 U2923 ( .A1(n2945), .A2(n2908), .A3(n2914), .ZN(n2985) );
  NAND2_X1 U2924 ( .A1(n3985), .A2(n2270), .ZN(n2480) );
  OAI211_X1 U2925 ( .C1(n3985), .C2(n2483), .A(n2481), .B(n2480), .ZN(n4871)
         );
  NOR2_X1 U2926 ( .A1(n3991), .A2(n5011), .ZN(n2487) );
  OAI211_X1 U2927 ( .C1(n2488), .C2(REG1_REG_10__SCAN_IN), .A(n4822), .B(n4870), .ZN(n4828) );
  NAND2_X1 U2928 ( .A1(n2492), .A2(n4806), .ZN(n2491) );
  NAND2_X1 U2929 ( .A1(n2491), .A2(n2494), .ZN(n2669) );
  MUX2_X1 U2930 ( .A(REG1_REG_1__SCAN_IN), .B(n2610), .S(n4766), .Z(n2612) );
  INV_X1 U2931 ( .A(n2506), .ZN(n3973) );
  INV_X1 U2932 ( .A(n2505), .ZN(n3977) );
  INV_X1 U2933 ( .A(n3326), .ZN(n2519) );
  NAND2_X1 U2934 ( .A1(n2875), .A2(n2265), .ZN(n2529) );
  NAND2_X1 U2935 ( .A1(n3024), .A2(n3025), .ZN(n2530) );
  NAND2_X1 U2936 ( .A1(n3645), .A2(n2292), .ZN(n2537) );
  OAI22_X1 U2937 ( .A1(n3626), .A2(n3627), .B1(n3583), .B2(n3584), .ZN(n3602)
         );
  NAND2_X1 U2938 ( .A1(n3645), .A2(n2300), .ZN(n2531) );
  INV_X1 U2939 ( .A(n3554), .ZN(n2536) );
  NAND2_X1 U2940 ( .A1(n2538), .A2(n2299), .ZN(n3435) );
  NAND2_X1 U2941 ( .A1(n2542), .A2(n2266), .ZN(n3314) );
  NAND2_X1 U2942 ( .A1(n2587), .A2(n2589), .ZN(n2570) );
  OAI22_X1 U2943 ( .A1(n2655), .A2(n4917), .B1(n2654), .B2(n2653), .ZN(n2692)
         );
  NOR2_X1 U2944 ( .A1(n2689), .A2(n2688), .ZN(n2687) );
  NAND2_X1 U2945 ( .A1(n4035), .A2(n4034), .ZN(n4036) );
  INV_X1 U2946 ( .A(n3962), .ZN(n2670) );
  AOI21_X2 U2947 ( .B1(n3732), .B2(n3734), .A(n3733), .ZN(n5029) );
  AND2_X1 U2948 ( .A1(n4051), .A2(n4050), .ZN(n2550) );
  OR2_X1 U2949 ( .A1(n2808), .A2(n3919), .ZN(n4991) );
  OR3_X1 U2950 ( .A1(n2808), .A2(n4755), .A3(n2806), .ZN(n5032) );
  OAI211_X1 U2951 ( .C1(n3607), .C2(n4505), .A(n3502), .B(n3501), .ZN(n4242)
         );
  AND2_X1 U2952 ( .A1(n3411), .A2(n3410), .ZN(n4003) );
  AND2_X1 U2953 ( .A1(n4757), .A2(REG2_REG_18__SCAN_IN), .ZN(n2551) );
  OR2_X1 U2954 ( .A1(n4224), .A2(n4060), .ZN(n2552) );
  AND2_X1 U2955 ( .A1(n3381), .A2(n3380), .ZN(n2553) );
  INV_X1 U2956 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3452) );
  AND2_X1 U2957 ( .A1(n2800), .A2(REG1_REG_3__SCAN_IN), .ZN(n2554) );
  INV_X1 U2958 ( .A(n4116), .ZN(n4425) );
  NOR2_X1 U2959 ( .A1(n4049), .A2(n4048), .ZN(n2555) );
  INV_X1 U2960 ( .A(n3203), .ZN(n3170) );
  INV_X1 U2961 ( .A(n4221), .ZN(n4058) );
  AND2_X1 U2962 ( .A1(n3674), .A2(n3708), .ZN(n2556) );
  OR2_X1 U2963 ( .A1(n4823), .A2(n4034), .ZN(n2557) );
  NOR2_X1 U2964 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2564)
         );
  NAND2_X1 U2965 ( .A1(n4070), .A2(n4069), .ZN(n4071) );
  INV_X1 U2966 ( .A(n3317), .ZN(n3295) );
  AND2_X1 U2967 ( .A1(n3863), .A2(n4163), .ZN(n4085) );
  INV_X1 U2968 ( .A(n2306), .ZN(n3122) );
  INV_X1 U2969 ( .A(n2786), .ZN(n3598) );
  AOI21_X1 U2970 ( .B1(n3382), .B2(n3634), .A(n2553), .ZN(n3397) );
  INV_X1 U2971 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4573) );
  INV_X1 U2972 ( .A(n4937), .ZN(n3083) );
  INV_X1 U2973 ( .A(n3123), .ZN(n3124) );
  NAND2_X1 U2974 ( .A1(n2261), .A2(DATAI_1_), .ZN(n2785) );
  NAND2_X1 U2975 ( .A1(n2788), .A2(n2787), .ZN(n2789) );
  NOR2_X1 U2976 ( .A1(n3679), .A2(n2556), .ZN(n3555) );
  INV_X1 U2977 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3093) );
  AND2_X1 U2978 ( .A1(n3305), .A2(n3304), .ZN(n3328) );
  OR2_X1 U2979 ( .A1(n3538), .A2(n4507), .ZN(n3556) );
  OR2_X1 U2980 ( .A1(n3227), .A2(n4684), .ZN(n3237) );
  AND2_X1 U2981 ( .A1(n2678), .A2(n4763), .ZN(n2679) );
  INV_X1 U2982 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4029) );
  NAND2_X1 U2983 ( .A1(n3498), .A2(REG3_REG_22__SCAN_IN), .ZN(n3509) );
  AND2_X1 U2984 ( .A1(n3419), .A2(REG3_REG_17__SCAN_IN), .ZN(n3436) );
  AND2_X1 U2985 ( .A1(n3402), .A2(REG3_REG_16__SCAN_IN), .ZN(n3419) );
  NOR2_X1 U2986 ( .A1(n2555), .A2(n2550), .ZN(n4052) );
  OR2_X1 U2987 ( .A1(n2756), .A2(n2755), .ZN(n2980) );
  INV_X1 U2988 ( .A(IR_REG_22__SCAN_IN), .ZN(n2589) );
  INV_X1 U2989 ( .A(n2620), .ZN(n2625) );
  INV_X1 U2990 ( .A(n3128), .ZN(n4940) );
  INV_X1 U2991 ( .A(n2959), .ZN(n2962) );
  AND2_X1 U2992 ( .A1(n2743), .A2(n2742), .ZN(n2758) );
  OR2_X1 U2993 ( .A1(n4120), .A2(n3603), .ZN(n3594) );
  OR2_X1 U2994 ( .A1(n3484), .A2(n4686), .ZN(n3499) );
  INV_X1 U2995 ( .A(n4967), .ZN(n3951) );
  INV_X1 U2996 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4684) );
  NAND2_X1 U2997 ( .A1(n3982), .A2(n3981), .ZN(n3985) );
  AND2_X1 U2998 ( .A1(n2756), .A2(n4767), .ZN(n2629) );
  INV_X1 U2999 ( .A(n3851), .ZN(n4086) );
  INV_X1 U3000 ( .A(n3761), .ZN(n4300) );
  NAND2_X1 U3001 ( .A1(n2262), .A2(n4876), .ZN(n4939) );
  NAND2_X1 U3002 ( .A1(n4755), .A2(n2917), .ZN(n4941) );
  OR2_X1 U3003 ( .A1(n3263), .A2(n4041), .ZN(n3265) );
  INV_X1 U3004 ( .A(n4878), .ZN(n4946) );
  XNOR2_X1 U3005 ( .A(n2590), .B(n2589), .ZN(n2720) );
  AND2_X1 U3006 ( .A1(n2648), .A2(IR_REG_31__SCAN_IN), .ZN(n2665) );
  AND2_X1 U3007 ( .A1(n2625), .A2(STATE_REG_SCAN_IN), .ZN(n2606) );
  INV_X1 U3008 ( .A(n5054), .ZN(n3750) );
  INV_X1 U3009 ( .A(n3774), .ZN(n3607) );
  INV_X1 U3010 ( .A(n4847), .ZN(n4864) );
  NAND2_X1 U3011 ( .A1(n4825), .A2(REG2_REG_10__SCAN_IN), .ZN(n4824) );
  NOR2_X1 U3012 ( .A1(n2699), .A2(n2637), .ZN(n4847) );
  NOR2_X1 U3013 ( .A1(n2699), .A2(n4755), .ZN(n4823) );
  OR2_X1 U3014 ( .A1(n4086), .A2(n3862), .ZN(n4143) );
  INV_X1 U3015 ( .A(n4941), .ZN(n4391) );
  INV_X1 U3016 ( .A(n4325), .ZN(n4365) );
  AND2_X1 U3017 ( .A1(n3807), .A2(n3824), .ZN(n3880) );
  NAND2_X1 U3018 ( .A1(n3794), .A2(n2916), .ZN(n4878) );
  NAND2_X1 U3019 ( .A1(n4397), .A2(n4983), .ZN(n5010) );
  INV_X1 U3020 ( .A(n5007), .ZN(n5020) );
  INV_X1 U3021 ( .A(n4983), .ZN(n4975) );
  INV_X1 U3022 ( .A(n2756), .ZN(n2742) );
  INV_X1 U3023 ( .A(n2720), .ZN(n3920) );
  AND2_X1 U3024 ( .A1(n2649), .A2(n2648), .ZN(n3027) );
  INV_X1 U3025 ( .A(n2606), .ZN(n3917) );
  INV_X1 U3026 ( .A(n5048), .ZN(n3753) );
  NAND2_X1 U3027 ( .A1(n3611), .A2(n3610), .ZN(n4111) );
  NAND2_X1 U3028 ( .A1(n3544), .A2(n3543), .ZN(n4209) );
  INV_X1 U3029 ( .A(n4870), .ZN(n4863) );
  INV_X1 U3030 ( .A(n4823), .ZN(n4875) );
  NAND2_X1 U3031 ( .A1(n2749), .A2(n4975), .ZN(n4950) );
  NAND2_X1 U3032 ( .A1(n5022), .A2(n5020), .ZN(n4487) );
  INV_X1 U3033 ( .A(n5022), .ZN(n5021) );
  NAND2_X1 U3034 ( .A1(n5025), .A2(n5020), .ZN(n4751) );
  INV_X1 U3035 ( .A(n5025), .ZN(n5023) );
  AND2_X2 U3036 ( .A1(n3003), .A2(n3002), .ZN(n5025) );
  INV_X2 U3037 ( .A(n4769), .ZN(n4800) );
  INV_X1 U3038 ( .A(n2918), .ZN(n4755) );
  INV_X1 U3039 ( .A(n3965), .ZN(n4970) );
  INV_X1 U3040 ( .A(n3027), .ZN(n4927) );
  NOR2_X1 U3041 ( .A1(n2715), .A2(n3917), .ZN(U4043) );
  NAND2_X1 U3042 ( .A1(n3189), .A2(n2561), .ZN(n3357) );
  INV_X1 U3043 ( .A(n3409), .ZN(n2566) );
  NAND2_X1 U3044 ( .A1(n2570), .A2(IR_REG_31__SCAN_IN), .ZN(n2577) );
  NAND2_X1 U3045 ( .A1(n2577), .A2(n2576), .ZN(n2579) );
  NAND2_X1 U3046 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2567) );
  INV_X1 U3047 ( .A(n2726), .ZN(n2573) );
  NAND2_X1 U3048 ( .A1(n2576), .A2(n2568), .ZN(n2569) );
  NAND2_X1 U3049 ( .A1(n2290), .A2(IR_REG_31__SCAN_IN), .ZN(n2571) );
  MUX2_X1 U3050 ( .A(IR_REG_31__SCAN_IN), .B(n2571), .S(IR_REG_25__SCAN_IN), 
        .Z(n2572) );
  NAND2_X1 U3051 ( .A1(n2572), .A2(n2264), .ZN(n2738) );
  NAND2_X1 U3052 ( .A1(n2264), .A2(IR_REG_31__SCAN_IN), .ZN(n2574) );
  OR2_X1 U3053 ( .A1(n2577), .A2(n2576), .ZN(n2578) );
  INV_X2 U3054 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3055 ( .A(DATAI_21_), .ZN(n4535) );
  NAND2_X1 U3056 ( .A1(n2580), .A2(IR_REG_31__SCAN_IN), .ZN(n2581) );
  NAND2_X1 U3057 ( .A1(n3797), .A2(STATE_REG_SCAN_IN), .ZN(n2582) );
  OAI21_X1 U3058 ( .B1(STATE_REG_SCAN_IN), .B2(n4535), .A(n2582), .ZN(U3331)
         );
  INV_X1 U3059 ( .A(DATAI_17_), .ZN(n4636) );
  NAND2_X1 U3060 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U3061 ( .A1(n3368), .A2(n2583), .ZN(n3392) );
  INV_X1 U3062 ( .A(IR_REG_17__SCAN_IN), .ZN(n2585) );
  XNOR2_X1 U3063 ( .A(n2596), .B(n2585), .ZN(n4020) );
  NAND2_X1 U3064 ( .A1(n4020), .A2(STATE_REG_SCAN_IN), .ZN(n2586) );
  OAI21_X1 U3065 ( .B1(STATE_REG_SCAN_IN), .B2(n4636), .A(n2586), .ZN(U3335)
         );
  INV_X1 U3066 ( .A(DATAI_22_), .ZN(n4519) );
  INV_X1 U3067 ( .A(n2587), .ZN(n2588) );
  NAND2_X1 U3068 ( .A1(n2588), .A2(IR_REG_31__SCAN_IN), .ZN(n2590) );
  NAND2_X1 U3069 ( .A1(n3920), .A2(STATE_REG_SCAN_IN), .ZN(n2591) );
  OAI21_X1 U3070 ( .B1(STATE_REG_SCAN_IN), .B2(n4519), .A(n2591), .ZN(U3330)
         );
  NAND2_X1 U3071 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2592) );
  OAI21_X1 U3072 ( .B1(n2738), .B2(U3149), .A(n2592), .ZN(U3327) );
  INV_X1 U3073 ( .A(DATAI_24_), .ZN(n4626) );
  NAND2_X1 U3074 ( .A1(n2726), .A2(STATE_REG_SCAN_IN), .ZN(n2593) );
  OAI21_X1 U3075 ( .B1(STATE_REG_SCAN_IN), .B2(n4626), .A(n2593), .ZN(U3328)
         );
  INV_X1 U3076 ( .A(DATAI_26_), .ZN(n4620) );
  NAND2_X1 U3077 ( .A1(n2737), .A2(STATE_REG_SCAN_IN), .ZN(n2594) );
  OAI21_X1 U3078 ( .B1(STATE_REG_SCAN_IN), .B2(n4620), .A(n2594), .ZN(U3326)
         );
  INV_X1 U3079 ( .A(DATAI_20_), .ZN(n4631) );
  NAND2_X1 U3080 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U3081 ( .A1(n2262), .A2(STATE_REG_SCAN_IN), .ZN(n2598) );
  OAI21_X1 U3082 ( .B1(STATE_REG_SCAN_IN), .B2(n4631), .A(n2598), .ZN(U3332)
         );
  INV_X1 U3083 ( .A(DATAI_29_), .ZN(n4614) );
  NAND2_X1 U3084 ( .A1(n2601), .A2(IR_REG_31__SCAN_IN), .ZN(n2600) );
  INV_X1 U3085 ( .A(n2704), .ZN(n3353) );
  NAND2_X1 U3086 ( .A1(n2707), .A2(STATE_REG_SCAN_IN), .ZN(n2603) );
  OAI21_X1 U3087 ( .B1(STATE_REG_SCAN_IN), .B2(n4614), .A(n2603), .ZN(U3323)
         );
  NAND2_X1 U3088 ( .A1(n2738), .A2(B_REG_SCAN_IN), .ZN(n2604) );
  MUX2_X1 U3089 ( .A(n2604), .B(B_REG_SCAN_IN), .S(n2726), .Z(n2605) );
  INV_X1 U3090 ( .A(D_REG_0__SCAN_IN), .ZN(n2608) );
  NOR3_X1 U3091 ( .A1(n2737), .A2(n3917), .A3(n2726), .ZN(n2607) );
  AOI21_X1 U3092 ( .B1(n4769), .B2(n2608), .A(n2607), .ZN(U3458) );
  INV_X1 U3093 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2610) );
  AND2_X1 U3094 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2611)
         );
  NAND2_X1 U3095 ( .A1(n2612), .A2(n2611), .ZN(n3936) );
  NAND2_X1 U3096 ( .A1(n4766), .A2(REG1_REG_1__SCAN_IN), .ZN(n2613) );
  INV_X1 U3097 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3001) );
  MUX2_X1 U3098 ( .A(n3001), .B(REG1_REG_2__SCAN_IN), .S(n4765), .Z(n2828) );
  INV_X1 U3099 ( .A(IR_REG_2__SCAN_IN), .ZN(n2614) );
  AND2_X1 U3100 ( .A1(n2615), .A2(n2614), .ZN(n2643) );
  NOR2_X1 U3101 ( .A1(n2643), .A2(n3190), .ZN(n2616) );
  NAND2_X1 U3102 ( .A1(n2616), .A2(IR_REG_3__SCAN_IN), .ZN(n2619) );
  INV_X1 U3103 ( .A(n2616), .ZN(n2618) );
  NAND2_X1 U3104 ( .A1(n2618), .A2(n2617), .ZN(n2651) );
  XNOR2_X1 U3105 ( .A(n2650), .B(REG1_REG_3__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3106 ( .A1(n2620), .A2(STATE_REG_SCAN_IN), .ZN(n4767) );
  NAND2_X1 U3107 ( .A1(n2622), .A2(IR_REG_27__SCAN_IN), .ZN(n2623) );
  NAND2_X1 U3108 ( .A1(n2625), .A2(n2917), .ZN(n2626) );
  NAND2_X1 U3109 ( .A1(n2261), .A2(n2626), .ZN(n2628) );
  OR2_X1 U3110 ( .A1(n2629), .A2(n2628), .ZN(n2699) );
  XNOR2_X1 U3111 ( .A(n2627), .B(n2316), .ZN(n4756) );
  NOR2_X2 U3112 ( .A1(n2699), .A2(n4756), .ZN(n4870) );
  INV_X1 U3113 ( .A(n2628), .ZN(n2630) );
  INV_X1 U3114 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4567) );
  NOR2_X1 U3115 ( .A1(STATE_REG_SCAN_IN), .A2(n4567), .ZN(n2860) );
  NAND2_X1 U3116 ( .A1(n2303), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  MUX2_X1 U3117 ( .A(IR_REG_31__SCAN_IN), .B(n2631), .S(IR_REG_28__SCAN_IN), 
        .Z(n2632) );
  NAND2_X1 U3118 ( .A1(n2632), .A2(n2601), .ZN(n2918) );
  NOR2_X1 U3119 ( .A1(n4875), .A2(n2478), .ZN(n2633) );
  AOI211_X1 U3120 ( .C1(n4869), .C2(ADDR_REG_3__SCAN_IN), .A(n2860), .B(n2633), 
        .ZN(n2640) );
  INV_X1 U3121 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2774) );
  XNOR2_X1 U3122 ( .A(n4765), .B(n2774), .ZN(n2831) );
  INV_X1 U3123 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2954) );
  NAND2_X1 U3124 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2815) );
  INV_X1 U3125 ( .A(n2815), .ZN(n3938) );
  NAND2_X1 U3126 ( .A1(n4766), .A2(REG2_REG_1__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U3127 ( .A1(n3937), .A2(n2634), .ZN(n2830) );
  NAND2_X1 U3128 ( .A1(n4765), .A2(REG2_REG_2__SCAN_IN), .ZN(n2635) );
  NAND2_X1 U3129 ( .A1(n2636), .A2(n2635), .ZN(n2675) );
  XNOR2_X1 U3130 ( .A(n2675), .B(n2478), .ZN(n2638) );
  NAND2_X1 U3131 ( .A1(n4755), .A2(n4756), .ZN(n2637) );
  NAND2_X1 U3132 ( .A1(n2638), .A2(REG2_REG_3__SCAN_IN), .ZN(n2677) );
  OAI211_X1 U3133 ( .C1(REG2_REG_3__SCAN_IN), .C2(n2638), .A(n4847), .B(n2677), 
        .ZN(n2639) );
  OAI211_X1 U3134 ( .C1(n2641), .C2(n4863), .A(n2640), .B(n2639), .ZN(U3243)
         );
  NOR2_X1 U3135 ( .A1(n4869), .A2(U4043), .ZN(U3148) );
  NOR2_X1 U3136 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2642)
         );
  NAND2_X1 U3137 ( .A1(n2656), .A2(n4599), .ZN(n2658) );
  INV_X1 U3138 ( .A(n2665), .ZN(n2644) );
  NAND2_X1 U3139 ( .A1(n2644), .A2(n4717), .ZN(n2666) );
  NAND2_X1 U3140 ( .A1(n2666), .A2(IR_REG_31__SCAN_IN), .ZN(n2645) );
  XNOR2_X1 U3141 ( .A(n2645), .B(IR_REG_8__SCAN_IN), .ZN(n4760) );
  NOR2_X1 U3142 ( .A1(STATE_REG_SCAN_IN), .A2(n4573), .ZN(n3143) );
  AOI21_X1 U3143 ( .B1(n4869), .B2(ADDR_REG_8__SCAN_IN), .A(n3143), .ZN(n2646)
         );
  INV_X1 U3144 ( .A(n2646), .ZN(n2674) );
  INV_X1 U3145 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2672) );
  NAND2_X1 U3146 ( .A1(n2658), .A2(IR_REG_31__SCAN_IN), .ZN(n2647) );
  MUX2_X1 U3147 ( .A(IR_REG_31__SCAN_IN), .B(n2647), .S(IR_REG_6__SCAN_IN), 
        .Z(n2649) );
  NAND2_X1 U31480 ( .A1(n2651), .A2(IR_REG_31__SCAN_IN), .ZN(n2652) );
  XNOR2_X1 U31490 ( .A(n2652), .B(IR_REG_4__SCAN_IN), .ZN(n4763) );
  XNOR2_X1 U3150 ( .A(n2654), .B(n4763), .ZN(n2812) );
  INV_X1 U3151 ( .A(n2812), .ZN(n2655) );
  INV_X1 U3152 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4917) );
  INV_X1 U3153 ( .A(n4763), .ZN(n2653) );
  INV_X1 U3154 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2661) );
  NOR2_X1 U3155 ( .A1(n2656), .A2(n3190), .ZN(n2657) );
  MUX2_X1 U3156 ( .A(n3190), .B(n2657), .S(IR_REG_5__SCAN_IN), .Z(n2660) );
  INV_X1 U3157 ( .A(n2658), .ZN(n2659) );
  MUX2_X1 U3158 ( .A(REG1_REG_5__SCAN_IN), .B(n2661), .S(n4762), .Z(n2693) );
  NAND2_X1 U3159 ( .A1(n4762), .A2(REG1_REG_5__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3160 ( .A1(n3027), .A2(n2663), .ZN(n2664) );
  NAND2_X1 U3161 ( .A1(n2665), .A2(IR_REG_7__SCAN_IN), .ZN(n2667) );
  AND2_X1 U3162 ( .A1(n4761), .A2(REG1_REG_7__SCAN_IN), .ZN(n2766) );
  INV_X1 U3163 ( .A(n4760), .ZN(n2668) );
  AOI211_X1 U3164 ( .C1(n2672), .C2(n2671), .A(n3961), .B(n4863), .ZN(n2673)
         );
  AOI211_X1 U3165 ( .C1(n4823), .C2(n4760), .A(n2674), .B(n2673), .ZN(n2686)
         );
  NAND2_X1 U3166 ( .A1(n2675), .A2(n4764), .ZN(n2676) );
  NAND2_X1 U3167 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  XNOR2_X1 U3168 ( .A(n2678), .B(n4763), .ZN(n2820) );
  INV_X1 U3169 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2821) );
  NOR2_X1 U3170 ( .A1(n2820), .A2(n2821), .ZN(n2819) );
  XNOR2_X1 U3171 ( .A(n4762), .B(REG2_REG_5__SCAN_IN), .ZN(n2688) );
  INV_X1 U3172 ( .A(REG2_REG_6__SCAN_IN), .ZN(n4803) );
  INV_X1 U3173 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2681) );
  XNOR2_X1 U3174 ( .A(n3947), .B(n4760), .ZN(n2684) );
  OAI211_X1 U3175 ( .C1(n2684), .C2(REG2_REG_8__SCAN_IN), .A(n4847), .B(n3949), 
        .ZN(n2685) );
  NAND2_X1 U3176 ( .A1(n2686), .A2(n2685), .ZN(U3248) );
  INV_X1 U3177 ( .A(n4762), .ZN(n2696) );
  AND2_X1 U3178 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n2902) );
  AOI211_X1 U3179 ( .C1(n2689), .C2(n2688), .A(n2687), .B(n4864), .ZN(n2690)
         );
  AOI211_X1 U3180 ( .C1(n4869), .C2(ADDR_REG_5__SCAN_IN), .A(n2902), .B(n2690), 
        .ZN(n2695) );
  OAI211_X1 U3181 ( .C1(n2693), .C2(n2692), .A(n4870), .B(n2691), .ZN(n2694)
         );
  OAI211_X1 U3182 ( .C1(n4875), .C2(n2696), .A(n2695), .B(n2694), .ZN(U3245)
         );
  INV_X1 U3183 ( .A(IR_REG_0__SCAN_IN), .ZN(n3934) );
  OAI21_X1 U3184 ( .B1(n4756), .B2(REG1_REG_0__SCAN_IN), .A(n3934), .ZN(n2697)
         );
  INV_X1 U3185 ( .A(n4756), .ZN(n3918) );
  INV_X1 U3186 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4889) );
  OAI21_X1 U3187 ( .B1(n3918), .B2(REG2_REG_0__SCAN_IN), .A(n4755), .ZN(n2817)
         );
  MUX2_X1 U3188 ( .A(n2697), .B(n3934), .S(n2817), .Z(n2700) );
  INV_X1 U3189 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2698) );
  OAI22_X1 U3190 ( .A1(n2700), .A2(n2699), .B1(STATE_REG_SCAN_IN), .B2(n2698), 
        .ZN(n2701) );
  AOI21_X1 U3191 ( .B1(n4869), .B2(ADDR_REG_0__SCAN_IN), .A(n2701), .ZN(n2703)
         );
  INV_X1 U3192 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4881) );
  NAND3_X1 U3193 ( .A1(n4870), .A2(IR_REG_0__SCAN_IN), .A3(n4881), .ZN(n2702)
         );
  NAND2_X1 U3194 ( .A1(n2703), .A2(n2702), .ZN(U3240) );
  NAND2_X1 U3195 ( .A1(n3774), .A2(REG0_REG_0__SCAN_IN), .ZN(n2712) );
  INV_X1 U3196 ( .A(n2706), .ZN(n4754) );
  AND2_X2 U3197 ( .A1(n4754), .A2(n2707), .ZN(n2797) );
  NAND2_X1 U3198 ( .A1(n2797), .A2(REG3_REG_0__SCAN_IN), .ZN(n2711) );
  AND2_X2 U3199 ( .A1(n2706), .A2(n2707), .ZN(n2800) );
  NAND2_X1 U3200 ( .A1(n2800), .A2(REG1_REG_0__SCAN_IN), .ZN(n2710) );
  NAND2_X2 U3201 ( .A1(n4754), .A2(n2708), .ZN(n2802) );
  AND2_X4 U3202 ( .A1(n2757), .A2(n2715), .ZN(n3477) );
  NAND2_X1 U3203 ( .A1(n2907), .A2(n3477), .ZN(n2717) );
  AND2_X4 U3204 ( .A1(n2715), .A2(n2928), .ZN(n2786) );
  NAND2_X1 U3205 ( .A1(n3795), .A2(n2786), .ZN(n2716) );
  INV_X1 U3206 ( .A(n2715), .ZN(n2721) );
  NAND2_X1 U3207 ( .A1(n2721), .A2(REG1_REG_0__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3208 ( .A1(n2782), .A2(n2718), .ZN(n2725) );
  NAND2_X2 U3209 ( .A1(n2786), .A2(n5007), .ZN(n3595) );
  NAND2_X1 U32100 ( .A1(n2907), .A2(n3548), .ZN(n2723) );
  AOI22_X1 U32110 ( .A1(n3795), .A2(n3477), .B1(n2721), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2722) );
  NAND2_X1 U32120 ( .A1(n2723), .A2(n2722), .ZN(n2724) );
  OAI21_X1 U32130 ( .B1(n2725), .B2(n2724), .A(n2784), .ZN(n2813) );
  INV_X1 U32140 ( .A(n3002), .ZN(n2984) );
  NOR4_X1 U32150 ( .A1(D_REG_27__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_25__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2735) );
  NOR4_X1 U32160 ( .A1(D_REG_23__SCAN_IN), .A2(D_REG_22__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_20__SCAN_IN), .ZN(n2734) );
  INV_X1 U32170 ( .A(D_REG_31__SCAN_IN), .ZN(n4799) );
  INV_X1 U32180 ( .A(D_REG_30__SCAN_IN), .ZN(n4798) );
  INV_X1 U32190 ( .A(D_REG_29__SCAN_IN), .ZN(n4797) );
  INV_X1 U32200 ( .A(D_REG_28__SCAN_IN), .ZN(n4796) );
  NAND4_X1 U32210 ( .A1(n4799), .A2(n4798), .A3(n4797), .A4(n4796), .ZN(n2732)
         );
  NOR4_X1 U32220 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n2730) );
  NOR4_X1 U32230 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2729) );
  NOR4_X1 U32240 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_6__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n2728) );
  NOR4_X1 U32250 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2727) );
  NAND4_X1 U32260 ( .A1(n2730), .A2(n2729), .A3(n2728), .A4(n2727), .ZN(n2731)
         );
  NOR4_X1 U32270 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(n2732), 
        .A4(n2731), .ZN(n2733) );
  AND3_X1 U32280 ( .A1(n2735), .A2(n2734), .A3(n2733), .ZN(n2736) );
  NOR2_X1 U32290 ( .A1(n2740), .A2(n2736), .ZN(n2924) );
  INV_X1 U32300 ( .A(n2737), .ZN(n2739) );
  NAND2_X1 U32310 ( .A1(n2739), .A2(n2738), .ZN(n4753) );
  OAI21_X1 U32320 ( .B1(n2740), .B2(D_REG_1__SCAN_IN), .A(n4753), .ZN(n2981)
         );
  NOR2_X1 U32330 ( .A1(n2924), .A2(n2981), .ZN(n2741) );
  NAND2_X1 U32340 ( .A1(n2984), .A2(n2741), .ZN(n2753) );
  INV_X1 U32350 ( .A(n2753), .ZN(n2743) );
  XNOR2_X1 U32360 ( .A(n2745), .B(n2744), .ZN(n2748) );
  AOI21_X1 U32370 ( .B1(n4936), .B2(n4876), .A(n2917), .ZN(n2746) );
  AND2_X1 U32380 ( .A1(n4939), .A2(n2746), .ZN(n2751) );
  INV_X1 U32390 ( .A(n2758), .ZN(n2747) );
  OR2_X1 U32400 ( .A1(n2747), .A2(n4939), .ZN(n2750) );
  NOR2_X1 U32410 ( .A1(n2756), .A2(n3797), .ZN(n2749) );
  NAND2_X1 U32420 ( .A1(n2753), .A2(n2751), .ZN(n2854) );
  OAI22_X1 U32430 ( .A1(n2756), .A2(n2928), .B1(n4939), .B2(U3149), .ZN(n2752)
         );
  NAND2_X1 U32440 ( .A1(n2753), .A2(n2752), .ZN(n2856) );
  NAND2_X1 U32450 ( .A1(n2719), .A2(n4034), .ZN(n2754) );
  NAND2_X1 U32460 ( .A1(n2754), .A2(n2917), .ZN(n2853) );
  INV_X1 U32470 ( .A(n2853), .ZN(n2755) );
  INV_X1 U32480 ( .A(n2980), .ZN(n2925) );
  NAND3_X1 U32490 ( .A1(n2854), .A2(n2856), .A3(n2925), .ZN(n3655) );
  AOI22_X1 U32500 ( .A1(n5050), .A2(n3795), .B1(n3655), .B2(
        REG3_REG_0__SCAN_IN), .ZN(n2764) );
  NAND2_X1 U32510 ( .A1(n2758), .A2(n2757), .ZN(n2808) );
  NAND2_X1 U32520 ( .A1(n3774), .A2(REG0_REG_1__SCAN_IN), .ZN(n2762) );
  NAND2_X1 U32530 ( .A1(n2800), .A2(REG1_REG_1__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U32540 ( .A1(n5040), .A2(n2906), .ZN(n2763) );
  OAI211_X1 U32550 ( .C1(n2813), .C2(n3753), .A(n2764), .B(n2763), .ZN(U3229)
         );
  MUX2_X1 U32560 ( .A(n2681), .B(REG2_REG_7__SCAN_IN), .S(n4761), .Z(n2765) );
  AOI21_X1 U32570 ( .B1(n2495), .B2(n2496), .A(n2766), .ZN(n2768) );
  AOI21_X1 U32580 ( .B1(n2768), .B2(n2769), .A(n4863), .ZN(n2767) );
  OAI21_X1 U32590 ( .B1(n2769), .B2(n2768), .A(n2767), .ZN(n2771) );
  INV_X1 U32600 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4665) );
  NOR2_X1 U32610 ( .A1(STATE_REG_SCAN_IN), .A2(n4665), .ZN(n3621) );
  AOI21_X1 U32620 ( .B1(n4869), .B2(ADDR_REG_7__SCAN_IN), .A(n3621), .ZN(n2770) );
  OAI211_X1 U32630 ( .C1(n4875), .C2(n2496), .A(n2771), .B(n2770), .ZN(n2772)
         );
  OR2_X1 U32640 ( .A1(n2773), .A2(n2772), .ZN(U3247) );
  MUX2_X1 U32650 ( .A(n4765), .B(DATAI_2_), .S(n2261), .Z(n2995) );
  NAND2_X1 U32660 ( .A1(n2995), .A2(n2786), .ZN(n2780) );
  NAND2_X1 U32670 ( .A1(n3774), .A2(REG0_REG_2__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U32680 ( .A1(n2797), .A2(REG3_REG_2__SCAN_IN), .ZN(n2777) );
  NAND2_X1 U32690 ( .A1(n2800), .A2(REG1_REG_2__SCAN_IN), .ZN(n2776) );
  NAND2_X1 U32700 ( .A1(n3931), .A2(n3477), .ZN(n2779) );
  NAND2_X1 U32710 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  NAND2_X4 U32720 ( .A1(n2928), .A2(n2806), .ZN(n3596) );
  XNOR2_X1 U32730 ( .A(n2781), .B(n3566), .ZN(n2845) );
  AOI22_X1 U32740 ( .A1(n3931), .A2(n3548), .B1(n3477), .B2(n2995), .ZN(n2844)
         );
  XNOR2_X1 U32750 ( .A(n2845), .B(n2844), .ZN(n2796) );
  NAND2_X1 U32760 ( .A1(n2782), .A2(n3566), .ZN(n2783) );
  NAND2_X1 U32770 ( .A1(n2784), .A2(n2783), .ZN(n3653) );
  NAND2_X1 U32780 ( .A1(n2906), .A2(n3477), .ZN(n2788) );
  NAND2_X1 U32790 ( .A1(n3653), .A2(n3654), .ZN(n3652) );
  INV_X1 U32800 ( .A(n2791), .ZN(n2792) );
  NAND2_X1 U32810 ( .A1(n2790), .A2(n2792), .ZN(n2793) );
  NAND2_X1 U32820 ( .A1(n3652), .A2(n2793), .ZN(n2795) );
  INV_X1 U32830 ( .A(n2847), .ZN(n2794) );
  AOI21_X1 U32840 ( .B1(n2796), .B2(n2795), .A(n2794), .ZN(n2811) );
  AOI22_X1 U32850 ( .A1(n5050), .A2(n2995), .B1(n3655), .B2(
        REG3_REG_2__SCAN_IN), .ZN(n2810) );
  INV_X2 U32860 ( .A(n5032), .ZN(n5040) );
  NAND2_X1 U32870 ( .A1(n2797), .A2(n4567), .ZN(n2799) );
  NAND2_X1 U32880 ( .A1(n3774), .A2(REG0_REG_3__SCAN_IN), .ZN(n2798) );
  NAND2_X1 U32890 ( .A1(n2799), .A2(n2798), .ZN(n2801) );
  NOR2_X1 U32900 ( .A1(n2801), .A2(n2554), .ZN(n2805) );
  INV_X1 U32910 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2803) );
  OR2_X1 U32920 ( .A1(n2802), .A2(n2803), .ZN(n2804) );
  INV_X1 U32930 ( .A(n2806), .ZN(n2807) );
  NAND2_X1 U32940 ( .A1(n4755), .A2(n2807), .ZN(n3919) );
  INV_X2 U32950 ( .A(n4991), .ZN(n5045) );
  AOI22_X1 U32960 ( .A1(n5040), .A2(n2843), .B1(n5045), .B2(n2906), .ZN(n2809)
         );
  OAI211_X1 U32970 ( .C1(n2811), .C2(n3753), .A(n2810), .B(n2809), .ZN(U3234)
         );
  XOR2_X1 U32980 ( .A(n4917), .B(n2812), .Z(n2826) );
  NOR2_X1 U32990 ( .A1(n2813), .A2(n4756), .ZN(n2814) );
  AOI211_X1 U33000 ( .C1(n4756), .C2(n2815), .A(n2918), .B(n2814), .ZN(n2816)
         );
  AOI211_X1 U33010 ( .C1(n3934), .C2(n2817), .A(n3932), .B(n2816), .ZN(n2839)
         );
  INV_X1 U33020 ( .A(n2839), .ZN(n2825) );
  AND2_X1 U33030 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n2938) );
  AOI21_X1 U33040 ( .B1(n4869), .B2(ADDR_REG_4__SCAN_IN), .A(n2938), .ZN(n2818) );
  INV_X1 U33050 ( .A(n2818), .ZN(n2823) );
  AOI211_X1 U33060 ( .C1(n2821), .C2(n2820), .A(n2819), .B(n4864), .ZN(n2822)
         );
  AOI211_X1 U33070 ( .C1(n4823), .C2(n4763), .A(n2823), .B(n2822), .ZN(n2824)
         );
  OAI211_X1 U33080 ( .C1(n4863), .C2(n2826), .A(n2825), .B(n2824), .ZN(U3244)
         );
  AOI211_X1 U33090 ( .C1(n2829), .C2(n2828), .A(n2827), .B(n4863), .ZN(n2838)
         );
  INV_X1 U33100 ( .A(n2830), .ZN(n2833) );
  INV_X1 U33110 ( .A(n2831), .ZN(n2832) );
  INV_X1 U33120 ( .A(n4765), .ZN(n2835) );
  AOI22_X1 U33130 ( .A1(n4869), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2834) );
  OAI21_X1 U33140 ( .B1(n4875), .B2(n2835), .A(n2834), .ZN(n2836) );
  OR4_X1 U33150 ( .A1(n2839), .A2(n2838), .A3(n2837), .A4(n2836), .ZN(U3242)
         );
  NAND2_X1 U33160 ( .A1(n2843), .A2(n3477), .ZN(n2841) );
  MUX2_X1 U33170 ( .A(n4764), .B(DATAI_3_), .S(n2261), .Z(n2959) );
  NAND2_X1 U33180 ( .A1(n2959), .A2(n2786), .ZN(n2840) );
  NAND2_X1 U33190 ( .A1(n2841), .A2(n2840), .ZN(n2842) );
  AOI22_X1 U33200 ( .A1(n2843), .A2(n3548), .B1(n3477), .B2(n2959), .ZN(n2867)
         );
  XNOR2_X1 U33210 ( .A(n2866), .B(n2867), .ZN(n2864) );
  NAND2_X1 U33220 ( .A1(n2845), .A2(n2844), .ZN(n2846) );
  XOR2_X1 U33230 ( .A(n2864), .B(n2865), .Z(n2863) );
  NAND2_X1 U33240 ( .A1(n3774), .A2(REG0_REG_4__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U33250 ( .A1(n2800), .A2(REG1_REG_4__SCAN_IN), .ZN(n2851) );
  INV_X1 U33260 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2848) );
  XNOR2_X1 U33270 ( .A(n2848), .B(REG3_REG_3__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U33280 ( .A1(n2797), .A2(n3020), .ZN(n2850) );
  OR2_X1 U33290 ( .A1(n2802), .A2(n2821), .ZN(n2849) );
  AOI22_X1 U33300 ( .A1(n5040), .A2(n3930), .B1(n5045), .B2(n3931), .ZN(n2862)
         );
  NAND3_X1 U33310 ( .A1(n2854), .A2(n2715), .A3(n2853), .ZN(n2855) );
  NAND2_X1 U33320 ( .A1(n2855), .A2(STATE_REG_SCAN_IN), .ZN(n2858) );
  AND2_X1 U33330 ( .A1(n2856), .A2(n4767), .ZN(n2857) );
  NOR2_X1 U33340 ( .A1(n3748), .A2(n2962), .ZN(n2859) );
  AOI211_X1 U33350 ( .C1(n4567), .C2(n3750), .A(n2860), .B(n2859), .ZN(n2861)
         );
  OAI211_X1 U33360 ( .C1(n2863), .C2(n3753), .A(n2862), .B(n2861), .ZN(U3215)
         );
  INV_X1 U33370 ( .A(n2866), .ZN(n2868) );
  NAND2_X1 U33380 ( .A1(n2868), .A2(n2867), .ZN(n2869) );
  NAND2_X1 U33390 ( .A1(n2870), .A2(n2869), .ZN(n2934) );
  INV_X1 U33400 ( .A(n2934), .ZN(n2875) );
  NAND2_X1 U33410 ( .A1(n3930), .A2(n3477), .ZN(n2872) );
  MUX2_X1 U33420 ( .A(n4763), .B(DATAI_4_), .S(n2261), .Z(n3019) );
  NAND2_X1 U33430 ( .A1(n3019), .A2(n2786), .ZN(n2871) );
  NAND2_X1 U33440 ( .A1(n2872), .A2(n2871), .ZN(n2873) );
  XNOR2_X1 U33450 ( .A(n2873), .B(n3566), .ZN(n2876) );
  AOI22_X1 U33460 ( .A1(n3930), .A2(n3548), .B1(n3477), .B2(n3019), .ZN(n2877)
         );
  XNOR2_X1 U33470 ( .A(n2876), .B(n2877), .ZN(n2937) );
  INV_X1 U33480 ( .A(n2937), .ZN(n2874) );
  INV_X1 U33490 ( .A(n2876), .ZN(n2879) );
  INV_X1 U33500 ( .A(n2877), .ZN(n2878) );
  NAND2_X1 U33510 ( .A1(n2879), .A2(n2878), .ZN(n2880) );
  NAND2_X1 U33520 ( .A1(n3774), .A2(REG0_REG_5__SCAN_IN), .ZN(n2888) );
  NAND2_X1 U3353 ( .A1(n2800), .A2(REG1_REG_5__SCAN_IN), .ZN(n2887) );
  INV_X1 U33540 ( .A(n2883), .ZN(n2882) );
  INV_X1 U3355 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2881) );
  NAND2_X1 U3356 ( .A1(n2882), .A2(n2881), .ZN(n2884) );
  NAND2_X1 U3357 ( .A1(n2883), .A2(REG3_REG_5__SCAN_IN), .ZN(n2895) );
  AND2_X1 U3358 ( .A1(n2884), .A2(n2895), .ZN(n2967) );
  NAND2_X1 U3359 ( .A1(n2797), .A2(n2967), .ZN(n2886) );
  INV_X1 U3360 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2969) );
  OR2_X1 U3361 ( .A1(n2802), .A2(n2969), .ZN(n2885) );
  NAND4_X1 U3362 ( .A1(n2888), .A2(n2887), .A3(n2886), .A4(n2885), .ZN(n3929)
         );
  NAND2_X1 U3363 ( .A1(n3929), .A2(n3548), .ZN(n2890) );
  MUX2_X1 U3364 ( .A(n4762), .B(DATAI_5_), .S(n2261), .Z(n3055) );
  NAND2_X1 U3365 ( .A1(n3055), .A2(n3477), .ZN(n2889) );
  NAND2_X1 U3366 ( .A1(n2890), .A2(n2889), .ZN(n3025) );
  NAND2_X1 U3367 ( .A1(n3929), .A2(n3477), .ZN(n2892) );
  NAND2_X1 U3368 ( .A1(n3055), .A2(n2786), .ZN(n2891) );
  NAND2_X1 U3369 ( .A1(n2892), .A2(n2891), .ZN(n2893) );
  XNOR2_X1 U3370 ( .A(n2893), .B(n3596), .ZN(n3024) );
  XOR2_X1 U3371 ( .A(n3025), .B(n3024), .Z(n2894) );
  XNOR2_X1 U3372 ( .A(n3026), .B(n2894), .ZN(n2905) );
  NAND2_X1 U3373 ( .A1(n3774), .A2(REG0_REG_6__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U3374 ( .A1(n2800), .A2(REG1_REG_6__SCAN_IN), .ZN(n2899) );
  AND2_X1 U3375 ( .A1(n2895), .A2(n3045), .ZN(n2896) );
  NOR2_X1 U3376 ( .A1(n3039), .A2(n2896), .ZN(n3038) );
  NAND2_X1 U3377 ( .A1(n2797), .A2(n3038), .ZN(n2898) );
  OR2_X1 U3378 ( .A1(n2802), .A2(n4803), .ZN(n2897) );
  NAND4_X1 U3379 ( .A1(n2900), .A2(n2899), .A3(n2898), .A4(n2897), .ZN(n3928)
         );
  AOI22_X1 U3380 ( .A1(n5040), .A2(n3928), .B1(n5045), .B2(n3930), .ZN(n2904)
         );
  INV_X1 U3381 ( .A(n3055), .ZN(n3051) );
  NOR2_X1 U3382 ( .A1(n3748), .A2(n3051), .ZN(n2901) );
  AOI211_X1 U3383 ( .C1(n2967), .C2(n3750), .A(n2902), .B(n2901), .ZN(n2903)
         );
  OAI211_X1 U3384 ( .C1(n2905), .C2(n3753), .A(n2904), .B(n2903), .ZN(U3224)
         );
  INV_X1 U3385 ( .A(n2906), .ZN(n2990) );
  NAND2_X1 U3386 ( .A1(n2990), .A2(n3656), .ZN(n2912) );
  INV_X1 U3387 ( .A(n3656), .ZN(n2947) );
  AND2_X1 U3388 ( .A1(n2907), .A2(n3795), .ZN(n2946) );
  NAND2_X1 U3389 ( .A1(n2906), .A2(n3656), .ZN(n2908) );
  INV_X1 U3390 ( .A(n2995), .ZN(n2909) );
  NAND2_X1 U3391 ( .A1(n3931), .A2(n2909), .ZN(n3802) );
  NAND2_X1 U3392 ( .A1(n2920), .A2(n2909), .ZN(n2910) );
  NAND2_X1 U3393 ( .A1(n2985), .A2(n2910), .ZN(n2961) );
  NAND2_X1 U3394 ( .A1(n2963), .A2(n2959), .ZN(n3804) );
  NAND2_X1 U3395 ( .A1(n2843), .A2(n2962), .ZN(n3801) );
  XNOR2_X1 U3396 ( .A(n2961), .B(n3892), .ZN(n4906) );
  XNOR2_X1 U3397 ( .A(n2928), .B(n3920), .ZN(n2911) );
  INV_X1 U3398 ( .A(n2907), .ZN(n2948) );
  NAND2_X1 U3399 ( .A1(n2948), .A2(n3795), .ZN(n3867) );
  NAND2_X1 U3400 ( .A1(n2989), .A2(n3884), .ZN(n2988) );
  NAND2_X1 U3401 ( .A1(n2988), .A2(n3799), .ZN(n2915) );
  NAND2_X1 U3402 ( .A1(n2915), .A2(n3892), .ZN(n2971) );
  OAI21_X1 U3403 ( .B1(n3892), .B2(n2915), .A(n2971), .ZN(n2922) );
  NAND2_X1 U3404 ( .A1(n2262), .A2(n3797), .ZN(n3794) );
  NAND2_X1 U3405 ( .A1(n4936), .A2(n3920), .ZN(n2916) );
  AOI22_X1 U3406 ( .A1(n3930), .A2(n4944), .B1(n4417), .B2(n2959), .ZN(n2919)
         );
  OAI21_X1 U3407 ( .B1(n2920), .B2(n4941), .A(n2919), .ZN(n2921) );
  AOI21_X1 U3408 ( .B1(n2922), .B2(n4878), .A(n2921), .ZN(n2923) );
  OAI21_X1 U3409 ( .B1(n4906), .B2(n4397), .A(n2923), .ZN(n4908) );
  INV_X1 U3410 ( .A(n4908), .ZN(n2933) );
  INV_X1 U3411 ( .A(n2981), .ZN(n2926) );
  INV_X1 U3412 ( .A(n2924), .ZN(n2983) );
  NAND4_X1 U3413 ( .A1(n2926), .A2(n2925), .A3(n2983), .A4(n3002), .ZN(n2927)
         );
  INV_X1 U3414 ( .A(n4906), .ZN(n2931) );
  NOR2_X1 U3415 ( .A1(n2928), .A2(n4034), .ZN(n4933) );
  NAND2_X1 U3416 ( .A1(n2260), .A2(n4933), .ZN(n4406) );
  INV_X1 U3417 ( .A(n4406), .ZN(n4900) );
  NAND2_X1 U3418 ( .A1(n2998), .A2(n2962), .ZN(n3018) );
  OAI21_X1 U3419 ( .B1(n2998), .B2(n2962), .A(n3018), .ZN(n4905) );
  NAND2_X1 U3420 ( .A1(n2260), .A2(n4034), .ZN(n4305) );
  OR2_X1 U3421 ( .A1(n4305), .A2(n5007), .ZN(n4338) );
  AOI22_X1 U3422 ( .A1(n5058), .A2(REG2_REG_3__SCAN_IN), .B1(n4897), .B2(n4567), .ZN(n2929) );
  OAI21_X1 U3423 ( .B1(n4905), .B2(n4338), .A(n2929), .ZN(n2930) );
  AOI21_X1 U3424 ( .B1(n2931), .B2(n4900), .A(n2930), .ZN(n2932) );
  OAI21_X1 U3425 ( .B1(n2933), .B2(n5058), .A(n2932), .ZN(U3287) );
  INV_X1 U3426 ( .A(n2935), .ZN(n2936) );
  AOI211_X1 U3427 ( .C1(n2937), .C2(n2934), .A(n3753), .B(n2936), .ZN(n2943)
         );
  INV_X1 U3428 ( .A(n3020), .ZN(n2941) );
  AOI22_X1 U3429 ( .A1(n5040), .A2(n3929), .B1(n5045), .B2(n2843), .ZN(n2940)
         );
  AOI21_X1 U3430 ( .B1(n5050), .B2(n3019), .A(n2938), .ZN(n2939) );
  OAI211_X1 U3431 ( .C1(n5054), .C2(n2941), .A(n2940), .B(n2939), .ZN(n2942)
         );
  OR2_X1 U3432 ( .A1(n2943), .A2(n2942), .ZN(U3227) );
  INV_X1 U3433 ( .A(n4397), .ZN(n4934) );
  NAND2_X1 U3434 ( .A1(n2260), .A2(n4934), .ZN(n2944) );
  OAI21_X1 U3435 ( .B1(n3882), .B2(n2946), .A(n2945), .ZN(n4892) );
  INV_X1 U3436 ( .A(n3867), .ZN(n3798) );
  XNOR2_X1 U3437 ( .A(n3882), .B(n3798), .ZN(n2951) );
  OAI22_X1 U3438 ( .A1(n2948), .A2(n4941), .B1(n2947), .B2(n4939), .ZN(n2949)
         );
  AOI21_X1 U3439 ( .B1(n4944), .B2(n3931), .A(n2949), .ZN(n2950) );
  OAI21_X1 U3440 ( .B1(n2951), .B2(n4946), .A(n2950), .ZN(n4894) );
  NAND2_X1 U3441 ( .A1(n4894), .A2(n2260), .ZN(n2958) );
  NAND2_X1 U3442 ( .A1(n3656), .A2(n3795), .ZN(n2952) );
  NAND2_X1 U3443 ( .A1(n2996), .A2(n2952), .ZN(n4891) );
  INV_X1 U3444 ( .A(n4891), .ZN(n2956) );
  INV_X1 U3445 ( .A(REG3_REG_1__SCAN_IN), .ZN(n2953) );
  OAI22_X1 U3446 ( .A1(n2260), .A2(n2954), .B1(n2953), .B2(n4950), .ZN(n2955)
         );
  AOI21_X1 U3447 ( .B1(n5059), .B2(n2956), .A(n2955), .ZN(n2957) );
  OAI211_X1 U3448 ( .C1(n4325), .C2(n4892), .A(n2958), .B(n2957), .ZN(U3289)
         );
  NAND2_X1 U3449 ( .A1(n2843), .A2(n2959), .ZN(n2960) );
  NAND2_X1 U3450 ( .A1(n2963), .A2(n2962), .ZN(n2964) );
  INV_X1 U3451 ( .A(n3930), .ZN(n2973) );
  NAND2_X1 U3452 ( .A1(n2973), .A2(n3019), .ZN(n3805) );
  INV_X1 U3453 ( .A(n3019), .ZN(n2965) );
  NAND2_X1 U3454 ( .A1(n3930), .A2(n2965), .ZN(n3808) );
  NAND2_X1 U3455 ( .A1(n3930), .A2(n3019), .ZN(n2966) );
  NAND2_X1 U3456 ( .A1(n3011), .A2(n2966), .ZN(n3054) );
  AND2_X1 U3457 ( .A1(n3929), .A2(n3051), .ZN(n3058) );
  INV_X1 U34580 ( .A(n3058), .ZN(n3807) );
  INV_X1 U34590 ( .A(n3929), .ZN(n3052) );
  NAND2_X1 U3460 ( .A1(n3052), .A2(n3055), .ZN(n3824) );
  XOR2_X1 U3461 ( .A(n3054), .B(n3880), .Z(n4920) );
  AOI21_X1 U3462 ( .B1(n3055), .B2(n3016), .A(n3063), .ZN(n4923) );
  INV_X1 U3463 ( .A(n2967), .ZN(n2968) );
  OAI22_X1 U3464 ( .A1(n2260), .A2(n2969), .B1(n2968), .B2(n4950), .ZN(n2970)
         );
  AOI21_X1 U3465 ( .B1(n4923), .B2(n5059), .A(n2970), .ZN(n2978) );
  INV_X1 U3466 ( .A(n3805), .ZN(n2972) );
  XNOR2_X1 U34670 ( .A(n3059), .B(n3880), .ZN(n2976) );
  OAI22_X1 U3468 ( .A1(n2973), .A2(n4941), .B1(n3051), .B2(n4939), .ZN(n2974)
         );
  AOI21_X1 U34690 ( .B1(n4944), .B2(n3928), .A(n2974), .ZN(n2975) );
  OAI21_X1 U3470 ( .B1(n2976), .B2(n4946), .A(n2975), .ZN(n4922) );
  NAND2_X1 U34710 ( .A1(n4922), .A2(n2260), .ZN(n2977) );
  OAI211_X1 U3472 ( .C1(n4920), .C2(n4325), .A(n2978), .B(n2977), .ZN(U3285)
         );
  NOR2_X1 U34730 ( .A1(n4983), .A2(n3797), .ZN(n2979) );
  NOR2_X1 U3474 ( .A1(n2980), .A2(n2979), .ZN(n2982) );
  INV_X1 U34750 ( .A(n2985), .ZN(n2986) );
  AOI21_X1 U3476 ( .B1(n3884), .B2(n2987), .A(n2986), .ZN(n4898) );
  OAI21_X1 U34770 ( .B1(n3884), .B2(n2989), .A(n2988), .ZN(n2994) );
  AOI22_X1 U3478 ( .A1(n2843), .A2(n4944), .B1(n2995), .B2(n4417), .ZN(n2991)
         );
  OAI21_X1 U34790 ( .B1(n2990), .B2(n4941), .A(n2991), .ZN(n2993) );
  NOR2_X1 U3480 ( .A1(n4898), .A2(n4397), .ZN(n2992) );
  AOI211_X1 U34810 ( .C1(n4878), .C2(n2994), .A(n2993), .B(n2992), .ZN(n4904)
         );
  OAI21_X1 U3482 ( .B1(n4898), .B2(n4983), .A(n4904), .ZN(n3004) );
  NAND2_X1 U34830 ( .A1(n3004), .A2(n5022), .ZN(n3000) );
  AND2_X1 U3484 ( .A1(n2996), .A2(n2995), .ZN(n2997) );
  NOR2_X1 U34850 ( .A1(n2998), .A2(n2997), .ZN(n4899) );
  INV_X1 U3486 ( .A(n4487), .ZN(n3113) );
  NAND2_X1 U34870 ( .A1(n4899), .A2(n3113), .ZN(n2999) );
  OAI211_X1 U3488 ( .C1(n5022), .C2(n3001), .A(n3000), .B(n2999), .ZN(U3520)
         );
  INV_X1 U34890 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3007) );
  NAND2_X1 U3490 ( .A1(n3004), .A2(n5025), .ZN(n3006) );
  INV_X1 U34910 ( .A(n4751), .ZN(n3117) );
  NAND2_X1 U3492 ( .A1(n3117), .A2(n4899), .ZN(n3005) );
  OAI211_X1 U34930 ( .C1(n5025), .C2(n3007), .A(n3006), .B(n3005), .ZN(U3471)
         );
  XNOR2_X1 U3494 ( .A(n3008), .B(n2268), .ZN(n3015) );
  NAND2_X1 U34950 ( .A1(n3009), .A2(n2268), .ZN(n3010) );
  NAND2_X1 U3496 ( .A1(n3011), .A2(n3010), .ZN(n4912) );
  AOI22_X1 U34970 ( .A1(n2843), .A2(n4391), .B1(n3019), .B2(n4417), .ZN(n3013)
         );
  NAND2_X1 U3498 ( .A1(n3929), .A2(n4944), .ZN(n3012) );
  OAI211_X1 U34990 ( .C1(n4912), .C2(n4397), .A(n3013), .B(n3012), .ZN(n3014)
         );
  AOI21_X1 U3500 ( .B1(n3015), .B2(n4878), .A(n3014), .ZN(n4913) );
  INV_X1 U35010 ( .A(n3016), .ZN(n3017) );
  AOI211_X1 U3502 ( .C1(n3019), .C2(n3018), .A(n5007), .B(n3017), .ZN(n4915)
         );
  AOI22_X1 U35030 ( .A1(n4915), .A2(n4034), .B1(n3020), .B2(n4897), .ZN(n3021)
         );
  AOI21_X1 U3504 ( .B1(n4913), .B2(n3021), .A(n5058), .ZN(n3023) );
  OAI22_X1 U35050 ( .A1(n4912), .A2(n4406), .B1(n2821), .B2(n2260), .ZN(n3022)
         );
  OR2_X1 U35060 ( .A1(n3023), .A2(n3022), .ZN(U3286) );
  NAND2_X1 U35070 ( .A1(n3928), .A2(n3477), .ZN(n3029) );
  MUX2_X1 U35080 ( .A(n3027), .B(DATAI_6_), .S(n2261), .Z(n3080) );
  NAND2_X1 U35090 ( .A1(n3080), .A2(n2786), .ZN(n3028) );
  NAND2_X1 U35100 ( .A1(n3029), .A2(n3028), .ZN(n3030) );
  XNOR2_X1 U35110 ( .A(n3030), .B(n3596), .ZN(n3033) );
  NAND2_X1 U35120 ( .A1(n3928), .A2(n3548), .ZN(n3032) );
  NAND2_X1 U35130 ( .A1(n3080), .A2(n3477), .ZN(n3031) );
  NAND2_X1 U35140 ( .A1(n3032), .A2(n3031), .ZN(n3034) );
  INV_X1 U35150 ( .A(n3033), .ZN(n3036) );
  INV_X1 U35160 ( .A(n3034), .ZN(n3035) );
  NAND2_X1 U35170 ( .A1(n3036), .A2(n3035), .ZN(n3123) );
  NAND2_X1 U35180 ( .A1(n2306), .A2(n3123), .ZN(n3037) );
  XNOR2_X1 U35190 ( .A(n3121), .B(n3037), .ZN(n3049) );
  INV_X1 U35200 ( .A(n3038), .ZN(n3073) );
  NAND2_X1 U35210 ( .A1(n3774), .A2(REG0_REG_7__SCAN_IN), .ZN(n3044) );
  NAND2_X1 U35220 ( .A1(n3039), .A2(REG3_REG_7__SCAN_IN), .ZN(n3084) );
  OR2_X1 U35230 ( .A1(n3039), .A2(REG3_REG_7__SCAN_IN), .ZN(n3040) );
  NAND2_X1 U35240 ( .A1(n3084), .A2(n3040), .ZN(n4951) );
  INV_X1 U35250 ( .A(n4951), .ZN(n3622) );
  NAND2_X1 U35260 ( .A1(n2797), .A2(n3622), .ZN(n3043) );
  NAND2_X1 U35270 ( .A1(n2800), .A2(REG1_REG_7__SCAN_IN), .ZN(n3042) );
  OR2_X1 U35280 ( .A1(n2802), .A2(n2681), .ZN(n3041) );
  NAND4_X1 U35290 ( .A1(n3044), .A2(n3043), .A3(n3042), .A4(n3041), .ZN(n3927)
         );
  AOI22_X1 U35300 ( .A1(n5040), .A2(n3927), .B1(n5045), .B2(n3929), .ZN(n3047)
         );
  NOR2_X1 U35310 ( .A1(STATE_REG_SCAN_IN), .A2(n3045), .ZN(n4804) );
  AOI21_X1 U35320 ( .B1(n5050), .B2(n3080), .A(n4804), .ZN(n3046) );
  OAI211_X1 U35330 ( .C1(n5054), .C2(n3073), .A(n3047), .B(n3046), .ZN(n3048)
         );
  AOI21_X1 U35340 ( .B1(n3049), .B2(n5048), .A(n3048), .ZN(n3050) );
  INV_X1 U35350 ( .A(n3050), .ZN(U3236) );
  NAND2_X1 U35360 ( .A1(n2466), .A2(n3080), .ZN(n3810) );
  NAND2_X1 U35370 ( .A1(n3928), .A2(n2465), .ZN(n3825) );
  AND2_X1 U35380 ( .A1(n3810), .A2(n3825), .ZN(n3890) );
  NAND2_X1 U35390 ( .A1(n3052), .A2(n3051), .ZN(n3053) );
  NAND2_X1 U35400 ( .A1(n3054), .A2(n3053), .ZN(n3057) );
  NAND2_X1 U35410 ( .A1(n3929), .A2(n3055), .ZN(n3056) );
  XOR2_X1 U35420 ( .A(n3890), .B(n3082), .Z(n3074) );
  XNOR2_X1 U35430 ( .A(n3090), .B(n3890), .ZN(n3062) );
  INV_X1 U35440 ( .A(n3927), .ZN(n3101) );
  AOI22_X1 U35450 ( .A1(n3929), .A2(n4391), .B1(n3080), .B2(n4417), .ZN(n3060)
         );
  OAI21_X1 U35460 ( .B1(n3101), .B2(n4880), .A(n3060), .ZN(n3061) );
  AOI21_X1 U35470 ( .B1(n3062), .B2(n4878), .A(n3061), .ZN(n3079) );
  OAI21_X1 U35480 ( .B1(n3074), .B2(n5015), .A(n3079), .ZN(n3070) );
  NOR2_X1 U35490 ( .A1(n3063), .A2(n2465), .ZN(n3064) );
  OR2_X1 U35500 ( .A1(n4929), .A2(n3064), .ZN(n3072) );
  INV_X1 U35510 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3065) );
  OAI22_X1 U35520 ( .A1(n3072), .A2(n4487), .B1(n5022), .B2(n3065), .ZN(n3066)
         );
  AOI21_X1 U35530 ( .B1(n3070), .B2(n5022), .A(n3066), .ZN(n3067) );
  INV_X1 U35540 ( .A(n3067), .ZN(U3524) );
  INV_X1 U35550 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3068) );
  OAI22_X1 U35560 ( .A1(n3072), .A2(n4751), .B1(n5025), .B2(n3068), .ZN(n3069)
         );
  AOI21_X1 U35570 ( .B1(n3070), .B2(n5025), .A(n3069), .ZN(n3071) );
  INV_X1 U35580 ( .A(n3071), .ZN(U3479) );
  INV_X1 U35590 ( .A(n3072), .ZN(n3077) );
  OAI22_X1 U35600 ( .A1(n2260), .A2(n4803), .B1(n3073), .B2(n4950), .ZN(n3076)
         );
  NOR2_X1 U35610 ( .A1(n3074), .A2(n4325), .ZN(n3075) );
  AOI211_X1 U35620 ( .C1(n3077), .C2(n5059), .A(n3076), .B(n3075), .ZN(n3078)
         );
  OAI21_X1 U35630 ( .B1(n5058), .B2(n3079), .A(n3078), .ZN(U3284) );
  AND2_X1 U35640 ( .A1(n3928), .A2(n3080), .ZN(n3081) );
  MUX2_X1 U35650 ( .A(n4761), .B(DATAI_7_), .S(n2261), .Z(n3128) );
  NAND2_X1 U35660 ( .A1(n3101), .A2(n3128), .ZN(n3811) );
  NAND2_X1 U35670 ( .A1(n3927), .A2(n4940), .ZN(n3823) );
  NAND2_X1 U35680 ( .A1(n3927), .A2(n3128), .ZN(n3208) );
  NAND2_X1 U35690 ( .A1(n2800), .A2(REG1_REG_8__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U35700 ( .A1(n3084), .A2(n4573), .ZN(n3085) );
  AND2_X1 U35710 ( .A1(n3094), .A2(n3085), .ZN(n3105) );
  NAND2_X1 U35720 ( .A1(n2797), .A2(n3105), .ZN(n3088) );
  NAND2_X1 U35730 ( .A1(n3774), .A2(REG0_REG_8__SCAN_IN), .ZN(n3087) );
  INV_X1 U35740 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3106) );
  OR2_X1 U35750 ( .A1(n2802), .A2(n3106), .ZN(n3086) );
  NAND4_X1 U35760 ( .A1(n3089), .A2(n3088), .A3(n3087), .A4(n3086), .ZN(n4943)
         );
  INV_X1 U35770 ( .A(n4943), .ZN(n3164) );
  MUX2_X1 U35780 ( .A(n4760), .B(DATAI_8_), .S(n2261), .Z(n3150) );
  NAND2_X1 U35790 ( .A1(n3164), .A2(n3150), .ZN(n3814) );
  INV_X1 U35800 ( .A(n3150), .ZN(n3151) );
  NAND2_X1 U35810 ( .A1(n4943), .A2(n3151), .ZN(n3826) );
  AND2_X1 U3582 ( .A1(n3814), .A2(n3826), .ZN(n3891) );
  XNOR2_X1 U3583 ( .A(n3251), .B(n3891), .ZN(n3112) );
  INV_X1 U3584 ( .A(n3112), .ZN(n3110) );
  INV_X1 U3585 ( .A(n3811), .ZN(n3092) );
  XNOR2_X1 U3586 ( .A(n3156), .B(n3891), .ZN(n3104) );
  NAND2_X1 U3587 ( .A1(n3774), .A2(REG0_REG_9__SCAN_IN), .ZN(n3100) );
  NAND2_X1 U3588 ( .A1(n2800), .A2(REG1_REG_9__SCAN_IN), .ZN(n3099) );
  AND2_X1 U3589 ( .A1(n3094), .A2(n3093), .ZN(n3095) );
  NOR2_X1 U3590 ( .A1(n3157), .A2(n3095), .ZN(n3183) );
  NAND2_X1 U3591 ( .A1(n2797), .A2(n3183), .ZN(n3098) );
  INV_X1 U3592 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3096) );
  OR2_X1 U3593 ( .A1(n2802), .A2(n3096), .ZN(n3097) );
  NAND4_X1 U3594 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .ZN(n3926)
         );
  OAI22_X1 U3595 ( .A1(n3101), .A2(n4941), .B1(n3151), .B2(n4939), .ZN(n3102)
         );
  AOI21_X1 U3596 ( .B1(n4944), .B2(n3926), .A(n3102), .ZN(n3103) );
  OAI21_X1 U3597 ( .B1(n3104), .B2(n4946), .A(n3103), .ZN(n3111) );
  NAND2_X1 U3598 ( .A1(n3111), .A2(n2260), .ZN(n3109) );
  AOI21_X1 U3599 ( .B1(n3150), .B2(n4928), .A(n3171), .ZN(n3118) );
  INV_X1 U3600 ( .A(n3105), .ZN(n3146) );
  OAI22_X1 U3601 ( .A1(n2260), .A2(n3106), .B1(n3146), .B2(n4950), .ZN(n3107)
         );
  AOI21_X1 U3602 ( .B1(n3118), .B2(n5059), .A(n3107), .ZN(n3108) );
  OAI211_X1 U3603 ( .C1(n4325), .C2(n3110), .A(n3109), .B(n3108), .ZN(U3282)
         );
  AOI21_X1 U3604 ( .B1(n3112), .B2(n5010), .A(n3111), .ZN(n3120) );
  AOI22_X1 U3605 ( .A1(n3118), .A2(n3113), .B1(n5021), .B2(REG1_REG_8__SCAN_IN), .ZN(n3114) );
  OAI21_X1 U3606 ( .B1(n3120), .B2(n5021), .A(n3114), .ZN(U3526) );
  INV_X1 U3607 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3115) );
  NOR2_X1 U3608 ( .A1(n5025), .A2(n3115), .ZN(n3116) );
  AOI21_X1 U3609 ( .B1(n3118), .B2(n3117), .A(n3116), .ZN(n3119) );
  OAI21_X1 U3610 ( .B1(n3120), .B2(n5023), .A(n3119), .ZN(U3483) );
  NAND2_X1 U3611 ( .A1(n3927), .A2(n3477), .ZN(n3126) );
  NAND2_X1 U3612 ( .A1(n3128), .A2(n2786), .ZN(n3125) );
  NAND2_X1 U3613 ( .A1(n3126), .A2(n3125), .ZN(n3127) );
  XNOR2_X1 U3614 ( .A(n3127), .B(n3596), .ZN(n3131) );
  AOI22_X1 U3615 ( .A1(n3927), .A2(n3548), .B1(n3477), .B2(n3128), .ZN(n3129)
         );
  XNOR2_X1 U3616 ( .A(n3131), .B(n3129), .ZN(n3619) );
  INV_X1 U3617 ( .A(n3129), .ZN(n3130) );
  NAND2_X1 U3618 ( .A1(n4943), .A2(n3477), .ZN(n3133) );
  NAND2_X1 U3619 ( .A1(n3150), .A2(n2786), .ZN(n3132) );
  NAND2_X1 U3620 ( .A1(n3133), .A2(n3132), .ZN(n3134) );
  XNOR2_X1 U3621 ( .A(n3134), .B(n3596), .ZN(n3137) );
  NAND2_X1 U3622 ( .A1(n4943), .A2(n3548), .ZN(n3136) );
  NAND2_X1 U3623 ( .A1(n3150), .A2(n3477), .ZN(n3135) );
  NAND2_X1 U3624 ( .A1(n3136), .A2(n3135), .ZN(n3138) );
  AND2_X1 U3625 ( .A1(n3137), .A2(n3138), .ZN(n3177) );
  INV_X1 U3626 ( .A(n3177), .ZN(n3141) );
  INV_X1 U3627 ( .A(n3137), .ZN(n3140) );
  INV_X1 U3628 ( .A(n3138), .ZN(n3139) );
  NAND2_X1 U3629 ( .A1(n3140), .A2(n3139), .ZN(n3176) );
  NAND2_X1 U3630 ( .A1(n3141), .A2(n3176), .ZN(n3142) );
  XNOR2_X1 U3631 ( .A(n3178), .B(n3142), .ZN(n3148) );
  AOI22_X1 U3632 ( .A1(n5040), .A2(n3926), .B1(n5045), .B2(n3927), .ZN(n3145)
         );
  AOI21_X1 U3633 ( .B1(n5050), .B2(n3150), .A(n3143), .ZN(n3144) );
  OAI211_X1 U3634 ( .C1(n5054), .C2(n3146), .A(n3145), .B(n3144), .ZN(n3147)
         );
  AOI21_X1 U3635 ( .B1(n3148), .B2(n5048), .A(n3147), .ZN(n3149) );
  INV_X1 U3636 ( .A(n3149), .ZN(U3218) );
  NAND2_X1 U3637 ( .A1(n4943), .A2(n3150), .ZN(n3205) );
  INV_X1 U3638 ( .A(n3205), .ZN(n3152) );
  NAND2_X1 U3639 ( .A1(n3164), .A2(n3151), .ZN(n3210) );
  OAI21_X1 U3640 ( .B1(n3251), .B2(n3152), .A(n3210), .ZN(n3155) );
  NAND2_X1 U3641 ( .A1(n3153), .A2(IR_REG_31__SCAN_IN), .ZN(n3154) );
  XNOR2_X1 U3642 ( .A(n3154), .B(IR_REG_9__SCAN_IN), .ZN(n4810) );
  MUX2_X1 U3643 ( .A(n4810), .B(DATAI_9_), .S(n2261), .Z(n3203) );
  AND2_X1 U3644 ( .A1(n3926), .A2(n3170), .ZN(n3820) );
  INV_X1 U3645 ( .A(n3820), .ZN(n3827) );
  INV_X1 U3646 ( .A(n3926), .ZN(n3202) );
  NAND2_X1 U3647 ( .A1(n3202), .A2(n3203), .ZN(n3815) );
  NAND2_X1 U3648 ( .A1(n3827), .A2(n3815), .ZN(n3871) );
  XNOR2_X1 U3649 ( .A(n3155), .B(n3871), .ZN(n3166) );
  INV_X1 U3650 ( .A(n3166), .ZN(n4960) );
  XOR2_X1 U3651 ( .A(n3871), .B(n3187), .Z(n3169) );
  NAND2_X1 U3652 ( .A1(n2800), .A2(REG1_REG_10__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U3653 ( .A1(n3774), .A2(REG0_REG_10__SCAN_IN), .ZN(n3162) );
  NOR2_X1 U3654 ( .A1(n3157), .A2(REG3_REG_10__SCAN_IN), .ZN(n3158) );
  OR2_X1 U3655 ( .A1(n3192), .A2(n3158), .ZN(n3322) );
  INV_X1 U3656 ( .A(n3322), .ZN(n3215) );
  NAND2_X1 U3657 ( .A1(n2797), .A2(n3215), .ZN(n3161) );
  INV_X1 U3658 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3159) );
  OR2_X1 U3659 ( .A1(n2802), .A2(n3159), .ZN(n3160) );
  NAND4_X1 U3660 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3925)
         );
  OAI22_X1 U3661 ( .A1(n3164), .A2(n4941), .B1(n4939), .B2(n3170), .ZN(n3165)
         );
  AOI21_X1 U3662 ( .B1(n4944), .B2(n3925), .A(n3165), .ZN(n3168) );
  NAND2_X1 U3663 ( .A1(n3166), .A2(n4934), .ZN(n3167) );
  OAI211_X1 U3664 ( .C1(n3169), .C2(n4946), .A(n3168), .B(n3167), .ZN(n4961)
         );
  NAND2_X1 U3665 ( .A1(n4961), .A2(n2260), .ZN(n3175) );
  AOI21_X1 U3666 ( .B1(n3203), .B2(n2323), .A(n2305), .ZN(n4963) );
  INV_X1 U3667 ( .A(n3183), .ZN(n3172) );
  OAI22_X1 U3668 ( .A1(n2260), .A2(n3096), .B1(n3172), .B2(n4950), .ZN(n3173)
         );
  AOI21_X1 U3669 ( .B1(n4963), .B2(n5059), .A(n3173), .ZN(n3174) );
  OAI211_X1 U3670 ( .C1(n4960), .C2(n4406), .A(n3175), .B(n3174), .ZN(U3281)
         );
  NAND2_X1 U3671 ( .A1(n3926), .A2(n3477), .ZN(n3180) );
  NAND2_X1 U3672 ( .A1(n3203), .A2(n2786), .ZN(n3179) );
  NAND2_X1 U3673 ( .A1(n3180), .A2(n3179), .ZN(n3181) );
  XNOR2_X1 U3674 ( .A(n3181), .B(n3596), .ZN(n3288) );
  AOI22_X1 U3675 ( .A1(n3926), .A2(n3548), .B1(n3477), .B2(n3203), .ZN(n3289)
         );
  XNOR2_X1 U3676 ( .A(n3288), .B(n3289), .ZN(n3286) );
  XOR2_X1 U3677 ( .A(n3287), .B(n3286), .Z(n3186) );
  AOI22_X1 U3678 ( .A1(n5040), .A2(n3925), .B1(n5045), .B2(n4943), .ZN(n3185)
         );
  AND2_X1 U3679 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4814) );
  NOR2_X1 U3680 ( .A1(n3748), .A2(n3170), .ZN(n3182) );
  AOI211_X1 U3681 ( .C1(n3183), .C2(n3750), .A(n4814), .B(n3182), .ZN(n3184)
         );
  OAI211_X1 U3682 ( .C1(n3186), .C2(n3753), .A(n3185), .B(n3184), .ZN(U3228)
         );
  INV_X1 U3683 ( .A(n3187), .ZN(n3188) );
  INV_X1 U3684 ( .A(n3925), .ZN(n3253) );
  OR2_X1 U3685 ( .A1(n3189), .A2(n3190), .ZN(n3191) );
  XNOR2_X1 U3686 ( .A(n3191), .B(IR_REG_10__SCAN_IN), .ZN(n4967) );
  MUX2_X1 U3687 ( .A(n4967), .B(DATAI_10_), .S(n2261), .Z(n3319) );
  NAND2_X1 U3688 ( .A1(n3253), .A2(n3319), .ZN(n3829) );
  NAND2_X1 U3689 ( .A1(n3925), .A2(n2320), .ZN(n3817) );
  NAND2_X1 U3690 ( .A1(n3829), .A2(n3817), .ZN(n3872) );
  XNOR2_X1 U3691 ( .A(n3220), .B(n3872), .ZN(n3201) );
  NAND2_X1 U3692 ( .A1(n2800), .A2(REG1_REG_11__SCAN_IN), .ZN(n3198) );
  OR2_X1 U3693 ( .A1(n3192), .A2(REG3_REG_11__SCAN_IN), .ZN(n3193) );
  AND2_X1 U3694 ( .A1(n3227), .A2(n3193), .ZN(n3273) );
  NAND2_X1 U3695 ( .A1(n2797), .A2(n3273), .ZN(n3197) );
  NAND2_X1 U3696 ( .A1(n3774), .A2(REG0_REG_11__SCAN_IN), .ZN(n3196) );
  INV_X1 U3697 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3194) );
  OR2_X1 U3698 ( .A1(n2802), .A2(n3194), .ZN(n3195) );
  NAND4_X1 U3699 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3924)
         );
  INV_X1 U3700 ( .A(n3924), .ZN(n3255) );
  OAI22_X1 U3701 ( .A1(n3255), .A2(n4880), .B1(n2320), .B2(n4939), .ZN(n3199)
         );
  AOI21_X1 U3702 ( .B1(n4391), .B2(n3926), .A(n3199), .ZN(n3200) );
  OAI21_X1 U3703 ( .B1(n3201), .B2(n4946), .A(n3200), .ZN(n3278) );
  INV_X1 U3704 ( .A(n3278), .ZN(n3219) );
  NAND2_X1 U3705 ( .A1(n3202), .A2(n3170), .ZN(n3209) );
  INV_X1 U3706 ( .A(n3209), .ZN(n3207) );
  NAND2_X1 U3707 ( .A1(n3926), .A2(n3203), .ZN(n3204) );
  AND2_X1 U3708 ( .A1(n3205), .A2(n3204), .ZN(n3206) );
  INV_X1 U3709 ( .A(n3252), .ZN(n3211) );
  AND2_X1 U3710 ( .A1(n3210), .A2(n3209), .ZN(n3249) );
  OR2_X1 U3711 ( .A1(n3211), .A2(n3249), .ZN(n3212) );
  NAND2_X1 U3712 ( .A1(n3213), .A2(n3212), .ZN(n3247) );
  XNOR2_X1 U3713 ( .A(n3247), .B(n3872), .ZN(n3279) );
  INV_X1 U3714 ( .A(n3272), .ZN(n3214) );
  OAI21_X1 U3715 ( .B1(n2305), .B2(n2320), .A(n3214), .ZN(n3285) );
  AOI22_X1 U3716 ( .A1(n5058), .A2(REG2_REG_10__SCAN_IN), .B1(n3215), .B2(
        n4897), .ZN(n3216) );
  OAI21_X1 U3717 ( .B1(n3285), .B2(n4338), .A(n3216), .ZN(n3217) );
  AOI21_X1 U3718 ( .B1(n3279), .B2(n4365), .A(n3217), .ZN(n3218) );
  OAI21_X1 U3719 ( .B1(n3219), .B2(n5058), .A(n3218), .ZN(U3280) );
  INV_X1 U3720 ( .A(IR_REG_10__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U3721 ( .A1(n3189), .A2(n3221), .ZN(n3222) );
  NAND2_X1 U3722 ( .A1(n3222), .A2(IR_REG_31__SCAN_IN), .ZN(n3224) );
  INV_X1 U3723 ( .A(IR_REG_11__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U3724 ( .A1(n3224), .A2(n3223), .ZN(n3234) );
  OR2_X1 U3725 ( .A1(n3224), .A2(n3223), .ZN(n3225) );
  MUX2_X1 U3726 ( .A(n3965), .B(DATAI_11_), .S(n2261), .Z(n3307) );
  NAND2_X1 U3727 ( .A1(n3924), .A2(n3271), .ZN(n3818) );
  NAND2_X1 U3728 ( .A1(n3262), .A2(n3818), .ZN(n3226) );
  NAND2_X1 U3729 ( .A1(n3255), .A2(n3307), .ZN(n3831) );
  NAND2_X1 U3730 ( .A1(n2800), .A2(REG1_REG_12__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U3731 ( .A1(n3227), .A2(n4684), .ZN(n3228) );
  AND2_X1 U3732 ( .A1(n3237), .A2(n3228), .ZN(n3343) );
  NAND2_X1 U3733 ( .A1(n2797), .A2(n3343), .ZN(n3232) );
  NAND2_X1 U3734 ( .A1(n3774), .A2(REG0_REG_12__SCAN_IN), .ZN(n3231) );
  INV_X1 U3735 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3229) );
  OR2_X1 U3736 ( .A1(n2802), .A2(n3229), .ZN(n3230) );
  NAND4_X1 U3737 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n4392)
         );
  NAND2_X1 U3738 ( .A1(n3234), .A2(IR_REG_31__SCAN_IN), .ZN(n3235) );
  XNOR2_X1 U3739 ( .A(n3235), .B(IR_REG_12__SCAN_IN), .ZN(n3967) );
  MUX2_X1 U3740 ( .A(n3967), .B(DATAI_12_), .S(n2261), .Z(n4040) );
  INV_X1 U3741 ( .A(n4040), .ZN(n4050) );
  NAND2_X1 U3742 ( .A1(n4392), .A2(n4050), .ZN(n4386) );
  INV_X1 U3743 ( .A(n4386), .ZN(n3236) );
  NOR2_X1 U3744 ( .A1(n4392), .A2(n4050), .ZN(n4387) );
  OR2_X1 U3745 ( .A1(n3236), .A2(n4387), .ZN(n3256) );
  INV_X1 U3746 ( .A(n3256), .ZN(n3881) );
  XNOR2_X1 U3747 ( .A(n4388), .B(n3881), .ZN(n3246) );
  NAND2_X1 U3748 ( .A1(n3924), .A2(n4391), .ZN(n3244) );
  NAND2_X1 U3749 ( .A1(n2800), .A2(REG1_REG_13__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U3750 ( .A1(n3237), .A2(n4699), .ZN(n3238) );
  AND2_X1 U3751 ( .A1(n3385), .A2(n3238), .ZN(n4400) );
  NAND2_X1 U3752 ( .A1(n2797), .A2(n4400), .ZN(n3241) );
  NAND2_X1 U3753 ( .A1(n3774), .A2(REG0_REG_13__SCAN_IN), .ZN(n3240) );
  INV_X1 U3754 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4402) );
  OR2_X1 U3755 ( .A1(n2802), .A2(n4402), .ZN(n3239) );
  NAND4_X1 U3756 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n4373)
         );
  NAND2_X1 U3757 ( .A1(n4373), .A2(n4944), .ZN(n3243) );
  OAI211_X1 U3758 ( .C1(n4939), .C2(n4050), .A(n3244), .B(n3243), .ZN(n3245)
         );
  AOI21_X1 U3759 ( .B1(n3246), .B2(n4878), .A(n3245), .ZN(n4485) );
  NAND2_X1 U3760 ( .A1(n3247), .A2(n3253), .ZN(n3248) );
  NAND2_X1 U3761 ( .A1(n3248), .A2(n3319), .ZN(n4047) );
  AND2_X1 U3762 ( .A1(n3249), .A2(n3925), .ZN(n3250) );
  NAND2_X1 U3763 ( .A1(n3251), .A2(n3250), .ZN(n4045) );
  OR2_X1 U3764 ( .A1(n3253), .A2(n3252), .ZN(n4042) );
  AND2_X1 U3765 ( .A1(n4045), .A2(n4042), .ZN(n3254) );
  NAND2_X1 U3766 ( .A1(n4047), .A2(n3254), .ZN(n3263) );
  NAND2_X1 U3767 ( .A1(n3255), .A2(n3271), .ZN(n4048) );
  NAND2_X1 U3768 ( .A1(n3265), .A2(n4048), .ZN(n3257) );
  XNOR2_X1 U3769 ( .A(n3257), .B(n3256), .ZN(n4483) );
  NAND2_X1 U3770 ( .A1(n3272), .A2(n3271), .ZN(n3270) );
  NAND2_X1 U3771 ( .A1(n3270), .A2(n4040), .ZN(n3258) );
  NAND2_X1 U3772 ( .A1(n2273), .A2(n3258), .ZN(n4752) );
  AOI22_X1 U3773 ( .A1(n5058), .A2(REG2_REG_12__SCAN_IN), .B1(n3343), .B2(
        n4897), .ZN(n3259) );
  OAI21_X1 U3774 ( .B1(n4752), .B2(n4338), .A(n3259), .ZN(n3260) );
  AOI21_X1 U3775 ( .B1(n4483), .B2(n4365), .A(n3260), .ZN(n3261) );
  OAI21_X1 U3776 ( .B1(n4485), .B2(n5058), .A(n3261), .ZN(U3278) );
  XOR2_X1 U3777 ( .A(n4041), .B(n3262), .Z(n3269) );
  NAND2_X1 U3778 ( .A1(n3263), .A2(n4041), .ZN(n3264) );
  NAND2_X1 U3779 ( .A1(n3265), .A2(n3264), .ZN(n4974) );
  INV_X1 U3780 ( .A(n4392), .ZN(n4051) );
  AOI22_X1 U3781 ( .A1(n3925), .A2(n4391), .B1(n4417), .B2(n3307), .ZN(n3266)
         );
  OAI21_X1 U3782 ( .B1(n4051), .B2(n4880), .A(n3266), .ZN(n3267) );
  AOI21_X1 U3783 ( .B1(n4974), .B2(n4934), .A(n3267), .ZN(n3268) );
  OAI21_X1 U3784 ( .B1(n3269), .B2(n4946), .A(n3268), .ZN(n4972) );
  INV_X1 U3785 ( .A(n4972), .ZN(n3277) );
  OAI21_X1 U3786 ( .B1(n3272), .B2(n3271), .A(n3270), .ZN(n4971) );
  NOR2_X1 U3787 ( .A1(n4971), .A2(n4338), .ZN(n3275) );
  INV_X1 U3788 ( .A(n3273), .ZN(n3310) );
  OAI22_X1 U3789 ( .A1(n2260), .A2(n3194), .B1(n3310), .B2(n4950), .ZN(n3274)
         );
  AOI211_X1 U3790 ( .C1(n4974), .C2(n4900), .A(n3275), .B(n3274), .ZN(n3276)
         );
  OAI21_X1 U3791 ( .B1(n3277), .B2(n5058), .A(n3276), .ZN(U3279) );
  INV_X1 U3792 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3280) );
  AOI21_X1 U3793 ( .B1(n5010), .B2(n3279), .A(n3278), .ZN(n3282) );
  MUX2_X1 U3794 ( .A(n3280), .B(n3282), .S(n5025), .Z(n3281) );
  OAI21_X1 U3795 ( .B1(n3285), .B2(n4751), .A(n3281), .ZN(U3487) );
  INV_X1 U3796 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3283) );
  MUX2_X1 U3797 ( .A(n3283), .B(n3282), .S(n5022), .Z(n3284) );
  OAI21_X1 U3798 ( .B1(n3285), .B2(n4487), .A(n3284), .ZN(U3528) );
  INV_X1 U3799 ( .A(n3288), .ZN(n3290) );
  NAND2_X1 U3800 ( .A1(n3290), .A2(n3289), .ZN(n3291) );
  NAND2_X1 U3801 ( .A1(n3925), .A2(n3477), .ZN(n3293) );
  NAND2_X1 U3802 ( .A1(n3319), .A2(n2786), .ZN(n3292) );
  NAND2_X1 U3803 ( .A1(n3293), .A2(n3292), .ZN(n3294) );
  XNOR2_X1 U3804 ( .A(n3294), .B(n3566), .ZN(n3296) );
  AOI22_X1 U3805 ( .A1(n3925), .A2(n3548), .B1(n3477), .B2(n3319), .ZN(n3297)
         );
  XNOR2_X1 U3806 ( .A(n3296), .B(n3297), .ZN(n3317) );
  INV_X1 U3807 ( .A(n3296), .ZN(n3299) );
  INV_X1 U3808 ( .A(n3297), .ZN(n3298) );
  NAND2_X1 U3809 ( .A1(n3299), .A2(n3298), .ZN(n3300) );
  NAND2_X1 U3810 ( .A1(n3924), .A2(n3477), .ZN(n3302) );
  NAND2_X1 U3811 ( .A1(n3307), .A2(n2786), .ZN(n3301) );
  NAND2_X1 U3812 ( .A1(n3302), .A2(n3301), .ZN(n3303) );
  XNOR2_X1 U3813 ( .A(n3303), .B(n3566), .ZN(n3327) );
  NAND2_X1 U3814 ( .A1(n3924), .A2(n3548), .ZN(n3305) );
  NAND2_X1 U3815 ( .A1(n3307), .A2(n3477), .ZN(n3304) );
  XNOR2_X1 U3816 ( .A(n3327), .B(n3328), .ZN(n3306) );
  XNOR2_X1 U3817 ( .A(n3326), .B(n3306), .ZN(n3312) );
  AOI22_X1 U3818 ( .A1(n5040), .A2(n4392), .B1(n5045), .B2(n3925), .ZN(n3309)
         );
  AND2_X1 U3819 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4834) );
  AOI21_X1 U3820 ( .B1(n5050), .B2(n3307), .A(n4834), .ZN(n3308) );
  OAI211_X1 U3821 ( .C1(n5054), .C2(n3310), .A(n3309), .B(n3308), .ZN(n3311)
         );
  AOI21_X1 U3822 ( .B1(n3312), .B2(n5048), .A(n3311), .ZN(n3313) );
  INV_X1 U3823 ( .A(n3313), .ZN(U3233) );
  INV_X1 U3824 ( .A(n3314), .ZN(n3315) );
  AOI211_X1 U3825 ( .C1(n3317), .C2(n3316), .A(n3753), .B(n3315), .ZN(n3324)
         );
  AOI22_X1 U3826 ( .A1(n5040), .A2(n3924), .B1(n5045), .B2(n3926), .ZN(n3321)
         );
  INV_X1 U3827 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3318) );
  NOR2_X1 U3828 ( .A1(STATE_REG_SCAN_IN), .A2(n3318), .ZN(n4821) );
  AOI21_X1 U3829 ( .B1(n5050), .B2(n3319), .A(n4821), .ZN(n3320) );
  OAI211_X1 U3830 ( .C1(n5054), .C2(n3322), .A(n3321), .B(n3320), .ZN(n3323)
         );
  OR2_X1 U3831 ( .A1(n3324), .A2(n3323), .ZN(U3214) );
  NAND2_X1 U3832 ( .A1(n3327), .A2(n3328), .ZN(n3325) );
  INV_X1 U3833 ( .A(n3327), .ZN(n3330) );
  INV_X1 U3834 ( .A(n3328), .ZN(n3329) );
  NAND2_X1 U3835 ( .A1(n3330), .A2(n3329), .ZN(n3331) );
  NAND2_X1 U3836 ( .A1(n4392), .A2(n3477), .ZN(n3333) );
  NAND2_X1 U3837 ( .A1(n4040), .A2(n2786), .ZN(n3332) );
  NAND2_X1 U3838 ( .A1(n3333), .A2(n3332), .ZN(n3334) );
  XNOR2_X1 U3839 ( .A(n3334), .B(n3596), .ZN(n3337) );
  NAND2_X1 U3840 ( .A1(n4392), .A2(n3548), .ZN(n3336) );
  NAND2_X1 U3841 ( .A1(n4040), .A2(n3477), .ZN(n3335) );
  NAND2_X1 U3842 ( .A1(n3336), .A2(n3335), .ZN(n3338) );
  AND2_X1 U3843 ( .A1(n3337), .A2(n3338), .ZN(n3355) );
  INV_X1 U3844 ( .A(n3355), .ZN(n3341) );
  INV_X1 U3845 ( .A(n3337), .ZN(n3340) );
  INV_X1 U3846 ( .A(n3338), .ZN(n3339) );
  NAND2_X1 U3847 ( .A1(n3340), .A2(n3339), .ZN(n3354) );
  NAND2_X1 U3848 ( .A1(n3341), .A2(n3354), .ZN(n3342) );
  XNOR2_X1 U3849 ( .A(n3356), .B(n3342), .ZN(n3348) );
  INV_X1 U3850 ( .A(n3343), .ZN(n3346) );
  AOI22_X1 U3851 ( .A1(n5040), .A2(n4373), .B1(n5045), .B2(n3924), .ZN(n3345)
         );
  NOR2_X1 U3852 ( .A1(STATE_REG_SCAN_IN), .A2(n4684), .ZN(n4844) );
  AOI21_X1 U3853 ( .B1(n5050), .B2(n4040), .A(n4844), .ZN(n3344) );
  OAI211_X1 U3854 ( .C1(n5054), .C2(n3346), .A(n3345), .B(n3344), .ZN(n3347)
         );
  AOI21_X1 U3855 ( .B1(n3348), .B2(n5048), .A(n3347), .ZN(n3349) );
  INV_X1 U3856 ( .A(n3349), .ZN(U3221) );
  NAND3_X1 U3857 ( .A1(n3350), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3352) );
  INV_X1 U3858 ( .A(DATAI_31_), .ZN(n3351) );
  OAI22_X1 U3859 ( .A1(n3353), .A2(n3352), .B1(STATE_REG_SCAN_IN), .B2(n3351), 
        .ZN(U3321) );
  NAND2_X1 U3860 ( .A1(n4373), .A2(n3477), .ZN(n3362) );
  NAND2_X1 U3861 ( .A1(n3357), .A2(IR_REG_31__SCAN_IN), .ZN(n3358) );
  MUX2_X1 U3862 ( .A(IR_REG_31__SCAN_IN), .B(n3358), .S(IR_REG_13__SCAN_IN), 
        .Z(n3360) );
  AND2_X1 U3863 ( .A1(n3360), .A2(n3359), .ZN(n4852) );
  MUX2_X1 U3864 ( .A(n4852), .B(DATAI_13_), .S(n2261), .Z(n4399) );
  NAND2_X1 U3865 ( .A1(n4399), .A2(n2786), .ZN(n3361) );
  NAND2_X1 U3866 ( .A1(n3362), .A2(n3361), .ZN(n3363) );
  XNOR2_X1 U3867 ( .A(n3363), .B(n3566), .ZN(n3715) );
  NAND2_X1 U3868 ( .A1(n3774), .A2(REG0_REG_14__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U3869 ( .A1(n2800), .A2(REG1_REG_14__SCAN_IN), .ZN(n3366) );
  XNOR2_X1 U3870 ( .A(n3385), .B(REG3_REG_14__SCAN_IN), .ZN(n4380) );
  NAND2_X1 U3871 ( .A1(n2797), .A2(n4380), .ZN(n3365) );
  INV_X1 U3872 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4382) );
  OR2_X1 U3873 ( .A1(n2802), .A2(n4382), .ZN(n3364) );
  NAND4_X1 U3874 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n4350)
         );
  NAND2_X1 U3875 ( .A1(n4350), .A2(n3477), .ZN(n3370) );
  XNOR2_X1 U3876 ( .A(n3368), .B(IR_REG_14__SCAN_IN), .ZN(n4759) );
  MUX2_X1 U3877 ( .A(n4759), .B(DATAI_14_), .S(n2261), .Z(n4378) );
  NAND2_X1 U3878 ( .A1(n4378), .A2(n2786), .ZN(n3369) );
  NAND2_X1 U3879 ( .A1(n3370), .A2(n3369), .ZN(n3371) );
  XNOR2_X1 U3880 ( .A(n3371), .B(n3596), .ZN(n3378) );
  NAND2_X1 U3881 ( .A1(n4350), .A2(n3548), .ZN(n3373) );
  NAND2_X1 U3882 ( .A1(n4378), .A2(n3477), .ZN(n3372) );
  NAND2_X1 U3883 ( .A1(n3373), .A2(n3372), .ZN(n3379) );
  AND2_X1 U3884 ( .A1(n3378), .A2(n3379), .ZN(n3635) );
  INV_X1 U3885 ( .A(n3374), .ZN(n3382) );
  NAND2_X1 U3886 ( .A1(n4373), .A2(n3548), .ZN(n3376) );
  NAND2_X1 U3887 ( .A1(n4399), .A2(n3477), .ZN(n3375) );
  NAND2_X1 U3888 ( .A1(n3376), .A2(n3375), .ZN(n3716) );
  NAND2_X1 U3889 ( .A1(n3377), .A2(n3716), .ZN(n3634) );
  INV_X1 U3890 ( .A(n3378), .ZN(n3381) );
  INV_X1 U3891 ( .A(n3379), .ZN(n3380) );
  NAND2_X1 U3892 ( .A1(n3774), .A2(REG0_REG_15__SCAN_IN), .ZN(n3391) );
  INV_X1 U3893 ( .A(n3385), .ZN(n3383) );
  AOI21_X1 U3894 ( .B1(n3383), .B2(REG3_REG_14__SCAN_IN), .A(
        REG3_REG_15__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U3895 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_15__SCAN_IN), .ZN(
        n3384) );
  OR2_X1 U3896 ( .A1(n3386), .A2(n3402), .ZN(n5004) );
  INV_X1 U3897 ( .A(n5004), .ZN(n3387) );
  NAND2_X1 U3898 ( .A1(n2797), .A2(n3387), .ZN(n3390) );
  NAND2_X1 U3899 ( .A1(n2800), .A2(REG1_REG_15__SCAN_IN), .ZN(n3389) );
  INV_X1 U3900 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4354) );
  OR2_X1 U3901 ( .A1(n2802), .A2(n4354), .ZN(n3388) );
  NAND4_X1 U3902 ( .A1(n3391), .A2(n3390), .A3(n3389), .A4(n3388), .ZN(n4329)
         );
  NAND2_X1 U3903 ( .A1(n4329), .A2(n3477), .ZN(n3395) );
  XNOR2_X1 U3904 ( .A(n3392), .B(n3393), .ZN(n4758) );
  MUX2_X1 U3905 ( .A(n4758), .B(DATAI_15_), .S(n2261), .Z(n4996) );
  NAND2_X1 U3906 ( .A1(n4996), .A2(n2786), .ZN(n3394) );
  NAND2_X1 U3907 ( .A1(n3395), .A2(n3394), .ZN(n3396) );
  XNOR2_X1 U3908 ( .A(n3396), .B(n3596), .ZN(n3398) );
  NAND2_X1 U3909 ( .A1(n3397), .A2(n3398), .ZN(n4998) );
  NAND2_X1 U3910 ( .A1(n4998), .A2(n5000), .ZN(n3401) );
  INV_X1 U3911 ( .A(n3397), .ZN(n3400) );
  INV_X1 U3912 ( .A(n3398), .ZN(n3399) );
  NAND2_X1 U3913 ( .A1(n3400), .A2(n3399), .ZN(n4997) );
  NAND2_X1 U3914 ( .A1(n3401), .A2(n4997), .ZN(n3689) );
  NAND2_X1 U3915 ( .A1(n3774), .A2(REG0_REG_16__SCAN_IN), .ZN(n3407) );
  NAND2_X1 U3916 ( .A1(n2800), .A2(REG1_REG_16__SCAN_IN), .ZN(n3406) );
  NOR2_X1 U3917 ( .A1(n3402), .A2(REG3_REG_16__SCAN_IN), .ZN(n3403) );
  OR2_X1 U3918 ( .A1(n3419), .A2(n3403), .ZN(n4339) );
  INV_X1 U3919 ( .A(n4339), .ZN(n3693) );
  NAND2_X1 U3920 ( .A1(n2797), .A2(n3693), .ZN(n3405) );
  INV_X1 U3921 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4340) );
  OR2_X1 U3922 ( .A1(n2802), .A2(n4340), .ZN(n3404) );
  NAND4_X1 U3923 ( .A1(n3407), .A2(n3406), .A3(n3405), .A4(n3404), .ZN(n4314)
         );
  NAND2_X1 U3924 ( .A1(n4314), .A2(n3477), .ZN(n3413) );
  OAI21_X1 U3925 ( .B1(n3392), .B2(IR_REG_15__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n3408) );
  MUX2_X1 U3926 ( .A(IR_REG_31__SCAN_IN), .B(n3408), .S(IR_REG_16__SCAN_IN), 
        .Z(n3411) );
  OR2_X1 U3927 ( .A1(n3392), .A2(n3409), .ZN(n3410) );
  MUX2_X1 U3928 ( .A(n4003), .B(DATAI_16_), .S(n2261), .Z(n4328) );
  NAND2_X1 U3929 ( .A1(n4328), .A2(n2786), .ZN(n3412) );
  NAND2_X1 U3930 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  XNOR2_X1 U3931 ( .A(n3414), .B(n3596), .ZN(n3415) );
  AOI22_X1 U3932 ( .A1(n4314), .A2(n3548), .B1(n3477), .B2(n4328), .ZN(n3416)
         );
  XNOR2_X1 U3933 ( .A(n3415), .B(n3416), .ZN(n3690) );
  INV_X1 U3934 ( .A(n3415), .ZN(n3417) );
  NAND2_X1 U3935 ( .A1(n3417), .A2(n3416), .ZN(n3418) );
  NAND2_X1 U3936 ( .A1(n3604), .A2(REG2_REG_17__SCAN_IN), .ZN(n3426) );
  NAND2_X1 U3937 ( .A1(n2800), .A2(REG1_REG_17__SCAN_IN), .ZN(n3425) );
  NOR2_X1 U3938 ( .A1(n3419), .A2(REG3_REG_17__SCAN_IN), .ZN(n3420) );
  OR2_X1 U3939 ( .A1(n3436), .A2(n3420), .ZN(n4320) );
  INV_X1 U3940 ( .A(n4320), .ZN(n3421) );
  NAND2_X1 U3941 ( .A1(n2797), .A2(n3421), .ZN(n3424) );
  INV_X1 U3942 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3422) );
  OR2_X1 U3943 ( .A1(n3607), .A2(n3422), .ZN(n3423) );
  NAND4_X1 U3944 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n4293)
         );
  NAND2_X1 U3945 ( .A1(n4293), .A2(n3477), .ZN(n3428) );
  MUX2_X1 U3946 ( .A(n4020), .B(DATAI_17_), .S(n2261), .Z(n4317) );
  NAND2_X1 U3947 ( .A1(n4317), .A2(n2786), .ZN(n3427) );
  NAND2_X1 U3948 ( .A1(n3428), .A2(n3427), .ZN(n3429) );
  XNOR2_X1 U3949 ( .A(n3429), .B(n3566), .ZN(n3699) );
  NAND2_X1 U3950 ( .A1(n4293), .A2(n3548), .ZN(n3431) );
  NAND2_X1 U3951 ( .A1(n4317), .A2(n3477), .ZN(n3430) );
  AND2_X1 U3952 ( .A1(n3431), .A2(n3430), .ZN(n3432) );
  INV_X1 U3953 ( .A(n3699), .ZN(n3433) );
  INV_X1 U3954 ( .A(n3432), .ZN(n3698) );
  NAND2_X1 U3955 ( .A1(n3433), .A2(n3698), .ZN(n3434) );
  NAND2_X1 U3956 ( .A1(n3435), .A2(n3434), .ZN(n3732) );
  NAND2_X1 U3957 ( .A1(n3604), .A2(REG2_REG_18__SCAN_IN), .ZN(n3441) );
  NAND2_X1 U3958 ( .A1(n2800), .A2(REG1_REG_18__SCAN_IN), .ZN(n3440) );
  OR2_X1 U3959 ( .A1(n3436), .A2(REG3_REG_18__SCAN_IN), .ZN(n3437) );
  AND2_X1 U3960 ( .A1(n3437), .A2(n3453), .ZN(n4303) );
  NAND2_X1 U3961 ( .A1(n2797), .A2(n4303), .ZN(n3439) );
  INV_X1 U3962 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4741) );
  OR2_X1 U3963 ( .A1(n3607), .A2(n4741), .ZN(n3438) );
  NAND4_X1 U3964 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(n5027)
         );
  NAND2_X1 U3965 ( .A1(n5027), .A2(n3477), .ZN(n3444) );
  INV_X1 U3966 ( .A(IR_REG_18__SCAN_IN), .ZN(n3442) );
  XNOR2_X1 U3967 ( .A(n2293), .B(n3442), .ZN(n4757) );
  MUX2_X1 U3968 ( .A(n4757), .B(DATAI_18_), .S(n2261), .Z(n3761) );
  NAND2_X1 U3969 ( .A1(n3761), .A2(n2786), .ZN(n3443) );
  NAND2_X1 U3970 ( .A1(n3444), .A2(n3443), .ZN(n3445) );
  XNOR2_X1 U3971 ( .A(n3445), .B(n3596), .ZN(n3451) );
  INV_X1 U3972 ( .A(n3451), .ZN(n3449) );
  NAND2_X1 U3973 ( .A1(n5027), .A2(n3548), .ZN(n3447) );
  NAND2_X1 U3974 ( .A1(n3761), .A2(n3477), .ZN(n3446) );
  NAND2_X1 U3975 ( .A1(n3447), .A2(n3446), .ZN(n3450) );
  INV_X1 U3976 ( .A(n3450), .ZN(n3448) );
  NAND2_X1 U3977 ( .A1(n3449), .A2(n3448), .ZN(n3734) );
  AND2_X1 U3978 ( .A1(n3451), .A2(n3450), .ZN(n3733) );
  NAND2_X1 U3979 ( .A1(n3774), .A2(REG0_REG_19__SCAN_IN), .ZN(n3459) );
  NAND2_X1 U3980 ( .A1(n3453), .A2(n3452), .ZN(n3454) );
  NAND2_X1 U3981 ( .A1(n3468), .A2(n3454), .ZN(n5038) );
  INV_X1 U3982 ( .A(n5038), .ZN(n4286) );
  NAND2_X1 U3983 ( .A1(n2797), .A2(n4286), .ZN(n3458) );
  NAND2_X1 U3984 ( .A1(n2800), .A2(REG1_REG_19__SCAN_IN), .ZN(n3457) );
  INV_X1 U3985 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3455) );
  OR2_X1 U3986 ( .A1(n2802), .A2(n3455), .ZN(n3456) );
  NAND2_X1 U3987 ( .A1(n5046), .A2(n3477), .ZN(n3461) );
  MUX2_X1 U3988 ( .A(n4936), .B(DATAI_19_), .S(n2261), .Z(n5026) );
  NAND2_X1 U3989 ( .A1(n5026), .A2(n2786), .ZN(n3460) );
  NAND2_X1 U3990 ( .A1(n3461), .A2(n3460), .ZN(n3462) );
  XNOR2_X1 U3991 ( .A(n3462), .B(n3596), .ZN(n3463) );
  AOI22_X1 U3992 ( .A1(n5046), .A2(n3548), .B1(n3477), .B2(n5026), .ZN(n3464)
         );
  XNOR2_X1 U3993 ( .A(n3463), .B(n3464), .ZN(n5030) );
  INV_X1 U3994 ( .A(n3463), .ZN(n3465) );
  NAND2_X1 U3995 ( .A1(n3465), .A2(n3464), .ZN(n3466) );
  INV_X1 U3996 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U3997 ( .A1(n3468), .A2(n4698), .ZN(n3469) );
  NAND2_X1 U3998 ( .A1(n3484), .A2(n3469), .ZN(n5053) );
  OR2_X1 U3999 ( .A1(n3603), .A2(n5053), .ZN(n3473) );
  NAND2_X1 U4000 ( .A1(n3604), .A2(REG2_REG_20__SCAN_IN), .ZN(n3472) );
  NAND2_X1 U4001 ( .A1(n2800), .A2(REG1_REG_20__SCAN_IN), .ZN(n3471) );
  NAND2_X1 U4002 ( .A1(n3774), .A2(REG0_REG_20__SCAN_IN), .ZN(n3470) );
  NAND4_X1 U4003 ( .A1(n3473), .A2(n3472), .A3(n3471), .A4(n3470), .ZN(n4279)
         );
  NAND2_X1 U4004 ( .A1(n4279), .A2(n3477), .ZN(n3475) );
  NAND2_X1 U4005 ( .A1(n2261), .A2(DATAI_20_), .ZN(n4057) );
  OR2_X1 U4006 ( .A1(n4057), .A2(n3598), .ZN(n3474) );
  NAND2_X1 U4007 ( .A1(n3475), .A2(n3474), .ZN(n3476) );
  XNOR2_X1 U4008 ( .A(n3476), .B(n3596), .ZN(n3480) );
  NAND2_X1 U4009 ( .A1(n4279), .A2(n3548), .ZN(n3479) );
  OR2_X1 U4010 ( .A1(n4057), .A2(n3533), .ZN(n3478) );
  NAND2_X1 U4011 ( .A1(n3479), .A2(n3478), .ZN(n3481) );
  INV_X1 U4012 ( .A(n3480), .ZN(n3483) );
  INV_X1 U4013 ( .A(n3481), .ZN(n3482) );
  NAND2_X1 U4014 ( .A1(n3483), .A2(n3482), .ZN(n5041) );
  NAND2_X1 U4015 ( .A1(n3484), .A2(n4686), .ZN(n3485) );
  NAND2_X1 U4016 ( .A1(n3499), .A2(n3485), .ZN(n4247) );
  NAND2_X1 U4017 ( .A1(n3604), .A2(REG2_REG_21__SCAN_IN), .ZN(n3487) );
  NAND2_X1 U4018 ( .A1(n2800), .A2(REG1_REG_21__SCAN_IN), .ZN(n3486) );
  AND2_X1 U4019 ( .A1(n3487), .A2(n3486), .ZN(n3489) );
  NAND2_X1 U4020 ( .A1(n3774), .A2(REG0_REG_21__SCAN_IN), .ZN(n3488) );
  NAND2_X1 U4021 ( .A1(n5039), .A2(n3477), .ZN(n3491) );
  NAND2_X1 U4022 ( .A1(n2261), .A2(DATAI_21_), .ZN(n4246) );
  OR2_X1 U4023 ( .A1(n4246), .A2(n3598), .ZN(n3490) );
  NAND2_X1 U4024 ( .A1(n3491), .A2(n3490), .ZN(n3492) );
  XNOR2_X1 U4025 ( .A(n3492), .B(n3566), .ZN(n3494) );
  NOR2_X1 U4026 ( .A1(n4246), .A2(n3533), .ZN(n3493) );
  AOI21_X1 U4027 ( .B1(n5039), .B2(n3548), .A(n3493), .ZN(n3495) );
  NAND2_X1 U4028 ( .A1(n3494), .A2(n3495), .ZN(n3660) );
  INV_X1 U4029 ( .A(n3494), .ZN(n3497) );
  INV_X1 U4030 ( .A(n3495), .ZN(n3496) );
  NAND2_X1 U4031 ( .A1(n3497), .A2(n3496), .ZN(n3661) );
  INV_X1 U4032 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4505) );
  INV_X1 U4033 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3726) );
  NAND2_X1 U4034 ( .A1(n3499), .A2(n3726), .ZN(n3500) );
  NAND2_X1 U4035 ( .A1(n3509), .A2(n3500), .ZN(n4228) );
  OR2_X1 U4036 ( .A1(n4228), .A2(n3603), .ZN(n3502) );
  AOI22_X1 U4037 ( .A1(n3604), .A2(REG2_REG_22__SCAN_IN), .B1(n2800), .B2(
        REG1_REG_22__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U4038 ( .A1(n4242), .A2(n3477), .ZN(n3504) );
  NAND2_X1 U4039 ( .A1(n2261), .A2(DATAI_22_), .ZN(n4221) );
  OR2_X1 U4040 ( .A1(n4221), .A2(n3598), .ZN(n3503) );
  NAND2_X1 U4041 ( .A1(n3504), .A2(n3503), .ZN(n3505) );
  XNOR2_X1 U4042 ( .A(n3505), .B(n3566), .ZN(n3508) );
  NOR2_X1 U40430 ( .A1(n4221), .A2(n3533), .ZN(n3506) );
  AOI21_X1 U4044 ( .B1(n4242), .B2(n3548), .A(n3506), .ZN(n3507) );
  XNOR2_X1 U4045 ( .A(n3508), .B(n3507), .ZN(n3725) );
  INV_X1 U4046 ( .A(n3644), .ZN(n3518) );
  NAND2_X1 U4047 ( .A1(n3509), .A2(n4514), .ZN(n3510) );
  NAND2_X1 U4048 ( .A1(n3536), .A2(n3510), .ZN(n4215) );
  AOI22_X1 U4049 ( .A1(n3604), .A2(REG2_REG_23__SCAN_IN), .B1(n2800), .B2(
        REG1_REG_23__SCAN_IN), .ZN(n3512) );
  NAND2_X1 U4050 ( .A1(n3774), .A2(REG0_REG_23__SCAN_IN), .ZN(n3511) );
  NAND2_X1 U4051 ( .A1(n4224), .A2(n3477), .ZN(n3514) );
  NAND2_X1 U4052 ( .A1(n2261), .A2(DATAI_23_), .ZN(n4213) );
  OR2_X1 U4053 ( .A1(n4213), .A2(n3598), .ZN(n3513) );
  NAND2_X1 U4054 ( .A1(n3514), .A2(n3513), .ZN(n3515) );
  XNOR2_X1 U4055 ( .A(n3515), .B(n3566), .ZN(n3520) );
  NOR2_X1 U4056 ( .A1(n4213), .A2(n3533), .ZN(n3516) );
  AOI21_X1 U4057 ( .B1(n4224), .B2(n3548), .A(n3516), .ZN(n3519) );
  XNOR2_X1 U4058 ( .A(n3520), .B(n3519), .ZN(n3647) );
  OR2_X1 U4059 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  NAND2_X1 U4060 ( .A1(n3538), .A2(n4507), .ZN(n3523) );
  NAND2_X1 U4061 ( .A1(n3556), .A2(n3523), .ZN(n3684) );
  INV_X1 U4062 ( .A(REG0_REG_25__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4063 ( .A1(n2800), .A2(REG1_REG_25__SCAN_IN), .ZN(n3525) );
  NAND2_X1 U4064 ( .A1(n3604), .A2(REG2_REG_25__SCAN_IN), .ZN(n3524) );
  OAI211_X1 U4065 ( .C1(n3607), .C2(n3526), .A(n3525), .B(n3524), .ZN(n3527)
         );
  INV_X1 U4066 ( .A(n3527), .ZN(n3528) );
  NAND2_X1 U4067 ( .A1(n4150), .A2(n3477), .ZN(n3531) );
  NAND2_X1 U4068 ( .A1(n2261), .A2(DATAI_25_), .ZN(n4173) );
  OR2_X1 U4069 ( .A1(n4173), .A2(n3598), .ZN(n3530) );
  NAND2_X1 U4070 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  XNOR2_X1 U4071 ( .A(n3532), .B(n3566), .ZN(n3551) );
  NOR2_X1 U4072 ( .A1(n4173), .A2(n3533), .ZN(n3534) );
  AOI21_X1 U4073 ( .B1(n4150), .B2(n3548), .A(n3534), .ZN(n3671) );
  NOR2_X1 U4074 ( .A1(n3551), .A2(n3671), .ZN(n3679) );
  INV_X1 U4075 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4076 ( .A1(n3536), .A2(n3535), .ZN(n3537) );
  NAND2_X1 U4077 ( .A1(n3538), .A2(n3537), .ZN(n4193) );
  INV_X1 U4078 ( .A(REG0_REG_24__SCAN_IN), .ZN(n3541) );
  NAND2_X1 U4079 ( .A1(n3604), .A2(REG2_REG_24__SCAN_IN), .ZN(n3540) );
  NAND2_X1 U4080 ( .A1(n2800), .A2(REG1_REG_24__SCAN_IN), .ZN(n3539) );
  OAI211_X1 U4081 ( .C1(n3541), .C2(n3607), .A(n3540), .B(n3539), .ZN(n3542)
         );
  INV_X1 U4082 ( .A(n3542), .ZN(n3543) );
  NAND2_X1 U4083 ( .A1(n4209), .A2(n3477), .ZN(n3546) );
  NAND2_X1 U4084 ( .A1(n2261), .A2(DATAI_24_), .ZN(n4100) );
  OR2_X1 U4085 ( .A1(n4100), .A2(n3598), .ZN(n3545) );
  NAND2_X1 U4086 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  XNOR2_X1 U4087 ( .A(n3547), .B(n3596), .ZN(n3674) );
  NAND2_X1 U4088 ( .A1(n4209), .A2(n3548), .ZN(n3550) );
  OR2_X1 U4089 ( .A1(n4100), .A2(n3533), .ZN(n3549) );
  NAND2_X1 U4090 ( .A1(n3550), .A2(n3549), .ZN(n3708) );
  INV_X1 U4091 ( .A(n3674), .ZN(n3676) );
  INV_X1 U4092 ( .A(n3708), .ZN(n3681) );
  AOI21_X1 U4093 ( .B1(n3676), .B2(n3681), .A(n3671), .ZN(n3553) );
  INV_X1 U4094 ( .A(n3551), .ZN(n3673) );
  NAND2_X1 U4095 ( .A1(n3671), .A2(n3681), .ZN(n3552) );
  OAI22_X1 U4096 ( .A1(n3553), .A2(n3673), .B1(n3674), .B2(n3552), .ZN(n3554)
         );
  INV_X1 U4097 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3747) );
  NAND2_X1 U4098 ( .A1(n3556), .A2(n3747), .ZN(n3557) );
  NAND2_X1 U4099 ( .A1(n4155), .A2(n2797), .ZN(n3563) );
  INV_X1 U4100 ( .A(REG0_REG_26__SCAN_IN), .ZN(n3560) );
  NAND2_X1 U4101 ( .A1(n3604), .A2(REG2_REG_26__SCAN_IN), .ZN(n3559) );
  NAND2_X1 U4102 ( .A1(n2800), .A2(REG1_REG_26__SCAN_IN), .ZN(n3558) );
  OAI211_X1 U4103 ( .C1(n3560), .C2(n3607), .A(n3559), .B(n3558), .ZN(n3561)
         );
  INV_X1 U4104 ( .A(n3561), .ZN(n3562) );
  NAND2_X1 U4105 ( .A1(n4065), .A2(n3477), .ZN(n3565) );
  NAND2_X1 U4106 ( .A1(n2261), .A2(DATAI_26_), .ZN(n4066) );
  OR2_X1 U4107 ( .A1(n4066), .A2(n3598), .ZN(n3564) );
  NAND2_X1 U4108 ( .A1(n3565), .A2(n3564), .ZN(n3567) );
  XNOR2_X1 U4109 ( .A(n3567), .B(n3566), .ZN(n3570) );
  NOR2_X1 U4110 ( .A1(n4066), .A2(n3533), .ZN(n3568) );
  AOI21_X1 U4111 ( .B1(n4065), .B2(n3548), .A(n3568), .ZN(n3569) );
  NOR2_X1 U4112 ( .A1(n3570), .A2(n3569), .ZN(n3745) );
  NAND2_X1 U4113 ( .A1(n3570), .A2(n3569), .ZN(n3743) );
  INV_X1 U4114 ( .A(n3572), .ZN(n3571) );
  NAND2_X1 U4115 ( .A1(n3571), .A2(REG3_REG_27__SCAN_IN), .ZN(n3587) );
  INV_X1 U4116 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U4117 ( .A1(n3572), .A2(n4671), .ZN(n3573) );
  NAND2_X1 U4118 ( .A1(n3587), .A2(n3573), .ZN(n3628) );
  INV_X1 U4119 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3576) );
  NAND2_X1 U4120 ( .A1(n3604), .A2(REG2_REG_27__SCAN_IN), .ZN(n3575) );
  NAND2_X1 U4121 ( .A1(n2800), .A2(REG1_REG_27__SCAN_IN), .ZN(n3574) );
  OAI211_X1 U4122 ( .C1(n3576), .C2(n3607), .A(n3575), .B(n3574), .ZN(n3577)
         );
  INV_X1 U4123 ( .A(n3577), .ZN(n3578) );
  NAND2_X1 U4124 ( .A1(n2261), .A2(DATAI_27_), .ZN(n4129) );
  OAI22_X1 U4125 ( .A1(n4152), .A2(n3533), .B1(n4129), .B2(n3598), .ZN(n3580)
         );
  XNOR2_X1 U4126 ( .A(n3580), .B(n3596), .ZN(n3582) );
  OAI22_X1 U4127 ( .A1(n4152), .A2(n3595), .B1(n4129), .B2(n3533), .ZN(n3581)
         );
  XNOR2_X1 U4128 ( .A(n3582), .B(n3581), .ZN(n3627) );
  INV_X1 U4129 ( .A(n3581), .ZN(n3584) );
  INV_X1 U4130 ( .A(n3582), .ZN(n3583) );
  INV_X1 U4131 ( .A(n3587), .ZN(n3585) );
  NAND2_X1 U4132 ( .A1(n3585), .A2(REG3_REG_28__SCAN_IN), .ZN(n4098) );
  INV_X1 U4133 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3586) );
  NAND2_X1 U4134 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  NAND2_X1 U4135 ( .A1(n4098), .A2(n3588), .ZN(n4120) );
  INV_X1 U4136 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3591) );
  NAND2_X1 U4137 ( .A1(n2800), .A2(REG1_REG_28__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4138 ( .A1(n3604), .A2(REG2_REG_28__SCAN_IN), .ZN(n3589) );
  OAI211_X1 U4139 ( .C1(n3607), .C2(n3591), .A(n3590), .B(n3589), .ZN(n3592)
         );
  INV_X1 U4140 ( .A(n3592), .ZN(n3593) );
  NAND2_X1 U4141 ( .A1(n2261), .A2(DATAI_28_), .ZN(n4119) );
  OAI22_X1 U4142 ( .A1(n4128), .A2(n3595), .B1(n3533), .B2(n4119), .ZN(n3597)
         );
  XNOR2_X1 U4143 ( .A(n3597), .B(n3596), .ZN(n3600) );
  OAI22_X1 U4144 ( .A1(n4128), .A2(n3533), .B1(n3598), .B2(n4119), .ZN(n3599)
         );
  XNOR2_X1 U4145 ( .A(n3600), .B(n3599), .ZN(n3601) );
  XNOR2_X1 U4146 ( .A(n3602), .B(n3601), .ZN(n3615) );
  OR2_X1 U4147 ( .A1(n4098), .A2(n3603), .ZN(n3611) );
  INV_X1 U4148 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3608) );
  NAND2_X1 U4149 ( .A1(n3604), .A2(REG2_REG_29__SCAN_IN), .ZN(n3606) );
  NAND2_X1 U4150 ( .A1(n2800), .A2(REG1_REG_29__SCAN_IN), .ZN(n3605) );
  OAI211_X1 U4151 ( .C1(n3608), .C2(n3607), .A(n3606), .B(n3605), .ZN(n3609)
         );
  INV_X1 U4152 ( .A(n3609), .ZN(n3610) );
  AOI22_X1 U4153 ( .A1(n5040), .A2(n4111), .B1(n4067), .B2(n5045), .ZN(n3613)
         );
  INV_X1 U4154 ( .A(n4119), .ZN(n4069) );
  AOI22_X1 U4155 ( .A1(n5050), .A2(n4069), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3612) );
  OAI211_X1 U4156 ( .C1(n5054), .C2(n4120), .A(n3613), .B(n3612), .ZN(n3614)
         );
  AOI21_X1 U4157 ( .B1(n3615), .B2(n5048), .A(n3614), .ZN(n3616) );
  INV_X1 U4158 ( .A(n3616), .ZN(U3217) );
  OAI211_X1 U4159 ( .C1(n3617), .C2(n3619), .A(n3618), .B(n5048), .ZN(n3625)
         );
  AOI22_X1 U4160 ( .A1(n5040), .A2(n4943), .B1(n5045), .B2(n3928), .ZN(n3624)
         );
  NOR2_X1 U4161 ( .A1(n3748), .A2(n4940), .ZN(n3620) );
  AOI211_X1 U4162 ( .C1(n3622), .C2(n3750), .A(n3621), .B(n3620), .ZN(n3623)
         );
  NAND3_X1 U4163 ( .A1(n3625), .A2(n3624), .A3(n3623), .ZN(U3210) );
  XNOR2_X1 U4164 ( .A(n3626), .B(n3627), .ZN(n3632) );
  AOI22_X1 U4165 ( .A1(n4070), .A2(n5040), .B1(n5045), .B2(n4065), .ZN(n3631)
         );
  INV_X1 U4166 ( .A(n3628), .ZN(n4137) );
  OAI22_X1 U4167 ( .A1(n3748), .A2(n4129), .B1(STATE_REG_SCAN_IN), .B2(n4671), 
        .ZN(n3629) );
  AOI21_X1 U4168 ( .B1(n4137), .B2(n3750), .A(n3629), .ZN(n3630) );
  OAI211_X1 U4169 ( .C1(n3632), .C2(n3753), .A(n3631), .B(n3630), .ZN(U3211)
         );
  OR2_X1 U4170 ( .A1(n3719), .A2(n3715), .ZN(n3633) );
  NAND2_X1 U4171 ( .A1(n3634), .A2(n3633), .ZN(n3637) );
  NOR2_X1 U4172 ( .A1(n2553), .A2(n3635), .ZN(n3636) );
  XNOR2_X1 U4173 ( .A(n3637), .B(n3636), .ZN(n3643) );
  NAND2_X1 U4174 ( .A1(n5050), .A2(n4378), .ZN(n3638) );
  NAND2_X1 U4175 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n3944) );
  NAND2_X1 U4176 ( .A1(n3638), .A2(n3944), .ZN(n3641) );
  INV_X1 U4177 ( .A(n4329), .ZN(n4371) );
  INV_X1 U4178 ( .A(n4373), .ZN(n3639) );
  OAI22_X1 U4179 ( .A1(n5032), .A2(n4371), .B1(n3639), .B2(n4991), .ZN(n3640)
         );
  AOI211_X1 U4180 ( .C1(n4380), .C2(n3750), .A(n3641), .B(n3640), .ZN(n3642)
         );
  OAI21_X1 U4181 ( .B1(n3643), .B2(n3753), .A(n3642), .ZN(U3212) );
  INV_X1 U4182 ( .A(n3645), .ZN(n3646) );
  AOI211_X1 U4183 ( .C1(n3647), .C2(n3644), .A(n3753), .B(n3646), .ZN(n3651)
         );
  AOI22_X1 U4184 ( .A1(n5040), .A2(n4209), .B1(n5045), .B2(n4242), .ZN(n3649)
         );
  INV_X1 U4185 ( .A(n4213), .ZN(n4060) );
  AOI22_X1 U4186 ( .A1(n5050), .A2(n4060), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3648) );
  OAI211_X1 U4187 ( .C1(n5054), .C2(n4215), .A(n3649), .B(n3648), .ZN(n3650)
         );
  OR2_X1 U4188 ( .A1(n3651), .A2(n3650), .ZN(U3213) );
  OAI211_X1 U4189 ( .C1(n3654), .C2(n3653), .A(n3652), .B(n5048), .ZN(n3659)
         );
  AOI22_X1 U4190 ( .A1(n5050), .A2(n3656), .B1(n3655), .B2(REG3_REG_1__SCAN_IN), .ZN(n3658) );
  AOI22_X1 U4191 ( .A1(n5040), .A2(n3931), .B1(n5045), .B2(n2907), .ZN(n3657)
         );
  NAND3_X1 U4192 ( .A1(n3659), .A2(n3658), .A3(n3657), .ZN(U3219) );
  NAND2_X1 U4193 ( .A1(n3661), .A2(n3660), .ZN(n3664) );
  INV_X1 U4194 ( .A(n5041), .ZN(n3662) );
  OAI21_X1 U4195 ( .B1(n5043), .B2(n3662), .A(n5042), .ZN(n3663) );
  XOR2_X1 U4196 ( .A(n3664), .B(n3663), .Z(n3669) );
  AOI22_X1 U4197 ( .A1(n5040), .A2(n4242), .B1(n5045), .B2(n4279), .ZN(n3668)
         );
  INV_X1 U4198 ( .A(n4247), .ZN(n3666) );
  OAI22_X1 U4199 ( .A1(n3748), .A2(n4246), .B1(STATE_REG_SCAN_IN), .B2(n4686), 
        .ZN(n3665) );
  AOI21_X1 U4200 ( .B1(n3666), .B2(n3750), .A(n3665), .ZN(n3667) );
  OAI211_X1 U4201 ( .C1(n3669), .C2(n3753), .A(n3668), .B(n3667), .ZN(U3220)
         );
  INV_X1 U4202 ( .A(n3671), .ZN(n3672) );
  NOR2_X1 U4203 ( .A1(n3673), .A2(n3672), .ZN(n3678) );
  INV_X1 U4204 ( .A(n3678), .ZN(n3683) );
  NAND2_X1 U4205 ( .A1(n3677), .A2(n3676), .ZN(n3707) );
  OAI21_X1 U4206 ( .B1(n3679), .B2(n3678), .A(n3707), .ZN(n3680) );
  AOI21_X1 U4207 ( .B1(n3681), .B2(n3706), .A(n3680), .ZN(n3682) );
  AOI21_X1 U4208 ( .B1(n2533), .B2(n3683), .A(n3682), .ZN(n3688) );
  AOI22_X1 U4209 ( .A1(n4065), .A2(n5040), .B1(n5045), .B2(n4209), .ZN(n3687)
         );
  INV_X1 U4210 ( .A(n3684), .ZN(n4174) );
  OAI22_X1 U4211 ( .A1(n3748), .A2(n4173), .B1(STATE_REG_SCAN_IN), .B2(n4507), 
        .ZN(n3685) );
  AOI21_X1 U4212 ( .B1(n4174), .B2(n3750), .A(n3685), .ZN(n3686) );
  OAI211_X1 U4213 ( .C1(n3688), .C2(n3753), .A(n3687), .B(n3686), .ZN(U3222)
         );
  XOR2_X1 U4214 ( .A(n3690), .B(n3689), .Z(n3696) );
  AOI22_X1 U4215 ( .A1(n5040), .A2(n4293), .B1(n5045), .B2(n4329), .ZN(n3695)
         );
  INV_X1 U4216 ( .A(REG3_REG_16__SCAN_IN), .ZN(n3691) );
  NOR2_X1 U4217 ( .A1(STATE_REG_SCAN_IN), .A2(n3691), .ZN(n4868) );
  INV_X1 U4218 ( .A(n4328), .ZN(n4336) );
  NOR2_X1 U4219 ( .A1(n3748), .A2(n4336), .ZN(n3692) );
  AOI211_X1 U4220 ( .C1(n3693), .C2(n3750), .A(n4868), .B(n3692), .ZN(n3694)
         );
  OAI211_X1 U4221 ( .C1(n3696), .C2(n3753), .A(n3695), .B(n3694), .ZN(U3223)
         );
  XNOR2_X1 U4222 ( .A(n3699), .B(n3698), .ZN(n3700) );
  XNOR2_X1 U4223 ( .A(n3697), .B(n3700), .ZN(n3704) );
  AOI22_X1 U4224 ( .A1(n5040), .A2(n5027), .B1(n5045), .B2(n4314), .ZN(n3702)
         );
  INV_X1 U4225 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4692) );
  NOR2_X1 U4226 ( .A1(STATE_REG_SCAN_IN), .A2(n4692), .ZN(n4009) );
  AOI21_X1 U4227 ( .B1(n5050), .B2(n4317), .A(n4009), .ZN(n3701) );
  OAI211_X1 U4228 ( .C1(n5054), .C2(n4320), .A(n3702), .B(n3701), .ZN(n3703)
         );
  AOI21_X1 U4229 ( .B1(n3704), .B2(n5048), .A(n3703), .ZN(n3705) );
  INV_X1 U4230 ( .A(n3705), .ZN(U3225) );
  NAND2_X1 U4231 ( .A1(n3707), .A2(n3706), .ZN(n3709) );
  XNOR2_X1 U4232 ( .A(n3709), .B(n3708), .ZN(n3713) );
  AOI22_X1 U4233 ( .A1(n4150), .A2(n5040), .B1(n5045), .B2(n4224), .ZN(n3711)
         );
  INV_X1 U4234 ( .A(n4100), .ZN(n4191) );
  AOI22_X1 U4235 ( .A1(n5050), .A2(n4191), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3710) );
  OAI211_X1 U4236 ( .C1(n5054), .C2(n4193), .A(n3711), .B(n3710), .ZN(n3712)
         );
  INV_X1 U4237 ( .A(n3714), .ZN(U3226) );
  INV_X1 U4238 ( .A(n3715), .ZN(n3717) );
  XNOR2_X1 U4239 ( .A(n3717), .B(n3716), .ZN(n3718) );
  XNOR2_X1 U4240 ( .A(n3719), .B(n3718), .ZN(n3723) );
  AOI22_X1 U4241 ( .A1(n5040), .A2(n4350), .B1(n5045), .B2(n4392), .ZN(n3722)
         );
  NOR2_X1 U4242 ( .A1(STATE_REG_SCAN_IN), .A2(n4699), .ZN(n4860) );
  INV_X1 U4243 ( .A(n4399), .ZN(n3756) );
  NOR2_X1 U4244 ( .A1(n3748), .A2(n3756), .ZN(n3720) );
  AOI211_X1 U4245 ( .C1(n4400), .C2(n3750), .A(n4860), .B(n3720), .ZN(n3721)
         );
  OAI211_X1 U4246 ( .C1(n3723), .C2(n3753), .A(n3722), .B(n3721), .ZN(U3231)
         );
  XOR2_X1 U4247 ( .A(n3725), .B(n3724), .Z(n3731) );
  AOI22_X1 U4248 ( .A1(n5040), .A2(n4224), .B1(n5045), .B2(n5039), .ZN(n3730)
         );
  INV_X1 U4249 ( .A(n4228), .ZN(n3728) );
  OAI22_X1 U4250 ( .A1(n3748), .A2(n4221), .B1(STATE_REG_SCAN_IN), .B2(n3726), 
        .ZN(n3727) );
  AOI21_X1 U4251 ( .B1(n3728), .B2(n3750), .A(n3727), .ZN(n3729) );
  OAI211_X1 U4252 ( .C1(n3731), .C2(n3753), .A(n3730), .B(n3729), .ZN(U3232)
         );
  INV_X1 U4253 ( .A(n3733), .ZN(n3735) );
  NAND2_X1 U4254 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  XNOR2_X1 U4255 ( .A(n3732), .B(n3736), .ZN(n3741) );
  INV_X1 U4256 ( .A(n4303), .ZN(n3739) );
  AOI22_X1 U4257 ( .A1(n5040), .A2(n5046), .B1(n5045), .B2(n4293), .ZN(n3738)
         );
  AND2_X1 U4258 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4024) );
  AOI21_X1 U4259 ( .B1(n5050), .B2(n3761), .A(n4024), .ZN(n3737) );
  OAI211_X1 U4260 ( .C1(n5054), .C2(n3739), .A(n3738), .B(n3737), .ZN(n3740)
         );
  AOI21_X1 U4261 ( .B1(n3741), .B2(n5048), .A(n3740), .ZN(n3742) );
  INV_X1 U4262 ( .A(n3742), .ZN(U3235) );
  INV_X1 U4263 ( .A(n3743), .ZN(n3744) );
  NOR2_X1 U4264 ( .A1(n3745), .A2(n3744), .ZN(n3746) );
  XNOR2_X1 U4265 ( .A(n3670), .B(n3746), .ZN(n3754) );
  AOI22_X1 U4266 ( .A1(n4067), .A2(n5040), .B1(n5045), .B2(n4150), .ZN(n3752)
         );
  OAI22_X1 U4267 ( .A1(n3748), .A2(n4066), .B1(STATE_REG_SCAN_IN), .B2(n3747), 
        .ZN(n3749) );
  AOI21_X1 U4268 ( .B1(n4155), .B2(n3750), .A(n3749), .ZN(n3751) );
  OAI211_X1 U4269 ( .C1(n3754), .C2(n3753), .A(n3752), .B(n3751), .ZN(U3237)
         );
  NAND2_X1 U4270 ( .A1(n4150), .A2(n4173), .ZN(n3863) );
  NAND2_X1 U4271 ( .A1(n4209), .A2(n4100), .ZN(n4163) );
  OR2_X1 U4272 ( .A1(n4242), .A2(n4221), .ZN(n4202) );
  OR2_X1 U4273 ( .A1(n5039), .A2(n4246), .ZN(n4199) );
  NAND2_X1 U4274 ( .A1(n4202), .A2(n4199), .ZN(n4083) );
  NAND2_X1 U4275 ( .A1(n4373), .A2(n3756), .ZN(n3755) );
  NOR2_X1 U4276 ( .A1(n4373), .A2(n3756), .ZN(n3757) );
  AOI21_X1 U4277 ( .B1(n3833), .B2(n4387), .A(n3757), .ZN(n3836) );
  INV_X1 U4278 ( .A(n4350), .ZN(n4992) );
  NAND2_X1 U4279 ( .A1(n4992), .A2(n4378), .ZN(n4076) );
  NAND2_X1 U4280 ( .A1(n4371), .A2(n4996), .ZN(n3894) );
  NAND2_X1 U4281 ( .A1(n4076), .A2(n3894), .ZN(n3832) );
  NAND2_X1 U4282 ( .A1(n4350), .A2(n4370), .ZN(n3883) );
  INV_X1 U4283 ( .A(n3883), .ZN(n3821) );
  NAND2_X1 U4284 ( .A1(n4329), .A2(n4351), .ZN(n4077) );
  INV_X1 U4285 ( .A(n4077), .ZN(n3822) );
  AOI21_X1 U4286 ( .B1(n3821), .B2(n3894), .A(n3822), .ZN(n3840) );
  AND2_X1 U4287 ( .A1(n4314), .A2(n4336), .ZN(n3844) );
  OAI211_X1 U4288 ( .C1(n4075), .C2(n3832), .A(n3840), .B(n4078), .ZN(n3759)
         );
  INV_X1 U4289 ( .A(n4314), .ZN(n4993) );
  NAND2_X1 U4290 ( .A1(n4993), .A2(n4328), .ZN(n3869) );
  AND2_X1 U4291 ( .A1(n3759), .A2(n3869), .ZN(n3766) );
  NAND2_X1 U4292 ( .A1(n5027), .A2(n4300), .ZN(n4276) );
  NAND2_X1 U4293 ( .A1(n5046), .A2(n4284), .ZN(n3760) );
  AND2_X1 U4294 ( .A1(n4276), .A2(n3760), .ZN(n3763) );
  INV_X1 U4295 ( .A(n4317), .ZN(n4311) );
  NAND2_X1 U4296 ( .A1(n4293), .A2(n4311), .ZN(n4270) );
  NAND2_X1 U4297 ( .A1(n3763), .A2(n4270), .ZN(n4079) );
  NAND2_X1 U4298 ( .A1(n4279), .A2(n4057), .ZN(n3888) );
  INV_X1 U4299 ( .A(n3888), .ZN(n4081) );
  OR2_X1 U4300 ( .A1(n4079), .A2(n4081), .ZN(n3843) );
  INV_X1 U4301 ( .A(n5027), .ZN(n4312) );
  NAND2_X1 U4302 ( .A1(n4312), .A2(n3761), .ZN(n4274) );
  INV_X1 U4303 ( .A(n4293), .ZN(n4332) );
  NAND2_X1 U4304 ( .A1(n4332), .A2(n4317), .ZN(n4272) );
  NAND2_X1 U4305 ( .A1(n4274), .A2(n4272), .ZN(n3764) );
  NOR2_X1 U4306 ( .A1(n5046), .A2(n4284), .ZN(n3762) );
  AOI21_X1 U4307 ( .B1(n3764), .B2(n3763), .A(n3762), .ZN(n4254) );
  INV_X1 U4308 ( .A(n4279), .ZN(n5031) );
  NAND2_X1 U4309 ( .A1(n5031), .A2(n5049), .ZN(n3889) );
  NAND2_X1 U4310 ( .A1(n4254), .A2(n3889), .ZN(n3765) );
  NAND2_X1 U4311 ( .A1(n3765), .A2(n3888), .ZN(n4080) );
  OAI21_X1 U4312 ( .B1(n3766), .B2(n3843), .A(n4080), .ZN(n3768) );
  NAND2_X1 U4313 ( .A1(n4224), .A2(n4213), .ZN(n3870) );
  NAND2_X1 U4314 ( .A1(n4242), .A2(n4221), .ZN(n4204) );
  NAND2_X1 U4315 ( .A1(n3870), .A2(n4204), .ZN(n3847) );
  NAND2_X1 U4316 ( .A1(n5039), .A2(n4246), .ZN(n3865) );
  INV_X1 U4317 ( .A(n3865), .ZN(n4200) );
  AND2_X1 U4318 ( .A1(n4202), .A2(n4200), .ZN(n3767) );
  NOR2_X1 U4319 ( .A1(n3847), .A2(n3767), .ZN(n4082) );
  OAI21_X1 U4320 ( .B1(n4083), .B2(n3768), .A(n4082), .ZN(n3769) );
  OR2_X1 U4321 ( .A1(n4209), .A2(n4100), .ZN(n3868) );
  OR2_X1 U4322 ( .A1(n4224), .A2(n4213), .ZN(n4181) );
  NAND2_X1 U4323 ( .A1(n3769), .A2(n4084), .ZN(n3781) );
  NAND2_X1 U4324 ( .A1(n4128), .A2(n4069), .ZN(n4090) );
  NAND2_X1 U4325 ( .A1(n4152), .A2(n4134), .ZN(n3782) );
  NAND2_X1 U4326 ( .A1(n4090), .A2(n3782), .ZN(n3786) );
  INV_X1 U4327 ( .A(n4111), .ZN(n3770) );
  NAND2_X1 U4328 ( .A1(n2261), .A2(DATAI_29_), .ZN(n4101) );
  INV_X1 U4329 ( .A(n4101), .ZN(n4093) );
  NAND2_X1 U4330 ( .A1(n3770), .A2(n4093), .ZN(n3780) );
  INV_X1 U4331 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4332 ( .A1(n2800), .A2(REG1_REG_30__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4333 ( .A1(n3774), .A2(REG0_REG_30__SCAN_IN), .ZN(n3771) );
  OAI211_X1 U4334 ( .C1(n2802), .C2(n3773), .A(n3772), .B(n3771), .ZN(n4094)
         );
  NAND2_X1 U4335 ( .A1(n2261), .A2(DATAI_30_), .ZN(n4407) );
  OR2_X1 U4336 ( .A1(n4094), .A2(n4407), .ZN(n3779) );
  INV_X1 U4337 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3777) );
  NAND2_X1 U4338 ( .A1(n2800), .A2(REG1_REG_31__SCAN_IN), .ZN(n3776) );
  NAND2_X1 U4339 ( .A1(n3774), .A2(REG0_REG_31__SCAN_IN), .ZN(n3775) );
  OAI211_X1 U4340 ( .C1(n2802), .C2(n3777), .A(n3776), .B(n3775), .ZN(n4410)
         );
  NAND2_X1 U4341 ( .A1(n2261), .A2(DATAI_31_), .ZN(n4408) );
  NAND2_X1 U4342 ( .A1(n4410), .A2(n4408), .ZN(n3855) );
  AND2_X1 U4343 ( .A1(n3779), .A2(n3855), .ZN(n3893) );
  NAND2_X1 U4344 ( .A1(n3780), .A2(n3893), .ZN(n3784) );
  AOI211_X1 U4345 ( .C1(n4085), .C2(n3781), .A(n3786), .B(n3784), .ZN(n3788)
         );
  NOR2_X1 U4346 ( .A1(n4065), .A2(n4066), .ZN(n3862) );
  NOR2_X1 U4347 ( .A1(n4150), .A2(n4173), .ZN(n4145) );
  NOR2_X1 U4348 ( .A1(n3862), .A2(n4145), .ZN(n4087) );
  INV_X1 U4349 ( .A(n3782), .ZN(n4088) );
  NOR2_X1 U4350 ( .A1(n4152), .A2(n4134), .ZN(n3853) );
  NAND2_X1 U4351 ( .A1(n4111), .A2(n4101), .ZN(n3783) );
  NAND2_X1 U4352 ( .A1(n4070), .A2(n4119), .ZN(n4089) );
  NAND2_X1 U4353 ( .A1(n4065), .A2(n4066), .ZN(n3851) );
  NAND4_X1 U4354 ( .A1(n4126), .A2(n3783), .A3(n4089), .A4(n3851), .ZN(n3787)
         );
  NAND2_X1 U4355 ( .A1(n3783), .A2(n4089), .ZN(n3852) );
  INV_X1 U4356 ( .A(n3852), .ZN(n3785) );
  AOI21_X1 U4357 ( .B1(n3786), .B2(n3785), .A(n3784), .ZN(n3854) );
  AOI22_X1 U4358 ( .A1(n3788), .A2(n4087), .B1(n3787), .B2(n3854), .ZN(n3792)
         );
  NOR2_X1 U4359 ( .A1(n4410), .A2(n4407), .ZN(n3791) );
  OR2_X1 U4360 ( .A1(n4410), .A2(n4408), .ZN(n3790) );
  NAND2_X1 U4361 ( .A1(n4094), .A2(n4407), .ZN(n3789) );
  NAND2_X1 U4362 ( .A1(n3790), .A2(n3789), .ZN(n3856) );
  INV_X1 U4363 ( .A(n3856), .ZN(n3874) );
  OAI22_X1 U4364 ( .A1(n3792), .A2(n3791), .B1(n3874), .B2(n4408), .ZN(n3793)
         );
  XNOR2_X1 U4365 ( .A(n3793), .B(n4936), .ZN(n3916) );
  INV_X1 U4366 ( .A(n3794), .ZN(n3915) );
  NAND2_X1 U4367 ( .A1(n2907), .A2(n2314), .ZN(n3866) );
  OAI211_X1 U4368 ( .C1(n3798), .C2(n3797), .A(n3866), .B(n3796), .ZN(n3800)
         );
  NAND3_X1 U4369 ( .A1(n3800), .A2(n3799), .A3(n2912), .ZN(n3803) );
  NAND3_X1 U4370 ( .A1(n3803), .A2(n3802), .A3(n3801), .ZN(n3806) );
  NAND3_X1 U4371 ( .A1(n3806), .A2(n3805), .A3(n3804), .ZN(n3809) );
  NAND4_X1 U4372 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3825), .ZN(n3812)
         );
  NAND3_X1 U4373 ( .A1(n3812), .A2(n3811), .A3(n3810), .ZN(n3813) );
  NAND3_X1 U4374 ( .A1(n3813), .A2(n3823), .A3(n3826), .ZN(n3816) );
  NAND3_X1 U4375 ( .A1(n3816), .A2(n3815), .A3(n3814), .ZN(n3842) );
  AND2_X1 U4376 ( .A1(n3818), .A2(n3817), .ZN(n3819) );
  NAND2_X1 U4377 ( .A1(n3833), .A2(n3819), .ZN(n3837) );
  NOR4_X1 U4378 ( .A1(n3837), .A2(n3822), .A3(n3821), .A4(n3820), .ZN(n3841)
         );
  NOR2_X1 U4379 ( .A1(n2425), .A2(n3824), .ZN(n3828) );
  NAND4_X1 U4380 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3830)
         );
  AND2_X1 U4381 ( .A1(n3830), .A2(n3829), .ZN(n3838) );
  INV_X1 U4382 ( .A(n3831), .ZN(n3834) );
  AOI21_X1 U4383 ( .B1(n3834), .B2(n3833), .A(n3832), .ZN(n3835) );
  OAI211_X1 U4384 ( .C1(n3838), .C2(n3837), .A(n3836), .B(n3835), .ZN(n3839)
         );
  AOI22_X1 U4385 ( .A1(n3842), .A2(n3841), .B1(n3840), .B2(n3839), .ZN(n3845)
         );
  AOI211_X1 U4386 ( .C1(n3869), .C2(n3845), .A(n3844), .B(n3843), .ZN(n3846)
         );
  AOI221_X1 U4387 ( .B1(n2414), .B2(n3865), .C1(n3846), .C2(n3865), .A(n4083), 
        .ZN(n3848) );
  OAI21_X1 U4388 ( .B1(n3848), .B2(n3847), .A(n4084), .ZN(n3849) );
  NAND2_X1 U4389 ( .A1(n3849), .A2(n4085), .ZN(n3850) );
  NAND2_X1 U4390 ( .A1(n3850), .A2(n4087), .ZN(n3860) );
  NOR4_X1 U4391 ( .A1(n3853), .A2(n4086), .A3(n3852), .A4(n3856), .ZN(n3859)
         );
  INV_X1 U4392 ( .A(n3854), .ZN(n3858) );
  NAND2_X1 U4393 ( .A1(n3856), .A2(n3855), .ZN(n3857) );
  AOI22_X1 U4394 ( .A1(n3860), .A2(n3859), .B1(n3858), .B2(n3857), .ZN(n3861)
         );
  NOR2_X1 U4395 ( .A1(n3861), .A2(n2262), .ZN(n3911) );
  INV_X1 U4396 ( .A(n3911), .ZN(n3907) );
  NAND2_X1 U4397 ( .A1(n4089), .A2(n4090), .ZN(n4110) );
  INV_X1 U4398 ( .A(n4110), .ZN(n3904) );
  XNOR2_X1 U4399 ( .A(n4111), .B(n4101), .ZN(n4092) );
  INV_X1 U4400 ( .A(n4092), .ZN(n3903) );
  INV_X1 U4401 ( .A(n4143), .ZN(n4148) );
  INV_X1 U4402 ( .A(n3863), .ZN(n3864) );
  OR2_X1 U4403 ( .A1(n3864), .A2(n4145), .ZN(n4165) );
  XNOR2_X1 U4404 ( .A(n5046), .B(n4284), .ZN(n4283) );
  NAND2_X1 U4405 ( .A1(n4199), .A2(n3865), .ZN(n4239) );
  NAND2_X1 U4406 ( .A1(n3867), .A2(n3866), .ZN(n4887) );
  NOR4_X1 U4407 ( .A1(n4165), .A2(n4283), .A3(n4239), .A4(n4887), .ZN(n3879)
         );
  NAND2_X1 U4408 ( .A1(n3868), .A2(n4163), .ZN(n4184) );
  NAND2_X1 U4409 ( .A1(n4181), .A2(n3870), .ZN(n4206) );
  NOR3_X1 U4410 ( .A1(n4206), .A2(n3872), .A3(n3871), .ZN(n3873) );
  NAND3_X1 U4411 ( .A1(n4333), .A2(n3874), .A3(n3873), .ZN(n3877) );
  AND2_X1 U4412 ( .A1(n4272), .A2(n4270), .ZN(n4309) );
  NAND2_X1 U4413 ( .A1(n4373), .A2(n4399), .ZN(n4358) );
  INV_X1 U4414 ( .A(n4358), .ZN(n3875) );
  NOR2_X1 U4415 ( .A1(n4373), .A2(n4399), .ZN(n4359) );
  OR2_X1 U4416 ( .A1(n3875), .A2(n4359), .ZN(n4390) );
  NAND2_X1 U4417 ( .A1(n4309), .A2(n4390), .ZN(n3876) );
  NOR3_X1 U4418 ( .A1(n4184), .A2(n3877), .A3(n3876), .ZN(n3878) );
  AND3_X1 U4419 ( .A1(n4148), .A2(n3879), .A3(n3878), .ZN(n3902) );
  NAND2_X1 U4420 ( .A1(n4274), .A2(n4276), .ZN(n4298) );
  INV_X1 U4421 ( .A(n4298), .ZN(n4291) );
  NAND4_X1 U4422 ( .A1(n3881), .A2(n4291), .A3(n4041), .A4(n3880), .ZN(n3887)
         );
  INV_X1 U4423 ( .A(n3882), .ZN(n3885) );
  NAND2_X1 U4424 ( .A1(n4076), .A2(n3883), .ZN(n4369) );
  INV_X1 U4425 ( .A(n4369), .ZN(n4074) );
  NAND4_X1 U4426 ( .A1(n3885), .A2(n4074), .A3(n2268), .A4(n3884), .ZN(n3886)
         );
  NOR2_X1 U4427 ( .A1(n3887), .A2(n3886), .ZN(n3898) );
  AND2_X1 U4428 ( .A1(n3889), .A2(n3888), .ZN(n4256) );
  AND4_X1 U4429 ( .A1(n3892), .A2(n4256), .A3(n3891), .A4(n3890), .ZN(n3897)
         );
  AND2_X1 U4430 ( .A1(n4937), .A2(n3893), .ZN(n3896) );
  NAND2_X1 U4431 ( .A1(n4202), .A2(n4204), .ZN(n4231) );
  NAND2_X1 U4432 ( .A1(n3894), .A2(n4077), .ZN(n4364) );
  NOR2_X1 U4433 ( .A1(n4231), .A2(n4364), .ZN(n3895) );
  NAND4_X1 U4434 ( .A1(n3898), .A2(n3897), .A3(n3896), .A4(n3895), .ZN(n3899)
         );
  NOR2_X1 U4435 ( .A1(n3900), .A2(n3899), .ZN(n3901) );
  NAND4_X1 U4436 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3909)
         );
  INV_X1 U4437 ( .A(n3909), .ZN(n3905) );
  NAND3_X1 U4438 ( .A1(n3905), .A2(n2262), .A3(n3908), .ZN(n3906) );
  NAND2_X1 U4439 ( .A1(n3907), .A2(n3906), .ZN(n3913) );
  AOI21_X1 U4440 ( .B1(n3909), .B2(n3908), .A(n2719), .ZN(n3910) );
  NOR2_X1 U4441 ( .A1(n3911), .A2(n3910), .ZN(n3912) );
  MUX2_X1 U4442 ( .A(n3913), .B(n3912), .S(n4936), .Z(n3914) );
  AOI21_X1 U4443 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3923) );
  NOR4_X1 U4444 ( .A1(n3533), .A2(n3919), .A3(n3918), .A4(n3917), .ZN(n3922)
         );
  OAI21_X1 U4445 ( .B1(n4767), .B2(n3920), .A(B_REG_SCAN_IN), .ZN(n3921) );
  OAI22_X1 U4446 ( .A1(n3923), .A2(n4767), .B1(n3922), .B2(n3921), .ZN(U3239)
         );
  MUX2_X1 U4447 ( .A(n4410), .B(DATAO_REG_31__SCAN_IN), .S(n3932), .Z(U3581)
         );
  MUX2_X1 U4448 ( .A(n4094), .B(DATAO_REG_30__SCAN_IN), .S(n3932), .Z(U3580)
         );
  MUX2_X1 U4449 ( .A(DATAO_REG_29__SCAN_IN), .B(n4111), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4450 ( .A(DATAO_REG_28__SCAN_IN), .B(n4070), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4451 ( .A(DATAO_REG_27__SCAN_IN), .B(n4067), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4452 ( .A(n4065), .B(DATAO_REG_26__SCAN_IN), .S(n3932), .Z(U3576)
         );
  MUX2_X1 U4453 ( .A(n4150), .B(DATAO_REG_25__SCAN_IN), .S(n3932), .Z(U3575)
         );
  MUX2_X1 U4454 ( .A(n4209), .B(DATAO_REG_24__SCAN_IN), .S(n3932), .Z(U3574)
         );
  MUX2_X1 U4455 ( .A(n4224), .B(DATAO_REG_23__SCAN_IN), .S(n3932), .Z(U3573)
         );
  MUX2_X1 U4456 ( .A(n4242), .B(DATAO_REG_22__SCAN_IN), .S(n3932), .Z(U3572)
         );
  MUX2_X1 U4457 ( .A(n5039), .B(DATAO_REG_21__SCAN_IN), .S(n3932), .Z(U3571)
         );
  MUX2_X1 U4458 ( .A(n4279), .B(DATAO_REG_20__SCAN_IN), .S(n3932), .Z(U3570)
         );
  MUX2_X1 U4459 ( .A(n5046), .B(DATAO_REG_19__SCAN_IN), .S(n3932), .Z(U3569)
         );
  MUX2_X1 U4460 ( .A(n5027), .B(DATAO_REG_18__SCAN_IN), .S(n3932), .Z(U3568)
         );
  MUX2_X1 U4461 ( .A(n4293), .B(DATAO_REG_17__SCAN_IN), .S(n3932), .Z(U3567)
         );
  MUX2_X1 U4462 ( .A(n4314), .B(DATAO_REG_16__SCAN_IN), .S(n3932), .Z(U3566)
         );
  MUX2_X1 U4463 ( .A(n4329), .B(DATAO_REG_15__SCAN_IN), .S(n3932), .Z(U3565)
         );
  MUX2_X1 U4464 ( .A(n4350), .B(DATAO_REG_14__SCAN_IN), .S(n3932), .Z(U3564)
         );
  MUX2_X1 U4465 ( .A(n4373), .B(DATAO_REG_13__SCAN_IN), .S(n3932), .Z(U3563)
         );
  MUX2_X1 U4466 ( .A(n4392), .B(DATAO_REG_12__SCAN_IN), .S(n3932), .Z(U3562)
         );
  MUX2_X1 U4467 ( .A(n3924), .B(DATAO_REG_11__SCAN_IN), .S(n3932), .Z(U3561)
         );
  MUX2_X1 U4468 ( .A(n3925), .B(DATAO_REG_10__SCAN_IN), .S(n3932), .Z(U3560)
         );
  MUX2_X1 U4469 ( .A(n3926), .B(DATAO_REG_9__SCAN_IN), .S(n3932), .Z(U3559) );
  MUX2_X1 U4470 ( .A(n4943), .B(DATAO_REG_8__SCAN_IN), .S(n3932), .Z(U3558) );
  MUX2_X1 U4471 ( .A(n3927), .B(DATAO_REG_7__SCAN_IN), .S(n3932), .Z(U3557) );
  MUX2_X1 U4472 ( .A(n3928), .B(DATAO_REG_6__SCAN_IN), .S(n3932), .Z(U3556) );
  MUX2_X1 U4473 ( .A(n3929), .B(DATAO_REG_5__SCAN_IN), .S(n3932), .Z(U3555) );
  MUX2_X1 U4474 ( .A(n3930), .B(DATAO_REG_4__SCAN_IN), .S(n3932), .Z(U3554) );
  MUX2_X1 U4475 ( .A(n2843), .B(DATAO_REG_3__SCAN_IN), .S(n3932), .Z(U3553) );
  MUX2_X1 U4476 ( .A(n3931), .B(DATAO_REG_2__SCAN_IN), .S(n3932), .Z(U3552) );
  MUX2_X1 U4477 ( .A(n2906), .B(DATAO_REG_1__SCAN_IN), .S(n3932), .Z(U3551) );
  MUX2_X1 U4478 ( .A(n2907), .B(DATAO_REG_0__SCAN_IN), .S(n3932), .Z(U3550) );
  AOI22_X1 U4479 ( .A1(n4869), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3943) );
  NAND2_X1 U4480 ( .A1(n4823), .A2(n4766), .ZN(n3942) );
  MUX2_X1 U4481 ( .A(n2610), .B(REG1_REG_1__SCAN_IN), .S(n4766), .Z(n3933) );
  OAI21_X1 U4482 ( .B1(n4881), .B2(n3934), .A(n3933), .ZN(n3935) );
  NAND3_X1 U4483 ( .A1(n4870), .A2(n3936), .A3(n3935), .ZN(n3941) );
  OAI211_X1 U4484 ( .C1(n3939), .C2(n3938), .A(n4847), .B(n3937), .ZN(n3940)
         );
  NAND4_X1 U4485 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(U3241)
         );
  INV_X1 U4486 ( .A(n3944), .ZN(n3945) );
  AOI21_X1 U4487 ( .B1(n4869), .B2(ADDR_REG_14__SCAN_IN), .A(n3945), .ZN(n3946) );
  INV_X1 U4488 ( .A(n3946), .ZN(n3960) );
  INV_X1 U4489 ( .A(n4759), .ZN(n3957) );
  NAND2_X1 U4490 ( .A1(n3965), .A2(REG2_REG_11__SCAN_IN), .ZN(n3954) );
  AOI22_X1 U4491 ( .A1(n3965), .A2(REG2_REG_11__SCAN_IN), .B1(n3194), .B2(
        n4970), .ZN(n4838) );
  AOI22_X1 U4492 ( .A1(n4810), .A2(REG2_REG_9__SCAN_IN), .B1(n3096), .B2(n4959), .ZN(n4818) );
  INV_X1 U4493 ( .A(n3947), .ZN(n3948) );
  NAND2_X1 U4494 ( .A1(n3948), .A2(n4760), .ZN(n3950) );
  NAND2_X1 U4495 ( .A1(n4967), .A2(n3952), .ZN(n3953) );
  NAND2_X1 U4496 ( .A1(n3953), .A2(n4824), .ZN(n4837) );
  NAND2_X1 U4497 ( .A1(n4838), .A2(n4837), .ZN(n4836) );
  NAND2_X1 U4498 ( .A1(n3967), .A2(n3955), .ZN(n3956) );
  INV_X1 U4499 ( .A(n3967), .ZN(n4980) );
  XNOR2_X1 U4500 ( .A(n3955), .B(n4980), .ZN(n4848) );
  NAND2_X1 U4501 ( .A1(REG2_REG_12__SCAN_IN), .A2(n4848), .ZN(n4846) );
  NAND2_X1 U4502 ( .A1(n3956), .A2(n4846), .ZN(n4856) );
  INV_X1 U4503 ( .A(n4852), .ZN(n4982) );
  NOR2_X1 U4504 ( .A1(n4982), .A2(n4402), .ZN(n4855) );
  AOI211_X1 U4505 ( .C1(n4382), .C2(n3958), .A(n3973), .B(n4864), .ZN(n3959)
         );
  AOI211_X1 U4506 ( .C1(n4823), .C2(n4759), .A(n3960), .B(n3959), .ZN(n3972)
         );
  INV_X1 U4507 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4976) );
  NOR2_X1 U4508 ( .A1(n4970), .A2(n4976), .ZN(n4830) );
  INV_X1 U4509 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4964) );
  AOI222_X1 U4510 ( .A1(n4813), .A2(n4959), .B1(n4813), .B2(n4964), .C1(n4959), 
        .C2(n4964), .ZN(n3963) );
  NAND2_X1 U4511 ( .A1(n4967), .A2(n3963), .ZN(n3964) );
  NOR2_X1 U4512 ( .A1(n4980), .A2(n3966), .ZN(n3968) );
  INV_X1 U4513 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4843) );
  NAND2_X1 U4514 ( .A1(n4852), .A2(REG1_REG_13__SCAN_IN), .ZN(n4851) );
  INV_X1 U4515 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4988) );
  NAND2_X1 U4516 ( .A1(n4982), .A2(n4988), .ZN(n3969) );
  NAND2_X1 U4517 ( .A1(REG1_REG_14__SCAN_IN), .A2(n3970), .ZN(n3982) );
  OAI211_X1 U4518 ( .C1(n3970), .C2(REG1_REG_14__SCAN_IN), .A(n4870), .B(n3982), .ZN(n3971) );
  NAND2_X1 U4519 ( .A1(n3972), .A2(n3971), .ZN(U3254) );
  INV_X1 U4520 ( .A(n4758), .ZN(n3991) );
  AND2_X1 U4521 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4995) );
  NAND2_X1 U4522 ( .A1(n4758), .A2(REG2_REG_15__SCAN_IN), .ZN(n4001) );
  OR2_X1 U4523 ( .A1(n4758), .A2(REG2_REG_15__SCAN_IN), .ZN(n3974) );
  NAND2_X1 U4524 ( .A1(n4001), .A2(n3974), .ZN(n3976) );
  INV_X1 U4525 ( .A(n4002), .ZN(n3975) );
  AOI211_X1 U4526 ( .C1(n3977), .C2(n3976), .A(n3975), .B(n4864), .ZN(n3978)
         );
  AOI211_X1 U4527 ( .C1(n4869), .C2(ADDR_REG_15__SCAN_IN), .A(n4995), .B(n3978), .ZN(n3989) );
  INV_X1 U4528 ( .A(n3979), .ZN(n3980) );
  NAND2_X1 U4529 ( .A1(n4759), .A2(n3980), .ZN(n3981) );
  NOR2_X1 U4530 ( .A1(n4758), .A2(REG1_REG_15__SCAN_IN), .ZN(n3983) );
  INV_X1 U4531 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5011) );
  AOI21_X1 U4532 ( .B1(n4758), .B2(n5011), .A(n3985), .ZN(n3986) );
  OAI21_X1 U4533 ( .B1(n5011), .B2(n4758), .A(n3986), .ZN(n3987) );
  NAND3_X1 U4534 ( .A1(n4870), .A2(n3990), .A3(n3987), .ZN(n3988) );
  OAI211_X1 U4535 ( .C1(n4875), .C2(n3991), .A(n3989), .B(n3988), .ZN(U3255)
         );
  INV_X1 U4536 ( .A(n4020), .ZN(n4012) );
  INV_X1 U4537 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3993) );
  OR2_X1 U4538 ( .A1(n4020), .A2(n3993), .ZN(n3995) );
  NAND2_X1 U4539 ( .A1(n4020), .A2(n3993), .ZN(n3994) );
  NAND2_X1 U4540 ( .A1(n3995), .A2(n3994), .ZN(n3997) );
  OAI21_X1 U4541 ( .B1(n2501), .B2(n3997), .A(n4014), .ZN(n3998) );
  NAND2_X1 U4542 ( .A1(n3998), .A2(n4870), .ZN(n4011) );
  INV_X1 U4543 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4321) );
  OR2_X1 U4544 ( .A1(n4020), .A2(REG2_REG_17__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U4545 ( .A1(n4020), .A2(REG2_REG_17__SCAN_IN), .ZN(n3999) );
  AND2_X1 U4546 ( .A1(n4000), .A2(n3999), .ZN(n4007) );
  NAND2_X1 U4547 ( .A1(n4004), .A2(n2485), .ZN(n4005) );
  NAND2_X1 U4548 ( .A1(n4019), .A2(n4007), .ZN(n4006) );
  AOI221_X1 U4549 ( .B1(n4007), .B2(n4006), .C1(n4019), .C2(n4006), .A(n4864), 
        .ZN(n4008) );
  AOI211_X1 U4550 ( .C1(n4869), .C2(ADDR_REG_17__SCAN_IN), .A(n4009), .B(n4008), .ZN(n4010) );
  OAI211_X1 U4551 ( .C1(n4012), .C2(n4875), .A(n4011), .B(n4010), .ZN(U3257)
         );
  INV_X1 U4552 ( .A(n4757), .ZN(n4027) );
  NAND2_X1 U4553 ( .A1(n4012), .A2(n3993), .ZN(n4013) );
  XNOR2_X1 U4554 ( .A(n4757), .B(REG1_REG_18__SCAN_IN), .ZN(n4015) );
  INV_X1 U4555 ( .A(n4015), .ZN(n4016) );
  OAI211_X1 U4556 ( .C1(n2283), .C2(n4016), .A(n4028), .B(n4870), .ZN(n4026)
         );
  INV_X1 U4557 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4018) );
  NOR2_X1 U4558 ( .A1(n4757), .A2(n4018), .ZN(n4017) );
  AOI21_X1 U4559 ( .B1(n4018), .B2(n4757), .A(n4017), .ZN(n4022) );
  AOI211_X1 U4560 ( .C1(n4022), .C2(n4021), .A(n2282), .B(n4864), .ZN(n4023)
         );
  AOI211_X1 U4561 ( .C1(n4869), .C2(ADDR_REG_18__SCAN_IN), .A(n4024), .B(n4023), .ZN(n4025) );
  OAI211_X1 U4562 ( .C1(n4027), .C2(n4875), .A(n4026), .B(n4025), .ZN(U3258)
         );
  INV_X1 U4563 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4471) );
  XNOR2_X1 U4564 ( .A(REG2_REG_19__SCAN_IN), .B(n4031), .ZN(n4032) );
  OAI22_X1 U4565 ( .A1(n4863), .A2(n4033), .B1(n4864), .B2(n4032), .ZN(n4037)
         );
  AOI22_X1 U4566 ( .A1(n4870), .A2(n4033), .B1(n4847), .B2(n4032), .ZN(n4035)
         );
  NOR2_X1 U4567 ( .A1(STATE_REG_SCAN_IN), .A2(n3452), .ZN(n5033) );
  AOI21_X1 U4568 ( .B1(n4869), .B2(ADDR_REG_19__SCAN_IN), .A(n5033), .ZN(n4038) );
  NAND2_X1 U4569 ( .A1(n4039), .A2(n4038), .ZN(U3259) );
  INV_X1 U4570 ( .A(n4065), .ZN(n4169) );
  AND2_X1 U4571 ( .A1(n4392), .A2(n4040), .ZN(n4049) );
  NOR2_X1 U4572 ( .A1(n4041), .A2(n4049), .ZN(n4043) );
  AND2_X1 U4573 ( .A1(n4043), .A2(n4042), .ZN(n4044) );
  AND2_X1 U4574 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  NAND2_X1 U4575 ( .A1(n4047), .A2(n4046), .ZN(n4053) );
  NAND2_X1 U4576 ( .A1(n4053), .A2(n4052), .ZN(n4357) );
  NAND2_X1 U4577 ( .A1(n4329), .A2(n4996), .ZN(n4055) );
  AND3_X1 U4578 ( .A1(n4369), .A2(n4055), .A3(n4358), .ZN(n4054) );
  NOR2_X1 U4579 ( .A1(n4350), .A2(n4378), .ZN(n4362) );
  AOI22_X1 U4580 ( .A1(n4362), .A2(n4055), .B1(n4371), .B2(n4351), .ZN(n4056)
         );
  AOI22_X1 U4581 ( .A1(n4299), .A2(n4298), .B1(n4300), .B2(n4312), .ZN(n4282)
         );
  INV_X1 U4582 ( .A(n5046), .ZN(n4259) );
  INV_X1 U4583 ( .A(n4246), .ZN(n4099) );
  AND2_X1 U4584 ( .A1(n5039), .A2(n4099), .ZN(n4232) );
  INV_X1 U4585 ( .A(n5039), .ZN(n4222) );
  NAND2_X1 U4586 ( .A1(n4222), .A2(n4246), .ZN(n4233) );
  INV_X1 U4587 ( .A(n4242), .ZN(n4207) );
  INV_X1 U4588 ( .A(n4224), .ZN(n4061) );
  INV_X1 U4589 ( .A(n4209), .ZN(n4063) );
  INV_X1 U4590 ( .A(n4173), .ZN(n4167) );
  INV_X1 U4591 ( .A(n4150), .ZN(n4186) );
  OAI22_X1 U4592 ( .A1(n4161), .A2(n4064), .B1(n4186), .B2(n4173), .ZN(n4144)
         );
  NAND2_X1 U4593 ( .A1(n4067), .A2(n4134), .ZN(n4068) );
  NAND2_X1 U4594 ( .A1(n4108), .A2(n4110), .ZN(n4072) );
  NAND2_X1 U4595 ( .A1(n4072), .A2(n4071), .ZN(n4073) );
  XNOR2_X1 U4596 ( .A(n4073), .B(n3903), .ZN(n4421) );
  INV_X1 U4597 ( .A(n4421), .ZN(n4107) );
  NAND2_X1 U4598 ( .A1(n4345), .A2(n4077), .ZN(n4327) );
  XOR2_X1 U4599 ( .A(n4092), .B(n4091), .Z(n4097) );
  AOI21_X1 U4600 ( .B1(B_REG_SCAN_IN), .B2(n4756), .A(n4880), .ZN(n4409) );
  AOI22_X1 U4601 ( .A1(n4094), .A2(n4409), .B1(n4417), .B2(n4093), .ZN(n4095)
         );
  OAI21_X1 U4602 ( .B1(n4128), .B2(n4941), .A(n4095), .ZN(n4096) );
  OAI21_X1 U4603 ( .B1(n4098), .B2(n4950), .A(n4422), .ZN(n4105) );
  INV_X1 U4604 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4103) );
  OAI22_X1 U4605 ( .A1(n4423), .A2(n4338), .B1(n4103), .B2(n2260), .ZN(n4104)
         );
  AOI21_X1 U4606 ( .B1(n4105), .B2(n2260), .A(n4104), .ZN(n4106) );
  OAI21_X1 U4607 ( .B1(n4107), .B2(n4325), .A(n4106), .ZN(U3354) );
  XNOR2_X1 U4608 ( .A(n4108), .B(n4110), .ZN(n4426) );
  XOR2_X1 U4609 ( .A(n4110), .B(n4109), .Z(n4115) );
  OAI22_X1 U4610 ( .A1(n4152), .A2(n4941), .B1(n4939), .B2(n4119), .ZN(n4113)
         );
  INV_X1 U4611 ( .A(n4117), .ZN(n4118) );
  OAI211_X1 U4612 ( .C1(n4133), .C2(n4119), .A(n4118), .B(n5020), .ZN(n4424)
         );
  INV_X1 U4613 ( .A(n4120), .ZN(n4121) );
  AOI22_X1 U4614 ( .A1(n4121), .A2(n4897), .B1(REG2_REG_28__SCAN_IN), .B2(
        n5058), .ZN(n4122) );
  OAI21_X1 U4615 ( .B1(n4424), .B2(n4305), .A(n4122), .ZN(n4123) );
  AOI21_X1 U4616 ( .B1(n4116), .B2(n2260), .A(n4123), .ZN(n4124) );
  OAI21_X1 U4617 ( .B1(n4426), .B2(n4325), .A(n4124), .ZN(U3262) );
  XNOR2_X1 U4618 ( .A(n4125), .B(n4126), .ZN(n4427) );
  INV_X1 U4619 ( .A(n4427), .ZN(n4142) );
  XNOR2_X1 U4620 ( .A(n4127), .B(n4126), .ZN(n4132) );
  NOR2_X1 U4621 ( .A1(n4128), .A2(n4880), .ZN(n4131) );
  OAI22_X1 U4622 ( .A1(n4169), .A2(n4941), .B1(n4129), .B2(n4939), .ZN(n4130)
         );
  AOI211_X1 U4623 ( .C1(n4132), .C2(n4878), .A(n4131), .B(n4130), .ZN(n4428)
         );
  INV_X1 U4624 ( .A(n4428), .ZN(n4140) );
  INV_X1 U4625 ( .A(n4133), .ZN(n4136) );
  NAND2_X1 U4626 ( .A1(n2274), .A2(n4134), .ZN(n4135) );
  NAND2_X1 U4627 ( .A1(n4136), .A2(n4135), .ZN(n4430) );
  AOI22_X1 U4628 ( .A1(n4137), .A2(n4897), .B1(REG2_REG_27__SCAN_IN), .B2(
        n5058), .ZN(n4138) );
  OAI21_X1 U4629 ( .B1(n4430), .B2(n4338), .A(n4138), .ZN(n4139) );
  AOI21_X1 U4630 ( .B1(n4140), .B2(n2260), .A(n4139), .ZN(n4141) );
  OAI21_X1 U4631 ( .B1(n4142), .B2(n4325), .A(n4141), .ZN(U3263) );
  XNOR2_X1 U4632 ( .A(n4144), .B(n4143), .ZN(n4434) );
  INV_X1 U4633 ( .A(n4145), .ZN(n4146) );
  NAND2_X1 U4634 ( .A1(n4147), .A2(n4146), .ZN(n4149) );
  XNOR2_X1 U4635 ( .A(n4149), .B(n4148), .ZN(n4154) );
  AOI22_X1 U4636 ( .A1(n4150), .A2(n4391), .B1(n4156), .B2(n4417), .ZN(n4151)
         );
  OAI21_X1 U4637 ( .B1(n4152), .B2(n4880), .A(n4151), .ZN(n4153) );
  AOI21_X1 U4638 ( .B1(n4154), .B2(n4878), .A(n4153), .ZN(n4433) );
  AOI22_X1 U4639 ( .A1(n4155), .A2(n4897), .B1(REG2_REG_26__SCAN_IN), .B2(
        n5058), .ZN(n4158) );
  NAND2_X1 U4640 ( .A1(n4172), .A2(n4156), .ZN(n4431) );
  NAND3_X1 U4641 ( .A1(n2274), .A2(n5059), .A3(n4431), .ZN(n4157) );
  OAI211_X1 U4642 ( .C1(n4433), .C2(n5058), .A(n4158), .B(n4157), .ZN(n4159)
         );
  INV_X1 U4643 ( .A(n4159), .ZN(n4160) );
  OAI21_X1 U4644 ( .B1(n4434), .B2(n4325), .A(n4160), .ZN(U3264) );
  INV_X1 U4645 ( .A(n4161), .ZN(n4162) );
  XOR2_X1 U4646 ( .A(n4165), .B(n4162), .Z(n4435) );
  INV_X1 U4647 ( .A(n4435), .ZN(n4179) );
  NAND2_X1 U4648 ( .A1(n4164), .A2(n4163), .ZN(n4166) );
  XNOR2_X1 U4649 ( .A(n4166), .B(n4165), .ZN(n4171) );
  AOI22_X1 U4650 ( .A1(n4209), .A2(n4391), .B1(n4417), .B2(n4167), .ZN(n4168)
         );
  OAI21_X1 U4651 ( .B1(n4169), .B2(n4880), .A(n4168), .ZN(n4170) );
  AOI21_X1 U4652 ( .B1(n4171), .B2(n4878), .A(n4170), .ZN(n4436) );
  INV_X1 U4653 ( .A(n4436), .ZN(n4177) );
  OAI21_X1 U4654 ( .B1(n4189), .B2(n4173), .A(n4172), .ZN(n4438) );
  AOI22_X1 U4655 ( .A1(n4174), .A2(n4897), .B1(REG2_REG_25__SCAN_IN), .B2(
        n5058), .ZN(n4175) );
  OAI21_X1 U4656 ( .B1(n4438), .B2(n4338), .A(n4175), .ZN(n4176) );
  AOI21_X1 U4657 ( .B1(n4177), .B2(n2260), .A(n4176), .ZN(n4178) );
  OAI21_X1 U4658 ( .B1(n4179), .B2(n4325), .A(n4178), .ZN(U3265) );
  XNOR2_X1 U4659 ( .A(n4180), .B(n4184), .ZN(n4443) );
  NAND2_X1 U4660 ( .A1(n4182), .A2(n4181), .ZN(n4183) );
  XOR2_X1 U4661 ( .A(n4184), .B(n4183), .Z(n4188) );
  AOI22_X1 U4662 ( .A1(n4224), .A2(n4391), .B1(n4417), .B2(n4191), .ZN(n4185)
         );
  OAI21_X1 U4663 ( .B1(n4186), .B2(n4880), .A(n4185), .ZN(n4187) );
  AOI21_X1 U4664 ( .B1(n4188), .B2(n4878), .A(n4187), .ZN(n4442) );
  INV_X1 U4665 ( .A(n4442), .ZN(n4196) );
  INV_X1 U4666 ( .A(n4189), .ZN(n4440) );
  INV_X1 U4667 ( .A(n4190), .ZN(n4212) );
  NAND2_X1 U4668 ( .A1(n4212), .A2(n4191), .ZN(n4439) );
  AND3_X1 U4669 ( .A1(n4440), .A2(n5059), .A3(n4439), .ZN(n4195) );
  INV_X1 U4670 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4192) );
  OAI22_X1 U4671 ( .A1(n4193), .A2(n4950), .B1(n4192), .B2(n2260), .ZN(n4194)
         );
  AOI211_X1 U4672 ( .C1(n4196), .C2(n2260), .A(n4195), .B(n4194), .ZN(n4197)
         );
  OAI21_X1 U4673 ( .B1(n4443), .B2(n4325), .A(n4197), .ZN(U3266) );
  XOR2_X1 U4674 ( .A(n4206), .B(n4198), .Z(n4445) );
  INV_X1 U4675 ( .A(n4445), .ZN(n4219) );
  INV_X1 U4676 ( .A(n4240), .ZN(n4201) );
  OAI21_X1 U4677 ( .B1(n4201), .B2(n4200), .A(n4199), .ZN(n4220) );
  INV_X1 U4678 ( .A(n4202), .ZN(n4203) );
  AOI21_X1 U4679 ( .B1(n4220), .B2(n4204), .A(n4203), .ZN(n4205) );
  XOR2_X1 U4680 ( .A(n4206), .B(n4205), .Z(n4211) );
  OAI22_X1 U4681 ( .A1(n4207), .A2(n4941), .B1(n4213), .B2(n4939), .ZN(n4208)
         );
  AOI21_X1 U4682 ( .B1(n4944), .B2(n4209), .A(n4208), .ZN(n4210) );
  OAI21_X1 U4683 ( .B1(n4211), .B2(n4946), .A(n4210), .ZN(n4444) );
  OAI21_X1 U4684 ( .B1(n4227), .B2(n4213), .A(n4212), .ZN(n4503) );
  NOR2_X1 U4685 ( .A1(n4503), .A2(n4338), .ZN(n4217) );
  INV_X1 U4686 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4214) );
  OAI22_X1 U4687 ( .A1(n4215), .A2(n4950), .B1(n2260), .B2(n4214), .ZN(n4216)
         );
  AOI211_X1 U4688 ( .C1(n4444), .C2(n2260), .A(n4217), .B(n4216), .ZN(n4218)
         );
  OAI21_X1 U4689 ( .B1(n4219), .B2(n4325), .A(n4218), .ZN(U3267) );
  XNOR2_X1 U4690 ( .A(n4220), .B(n4231), .ZN(n4226) );
  OAI22_X1 U4691 ( .A1(n4222), .A2(n4941), .B1(n4221), .B2(n4939), .ZN(n4223)
         );
  AOI21_X1 U4692 ( .B1(n4944), .B2(n4224), .A(n4223), .ZN(n4225) );
  OAI21_X1 U4693 ( .B1(n4226), .B2(n4946), .A(n4225), .ZN(n4451) );
  INV_X1 U4694 ( .A(n4451), .ZN(n4237) );
  AOI21_X1 U4695 ( .B1(n4058), .B2(n4245), .A(n4227), .ZN(n4452) );
  INV_X1 U4696 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4229) );
  OAI22_X1 U4697 ( .A1(n2260), .A2(n4229), .B1(n4228), .B2(n4950), .ZN(n4235)
         );
  INV_X1 U4698 ( .A(n4230), .ZN(n4449) );
  AOI211_X1 U4699 ( .C1(n4238), .C2(n4233), .A(n4232), .B(n4231), .ZN(n4448)
         );
  NOR3_X1 U4700 ( .A1(n4449), .A2(n4448), .A3(n4325), .ZN(n4234) );
  AOI211_X1 U4701 ( .C1(n4452), .C2(n5059), .A(n4235), .B(n4234), .ZN(n4236)
         );
  OAI21_X1 U4702 ( .B1(n5058), .B2(n4237), .A(n4236), .ZN(U3268) );
  XOR2_X1 U4703 ( .A(n4239), .B(n4238), .Z(n4455) );
  INV_X1 U4704 ( .A(n4455), .ZN(n4252) );
  XNOR2_X1 U4705 ( .A(n4240), .B(n4239), .ZN(n4244) );
  OAI22_X1 U4706 ( .A1(n5031), .A2(n4941), .B1(n4246), .B2(n4939), .ZN(n4241)
         );
  AOI21_X1 U4707 ( .B1(n4944), .B2(n4242), .A(n4241), .ZN(n4243) );
  OAI21_X1 U4708 ( .B1(n4244), .B2(n4946), .A(n4243), .ZN(n4454) );
  OAI21_X1 U4709 ( .B1(n2328), .B2(n4246), .A(n4245), .ZN(n4731) );
  NOR2_X1 U4710 ( .A1(n4731), .A2(n4338), .ZN(n4250) );
  INV_X1 U4711 ( .A(REG2_REG_21__SCAN_IN), .ZN(n4248) );
  OAI22_X1 U4712 ( .A1(n2260), .A2(n4248), .B1(n4247), .B2(n4950), .ZN(n4249)
         );
  AOI211_X1 U4713 ( .C1(n4454), .C2(n2260), .A(n4250), .B(n4249), .ZN(n4251)
         );
  OAI21_X1 U4714 ( .B1(n4252), .B2(n4325), .A(n4251), .ZN(U3269) );
  XOR2_X1 U4715 ( .A(n4256), .B(n4253), .Z(n4458) );
  NAND2_X1 U4716 ( .A1(n4255), .A2(n4254), .ZN(n4257) );
  XNOR2_X1 U4717 ( .A(n4257), .B(n4256), .ZN(n4261) );
  AOI22_X1 U4718 ( .A1(n5039), .A2(n4944), .B1(n4417), .B2(n5049), .ZN(n4258)
         );
  OAI21_X1 U4719 ( .B1(n4259), .B2(n4941), .A(n4258), .ZN(n4260) );
  AOI21_X1 U4720 ( .B1(n4261), .B2(n4878), .A(n4260), .ZN(n4262) );
  OAI21_X1 U4721 ( .B1(n4458), .B2(n4397), .A(n4262), .ZN(n4459) );
  NAND2_X1 U4722 ( .A1(n4459), .A2(n2260), .ZN(n4269) );
  NAND2_X1 U4723 ( .A1(n2302), .A2(n5049), .ZN(n4263) );
  NAND2_X1 U4724 ( .A1(n4264), .A2(n4263), .ZN(n4735) );
  INV_X1 U4725 ( .A(n4735), .ZN(n4267) );
  INV_X1 U4726 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4265) );
  OAI22_X1 U4727 ( .A1(n2260), .A2(n4265), .B1(n5053), .B2(n4950), .ZN(n4266)
         );
  AOI21_X1 U4728 ( .B1(n4267), .B2(n5059), .A(n4266), .ZN(n4268) );
  OAI211_X1 U4729 ( .C1(n4458), .C2(n4406), .A(n4269), .B(n4268), .ZN(U3270)
         );
  INV_X1 U4730 ( .A(n4270), .ZN(n4271) );
  OR2_X1 U4731 ( .A1(n4310), .A2(n4271), .ZN(n4273) );
  NAND2_X1 U4732 ( .A1(n4273), .A2(n4272), .ZN(n4292) );
  INV_X1 U4733 ( .A(n4274), .ZN(n4275) );
  AOI21_X1 U4734 ( .B1(n4292), .B2(n4276), .A(n4275), .ZN(n4277) );
  XOR2_X1 U4735 ( .A(n4283), .B(n4277), .Z(n4281) );
  OAI22_X1 U4736 ( .A1(n4312), .A2(n4941), .B1(n4284), .B2(n4939), .ZN(n4278)
         );
  AOI21_X1 U4737 ( .B1(n4944), .B2(n4279), .A(n4278), .ZN(n4280) );
  OAI21_X1 U4738 ( .B1(n4281), .B2(n4946), .A(n4280), .ZN(n4463) );
  INV_X1 U4739 ( .A(n4463), .ZN(n4290) );
  XOR2_X1 U4740 ( .A(n4283), .B(n4282), .Z(n4464) );
  OR2_X1 U4741 ( .A1(n4301), .A2(n4284), .ZN(n4285) );
  NAND2_X1 U4742 ( .A1(n2302), .A2(n4285), .ZN(n4739) );
  AOI22_X1 U4743 ( .A1(n5058), .A2(REG2_REG_19__SCAN_IN), .B1(n4286), .B2(
        n4897), .ZN(n4287) );
  OAI21_X1 U4744 ( .B1(n4739), .B2(n4338), .A(n4287), .ZN(n4288) );
  AOI21_X1 U4745 ( .B1(n4464), .B2(n4365), .A(n4288), .ZN(n4289) );
  OAI21_X1 U4746 ( .B1(n4290), .B2(n5058), .A(n4289), .ZN(U3271) );
  XNOR2_X1 U4747 ( .A(n4292), .B(n4291), .ZN(n4297) );
  NAND2_X1 U4748 ( .A1(n4293), .A2(n4391), .ZN(n4295) );
  NAND2_X1 U4749 ( .A1(n5046), .A2(n4944), .ZN(n4294) );
  OAI211_X1 U4750 ( .C1(n4300), .C2(n4939), .A(n4295), .B(n4294), .ZN(n4296)
         );
  AOI21_X1 U4751 ( .B1(n4297), .B2(n4878), .A(n4296), .ZN(n4470) );
  XNOR2_X1 U4752 ( .A(n4299), .B(n4298), .ZN(n4468) );
  OAI21_X1 U4753 ( .B1(n4319), .B2(n4300), .A(n5020), .ZN(n4302) );
  OR2_X1 U4754 ( .A1(n4302), .A2(n4301), .ZN(n4466) );
  AOI22_X1 U4755 ( .A1(n5058), .A2(REG2_REG_18__SCAN_IN), .B1(n4303), .B2(
        n4897), .ZN(n4304) );
  OAI21_X1 U4756 ( .B1(n4466), .B2(n4305), .A(n4304), .ZN(n4306) );
  AOI21_X1 U4757 ( .B1(n4468), .B2(n4365), .A(n4306), .ZN(n4307) );
  OAI21_X1 U4758 ( .B1(n4470), .B2(n5058), .A(n4307), .ZN(U3272) );
  XOR2_X1 U4759 ( .A(n4309), .B(n4308), .Z(n5016) );
  XNOR2_X1 U4760 ( .A(n4310), .B(n4309), .ZN(n4316) );
  OAI22_X1 U4761 ( .A1(n4312), .A2(n4880), .B1(n4311), .B2(n4939), .ZN(n4313)
         );
  AOI21_X1 U4762 ( .B1(n4391), .B2(n4314), .A(n4313), .ZN(n4315) );
  OAI21_X1 U4763 ( .B1(n4316), .B2(n4946), .A(n4315), .ZN(n5018) );
  NAND2_X1 U4764 ( .A1(n5018), .A2(n2260), .ZN(n4324) );
  AND2_X1 U4765 ( .A1(n4335), .A2(n4317), .ZN(n4318) );
  NOR2_X1 U4766 ( .A1(n4319), .A2(n4318), .ZN(n5019) );
  OAI22_X1 U4767 ( .A1(n2260), .A2(n4321), .B1(n4320), .B2(n4950), .ZN(n4322)
         );
  AOI21_X1 U4768 ( .B1(n5019), .B2(n5059), .A(n4322), .ZN(n4323) );
  OAI211_X1 U4769 ( .C1(n4325), .C2(n5016), .A(n4324), .B(n4323), .ZN(U3273)
         );
  OAI211_X1 U4770 ( .C1(n4327), .C2(n4333), .A(n4326), .B(n4878), .ZN(n4331)
         );
  AOI22_X1 U4771 ( .A1(n4329), .A2(n4391), .B1(n4417), .B2(n4328), .ZN(n4330)
         );
  OAI211_X1 U4772 ( .C1(n4332), .C2(n4880), .A(n4331), .B(n4330), .ZN(n4473)
         );
  INV_X1 U4773 ( .A(n4473), .ZN(n4344) );
  XOR2_X1 U4774 ( .A(n4334), .B(n4333), .Z(n4474) );
  INV_X1 U4775 ( .A(n4353), .ZN(n4337) );
  OAI21_X1 U4776 ( .B1(n4337), .B2(n4336), .A(n4335), .ZN(n4746) );
  NOR2_X1 U4777 ( .A1(n4746), .A2(n4338), .ZN(n4342) );
  OAI22_X1 U4778 ( .A1(n2260), .A2(n4340), .B1(n4339), .B2(n4950), .ZN(n4341)
         );
  AOI211_X1 U4779 ( .C1(n4474), .C2(n4365), .A(n4342), .B(n4341), .ZN(n4343)
         );
  OAI21_X1 U4780 ( .B1(n5058), .B2(n4344), .A(n4343), .ZN(U3274) );
  OAI22_X1 U4781 ( .A1(n4993), .A2(n4880), .B1(n4351), .B2(n4939), .ZN(n4349)
         );
  INV_X1 U4782 ( .A(n4345), .ZN(n4346) );
  AOI211_X1 U4783 ( .C1(n4347), .C2(n4364), .A(n4946), .B(n4346), .ZN(n4348)
         );
  AOI211_X1 U4784 ( .C1(n4391), .C2(n4350), .A(n4349), .B(n4348), .ZN(n5005)
         );
  OR2_X1 U4785 ( .A1(n4377), .A2(n4351), .ZN(n4352) );
  NAND2_X1 U4786 ( .A1(n4353), .A2(n4352), .ZN(n5006) );
  INV_X1 U4787 ( .A(n5006), .ZN(n4356) );
  OAI22_X1 U4788 ( .A1(n2260), .A2(n4354), .B1(n5004), .B2(n4950), .ZN(n4355)
         );
  AOI21_X1 U4789 ( .B1(n4356), .B2(n5059), .A(n4355), .ZN(n4367) );
  NAND2_X1 U4790 ( .A1(n4357), .A2(n4358), .ZN(n4361) );
  INV_X1 U4791 ( .A(n4359), .ZN(n4360) );
  NAND2_X1 U4792 ( .A1(n4361), .A2(n4360), .ZN(n4368) );
  AOI21_X1 U4793 ( .B1(n4368), .B2(n4369), .A(n4362), .ZN(n4363) );
  XOR2_X1 U4794 ( .A(n4364), .B(n4363), .Z(n5009) );
  NAND2_X1 U4795 ( .A1(n5009), .A2(n4365), .ZN(n4366) );
  OAI211_X1 U4796 ( .C1(n5005), .C2(n5058), .A(n4367), .B(n4366), .ZN(U3275)
         );
  XNOR2_X1 U4797 ( .A(n4368), .B(n4369), .ZN(n4477) );
  XNOR2_X1 U4798 ( .A(n4075), .B(n4369), .ZN(n4375) );
  OAI22_X1 U4799 ( .A1(n4371), .A2(n4880), .B1(n4370), .B2(n4939), .ZN(n4372)
         );
  AOI21_X1 U4800 ( .B1(n4391), .B2(n4373), .A(n4372), .ZN(n4374) );
  OAI21_X1 U4801 ( .B1(n4375), .B2(n4946), .A(n4374), .ZN(n4376) );
  AOI21_X1 U4802 ( .B1(n4477), .B2(n4934), .A(n4376), .ZN(n4481) );
  INV_X1 U4803 ( .A(n4377), .ZN(n4479) );
  INV_X1 U4804 ( .A(n4398), .ZN(n4379) );
  NAND2_X1 U4805 ( .A1(n4379), .A2(n4378), .ZN(n4478) );
  AND3_X1 U4806 ( .A1(n4479), .A2(n5059), .A3(n4478), .ZN(n4384) );
  INV_X1 U4807 ( .A(n4380), .ZN(n4381) );
  OAI22_X1 U4808 ( .A1(n2260), .A2(n4382), .B1(n4381), .B2(n4950), .ZN(n4383)
         );
  AOI211_X1 U4809 ( .C1(n4477), .C2(n4900), .A(n4384), .B(n4383), .ZN(n4385)
         );
  OAI21_X1 U4810 ( .B1(n4481), .B2(n5058), .A(n4385), .ZN(U3276) );
  XNOR2_X1 U4811 ( .A(n4357), .B(n4390), .ZN(n4984) );
  OAI21_X1 U4812 ( .B1(n4388), .B2(n4387), .A(n4386), .ZN(n4389) );
  XOR2_X1 U4813 ( .A(n4390), .B(n4389), .Z(n4395) );
  AOI22_X1 U4814 ( .A1(n4392), .A2(n4391), .B1(n4399), .B2(n4417), .ZN(n4393)
         );
  OAI21_X1 U4815 ( .B1(n4992), .B2(n4880), .A(n4393), .ZN(n4394) );
  AOI21_X1 U4816 ( .B1(n4395), .B2(n4878), .A(n4394), .ZN(n4396) );
  OAI21_X1 U4817 ( .B1(n4397), .B2(n4984), .A(n4396), .ZN(n4985) );
  NAND2_X1 U4818 ( .A1(n4985), .A2(n2260), .ZN(n4405) );
  AOI21_X1 U4819 ( .B1(n4399), .B2(n2273), .A(n4398), .ZN(n4987) );
  INV_X1 U4820 ( .A(n4400), .ZN(n4401) );
  OAI22_X1 U4821 ( .A1(n2260), .A2(n4402), .B1(n4401), .B2(n4950), .ZN(n4403)
         );
  AOI21_X1 U4822 ( .B1(n4987), .B2(n5059), .A(n4403), .ZN(n4404) );
  OAI211_X1 U4823 ( .C1(n4984), .C2(n4406), .A(n4405), .B(n4404), .ZN(U3277)
         );
  XOR2_X1 U4824 ( .A(n4408), .B(n4414), .Z(n5060) );
  INV_X1 U4825 ( .A(n5060), .ZN(n4490) );
  INV_X1 U4826 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4412) );
  INV_X1 U4827 ( .A(n4408), .ZN(n4411) );
  AND2_X1 U4828 ( .A1(n4410), .A2(n4409), .ZN(n4416) );
  AOI21_X1 U4829 ( .B1(n4411), .B2(n4417), .A(n4416), .ZN(n5062) );
  MUX2_X1 U4830 ( .A(n4412), .B(n5062), .S(n5022), .Z(n4413) );
  OAI21_X1 U4831 ( .B1(n4490), .B2(n4487), .A(n4413), .ZN(U3549) );
  AOI21_X1 U4832 ( .B1(n4418), .B2(n4415), .A(n4414), .ZN(n5055) );
  INV_X1 U4833 ( .A(n5055), .ZN(n4493) );
  INV_X1 U4834 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4419) );
  AOI21_X1 U4835 ( .B1(n4418), .B2(n4417), .A(n4416), .ZN(n5057) );
  MUX2_X1 U4836 ( .A(n4419), .B(n5057), .S(n5022), .Z(n4420) );
  OAI21_X1 U4837 ( .B1(n4493), .B2(n4487), .A(n4420), .ZN(U3548) );
  OAI211_X1 U4838 ( .C1(n4426), .C2(n5015), .A(n4425), .B(n4424), .ZN(n4495)
         );
  MUX2_X1 U4839 ( .A(REG1_REG_28__SCAN_IN), .B(n4495), .S(n5022), .Z(U3546) );
  NAND2_X1 U4840 ( .A1(n4427), .A2(n5010), .ZN(n4429) );
  OAI211_X1 U4841 ( .C1(n5007), .C2(n4430), .A(n4429), .B(n4428), .ZN(n4496)
         );
  MUX2_X1 U4842 ( .A(REG1_REG_27__SCAN_IN), .B(n4496), .S(n5022), .Z(U3545) );
  NAND3_X1 U4843 ( .A1(n2274), .A2(n5020), .A3(n4431), .ZN(n4432) );
  OAI211_X1 U4844 ( .C1(n4434), .C2(n5015), .A(n4433), .B(n4432), .ZN(n4497)
         );
  MUX2_X1 U4845 ( .A(REG1_REG_26__SCAN_IN), .B(n4497), .S(n5022), .Z(U3544) );
  NAND2_X1 U4846 ( .A1(n4435), .A2(n5010), .ZN(n4437) );
  OAI211_X1 U4847 ( .C1(n5007), .C2(n4438), .A(n4437), .B(n4436), .ZN(n4498)
         );
  MUX2_X1 U4848 ( .A(REG1_REG_25__SCAN_IN), .B(n4498), .S(n5022), .Z(U3543) );
  NAND3_X1 U4849 ( .A1(n4440), .A2(n5020), .A3(n4439), .ZN(n4441) );
  OAI211_X1 U4850 ( .C1(n4443), .C2(n5015), .A(n4442), .B(n4441), .ZN(n4499)
         );
  MUX2_X1 U4851 ( .A(REG1_REG_24__SCAN_IN), .B(n4499), .S(n5022), .Z(U3542) );
  INV_X1 U4852 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4446) );
  AOI21_X1 U4853 ( .B1(n4445), .B2(n5010), .A(n4444), .ZN(n4500) );
  MUX2_X1 U4854 ( .A(n4446), .B(n4500), .S(n5022), .Z(n4447) );
  OAI21_X1 U4855 ( .B1(n4503), .B2(n4487), .A(n4447), .ZN(U3541) );
  NOR3_X1 U4856 ( .A1(n4449), .A2(n4448), .A3(n5015), .ZN(n4450) );
  AOI211_X1 U4857 ( .C1(n5020), .C2(n4452), .A(n4451), .B(n4450), .ZN(n4504)
         );
  NAND2_X1 U4858 ( .A1(n5021), .A2(REG1_REG_22__SCAN_IN), .ZN(n4453) );
  OAI21_X1 U4859 ( .B1(n4504), .B2(n5021), .A(n4453), .ZN(U3540) );
  INV_X1 U4860 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4456) );
  AOI21_X1 U4861 ( .B1(n4455), .B2(n5010), .A(n4454), .ZN(n4728) );
  MUX2_X1 U4862 ( .A(n4456), .B(n4728), .S(n5022), .Z(n4457) );
  OAI21_X1 U4863 ( .B1(n4487), .B2(n4731), .A(n4457), .ZN(U3539) );
  INV_X1 U4864 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4461) );
  INV_X1 U4865 ( .A(n4458), .ZN(n4460) );
  AOI21_X1 U4866 ( .B1(n4975), .B2(n4460), .A(n4459), .ZN(n4732) );
  MUX2_X1 U4867 ( .A(n4461), .B(n4732), .S(n5022), .Z(n4462) );
  OAI21_X1 U4868 ( .B1(n4487), .B2(n4735), .A(n4462), .ZN(U3538) );
  AOI21_X1 U4869 ( .B1(n4464), .B2(n5010), .A(n4463), .ZN(n4736) );
  MUX2_X1 U4870 ( .A(n4029), .B(n4736), .S(n5022), .Z(n4465) );
  OAI21_X1 U4871 ( .B1(n4487), .B2(n4739), .A(n4465), .ZN(U3537) );
  INV_X1 U4872 ( .A(n4466), .ZN(n4467) );
  AOI21_X1 U4873 ( .B1(n4468), .B2(n5010), .A(n4467), .ZN(n4469) );
  AND2_X1 U4874 ( .A1(n4470), .A2(n4469), .ZN(n4740) );
  MUX2_X1 U4875 ( .A(n4471), .B(n4740), .S(n5022), .Z(n4472) );
  INV_X1 U4876 ( .A(n4472), .ZN(U3536) );
  INV_X1 U4877 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4475) );
  AOI21_X1 U4878 ( .B1(n5010), .B2(n4474), .A(n4473), .ZN(n4743) );
  MUX2_X1 U4879 ( .A(n4475), .B(n4743), .S(n5022), .Z(n4476) );
  OAI21_X1 U4880 ( .B1(n4746), .B2(n4487), .A(n4476), .ZN(U3534) );
  INV_X1 U4881 ( .A(n4477), .ZN(n4482) );
  NAND3_X1 U4882 ( .A1(n4479), .A2(n5020), .A3(n4478), .ZN(n4480) );
  OAI211_X1 U4883 ( .C1(n4482), .C2(n4983), .A(n4481), .B(n4480), .ZN(n4747)
         );
  MUX2_X1 U4884 ( .A(REG1_REG_14__SCAN_IN), .B(n4747), .S(n5022), .Z(U3532) );
  NAND2_X1 U4885 ( .A1(n4483), .A2(n5010), .ZN(n4484) );
  AND2_X1 U4886 ( .A1(n4485), .A2(n4484), .ZN(n4749) );
  MUX2_X1 U4887 ( .A(n4843), .B(n4749), .S(n5022), .Z(n4486) );
  OAI21_X1 U4888 ( .B1(n4752), .B2(n4487), .A(n4486), .ZN(U3530) );
  INV_X1 U4889 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4488) );
  MUX2_X1 U4890 ( .A(n4488), .B(n5062), .S(n5025), .Z(n4489) );
  OAI21_X1 U4891 ( .B1(n4490), .B2(n4751), .A(n4489), .ZN(U3517) );
  INV_X1 U4892 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4491) );
  MUX2_X1 U4893 ( .A(n4491), .B(n5057), .S(n5025), .Z(n4492) );
  OAI21_X1 U4894 ( .B1(n4493), .B2(n4751), .A(n4492), .ZN(U3516) );
  MUX2_X1 U4895 ( .A(REG0_REG_29__SCAN_IN), .B(n4494), .S(n5025), .Z(U3515) );
  MUX2_X1 U4896 ( .A(REG0_REG_28__SCAN_IN), .B(n4495), .S(n5025), .Z(U3514) );
  MUX2_X1 U4897 ( .A(REG0_REG_27__SCAN_IN), .B(n4496), .S(n5025), .Z(U3513) );
  MUX2_X1 U4898 ( .A(REG0_REG_26__SCAN_IN), .B(n4497), .S(n5025), .Z(U3512) );
  MUX2_X1 U4899 ( .A(REG0_REG_25__SCAN_IN), .B(n4498), .S(n5025), .Z(U3511) );
  MUX2_X1 U4900 ( .A(REG0_REG_24__SCAN_IN), .B(n4499), .S(n5025), .Z(U3510) );
  INV_X1 U4901 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4501) );
  MUX2_X1 U4902 ( .A(n4501), .B(n4500), .S(n5025), .Z(n4502) );
  OAI21_X1 U4903 ( .B1(n4503), .B2(n4751), .A(n4502), .ZN(U3509) );
  MUX2_X1 U4904 ( .A(n4505), .B(n4504), .S(n5025), .Z(n4727) );
  OAI22_X1 U4905 ( .A1(n4507), .A2(keyinput_45), .B1(REG3_REG_16__SCAN_IN), 
        .B2(keyinput_46), .ZN(n4506) );
  AOI221_X1 U4906 ( .B1(n4507), .B2(keyinput_45), .C1(keyinput_46), .C2(
        REG3_REG_16__SCAN_IN), .A(n4506), .ZN(n4510) );
  OAI22_X1 U4907 ( .A1(n4684), .A2(keyinput_44), .B1(keyinput_43), .B2(
        REG3_REG_21__SCAN_IN), .ZN(n4508) );
  AOI221_X1 U4908 ( .B1(n4684), .B2(keyinput_44), .C1(REG3_REG_21__SCAN_IN), 
        .C2(keyinput_43), .A(n4508), .ZN(n4509) );
  OAI211_X1 U4909 ( .C1(REG3_REG_5__SCAN_IN), .C2(keyinput_47), .A(n4510), .B(
        n4509), .ZN(n4511) );
  AOI21_X1 U4910 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_47), .A(n4511), .ZN(
        n4582) );
  AOI22_X1 U4911 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_39), .B1(n4671), 
        .B2(keyinput_34), .ZN(n4512) );
  OAI221_X1 U4912 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_39), .C1(n4671), 
        .C2(keyinput_34), .A(n4512), .ZN(n4576) );
  OAI22_X1 U4913 ( .A1(n4514), .A2(keyinput_36), .B1(n3586), .B2(keyinput_40), 
        .ZN(n4513) );
  AOI221_X1 U4914 ( .B1(n4514), .B2(keyinput_36), .C1(keyinput_40), .C2(n3586), 
        .A(n4513), .ZN(n4571) );
  OAI22_X1 U4915 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_37), .B1(
        keyinput_35), .B2(REG3_REG_14__SCAN_IN), .ZN(n4515) );
  AOI221_X1 U4916 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_37), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_35), .A(n4515), .ZN(n4570) );
  INV_X1 U4917 ( .A(keyinput_23), .ZN(n4553) );
  INV_X1 U4918 ( .A(DATAI_8_), .ZN(n4652) );
  INV_X1 U4919 ( .A(keyinput_22), .ZN(n4551) );
  INV_X1 U4920 ( .A(DATAI_9_), .ZN(n4958) );
  INV_X1 U4921 ( .A(DATAI_12_), .ZN(n4979) );
  OAI22_X1 U4922 ( .A1(n4979), .A2(keyinput_19), .B1(keyinput_21), .B2(
        DATAI_10_), .ZN(n4516) );
  AOI221_X1 U4923 ( .B1(n4979), .B2(keyinput_19), .C1(DATAI_10_), .C2(
        keyinput_21), .A(n4516), .ZN(n4548) );
  INV_X1 U4924 ( .A(DATAI_13_), .ZN(n4981) );
  INV_X1 U4925 ( .A(keyinput_18), .ZN(n4546) );
  INV_X1 U4926 ( .A(DATAI_14_), .ZN(n4642) );
  INV_X1 U4927 ( .A(DATAI_19_), .ZN(n4610) );
  OAI22_X1 U4928 ( .A1(n4610), .A2(keyinput_12), .B1(keyinput_13), .B2(
        DATAI_18_), .ZN(n4517) );
  AOI221_X1 U4929 ( .B1(n4610), .B2(keyinput_12), .C1(DATAI_18_), .C2(
        keyinput_13), .A(n4517), .ZN(n4539) );
  INV_X1 U4930 ( .A(keyinput_11), .ZN(n4537) );
  OAI22_X1 U4931 ( .A1(n4519), .A2(keyinput_9), .B1(DATAI_23_), .B2(keyinput_8), .ZN(n4518) );
  AOI221_X1 U4932 ( .B1(n4519), .B2(keyinput_9), .C1(keyinput_8), .C2(
        DATAI_23_), .A(n4518), .ZN(n4533) );
  INV_X1 U4933 ( .A(keyinput_7), .ZN(n4531) );
  INV_X1 U4934 ( .A(DATAI_25_), .ZN(n4529) );
  INV_X1 U4935 ( .A(keyinput_3), .ZN(n4524) );
  INV_X1 U4936 ( .A(DATAI_28_), .ZN(n4618) );
  INV_X1 U4937 ( .A(keyinput_2), .ZN(n4522) );
  OAI22_X1 U4938 ( .A1(DATAI_31_), .A2(keyinput_0), .B1(DATAI_30_), .B2(
        keyinput_1), .ZN(n4520) );
  AOI221_X1 U4939 ( .B1(DATAI_31_), .B2(keyinput_0), .C1(keyinput_1), .C2(
        DATAI_30_), .A(n4520), .ZN(n4521) );
  AOI221_X1 U4940 ( .B1(DATAI_29_), .B2(n4522), .C1(n4614), .C2(keyinput_2), 
        .A(n4521), .ZN(n4523) );
  AOI221_X1 U4941 ( .B1(DATAI_28_), .B2(n4524), .C1(n4618), .C2(keyinput_3), 
        .A(n4523), .ZN(n4527) );
  AOI22_X1 U4942 ( .A1(DATAI_27_), .A2(keyinput_4), .B1(n4620), .B2(keyinput_5), .ZN(n4525) );
  OAI221_X1 U4943 ( .B1(DATAI_27_), .B2(keyinput_4), .C1(n4620), .C2(
        keyinput_5), .A(n4525), .ZN(n4526) );
  AOI211_X1 U4944 ( .C1(n4529), .C2(keyinput_6), .A(n4527), .B(n4526), .ZN(
        n4528) );
  OAI21_X1 U4945 ( .B1(n4529), .B2(keyinput_6), .A(n4528), .ZN(n4530) );
  OAI221_X1 U4946 ( .B1(DATAI_24_), .B2(keyinput_7), .C1(n4626), .C2(n4531), 
        .A(n4530), .ZN(n4532) );
  AOI22_X1 U4947 ( .A1(keyinput_10), .A2(n4535), .B1(n4533), .B2(n4532), .ZN(
        n4534) );
  OAI21_X1 U4948 ( .B1(n4535), .B2(keyinput_10), .A(n4534), .ZN(n4536) );
  OAI221_X1 U4949 ( .B1(DATAI_20_), .B2(keyinput_11), .C1(n4631), .C2(n4537), 
        .A(n4536), .ZN(n4538) );
  OAI211_X1 U4950 ( .C1(n4636), .C2(keyinput_14), .A(n4539), .B(n4538), .ZN(
        n4540) );
  AOI21_X1 U4951 ( .B1(n4636), .B2(keyinput_14), .A(n4540), .ZN(n4543) );
  INV_X1 U4952 ( .A(DATAI_15_), .ZN(n4638) );
  INV_X1 U4953 ( .A(DATAI_16_), .ZN(n5014) );
  AOI22_X1 U4954 ( .A1(n4638), .A2(keyinput_16), .B1(n5014), .B2(keyinput_15), 
        .ZN(n4541) );
  OAI221_X1 U4955 ( .B1(n4638), .B2(keyinput_16), .C1(n5014), .C2(keyinput_15), 
        .A(n4541), .ZN(n4542) );
  AOI211_X1 U4956 ( .C1(n4642), .C2(keyinput_17), .A(n4543), .B(n4542), .ZN(
        n4544) );
  OAI21_X1 U4957 ( .B1(n4642), .B2(keyinput_17), .A(n4544), .ZN(n4545) );
  OAI221_X1 U4958 ( .B1(DATAI_13_), .B2(keyinput_18), .C1(n4981), .C2(n4546), 
        .A(n4545), .ZN(n4547) );
  OAI211_X1 U4959 ( .C1(DATAI_11_), .C2(keyinput_20), .A(n4548), .B(n4547), 
        .ZN(n4549) );
  AOI21_X1 U4960 ( .B1(DATAI_11_), .B2(keyinput_20), .A(n4549), .ZN(n4550) );
  AOI221_X1 U4961 ( .B1(DATAI_9_), .B2(n4551), .C1(n4958), .C2(keyinput_22), 
        .A(n4550), .ZN(n4552) );
  AOI221_X1 U4962 ( .B1(DATAI_8_), .B2(n4553), .C1(n4652), .C2(keyinput_23), 
        .A(n4552), .ZN(n4561) );
  INV_X1 U4963 ( .A(DATAI_6_), .ZN(n4926) );
  INV_X1 U4964 ( .A(DATAI_7_), .ZN(n4654) );
  AOI22_X1 U4965 ( .A1(n4926), .A2(keyinput_25), .B1(n4654), .B2(keyinput_24), 
        .ZN(n4554) );
  OAI221_X1 U4966 ( .B1(n4926), .B2(keyinput_25), .C1(n4654), .C2(keyinput_24), 
        .A(n4554), .ZN(n4560) );
  OAI22_X1 U4967 ( .A1(DATAI_5_), .A2(keyinput_26), .B1(keyinput_28), .B2(
        DATAI_3_), .ZN(n4555) );
  AOI221_X1 U4968 ( .B1(DATAI_5_), .B2(keyinput_26), .C1(DATAI_3_), .C2(
        keyinput_28), .A(n4555), .ZN(n4559) );
  XOR2_X1 U4969 ( .A(DATAI_2_), .B(keyinput_29), .Z(n4557) );
  XNOR2_X1 U4970 ( .A(DATAI_4_), .B(keyinput_27), .ZN(n4556) );
  NOR2_X1 U4971 ( .A1(n4557), .A2(n4556), .ZN(n4558) );
  OAI211_X1 U4972 ( .C1(n4561), .C2(n4560), .A(n4559), .B(n4558), .ZN(n4566)
         );
  OAI22_X1 U4973 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_33), .B1(keyinput_30), .B2(DATAI_1_), .ZN(n4562) );
  AOI221_X1 U4974 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_33), .C1(DATAI_1_), 
        .C2(keyinput_30), .A(n4562), .ZN(n4565) );
  XNOR2_X1 U4975 ( .A(STATE_REG_SCAN_IN), .B(keyinput_32), .ZN(n4564) );
  XNOR2_X1 U4976 ( .A(DATAI_0_), .B(keyinput_31), .ZN(n4563) );
  NAND4_X1 U4977 ( .A1(n4566), .A2(n4565), .A3(n4564), .A4(n4563), .ZN(n4569)
         );
  XOR2_X1 U4978 ( .A(n4567), .B(keyinput_38), .Z(n4568) );
  NAND4_X1 U4979 ( .A1(n4571), .A2(n4570), .A3(n4569), .A4(n4568), .ZN(n4575)
         );
  OAI22_X1 U4980 ( .A1(n4573), .A2(keyinput_41), .B1(keyinput_42), .B2(
        REG3_REG_1__SCAN_IN), .ZN(n4572) );
  AOI221_X1 U4981 ( .B1(n4573), .B2(keyinput_41), .C1(REG3_REG_1__SCAN_IN), 
        .C2(keyinput_42), .A(n4572), .ZN(n4574) );
  OAI21_X1 U4982 ( .B1(n4576), .B2(n4575), .A(n4574), .ZN(n4581) );
  AOI22_X1 U4983 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_51), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput_50), .ZN(n4577) );
  OAI221_X1 U4984 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_51), .C1(
        REG3_REG_4__SCAN_IN), .C2(keyinput_50), .A(n4577), .ZN(n4580) );
  AOI22_X1 U4985 ( .A1(REG3_REG_24__SCAN_IN), .A2(keyinput_49), .B1(
        REG3_REG_17__SCAN_IN), .B2(keyinput_48), .ZN(n4578) );
  OAI221_X1 U4986 ( .B1(REG3_REG_24__SCAN_IN), .B2(keyinput_49), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_48), .A(n4578), .ZN(n4579) );
  AOI211_X1 U4987 ( .C1(n4582), .C2(n4581), .A(n4580), .B(n4579), .ZN(n4586)
         );
  AOI22_X1 U4988 ( .A1(n4698), .A2(keyinput_53), .B1(n4699), .B2(keyinput_54), 
        .ZN(n4583) );
  OAI221_X1 U4989 ( .B1(n4698), .B2(keyinput_53), .C1(n4699), .C2(keyinput_54), 
        .A(n4583), .ZN(n4585) );
  XOR2_X1 U4990 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .Z(n4584) );
  NOR3_X1 U4991 ( .A1(n4586), .A2(n4585), .A3(n4584), .ZN(n4592) );
  INV_X1 U4992 ( .A(keyinput_55), .ZN(n4587) );
  MUX2_X1 U4993 ( .A(keyinput_55), .B(n4587), .S(IR_REG_0__SCAN_IN), .Z(n4588)
         );
  INV_X1 U4994 ( .A(n4588), .ZN(n4591) );
  INV_X1 U4995 ( .A(keyinput_56), .ZN(n4589) );
  MUX2_X1 U4996 ( .A(keyinput_56), .B(n4589), .S(IR_REG_1__SCAN_IN), .Z(n4590)
         );
  OAI21_X1 U4997 ( .B1(n4592), .B2(n4591), .A(n4590), .ZN(n4598) );
  INV_X1 U4998 ( .A(keyinput_57), .ZN(n4593) );
  MUX2_X1 U4999 ( .A(n4593), .B(keyinput_57), .S(IR_REG_2__SCAN_IN), .Z(n4597)
         );
  XNOR2_X1 U5000 ( .A(n4594), .B(keyinput_59), .ZN(n4596) );
  XNOR2_X1 U5001 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_58), .ZN(n4595) );
  AOI211_X1 U5002 ( .C1(n4598), .C2(n4597), .A(n4596), .B(n4595), .ZN(n4603)
         );
  XNOR2_X1 U5003 ( .A(n4599), .B(keyinput_60), .ZN(n4602) );
  INV_X1 U5004 ( .A(keyinput_61), .ZN(n4600) );
  MUX2_X1 U5005 ( .A(keyinput_61), .B(n4600), .S(IR_REG_6__SCAN_IN), .Z(n4601)
         );
  OAI21_X1 U5006 ( .B1(n4603), .B2(n4602), .A(n4601), .ZN(n4606) );
  INV_X1 U5007 ( .A(keyinput_62), .ZN(n4604) );
  MUX2_X1 U5008 ( .A(n4604), .B(keyinput_62), .S(IR_REG_7__SCAN_IN), .Z(n4605)
         );
  NAND2_X1 U5009 ( .A1(n4606), .A2(n4605), .ZN(n4725) );
  INV_X1 U5010 ( .A(keyinput_63), .ZN(n4607) );
  MUX2_X1 U5011 ( .A(keyinput_63), .B(n4607), .S(keyinput_127), .Z(n4724) );
  INV_X1 U5012 ( .A(keyinput_87), .ZN(n4651) );
  INV_X1 U5013 ( .A(keyinput_86), .ZN(n4649) );
  INV_X1 U5014 ( .A(DATAI_10_), .ZN(n4968) );
  OAI22_X1 U5015 ( .A1(n4979), .A2(keyinput_83), .B1(DATAI_11_), .B2(
        keyinput_84), .ZN(n4608) );
  AOI221_X1 U5016 ( .B1(n4979), .B2(keyinput_83), .C1(keyinput_84), .C2(
        DATAI_11_), .A(n4608), .ZN(n4646) );
  INV_X1 U5017 ( .A(keyinput_82), .ZN(n4644) );
  OAI22_X1 U5018 ( .A1(n4610), .A2(keyinput_76), .B1(DATAI_18_), .B2(
        keyinput_77), .ZN(n4609) );
  AOI221_X1 U5019 ( .B1(n4610), .B2(keyinput_76), .C1(keyinput_77), .C2(
        DATAI_18_), .A(n4609), .ZN(n4634) );
  INV_X1 U5020 ( .A(keyinput_75), .ZN(n4632) );
  OAI22_X1 U5021 ( .A1(DATAI_23_), .A2(keyinput_72), .B1(keyinput_73), .B2(
        DATAI_22_), .ZN(n4611) );
  AOI221_X1 U5022 ( .B1(DATAI_23_), .B2(keyinput_72), .C1(DATAI_22_), .C2(
        keyinput_73), .A(n4611), .ZN(n4628) );
  INV_X1 U5023 ( .A(keyinput_71), .ZN(n4625) );
  INV_X1 U5024 ( .A(keyinput_67), .ZN(n4617) );
  INV_X1 U5025 ( .A(keyinput_66), .ZN(n4615) );
  OAI22_X1 U5026 ( .A1(DATAI_31_), .A2(keyinput_64), .B1(DATAI_30_), .B2(
        keyinput_65), .ZN(n4612) );
  AOI221_X1 U5027 ( .B1(DATAI_31_), .B2(keyinput_64), .C1(keyinput_65), .C2(
        DATAI_30_), .A(n4612), .ZN(n4613) );
  AOI221_X1 U5028 ( .B1(DATAI_29_), .B2(n4615), .C1(n4614), .C2(keyinput_66), 
        .A(n4613), .ZN(n4616) );
  AOI221_X1 U5029 ( .B1(DATAI_28_), .B2(keyinput_67), .C1(n4618), .C2(n4617), 
        .A(n4616), .ZN(n4622) );
  AOI22_X1 U5030 ( .A1(DATAI_27_), .A2(keyinput_68), .B1(n4620), .B2(
        keyinput_69), .ZN(n4619) );
  OAI221_X1 U5031 ( .B1(DATAI_27_), .B2(keyinput_68), .C1(n4620), .C2(
        keyinput_69), .A(n4619), .ZN(n4621) );
  AOI211_X1 U5032 ( .C1(DATAI_25_), .C2(keyinput_70), .A(n4622), .B(n4621), 
        .ZN(n4623) );
  OAI21_X1 U5033 ( .B1(DATAI_25_), .B2(keyinput_70), .A(n4623), .ZN(n4624) );
  OAI221_X1 U5034 ( .B1(DATAI_24_), .B2(keyinput_71), .C1(n4626), .C2(n4625), 
        .A(n4624), .ZN(n4627) );
  AOI22_X1 U5035 ( .A1(n4628), .A2(n4627), .B1(keyinput_74), .B2(DATAI_21_), 
        .ZN(n4629) );
  OAI21_X1 U5036 ( .B1(keyinput_74), .B2(DATAI_21_), .A(n4629), .ZN(n4630) );
  OAI221_X1 U5037 ( .B1(DATAI_20_), .B2(n4632), .C1(n4631), .C2(keyinput_75), 
        .A(n4630), .ZN(n4633) );
  OAI211_X1 U5038 ( .C1(n4636), .C2(keyinput_78), .A(n4634), .B(n4633), .ZN(
        n4635) );
  AOI21_X1 U5039 ( .B1(n4636), .B2(keyinput_78), .A(n4635), .ZN(n4640) );
  AOI22_X1 U5040 ( .A1(DATAI_16_), .A2(keyinput_79), .B1(n4638), .B2(
        keyinput_80), .ZN(n4637) );
  OAI221_X1 U5041 ( .B1(DATAI_16_), .B2(keyinput_79), .C1(n4638), .C2(
        keyinput_80), .A(n4637), .ZN(n4639) );
  AOI211_X1 U5042 ( .C1(n4642), .C2(keyinput_81), .A(n4640), .B(n4639), .ZN(
        n4641) );
  OAI21_X1 U5043 ( .B1(n4642), .B2(keyinput_81), .A(n4641), .ZN(n4643) );
  OAI221_X1 U5044 ( .B1(DATAI_13_), .B2(keyinput_82), .C1(n4981), .C2(n4644), 
        .A(n4643), .ZN(n4645) );
  OAI211_X1 U5045 ( .C1(n4968), .C2(keyinput_85), .A(n4646), .B(n4645), .ZN(
        n4647) );
  AOI21_X1 U5046 ( .B1(n4968), .B2(keyinput_85), .A(n4647), .ZN(n4648) );
  AOI221_X1 U5047 ( .B1(DATAI_9_), .B2(n4649), .C1(n4958), .C2(keyinput_86), 
        .A(n4648), .ZN(n4650) );
  AOI221_X1 U5048 ( .B1(DATAI_8_), .B2(keyinput_87), .C1(n4652), .C2(n4651), 
        .A(n4650), .ZN(n4663) );
  AOI22_X1 U5049 ( .A1(n4926), .A2(keyinput_89), .B1(n4654), .B2(keyinput_88), 
        .ZN(n4653) );
  OAI221_X1 U5050 ( .B1(n4926), .B2(keyinput_89), .C1(n4654), .C2(keyinput_88), 
        .A(n4653), .ZN(n4662) );
  INV_X1 U5051 ( .A(DATAI_4_), .ZN(n4656) );
  OAI22_X1 U5052 ( .A1(n4656), .A2(keyinput_91), .B1(DATAI_3_), .B2(
        keyinput_92), .ZN(n4655) );
  AOI221_X1 U5053 ( .B1(n4656), .B2(keyinput_91), .C1(keyinput_92), .C2(
        DATAI_3_), .A(n4655), .ZN(n4661) );
  XOR2_X1 U5054 ( .A(DATAI_2_), .B(keyinput_93), .Z(n4659) );
  INV_X1 U5055 ( .A(DATAI_5_), .ZN(n4657) );
  XNOR2_X1 U5056 ( .A(keyinput_90), .B(n4657), .ZN(n4658) );
  NOR2_X1 U5057 ( .A1(n4659), .A2(n4658), .ZN(n4660) );
  OAI211_X1 U5058 ( .C1(n4663), .C2(n4662), .A(n4661), .B(n4660), .ZN(n4679)
         );
  AOI22_X1 U5059 ( .A1(U3149), .A2(keyinput_96), .B1(keyinput_97), .B2(n4665), 
        .ZN(n4664) );
  OAI221_X1 U5060 ( .B1(U3149), .B2(keyinput_96), .C1(n4665), .C2(keyinput_97), 
        .A(n4664), .ZN(n4668) );
  XOR2_X1 U5061 ( .A(DATAI_1_), .B(keyinput_94), .Z(n4667) );
  XNOR2_X1 U5062 ( .A(DATAI_0_), .B(keyinput_95), .ZN(n4666) );
  NOR3_X1 U5063 ( .A1(n4668), .A2(n4667), .A3(n4666), .ZN(n4678) );
  OAI22_X1 U5064 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_100), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_104), .ZN(n4669) );
  AOI221_X1 U5065 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_100), .C1(
        keyinput_104), .C2(REG3_REG_28__SCAN_IN), .A(n4669), .ZN(n4674) );
  AOI22_X1 U5066 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_102), .B1(n4671), 
        .B2(keyinput_98), .ZN(n4670) );
  OAI221_X1 U5067 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_102), .C1(n4671), 
        .C2(keyinput_98), .A(n4670), .ZN(n4672) );
  AOI21_X1 U5068 ( .B1(keyinput_103), .B2(n3452), .A(n4672), .ZN(n4673) );
  OAI211_X1 U5069 ( .C1(keyinput_103), .C2(n3452), .A(n4674), .B(n4673), .ZN(
        n4677) );
  AOI22_X1 U5070 ( .A1(REG3_REG_14__SCAN_IN), .A2(keyinput_99), .B1(
        REG3_REG_10__SCAN_IN), .B2(keyinput_101), .ZN(n4675) );
  OAI221_X1 U5071 ( .B1(REG3_REG_14__SCAN_IN), .B2(keyinput_99), .C1(
        REG3_REG_10__SCAN_IN), .C2(keyinput_101), .A(n4675), .ZN(n4676) );
  AOI211_X1 U5072 ( .C1(n4679), .C2(n4678), .A(n4677), .B(n4676), .ZN(n4682)
         );
  XOR2_X1 U5073 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_106), .Z(n4681) );
  XNOR2_X1 U5074 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_105), .ZN(n4680) );
  NOR3_X1 U5075 ( .A1(n4682), .A2(n4681), .A3(n4680), .ZN(n4696) );
  OAI22_X1 U5076 ( .A1(n4684), .A2(keyinput_108), .B1(keyinput_109), .B2(
        REG3_REG_25__SCAN_IN), .ZN(n4683) );
  AOI221_X1 U5077 ( .B1(n4684), .B2(keyinput_108), .C1(REG3_REG_25__SCAN_IN), 
        .C2(keyinput_109), .A(n4683), .ZN(n4689) );
  OAI22_X1 U5078 ( .A1(n4686), .A2(keyinput_107), .B1(REG3_REG_16__SCAN_IN), 
        .B2(keyinput_110), .ZN(n4685) );
  AOI221_X1 U5079 ( .B1(n4686), .B2(keyinput_107), .C1(keyinput_110), .C2(
        REG3_REG_16__SCAN_IN), .A(n4685), .ZN(n4688) );
  XOR2_X1 U5080 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_111), .Z(n4687) );
  NAND3_X1 U5081 ( .A1(n4689), .A2(n4688), .A3(n4687), .ZN(n4695) );
  OAI22_X1 U5082 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_114), .B1(
        keyinput_113), .B2(REG3_REG_24__SCAN_IN), .ZN(n4690) );
  AOI221_X1 U5083 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_114), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_113), .A(n4690), .ZN(n4694) );
  OAI22_X1 U5084 ( .A1(n4692), .A2(keyinput_112), .B1(keyinput_115), .B2(
        REG3_REG_9__SCAN_IN), .ZN(n4691) );
  AOI221_X1 U5085 ( .B1(n4692), .B2(keyinput_112), .C1(REG3_REG_9__SCAN_IN), 
        .C2(keyinput_115), .A(n4691), .ZN(n4693) );
  OAI211_X1 U5086 ( .C1(n4696), .C2(n4695), .A(n4694), .B(n4693), .ZN(n4702)
         );
  OAI22_X1 U5087 ( .A1(n4699), .A2(keyinput_118), .B1(n4698), .B2(keyinput_117), .ZN(n4697) );
  AOI221_X1 U5088 ( .B1(n4699), .B2(keyinput_118), .C1(keyinput_117), .C2(
        n4698), .A(n4697), .ZN(n4701) );
  XNOR2_X1 U5089 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_116), .ZN(n4700) );
  NAND3_X1 U5090 ( .A1(n4702), .A2(n4701), .A3(n4700), .ZN(n4708) );
  INV_X1 U5091 ( .A(keyinput_119), .ZN(n4703) );
  MUX2_X1 U5092 ( .A(keyinput_119), .B(n4703), .S(IR_REG_0__SCAN_IN), .Z(n4704) );
  INV_X1 U5093 ( .A(n4704), .ZN(n4707) );
  INV_X1 U5094 ( .A(keyinput_120), .ZN(n4705) );
  MUX2_X1 U5095 ( .A(keyinput_120), .B(n4705), .S(IR_REG_1__SCAN_IN), .Z(n4706) );
  AOI21_X1 U5096 ( .B1(n4708), .B2(n4707), .A(n4706), .ZN(n4713) );
  INV_X1 U5097 ( .A(keyinput_121), .ZN(n4709) );
  MUX2_X1 U5098 ( .A(n4709), .B(keyinput_121), .S(IR_REG_2__SCAN_IN), .Z(n4712) );
  XNOR2_X1 U5099 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_123), .ZN(n4711) );
  XNOR2_X1 U5100 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n4710) );
  OAI211_X1 U5101 ( .C1(n4713), .C2(n4712), .A(n4711), .B(n4710), .ZN(n4715)
         );
  XNOR2_X1 U5102 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_124), .ZN(n4714) );
  NAND2_X1 U5103 ( .A1(n4715), .A2(n4714), .ZN(n4720) );
  INV_X1 U5104 ( .A(IR_REG_6__SCAN_IN), .ZN(n4716) );
  XNOR2_X1 U5105 ( .A(n4716), .B(keyinput_125), .ZN(n4719) );
  XNOR2_X1 U5106 ( .A(n4717), .B(keyinput_126), .ZN(n4718) );
  AOI21_X1 U5107 ( .B1(n4720), .B2(n4719), .A(n4718), .ZN(n4723) );
  XNOR2_X1 U5108 ( .A(n4721), .B(keyinput_127), .ZN(n4722) );
  AOI211_X1 U5109 ( .C1(n4725), .C2(n4724), .A(n4723), .B(n4722), .ZN(n4726)
         );
  XNOR2_X1 U5110 ( .A(n4727), .B(n4726), .ZN(U3508) );
  INV_X1 U5111 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4729) );
  MUX2_X1 U5112 ( .A(n4729), .B(n4728), .S(n5025), .Z(n4730) );
  OAI21_X1 U5113 ( .B1(n4731), .B2(n4751), .A(n4730), .ZN(U3507) );
  INV_X1 U5114 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4733) );
  MUX2_X1 U5115 ( .A(n4733), .B(n4732), .S(n5025), .Z(n4734) );
  OAI21_X1 U5116 ( .B1(n4735), .B2(n4751), .A(n4734), .ZN(U3506) );
  INV_X1 U5117 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4737) );
  MUX2_X1 U5118 ( .A(n4737), .B(n4736), .S(n5025), .Z(n4738) );
  OAI21_X1 U5119 ( .B1(n4739), .B2(n4751), .A(n4738), .ZN(U3505) );
  MUX2_X1 U5120 ( .A(n4741), .B(n4740), .S(n5025), .Z(n4742) );
  INV_X1 U5121 ( .A(n4742), .ZN(U3503) );
  INV_X1 U5122 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4744) );
  MUX2_X1 U5123 ( .A(n4744), .B(n4743), .S(n5025), .Z(n4745) );
  OAI21_X1 U5124 ( .B1(n4746), .B2(n4751), .A(n4745), .ZN(U3499) );
  MUX2_X1 U5125 ( .A(REG0_REG_14__SCAN_IN), .B(n4747), .S(n5025), .Z(U3495) );
  INV_X1 U5126 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4748) );
  MUX2_X1 U5127 ( .A(n4749), .B(n4748), .S(n5023), .Z(n4750) );
  OAI21_X1 U5128 ( .B1(n4752), .B2(n4751), .A(n4750), .ZN(U3491) );
  MUX2_X1 U5129 ( .A(n4753), .B(D_REG_1__SCAN_IN), .S(n4769), .Z(U3459) );
  MUX2_X1 U5130 ( .A(DATAI_30_), .B(n4754), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5131 ( .A(n4755), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U5132 ( .A(DATAI_27_), .B(n4756), .S(STATE_REG_SCAN_IN), .Z(U3325)
         );
  MUX2_X1 U5133 ( .A(n4936), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U5134 ( .A(DATAI_18_), .B(n4757), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5135 ( .A(n4758), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5136 ( .A(n4759), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5137 ( .A(n4760), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U5138 ( .A(n4761), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5139 ( .A(DATAI_5_), .B(n4762), .S(STATE_REG_SCAN_IN), .Z(U3347) );
  MUX2_X1 U5140 ( .A(n4763), .B(DATAI_4_), .S(U3149), .Z(U3348) );
  MUX2_X1 U5141 ( .A(n4764), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5142 ( .A(n4765), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5143 ( .A(n4766), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5144 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5145 ( .A(DATAI_23_), .ZN(n4768) );
  OAI21_X1 U5146 ( .B1(STATE_REG_SCAN_IN), .B2(n4768), .A(n4767), .ZN(U3329)
         );
  INV_X1 U5147 ( .A(D_REG_2__SCAN_IN), .ZN(n4770) );
  NOR2_X1 U5148 ( .A1(n4800), .A2(n4770), .ZN(U3320) );
  INV_X1 U5149 ( .A(D_REG_3__SCAN_IN), .ZN(n4771) );
  NOR2_X1 U5150 ( .A1(n4800), .A2(n4771), .ZN(U3319) );
  INV_X1 U5151 ( .A(D_REG_4__SCAN_IN), .ZN(n4772) );
  NOR2_X1 U5152 ( .A1(n4800), .A2(n4772), .ZN(U3318) );
  INV_X1 U5153 ( .A(D_REG_5__SCAN_IN), .ZN(n4773) );
  NOR2_X1 U5154 ( .A1(n4800), .A2(n4773), .ZN(U3317) );
  INV_X1 U5155 ( .A(D_REG_6__SCAN_IN), .ZN(n4774) );
  NOR2_X1 U5156 ( .A1(n4800), .A2(n4774), .ZN(U3316) );
  INV_X1 U5157 ( .A(D_REG_7__SCAN_IN), .ZN(n4775) );
  NOR2_X1 U5158 ( .A1(n4800), .A2(n4775), .ZN(U3315) );
  INV_X1 U5159 ( .A(D_REG_8__SCAN_IN), .ZN(n4776) );
  NOR2_X1 U5160 ( .A1(n4800), .A2(n4776), .ZN(U3314) );
  INV_X1 U5161 ( .A(D_REG_9__SCAN_IN), .ZN(n4777) );
  NOR2_X1 U5162 ( .A1(n4800), .A2(n4777), .ZN(U3313) );
  INV_X1 U5163 ( .A(D_REG_10__SCAN_IN), .ZN(n4778) );
  NOR2_X1 U5164 ( .A1(n4800), .A2(n4778), .ZN(U3312) );
  INV_X1 U5165 ( .A(D_REG_11__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5166 ( .A1(n4800), .A2(n4779), .ZN(U3311) );
  INV_X1 U5167 ( .A(D_REG_12__SCAN_IN), .ZN(n4780) );
  NOR2_X1 U5168 ( .A1(n4800), .A2(n4780), .ZN(U3310) );
  INV_X1 U5169 ( .A(D_REG_13__SCAN_IN), .ZN(n4781) );
  NOR2_X1 U5170 ( .A1(n4800), .A2(n4781), .ZN(U3309) );
  INV_X1 U5171 ( .A(D_REG_14__SCAN_IN), .ZN(n4782) );
  NOR2_X1 U5172 ( .A1(n4800), .A2(n4782), .ZN(U3308) );
  INV_X1 U5173 ( .A(D_REG_15__SCAN_IN), .ZN(n4783) );
  NOR2_X1 U5174 ( .A1(n4800), .A2(n4783), .ZN(U3307) );
  INV_X1 U5175 ( .A(D_REG_16__SCAN_IN), .ZN(n4784) );
  NOR2_X1 U5176 ( .A1(n4800), .A2(n4784), .ZN(U3306) );
  INV_X1 U5177 ( .A(D_REG_17__SCAN_IN), .ZN(n4785) );
  NOR2_X1 U5178 ( .A1(n4800), .A2(n4785), .ZN(U3305) );
  INV_X1 U5179 ( .A(D_REG_18__SCAN_IN), .ZN(n4786) );
  NOR2_X1 U5180 ( .A1(n4800), .A2(n4786), .ZN(U3304) );
  INV_X1 U5181 ( .A(D_REG_19__SCAN_IN), .ZN(n4787) );
  NOR2_X1 U5182 ( .A1(n4800), .A2(n4787), .ZN(U3303) );
  INV_X1 U5183 ( .A(D_REG_20__SCAN_IN), .ZN(n4788) );
  NOR2_X1 U5184 ( .A1(n4800), .A2(n4788), .ZN(U3302) );
  INV_X1 U5185 ( .A(D_REG_21__SCAN_IN), .ZN(n4789) );
  NOR2_X1 U5186 ( .A1(n4800), .A2(n4789), .ZN(U3301) );
  INV_X1 U5187 ( .A(D_REG_22__SCAN_IN), .ZN(n4790) );
  NOR2_X1 U5188 ( .A1(n4800), .A2(n4790), .ZN(U3300) );
  INV_X1 U5189 ( .A(D_REG_23__SCAN_IN), .ZN(n4791) );
  NOR2_X1 U5190 ( .A1(n4800), .A2(n4791), .ZN(U3299) );
  INV_X1 U5191 ( .A(D_REG_24__SCAN_IN), .ZN(n4792) );
  NOR2_X1 U5192 ( .A1(n4800), .A2(n4792), .ZN(U3298) );
  INV_X1 U5193 ( .A(D_REG_25__SCAN_IN), .ZN(n4793) );
  NOR2_X1 U5194 ( .A1(n4800), .A2(n4793), .ZN(U3297) );
  INV_X1 U5195 ( .A(D_REG_26__SCAN_IN), .ZN(n4794) );
  NOR2_X1 U5196 ( .A1(n4800), .A2(n4794), .ZN(U3296) );
  INV_X1 U5197 ( .A(D_REG_27__SCAN_IN), .ZN(n4795) );
  NOR2_X1 U5198 ( .A1(n4800), .A2(n4795), .ZN(U3295) );
  NOR2_X1 U5199 ( .A1(n4800), .A2(n4796), .ZN(U3294) );
  NOR2_X1 U5200 ( .A1(n4800), .A2(n4797), .ZN(U3293) );
  NOR2_X1 U5201 ( .A1(n4800), .A2(n4798), .ZN(U3292) );
  NOR2_X1 U5202 ( .A1(n4800), .A2(n4799), .ZN(U3291) );
  AOI211_X1 U5203 ( .C1(n4803), .C2(n4802), .A(n4801), .B(n4864), .ZN(n4805)
         );
  AOI211_X1 U5204 ( .C1(n4869), .C2(ADDR_REG_6__SCAN_IN), .A(n4805), .B(n4804), 
        .ZN(n4809) );
  OAI211_X1 U5205 ( .C1(REG1_REG_6__SCAN_IN), .C2(n4807), .A(n4870), .B(n4806), 
        .ZN(n4808) );
  OAI211_X1 U5206 ( .C1(n4875), .C2(n4927), .A(n4809), .B(n4808), .ZN(U3246)
         );
  AOI22_X1 U5207 ( .A1(n4810), .A2(n4964), .B1(REG1_REG_9__SCAN_IN), .B2(n4959), .ZN(n4812) );
  OAI21_X1 U5208 ( .B1(n4813), .B2(n4812), .A(n4870), .ZN(n4811) );
  AOI21_X1 U5209 ( .B1(n4813), .B2(n4812), .A(n4811), .ZN(n4815) );
  AOI211_X1 U5210 ( .C1(n4869), .C2(ADDR_REG_9__SCAN_IN), .A(n4815), .B(n4814), 
        .ZN(n4820) );
  OAI211_X1 U5211 ( .C1(n4818), .C2(n4817), .A(n4847), .B(n4816), .ZN(n4819)
         );
  OAI211_X1 U5212 ( .C1(n4875), .C2(n4959), .A(n4820), .B(n4819), .ZN(U3249)
         );
  AOI21_X1 U5213 ( .B1(n4869), .B2(ADDR_REG_10__SCAN_IN), .A(n4821), .ZN(n4829) );
  NAND2_X1 U5214 ( .A1(n4967), .A2(n4823), .ZN(n4827) );
  OAI211_X1 U5215 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4825), .A(n4847), .B(n4824), .ZN(n4826) );
  NAND4_X1 U5216 ( .A1(n4829), .A2(n4828), .A3(n4827), .A4(n4826), .ZN(U3250)
         );
  AOI21_X1 U5217 ( .B1(n4970), .B2(n4976), .A(n4830), .ZN(n4833) );
  OAI21_X1 U5218 ( .B1(n4833), .B2(n4832), .A(n4870), .ZN(n4831) );
  AOI21_X1 U5219 ( .B1(n4833), .B2(n4832), .A(n4831), .ZN(n4835) );
  AOI211_X1 U5220 ( .C1(n4869), .C2(ADDR_REG_11__SCAN_IN), .A(n4835), .B(n4834), .ZN(n4840) );
  OAI211_X1 U5221 ( .C1(n4838), .C2(n4837), .A(n4847), .B(n4836), .ZN(n4839)
         );
  OAI211_X1 U5222 ( .C1(n4875), .C2(n4970), .A(n4840), .B(n4839), .ZN(U3251)
         );
  AOI211_X1 U5223 ( .C1(n4843), .C2(n4842), .A(n4841), .B(n4863), .ZN(n4845)
         );
  AOI211_X1 U5224 ( .C1(n4869), .C2(ADDR_REG_12__SCAN_IN), .A(n4845), .B(n4844), .ZN(n4850) );
  OAI211_X1 U5225 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4848), .A(n4847), .B(n4846), .ZN(n4849) );
  OAI211_X1 U5226 ( .C1(n4875), .C2(n4980), .A(n4850), .B(n4849), .ZN(U3252)
         );
  OAI21_X1 U5227 ( .B1(n4852), .B2(REG1_REG_13__SCAN_IN), .A(n4851), .ZN(n4854) );
  XNOR2_X1 U5228 ( .A(n4854), .B(n4853), .ZN(n4862) );
  AOI21_X1 U5229 ( .B1(n4982), .B2(n4402), .A(n4855), .ZN(n4857) );
  XNOR2_X1 U5230 ( .A(n4857), .B(n4856), .ZN(n4858) );
  OAI22_X1 U5231 ( .A1(n4982), .A2(n4875), .B1(n4864), .B2(n4858), .ZN(n4859)
         );
  AOI211_X1 U5232 ( .C1(n4869), .C2(ADDR_REG_13__SCAN_IN), .A(n4860), .B(n4859), .ZN(n4861) );
  OAI21_X1 U5233 ( .B1(n4863), .B2(n4862), .A(n4861), .ZN(U3253) );
  AOI221_X1 U5234 ( .B1(n4866), .B2(n4865), .C1(n4340), .C2(n4865), .A(n4864), 
        .ZN(n4867) );
  AOI211_X1 U5235 ( .C1(n4869), .C2(ADDR_REG_16__SCAN_IN), .A(n4868), .B(n4867), .ZN(n4874) );
  OAI221_X1 U5236 ( .B1(n4872), .B2(REG1_REG_16__SCAN_IN), .C1(n4872), .C2(
        n4871), .A(n4870), .ZN(n4873) );
  OAI211_X1 U5237 ( .C1(n4875), .C2(n2485), .A(n4874), .B(n4873), .ZN(U3256)
         );
  INV_X1 U5238 ( .A(n4876), .ZN(n4877) );
  NOR2_X1 U5239 ( .A1(n2314), .A2(n4877), .ZN(n4886) );
  OAI21_X1 U5240 ( .B1(n4934), .B2(n4878), .A(n4887), .ZN(n4879) );
  OAI21_X1 U5241 ( .B1(n2990), .B2(n4880), .A(n4879), .ZN(n4884) );
  AOI211_X1 U5242 ( .C1(n4975), .C2(n4887), .A(n4886), .B(n4884), .ZN(n4883)
         );
  AOI22_X1 U5243 ( .A1(n5022), .A2(n4883), .B1(n4881), .B2(n5021), .ZN(U3518)
         );
  INV_X1 U5244 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4882) );
  AOI22_X1 U5245 ( .A1(n5025), .A2(n4883), .B1(n4882), .B2(n5023), .ZN(U3467)
         );
  AOI21_X1 U5246 ( .B1(n4886), .B2(n4885), .A(n4884), .ZN(n4890) );
  AOI22_X1 U5247 ( .A1(n4887), .A2(n4900), .B1(REG3_REG_0__SCAN_IN), .B2(n4897), .ZN(n4888) );
  OAI221_X1 U5248 ( .B1(n5058), .B2(n4890), .C1(n2260), .C2(n4889), .A(n4888), 
        .ZN(U3290) );
  OAI22_X1 U5249 ( .A1(n4892), .A2(n5015), .B1(n5007), .B2(n4891), .ZN(n4893)
         );
  NOR2_X1 U5250 ( .A1(n4894), .A2(n4893), .ZN(n4896) );
  AOI22_X1 U5251 ( .A1(n5022), .A2(n4896), .B1(n2610), .B2(n5021), .ZN(U3519)
         );
  INV_X1 U5252 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4895) );
  AOI22_X1 U5253 ( .A1(n5025), .A2(n4896), .B1(n4895), .B2(n5023), .ZN(U3469)
         );
  AOI22_X1 U5254 ( .A1(REG2_REG_2__SCAN_IN), .A2(n5058), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4897), .ZN(n4903) );
  INV_X1 U5255 ( .A(n4898), .ZN(n4901) );
  AOI22_X1 U5256 ( .A1(n4901), .A2(n4900), .B1(n5059), .B2(n4899), .ZN(n4902)
         );
  OAI211_X1 U5257 ( .C1(n5058), .C2(n4904), .A(n4903), .B(n4902), .ZN(U3288)
         );
  OAI22_X1 U5258 ( .A1(n4906), .A2(n4983), .B1(n5007), .B2(n4905), .ZN(n4907)
         );
  NOR2_X1 U5259 ( .A1(n4908), .A2(n4907), .ZN(n4911) );
  INV_X1 U5260 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4909) );
  AOI22_X1 U5261 ( .A1(n5022), .A2(n4911), .B1(n4909), .B2(n5021), .ZN(U3521)
         );
  INV_X1 U5262 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4910) );
  AOI22_X1 U5263 ( .A1(n5025), .A2(n4911), .B1(n4910), .B2(n5023), .ZN(U3473)
         );
  INV_X1 U5264 ( .A(n4912), .ZN(n4916) );
  INV_X1 U5265 ( .A(n4913), .ZN(n4914) );
  AOI211_X1 U5266 ( .C1(n4916), .C2(n4975), .A(n4915), .B(n4914), .ZN(n4919)
         );
  AOI22_X1 U5267 ( .A1(n5022), .A2(n4919), .B1(n4917), .B2(n5021), .ZN(U3522)
         );
  INV_X1 U5268 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4918) );
  AOI22_X1 U5269 ( .A1(n5025), .A2(n4919), .B1(n4918), .B2(n5023), .ZN(U3475)
         );
  NOR2_X1 U5270 ( .A1(n4920), .A2(n5015), .ZN(n4921) );
  AOI211_X1 U5271 ( .C1(n5020), .C2(n4923), .A(n4922), .B(n4921), .ZN(n4925)
         );
  AOI22_X1 U5272 ( .A1(n5022), .A2(n4925), .B1(n2661), .B2(n5021), .ZN(U3523)
         );
  INV_X1 U5273 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4924) );
  AOI22_X1 U5274 ( .A1(n5025), .A2(n4925), .B1(n4924), .B2(n5023), .ZN(U3477)
         );
  AOI22_X1 U5275 ( .A1(STATE_REG_SCAN_IN), .A2(n4927), .B1(n4926), .B2(U3149), 
        .ZN(U3346) );
  OAI211_X1 U5276 ( .C1(n4929), .C2(n4940), .A(n5020), .B(n4928), .ZN(n4952)
         );
  INV_X1 U5277 ( .A(n4930), .ZN(n4931) );
  AOI21_X1 U5278 ( .B1(n4937), .B2(n4932), .A(n4931), .ZN(n4955) );
  OAI21_X1 U5279 ( .B1(n4934), .B2(n4933), .A(n4955), .ZN(n4935) );
  OAI211_X1 U5280 ( .C1(n4936), .C2(n4952), .A(n4935), .B(n2260), .ZN(n4948)
         );
  XOR2_X1 U5281 ( .A(n4938), .B(n4937), .Z(n4947) );
  OAI22_X1 U5282 ( .A1(n2466), .A2(n4941), .B1(n4940), .B2(n4939), .ZN(n4942)
         );
  AOI21_X1 U5283 ( .B1(n4944), .B2(n4943), .A(n4942), .ZN(n4945) );
  OAI21_X1 U5284 ( .B1(n4947), .B2(n4946), .A(n4945), .ZN(n4953) );
  OAI22_X1 U5285 ( .A1(n4948), .A2(n4953), .B1(REG2_REG_7__SCAN_IN), .B2(n2260), .ZN(n4949) );
  OAI21_X1 U5286 ( .B1(n4951), .B2(n4950), .A(n4949), .ZN(U3283) );
  INV_X1 U5287 ( .A(n4952), .ZN(n4954) );
  AOI211_X1 U5288 ( .C1(n4955), .C2(n5010), .A(n4954), .B(n4953), .ZN(n4957)
         );
  AOI22_X1 U5289 ( .A1(n5022), .A2(n4957), .B1(n2495), .B2(n5021), .ZN(U3525)
         );
  INV_X1 U5290 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4956) );
  AOI22_X1 U5291 ( .A1(n5025), .A2(n4957), .B1(n4956), .B2(n5023), .ZN(U3481)
         );
  AOI22_X1 U5292 ( .A1(STATE_REG_SCAN_IN), .A2(n4959), .B1(n4958), .B2(U3149), 
        .ZN(U3343) );
  NOR2_X1 U5293 ( .A1(n4960), .A2(n4983), .ZN(n4962) );
  AOI211_X1 U5294 ( .C1(n5020), .C2(n4963), .A(n4962), .B(n4961), .ZN(n4966)
         );
  AOI22_X1 U5295 ( .A1(n5022), .A2(n4966), .B1(n4964), .B2(n5021), .ZN(U3527)
         );
  INV_X1 U5296 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4965) );
  AOI22_X1 U5297 ( .A1(n5025), .A2(n4966), .B1(n4965), .B2(n5023), .ZN(U3485)
         );
  AOI22_X1 U5298 ( .A1(STATE_REG_SCAN_IN), .A2(n3951), .B1(n4968), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5299 ( .A(DATAI_11_), .ZN(n4969) );
  AOI22_X1 U5300 ( .A1(STATE_REG_SCAN_IN), .A2(n4970), .B1(n4969), .B2(U3149), 
        .ZN(U3341) );
  NOR2_X1 U5301 ( .A1(n4971), .A2(n5007), .ZN(n4973) );
  AOI211_X1 U5302 ( .C1(n4975), .C2(n4974), .A(n4973), .B(n4972), .ZN(n4978)
         );
  AOI22_X1 U5303 ( .A1(n5022), .A2(n4978), .B1(n4976), .B2(n5021), .ZN(U3529)
         );
  INV_X1 U5304 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4977) );
  AOI22_X1 U5305 ( .A1(n5025), .A2(n4978), .B1(n4977), .B2(n5023), .ZN(U3489)
         );
  AOI22_X1 U5306 ( .A1(STATE_REG_SCAN_IN), .A2(n4980), .B1(n4979), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5307 ( .A1(STATE_REG_SCAN_IN), .A2(n4982), .B1(n4981), .B2(U3149), 
        .ZN(U3339) );
  NOR2_X1 U5308 ( .A1(n4984), .A2(n4983), .ZN(n4986) );
  AOI211_X1 U5309 ( .C1(n5020), .C2(n4987), .A(n4986), .B(n4985), .ZN(n4990)
         );
  AOI22_X1 U5310 ( .A1(n5022), .A2(n4990), .B1(n4988), .B2(n5021), .ZN(U3531)
         );
  INV_X1 U5311 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4989) );
  AOI22_X1 U5312 ( .A1(n5025), .A2(n4990), .B1(n4989), .B2(n5023), .ZN(U3493)
         );
  OAI22_X1 U5313 ( .A1(n5032), .A2(n4993), .B1(n4992), .B2(n4991), .ZN(n4994)
         );
  AOI211_X1 U5314 ( .C1(n4996), .C2(n5050), .A(n4995), .B(n4994), .ZN(n5003)
         );
  NAND2_X1 U5315 ( .A1(n4998), .A2(n4997), .ZN(n4999) );
  XOR2_X1 U5316 ( .A(n5000), .B(n4999), .Z(n5001) );
  NAND2_X1 U5317 ( .A1(n5001), .A2(n5048), .ZN(n5002) );
  OAI211_X1 U5318 ( .C1(n5054), .C2(n5004), .A(n5003), .B(n5002), .ZN(U3238)
         );
  OAI21_X1 U5319 ( .B1(n5007), .B2(n5006), .A(n5005), .ZN(n5008) );
  AOI21_X1 U5320 ( .B1(n5010), .B2(n5009), .A(n5008), .ZN(n5013) );
  AOI22_X1 U5321 ( .A1(n5022), .A2(n5013), .B1(n5011), .B2(n5021), .ZN(U3533)
         );
  INV_X1 U5322 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5012) );
  AOI22_X1 U5323 ( .A1(n5025), .A2(n5013), .B1(n5012), .B2(n5023), .ZN(U3497)
         );
  AOI22_X1 U5324 ( .A1(STATE_REG_SCAN_IN), .A2(n2485), .B1(n5014), .B2(U3149), 
        .ZN(U3336) );
  NOR2_X1 U5325 ( .A1(n5016), .A2(n5015), .ZN(n5017) );
  AOI211_X1 U5326 ( .C1(n5020), .C2(n5019), .A(n5018), .B(n5017), .ZN(n5024)
         );
  AOI22_X1 U5327 ( .A1(n5022), .A2(n5024), .B1(n3993), .B2(n5021), .ZN(U3535)
         );
  AOI22_X1 U5328 ( .A1(n5025), .A2(n5024), .B1(n3422), .B2(n5023), .ZN(U3501)
         );
  AOI22_X1 U5329 ( .A1(n5045), .A2(n5027), .B1(n5026), .B2(n5050), .ZN(n5037)
         );
  OAI21_X1 U5330 ( .B1(n5030), .B2(n5029), .A(n5028), .ZN(n5035) );
  NOR2_X1 U5331 ( .A1(n5032), .A2(n5031), .ZN(n5034) );
  AOI211_X1 U5332 ( .C1(n5035), .C2(n5048), .A(n5034), .B(n5033), .ZN(n5036)
         );
  OAI211_X1 U5333 ( .C1(n5054), .C2(n5038), .A(n5037), .B(n5036), .ZN(U3216)
         );
  AOI22_X1 U5334 ( .A1(n5040), .A2(n5039), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n5052) );
  NAND2_X1 U5335 ( .A1(n5042), .A2(n5041), .ZN(n5044) );
  XOR2_X1 U5336 ( .A(n5044), .B(n5043), .Z(n5047) );
  AOI222_X1 U5337 ( .A1(n5050), .A2(n5049), .B1(n5048), .B2(n5047), .C1(n5046), 
        .C2(n5045), .ZN(n5051) );
  OAI211_X1 U5338 ( .C1(n5054), .C2(n5053), .A(n5052), .B(n5051), .ZN(U3230)
         );
  AOI22_X1 U5339 ( .A1(n5055), .A2(n5059), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5058), .ZN(n5056) );
  OAI21_X1 U5340 ( .B1(n5058), .B2(n5057), .A(n5056), .ZN(U3261) );
  AOI22_X1 U5341 ( .A1(n5060), .A2(n5059), .B1(n5058), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5061) );
  OAI21_X1 U5342 ( .B1(n5058), .B2(n5062), .A(n5061), .ZN(U3260) );
endmodule

