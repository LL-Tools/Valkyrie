
module b20_C_2inp_gates_syn ( 
    P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
    P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
    P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
    P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
    P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
    P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
    P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
    P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
    P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
    P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
    P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
    P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
    P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
    P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
    P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
    P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
    P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
    P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465,
    P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486,
    P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507,
    P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
    P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
    P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
    P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
    P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
    P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
    P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554,
    P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
    P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
    P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
    P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
    P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290,
    P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283,
    P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276,
    P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269,
    P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377,
    P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257,
    P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250,
    P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243,
    P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236,
    P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402,
    P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423,
    P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444,
    P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452,
    P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459,
    P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466,
    P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473,
    P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480,
    P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487,
    P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230,
    P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223,
    P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216,
    P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491,
    P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498,
    P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505,
    P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
    P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
    P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179,
    P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
    P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
    P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
    P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150,
    P2_U3893  );
  input  P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
    P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
    P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
    P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
    P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
    P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
    P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
    P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
    P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
    P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
    P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
    P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
    P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
    P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
    P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
    P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
    P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
    P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465,
    P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486,
    P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507,
    P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
    P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
    P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
    P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
    P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
    P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
    P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554,
    P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
    P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
    P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
    P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
    P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290,
    P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283,
    P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276,
    P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269,
    P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377,
    P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257,
    P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250,
    P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243,
    P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236,
    P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402,
    P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423,
    P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444,
    P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452,
    P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459,
    P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466,
    P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473,
    P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480,
    P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487,
    P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230,
    P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223,
    P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216,
    P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491,
    P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498,
    P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505,
    P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
    P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
    P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179,
    P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
    P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
    P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
    P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150,
    P2_U3893;
  wire n11337, n11099, n14839, n10624, n10370, n15659, n17009, n15734,
    n13122, n11905, n11910, n10007, n9875, n10438, n8909, n10803, n12871,
    n13336, n10121, n12266, n12623, n10861, n8876, n8891, n14961, n16271,
    n10119, n12865, n13837, n15167, n9833, n15615, n16315, n11282, n12580,
    n14362, n12072, n11906, n16202, n11800, n16279, n11071, n16936, n9368,
    n9663, n9555, n11997, n11149, n10996, n9116, n8873, n10995, n10864,
    n8877, n8878, n8880, n16028, n12290, n16901, n10361, n10422, n8881,
    n13256, n8896, n9906, n9898, n8882, n12847, n13278, n8884, n8885,
    n10387, n8886, n8887, n10286, n9444, n9635, n9668, n9763, n16612,
    n16543, n9110, n16666, n9103, n16634, n9605, n9260, n9400, n14620,
    n15050, n9335, n9136, n9589, n11899, n9591, n9590, n14539, n12529,
    n13785, n9294, n9126, n11998, n9487, n13854, n14484, n14704, n9443,
    n16899, n9346, n9445, n16861, n12345, n9130, n14155, n14756, n14165,
    n11091, n13327, n9704, n14778, n12911, n14802, n9271, n14876, n14822,
    n15124, n15102, n13895, n10315, n13134, n9767, n9689, n13307, n15024,
    n15613, n10752, n14269, n16826, n11077, n15638, n8904, n16054, n16068,
    n12430, n16805, n15818, n15637, n9546, n15709, n14290, n10552, n10337,
    n17451, n16442, n9282, n15344, n16774, n16258, n15819, n12348, n17200,
    n13286, n13395, n15785, n15722, n15823, n13401, n13398, n13047, n13846,
    n15729, n17102, n15844, n11964, n15876, n17175, n11903, n16507, n11055,
    n9467, n17036, n9802, n16216, n16466, n12644, n17151, n9913, n17053,
    n11128, n13263, n9862, n15930, n9234, n16173, n9520, n9109, n11531,
    n12881, n12848, n9907, n11990, n12205, n8889, n8890, n11486, n17319,
    n16029, n9920, n11878, n9914, n10557, n10906, n11172, n10261, n12051,
    n9995, n11068, n10540, n11406, n10036, n11018, n10230, n10153, n10161,
    n9248, n16154, n11403, n8905, n10039, n11165, n17341, n17338, n9360,
    n17335, n11572, n9848, n10978, n10967, n9837, n11045, n9990, n9818,
    n10965, n10053, n10168, n9876, n9823, n9820, n9851, n9852, n9819,
    n9881, n9835, n9834, n13440, n13375, n9363, n9890, n9301, n8892, n8893,
    n10596, n16676, n8894, n8897, n12595, n9795, n10128, n10475, n14043,
    n12509, n16295, n12724, n9640, n13254, n12855, n9526, n13034, n9583,
    n9244, n9246, n9408, n15935, n9525, n9321, n12831, n12451, n14730,
    n11985, n13091, n9560, n11955, n9229, n11991, n9540, n12481, n9731,
    n9456, n11513, n9499, n9500, n12184, n12534, n17015, n9439, n9440,
    n9737, n9530, n9531, n10980, n9462, n9867, n10849, n11933, n9564,
    n14755, n14817, n9774, n9775, n9776, n11931, n11929, n9766, n10227,
    n10190, n13601, n13739, n12936, n12566, n9430, n9127, n9431, n14068,
    n17365, n9100, n11766, n9156, n9157, n10520, n9119, n9765, n15052,
    n9921, n12402, n9221, n9218, n15732, n9212, n9214, n13382, n13051,
    n9743, n9184, n9619, n9620, n9628, n9629, n9287, n13205, n9746, n9378,
    n12805, n9505, n9257, n9751, n9411, n9412, n9413, n11971, n9084, n9086,
    n12944, n10964, n9258, n9814, n9242, n9676, n9238, n9384, n9385, n9822,
    n9882, n9878, n9879, n9732, n9727, n9598, n9647, n9652, n9610, n9615,
    n9485, n9115, n9479, n9480, n9280, n9279, n9508, n9509, n9580, n9067,
    n12464, n13972, n12435, n12434, n9071, n9070, n9077, n12961, n12450,
    n12634, n12636, n17075, n9060, n9062, n10429, n11004, n11953, n13354,
    n9664, n9666, n9388, n9199, n13335, n9779, n13418, n11973, n15842,
    n11962, n9292, n15871, n9317, n9318, n9787, n9788, n9331, n9332,
    n10681, n10683, n10590, n10421, n9713, n12123, n9735, n9736, n9725,
    n9414, n9415, n9416, n12979, n9418, n9304, n9091, n9092, n9512, n9513,
    n9517, n11413, n11038, n9468, n9653, n9458, n9460, n9475, n9473, n9474,
    n9139, n16831, n9518, n12255, n11536, n11411, n11495, n17029, n11512,
    n17155, n13833, n13879, n12897, n17464, n9074, n10979, n11005, n9357,
    n11025, n9688, n9936, n14587, n10277, n9178, n9167, n9177, n15369,
    n9052, n9056, n10666, n9773, n9561, n9210, n9551, n15071, n9196, n9195,
    n15135, n9554, n14994, n9202, n11921, n15788, n9896, n10842, n9539,
    n9858, n16087, n9329, n10225, n10120, n10146, n16555, n9141, n13505,
    n9143, n9144, n14186, n13518, n9148, n13604, n13886, n12055, n9152,
    n11414, n16660, n9454, n16772, n16846, n16904, n11145, n16943, n11112,
    n11113, n9658, n14146, n13776, n13828, n13871, n13919, n9449, n9450,
    n13909, n14249, n14032, n14067, n9345, n11410, n9496, n16522, n9645,
    n13500, n12576, n9108, n9296, n17452, n11014, n9322, n10987, n9718,
    n9722, n10479, n9338, n9696, n9697, n14773, n14865, n15882, n15011,
    n14998, n14455, n10204, n10194, n14705, n13261, n9556, n9557, n9791,
    n14720, n15056, n10451, n10408, n13105, n15697, n9565, n10199, n9235,
    n9236, n15036, n13273, n9399, n9228, n9225, n16225, n12392, n11873,
    n14196, n16496, n13609, n13693, n16610, n9364, n17544, n17529, n12262,
    n11896, n17120, n12296, n10813, n9538, n9544, n10531, n15917, n17560,
    n11849, n17608, n13025, n13084, n9250, n13142, n9660, n12682, n9742,
    n13159, n12707, n9618, n9625, n9627, n9314, n13213, n9642, n9643,
    n9373, n9376, n9528, n9423, n9504, n9350, n9351, n12914, n12862, n9529,
    n9348, n9255, n9259, n9753, n10658, n12971, n9410, n9082, n9638,
    n12471, n12472, n12431, n9681, n9247, n9669, n9197, n9201, n9670,
    n9671, n13412, n13292, n9545, n10234, n9522, n12122, n9419, n9420,
    n9421, n11040, n9457, n9435, n9516, n9495, n9507, n9576, n12920,
    n12919, n9447, n12912, n9584, n9585, n9441, n9437, n9438, n12606,
    n17096, n9738, n9534, n9535, n10966, n9702, n9865, n9169, n9172, n9176,
    n9173, n9174, n9694, n9175, n9761, n9053, n9057, n13323, n13236,
    n13242, n14744, n13343, n9569, n9571, n14889, n9240, n9243, n14909,
    n14936, n9203, n9204, n9205, n9206, n15616, n9673, n9237, n9394, n9395,
    n9796, n13414, n9261, n15725, n15763, n10522, n10442, n9381, n9382,
    n9824, n9847, n10150, n10049, n10148, n10125, n9521, n9734, n9145,
    n9716, n9717, n9146, n9147, n9728, n11471, n9506, n11534, n16645,
    n16665, n9290, n9275, n9273, n11133, n9359, n9649, n9455, n9616, n9483,
    n9482, n11142, n9133, n9477, n9476, n9276, n12358, n9432, n9124, n9125,
    n12314, n9514, n9515, n12234, n12220, n11590, n11438, n12506, n11581,
    n9061, n9646, n9065, n13753, n9063, n9066, n13835, n13924, n12511,
    n13948, n13996, n9069, n14099, n9075, n9076, n9343, n14125, n16987,
    n12443, n17081, n12497, n9102, n17126, n17129, n10973, n10976, n9719,
    n9720, n9721, n10436, n9121, n10471, n11072, n11024, n11031, n9698,
    n10725, n9165, n9166, n10795, n10863, n13369, n9324, n10106, n13367,
    n9559, n9792, n13349, n9219, n9220, n9222, n9223, n10827, n14801,
    n9567, n9568, n10764, n10627, n13173, n10600, n14938, n9552, n10455,
    n16304, n9562, n9783, n9784, n9215, n9406, n13285, n15974, n9316,
    n13012, n9558, n9793, n9794, n14731, n14779, n15082, n14815, n9390,
    n14923, n14970, n15643, n11920, n15786, n9549, n9230, n13282, n9045,
    n9044, n9901, n9902, n10935, n9874, n9871, n9843, n10648, n10652,
    n9690, n9691, n10551, n10224, n12161, n9160, n14231, n13533, n12203,
    n12053, n14258, n11781, n12226, n13862, n16580, n13691, n9724, n12987,
    n9094, n9087, n9088, n12289, n14050, n13644, n9428, n16638, n9630,
    n9631, n9633, n16697, n16722, n9465, n16735, n16758, n16792, n9263,
    n9471, n9470, n11139, n16849, n9268, n9269, n9272, n16922, n9593,
    n9594, n9595, n9592, n13740, n12313, n12298, n14221, n12215, n13961,
    n14008, n17463, n11493, n17166, n17147, n14142, n13880, n13970, n9095,
    n9096, n17422, n17414, n12584, n12869, n12841, n9059, n9073, n9622,
    n9623, n9463, n9464, n11013, n9104, n9541, n9543, n9047, n9050, n16768,
    n11069, n12077, n9137, n9323, n15268, n10917, n9162, n14446, n14449,
    n9708, n9709, n9693, n14553, n9707, n14570, n16094, n15347, n9758,
    n15012, n14457, n10081, n9956, n10167, n10237, n9772, n15022, n9208,
    n10341, n9563, n15708, n15746, n10200, n15975, n15977, n15968, n15992,
    n15043, n9771, n14982, n10006, n15233, n9043, n9036, n9040, n9041,
    n9042, n9046, n11868, n15431, n17219, n10332, n10030, n12066, n9403,
    n13931, n16473, n14175, n13560, n9726, n13607, n13655, n16574, n9149,
    n9151, n9150, n16609, n13707, n17547, n17541, n17538, n9511, n17535,
    n17532, n17522, n17519, n17516, n13904, n14270, n14291, n17465, n9099,
    n9574, n16756, n16917, n9657, n14136, n13805, n13801, n13824, n14061,
    n14094, n17196, n11504, n9498, n11561, n17197, n13501, n14150, n17350,
    n11405, n15241, n11407, n17214, n11323, n17232, n11003, n17243, n9337,
    n17307, n17325, n16135, n9342, n15254, n14721, n14924, n10537, n15381,
    n14610, n10561, n10792, n9319, n9320, n15333, n16415, n16412, n16409,
    n16406, n16403, n16400, n16394, n16391, n16388, n13151, n15661, n15711,
    n9306, n9310, n15035, n14706, n12006, n15695, n9566, n16004, n9398,
    n15076, n15232, n9037, n9039, n9038, n17562, n17558, n11851, n17604,
    n17596, n9186, n9134, n9135, n9295, n15737, n8898, n8899, n8900,
    n15674, n8901, n8902, n8903, n8906, n8907, n8908, n13419, n11940,
    n10720, n13283, n13149, n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n13855, n13998, n11458, n8917, n8918, n8919, n8920, n8921,
    n12303, n8922, n9899, n8923, n16292, n9297, n10124, n8924, n9200,
    n16227, n8925, n8926, n12985, n9417, n8927, n9325, n14741, n14835,
    n14072, n14908, n14960, n14887, n9198, n10482, n8928, n8929, n8930,
    n14997, n8931, n8932, n9782, n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n10611, n10682, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n9699, n8951, n8952, n8953, n8954, n8955,
    n8956, n10292, n9828, n9665, n8957, n8958, n8959, n8960, n8961, n9459,
    n15092, n9433, n9434, n8962, n9581, n9582, n8963, n9570, n14559, n9305,
    n8964, n12263, n11058, n9356, n8965, n10716, n9051, n8966, n8967,
    n8968, n8969, n8970, n17330, n8971, n8972, n13397, n8973, n8974,
    n12399, n8975, n8976, n8977, n9872, n8978, n8979, n8980, n15157, n9049,
    n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n15061, n8993, n8994, n8995, n8996, n8997, n8998, n12594,
    n13179, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n12692, n9344, n9010, n9011, n9012, n9756, n9013, n9014,
    n9015, n9714, n12173, n9016, n10545, n9017, n9018, n9692, n13009,
    n9019, n17051, n15007, n9020, n9501, n9502, n9021, n9022, n9510, n9608,
    n9497, n9023, n17449, n9107, n9024, n9025, n9026, n9027, n9028, n9596,
    n17238, n13376, n16034, n9494, n9029, n17294, n9307, n9030, n9031,
    n9032, n9033, n9034, n16385, n16165, n16008, n9527, n17205, n12808,
    n16338, n9035, n9048, n10750, n10718, n9054, n9055, n9058, n12842,
    n12484, n17097, n12444, n9579, n13752, n9064, n9575, n13770, n9586,
    n9068, n13995, n9452, n9072, n9078, n9079, n12935, n9080, n9081, n9083,
    n9085, n9089, n9090, n9093, n12992, n9098, n12910, n9097, n9101, n9429,
    n10981, n9105, n9106, n13748, n9111, n9112, n9113, n16844, n9114,
    n9603, n9117, n10437, n9118, n9120, n9122, n9123, n9129, n9131, n9128,
    n16881, n9132, n11051, n9138, n11023, n16787, n11136, n9140, n12344,
    n12321, n9142, n16581, n9153, n9155, n9154, n11001, n9158, n16459,
    n16458, n9159, n9161, n9164, n9163, n12020, n10747, n9170, n14571,
    n9168, n10738, n10646, n9171, n14409, n10305, n9181, n9179, n12860,
    n9180, n9182, n9183, n9617, n9187, n9185, n9191, n9188, n9189, n9190,
    n12753, n12740, n9192, n9389, n9193, n9194, n15614, n9207, n9213,
    n9216, n9209, n9211, n9786, n9785, n9409, n15969, n11907, n9217,
    n14767, n9224, n9226, n9227, n9233, n9232, n9231, n9239, n9241, n9245,
    n14947, n11976, n11981, n9680, n9402, n9252, n9249, n13082, n9251,
    n15889, n9253, n9254, n9256, n13258, n16940, n9262, n16751, n9264,
    n16789, n9265, n9266, n9267, n9270, n11043, n11050, n16693, n9274,
    n9277, n11107, n9278, n9341, n9745, n9281, n9391, n9349, n13042, n9283,
    n10054, n16182, n9953, n9284, n9285, n13190, n9286, n9573, n11028,
    n9288, n9339, n9291, n9289, n13036, n11150, n16864, n11124, n16662,
    n17343, n9358, n13126, n9299, n15872, n9293, n12838, n9759, n12894,
    n12893, n9532, n13039, n14863, n13007, n13136, n13760, n13755, n13054,
    n9300, n13406, n9983, n14382, n10257, n9503, n12244, n12267, n13031,
    n9298, n9302, n13423, n12898, n12924, n9436, n12918, n9957, n9427,
    n12946, n10085, n9405, n9798, n9880, n9303, n13448, n15678, n14467,
    n17058, n17168, n9315, n9404, n15892, n15745, n12401, n13023, n13085,
    n10382, n10824, n9374, n15346, n9492, n12602, n9308, n17167, n9353,
    n10677, n13052, n9309, n10358, n9311, n9312, n10702, n9313, n9748,
    n13422, n16828, n11111, n9939, n9930, n14995, n12409, n9868, n14633,
    n13148, n9553, n9973, n9996, n13099, n13314, n9599, n16714, n9326,
    n9347, n17174, n9396, n9407, n10283, n9327, n9328, n9372, n9426, n9362,
    n11974, n13040, n10226, n16962, n12504, n17127, n10285, n9330, n9686,
    n12021, n9334, n9684, n13623, n9672, n9386, n9962, n9333, n9695,
    n17154, n9710, n16590, n17259, n9706, n9519, n13264, n9655, n13269,
    n9336, n9369, n9840, n9355, n9340, n12129, n11120, n9685, n10483,
    n11129, n13313, n9760, n13309, n13161, n9352, n9747, n9354, n9361,
    n9611, n9639, n13491, n9370, n9894, n9764, n9365, n9366, n9367, n9998,
    n9972, n10326, n10157, n10191, n9371, n12826, n9375, n9377, n9379,
    n9383, n9380, n10389, n9387, n11947, n9392, n9397, n9393, n15660,
    n15639, n15195, n15193, n9401, n15813, n15794, n9422, n9424, n9425,
    n17141, n17143, n12494, n17388, n9442, n17027, n9446, n9448, n9451,
    n12514, n13941, n11809, n11201, n9453, n9461, n9469, n9466, n16705,
    n16816, n9472, n16942, n9478, n9481, n16868, n9484, n9486, n12863,
    n9488, n9489, n9490, n9491, n9606, n9493, n12299, n10045, n10073,
    n10123, n12090, n9938, n9886, n9523, n9524, n9533, n9536, n9537,
    n10815, n10783, n9542, n10685, n15884, n9547, n9548, n9550, n14984,
    n14703, n14875, n9572, n13729, n12483, n9577, n9578, n12476, n13834,
    n9587, n9588, n11153, n16738, n9597, n11132, n9600, n16696, n9601,
    n9602, n9604, n16821, n9607, n9609, n16683, n9614, n9612, n9613, n9621,
    n9624, n9626, n16639, n9632, n9634, n9636, n9637, n9641, n9644, n9651,
    n16741, n9648, n9650, n16718, n11118, n9654, n9656, n9659, n12675,
    n9661, n9662, n14837, n9667, n9678, n9674, n15644, n9675, n9677, n9679,
    n15710, n14742, n9682, n9683, n9687, n11298, n10145, n14468, n14556,
    n9700, n9701, n9703, n14447, n9705, n10189, n11721, n13586, n9711,
    n9712, n9715, n10990, n10968, n9723, n9733, n9729, n9730, n13547,
    n11728, n11730, n9739, n9740, n9741, n9744, n13221, n9749, n9750,
    n9752, n9754, n9755, n9757, n10262, n9762, n10001, n10476, n12213,
    n9769, n9768, n9870, n11935, n9770, n14981, n9777, n14860, n9778,
    n9780, n9781, n15793, n15758, n9849, n9789, n9790, n9799, n9797,
    n12311, n10823, n9800, n9801, n9803, n9804, n9805, n9806, n9807, n9808,
    n11081, n13390, n9809, n9810, n9811, n9812, n9813, n9815, n9816, n9817,
    n13459, n11923, n11943, n10322, n11948, n10433, n10325, n11017, n12086,
    n11185, n12233, n12438, n12887, n17172, n12398, n10705, n10564, n9827,
    n15178, n12012, n10717, n10528, n13638, n16539, n12221, n13932, n12969,
    n16993, n17083, n17373, n17356, n14972, n14622, n14891, n14625, n14679,
    n10108, n16170, n10156, n16605, n17185, n13719, n10918, n10761, n10268,
    n10612, n16616, n16542, n13625, n16573, n16618, n13951, n16949, n17396,
    n11772, n15311, n12394, n11837, n16577, n16595, n17551, n14097, n17349,
    n15361, n15376, n16418, n16397, n15640, n15896, n15991, n11847, n11853,
    n10956, n17564, n17600, n9821, n9826, n9825, n9829, n10446, n9830,
    n9831, n10556, n9832, n11959, n9836, n9845, n9838, n9839, n9841,
    n14848, n9842, n9844, n9846, n11802, n9850, n16009, n9857, n9853,
    n9854, n9855, n9856, n16015, n11296, n9863, n13477, n9860, n9859,
    n9861, n10905, n13484, n10500, n9864, n9866, n13008, n9869, n9873,
    n15386, n9877, n16148, n9893, n9883, n9885, n9884, n9887, n9888, n9994,
    n9889, n9891, n12056, n9892, n11909, n10164, n9895, n11908, n16193,
    n9916, n9897, n15236, n9900, n9904, n9903, n9905, n9909, n9910, n9908,
    n9912, n9911, n10118, n10093, n9915, n9917, n9967, n9919, n10013,
    n9918, n9968, n15345, n15423, n9924, n9922, n11316, n9923, n9926,
    n9925, n9928, n9927, n9929, n15980, n9931, n11604, n9935, n9933, n9932,
    n9934, n11720, n9937, n9941, n9940, n12043, n17342, n9949, n9947,
    n9942, n9945, n9943, n9944, n9946, n16155, n9948, n9952, n9950, n9951,
    n9959, n9954, n9955, n9958, n9960, n9961, n9964, n9963, n9966, n9965,
    n11300, n9970, n9969, n9971, n9997, n9974, n9975, n16142, n9977, n9985,
    n9980, n9978, n9979, n9982, n9981, n9984, n9986, n10019, n9988, n9987,
    n10020, n15266, n15307, n9989, n9993, n9991, n16136, n9992, n10000,
    n9999, n10035, n10003, n10002, n10071, n10004, n10005, n10015, n10008,
    n10009, n15865, n10011, n10010, n10012, n10014, n10016, n10024, n10018,
    n10017, n10025, n15308, n10022, n10021, n15306, n10023, n10028, n10026,
    n10027, n10029, n10034, n10067, n10031, n10032, n15477, n10033, n10052,
    n10074, n10038, n10037, n10046, n10076, n10043, n10041, n10040, n10042,
    n10044, n10048, n10047, n10050, n10051, n10062, n10056, n15380, n10055,
    n10060, n10058, n10057, n10059, n10061, n10063, n10099, n10065, n10064,
    n10100, n15373, n10066, n10070, n10068, n16128, n10069, n10079, n10072,
    n10075, n10077, n16127, n10078, n10091, n10080, n10089, n10083, n10082,
    n10084, n15858, n10087, n10086, n10088, n10090, n10092, n15368, n10095,
    n10094, n15366, n10096, n10097, n10098, n10103, n10102, n10101, n15372,
    n10104, n10105, n10117, n10107, n10113, n10109, n10111, n10110, n10112,
    n15781, n10115, n10114, n10116, n10138, n10122, n10147, n10126, n10127,
    n17312, n10136, n10129, n10134, n10130, n10131, n10132, n11672, n10133,
    n10135, n10137, n10139, n10144, n10141, n10140, n10143, n15251, n10142,
    n15250, n15284, n10149, n10151, n10152, n10154, n10155, n10159, n10158,
    n10160, n10162, n10163, n17300, n10173, n10193, n10165, n10171, n10166,
    n10236, n10169, n11717, n10170, n10172, n10185, n10179, n10174, n11711,
    n10176, n10175, n15741, n10177, n10178, n10183, n10181, n10180, n10182,
    n15771, n10184, n10186, n15328, n10188, n10187, n10216, n10214, n17306,
    n10192, n10197, n10195, n11699, n10196, n10198, n10209, n10203, n15754,
    n10201, n10202, n10207, n10205, n10206, n10208, n10210, n15324, n10212,
    n10211, n15322, n10213, n10215, n10223, n15285, n15286, n10217, n15327,
    n10218, n10221, n10219, n10220, n10222, n14395, n10229, n10228, n10320,
    n10232, n10231, n10233, n10323, n10235, n10321, n10284, n10245, n10264,
    n10238, n10239, n10240, n16095, n10243, n10241, n10242, n10244, n10850,
    n10251, n10246, n14597, n10248, n10247, n15691, n10249, n10250, n10255,
    n10253, n10252, n10254, n10256, n10258, n10309, n10260, n10259, n10310,
    n14591, n10263, n10266, n16101, n10265, n10267, n10271, n15705, n10269,
    n10270, n10275, n10273, n10272, n10274, n10276, n10278, n10280, n10279,
    n14585, n10281, n10282, n10290, n10288, n10287, n10327, n10289, n10324,
    n10297, n10291, n10295, n10293, n16088, n10294, n10296, n10299, n15656,
    n14454, n10298, n10303, n10301, n10300, n10302, n10304, n10316, n10307,
    n10306, n10317, n10314, n10308, n10313, n10312, n10311, n14590, n10319,
    n10318, n14448, n10419, n10329, n10328, n10362, n10359, n10330, n17276,
    n10331, n10335, n10333, n16081, n10334, n10336, n10350, n10344, n10339,
    n10338, n10342, n10340, n15634, n14558, n10343, n10348, n10346, n10345,
    n10347, n10349, n10351, n10354, n10353, n10352, n10355, n14554, n10357,
    n10356, n10360, n10426, n10420, n10364, n10363, n10430, n10423, n10365,
    n12157, n10366, n10368, n10395, n16075, n10367, n10369, n10378, n10372,
    n10404, n15610, n14372, n10371, n10376, n10374, n10373, n10375, n10377,
    n10379, n10383, n14367, n10381, n10380, n14370, n10386, n10385, n10384,
    n14368, n10388, n10391, n10390, n10392, n10401, n10393, n10399, n10394,
    n10396, n10397, n16069, n10398, n10400, n10415, n10403, n10402, n10413,
    n10406, n10405, n10409, n10407, n15025, n10411, n10410, n10412, n10414,
    n10416, n14481, n10418, n10417, n10507, n10466, n10424, n10425, n10427,
    n10428, n10432, n10431, n10435, n10434, n10440, n10439, n10441, n10477,
    n10443, n10444, n10445, n10449, n10447, n16062, n10448, n10450, n10462,
    n10453, n10452, n10460, n10454, n10456, n14987, n10458, n10457, n10459,
    n10461, n10463, n10503, n10465, n10464, n10504, n14486, n10467, n10512,
    n10469, n10468, n10470, n10519, n10472, n10473, n10474, n10480, n10478,
    n10489, n10481, n10487, n10484, n10485, n16056, n10486, n10488, n10498,
    n10490, n14962, n10492, n10491, n10496, n10494, n10493, n10495, n10497,
    n10499, n10513, n10502, n10501, n10514, n14503, n10506, n10505, n14501,
    n10510, n14483, n14636, n10508, n10509, n10511, n10516, n10515, n14504,
    n10518, n10517, n10523, n10553, n10521, n10524, n10526, n10525, n10527,
    n10615, n10529, n10530, n17248, n10535, n10532, n10534, n10536, n10547,
    n10539, n10538, n10544, n14925, n10542, n10541, n10543, n10546, n10548,
    n14413, n10550, n10549, n14412, n14415, n10554, n17253, n10555, n10559,
    n16049, n10558, n10560, n10571, n10563, n10562, n10569, n10565, n14939,
    n10567, n10566, n10568, n10570, n10572, n10577, n10574, n10573, n10578,
    n10575, n10576, n14408, n14607, n10580, n10579, n10581, n10584, n10582,
    n10583, n10585, n10586, n10593, n10588, n10587, n10589, n10614, n10591,
    n10613, n10592, n10594, n10595, n10607, n10598, n10597, n10605, n10599,
    n10601, n14898, n10603, n10602, n10604, n10606, n10608, n10641, n10610,
    n10609, n10640, n14428, n10618, n10617, n10616, n10621, n10620, n10619,
    n10647, n10650, n10622, n10623, n15113, n10634, n10626, n10625, n10632,
    n10628, n14877, n10630, n10629, n10631, n10633, n10635, n14432, n10638,
    n10637, n10636, n10639, n14431, n10644, n10642, n14430, n10643, n10645,
    n10649, n10654, n10653, n10651, n10656, n10655, n10657, n10686, n10659,
    n10660, n10684, n10663, n10661, n10662, n10673, n10665, n10664, n10671,
    n10667, n14851, n10669, n10668, n10670, n10672, n10674, n10678, n10676,
    n10675, n14572, n10679, n10680, n10688, n10687, n10690, n10689, n10693,
    n10691, n10692, n10695, n10694, n10697, n10696, n10751, n10698, n10699,
    n10748, n10700, n10701, n10712, n10704, n10703, n10710, n10706, n14803,
    n10708, n10707, n10709, n10711, n10713, n10741, n10715, n10714, n10742,
    n14524, n10719, n16021, n10722, n16022, n10721, n10732, n10724, n10723,
    n10730, n10726, n14824, n10728, n10727, n10729, n10731, n10733, n14520,
    n10735, n10734, n14518, n10736, n10737, n14517, n10739, n10740, n10745,
    n10744, n10743, n14523, n10746, n10749, n10754, n10753, n10756, n10755,
    n10784, n10757, n10758, n10781, n17213, n10759, n10760, n10771, n10763,
    n10762, n10769, n10765, n14781, n10767, n10766, n10768, n10770, n10772,
    n10776, n10774, n10773, n10777, n10775, n10780, n10778, n10779, n14466,
    n10782, n10786, n10785, n10788, n10787, n10814, n10789, n10790, n10811,
    n11804, n10791, n10802, n10794, n10793, n10800, n10796, n14757, n10798,
    n10797, n10799, n10801, n10804, n10807, n10806, n10805, n10808, n14621,
    n10809, n10810, n10812, n10817, n10816, n10819, n10818, n10843, n10820,
    n10821, n10840, n11814, n10822, n10833, n10826, n10825, n10831, n10853,
    n14722, n10829, n10828, n10830, n10832, n10834, n10838, n10836, n10835,
    n10837, n10839, n12019, n10841, n10845, n10844, n10846, n11869, n10847,
    n11866, n11825, n10848, n10860, n10852, n10851, n10858, n12023, n10936,
    n10854, n12001, n10856, n10855, n10857, n10859, n10862, n10868, n10866,
    n10865, n10867, n10915, n10920, n16174, n16329, n10927, n10912, n10869,
    n10871, n10870, n10872, n16007, n10878, n10876, n10874, n10873, n10875,
    n10877, n10894, n10880, n10879, n10884, n10882, n10881, n10883, n10892,
    n10886, n10885, n10890, n10888, n10887, n10889, n10891, n10893, n10899,
    n10896, n10895, n10897, n10898, n10900, n10901, n12010, n10902, n16166,
    n10903, n16162, n10904, n10934, n10907, n10909, n10908, n13383, n11600,
    n10910, n10921, n10911, n15293, n10913, n10914, n10957, n10916, n10955,
    n10919, n10954, n15902, n10923, n10922, n10952, n13479, n10924, n10926,
    n10925, n12009, n10928, n10929, n11304, n10933, n11958, n10930, n13483,
    n10931, n10932, n11302, n10950, n10946, n15319, n10939, n13013, n10937,
    n10938, n10943, n10941, n10940, n10942, n16421, n10945, n10944, n10948,
    n15426, n15332, n10947, n10949, n10951, n10953, n10958, n10959, n10960,
    n10972, n11765, n11102, n10961, n10962, n11007, n10992, n10963, n11009,
    n10969, n10970, n10971, n10974, n10975, n10977, n10982, n10984, n10983,
    n10985, n10989, n10986, n10988, n10991, n12999, n11289, n10994, n10993,
    n10998, n10997, n10999, n11020, n11000, n11002, n11074, n11006, n11089,
    n11008, n11010, n12892, n11011, n12993, n11292, n11012, n11015, n11016,
    n12179, n11019, n11021, n17254, n11115, n11265, n11251, n11234, n11022,
    n11225, n16984, n11027, n11026, n11029, n11030, n11034, n11032, n11033,
    n11036, n11035, n16625, n11037, n11039, n11041, n11044, n11042, n12064,
    n11047, n11046, n11049, n11048, n16694, n11054, n11053, n11052, n11056,
    n17070, n11057, n11063, n11059, n11062, n11060, n11061, n11064, n16731,
    n11186, n11065, n11066, n16740, n11067, n11197, n11193, n17022, n11070,
    n16777, n11073, n11211, n11078, n11075, n11217, n17295, n16822, n11076,
    n11079, n11080, n11082, n11221, n17289, n11085, n11083, n11084, n11231,
    n17283, n11087, n11086, n11088, n11093, n11090, n11238, n17277, n11092,
    n11243, n11095, n11094, n11096, n11105, n16888, n17271, n16883, n11097,
    n11098, n12165, n17266, n11100, n11259, n11101, n11103, n11104, n11108,
    n17260, n16919, n16925, n11106, n11109, n11110, n12185, n16948, n11888,
    n13958, n11114, n11898, n11116, n11117, n11281, n11833, n16628, n16939,
    n16862, n11154, n11252, n16865, n16937, n11283, n11152, n11897, n11148,
    n16916, n11144, n16880, n11141, n16843, n11138, n16804, n17301, n11135,
    n16775, n17313, n11119, n11121, n11122, n16663, n11123, n11125, n11126,
    n11173, n11127, n16737, n11130, n11131, n11134, n11137, n11140, n11143,
    n11147, n11146, n11151, n11156, n11155, n11157, n11158, n11161, n11160,
    n11159, n16629, n16644, n16643, n16658, n11163, n11162, n11164, n16657,
    n11166, n11167, n16681, n11169, n11168, n11170, n16680, n11171, n12994,
    n17115, n11175, n11174, n11176, n11179, n11177, n16701, n11178, n16704,
    n11181, n16713, n11180, n11182, n11184, n11183, n16723, n11189, n11187,
    n11188, n11190, n16734, n11191, n11192, n11196, n11194, n11195, n11198,
    n16755, n11199, n11200, n11204, n11202, n11203, n11205, n16771, n11206,
    n11207, n11210, n11208, n11209, n11212, n16791, n11213, n11214, n11216,
    n11215, n11218, n16814, n11220, n11219, n16813, n11224, n11222, n11223,
    n11226, n16830, n11227, n11228, n11230, n11229, n11232, n16848, n11233,
    n11237, n11235, n11236, n11239, n16867, n11242, n11240, n11241, n16886,
    n11246, n11244, n11245, n11247, n16885, n11250, n11248, n11249, n11255,
    n11253, n11254, n11256, n16903, n11257, n11258, n11262, n11260, n11261,
    n11263, n16921, n11264, n11268, n11266, n11267, n11269, n16941, n11272,
    n11270, n11271, n11276, n11275, n11274, n11277, n11884, n11279, n11278,
    n11883, n11280, n11287, n11285, n11284, n11286, n11288, n12995, n16817,
    n16945, n11290, n11294, n11822, n11291, n11293, n16924, n11770, n11295,
    n13535, n11297, n11299, n11301, n11306, n11303, n15355, n11305, n11312,
    n11308, n13035, n11307, n11310, n15360, n11309, n11311, n11313, n11787,
    n11315, n11314, n11318, n11317, n11830, n11322, n11320, n17226, n12071,
    n11319, n11321, n11368, n11326, n11325, n17348, n11374, n11327, n11328,
    n11329, n11330, n11331, n11332, n11334, n11333, n11336, n11335, n11339,
    n11338, n11341, n11340, n11343, n11342, n11977, n11345, n11344, n11347,
    n11346, n11349, n11348, n11351, n11350, n11353, n11352, n11355, n11354,
    n11357, n11356, n15618, n11359, n11358, n11361, n11360, n11363, n11362,
    n11365, n11364, n11367, n11366, n11373, n11371, n11369, n11370, n11372,
    n11397, n11375, n11376, n11377, n11378, n11732, n11379, n11380, n11381,
    n11382, n11383, n11384, n11731, n11385, n11386, n11387, n11388, n11389,
    n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11402, n11398,
    n11400, n11399, n11401, n11404, n14354, n12327, n11409, n12216, n11408,
    n11418, n12219, n11412, n16958, n11416, n11415, n11417, n14116, n11420,
    n17550, n11419, n11422, n11421, n11426, n11424, n11423, n11425, n11428,
    n11427, n11430, n11429, n11435, n11433, n11563, n17071, n11431, n11432,
    n11434, n11437, n11436, n11580, n11470, n13574, n11448, n11439, n14009,
    n11441, n11440, n11445, n11443, n11442, n11444, n11447, n11446, n11449,
    n13984, n11455, n11451, n11450, n11453, n11452, n11454, n14259, n11457,
    n11456, n11459, n17112, n11461, n11460, n11465, n11463, n11462, n11464,
    n17132, n11467, n11466, n11469, n11468, n11476, n11472, n14076, n11474,
    n11473, n11475, n11478, n11477, n11480, n11479, n11482, n11481, n11484,
    n11483, n11485, n11488, n11487, n11490, n11489, n11492, n11491, n11499,
    n11497, n11494, n16449, n11496, n11498, n16989, n11501, n11500, n11503,
    n11502, n11509, n11507, n17046, n11505, n11506, n11508, n11511, n11510,
    n11516, n11514, n17019, n11515, n11520, n11518, n11517, n11519, n11522,
    n11521, n11524, n11523, n11526, n11525, n11528, n14033, n11527, n14280,
    n11530, n11529, n11533, n11532, n11540, n11535, n14053, n11538, n11537,
    n11539, n11542, n11541, n11544, n11543, n11548, n11546, n11545, n11547,
    n17150, n11550, n11549, n13677, n12256, n11556, n11552, n11551, n11554,
    n11553, n11555, n13926, n11558, n11557, n11560, n11559, n11567, n11565,
    n17065, n11562, n11564, n11566, n17078, n11569, n11568, n11571, n11570,
    n11577, n11575, n16983, n11573, n11574, n11576, n11579, n11578, n16510,
    n11583, n11582, n11587, n11585, n11584, n11586, n16974, n11589, n11588,
    n13933, n11596, n11592, n11591, n11594, n11593, n11595, n11598, n11597,
    n14397, n11599, n11631, n16026, n11601, n11630, n11602, n15607, n11603,
    n11658, n14650, n15408, n15407, n15406, n11605, n15416, n15417, n11607,
    n11606, n11676, n11608, n11677, n11610, n11609, n15445, n11611, n15446,
    n11613, n11612, n15470, n11614, n15471, n11616, n11615, n15478, n11617,
    n15479, n11619, n11618, n11662, n11620, n11663, n11622, n11621, n11689,
    n11623, n11690, n11625, n11624, n11707, n16107, n11626, n11628, n11627,
    n11706, n11705, n11629, n14651, n11632, n15392, n15432, n15591, n11656,
    n14676, n15399, n15995, n15400, n11634, n11633, n15438, n15437, n11636,
    n11635, n11679, n11637, n11680, n11639, n11638, n15453, n15452, n11641,
    n11640, n15460, n15459, n11643, n11642, n15485, n15486, n11645, n16122,
    n15825, n11644, n11665, n11666, n11647, n16117, n15780, n11646, n11692,
    n11693, n11650, n16112, n11648, n11649, n11702, n11652, n11651, n11703,
    n11653, n14677, n11654, n13482, n15596, n15574, n11655, n11657, n11660,
    n15604, n11659, n15258, n11661, n11671, n11664, n11669, n11667, n11668,
    n11670, n11674, n11673, n15272, n11675, n11685, n11678, n11683, n11681,
    n11682, n11684, n11687, n11686, n15278, n11688, n11698, n11691, n11696,
    n11694, n11695, n11697, n11701, n11700, n11704, n11716, n11709, n11708,
    n11710, n11714, n15320, n11712, n11713, n11715, n11719, n11718, n11727,
    n15434, n11725, n15358, n11723, n11722, n11724, n11726, n11729, n12034,
    n11738, n11736, n11734, n11733, n11735, n11737, n11754, n11740, n11739,
    n11744, n11742, n11741, n11743, n11752, n11746, n11745, n11750, n11748,
    n11747, n11749, n11751, n11753, n11759, n11756, n11755, n11757, n11758,
    n11760, n11761, n12552, n11764, n11763, n11762, n12585, n12488, n11767,
    n11782, n11777, n12896, n12557, n11775, n11768, n11769, n12583, n12575,
    n12895, n11771, n11783, n11773, n11774, n11776, n11778, n11780, n12997,
    n11779, n16601, n11799, n11795, n12581, n11786, n11784, n11785, n11789,
    n11788, n17195, n17171, n11790, n17358, n11794, n11791, n11792, n13492,
    n11793, n11797, n12335, n12544, n17204, n11796, n11798, n11801, n16134,
    n11808, n11803, n11806, n16023, n11805, n11807, n11813, n11811, n11810,
    n11812, n11819, n11818, n11816, n11815, n11817, n11824, n11820, n11821,
    n11823, n11831, n11829, n11827, n11826, n11828, n11835, n11832, n11834,
    n17573, n17578, n17577, n17582, n17581, n17586, n17585, n17590, n17589,
    n17594, n17593, n17598, n17597, n17602, n17601, n17606, n17605, n11854,
    n11852, n11850, n11848, n11846, n11844, n11842, n17570, n11840, n11836,
    n17555, n17554, n11838, n17572, n17571, n11839, n17569, n11841, n17568,
    n17567, n11843, n17566, n17565, n11845, n17563, n17561, n17559, n17557,
    n11855, n11856, n11857, n11858, n17592, n11859, n17588, n11860, n17584,
    n11861, n17580, n11862, n17575, n17574, n11863, n11865, n11864, n11867,
    n11871, n11870, n12839, n11872, n11877, n11875, n12405, n11874, n11876,
    n11882, n11880, n11879, n11881, n11886, n11885, n11892, n11887, n11890,
    n11889, n11891, n11895, n13678, n11893, n11894, n11900, n11902, n11901,
    n13352, n13319, n11904, n15908, n15890, n15966, n15907, n13393, n11911,
    n15723, n11912, n15814, n11914, n15801, n11913, n11915, n11917, n11963,
    n11916, n15795, n11918, n13075, n11968, n14399, n13294, n11919, n15318,
    n15677, n11922, n11924, n11925, n11926, n11927, n11928, n11930, n11932,
    n11934, n14937, n11936, n15146, n11937, n14951, n11938, n11939, n14866,
    n11941, n11942, n11944, n11945, n11946, n14813, n11950, n11949, n14792,
    n11951, n11952, n11954, n11956, n11957, n12379, n15998, n11960, n11961,
    n15983, n15853, n12008, n15993, n15904, n13402, n15790, n15759, n11966,
    n11965, n11967, n15757, n15760, n11969, n13076, n11970, n13409, n11972,
    n13298, n13416, n13426, n13427, n15009, n13432, n11975, n14946, n13310,
    n11978, n13438, n14935, n11979, n13446, n13325, n13326, n14861, n13330,
    n13338, n14814, n11980, n14768, n13341, n14793, n13455, n11983, n14743,
    n13346, n11982, n11984, n13460, n11986, n13351, n11989, n11988, n11987,
    n11995, n15933, n11993, n15979, n15875, n11992, n11994, n12383, n15931,
    n15924, n11996, n14921, n11999, n16327, n12000, n12381, n12005, n15927,
    n12003, n16000, n12002, n12004, n12007, n12016, n12011, n12389, n12014,
    n12386, n12013, n12015, n12018, n15961, n12017, n12022, n12033, n12031,
    n12029, n12025, n12024, n12027, n12026, n12028, n12030, n12032, n12035,
    n12036, n12536, n12038, n12037, n12039, n12040, n12047, n12041, n12042,
    n12045, n12044, n12046, n12049, n12048, n12050, n12052, n17353, n16495,
    n12054, n16594, n12060, n12058, n12057, n12059, n12061, n16593, n12062,
    n12063, n12065, n16141, n12067, n12070, n12068, n12069, n16460, n12074,
    n12073, n12076, n12075, n17389, n12082, n16538, n12079, n12078, n12081,
    n12080, n12084, n16531, n12083, n16528, n12085, n12087, n12089, n12088,
    n12092, n17318, n12091, n17062, n12093, n12096, n12094, n12095, n16608,
    n12101, n12097, n12099, n12098, n12100, n12119, n16477, n12106, n12102,
    n12104, n12103, n12105, n12118, n12107, n12447, n16485, n12120, n16554,
    n12112, n12108, n12110, n12109, n12111, n16566, n12114, n12117, n12121,
    n12113, n12115, n16472, n12116, n16557, n16479, n16478, n16483, n16556,
    n16560, n16444, n12132, n12124, n12130, n12125, n12127, n12126, n12128,
    n16445, n12131, n12137, n12133, n12135, n12134, n12136, n12138, n12139,
    n12140, n16582, n12145, n12141, n12143, n12142, n12144, n12147, n13640,
    n12146, n12148, n13639, n12153, n12149, n12151, n12150, n12152, n12155,
    n13636, n12154, n12156, n13637, n12159, n12158, n12160, n12162, n13504,
    n12164, n12163, n12169, n12167, n12166, n12168, n12170, n12171, n12172,
    n13706, n12177, n12175, n12174, n12176, n12196, n13585, n12183, n12178,
    n12181, n12180, n12182, n12190, n13674, n12195, n12189, n12187, n12186,
    n12188, n13589, n13672, n12194, n12192, n12191, n12193, n12202, n12200,
    n13670, n12198, n12197, n13587, n12199, n12201, n12209, n12204, n12207,
    n12206, n12208, n12210, n13530, n12212, n12211, n13531, n12214, n13621,
    n12218, n12217, n12225, n13910, n12223, n12222, n12224, n12227, n12228,
    n12230, n12229, n13545, n12232, n12231, n12238, n13896, n12236, n12235,
    n12237, n12239, n12241, n12240, n13656, n12243, n12242, n12248, n13872,
    n12246, n12245, n12247, n12250, n12249, n13654, n12251, n12252, n12254,
    n12253, n13605, n13817, n12258, n12257, n12260, n12259, n12261, n12275,
    n12265, n12264, n13602, n12273, n12269, n12268, n12271, n12270, n12272,
    n17525, n12274, n12276, n12279, n12281, n12277, n12278, n12283, n12280,
    n12282, n12284, n12286, n12285, n12295, n12288, n12287, n12294, n13610,
    n13792, n12292, n12291, n12293, n13559, n12297, n12308, n12300, n13777,
    n12302, n12301, n12307, n12305, n12304, n12306, n13688, n12310, n12309,
    n13689, n12312, n12353, n13695, n12326, n13756, n12315, n12317, n12316,
    n12318, n12349, n12319, n12320, n12322, n12323, n12343, n12341, n12339,
    n12325, n12324, n12331, n13741, n12329, n12328, n12330, n12931, n12333,
    n12332, n12337, n12334, n12336, n12338, n12340, n12342, n12376, n12347,
    n12346, n12482, n12374, n12350, n12351, n12373, n12355, n12352, n12354,
    n12371, n12854, n12369, n12367, n12357, n12356, n12365, n12880, n12359,
    n12363, n12361, n12360, n12362, n12364, n12366, n12368, n12370, n12372,
    n12378, n12375, n12377, n12385, n12380, n12382, n12384, n12395, n12387,
    n12388, n16383, n12391, n12390, n12393, n16326, n12397, n12396, n12400,
    n12404, n12403, n12408, n12407, n12406, n13322, n13004, n12426, n12410,
    n12411, n12412, n12421, n12414, n12413, n12416, n12415, n16424, n12417,
    n14707, n12419, n12418, n12420, n13005, n13011, n12423, n12422, n12424,
    n12425, n12572, n12428, n12427, n12492, n12429, n12462, n12491, n14084,
    n14022, n12460, n14045, n12968, n14021, n12432, n12433, n12461, n12437,
    n17184, n12436, n12607, n17381, n17098, n17095, n12439, n17111, n17074,
    n12441, n12440, n12442, n17082, n17406, n12445, n17028, n17043, n12499,
    n17004, n12959, n12446, n12449, n12958, n17005, n12448, n12452, n16969,
    n17429, n14124, n12453, n12454, n16967, n12455, n12456, n12457, n12459,
    n12458, n14020, n12901, n12903, n13969, n12463, n13945, n13944, n13923,
    n13922, n12909, n13918, n12915, n13883, n13856, n12799, n12465, n12916,
    n13859, n12467, n12466, n12470, n13881, n12468, n12763, n13857, n12469,
    n13810, n12779, n12474, n12473, n13827, n13811, n12475, n12781, n12948,
    n12949, n13694, n12477, n13751, n12478, n12479, n12832, n13768, n12480,
    n12487, n12486, n12485, n12490, n12489, n12551, n12733, n12493, n12720,
    n14017, n12725, n13992, n12732, n13971, n17142, n12495, n17177, n12615,
    n12496, n12498, n12642, n12643, n17030, n12667, n14090, n16992, n12960,
    n16961, n12684, n14093, n12500, n12505, n12962, n12963, n12502, n12501,
    n14119, n12503, n12964, n12508, n12507, n14091, n14066, n14042, n12708,
    n14016, n13991, n12510, n12512, n13947, n13974, n12899, n12904, n12906,
    n12513, n12900, n12975, n13853, n12515, n12950, n12923, n12791, n13804,
    n12925, n12926, n13765, n12518, n12516, n12517, n12929, n12521, n13735,
    n12519, n12531, n12520, n12522, n12527, n13764, n12523, n13736, n12524,
    n12525, n12526, n12528, n12535, n12530, n12532, n12533, n12564, n12537,
    n12538, n12555, n17178, n12549, n14049, n12547, n12539, n12543, n12541,
    n12540, n12542, n17203, n12545, n13718, n12546, n12548, n12550, n12554,
    n12553, n13495, n12556, n13493, n13496, n12560, n12558, n12559, n12561,
    n12565, n17209, n12563, n12562, n12571, n17088, n17183, n13983, n12569,
    n17123, n12567, n13720, n12568, n12570, n12574, n12573, n13000, n17440,
    n12578, n12933, n12577, n12579, n12582, n12587, n12586, n12588, n17460,
    n17472, n12590, n12589, n12592, n12591, n12593, n12604, n12597, n12596,
    n12598, n12989, n12600, n12599, n12601, n12603, n12612, n12605, n12610,
    n12608, n12609, n12611, n12626, n12614, n12613, n12617, n12624, n12616,
    n12621, n12627, n12618, n12619, n12620, n12622, n12633, n12625, n12630,
    n12628, n12629, n12631, n12632, n12635, n12640, n12638, n12637, n12639,
    n12641, n17059, n12646, n12645, n12647, n12648, n12649, n12651, n12650,
    n12663, n12655, n12653, n12652, n12654, n12669, n12656, n12657, n12658,
    n12662, n12659, n12660, n12661, n12673, n12664, n12666, n12665, n12671,
    n12668, n12670, n12672, n12674, n12679, n17442, n12676, n12678, n12677,
    n12681, n12680, n12683, n12686, n12685, n12687, n12689, n12688, n12690,
    n12691, n12694, n12693, n12703, n12698, n12695, n12697, n12696, n12704,
    n12702, n12700, n12699, n12701, n12714, n12705, n12706, n12712, n12710,
    n12709, n12711, n12713, n12719, n12716, n12715, n12717, n12718, n12723,
    n12722, n12721, n12727, n12726, n12728, n12730, n12729, n12731, n12735,
    n12734, n12736, n12738, n12737, n12739, n12742, n12741, n12743, n12745,
    n12744, n12746, n12748, n12747, n12749, n12750, n12752, n12751, n12755,
    n12754, n12756, n12757, n12759, n12758, n12760, n12762, n12761, n12772,
    n12767, n12765, n12764, n12766, n12768, n12770, n12769, n12798, n12771,
    n12776, n12774, n12773, n12775, n12825, n12778, n12777, n12782, n12780,
    n12803, n12787, n12783, n12785, n12784, n12786, n12788, n12818, n12789,
    n12790, n12793, n12792, n12817, n12795, n12794, n12807, n12806, n12797,
    n12796, n12802, n12800, n12801, n12804, n12828, n12814, n12809, n12816,
    n12820, n12811, n12810, n12812, n12819, n12813, n12815, n12827, n12821,
    n12823, n12822, n12824, n12830, n12829, n12834, n12833, n12835, n12837,
    n12836, n12859, n12840, n12844, n12843, n12845, n12870, n12846, n12868,
    n12850, n12849, n14141, n12939, n12851, n12852, n12853, n12856, n12857,
    n12947, n12858, n12861, n12984, n12864, n12867, n12866, n12873, n12872,
    n12874, n12875, n12877, n12876, n12878, n12879, n12885, n12883, n12882,
    n12884, n12890, n12886, n12986, n12888, n12889, n12891, n12907, n12902,
    n12972, n12905, n12970, n12908, n12913, n12917, n12922, n12921, n12927,
    n12928, n12930, n12932, n12934, n12938, n12937, n12940, n12941, n12942,
    n12943, n12945, n12983, n12980, n13806, n13829, n12952, n12951, n12953,
    n17107, n12955, n12954, n12957, n12956, n17014, n14126, n16972, n12965,
    n14098, n12967, n12966, n14071, n14024, n12974, n12973, n12976, n12977,
    n12978, n12981, n13786, n12982, n12988, n12990, n12991, n12996, n12998,
    n13002, n17229, n13001, n13003, n13021, n13006, n13019, n13010, n13017,
    n15023, n13015, n13014, n13016, n13018, n13020, n13022, n13038, n13024,
    n13027, n13026, n13044, n13028, n13030, n13029, n13033, n13032, n13388,
    n13037, n13041, n15934, n13043, n13046, n13045, n13050, n13049, n13048,
    n13062, n13053, n13060, n13055, n13058, n13057, n13059, n13061, n13064,
    n13063, n13066, n13068, n13067, n13069, n13071, n13070, n13072, n13074,
    n13073, n13090, n13080, n13078, n13077, n13079, n13081, n13097, n13083,
    n13103, n13087, n13086, n13089, n13088, n13098, n13094, n13092, n13093,
    n13095, n13096, n13101, n13100, n13102, n13109, n13104, n13107, n13106,
    n13108, n13114, n13110, n13112, n13111, n13113, n13115, n13117, n13116,
    n13118, n13120, n13119, n13121, n13124, n13123, n13125, n13130, n13128,
    n13127, n13129, n13135, n13132, n13131, n13133, n13141, n13430, n13139,
    n13137, n13138, n13140, n13145, n13144, n13143, n13147, n13146, n13150,
    n13153, n13152, n13154, n13156, n13155, n13157, n13158, n13160, n13165,
    n13163, n13162, n13164, n13170, n13166, n13168, n13167, n13169, n13178,
    n13172, n13171, n13176, n13175, n13174, n13177, n13186, n13180, n13182,
    n13181, n13185, n13183, n13184, n13188, n13187, n13189, n13195, n13191,
    n13193, n13192, n13194, n13197, n13196, n13199, n13198, n13201, n13206,
    n13200, n13204, n13203, n13202, n13208, n13207, n13210, n13209, n13211,
    n13212, n13214, n13216, n13215, n13217, n13219, n13218, n13220, n13226,
    n13222, n13224, n13223, n13225, n13230, n13228, n13227, n13229, n13235,
    n13231, n13233, n13232, n13234, n13240, n13238, n13237, n13239, n13246,
    n13241, n13244, n13243, n13245, n13250, n13248, n13247, n13249, n13252,
    n13251, n13253, n13255, n13257, n15243, n13260, n13262, n13266, n13265,
    n13268, n13267, n16427, n13275, n13363, n13270, n13272, n13274, n13324,
    n13276, n13277, n14746, n14770, n14862, n13280, n13279, n13435, n13281,
    n15664, n13387, n16171, n13284, n15850, n13291, n15893, n13289, n13287,
    n13288, n13290, n13293, n13295, n13296, n13297, n13299, n15680, n13300,
    n13304, n13302, n13301, n13303, n13306, n13305, n15008, n13308, n13311,
    n14911, n13312, n14888, n14836, n13315, n13316, n13317, n13318, n13320,
    n13321, n13474, n13472, n13334, n13328, n13329, n13332, n13331, n13333,
    n13452, n13345, n13337, n13339, n13340, n13342, n13344, n13386, n13348,
    n13347, n13350, n13385, n13353, n13463, n13356, n13355, n13466, n13358,
    n13357, n13362, n13359, n13361, n13360, n13467, n13365, n13364, n13366,
    n13368, n13371, n13370, n13372, n13373, n16044, n13374, n13380, n13378,
    n13377, n13379, n13381, n16039, n13384, n13458, n13454, n13389, n13391,
    n13392, n13394, n13396, n13400, n13399, n13405, n13403, n13404, n13407,
    n13408, n13411, n13410, n13413, n13415, n13417, n13421, n13420, n13425,
    n13424, n13429, n13428, n13431, n13434, n13433, n13437, n13436, n13439,
    n13445, n13443, n13441, n13442, n13444, n13447, n13449, n13450, n13451,
    n13453, n13456, n13457, n13462, n13461, n13464, n13465, n13469, n13468,
    n13471, n13470, n13473, n13475, n13476, n13481, n13478, n13480, n13489,
    n13487, n13485, n13486, n13488, n13490, n13494, n13498, n13497, n13499,
    n17511, n17512, n13503, n13502, n13506, n13517, n13515, n13513, n13509,
    n13507, n16892, n13508, n13511, n13510, n13512, n13514, n13516, n13519,
    n13529, n13525, n13523, n13521, n13520, n13522, n13524, n13527, n13526,
    n13528, n13532, n13534, n13544, n13542, n13540, n13536, n13538, n13537,
    n13539, n13541, n13543, n13546, n13548, n13558, n14213, n13556, n13554,
    n13550, n13549, n13552, n13551, n13553, n13555, n13557, n13561, n13571,
    n13569, n13567, n13565, n13563, n13562, n13564, n13566, n13568, n13570,
    n13572, n13573, n13584, n13582, n13580, n13576, n16929, n13575, n13578,
    n13577, n13579, n13581, n13583, n13588, n13671, n13590, n13591, n13600,
    n13598, n13596, n13592, n16947, n13594, n13593, n13595, n13597, n13599,
    n13603, n13606, n13608, n13620, n13618, n13616, n16604, n13614, n13612,
    n13611, n13613, n13615, n13617, n13619, n13622, n13624, n13635, n13633,
    n13631, n13629, n13627, n13626, n13628, n13630, n13632, n13634, n13642,
    n16514, n16513, n16516, n13641, n13643, n13653, n13651, n13649, n13645,
    n16871, n13647, n13646, n13648, n13650, n13652, n13658, n13657, n13659,
    n13669, n14205, n13667, n13663, n13661, n13660, n13662, n13665, n13664,
    n13666, n13668, n13673, n13675, n13676, n13687, n13962, n13683, n13679,
    n13681, n13680, n13682, n13685, n14241, n13684, n13686, n13690, n13692,
    n13705, n13703, n13701, n13697, n13696, n13699, n13698, n13700, n13702,
    n13704, n13708, n13717, n13715, n13713, n13709, n16907, n13711, n13710,
    n13712, n13714, n13716, n13724, n13722, n13721, n13725, n13723, n13728,
    n13726, n13727, n13730, n13732, n13731, n14151, n13734, n13733, n13750,
    n13737, n13738, n17108, n17128, n13746, n14085, n13744, n13742, n13743,
    n13745, n13747, n13749, n13754, n14159, n13757, n13758, n13759, n13763,
    n13762, n14107, n13761, n13766, n13767, n14160, n13769, n13772, n13771,
    n14169, n13775, n13773, n13774, n13784, n13782, n13780, n13778, n13779,
    n13781, n13783, n13788, n14170, n13787, n13789, n13791, n13790, n14179,
    n13796, n13793, n13794, n13795, n13797, n13800, n13798, n13799, n13803,
    n13802, n13809, n13807, n14180, n13808, n13812, n13813, n13814, n13816,
    n13815, n14190, n13820, n13818, n13819, n13821, n13823, n13822, n13826,
    n13825, n13832, n13830, n14185, n13831, n14195, n13843, n13836, n13841,
    n13839, n13838, n13840, n13842, n14201, n13845, n13844, n13852, n13850,
    n13848, n13847, n13849, n13851, n14204, n13868, n13858, n13860, n13861,
    n13866, n13864, n13863, n13865, n13867, n14209, n13870, n13869, n13878,
    n13876, n13874, n13873, n13875, n13877, n14212, n13892, n13882, n13884,
    n13885, n13890, n13888, n13887, n13889, n13891, n14217, n13894, n13893,
    n13902, n13900, n13898, n13897, n13899, n13901, n13903, n13906, n13905,
    n14225, n13908, n13907, n13917, n13915, n13913, n13911, n13912, n13914,
    n13916, n13921, n14220, n13920, n13940, n13925, n13928, n13927, n14235,
    n13930, n13929, n13939, n13937, n13935, n13934, n13936, n13938, n13943,
    n14230, n13942, n13946, n13949, n14240, n13957, n13950, n13955, n13953,
    n13952, n13954, n13956, n14245, n13960, n13959, n13968, n13966, n13964,
    n13963, n13965, n13967, n14248, n13980, n13973, n13978, n13976, n13975,
    n13977, n13979, n14254, n13982, n13981, n13990, n13988, n13986, n13985,
    n13987, n13989, n13993, n13994, n14257, n14015, n13997, n13999, n14000,
    n14001, n14003, n14002, n14263, n14004, n14005, n14007, n14006, n14013,
    n14011, n14010, n14012, n14014, n14018, n14019, n14268, n14041, n14046,
    n14023, n14025, n14026, n14028, n14027, n14274, n14030, n14029, n14039,
    n14031, n14037, n14035, n14034, n14036, n14038, n14040, n14044, n14279,
    n14065, n14047, n14048, n14052, n14051, n14284, n14057, n14054, n14055,
    n14056, n14058, n14060, n14059, n14063, n14062, n14064, n14069, n14070,
    n14289, n14089, n14073, n14075, n14074, n14295, n14080, n14077, n14078,
    n14079, n14081, n14083, n14082, n14087, n14086, n14088, n14092, n14095,
    n14096, n17461, n14113, n14100, n14102, n14101, n17469, n14103, n14104,
    n14106, n14105, n14111, n14109, n14108, n14110, n14112, n14115, n14114,
    n14133, n14118, n14117, n14123, n14120, n14121, n17441, n14122, n14129,
    n16968, n14127, n14128, n17439, n14130, n14131, n14132, n14135, n14134,
    n14137, n17462, n14138, n14300, n14140, n14139, n14143, n14303, n14145,
    n14144, n14148, n14147, n14149, n14152, n14306, n14154, n14153, n14157,
    n14156, n14158, n14162, n14161, n14309, n14164, n14163, n14167, n14166,
    n14168, n14172, n14171, n14312, n14174, n14173, n14177, n14176, n14178,
    n14182, n14181, n14315, n14184, n14183, n14192, n14188, n14187, n14189,
    n14191, n14318, n14194, n14193, n14199, n14197, n14198, n14200, n14321,
    n14203, n14202, n14207, n14206, n14208, n14324, n14211, n14210, n14215,
    n14214, n14216, n14327, n14219, n14218, n14227, n14223, n14222, n14224,
    n14226, n14330, n14229, n14228, n14237, n14233, n14232, n14234, n14236,
    n14333, n14239, n14238, n14243, n14242, n14244, n14336, n14247, n14246,
    n14252, n14250, n14251, n14253, n14339, n14256, n14255, n14265, n14261,
    n14260, n14262, n14264, n14342, n14267, n14266, n14276, n14272, n14271,
    n14273, n14275, n14345, n14278, n14277, n14286, n14282, n14281, n14283,
    n14285, n14348, n14288, n14287, n14297, n14293, n14292, n14294, n14296,
    n14351, n14299, n14298, n14302, n14301, n14305, n14304, n14308, n14307,
    n14311, n14310, n14314, n14313, n14317, n14316, n14320, n14319, n14323,
    n14322, n14326, n14325, n14329, n14328, n14332, n14331, n14335, n14334,
    n14338, n14337, n14341, n14340, n14344, n14343, n14347, n14346, n14350,
    n14349, n14353, n14352, n14361, n14357, n14355, n14356, n14359, n14358,
    n14360, n14366, n14364, n14363, n14365, n14369, n14371, n14381, n14379,
    n14377, n14373, n15533, n14375, n14374, n14376, n14378, n14380, n14383,
    n14384, n14394, n14392, n14390, n14386, n14385, n14388, n14387, n14389,
    n14391, n14393, n14586, n14396, n14403, n14398, n14401, n14400, n14402,
    n14405, n14404, n14407, n14406, n14608, n14411, n14410, n14417, n14414,
    n14416, n14418, n14427, n14425, n14423, n14419, n14649, n14421, n14420,
    n14422, n14424, n14426, n14429, n14538, n14541, n14434, n14433, n14435,
    n14445, n14443, n14441, n14437, n14436, n14439, n14438, n14440, n14442,
    n14444, n14452, n14450, n14451, n14453, n14465, n14463, n14461, n14456,
    n15508, n14459, n14458, n14460, n14462, n14464, n14469, n14470, n14480,
    n14478, n14476, n14472, n14471, n14474, n14473, n14475, n14477, n14479,
    n14482, n14635, n14485, n14634, n14488, n14487, n14502, n14490, n14489,
    n14491, n14500, n14498, n14496, n14492, n15562, n14494, n14493, n14495,
    n14497, n14499, n14506, n14505, n14507, n14516, n14512, n14508, n15577,
    n14510, n14509, n14511, n14514, n14513, n14515, n14519, n14522, n14521,
    n14526, n14525, n14527, n14537, n14535, n14533, n14529, n14528, n14531,
    n14530, n14532, n14534, n14536, n14540, n14542, n14552, n14550, n14548,
    n14544, n14543, n14546, n14545, n14547, n14549, n14551, n14555, n14557,
    n14569, n14567, n14565, n14561, n15519, n14560, n14563, n14562, n14564,
    n14566, n14568, n14573, n14574, n14584, n14582, n14580, n14576, n14575,
    n14578, n14577, n14579, n14581, n14583, n14589, n14588, n14594, n14593,
    n14592, n14596, n14595, n14602, n15491, n14599, n14598, n14600, n14601,
    n14604, n14603, n14606, n14605, n14609, n14619, n14617, n14615, n14611,
    n15588, n14613, n14612, n14614, n14616, n14618, n14631, n14629, n14624,
    n14623, n14627, n14626, n14628, n14630, n14632, n14637, n14638, n14647,
    n14645, n14643, n14639, n15547, n14641, n14640, n14642, n14644, n14646,
    n14648, n14675, n14672, n15603, n14670, n15590, n14668, n14666, n14661,
    n15535, n14659, n14657, n15510, n14655, n15496, n14653, n14652, n15495,
    n14654, n15509, n14656, n15524, n15523, n14658, n15534, n14660, n14662,
    n14664, n15550, n14663, n15559, n15558, n14665, n15578, n15579, n14667,
    n15589, n14669, n14671, n14673, n14674, n14700, n15594, n14694, n14692,
    n15564, n14687, n15538, n14685, n14683, n14681, n15493, n14678, n15492,
    n14680, n15505, n15504, n14682, n15520, n15521, n14684, n15537, n14686,
    n14688, n14690, n15548, n14689, n15563, n14691, n15573, n15572, n14693,
    n15593, n15597, n14695, n14697, n14696, n14698, n14699, n14702, n14701,
    n14713, n14711, n14709, n14708, n15044, n14714, n14710, n14712, n15042,
    n14719, n14717, n14715, n14716, n14718, n15747, n14729, n15051, n14727,
    n14725, n14723, n14724, n14726, n14728, n14740, n14732, n14736, n14734,
    n14733, n14735, n14738, n14737, n14739, n15059, n14766, n14745, n14747,
    n14748, n14752, n14750, n14749, n14751, n15065, n14754, n14753, n14764,
    n15060, n14762, n14760, n14758, n14759, n14761, n14763, n14765, n15070,
    n14788, n14769, n14771, n14772, n14777, n14775, n14774, n14776, n15075,
    n14780, n16289, n15073, n14785, n14783, n14782, n14784, n14786, n14787,
    n14789, n14791, n14790, n15080, n14812, n14794, n14798, n14796, n14795,
    n14797, n15086, n14800, n14799, n14810, n15081, n14808, n14806, n14804,
    n14805, n14807, n14809, n14811, n15091, n14831, n14816, n14821, n14819,
    n14818, n14820, n15096, n14823, n15094, n14828, n14826, n14825, n14827,
    n14829, n14830, n14832, n14834, n14833, n15101, n14845, n14838, n14843,
    n14841, n14840, n14842, n14844, n15108, n14847, n14846, n14859, n15675,
    n15954, n14857, n14849, n14850, n15104, n14986, n14855, n14853, n14852,
    n14854, n14856, n14858, n15111, n14872, n14864, n14870, n14868, n14867,
    n14869, n14871, n15119, n14874, n14873, n14886, n14884, n15112, n14882,
    n14880, n14878, n14879, n14881, n14883, n14885, n15122, n14907, n14890,
    n14895, n14893, n14892, n14894, n15128, n14897, n14896, n14905, n15123,
    n14903, n14901, n14899, n14900, n14902, n14904, n14906, n15133, n14934,
    n14910, n14913, n14912, n14914, n14918, n14916, n14915, n14917, n15139,
    n14920, n14919, n14932, n14922, n15134, n14930, n14928, n14926, n14927,
    n14929, n14931, n14933, n14948, n15144, n14945, n15145, n14943, n14941,
    n14940, n14942, n14944, n14959, n14949, n14950, n14955, n14953, n14952,
    n14954, n15150, n14957, n14956, n14958, n14969, n15155, n14968, n15156,
    n14966, n14964, n14963, n14965, n14967, n14980, n14971, n14976, n14974,
    n14973, n14975, n15161, n14978, n14977, n14979, n15166, n14993, n14983,
    n14985, n15169, n14991, n14989, n14988, n14990, n14992, n15006, n14996,
    n15002, n15000, n14999, n15001, n15171, n15004, n15003, n15005, n15176,
    n15018, n15010, n15016, n15014, n15013, n15015, n15017, n15184, n15021,
    n15019, n15020, n15034, n15032, n15177, n15030, n15028, n15026, n15027,
    n15029, n15031, n15033, n15039, n16291, n15037, n15038, n15187, n15041,
    n15040, n15047, n15045, n15046, n15190, n15049, n15048, n16318, n15054,
    n15053, n15055, n15058, n15057, n15067, n15063, n15062, n15064, n15066,
    n15196, n15069, n15068, n15077, n15072, n15074, n15199, n15079, n15078,
    n15088, n15084, n15083, n15085, n15087, n15202, n15090, n15089, n15098,
    n15093, n15095, n15097, n15205, n15100, n15099, n15106, n15103, n15105,
    n15107, n15208, n15110, n15109, n15117, n15115, n15114, n15116, n15118,
    n15211, n15121, n15120, n15130, n15126, n15125, n15127, n15129, n15214,
    n15132, n15131, n15141, n15137, n15136, n15138, n15140, n15217, n15143,
    n15142, n15152, n15148, n15147, n15149, n15151, n15220, n15154, n15153,
    n15163, n15159, n15158, n15160, n15162, n15223, n15165, n15164, n15173,
    n15168, n15170, n15172, n15226, n15175, n15174, n15182, n15180, n15179,
    n15181, n15183, n15229, n15186, n15185, n15189, n15188, n15192, n15191,
    n15194, n15198, n15197, n15201, n15200, n15204, n15203, n15207, n15206,
    n15210, n15209, n15213, n15212, n15216, n15215, n15219, n15218, n15222,
    n15221, n15225, n15224, n15228, n15227, n15231, n15230, n15240, n15234,
    n15235, n15238, n16159, n15237, n15239, n15242, n15247, n15245, n15244,
    n15246, n15249, n15248, n15257, n15252, n15253, n15255, n15256, n15263,
    n15261, n15259, n15260, n15262, n15265, n15264, n15271, n15267, n15269,
    n15270, n15277, n15273, n15275, n15274, n15276, n15279, n15283, n15281,
    n15280, n15282, n15291, n15323, n15287, n15289, n15288, n15290, n15292,
    n15464, n15302, n15367, n15294, n15300, n15298, n15901, n15296, n15295,
    n15297, n15299, n15301, n15304, n15303, n15317, n15305, n15444, n15315,
    n15309, n15310, n15313, n15312, n15314, n15316, n15321, n15341, n15326,
    n15325, n15330, n15329, n15331, n15337, n15335, n15334, n15336, n15339,
    n15338, n15340, n15343, n15342, n15354, n15349, n15348, n15350, n15352,
    n15351, n15353, n15357, n15356, n15359, n15476, n15365, n15363, n15362,
    n15364, n15385, n15371, n15370, n15375, n15374, n15379, n15377, n15378,
    n15383, n15826, n15382, n15384, n15388, n15387, n15389, n15390, n15391,
    n15394, n15393, n15396, n15395, n15398, n15397, n15405, n15401, n15403,
    n15402, n15404, n15413, n15410, n15409, n15411, n15412, n15415, n15414,
    n15422, n15420, n15418, n15419, n15421, n15442, n15424, n15425, n15429,
    n15427, n15428, n15430, n15436, n15433, n15435, n15456, n15439, n15440,
    n15441, n15443, n15451, n15449, n15447, n15448, n15450, n15458, n15454,
    n15455, n15457, n15461, n15469, n15463, n15462, n15465, n15467, n15466,
    n15468, n15474, n15472, n15473, n15475, n15484, n15482, n15480, n15481,
    n15483, n15489, n15487, n15488, n15490, n15503, n15494, n15501, n15497,
    n15499, n15498, n15500, n15502, n15506, n15517, n15507, n15515, n15513,
    n15511, n15512, n15514, n15516, n15518, n15531, n15522, n15529, n15525,
    n15527, n15526, n15528, n15530, n15532, n15543, n15536, n15541, n15539,
    n15540, n15542, n15545, n15544, n15546, n15557, n15549, n15555, n15551,
    n15553, n15552, n15554, n15556, n15560, n15571, n15561, n15569, n15565,
    n15567, n15566, n15568, n15570, n15575, n15586, n15576, n15584, n15580,
    n15582, n15581, n15583, n15585, n15587, n15602, n15592, n15600, n15595,
    n15598, n15599, n15601, n15606, n15605, n15609, n15608, n15612, n15611,
    n15631, n16328, n15626, n15627, n16335, n15942, n15624, n15617, n15622,
    n15620, n15619, n15621, n15623, n16333, n15625, n15629, n15628, n15630,
    n15633, n15632, n15636, n15635, n15653, n16314, n15651, n16319, n15649,
    n15642, n15641, n15647, n15645, n15646, n16323, n15648, n15650, n15652,
    n15655, n15654, n15658, n15657, n15673, n16303, n15671, n16307, n15669,
    n15663, n15662, n15667, n15665, n15666, n16311, n15668, n15670, n15672,
    n16296, n15676, n15690, n15679, n15681, n15687, n15683, n15682, n15685,
    n15684, n15686, n16298, n15688, n15689, n15693, n15692, n15694, n15700,
    n15696, n16290, n15698, n15699, n15702, n15701, n15704, n15703, n15707,
    n15706, n15721, n16278, n15719, n16282, n15717, n15715, n15713, n15712,
    n15714, n16286, n15716, n15718, n15720, n15724, n15791, n15764, n15726,
    n15727, n15728, n15731, n15730, n16270, n15733, n15736, n15735, n16273,
    n15739, n15738, n15740, n15743, n15742, n15744, n15749, n16268, n15748,
    n15751, n15750, n15753, n15752, n15756, n15755, n15779, n16257, n15762,
    n15766, n16261, n15768, n15971, n15761, n15777, n15765, n15767, n15770,
    n15769, n15775, n15773, n15772, n15774, n16265, n15776, n15778, n15784,
    n15782, n15783, n15812, n15787, n15789, n16252, n15806, n15800, n15792,
    n15798, n15796, n16248, n15797, n15799, n15803, n15802, n16254, n15804,
    n15805, n15807, n15810, n15808, n15809, n15811, n15849, n15815, n15833,
    n15817, n15816, n15822, n15820, n15821, n16245, n16237, n15824, n15832,
    n15828, n15827, n15830, n15829, n15831, n15835, n16241, n15834, n15837,
    n16238, n15836, n15838, n15839, n16231, n15841, n15840, n15856, n15843,
    n15848, n15846, n15845, n15847, n16233, n15852, n15851, n16226, n15854,
    n15855, n15857, n15861, n15859, n15860, n15863, n15862, n15864, n15868,
    n15866, n15867, n15870, n15869, n15900, n15873, n15874, n15881, n15879,
    n15877, n15878, n15880, n16220, n15883, n15886, n15885, n16221, n15887,
    n15888, n15898, n15891, n15895, n15894, n16215, n15897, n15899, n16204,
    n15903, n15915, n15938, n15905, n15906, n15914, n15941, n15909, n16208,
    n15910, n15912, n15911, n15913, n16212, n15916, n15921, n15919, n15918,
    n15920, n15923, n15922, n15926, n16205, n15925, n15929, n15928, n15951,
    n15932, n16197, n15949, n15946, n15936, n15937, n15939, n15944, n15940,
    n15953, n16192, n15943, n15945, n15948, n15947, n16199, n15950, n15952,
    n15956, n15955, n15958, n15957, n15960, n16181, n15959, n15965, n15963,
    n15962, n15964, n15973, n15967, n15970, n16187, n15972, n15990, n15976,
    n15978, n15988, n15982, n15981, n15986, n15984, n15985, n15987, n16186,
    n15989, n15994, n15997, n15996, n16006, n15999, n16176, n16002, n16001,
    n16003, n16005, n16012, n16010, n16011, n16014, n16013, n16018, n16016,
    n16017, n16020, n16019, n17224, n16025, n16024, n16027, n17231, n16031,
    n16030, n16033, n16032, n16036, n16035, n16038, n16037, n16041, n16040,
    n16043, n16042, n16046, n16045, n16048, n16047, n16051, n16050, n16053,
    n16052, n16055, n16059, n16057, n16058, n16061, n16060, n16065, n16063,
    n16064, n16067, n16066, n17265, n16072, n16070, n16071, n16074, n16073,
    n16078, n16076, n16077, n16080, n16079, n16084, n16082, n16083, n16086,
    n16085, n17282, n16091, n16089, n16090, n16093, n16092, n17288, n16098,
    n16096, n16097, n16100, n16099, n16104, n16102, n16103, n16106, n16105,
    n16109, n16108, n16111, n16110, n16114, n16113, n16116, n16115, n16119,
    n16118, n16121, n16120, n16124, n16123, n16126, n16125, n17324, n16131,
    n16129, n16130, n16133, n16132, n16138, n16137, n16140, n16139, n16145,
    n16143, n16144, n16147, n16146, n16151, n16149, n16150, n16153, n16152,
    n16158, n16156, n16157, n16161, n16160, n16164, n16167, n16163, n16169,
    n16168, n16180, n16172, n16178, n16175, n16177, n16341, n16179, n16191,
    n16184, n16183, n16185, n16189, n16334, n16188, n16344, n16190, n16201,
    n16195, n16194, n16196, n16198, n16347, n16200, n16214, n16203, n16207,
    n16206, n16210, n16209, n16211, n16350, n16213, n16224, n16218, n16217,
    n16219, n16222, n16353, n16223, n16235, n16229, n16228, n16230, n16232,
    n16356, n16234, n16247, n16236, n16240, n16239, n16243, n16242, n16244,
    n16359, n16246, n16256, n16250, n16249, n16251, n16253, n16362, n16255,
    n16267, n16260, n16259, n16263, n16262, n16264, n16365, n16266, n16277,
    n16269, n16275, n16272, n16274, n16368, n16276, n16288, n16281, n16280,
    n16284, n16283, n16285, n16371, n16287, n16302, n16294, n16293, n16300,
    n16297, n16299, n16374, n16301, n16313, n16306, n16305, n16309, n16308,
    n16310, n16377, n16312, n16325, n16317, n16316, n16321, n16320, n16322,
    n16380, n16324, n16340, n16331, n16330, n16332, n16337, n16336, n16384,
    n16339, n16343, n16342, n16346, n16345, n16349, n16348, n16352, n16351,
    n16355, n16354, n16358, n16357, n16361, n16360, n16364, n16363, n16367,
    n16366, n16370, n16369, n16373, n16372, n16376, n16375, n16379, n16378,
    n16382, n16381, n16387, n16386, n16390, n16389, n16393, n16392, n16396,
    n16395, n16399, n16398, n16402, n16401, n16405, n16404, n16408, n16407,
    n16411, n16410, n16414, n16413, n16417, n16416, n16420, n16419, n16423,
    n16422, n16426, n16425, n16429, n16428, n16430, n16753, n16434, n16432,
    n16431, n16433, n16439, n16435, n16437, n16436, n16438, n16441, n16440,
    n16455, n16443, n16808, n16453, n16447, n16446, n16448, n16451, n16450,
    n16452, n16454, n16457, n16456, n16465, n16463, n16461, n16462, n16464,
    n16471, n16467, n16678, n16469, n16468, n16470, n16475, n16474, n16494,
    n17018, n16476, n16770, n16492, n16484, n16481, n16480, n16482, n16488,
    n16486, n16487, n16490, n16489, n16491, n16493, n16497, n16505, n16499,
    n16498, n16503, n16501, n16500, n16502, n16504, n16506, n16852, n16509,
    n16508, n16521, n16512, n16511, n16519, n16515, n16517, n16518, n16520,
    n16523, n16720, n16527, n16525, n16524, n16526, n16536, n16529, n16530,
    n16532, n16534, n16533, n16535, n16537, n16702, n16549, n16540, n16547,
    n16541, n16545, n16544, n16546, n16548, n16551, n16550, n16553, n16552,
    n16565, n16561, n16558, n16559, n16563, n16562, n16564, n16571, n16567,
    n16795, n16569, n16568, n16570, n16572, n16834, n16576, n16575, n16589,
    n16579, n16578, n16587, n16585, n16583, n16584, n16586, n16588, n16592,
    n16591, n16600, n16596, n16598, n16597, n16599, n16603, n16602, n16607,
    n16606, n16615, n16611, n16613, n16614, n16622, n16617, n16732, n16620,
    n16619, n16621, n16624, n16623, n16627, n16626, n16633, n16631, n16630,
    n16632, n16637, n16635, n16636, n16654, n16640, n16642, n16641, n16652,
    n16650, n16647, n16646, n16648, n16649, n16651, n16653, n16656, n16655,
    n16673, n16659, n16661, n16671, n16664, n16669, n16667, n16668, n16670,
    n16672, n16675, n16674, n16677, n16679, n16690, n16682, n16688, n16686,
    n16684, n16685, n16687, n16689, n16692, n16691, n16695, n16700, n16698,
    n16699, n16712, n16703, n16710, n16708, n16706, n16707, n16709, n16711,
    n16715, n16717, n16716, n16730, n16719, n16721, n16728, n16726, n16724,
    n16725, n16727, n16729, n16733, n16748, n16736, n16746, n16739, n16744,
    n16742, n16743, n16745, n16747, n16750, n16749, n16752, n16754, n16765,
    n16757, n16763, n16759, n16761, n16760, n16762, n16764, n16767, n16766,
    n16769, n16784, n16773, n16782, n16776, n16780, n16778, n16779, n16781,
    n16783, n16786, n16785, n16788, n16803, n16790, n16801, n16793, n16799,
    n16794, n16797, n16796, n16798, n16800, n16802, n16806, n16812, n16807,
    n16810, n16809, n16811, n16820, n16815, n16818, n16819, n16825, n16823,
    n16824, n16827, n16842, n16829, n16840, n16832, n16838, n16833, n16836,
    n16835, n16837, n16839, n16841, n16845, n16860, n16847, n16858, n16850,
    n16856, n16851, n16854, n16853, n16855, n16857, n16859, n16863, n16879,
    n16866, n16877, n16869, n16875, n16870, n16873, n16872, n16874, n16876,
    n16878, n16882, n16898, n16884, n16896, n16887, n16894, n16890, n16889,
    n16891, n16893, n16895, n16897, n16900, n16915, n16902, n16913, n16905,
    n16911, n16906, n16909, n16908, n16910, n16912, n16914, n16918, n16935,
    n16920, n16933, n16923, n16931, n16927, n16926, n16928, n16930, n16932,
    n16934, n16938, n16957, n16955, n16944, n16953, n16946, n16951, n16950,
    n16952, n16954, n16956, n16960, n16959, n16966, n16963, n16964, n17450,
    n16965, n16982, n16970, n16971, n16973, n16978, n16976, n16975, n16977,
    n17457, n16979, n16980, n16981, n16986, n16985, n17003, n16988, n16997,
    n16991, n16990, n16995, n17432, n16994, n16996, n17431, n16998, n16999,
    n17001, n17000, n17002, n17006, n17007, n17008, n17013, n17011, n17010,
    n17012, n17426, n17421, n17016, n17017, n17026, n17021, n17020, n17024,
    n17023, n17025, n17413, n17033, n17041, n17031, n17032, n17035, n17034,
    n17040, n17038, n17037, n17039, n17418, n17042, n17050, n17045, n17044,
    n17048, n17047, n17049, n17052, n17057, n17055, n17054, n17056, n17410,
    n17405, n17060, n17061, n17069, n17064, n17063, n17067, n17066, n17068,
    n17073, n17072, n17094, n17076, n17077, n17087, n17080, n17079, n17085,
    n17399, n17084, n17086, n17398, n17089, n17090, n17092, n17091, n17093,
    n17130, n17099, n17100, n17101, n17106, n17104, n17103, n17105, n17393,
    n17109, n17110, n17119, n17114, n17113, n17117, n17116, n17118, n17122,
    n17121, n17125, n17124, n17140, n17380, n17138, n17131, n17136, n17134,
    n17133, n17135, n17385, n17137, n17139, n17144, n17372, n17157, n17146,
    n17145, n17149, n17148, n17162, n17153, n17152, n17161, n17156, n17159,
    n17158, n17160, n17377, n17163, n17165, n17164, n17170, n17169, n17182,
    n17173, n17180, n17176, n17363, n17179, n17181, n17369, n17189, n17187,
    n17186, n17188, n17190, n17192, n17191, n17194, n17193, n17199, n17198,
    n17202, n17201, n17212, n17355, n17208, n17206, n17207, n17210, n17211,
    n17216, n17215, n17218, n17217, n17221, n17220, n17223, n17222, n17228,
    n17225, n17227, n17230, n17234, n17233, n17236, n17235, n17240, n17239,
    n17242, n17241, n17245, n17244, n17247, n17246, n17250, n17249, n17252,
    n17251, n17256, n17255, n17258, n17257, n17262, n17261, n17264, n17263,
    n17268, n17267, n17270, n17269, n17273, n17272, n17275, n17274, n17279,
    n17278, n17281, n17280, n17285, n17284, n17287, n17286, n17291, n17290,
    n17293, n17292, n17297, n17296, n17299, n17298, n17303, n17302, n17305,
    n17304, n17309, n17308, n17311, n17310, n17315, n17314, n17317, n17316,
    n17321, n17320, n17323, n17322, n17327, n17326, n17329, n17328, n17332,
    n17331, n17334, n17333, n17337, n17336, n17340, n17339, n17345, n17344,
    n17347, n17346, n17352, n17351, n17362, n17354, n17360, n17357, n17359,
    n17475, n17361, n17371, n17364, n17367, n17366, n17368, n17478, n17370,
    n17379, n17375, n17374, n17376, n17481, n17378, n17387, n17383, n17382,
    n17384, n17484, n17386, n17395, n17391, n17390, n17392, n17487, n17394,
    n17404, n17397, n17402, n17400, n17433, n17401, n17490, n17403, n17412,
    n17408, n17407, n17409, n17493, n17411, n17420, n17416, n17415, n17417,
    n17496, n17419, n17428, n17424, n17423, n17425, n17499, n17427, n17438,
    n17430, n17436, n17434, n17435, n17502, n17437, n17448, n17446, n17444,
    n17443, n17445, n17505, n17447, n17459, n17455, n17453, n17454, n17456,
    n17508, n17458, n17474, n17471, n17467, n17466, n17468, n17470, n17513,
    n17473, n17477, n17476, n17480, n17479, n17483, n17482, n17486, n17485,
    n17489, n17488, n17492, n17491, n17495, n17494, n17498, n17497, n17501,
    n17500, n17504, n17503, n17507, n17506, n17510, n17509, n17515, n17514,
    n17518, n17517, n17521, n17520, n17524, n17523, n17528, n17527, n17531,
    n17530, n17534, n17533, n17537, n17536, n17540, n17539, n17543, n17542,
    n17546, n17545, n17549, n17548, n17553, n17552, n17556, n17576, n17579,
    n17583, n17587, n17591, n17595, n17599, n17603, n17607, n13271, n9976,
    n11273, n13056, n13065, n17237;
  assign n11337 = ~n13383 | ~n11297;
  assign n11099 = n9635 & n9358;
  assign n14839 = ~n16403;
  assign n10624 = n17237 | n8880;
  assign n10370 = n12157 | n8880;
  assign n15659 = ~n16304;
  assign n17009 = n11577 | n11576;
  assign n15734 = n10275 | n10274;
  assign n13122 = n13085;
  assign n11905 = ~n9983 | ~n8917;
  assign n11910 = ~n9802 | ~n9913;
  assign n10007 = n9906 & n11873;
  assign n9875 = ~n9873 | ~P1_IR_REG_31__SCAN_IN;
  assign n10438 = n9525;
  assign n8909 = n13369 & n13472;
  assign n10803 = ~n10861;
  assign n12871 = ~n9525;
  assign n13336 = ~n15092 | ~n14839;
  assign n10121 = ~n10050 | ~n10049;
  assign n12266 = ~n12348;
  assign n12623 = ~n16466 | ~n16543;
  assign n10861 = ~n9867 | ~n11296;
  assign n8876 = n10864;
  assign n8891 = n10596;
  assign n14961 = ~n15157;
  assign n16271 = n10173 & n10172;
  assign n10119 = ~n10121 ^ SI_6_;
  assign n12865 = ~n12892;
  assign n13837 = ~n17529;
  assign n15167 = ~n10451 | ~n10450;
  assign n9833 = ~n9832 | ~P1_IR_REG_31__SCAN_IN;
  assign n15615 = ~n13427 | ~n13136;
  assign n16315 = ~n15637;
  assign n11282 = ~n11172;
  assign n12580 = ~n12551 & ~n12550;
  assign n14362 = ~n11405 ^ P2_IR_REG_30__SCAN_IN;
  assign n12072 = ~n11047 ^ n11046;
  assign n11906 = ~n9957 | ~n9956;
  assign n16202 = n9234 & n9235;
  assign n11800 = ~n10438;
  assign n16279 = ~n9282 | ~n10267;
  assign n11071 = ~P2_IR_REG_31__SCAN_IN;
  assign n16936 = ~n11149 ^ n12185;
  assign n9368 = ~n9890 | ~n9889;
  assign n9663 = ~n9826 & ~n9825;
  assign n9555 = ~n11997;
  assign n11997 = n10370 & n10369;
  assign n11149 = ~n9105 | ~n11148;
  assign n10996 = ~P2_IR_REG_12__SCAN_IN & ~P2_IR_REG_17__SCAN_IN;
  assign n9116 = n9117 | n16826;
  assign n8873 = ~n9920 | ~n13271;
  assign n10995 = ~P2_IR_REG_11__SCAN_IN & ~P2_IR_REG_13__SCAN_IN;
  assign n10864 = ~n10500;
  assign n8877 = ~n10128;
  assign n8878 = ~n8877;
  assign n8880 = ~n8877;
  assign n16028 = ~n9285 ^ n10680;
  assign n12290 = n11486;
  assign n16901 = ~n11099 ^ n12165;
  assign n10361 = ~n10422 | ~n10419;
  assign n10422 = ~n10326 | ~n10325;
  assign n8881 = n11959 & n16029;
  assign n13256 = ~n13085;
  assign n8896 = ~n13122;
  assign n9906 = ~n9898 ^ n15233;
  assign n9898 = n9899 | n9897;
  assign n8882 = ~n12847;
  assign n12847 = ~n12179 | ~n13271;
  assign n13278 = ~n15167 | ~n15011;
  assign n8884 = n11172;
  assign n8885 = ~n9867 | ~n11296;
  assign n10387 = ~n9386 | ~n10420;
  assign n8886 = ~n9894;
  assign n8887 = ~n9894;
  assign n10286 = ~n9894;
  assign n9444 = n9445 & n12912;
  assign n9635 = n16861 | n9636;
  assign n9668 = n9669 & n13330;
  assign n9763 = ~n10401 | ~n10400;
  assign n16612 = ~n9152 | ~n9149;
  assign n16543 = n11548 & n11547;
  assign n9110 = n9111 & n16697;
  assign n16666 = n11030 & n11040;
  assign n9103 = ~n9624 & ~n8965;
  assign n16634 = n11120 & n11121;
  assign P1_U3086 = ~P1_STATE_REG_SCAN_IN;
  assign n9605 = n12894 & n12575;
  assign n9260 = ~n13250 | ~n13249;
  assign n9400 = n15050 | n16318;
  assign n14620 = n14468 & n10780;
  assign n15050 = n9227 & n9226;
  assign n9335 = n11153 & n8903;
  assign n9136 = ~n8906 & ~n8951;
  assign n9589 = ~n9590 & ~n9027;
  assign n11899 = ~n11113 & ~n11112;
  assign n9591 = n11896 | n9034;
  assign n9590 = n11896 & n9594;
  assign n14539 = ~n8955 & ~n9693;
  assign n12529 = n13785 | n12517;
  assign n13785 = ~n9127 | ~n9430;
  assign n9294 = n14863 | n9666;
  assign n9126 = ~n13854 | ~n13853;
  assign n11998 = n14755 | n9558;
  assign n9487 = n11288 | n16817;
  assign n13854 = ~n9443 | ~n9444;
  assign n14484 = n10386 & n14368;
  assign n14704 = ~n13012;
  assign n9443 = ~n13919 | ~n9447;
  assign n16899 = ~n11145 ^ n12165;
  assign n9346 = ~n13312 & ~n9347;
  assign n9445 = ~n9447 | ~n9448;
  assign n16861 = ~n11091 ^ n11238;
  assign n12345 = ~n11868 ^ n11866;
  assign n9130 = n9133 & n16880;
  assign n14155 = ~n12313 | ~n12312;
  assign n14756 = n10792 & n10791;
  assign n14165 = ~n12298 | ~n12297;
  assign n11091 = ~n9269 | ~n9268;
  assign n13327 = n15113 | n14891;
  assign n9704 = n9705 & n14448;
  assign n14778 = n10761 & n10760;
  assign n12911 = ~n13625 | ~n17516;
  assign n14802 = n10702 & n10701;
  assign n9271 = n16828 | n11221;
  assign n14876 = n10624 & n10623;
  assign n14822 = n10722 & n10721;
  assign n15124 = ~n9767 | ~n10595;
  assign n15102 = ~n10663 | ~n10662;
  assign n13895 = ~n12230 | ~n12229;
  assign n10315 = n10314 & n14446;
  assign n13134 = ~n15615 & ~n13133;
  assign n9767 = n12213 | n8880;
  assign n9689 = ~n15369 | ~n10097;
  assign n13307 = ~n9763 | ~n14997;
  assign n15024 = ~n9763;
  assign n15613 = ~n15638 & ~n16315;
  assign n10752 = ~n9050 | ~n9047;
  assign n14269 = ~n12169 | ~n12168;
  assign n16826 = ~n11139 ^ n11225;
  assign n11077 = ~n9263 | ~n9265;
  assign n15638 = ~n9561 | ~n9564;
  assign n8904 = n9796 & n8996;
  assign n16054 = ~n9315 | ~n10480;
  assign n16068 = ~n9281 ^ n10392;
  assign n12430 = ~n12161 | ~n12160;
  assign n16805 = ~n9139 | ~n11137;
  assign n15818 = ~n9232 | ~n8992;
  assign n15637 = n10337 & n10336;
  assign n9546 = ~n10552 | ~n10522;
  assign n15709 = n13414 & n15677;
  assign n14290 = ~n12153 | ~n12152;
  assign n10552 = ~n9122 | ~n9119;
  assign n10337 = n17276 | n8880;
  assign n17451 = ~n12137 | ~n12136;
  assign n16442 = ~n12129 | ~n12128;
  assign n9282 = ~n9283 | ~n10720;
  assign n15344 = n9970 | n9969;
  assign n16774 = ~n9106 | ~n11134;
  assign n16258 = ~n10199 | ~n10198;
  assign n15819 = ~n15722 | ~n15723;
  assign n12348 = ~n9142 | ~n12896;
  assign n17200 = n12565 & n17120;
  assign n13286 = ~n13395 | ~n13397;
  assign n13395 = n16202 | n11905;
  assign n15785 = n10136 & n10135;
  assign n15722 = n13065 | n15844;
  assign n15823 = ~n11964;
  assign n13401 = n15882 | n11903;
  assign n13398 = ~n11903 | ~n15882;
  assign n13047 = n13056 | n15876;
  assign n13846 = ~P2_REG3_REG_23__SCAN_IN ^ n12267;
  assign n15729 = n10206 | n10207;
  assign n17102 = n11435 | n11434;
  assign n15844 = n10060 | n10059;
  assign n11964 = n10117 & n10116;
  assign n15876 = n10088 | n10089;
  assign n17175 = ~n12595 | ~n12594;
  assign n11903 = ~n9306 | ~n10008;
  assign n16507 = n11418 & n11417;
  assign n11055 = ~n11053 | ~n12077;
  assign n9467 = n16704 | n9468;
  assign n17036 = n11520 | n11519;
  assign n9802 = n9909 & n9908;
  assign n16216 = ~n10006 | ~n10005;
  assign n16466 = ~n9645 | ~n9079;
  assign n12644 = n11567 & n11566;
  assign n17151 = ~n8920 | ~n9099;
  assign n9913 = n9912 & n9911;
  assign n17053 = n11509 | n11508;
  assign n11128 = ~n9109 | ~n11127;
  assign n13263 = n10007;
  assign n9862 = n13009 | n13484;
  assign n15930 = n11909 & n11908;
  assign P2_U3893 = n11289 & P2_STATE_REG_SCAN_IN;
  assign n9234 = n9236 & n9977;
  assign n16173 = ~n9924 | ~n9923;
  assign n9520 = ~n10048 | ~n10047;
  assign n9109 = ~n9112 | ~n9110;
  assign n11531 = n11414 & n11878;
  assign n12881 = n11414 & n11413;
  assign n12848 = ~n12205;
  assign n9907 = ~n11873;
  assign n11990 = ~n11991 & ~n15426;
  assign n12205 = ~n12179 | ~n11800;
  assign n8889 = n12219;
  assign n8890 = ~n9800;
  assign n11486 = n14362 & n11413;
  assign n17319 = ~n11064 | ~n11068;
  assign n16029 = ~n10906 ^ n10905;
  assign n9920 = ~n15386 | ~n10935;
  assign n11878 = ~n11407 ^ P2_IR_REG_29__SCAN_IN;
  assign n9914 = n13376 & n13382;
  assign n10557 = ~n9831 | ~P1_IR_REG_31__SCAN_IN;
  assign n10906 = ~n9861 | ~P1_IR_REG_31__SCAN_IN;
  assign n11172 = ~n11403 | ~n11018;
  assign n10261 = ~n10230 ^ SI_10_;
  assign n12051 = ~n11014 ^ P2_IR_REG_28__SCAN_IN;
  assign n9995 = n9994 & n9248;
  assign n11068 = n11063 | P2_IR_REG_6__SCAN_IN;
  assign n10540 = ~n10455 & ~n10454;
  assign n11406 = ~n11403 & ~P2_IR_REG_28__SCAN_IN;
  assign n10036 = n10074 & n10035;
  assign n11018 = ~n9073 | ~n9072;
  assign n10230 = ~n10229 | ~n10228;
  assign n10153 = n10151 & n10150;
  assign n10161 = n10159 & n10158;
  assign n9248 = ~n9368 | ~SI_2_;
  assign n16154 = ~n11800 | ~P1_U3086;
  assign n11403 = ~n8946 | ~n9103;
  assign n8905 = n9828 & n9690;
  assign n10039 = ~n10003 | ~n10002;
  assign n11165 = ~n17335;
  assign n17341 = ~n9525 | ~P2_U3151;
  assign n17338 = n11800 & P2_U3151;
  assign n9360 = n17335;
  assign n17335 = ~n11028 | ~n11045;
  assign n11572 = n11513 & n11512;
  assign n9848 = ~n9846 & ~n9845;
  assign n10978 = ~n10967 | ~n10966;
  assign n10967 = n10965 & n10964;
  assign n9837 = n9835 & n9834;
  assign n11045 = ~n11023 | ~n11025;
  assign n9990 = ~n9876 | ~n9818;
  assign n9818 = ~P1_IR_REG_2__SCAN_IN;
  assign n10965 = ~P2_IR_REG_5__SCAN_IN & ~P2_IR_REG_4__SCAN_IN;
  assign P2_U3151 = ~P2_STATE_REG_SCAN_IN;
  assign n10053 = P1_REG3_REG_4__SCAN_IN & P1_REG3_REG_5__SCAN_IN;
  assign n10168 = ~P1_IR_REG_8__SCAN_IN;
  assign n9876 = ~P1_IR_REG_1__SCAN_IN & ~P1_IR_REG_0__SCAN_IN;
  assign n9823 = ~P1_IR_REG_5__SCAN_IN & ~P1_IR_REG_4__SCAN_IN;
  assign n9820 = ~P1_IR_REG_3__SCAN_IN & ~P1_IR_REG_6__SCAN_IN;
  assign n9851 = ~P1_IR_REG_21__SCAN_IN & ~P1_IR_REG_20__SCAN_IN;
  assign n9852 = ~P1_IR_REG_22__SCAN_IN & ~P1_IR_REG_23__SCAN_IN;
  assign n9819 = ~P1_IR_REG_10__SCAN_IN & ~P1_IR_REG_9__SCAN_IN;
  assign n9881 = P2_ADDR_REG_19__SCAN_IN & P1_ADDR_REG_19__SCAN_IN;
  assign n9835 = ~P1_IR_REG_17__SCAN_IN & ~P1_IR_REG_19__SCAN_IN;
  assign n9834 = ~P1_IR_REG_16__SCAN_IN & ~P1_IR_REG_15__SCAN_IN;
  assign n13440 = ~n13149 | ~n13151;
  assign n13375 = ~n9055 | ~n9052;
  assign n9363 = ~n9879 | ~n9878;
  assign n9890 = ~n8886 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n9301 = n13256;
  assign n8892 = n10596;
  assign n8893 = n10596;
  assign n10596 = n9906 & n9907;
  assign n16676 = ~n11125 ^ n12064;
  assign n8894 = ~n9920;
  assign n8897 = n9907 & n9910;
  assign n12595 = n17151 | n17365;
  assign n9795 = ~n14741 | ~n11955;
  assign n10128 = ~n9920 | ~n12871;
  assign n10475 = n10477 & n10444;
  assign n14043 = ~n14067 | ~n12509;
  assign n12509 = n12508 & n14066;
  assign n16295 = ~n13122 | ~n13382;
  assign n12724 = n14269 | n8890;
  assign n9640 = n9641 & n12768;
  assign n13254 = ~n14704 & ~n9301;
  assign n12855 = ~n8976 | ~n9526;
  assign n9526 = ~n12486 | ~n9527;
  assign n13034 = n13035 | n11906;
  assign n9583 = n12450 | n12452;
  assign n9244 = n11978 & n9245;
  assign n9246 = ~n13440;
  assign n9408 = ~n11904 | ~n15889;
  assign n15935 = ~n15975 | ~n13034;
  assign n9525 = ~n9894;
  assign n9321 = n12942 & n12984;
  assign n12831 = ~n17538 | ~n9510;
  assign n12451 = ~n17029 | ~n12446;
  assign n14730 = n9680 & n11985;
  assign n11985 = ~n9814 & ~n11984;
  assign n13091 = n16258 | n15729;
  assign n9560 = n14721 & n14756;
  assign n11955 = ~n14756 | ~n14773;
  assign n9229 = n15872 & n13047;
  assign n11991 = n16034 | n16029;
  assign n9540 = ~n9541 | ~n10781;
  assign n12481 = n14146 | n17541;
  assign n9731 = ~n9732 & ~n12228;
  assign n9456 = ~n9458 | ~n9457;
  assign n11513 = ~n9500 & ~n9499;
  assign n9499 = ~n9502 | ~n11410;
  assign n9500 = ~n11458 | ~n9501;
  assign n12184 = ~n12179;
  assign n12534 = n13785 & n12533;
  assign n17015 = ~n9436 | ~n9439;
  assign n9439 = n9440 & n12667;
  assign n9440 = ~n9441 | ~n17030;
  assign n9737 = n11368 & n9738;
  assign n9530 = n9531 & n11869;
  assign n9531 = ~n9534 | ~n9536;
  assign n10980 = n9462 & n10959;
  assign n9462 = n10996 & n10958;
  assign n9867 = ~n9866 | ~n13008;
  assign n10849 = n12345 | n8880;
  assign n11933 = ~n14961 | ~n14998;
  assign n9564 = ~n15732;
  assign n14755 = ~n14779 | ~n14778;
  assign n14817 = ~n16406;
  assign n9774 = n9775 & n11932;
  assign n9775 = ~n9776 | ~n14994;
  assign n9776 = ~n11930;
  assign n11931 = ~n15007 | ~n11929;
  assign n11929 = ~n15024 | ~n14997;
  assign n9766 = ~n10437 | ~n10436;
  assign n10227 = ~n10161 | ~n10160;
  assign n10190 = n10156 & n10155;
  assign n13601 = ~n13518 ^ n13602;
  assign n13739 = ~n12481 | ~n12482;
  assign n12936 = ~n12486 | ~n12485;
  assign n12566 = ~P2_REG3_REG_28__SCAN_IN & ~n12358;
  assign n9430 = n9431 & n12926;
  assign n9127 = ~n9126 | ~n9124;
  assign n9431 = ~n9433 | ~n9432;
  assign n14068 = n12504 & n12964;
  assign n17365 = n9100 & n12047;
  assign n9100 = n9101 & n12046;
  assign n11766 = n9156 | n11071;
  assign n9156 = ~n11020 & ~n9157;
  assign n9157 = ~n11000 | ~n9158;
  assign n10520 = n10474 | n10477;
  assign n9119 = n9765 & n9120;
  assign n9765 = n8948 & n10436;
  assign n15052 = ~n10823 | ~n10822;
  assign n9921 = n9920;
  assign n12402 = ~n12399;
  assign n9221 = n11954 & n9222;
  assign n9218 = ~n14792 | ~n9219;
  assign n15732 = n15788 | n16258;
  assign n9212 = n9213 & n9783;
  assign n9214 = ~n9211 | ~n9210;
  assign n13382 = ~n9841 ^ n9692;
  assign n13051 = n13054 & n13050;
  assign n9743 = ~n9744 & ~n13148;
  assign n9184 = n9621 & n12687;
  assign n9619 = ~n9184 | ~n9620;
  assign n9620 = ~n12682;
  assign n9628 = ~n12728;
  assign n9629 = n9371 & n12731;
  assign n9287 = ~n9293 | ~n13185;
  assign n13205 = n9284 & n13204;
  assign n9746 = n9748 & n13217;
  assign n9378 = ~n9643;
  assign n12805 = n12818 | n12828;
  assign n9505 = ~n12821 & ~n12824;
  assign n9257 = n9751 & n13253;
  assign n9751 = ~n13255 & ~n9756;
  assign n9411 = ~n9412 | ~n12969;
  assign n9412 = ~n13998 & ~n9413;
  assign n9413 = ~n14071;
  assign n11971 = n11968 & n15760;
  assign n9084 = n12930 & n9085;
  assign n9086 = ~n12925;
  assign n12944 = ~n14136 & ~n17551;
  assign n10964 = ~P2_IR_REG_6__SCAN_IN & ~P2_IR_REG_3__SCAN_IN;
  assign n9258 = n9255 & n9260;
  assign n9814 = ~n13459 & ~n14744;
  assign n9242 = ~n9670;
  assign n9676 = n9677 & n13426;
  assign n9238 = n9676 & n13418;
  assign n9384 = ~n9385 & ~SI_14_;
  assign n9385 = ~n10420;
  assign n9822 = ~P1_IR_REG_7__SCAN_IN;
  assign n9882 = ~n9881 | ~n9880;
  assign n9878 = ~P2_ADDR_REG_19__SCAN_IN;
  assign n9879 = ~P1_ADDR_REG_19__SCAN_IN & ~P1_RD_REG_SCAN_IN;
  assign n9732 = ~n12239;
  assign n9727 = ~n12284;
  assign n9598 = ~n11129 | ~n16713;
  assign n9647 = n11055 & n9652;
  assign n9652 = ~n16740;
  assign n9610 = n9611 & n9615;
  assign n9615 = ~n16777;
  assign n9485 = n16848 | n16830;
  assign n9115 = ~n11140 | ~n11222;
  assign n9479 = n9480 | n16921;
  assign n9480 = ~n11258;
  assign n9280 = ~n16919;
  assign n9279 = n16919 | n11251;
  assign n9508 = n11411 & n9509;
  assign n9509 = ~P2_REG3_REG_10__SCAN_IN;
  assign n9580 = ~n12480 | ~n8968;
  assign n9067 = ~n9584 | ~n8967;
  assign n12464 = ~n13972 | ~n13969;
  assign n13972 = ~n8922 | ~n12462;
  assign n12435 = ~n12434 & ~n9810;
  assign n12434 = n12460 | n12433;
  assign n9071 = ~n9810;
  assign n9070 = ~n13998 | ~n12458;
  assign n9077 = ~n8923 | ~n12452;
  assign n12961 = n16442 | n16573;
  assign n12450 = n12449 | n12448;
  assign n12634 = n17102 | n17396;
  assign n12636 = ~n17102 | ~n17396;
  assign n17075 = ~n9062 | ~n9060;
  assign n9060 = ~n8980 & ~n9061;
  assign n9062 = ~n17096 | ~n12439;
  assign n10429 = ~n10433 & ~SI_15_;
  assign n11004 = ~P2_IR_REG_9__SCAN_IN;
  assign n11953 = ~n14778 | ~n14622;
  assign n13354 = n12402 | n12398;
  assign n9664 = ~n9668 | ~n9665;
  assign n9666 = ~n9668;
  assign n9388 = ~n9390 | ~n9392;
  assign n9199 = ~n9200 | ~n11938;
  assign n13335 = n15102 | n14865;
  assign n9779 = n9780 & n11943;
  assign n13418 = n9297 | n14457;
  assign n11973 = ~n15818 | ~n11967;
  assign n15842 = ~n13047 | ~n13406;
  assign n11962 = n15871 & n13401;
  assign n9292 = n15904 & n13397;
  assign n15871 = n13395 & n9317;
  assign n9317 = ~n13397 | ~n9318;
  assign n9318 = ~n13390;
  assign n9787 = n9788 & n9847;
  assign n9788 = n9663 & n9789;
  assign n9331 = ~n8940 & ~n9332;
  assign n9332 = ~n10686;
  assign n10681 = n10648 & n10649;
  assign n10683 = n10653 | n8934;
  assign n10590 = n10588 & n10587;
  assign n10421 = n10420 & n10419;
  assign n9713 = ~n9716 & ~n9714;
  assign n12123 = ~n16612 | ~n9735;
  assign n9735 = ~n12113 & ~n9736;
  assign n9736 = ~n12096;
  assign n9725 = n9727 & n8914;
  assign n9414 = n9415 & n12984;
  assign n9415 = ~n12983 & ~n9416;
  assign n9416 = ~n9417 | ~n13739;
  assign n12979 = n12978 & n9418;
  assign n9418 = ~n13806 & ~n9419;
  assign n9304 = n9321 & n12937;
  assign n9091 = ~n12946 | ~n9092;
  assign n9092 = n12945 & n11770;
  assign n9512 = ~n9516 | ~n9513;
  assign n9513 = ~P2_REG3_REG_22__SCAN_IN;
  assign n9517 = ~P2_REG3_REG_23__SCAN_IN;
  assign n11413 = ~n11878;
  assign n11038 = n17343 | n11037;
  assign n9468 = ~n11171;
  assign n9653 = n11056 & P2_REG2_REG_5__SCAN_IN;
  assign n9458 = n9460 & n11184;
  assign n9460 = ~n16734;
  assign n9475 = n16771 | n16791;
  assign n9473 = n11207 & n9474;
  assign n9474 = ~n16791;
  assign n9139 = ~n16787 | ~P2_REG1_REG_9__SCAN_IN;
  assign n16831 = ~n11220 & ~n16813;
  assign n9518 = ~n12255 & ~P2_REG3_REG_22__SCAN_IN;
  assign n12255 = P2_REG3_REG_21__SCAN_IN | n12244;
  assign n11536 = n11534 | P2_REG3_REG_14__SCAN_IN;
  assign n11411 = ~P2_REG3_REG_9__SCAN_IN;
  assign n11495 = ~n11572 | ~n9508;
  assign n17029 = n17051 | n12445;
  assign n11512 = ~P2_REG3_REG_8__SCAN_IN;
  assign n17155 = ~n12437 | ~n12436;
  assign n13833 = ~n9126 | ~n12919;
  assign n13879 = ~n13883;
  assign n12897 = n12493 | n9801;
  assign n17464 = ~n17203;
  assign n9074 = n11017 & n9622;
  assign n10979 = ~n10978;
  assign n11005 = ~P2_IR_REG_10__SCAN_IN;
  assign n9357 = ~n11051;
  assign n11025 = ~P2_IR_REG_2__SCAN_IN;
  assign n9688 = ~n11300;
  assign n9936 = n9710 & n9931;
  assign n14587 = ~n10278 ^ n10861;
  assign n10277 = ~n10824 | ~n16279;
  assign n9178 = ~n16304 | ~n10824;
  assign n9167 = ~n10677;
  assign n9177 = ~n10512 | ~n10511;
  assign n15369 = ~n10028 | ~n10027;
  assign n9052 = ~n9053 | ~n8925;
  assign n9056 = ~n8971 | ~n13277;
  assign n10666 = n10627 & P1_REG3_REG_20__SCAN_IN;
  assign n9773 = ~n9774 | ~n9777;
  assign n9561 = ~n9563 & ~n9562;
  assign n9210 = ~n15813;
  assign n9551 = ~n15924;
  assign n15071 = ~n14778;
  assign n9196 = n14937 | n9200;
  assign n9195 = ~n11937 | ~n9198;
  assign n15135 = ~n14924;
  assign n9554 = ~n15178 & ~n9555;
  assign n14994 = ~n13440 | ~n13278;
  assign n9202 = ~n15639 | ~n9203;
  assign n11921 = ~n16292 | ~n14457;
  assign n15788 = ~n15786 | ~n15785;
  assign n9896 = ~P1_IR_REG_28__SCAN_IN;
  assign n10842 = ~n10815 | ~n10814;
  assign n9539 = n9540 & n10812;
  assign n9858 = ~n8974 | ~n8905;
  assign n16087 = ~n10290 ^ n10324;
  assign n9329 = ~n10284;
  assign n10225 = ~n10224;
  assign n10120 = ~n10119;
  assign n10146 = ~n10148 ^ n10127;
  assign n16555 = ~n16612 | ~n12096;
  assign n9141 = ~n12310 | ~n13689;
  assign n13505 = ~n9144 | ~n9143;
  assign n9143 = ~n8977 | ~n13637;
  assign n9144 = ~n16581 | ~n9145;
  assign n14186 = ~n12254 | ~n12253;
  assign n13518 = ~n9148 | ~n8972;
  assign n9148 = ~n9146 | ~n9730;
  assign n13604 = ~n13601 & ~n17525;
  assign n13886 = ~n17522;
  assign n12055 = n16496 | n16495;
  assign n9152 = ~n9153 | ~n8954;
  assign n11414 = ~n14362;
  assign n16660 = ~n16658 & ~n16657;
  assign n9454 = ~n9461 | ~n9458;
  assign n16772 = ~n11201 & ~n11200;
  assign n16846 = n11085 ^ n17283;
  assign n16904 = ~n11250 & ~n11249;
  assign n11145 = ~n9131 | ~n11144;
  assign n16943 = ~n16817;
  assign n11112 = ~n12185 & ~n11111;
  assign n11113 = ~n9262 & ~n11265;
  assign n9658 = n11112 & n9659;
  assign n14146 = ~n12347 | ~n12346;
  assign n13776 = ~n17538;
  assign n13828 = n13833 | n12515;
  assign n13871 = ~n12241 | ~n12240;
  assign n13919 = ~n12514 | ~n12900;
  assign n9449 = ~n12906 & ~n9450;
  assign n9450 = ~n12904;
  assign n13909 = ~n17519;
  assign n14249 = ~n12189 | ~n12188;
  assign n14032 = ~n14270;
  assign n14067 = ~n17015 | ~n12500;
  assign n9345 = ~n12503 & ~n12962;
  assign n11410 = ~P2_REG3_REG_5__SCAN_IN;
  assign n9496 = ~P2_REG3_REG_4__SCAN_IN;
  assign n16522 = ~n12081 | ~n12080;
  assign n9645 = n12065 & n8924;
  assign n13500 = n12554 & n12553;
  assign n12576 = ~n12564;
  assign n9108 = ~n13738 ^ n13739;
  assign n9296 = ~n13753 ^ n12980;
  assign n17452 = ~n17238 | ~n17232;
  assign n11014 = ~n11403 | ~P2_IR_REG_31__SCAN_IN;
  assign n9322 = ~n10971 & ~n10972;
  assign n10987 = ~n10968 | ~P2_IR_REG_31__SCAN_IN;
  assign n9718 = ~n11007 & ~P2_IR_REG_23__SCAN_IN;
  assign n9722 = ~n11007;
  assign n10479 = n10519 & n10473;
  assign n9338 = ~n10477;
  assign n9696 = n9697 & n10810;
  assign n9697 = ~n9699 | ~n9698;
  assign n14773 = ~n16412;
  assign n14865 = ~n16400;
  assign n15882 = ~n16216;
  assign n15011 = ~n13151;
  assign n14998 = n10496 & n10495;
  assign n14455 = n10348 & n10347;
  assign n10204 = ~n8893 | ~P1_REG1_REG_8__SCAN_IN;
  assign n10194 = n10167 & n10166;
  assign n14705 = ~n13261 | ~n13260;
  assign n13261 = n15241 | n10128;
  assign n9556 = ~n14704 | ~n9557;
  assign n9557 = ~n9559;
  assign n9791 = ~n11957 & ~n9792;
  assign n14720 = ~n14755 & ~n15061;
  assign n15056 = ~n14736 & ~n14735;
  assign n10451 = n17259 | n8880;
  assign n10408 = ~n10341 | ~n10340;
  assign n13105 = ~n16279;
  assign n15697 = ~n9564 | ~n9565;
  assign n9565 = ~n9562;
  assign n10199 = n17306 | n8880;
  assign n9235 = n10128 | n12066;
  assign n9236 = n10482 | n9974;
  assign n15036 = ~n13274 | ~n9921;
  assign n13273 = n15232 | n13271;
  assign n9399 = ~n15056;
  assign n9228 = ~n9795 | ~n11956;
  assign n9225 = ~n14792 | ~n11951;
  assign n16225 = ~n15983 | ~n16295;
  assign n12392 = n10903 & n16162;
  assign n11873 = ~n9905 | ~n15236;
  assign n14196 = ~n12265 | ~n12264;
  assign n16496 = ~n12053 ^ n17151;
  assign n13609 = ~n14186;
  assign n13693 = n11792 & n17120;
  assign n16610 = n11786 & n11785;
  assign n9364 = n12992 | n17243;
  assign n17544 = n12363 | n12362;
  assign n17529 = ~n12262 | ~n12261;
  assign n12262 = n13817 | n12256;
  assign n11896 = ~n11150 | ~n11151;
  assign n17120 = ~n13492 | ~n17350;
  assign n12296 = ~n10813 ^ n10811;
  assign n10813 = ~n9538 | ~n9541;
  assign n9538 = ~n9544 | ~n10782;
  assign n9544 = ~n10752;
  assign n10531 = n11959;
  assign n15917 = n16295 | n10922;
  assign n17560 = ~n11850 & ~n11849;
  assign n11849 = ~n17562 & ~n17561;
  assign n17608 = ~n11854 & ~n11853;
  assign n13025 = n11910 | n8881;
  assign n13084 = ~n13414 | ~n9301;
  assign n9250 = n9251 & n13072;
  assign n13142 = n9763 | n9301;
  assign n9660 = n12649 & n12656;
  assign n12682 = ~n12681 | ~n12680;
  assign n9742 = n9336 & n9341;
  assign n13159 = n9672 | n13157;
  assign n12707 = ~n9617 | ~n9618;
  assign n9618 = n9619 & n12690;
  assign n9625 = n9627 & n12736;
  assign n9627 = ~n9629 | ~n9628;
  assign n9314 = n9750 & n9749;
  assign n13213 = n13212 & n14768;
  assign n9642 = ~n12757;
  assign n9643 = n12760 & n9644;
  assign n9373 = ~n9376 | ~n12805;
  assign n9376 = ~n12790 | ~n9377;
  assign n9528 = ~n12485;
  assign n9423 = ~n14126;
  assign n9504 = n9505 & n8931;
  assign n9350 = n13435 & n9351;
  assign n9351 = ~n15008;
  assign n12914 = n12910 & n12909;
  assign n12862 = ~n8969 | ~n9529;
  assign n9529 = ~n12855;
  assign n9348 = ~n14888;
  assign n9255 = ~n9752 & ~n9256;
  assign n9259 = ~n9254 | ~n9753;
  assign n9753 = n9755 & n9754;
  assign n10658 = n10656 & n10655;
  assign n12971 = n12967 & n9410;
  assign n9410 = ~n14024 & ~n9411;
  assign n9082 = ~n12928;
  assign n9638 = ~n16883;
  assign n12471 = n12470 | n12469;
  assign n12472 = ~n9067 | ~n8966;
  assign n12431 = n14269 & n14280;
  assign n9681 = n9815 & n13336;
  assign n9247 = n8928 & n11980;
  assign n9669 = ~n14861 | ~n13327;
  assign n9197 = ~n9201 & ~n9198;
  assign n9201 = ~n11938;
  assign n9670 = ~n9672 & ~n9671;
  assign n9671 = ~n13278;
  assign n13412 = n11969 & n13294;
  assign n13292 = ~n15759 | ~n15763;
  assign n9545 = n9807 & n10524;
  assign n10234 = n10232 & n10231;
  assign n9522 = ~n10124 | ~n8984;
  assign n12122 = n12121 | n16560;
  assign n9419 = ~n13829 | ~n9420;
  assign n9420 = ~n9421 & ~n13859;
  assign n9421 = ~n13835;
  assign n11040 = ~n17335 | ~P2_REG2_REG_2__SCAN_IN;
  assign n9457 = ~n16755;
  assign n9435 = ~n12923 | ~n12515;
  assign n9516 = n13610 & n9517;
  assign n9495 = ~n11448 & ~P2_REG3_REG_17__SCAN_IN;
  assign n9507 = ~P2_REG3_REG_11__SCAN_IN;
  assign n9576 = n9581 | n9577;
  assign n12920 = n14196 | n13862;
  assign n12919 = n13871 | n13886;
  assign n9447 = n9140 & n13879;
  assign n12912 = n13895 | n13909;
  assign n9584 = ~n12464 | ~n8991;
  assign n9585 = ~n13945;
  assign n9441 = ~n12643;
  assign n9437 = ~n12956 & ~n9438;
  assign n9438 = ~n12642;
  assign n12606 = ~n12438 | ~n16590;
  assign n17096 = ~n17155 | ~n17154;
  assign n9738 = ~P2_D_REG_0__SCAN_IN;
  assign n9534 = n9535 & n11867;
  assign n9535 = ~n10840 | ~n10843;
  assign n10966 = ~P2_IR_REG_8__SCAN_IN & ~P2_IR_REG_7__SCAN_IN;
  assign n9702 = ~n10315;
  assign n9865 = n11959 | n13376;
  assign n9169 = ~n14572;
  assign n9172 = ~n9176 & ~n9173;
  assign n9176 = ~n10576;
  assign n9173 = ~n10511;
  assign n9174 = ~n10576 | ~n9175;
  assign n9694 = n9817 & n10585;
  assign n9175 = ~n14504;
  assign n9761 = ~n10261;
  assign n9053 = ~n9054 | ~n13262;
  assign n9057 = ~n8898 | ~n9058;
  assign n13323 = n15036 & n16427;
  assign n13236 = ~n15052 & ~n14625;
  assign n13242 = n15052 & n14625;
  assign n14744 = n11983 | n11982;
  assign n13343 = n15071 | n14622;
  assign n9569 = ~n9571 | ~n9570;
  assign n9571 = ~n9572;
  assign n14889 = ~n9243 | ~n9240;
  assign n9240 = n9241 & n8989;
  assign n9243 = ~n14995 | ~n9244;
  assign n14909 = n14936 & n14946;
  assign n14936 = n15146 | n14972;
  assign n9203 = ~n9207 & ~n9204;
  assign n9204 = ~n11925;
  assign n9205 = ~n11927 | ~n9206;
  assign n9206 = ~n11926;
  assign n15616 = ~n9673 | ~n9237;
  assign n9673 = n9674 & n13422;
  assign n9237 = ~n9238 | ~n9239;
  assign n9394 = ~n11923 | ~n9395;
  assign n9395 = ~n11922;
  assign n9796 = ~n9799 | ~n11919;
  assign n13414 = ~n9282 | ~n9261;
  assign n9261 = n15734 & n10267;
  assign n15725 = ~n13292;
  assign n15763 = ~n11964 | ~n11963;
  assign n10522 = n10521 & n10551;
  assign n10442 = n10440 & n10439;
  assign n9381 = ~n9384 | ~n9382;
  assign n9382 = ~n10426;
  assign n9824 = ~P1_IR_REG_11__SCAN_IN;
  assign n9847 = ~n9990 & ~n9821;
  assign n10150 = ~n12871 | ~P2_DATAO_REG_8__SCAN_IN;
  assign n10049 = ~n12871 | ~P2_DATAO_REG_6__SCAN_IN;
  assign n10148 = ~n10126 | ~n10125;
  assign n10125 = ~n12871 | ~P2_DATAO_REG_7__SCAN_IN;
  assign n9521 = ~n10124 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n9734 = ~n16582 | ~n12146;
  assign n9145 = n13637 & n12146;
  assign n9716 = ~n9717 & ~n8926;
  assign n9717 = ~n13706;
  assign n9146 = ~n12212;
  assign n9147 = ~n9730 | ~n8973;
  assign n9728 = ~n9732 & ~n9729;
  assign n11471 = n11572 & n9506;
  assign n9506 = n8945 & n11580;
  assign n11534 = ~n11471 | ~n11470;
  assign n16645 = n11158 & n11161;
  assign n16665 = ~n16638 | ~n11039;
  assign n9290 = ~P2_REG1_REG_2__SCAN_IN;
  assign n9275 = ~n9273 | ~n12064;
  assign n9273 = ~n11044;
  assign n11133 = ~n11132 | ~n11131;
  assign n9359 = ~n8899 | ~n11066;
  assign n9649 = ~n9652 | ~n9650;
  assign n9455 = ~n9457 | ~n11192;
  assign n9616 = ~n9359 | ~n17313;
  assign n9483 = n8981 | n11233;
  assign n9482 = ~n16831 & ~n9485;
  assign n11142 = ~n9603 | ~n11141;
  assign n9133 = ~n11143 | ~n11235;
  assign n9477 = ~n9479 | ~n9019;
  assign n9476 = ~n16904 & ~n9481;
  assign n9276 = ~n11100 | ~n9280;
  assign n12358 = P2_REG3_REG_27__SCAN_IN | n12326;
  assign n9432 = ~n12923;
  assign n9124 = ~n9434 & ~n9125;
  assign n9125 = ~n12919;
  assign n12314 = ~n12255 & ~n9514;
  assign n9514 = ~n9516 | ~n9515;
  assign n9515 = ~P2_REG3_REG_22__SCAN_IN & ~P2_REG3_REG_25__SCAN_IN;
  assign n12234 = ~n12220 & ~P2_REG3_REG_19__SCAN_IN;
  assign n12220 = ~n9495 | ~n9494;
  assign n11590 = ~n9495;
  assign n11438 = ~n11536 & ~P2_REG3_REG_15__SCAN_IN;
  assign n12506 = n14093 & n9344;
  assign n11581 = n11572 & n8945;
  assign n9061 = ~n17381 & ~n16543;
  assign n9646 = ~P1_DATAO_REG_3__SCAN_IN;
  assign n9065 = ~n9582 & ~n9064;
  assign n13753 = ~n13752 | ~n13751;
  assign n9063 = ~n9066 & ~n9064;
  assign n9066 = ~n12477;
  assign n13835 = n12920 & n13827;
  assign n13924 = n9584 & n13944;
  assign n12511 = n12897 & n13971;
  assign n13948 = ~n12464 | ~n12463;
  assign n13996 = ~n12435;
  assign n9069 = ~n13995 & ~n9070;
  assign n14099 = ~n9075 | ~n12456;
  assign n9075 = ~n9078 | ~n9076;
  assign n9076 = n9077 & n12455;
  assign n9343 = ~n12961 | ~n14119;
  assign n14125 = n16987 | n12452;
  assign n16987 = n12451 & n12450;
  assign n12443 = n12442 | n17082;
  assign n17081 = ~n12497 | ~n12496;
  assign n12497 = ~n9102 | ~n8997;
  assign n9102 = ~n17127 | ~n17129;
  assign n17126 = ~n12615 | ~n12623;
  assign n17129 = ~n17126;
  assign n10973 = ~P2_IR_REG_20__SCAN_IN & ~P2_IR_REG_23__SCAN_IN;
  assign n10976 = ~n10963 | ~n11009;
  assign n9719 = n9720 & n9721;
  assign n9720 = ~n10976 & ~n10978;
  assign n9721 = ~n11045;
  assign n10436 = n10435 & n10434;
  assign n9121 = ~n10421;
  assign n10471 = n10469 & n10468;
  assign n11072 = ~n10978 & ~n11045;
  assign n11024 = n11023 | n11071;
  assign n11031 = ~P2_IR_REG_0__SCAN_IN | ~P2_IR_REG_31__SCAN_IN;
  assign n9698 = ~n14466;
  assign n10725 = n10705 & P1_REG3_REG_22__SCAN_IN;
  assign n9165 = ~n9167 | ~n9166;
  assign n9166 = ~n10678 | ~n9169;
  assign n10795 = n10764 & P1_REG3_REG_24__SCAN_IN;
  assign n10863 = ~n10118;
  assign n13369 = n13321 & n9324;
  assign n9324 = ~n9349 & ~n9325;
  assign n10106 = ~n8892 | ~P1_REG1_REG_7__SCAN_IN;
  assign n13367 = ~n11991;
  assign n9559 = ~n12399 | ~n9560;
  assign n9792 = ~n11955;
  assign n13349 = n15061 | n14773;
  assign n9219 = ~n9224 & ~n9220;
  assign n9220 = ~n11951;
  assign n9222 = ~n9223 | ~n11953;
  assign n9223 = ~n11952;
  assign n10827 = n10795 & P1_REG3_REG_25__SCAN_IN;
  assign n14801 = ~n14923 & ~n9567;
  assign n9567 = ~n9568 | ~n14822;
  assign n9568 = ~n9569;
  assign n10764 = n10725 & P1_REG3_REG_23__SCAN_IN;
  assign n10627 = ~n10600 & ~n10599;
  assign n13173 = ~n15124 | ~n14866;
  assign n10600 = ~n10564 | ~P1_REG3_REG_18__SCAN_IN;
  assign n14938 = n8978 & n9552;
  assign n9552 = n15613 & n14961;
  assign n10455 = n10408 | n10407;
  assign n16304 = ~n10297 | ~n10296;
  assign n9562 = ~n16271 | ~n8970;
  assign n9783 = ~n9784 & ~n11918;
  assign n9784 = ~n13091;
  assign n9215 = ~n11915;
  assign n9406 = n13285 & n13286;
  assign n13285 = ~n13390 | ~n13393;
  assign n15974 = ~n9316 | ~n16173;
  assign n9316 = ~n15980;
  assign n13012 = ~n12407 | ~n12406;
  assign n9558 = ~n9560;
  assign n9793 = ~n14731 & ~n9794;
  assign n9794 = ~n11956;
  assign n14731 = ~n13236 & ~n13242;
  assign n14779 = n14801 & n14802;
  assign n15082 = ~n14802;
  assign n14815 = ~n9294 | ~n8928;
  assign n9390 = n9391 & n11944;
  assign n14923 = n14921 | n15135;
  assign n14970 = ~n11976 | ~n13278;
  assign n15643 = ~n13302 & ~n13301;
  assign n11920 = ~n15745 & ~n15746;
  assign n15786 = ~n9548 & ~n11996;
  assign n9549 = ~n16227 & ~n9550;
  assign n9230 = ~n13047 | ~n9231;
  assign n13282 = ~n15974;
  assign n9045 = ~n12870;
  assign n9044 = n9045 | n12875;
  assign n9901 = ~n9769 & ~P1_IR_REG_28__SCAN_IN;
  assign n9902 = ~P1_IR_REG_29__SCAN_IN;
  assign n10935 = ~n9870 ^ n9896;
  assign n9874 = ~P1_IR_REG_27__SCAN_IN;
  assign n9871 = ~P1_IR_REG_26__SCAN_IN;
  assign n9843 = n9852 & n9851;
  assign n10648 = n10612 & n10613;
  assign n10652 = n10617 | n10616;
  assign n9690 = n9827 & n9691;
  assign n9691 = ~P1_IR_REG_13__SCAN_IN;
  assign n10551 = n10520 & n10519;
  assign n10224 = ~n10227 | ~n10163;
  assign n12161 = n12157 | n12847;
  assign n9160 = ~n12063;
  assign n14231 = ~n12209 | ~n12208;
  assign n13533 = ~n9155 | ~n8993;
  assign n12203 = n12202 | n12201;
  assign n12053 = ~n12348 ^ n17365;
  assign n14258 = ~n12177 | ~n12176;
  assign n11781 = n11764 | n17349;
  assign n12226 = n12212 & n13531;
  assign n13862 = ~n17525;
  assign n16580 = n16581 | n16582;
  assign n13691 = ~n9723 | ~n9724;
  assign n9724 = ~n8908 | ~n8914;
  assign n12987 = n12982 & n9414;
  assign n9094 = ~n9093 & ~n9087;
  assign n9087 = ~n9091 | ~n9088;
  assign n9088 = n9089 & n12989;
  assign n12289 = n9518 & n9517;
  assign n14050 = n11476 & n11475;
  assign n13644 = n11587 & n11586;
  assign n9428 = n11482 & n11481;
  assign n16638 = ~n11038 | ~n9630;
  assign n9630 = ~n9631 & ~n9632;
  assign n9631 = ~n11039;
  assign n9633 = ~n11038 | ~n11039;
  assign n16697 = ~n12072 ^ n11173;
  assign n16722 = ~n9466 | ~n9465;
  assign n9465 = ~n9467 | ~n11179;
  assign n16735 = ~n9461 | ~n11184;
  assign n16758 = ~n11133 ^ n11197;
  assign n16792 = ~n9472 & ~n11207;
  assign n9263 = ~n9264 | ~P2_REG2_REG_9__SCAN_IN;
  assign n9471 = n9473 | n11214;
  assign n9470 = ~n16772 & ~n9475;
  assign n11139 = ~n9604 | ~n11138;
  assign n16849 = ~n9484 & ~n11228;
  assign n9268 = n9272 | n9024;
  assign n9269 = ~n9271 | ~n9270;
  assign n9272 = ~n16846;
  assign n16922 = ~n9478 & ~n11258;
  assign n9593 = ~n11152;
  assign n9594 = ~n11283 & ~n9595;
  assign n9595 = ~n11897;
  assign n9592 = ~n9596 | ~n11152;
  assign n13740 = ~n17544;
  assign n12313 = n12311 | n12847;
  assign n12298 = n12296 | n12847;
  assign n14221 = ~n12215 | ~n12214;
  assign n12215 = n12213 | n12847;
  assign n13961 = ~n12183 | ~n12182;
  assign n14008 = ~n14259;
  assign n17463 = ~n12145 | ~n12144;
  assign n11493 = ~n11572 | ~n11411;
  assign n17166 = ~n14049;
  assign n17147 = n17452 | n12895;
  assign n14142 = n13719 | n13718;
  assign n13880 = ~n9446 | ~n12911;
  assign n13970 = ~n9096 & ~n9095;
  assign n9095 = ~n12897;
  assign n9096 = ~n12898;
  assign n17422 = n12106 & n12105;
  assign n17414 = n12101 & n12100;
  assign n12584 = n17185 | n11783;
  assign n12869 = ~n12842 | ~n12841;
  assign n12841 = n12838 | n12840;
  assign n9059 = ~n12838 ^ n12839;
  assign n9073 = ~n9074 | ~n8946;
  assign n9622 = n9623 & n10979;
  assign n9623 = n9463 & n10959;
  assign n9463 = n9464 & n10996;
  assign n9464 = n10958 & n11013;
  assign n11013 = ~P2_IR_REG_26__SCAN_IN;
  assign n9104 = ~n9624;
  assign n9541 = n9542 & n10784;
  assign n9543 = ~n10751;
  assign n9047 = n9048 & n10749;
  assign n9050 = ~n9051 | ~n10693;
  assign n16768 = ~n11070 ^ P2_IR_REG_8__SCAN_IN;
  assign n11069 = n11068 | P2_IR_REG_7__SCAN_IN;
  assign n12077 = ~n11052 ^ P2_IR_REG_5__SCAN_IN;
  assign n9137 = n11025 & n9138;
  assign n9323 = ~n16202;
  assign n15268 = ~n9682 | ~n9684;
  assign n10917 = n9695 & n9162;
  assign n9162 = ~n12019 & ~n9163;
  assign n14446 = n10313 & n14590;
  assign n14449 = n10316 & n10317;
  assign n9708 = ~n9709 & ~n8963;
  assign n9709 = ~n9931;
  assign n9693 = ~n10585;
  assign n14553 = n10357 | n10356;
  assign n9707 = ~n14395;
  assign n14570 = ~n9167 | ~n10679;
  assign n16094 = ~n10283 ^ n10284;
  assign n15347 = ~n11298 | ~n11300;
  assign n9758 = n9759 & n10531;
  assign n15012 = n10376 & n10375;
  assign n14457 = n10255 & n10254;
  assign n10081 = ~n8892 | ~P1_REG1_REG_5__SCAN_IN;
  assign n9956 = ~n8892 | ~P1_REG1_REG_1__SCAN_IN;
  assign n10167 = n10067 & n10031;
  assign n10237 = n10236 | P1_IR_REG_9__SCAN_IN;
  assign n9772 = n9773 & n11933;
  assign n15022 = ~n15613 | ~n11997;
  assign n9208 = ~n15639 | ~n11925;
  assign n10341 = n10268 & n10247;
  assign n9563 = n16304;
  assign n15708 = ~n15732 & ~n15737;
  assign n15746 = n11968 & n13294;
  assign n10200 = ~n10108 & ~n10107;
  assign n15975 = ~n15968 | ~n13282;
  assign n15977 = ~n16170;
  assign n15968 = ~n13283;
  assign n15992 = ~n15023;
  assign n15043 = ~n14705;
  assign n9771 = n11931 | n9777;
  assign n14982 = ~n15613 | ~n9554;
  assign n10006 = n9993 & n9992;
  assign n15233 = ~P1_IR_REG_30__SCAN_IN;
  assign n9043 = n12869 & n9036;
  assign n9036 = ~n9044;
  assign n9040 = ~n9042 | ~n9041;
  assign n9041 = ~n9045 | ~n12875;
  assign n9042 = n12868 | n9044;
  assign n9046 = ~n12869;
  assign n11868 = ~n9533 | ~n10843;
  assign n15431 = n10935;
  assign n17219 = ~n10750 ^ n10748;
  assign n10332 = ~n9828 | ~n9827;
  assign n10030 = n9990 | P1_IR_REG_3__SCAN_IN;
  assign n12066 = ~n9402 ^ n9401;
  assign n9403 = ~n9973 | ~n9972;
  assign n13931 = ~n14231;
  assign n16473 = ~n17053;
  assign n14175 = ~n12286 | ~n12285;
  assign n13560 = ~n9726 & ~n12284;
  assign n9726 = ~n13518 & ~n12276;
  assign n13607 = ~n13604 & ~n13603;
  assign n13655 = ~n13547 | ~n12239;
  assign n16574 = n12335 | n12334;
  assign n9149 = ~n9151 & ~n9150;
  assign n9151 = ~n16608;
  assign n9150 = ~n12086;
  assign n16609 = n9152 & n12086;
  assign n13707 = ~n9715 & ~n8926;
  assign n17547 = n12543 & n12542;
  assign n17541 = n12331 | n12330;
  assign n17538 = ~n12315 | ~n9511;
  assign n9511 = ~n12318 & ~n9023;
  assign n17535 = n12307 | n12306;
  assign n17532 = n12294 | n12293;
  assign n17522 = n12248 | n12247;
  assign n17519 = n12238 | n12237;
  assign n17516 = n12225 | n12224;
  assign n13904 = ~n13951;
  assign n14270 = n11445 | n11444;
  assign n14291 = n11540 | n11539;
  assign n17465 = ~n14050;
  assign n9099 = n11485 & n9574;
  assign n9574 = ~n8975 | ~n11414;
  assign n16756 = n9454 & n9459;
  assign n16917 = ~n11146 | ~n11147;
  assign n9657 = ~n11115;
  assign n14136 = ~n12878 | ~n12179;
  assign n13805 = ~n13828 | ~n12923;
  assign n13801 = ~n17535;
  assign n13824 = ~n17532;
  assign n14061 = n11528 & n11527;
  assign n14094 = ~n9345;
  assign n17196 = ~n17123;
  assign n11504 = ~n9498 | ~n9502;
  assign n9498 = n11458 & n11410;
  assign n11561 = ~n11458 | ~n11410;
  assign n17197 = ~n17120;
  assign n13501 = ~n12580 | ~n12579;
  assign n14150 = n9108 & n9107;
  assign n17350 = n11772 & n11325;
  assign n11405 = ~n14354 | ~P2_IR_REG_31__SCAN_IN;
  assign n15241 = ~n12869 ^ n12868;
  assign n11407 = n11406 | n11071;
  assign n17214 = ~n10988 ^ P2_IR_REG_25__SCAN_IN;
  assign n11323 = ~n10987 ^ n10969;
  assign n17232 = ~n11010 ^ n11009;
  assign n11003 = ~n11001 | ~P2_IR_REG_31__SCAN_IN;
  assign n17243 = ~n11766 ^ n11765;
  assign n9337 = ~n10479 & ~n9338;
  assign n17307 = ~n16768;
  assign n17325 = ~n12077;
  assign n16135 = ~n10073 ^ n10071;
  assign n9342 = n17343;
  assign n15254 = ~n9689 | ~n10104;
  assign n14721 = ~n15052;
  assign n14924 = n10537 & n10536;
  assign n10537 = n17248 | n8880;
  assign n15381 = ~n15311;
  assign n14610 = n10561 & n10560;
  assign n10561 = n17253 | n8880;
  assign n10792 = n12296 | n8880;
  assign n9319 = ~n14620 ^ n9320;
  assign n9320 = ~n14621;
  assign n15333 = n10923 & n15917;
  assign n16415 = n10831 | n10830;
  assign n16412 = n10800 | n10799;
  assign n16409 = n10769 | n10768;
  assign n16406 = n10710 | n10709;
  assign n16403 = n10730 | n10729;
  assign n16400 = n10671 | n10670;
  assign n16394 = n10605 | n10604;
  assign n16391 = n10544 | n10543;
  assign n16388 = n10569 | n10568;
  assign n13151 = n10460 | n10459;
  assign n15661 = ~n14455;
  assign n15711 = ~n14457;
  assign n9306 = ~n10012 & ~n8916;
  assign n9310 = n11906;
  assign n15035 = ~n14706 ^ n9035;
  assign n14706 = ~n8918 & ~n14705;
  assign n12006 = n12005 | n12004;
  assign n15695 = ~n15732 & ~n9566;
  assign n9566 = ~n16271 | ~n13105;
  assign n16004 = ~n12015 | ~n15917;
  assign n9398 = ~n9399 & ~n15055;
  assign n15076 = ~n15075 & ~n15074;
  assign n15232 = ~n9039 | ~n9037;
  assign n9037 = ~n9046 | ~n9038;
  assign n9039 = ~n9043 & ~n9040;
  assign n9038 = n12868 & n12875;
  assign n17562 = ~n11848 & ~n11847;
  assign n17558 = ~n11852 & ~n11851;
  assign n11851 = ~n17560 & ~n17559;
  assign n17604 = ~n17606 & ~n11855;
  assign n17596 = ~n17598 & ~n11857;
  assign n9186 = ~n8911 | ~n9018;
  assign n9134 = ~n9135 | ~n16937;
  assign n9135 = ~n11896 ^ n11897;
  assign n9295 = ~n13769 | ~n8964;
  assign n15737 = ~n16271;
  assign n8898 = ~n9253 & ~n8998;
  assign n8899 = n9651 & n9649;
  assign n8900 = n14704 | n13122;
  assign n15674 = ~n9797 & ~n9017;
  assign n8901 = n9634 & n9639;
  assign n8902 = n16680 & n11179;
  assign n8903 = n9487 & n9028;
  assign n8906 = n11900 & n16862;
  assign n8907 = n12597 & n9800;
  assign n8908 = n13559 | n8962;
  assign n13419 = ~n15659 | ~n9305;
  assign n11940 = ~n9196 | ~n8949;
  assign n10720 = ~n8878;
  assign n13283 = n11907 & n9217;
  assign n13149 = ~n15167;
  assign n8910 = n11924 & n9394;
  assign n8911 = n13003 | P2_STATE_REG_SCAN_IN;
  assign n8912 = n8911 & n12999;
  assign n8913 = n9031 & n9592;
  assign n8914 = n12295 | n17532;
  assign n8915 = ~n15157 | ~n14998;
  assign n8916 = n8891 & P1_REG1_REG_4__SCAN_IN;
  assign n13855 = n9067 & n13922;
  assign n13998 = n12429 & n12462;
  assign n11458 = n9497 & n9496;
  assign n8917 = n9981 & n9982;
  assign n8918 = n14755 | n9556;
  assign n8919 = n16279 | n15734;
  assign n8920 = n11488 & n11487;
  assign n8921 = n17132 | n17389;
  assign n12303 = n11531;
  assign n8922 = n12461 & n9068;
  assign n9899 = n9869 & n9768;
  assign n8923 = n9583 & n12453;
  assign n16292 = ~n9297;
  assign n9297 = ~n10245 | ~n10244;
  assign n10124 = ~n9894;
  assign n8924 = n12205 | n9646;
  assign n9200 = ~n11937;
  assign n16227 = ~n13056;
  assign n8925 = n13276 & n13363;
  assign n8926 = ~n12163 & ~n14291;
  assign n12985 = ~n12936 ^ n13740;
  assign n9417 = ~n12985;
  assign n8927 = n11479 & n9428;
  assign n9325 = ~n13322;
  assign n14741 = ~n9218 | ~n9221;
  assign n14835 = ~n9387 | ~n9390;
  assign n14072 = ~n12459 | ~n12458;
  assign n14908 = ~n9194 | ~n11937;
  assign n14960 = ~n9771 | ~n9774;
  assign n14887 = ~n11940 | ~n11939;
  assign n9198 = ~n11936;
  assign n10482 = ~n9920 | ~n13271;
  assign n8928 = n9664 & n13335;
  assign n8929 = n14705 ^ n16424;
  assign n8930 = n16768 | n17022;
  assign n14997 = n10413 & n10412;
  assign n8931 = n12820 | n12819;
  assign n8932 = ~n12085 & ~n17102;
  assign n9782 = ~n15795;
  assign n8933 = n10085 & P1_REG2_REG_1__SCAN_IN;
  assign n8934 = n10652 & n10651;
  assign n8935 = n13040 & n13041;
  assign n8936 = n12862 & n12854;
  assign n8937 = n12805 & n9640;
  assign n8938 = n9390 & n9199;
  assign n8939 = n9260 & n13253;
  assign n8940 = ~n10684 & ~n10683;
  assign n8941 = n10190 & n10149;
  assign n8942 = n13197 & n13196;
  assign n10611 = ~n9546 | ~n10524;
  assign n10682 = ~n10611;
  assign n8943 = n9598 & n11130;
  assign n8944 = n13213 & n9750;
  assign n8945 = n9508 & n9507;
  assign n8946 = n10977 & n9322;
  assign n8947 = n9388 & n11945;
  assign n8948 = n10475 & n10479;
  assign n8949 = n9195 & n11938;
  assign n8950 = n13306 & n13305;
  assign n9699 = n14621 & n10780;
  assign n8951 = n11895 | n11894;
  assign n8952 = n11972 & n15709;
  assign n8953 = n12722 & n12721;
  assign n8954 = ~n16538 & ~n12083;
  assign n8955 = n14409 & n10576;
  assign n8956 = n9328 & n12986;
  assign n10292 = ~n9663 | ~n9847;
  assign n9828 = ~n10292;
  assign n9665 = ~n13327;
  assign n8957 = n13064 & n13063;
  assign n8958 = n9882 & P1_DATAO_REG_3__SCAN_IN;
  assign n8959 = n13144 & n13143;
  assign n8960 = n9379 & n12889;
  assign n8961 = n9625 & n9192;
  assign n9459 = ~n11192;
  assign n15092 = ~n14822;
  assign n9433 = ~n9434;
  assign n9434 = ~n12925 | ~n9435;
  assign n8962 = n9727 & n12276;
  assign n9581 = ~n9582;
  assign n9582 = ~n12480 | ~n12477;
  assign n8963 = ~n11296 & ~n11604;
  assign n9570 = ~n15102;
  assign n14559 = n10303 & n10302;
  assign n9305 = ~n14559;
  assign n8964 = n13762 & n13761;
  assign n12263 = ~n12847;
  assign n11058 = ~n9356;
  assign n9356 = ~n9357 | ~n11046;
  assign n8965 = ~n11013 | ~n11012;
  assign n10716 = ~n10685 | ~n9331;
  assign n9051 = ~n10716;
  assign n8966 = n12466 & n13922;
  assign n8967 = n13923 & n13944;
  assign n8968 = ~n13751 | ~n12478;
  assign n8969 = ~n12936 | ~n17544;
  assign n8970 = n16292 & n13105;
  assign n17330 = ~n12064;
  assign n8971 = ~n13276 | ~n13270;
  assign n8972 = n9147 & n12252;
  assign n13397 = ~n16202 | ~n11905;
  assign n8973 = ~n9728 | ~n13531;
  assign n8974 = n9838 & n9692;
  assign n12399 = n10849 & n10848;
  assign n8975 = n11413 & P2_REG0_REG_1__SCAN_IN;
  assign n8976 = n17544 | n12887;
  assign n8977 = ~n9734 | ~n12154;
  assign n9872 = ~n9868 | ~P1_IR_REG_31__SCAN_IN;
  assign n8978 = n9554 & n13149;
  assign n8979 = n9793 | n11957;
  assign n8980 = n17111 & n17132;
  assign n15157 = ~n10489 | ~n10488;
  assign n9049 = ~n10717;
  assign n8981 = ~n16848 & ~n9486;
  assign n8982 = n9115 & n16843;
  assign n8983 = ~n14020 & ~n12460;
  assign n8984 = SI_0_ & P1_DATAO_REG_1__SCAN_IN;
  assign n8985 = n14923 | n9569;
  assign n8986 = n12957 | n9422;
  assign n8987 = ~n11100 & ~n9278;
  assign n8988 = n12862 & n12931;
  assign n8989 = n11979 & n13446;
  assign n8990 = n11020 | P2_IR_REG_18__SCAN_IN;
  assign n8991 = n9585 & n12463;
  assign n8992 = n9230 & n13406;
  assign n15061 = ~n14756;
  assign n8993 = n9154 & n12203;
  assign n8994 = n11928 & n9205;
  assign n8995 = n12897 & n12972;
  assign n8996 = n8919 & n11921;
  assign n8997 = n8921 & n12623;
  assign n8998 = n14705 & n13122;
  assign n12594 = ~n17151 | ~n17365;
  assign n13179 = ~n13174 | ~n13175;
  assign n8999 = n9813 & n12948;
  assign n9000 = n10104 & n10142;
  assign n9001 = n9586 & n9813;
  assign n9002 = n12867 & n12866;
  assign n9003 = ~n12924 | ~n12923;
  assign n9004 = n12678 & n12677;
  assign n9005 = n12752 & n12751;
  assign n9006 = n14923 | n9572;
  assign n9007 = ~n12250 | ~n13654;
  assign n9008 = ~n12192 | ~n12193;
  assign n9009 = ~P2_IR_REG_31__SCAN_IN | ~n11015;
  assign n12692 = n17463 & n13644;
  assign n9344 = ~n12692;
  assign n9010 = n9761 & n10227;
  assign n9011 = n10737 & n9168;
  assign n9012 = n9694 & n9174;
  assign n9756 = ~n16421;
  assign n9013 = n9576 & n12481;
  assign n9014 = ~n11942 | ~n11939;
  assign n9015 = n9381 & n10430;
  assign n9714 = ~n12173;
  assign n12173 = n12170 | n14061;
  assign n9016 = n9902 & n9896;
  assign n10545 = ~n10118;
  assign n9017 = ~n9796 | ~n8919;
  assign n9018 = ~n13002 & ~n13001;
  assign n9692 = ~P1_IR_REG_20__SCAN_IN;
  assign n13009 = n11959 | n13477;
  assign n9019 = n17260 | n11264;
  assign n17051 = n12444 & n12443;
  assign n15007 = ~n9202 | ~n8994;
  assign n9020 = n9271 & n9267;
  assign n9501 = ~P2_REG3_REG_7__SCAN_IN;
  assign n9502 = ~P2_REG3_REG_6__SCAN_IN;
  assign n9021 = n9233 & n13398;
  assign n9022 = n16888 | n11243;
  assign n9510 = ~n14155;
  assign n9608 = ~P2_REG2_REG_3__SCAN_IN;
  assign n9497 = ~P2_REG3_REG_3__SCAN_IN;
  assign n9023 = n12327 & P2_REG2_REG_27__SCAN_IN;
  assign n17449 = n17083 & n17440;
  assign n9107 = ~n17449;
  assign n9024 = ~n11231 & ~n11085;
  assign n9025 = n9239 & n13418;
  assign n9026 = ~n11920 & ~n11919;
  assign n9027 = n16865 | n8913;
  assign n9028 = n9805 & n11290;
  assign n9596 = ~n11283;
  assign n17238 = ~n11003 ^ n11002;
  assign n13376 = ~n9839 ^ P1_IR_REG_21__SCAN_IN;
  assign n16034 = ~n13376;
  assign n9494 = ~P2_REG3_REG_18__SCAN_IN;
  assign n9029 = n9613 & n9616;
  assign n17294 = ~n10262 ^ n10261;
  assign n9307 = ~n11910;
  assign n9030 = ~n11897 & ~n9593;
  assign n9031 = n9596 | n9030;
  assign n9032 = ~n9547 & ~n11996;
  assign n9033 = ~n13484 & ~n16034;
  assign n9034 = n9596 | n9593;
  assign n16385 = ~n16383;
  assign n16165 = ~n16008 | ~n16007;
  assign n16008 = n13383 & n11600;
  assign n9527 = ~n12865 & ~n9528;
  assign n17205 = ~n12865 & ~n12896;
  assign n12808 = n14165 | n12865;
  assign n16338 = ~n16326;
  assign n9035 = ~n15036;
  assign n9048 = ~n9049 | ~n10693;
  assign n10750 = ~n10718 | ~n10693;
  assign n10718 = ~n10716 | ~n10717;
  assign n9054 = ~n13269 | ~n14705;
  assign n9055 = ~n9057 | ~n9056;
  assign n9058 = ~n13269 | ~n15043;
  assign n12842 = ~n9059 | ~SI_29_;
  assign n12484 = ~n9059 ^ SI_29_;
  assign n17097 = ~n9061;
  assign n12444 = ~n17075 | ~n12440;
  assign n9579 = ~n12476 | ~n12949;
  assign n13752 = ~n12476 | ~n9063;
  assign n9064 = ~n12949;
  assign n9575 = ~n12476 | ~n9065;
  assign n13770 = ~n9579 ^ n13786;
  assign n9586 = ~n9587 | ~n12472;
  assign n9068 = ~n12459 | ~n9069;
  assign n13995 = ~n8983 | ~n9071;
  assign n9452 = ~n8946 | ~n9622;
  assign n9072 = ~n9009 | ~n11017;
  assign n9078 = ~n12451 | ~n8923;
  assign n9079 = ~n16141 | ~n8882;
  assign n12935 = ~n9083 | ~n9080;
  assign n9080 = n9081 & n12932;
  assign n9081 = ~n9084 | ~n9082;
  assign n9083 = ~n9003 | ~n9084;
  assign n9085 = ~n12928 | ~n9086;
  assign n9089 = ~n9090 | ~n11117;
  assign n9090 = ~n12945;
  assign n9093 = ~n12946 & ~n11770;
  assign n12992 = ~n12991 & ~n9094;
  assign n9098 = ~n12898 | ~n8995;
  assign n12910 = ~n9097 | ~n12908;
  assign n9097 = ~n9098 | ~n12970;
  assign n9101 = ~n12050 | ~n12051;
  assign n9429 = ~n9102 | ~n12623;
  assign n10981 = ~n8946 | ~n9104;
  assign n9105 = ~n16917 | ~n16916;
  assign n9106 = ~n16758 | ~P2_REG1_REG_7__SCAN_IN;
  assign n13748 = n9108 & n14097;
  assign n9111 = ~n11126 | ~n9602;
  assign n9112 = ~n9113 | ~n11126;
  assign n9113 = ~n16676;
  assign n16844 = ~n9114 | ~n11140;
  assign n9114 = ~n16826 | ~P2_REG1_REG_11__SCAN_IN;
  assign n9603 = ~n9116 | ~n8982;
  assign n9117 = ~n11140;
  assign n10437 = ~n9118 | ~n10428;
  assign n9118 = ~n10422 | ~n10421;
  assign n9120 = ~n10428 | ~n9121;
  assign n9122 = ~n9123 | ~n10428;
  assign n9123 = ~n10422;
  assign n9129 = ~n16864;
  assign n9131 = ~n9130 | ~n9128;
  assign n9128 = ~n9129 | ~n11143;
  assign n16881 = ~n9132 | ~n11143;
  assign n9132 = ~n16864 | ~P2_REG1_REG_13__SCAN_IN;
  assign P2_U3200 = ~n9136 | ~n9134;
  assign n11051 = ~n9137 | ~n11023;
  assign n9138 = ~P2_IR_REG_3__SCAN_IN;
  assign n11023 = ~P2_IR_REG_1__SCAN_IN & ~P2_IR_REG_0__SCAN_IN;
  assign n16787 = ~n11136 ^ n11211;
  assign n11136 = ~n9600 | ~n11135;
  assign n9140 = ~n13918 | ~n12911;
  assign n12344 = ~n9141 | ~n12322;
  assign n12321 = ~n9141 & ~n12322;
  assign n9142 = ~n12038 | ~n12037;
  assign n16581 = ~n12132 | ~n12131;
  assign n9153 = ~n16539;
  assign n9155 = ~n12164 | ~n9712;
  assign n9154 = ~n9712 | ~n9714;
  assign n11001 = ~n11766 | ~n11765;
  assign n9158 = ~P2_IR_REG_18__SCAN_IN;
  assign n16459 = ~n9161 | ~n12063;
  assign n16458 = ~n9161 | ~n9159;
  assign n9159 = ~n16460 & ~n9160;
  assign n9161 = ~n16594 | ~n16593;
  assign n9164 = ~n9695 | ~n9696;
  assign n9163 = ~n9696;
  assign n12020 = ~n9164 | ~n12019;
  assign n10747 = ~n9165 | ~n9011;
  assign n9170 = ~n14571 | ~n14572;
  assign n14571 = ~n10677 | ~n10678;
  assign n9168 = n10678 | n9169;
  assign n10738 = n14570 & n9170;
  assign n10646 = ~n9171 | ~n9012;
  assign n9171 = ~n10512 | ~n9172;
  assign n14409 = ~n9177 | ~n14504;
  assign n10305 = ~n9178 | ~n10304;
  assign n9181 = ~n9179 | ~n12815;
  assign n9179 = ~n9503 | ~n12806;
  assign n12860 = ~n9180 | ~n12835;
  assign n9180 = ~n9182 | ~n9181;
  assign n9182 = ~n9183 | ~n9504;
  assign n9183 = ~n12830 | ~n12829;
  assign n9617 = ~n12679 | ~n9184;
  assign n9187 = ~n9185 | ~n8912;
  assign n9185 = ~n9365 | ~n9364;
  assign P2_U3296 = ~n9187 | ~n9186;
  assign n9191 = ~n9190 | ~n9188;
  assign n9188 = n9189 & n12746;
  assign n9189 = ~n8961 | ~n9626;
  assign n9190 = ~n9362 | ~n12743;
  assign n12753 = ~n9191 | ~n12750;
  assign n12740 = ~n9626 | ~n9625;
  assign n9192 = ~n12739;
  assign n9389 = ~n9193 | ~n8938;
  assign n9193 = ~n14937 | ~n9197;
  assign n9194 = ~n14937 | ~n11936;
  assign n15614 = ~n9208 | ~n11926;
  assign n9207 = ~n11927;
  assign n9213 = ~n11915 | ~n9782;
  assign n9216 = ~n9210 | ~n9209;
  assign n9209 = ~n11912;
  assign n9211 = ~n11912 & ~n15795;
  assign n9786 = ~n9214 | ~n9212;
  assign n9785 = ~n9409 | ~n9782;
  assign n9409 = ~n9216 | ~n9215;
  assign n15969 = ~n15966 | ~n13283;
  assign n11907 = ~n9303 | ~n13035;
  assign n9217 = ~n11906 | ~n16182;
  assign n14767 = ~n9225 | ~n11952;
  assign n9224 = ~n11953;
  assign n9226 = ~n9795 | ~n9793;
  assign n9227 = ~n9228 | ~n14731;
  assign n9233 = ~n11962 | ~n15872;
  assign n9232 = ~n9229 | ~n11962;
  assign n9231 = ~n13398;
  assign n9239 = ~n15678 | ~n13416;
  assign n9241 = ~n9244 | ~n9242;
  assign n9245 = ~n9670 | ~n9246;
  assign n14947 = ~n11976 | ~n9670;
  assign n11976 = ~n14995 | ~n13440;
  assign n11981 = ~n9294 | ~n9247;
  assign n9680 = ~n11981 | ~n9681;
  assign n9402 = ~n9403 | ~n9248;
  assign n9252 = ~n9249 | ~n13062;
  assign n9249 = n13061 & n13069;
  assign n13082 = ~n9252 | ~n9250;
  assign n9251 = ~n8957 | ~n13069;
  assign n15889 = ~n15934 | ~n16202;
  assign n9253 = ~n13277;
  assign n9254 = ~n9260 | ~n9257;
  assign n9256 = ~n13253;
  assign n13258 = ~n9259 & ~n9258;
  assign n16940 = ~n9262 ^ P2_REG2_REG_17__SCAN_IN;
  assign n9262 = ~n11111 ^ n12185;
  assign n16751 = ~n9359 ^ n17313;
  assign n9264 = ~n16789;
  assign n16789 = ~n9266 ^ n17301;
  assign n9265 = ~n9266 | ~n17301;
  assign n9266 = ~n9614 | ~n8930;
  assign n9267 = ~n11082;
  assign n9270 = ~n11082 & ~n9024;
  assign n11043 = ~n9275;
  assign n11050 = ~n16693 | ~n16694;
  assign n16693 = ~n9274 | ~n9607;
  assign n9274 = ~n9275 | ~P2_REG2_REG_3__SCAN_IN;
  assign n9277 = n16901 | n9279;
  assign n11107 = ~n9277 | ~n9276;
  assign n9278 = ~n16901 & ~n11251;
  assign n9341 = ~n9745 | ~n9743;
  assign n9745 = ~n8959 | ~n13148;
  assign n9281 = ~n10388 | ~n10389;
  assign n9391 = ~n9779 | ~n9014;
  assign n9349 = ~n13474 | ~n8929;
  assign n13042 = n13033 & n13032;
  assign n9283 = ~n17294;
  assign n10054 = n9907 & n9910;
  assign n16182 = ~n9952 | ~n9951;
  assign n9953 = ~n10007 | ~P1_REG0_REG_1__SCAN_IN;
  assign n9284 = ~n13203 | ~n13202;
  assign n9285 = ~n10654 | ~n10683;
  assign n13190 = ~n13186 | ~n9286;
  assign n9286 = ~n9287 | ~n13179;
  assign n9573 = ~n15124;
  assign n11028 = ~n11027 | ~n11026;
  assign n9288 = P2_IR_REG_0__SCAN_IN;
  assign n9339 = ~n13037 ^ n13122;
  assign n9291 = ~n9289 | ~n13115;
  assign n9289 = ~n13097 | ~n13096;
  assign n13036 = ~n15974 | ~n13034;
  assign n11150 = ~n16936 | ~P2_REG1_REG_17__SCAN_IN;
  assign n16864 = ~n11142 ^ n11238;
  assign n11124 = ~n16663 | ~n16662;
  assign n16662 = ~n17335 ^ n9290;
  assign n17343 = ~n11036 | ~n11035;
  assign n9358 = n9637 & n9022;
  assign n13126 = ~n9291 | ~n9353;
  assign n9299 = ~n13038;
  assign n15872 = ~n9292 | ~n15935;
  assign n9293 = ~n9302 | ~n13184;
  assign n12838 = ~n9532 | ~n9530;
  assign n9759 = ~n9760 | ~n16034;
  assign n12894 = ~n12893 | ~n12892;
  assign n12893 = ~n8960 | ~n9327;
  assign n9532 = ~n10842 | ~n9534;
  assign n13039 = ~n9300;
  assign n14863 = ~n13325 | ~n13173;
  assign n13007 = ~n13005 & ~n15961;
  assign n13136 = ~n9555 | ~n15012;
  assign P2_U3206 = n13763 | n9295;
  assign n13760 = ~n14159 & ~n13758;
  assign n13755 = ~n9296 | ~n17172;
  assign n13054 = ~n13049 | ~n13048;
  assign n9300 = ~n13025 | ~n13024;
  assign n13406 = ~n15876 | ~n13056;
  assign n9983 = n9980 & n9979;
  assign n14382 = ~n10738;
  assign n10257 = ~n10824 | ~n9297;
  assign n9503 = ~n9374 | ~n9373;
  assign n12244 = ~n12234 | ~n12233;
  assign n12267 = ~n9518;
  assign n13031 = ~n13028 | ~n9298;
  assign n9298 = ~n9300 | ~n9299;
  assign n9302 = ~n13448 | ~n13183;
  assign n13423 = ~n16304 | ~n14559;
  assign n12898 = ~n14043 | ~n12510;
  assign n12924 = n12922 | n12921;
  assign n9436 = ~n17058 | ~n9437;
  assign n12918 = ~n12914 & ~n12913;
  assign n9957 = ~n9955 & ~n8933;
  assign n9427 = ~n17167;
  assign n12946 = ~n12938 | ~n9304;
  assign n10085 = n9910 & n11873;
  assign n9405 = ~n9407 & ~n9408;
  assign n9798 = ~n11920 | ~n9799;
  assign n9880 = ~P2_RD_REG_SCAN_IN;
  assign n9303 = ~n11906;
  assign n13448 = ~n9573 | ~n16394;
  assign n15678 = ~n8952 | ~n11973;
  assign n14467 = ~n10747 | ~n10746;
  assign n17058 = ~n12498 | ~n12636;
  assign n17168 = n11426 | n11425;
  assign n9315 = ~n10478 | ~n9337;
  assign n9404 = ~n9405 | ~n15892;
  assign n15892 = ~n15907 | ~n9406;
  assign n15745 = ~n9786 | ~n13075;
  assign n12401 = ~n9790 | ~n8979;
  assign n13023 = ~n9307 | ~n8881;
  assign n13085 = n11959 & n16029;
  assign n10382 = ~n10358 | ~n14553;
  assign n10824 = n10189;
  assign n9374 = ~n9372 | ~n8937;
  assign n15346 = ~n9962 | ~n9961;
  assign n9492 = ~n12860 | ~n12859;
  assign n12602 = ~n9308 | ~n12596;
  assign n9308 = ~n8907 | ~n12594;
  assign n17167 = ~n8927 | ~n11480;
  assign n9353 = n9312 & n13118;
  assign n10677 = ~n10646 | ~n10645;
  assign n13052 = ~n13042 | ~n9309;
  assign n9309 = ~n9339 | ~n8935;
  assign n10358 = ~n9703 | ~n9311;
  assign n9311 = n9701 & n14554;
  assign n9312 = ~n13119 | ~n13120;
  assign n10702 = ~n9313 | ~n10720;
  assign n9313 = ~n17219;
  assign n9748 = ~n9314 | ~n13213;
  assign n13422 = ~n16315 | ~n14455;
  assign n16828 = ~n11081 ^ n17289;
  assign n11111 = ~n11107 & ~n11106;
  assign n9939 = ~n9885 | ~n9884;
  assign n9930 = ~n9926 | ~n9925;
  assign n14995 = ~n11975 | ~n13307;
  assign n12409 = ~n11986 | ~n13351;
  assign n9868 = ~n9787 | ~n9848;
  assign n14633 = ~n9319 | ~n15376;
  assign n13148 = ~n13147 | ~n13146;
  assign n9553 = ~n15167;
  assign n9973 = ~n9994 | ~n9996;
  assign n9996 = n9887 & n9812;
  assign n13099 = n13087 & n13086;
  assign n13314 = ~n14814 & ~n13313;
  assign n9599 = n9326 | n16714;
  assign n16714 = ~n11128 ^ n12077;
  assign n9326 = ~n11129;
  assign n9347 = ~n14862 | ~n9348;
  assign n17174 = ~n9427 | ~n17195;
  assign n9396 = ~n9798 | ~n9393;
  assign n9407 = ~n15890;
  assign n10283 = ~n9369 | ~n10320;
  assign n9327 = ~n8956 | ~n12863;
  assign n9328 = ~n12861 | ~n12862;
  assign n9372 = ~n12753;
  assign n9426 = ~n17177 | ~n12595;
  assign n9362 = ~n12740 | ~n12739;
  assign n11974 = ~n15616 | ~n13427;
  assign n13040 = ~n13030 | ~n13029;
  assign n10226 = ~n10157 | ~n10156;
  assign n16962 = ~n12960 | ~n9343;
  assign n12504 = ~n9345 | ~n9344;
  assign n17127 = ~n17141 | ~n12606;
  assign n10285 = ~n9330 | ~n9329;
  assign n9330 = ~n10283;
  assign n9686 = ~n15344;
  assign n12021 = ~n10917;
  assign n9334 = ~n14467;
  assign n9684 = ~n9687 | ~n9685;
  assign n13623 = ~n12226;
  assign n9672 = ~n8915;
  assign n9386 = ~n10361 | ~n10426;
  assign n9962 = n9333 & n9937;
  assign n9333 = ~n9936 | ~n10803;
  assign n9695 = ~n9334 | ~n9699;
  assign P2_U3201 = ~n11154 | ~n9335;
  assign n17154 = ~n12607 | ~n12606;
  assign n9710 = ~n10189 | ~n16173;
  assign n16590 = ~n12060 | ~n12059;
  assign n17259 = ~n9766 ^ n10475;
  assign n9706 = ~n10282;
  assign n9519 = ~n10000 | ~n9999;
  assign n13264 = n10085;
  assign n9655 = ~n9658 & ~n9657;
  assign n13269 = ~n13258 & ~n13257;
  assign n9336 = ~n13156 | ~n13155;
  assign n9369 = ~n9762 | ~n9010;
  assign n9840 = ~n8905 | ~n9838;
  assign n9355 = ~n9340 | ~n13374;
  assign n9340 = ~n9757 | ~n9758;
  assign n12129 = ~n9283 | ~n12263;
  assign n11120 = n17343 | n11119;
  assign n9685 = ~n9686 & ~n9688;
  assign n10483 = ~n10446 & ~P1_IR_REG_16__SCAN_IN;
  assign n11129 = ~n11128 | ~n17325;
  assign n13313 = ~n9346;
  assign n9760 = ~n9033 & ~n8909;
  assign n13309 = ~n8950 | ~n9350;
  assign n13161 = ~n9352 | ~n9742;
  assign n9352 = ~n13145 | ~n9741;
  assign n9747 = ~n9354 | ~n8944;
  assign n9354 = ~n13195 | ~n13194;
  assign n9361 = ~n9355 | ~n13381;
  assign n9611 = ~n9616 | ~n11193;
  assign n9639 = ~n11092;
  assign n13491 = ~n9361 | ~n13384;
  assign n9370 = ~n10147 | ~n10146;
  assign n9894 = ~n9363 | ~n9882;
  assign n9764 = ~n8958 | ~n9363;
  assign n9365 = ~n9367 | ~n9366;
  assign n9366 = ~n9605 | ~n9493;
  assign n9367 = ~n9606 | ~n12896;
  assign n9998 = ~n9368 & ~SI_2_;
  assign n9972 = ~n9368 ^ n9891;
  assign n10326 = ~n9369 | ~n10322;
  assign n10157 = ~n9370 | ~n8941;
  assign n10191 = ~n9370 | ~n10149;
  assign n9371 = ~n8953 | ~n12728;
  assign n12826 = ~n9375 | ~n9640;
  assign n9375 = ~n12753 | ~n9643;
  assign n9377 = ~n9640 | ~n9378;
  assign n9379 = ~n12986 | ~n9002;
  assign n9383 = ~n9380 | ~n9384;
  assign n9380 = ~n10361;
  assign n10389 = ~n9383 | ~n9015;
  assign n9387 = n11940 | n9392;
  assign n11947 = ~n9389 | ~n8947;
  assign n9392 = ~n9779;
  assign n9397 = ~n9798 | ~n8904;
  assign n9393 = n8904 & n11923;
  assign n15660 = ~n9397 | ~n11922;
  assign n15639 = ~n9396 | ~n8910;
  assign n15195 = ~n15193 | ~n16338;
  assign n15193 = ~n9400 | ~n9398;
  assign n9401 = ~n9997;
  assign n15813 = ~n9404 | ~n11911;
  assign n15794 = ~n9409;
  assign n9422 = ~n9424 | ~n9423;
  assign n9424 = ~n12956 & ~n9425;
  assign n9425 = ~n17014 | ~n16992;
  assign n17141 = ~n17142 | ~n9426;
  assign n17143 = ~n17142 & ~n9426;
  assign n12494 = ~n17174;
  assign n17388 = ~n9429 ^ n17107;
  assign n9442 = ~n17058 | ~n12642;
  assign n17027 = ~n9442 | ~n12643;
  assign n9446 = ~n13919 | ~n12975;
  assign n9448 = ~n12911;
  assign n9451 = ~n13947 | ~n12899;
  assign n12514 = ~n9451 | ~n9449;
  assign n13941 = ~n9451 | ~n12904;
  assign n11809 = ~n10985 | ~n9452;
  assign n11201 = ~n9453 | ~n9455;
  assign n9453 = n11185 | n9456;
  assign n9461 = ~n11185;
  assign n9469 = ~n16681 | ~n16680;
  assign n9466 = ~n16681 | ~n8902;
  assign n16705 = ~n9469 | ~n11171;
  assign n16816 = ~n9470 & ~n9471;
  assign n9472 = ~n16772 & ~n16771;
  assign n16942 = ~n9476 & ~n9477;
  assign n9478 = ~n16904 & ~n16903;
  assign n9481 = n16921 | n16903;
  assign n16868 = ~n9482 & ~n9483;
  assign n9484 = ~n16831 & ~n16830;
  assign n9486 = ~n11228;
  assign n12863 = ~n9490 | ~n9488;
  assign n9488 = ~n9489 | ~n12858;
  assign n9489 = ~n9492 | ~n8936;
  assign n9490 = ~n9491 | ~n12853;
  assign n9491 = ~n9492 | ~n8988;
  assign n9606 = ~n9493 | ~n12894;
  assign n9493 = ~n12891 | ~n9804;
  assign n12299 = n12255 | n9512;
  assign n10045 = ~n9519 | ~n10036;
  assign n10073 = ~n9519 | ~n10035;
  assign n10123 = ~n9520 | ~n10120;
  assign n12090 = ~n9520 ^ n10119;
  assign n9938 = ~n9883 | ~n9521;
  assign n9886 = ~n9523 | ~n9522;
  assign n9523 = ~n9524 | ~SI_0_;
  assign n9524 = ~n9883;
  assign n9533 = ~n10842 | ~n10841;
  assign n9536 = ~n10843;
  assign n9537 = ~n10752 | ~n9541;
  assign n10815 = ~n9537 | ~n9539;
  assign n10783 = ~n10752 | ~n10751;
  assign n9542 = ~n9543 | ~n10782;
  assign n10685 = ~n9546 | ~n9545;
  assign n15884 = n11996 | n15924;
  assign n9547 = ~n9551 | ~n13056;
  assign n9548 = ~n9551 | ~n9549;
  assign n9550 = ~n13065;
  assign n14984 = ~n8978 | ~n15613;
  assign n14703 = ~n14755 & ~n9559;
  assign n14875 = ~n14923 & ~n15124;
  assign n9572 = ~n9573 | ~n14876;
  assign n13729 = ~n9575 | ~n9580;
  assign n12483 = ~n9578 | ~n9013;
  assign n9577 = ~n9580;
  assign n9578 = ~n9579 | ~n9580;
  assign n12476 = ~n9586 | ~n8999;
  assign n13834 = ~n12472 | ~n12471;
  assign n9587 = ~n9588 & ~n12473;
  assign n9588 = ~n12471;
  assign n11153 = ~n9589 | ~n9591;
  assign n16738 = ~n9597 | ~n11129;
  assign n9597 = ~n16714 | ~P2_REG1_REG_5__SCAN_IN;
  assign n11132 = ~n9599 | ~n8943;
  assign n9600 = ~n16774 | ~n16775;
  assign n16696 = ~n9601 | ~n11126;
  assign n9601 = ~n16676 | ~P2_REG1_REG_3__SCAN_IN;
  assign n9602 = ~P2_REG1_REG_3__SCAN_IN;
  assign n9604 = ~n16805 | ~n16804;
  assign n16821 = ~n11077;
  assign n9607 = ~n9609;
  assign n9609 = n11044 & n17330;
  assign n16683 = ~n11043 & ~n9609;
  assign n9614 = ~n9612 | ~n9610;
  assign n9612 = ~n16751 | ~n9616;
  assign n9613 = n16751 | n11193;
  assign n9621 = ~n12682 | ~n9004;
  assign n9624 = ~n10979 | ~n10980;
  assign n9626 = ~n12723 | ~n9629;
  assign n16639 = ~n9633 | ~n9632;
  assign n9632 = ~P2_REG2_REG_1__SCAN_IN;
  assign n9634 = n16861 | n11234;
  assign n9636 = ~n9638 | ~P2_REG2_REG_13__SCAN_IN;
  assign n9637 = ~n11092 | ~n9638;
  assign n9641 = ~n9643 | ~n9642;
  assign n9644 = ~n9005 | ~n12757;
  assign n9651 = ~n9647 | ~n9653;
  assign n16741 = n9648 & n11056;
  assign n9648 = ~n9653 | ~n11055;
  assign n9650 = ~n11056;
  assign n16718 = ~n11055 | ~n11056;
  assign n11118 = ~n9654 ^ n11281;
  assign n9654 = ~n9656 | ~n9655;
  assign n9656 = ~n11113 | ~n9659;
  assign n9659 = ~n11898;
  assign n12675 = ~n9661 | ~n9660;
  assign n9661 = ~n9662 | ~n12641;
  assign n9662 = ~n12632 | ~n12633;
  assign n14837 = ~n9667 | ~n13327;
  assign n9667 = n14863 | n14861;
  assign n9678 = ~n13419;
  assign n9674 = ~n9676 | ~n13281;
  assign n15644 = ~n9675 | ~n13423;
  assign n9675 = ~n9025 | ~n13419;
  assign n9677 = ~n9678 | ~n13423;
  assign n9679 = ~n11973 | ~n11972;
  assign n15710 = ~n9679 ^ n15709;
  assign n14742 = ~n11981 | ~n13336;
  assign n9682 = ~n9683 | ~n15344;
  assign n9683 = ~n15346 | ~n15345;
  assign n9687 = ~n9963 | ~n9964;
  assign n11298 = ~n9963 | ~n9964;
  assign n10145 = ~n9689 | ~n9000;
  assign n14468 = ~n14467 | ~n14466;
  assign n14556 = ~n9700 | ~n9704;
  assign n9700 = ~n9707 | ~n10315;
  assign n9701 = ~n9704 | ~n9702;
  assign n9703 = ~n14395 | ~n9704;
  assign n14447 = ~n14395 | ~n10282;
  assign n9705 = ~n10315 | ~n9706;
  assign n10189 = ~n10500 | ~n8885;
  assign n11721 = ~n9708 | ~n9710;
  assign n13586 = ~n9711 | ~n12173;
  assign n9711 = ~n12164 | ~n9716;
  assign n9712 = ~n9713 & ~n9008;
  assign n9715 = ~n12164;
  assign n10990 = ~n9719 | ~n9722;
  assign n10968 = ~n9719 | ~n9718;
  assign n9723 = ~n13518 | ~n9725;
  assign n9733 = ~n12226 | ~n9808;
  assign n9729 = ~n9808;
  assign n9730 = ~n9007 & ~n9731;
  assign n13547 = ~n9733 | ~n12228;
  assign n11728 = ~n9739 | ~n11368;
  assign n11730 = ~n9739 | ~n9737;
  assign n9739 = ~n9740 | ~n17214;
  assign n9740 = ~n11323 ^ P2_B_REG_SCAN_IN;
  assign n9741 = n13154 & n9745;
  assign n9744 = ~n13154;
  assign n13221 = ~n9747 | ~n9746;
  assign n9749 = ~n13205;
  assign n9750 = ~n13205 | ~n8942;
  assign n9752 = ~n8900 | ~n9756;
  assign n9754 = ~n16421 | ~n9301;
  assign n9755 = ~n13254 | ~n9756;
  assign n9757 = ~n13375 | ~n9760;
  assign n10262 = ~n9762 | ~n10227;
  assign n9762 = ~n10226 | ~n10225;
  assign n10001 = ~n9971 | ~n9764;
  assign n10476 = ~n9766;
  assign n12213 = ~n10593 ^ n10592;
  assign n9769 = ~n9869 | ~n9803;
  assign n9768 = n9016 & n9803;
  assign n9870 = ~n9769 | ~P1_IR_REG_31__SCAN_IN;
  assign n11935 = ~n9770 | ~n9772;
  assign n9770 = ~n11931 | ~n9774;
  assign n14981 = ~n11931 | ~n11930;
  assign n9777 = ~n14994;
  assign n14860 = ~n9778 | ~n11942;
  assign n9778 = ~n14887 | ~n11941;
  assign n9780 = ~n11942 | ~n9781;
  assign n9781 = ~n11941;
  assign n15793 = ~n9785;
  assign n15758 = ~n15793 & ~n11918;
  assign n9849 = ~n9848 | ~n9828;
  assign n9789 = ~P1_IR_REG_25__SCAN_IN;
  assign n9790 = ~n14741 | ~n9791;
  assign n9799 = ~n15709;
  assign n9797 = ~n9798;
  assign n12311 = ~n10842 ^ n10840;
  assign n10823 = n12311 | n10128;
  assign n9800 = ~n17238 & ~n17232;
  assign n9801 = n13992 & n12732;
  assign n9803 = n9871 & n9874;
  assign n9804 = n12890 & n8890;
  assign n9805 = n11295 & n13535;
  assign n9806 = ~n12083 & ~n16528;
  assign n9807 = n10681 & n10680;
  assign n9808 = ~n13621 | ~n17516;
  assign n11081 = ~n11079 | ~n9816;
  assign n13390 = n15930 | n11910;
  assign n9809 = ~n12720 | ~n14017;
  assign n9810 = ~n14269 & ~n14280;
  assign n9811 = n10954 & n10953;
  assign n9812 = ~n9938 | ~SI_1_;
  assign n9813 = n12475 & n12781;
  assign n9815 = ~n14743 & ~n13459;
  assign n9816 = n11217 | n11078;
  assign n9817 = ~n14428 & ~n10644;
  assign n13459 = ~n13346;
  assign n11923 = ~n15659 | ~n14559;
  assign n11943 = ~n14876 | ~n14891;
  assign n10322 = n10321 & n10320;
  assign n11948 = ~n14822 | ~n14839;
  assign n10433 = ~n10391 | ~n10390;
  assign n10325 = n10324 & n10323;
  assign n11017 = n11016 | P2_IR_REG_27__SCAN_IN;
  assign n12086 = ~n9806 & ~n8932;
  assign n11185 = ~n16722 & ~n16723;
  assign n12233 = ~P2_REG3_REG_20__SCAN_IN;
  assign n12438 = ~n17168;
  assign n12887 = n9800;
  assign n17172 = ~n17356;
  assign n12398 = ~n16418;
  assign n10705 = n10666 & P1_REG3_REG_21__SCAN_IN;
  assign n10564 = n10540 & P1_REG3_REG_17__SCAN_IN;
  assign n9827 = ~P1_IR_REG_12__SCAN_IN;
  assign n15178 = ~n15024;
  assign n12012 = n10902 & n16166;
  assign n10717 = n10693 & n10692;
  assign n10528 = n10526 & n10525;
  assign n13638 = n12138 | n16507;
  assign n16539 = ~n16458 | ~n12070;
  assign n12221 = ~n12234;
  assign n13932 = ~n17516;
  assign n12969 = ~n14022 | ~n12968;
  assign n16993 = ~n14092 | ~n14091;
  assign n17083 = n17205 | n12555;
  assign n17373 = ~n16590;
  assign n17356 = n12489 & n12488;
  assign n14972 = ~n16388;
  assign n14622 = ~n16409;
  assign n14891 = ~n16397;
  assign n14625 = ~n16415;
  assign n14679 = n14677 | n14676;
  assign n10108 = ~n10053 | ~P1_REG3_REG_3__SCAN_IN;
  assign n16170 = n11988 & n11987;
  assign n10156 = ~n10153 | ~n10152;
  assign n16605 = ~n16542;
  assign n17185 = ~n17147;
  assign n13719 = ~n17551;
  assign n10918 = n10838 | n10837;
  assign n10761 = n17213 | n8878;
  assign n10268 = n10200 & n10175;
  assign n10612 = n10615 & n10530;
  assign n16616 = ~n13693;
  assign n16542 = n12335 | n12544;
  assign n13625 = ~n14221;
  assign n16573 = ~n16989;
  assign n16618 = ~n16577;
  assign n13951 = n11596 & n11595;
  assign n16949 = n11294 & n11293;
  assign n17396 = ~n16522;
  assign n11772 = n10989 | n17214;
  assign n15311 = n10933 | n11302;
  assign n12394 = ~n12389 & ~n12388;
  assign n11837 = ~P1_ADDR_REG_1__SCAN_IN;
  assign n16577 = n11780 | n11779;
  assign n16595 = ~n16610;
  assign n17551 = n12885 | n12884;
  assign n14097 = ~n17128;
  assign n17349 = n11763 & n11762;
  assign n15361 = ~n15333;
  assign n15376 = ~n15293;
  assign n16418 = n10858 | n10857;
  assign n16397 = n10632 | n10631;
  assign n15640 = ~n15012;
  assign n15896 = n16004 & n15853;
  assign n15991 = n16004 & n13010;
  assign n11847 = ~n17564 & ~n17563;
  assign n11853 = ~n17558 & ~n17557;
  assign n10956 = n10955 & n9811;
  assign n17564 = ~n11846 & ~n11845;
  assign n17600 = ~n17602 & ~n11856;
  assign n9821 = ~n9820 | ~n9819;
  assign n9826 = ~n9823 | ~n9822;
  assign n9825 = ~n10168 | ~n9824;
  assign n9829 = ~P1_IR_REG_15__SCAN_IN & ~P1_IR_REG_14__SCAN_IN;
  assign n10446 = ~n8905 | ~n9829;
  assign n9830 = ~P1_IR_REG_17__SCAN_IN;
  assign n9831 = ~n10483 | ~n9830;
  assign n10556 = ~P1_IR_REG_18__SCAN_IN;
  assign n9832 = ~n10557 | ~n10556;
  assign n11959 = ~n9833 ^ P1_IR_REG_19__SCAN_IN;
  assign n9836 = ~P1_IR_REG_14__SCAN_IN & ~P1_IR_REG_18__SCAN_IN;
  assign n9845 = ~n9837 | ~n9836;
  assign n9838 = ~n9845;
  assign n9839 = ~n9858 | ~P1_IR_REG_31__SCAN_IN;
  assign n9841 = ~n9840 | ~P1_IR_REG_31__SCAN_IN;
  assign n14848 = ~n11959 | ~n9914;
  assign n9842 = ~P1_IR_REG_13__SCAN_IN & ~P1_IR_REG_24__SCAN_IN;
  assign n9844 = n9842 & n9827;
  assign n9846 = ~n9844 | ~n9843;
  assign n11802 = ~n9872 ^ P1_IR_REG_26__SCAN_IN;
  assign n9850 = ~n9849 | ~P1_IR_REG_31__SCAN_IN;
  assign n16009 = ~n9850 ^ P1_IR_REG_25__SCAN_IN;
  assign n9857 = n11802 & n16009;
  assign n9853 = ~n9852 | ~n9851;
  assign n9854 = ~n9845 & ~n9853;
  assign n9855 = ~n8905 | ~n9854;
  assign n9856 = ~n9855 | ~P1_IR_REG_31__SCAN_IN;
  assign n16015 = ~n9856 ^ P1_IR_REG_24__SCAN_IN;
  assign n11296 = ~n9857 | ~n16015;
  assign n9863 = n14848 & n11296;
  assign n13477 = ~n13382;
  assign n9860 = ~n9858;
  assign n9859 = ~P1_IR_REG_21__SCAN_IN;
  assign n9861 = ~n9860 | ~n9859;
  assign n10905 = ~P1_IR_REG_22__SCAN_IN;
  assign n13484 = ~n16029;
  assign n10500 = ~n9862 | ~n9863;
  assign n9864 = ~n9914;
  assign n9866 = ~n9865 | ~n9864;
  assign n13008 = ~n16029 | ~n16034;
  assign n9869 = ~n9868;
  assign n9873 = ~n9872 | ~n9871;
  assign n15386 = ~n9875 ^ n9874;
  assign n9877 = n9876 | n9897;
  assign n16148 = ~n9877 ^ P1_IR_REG_2__SCAN_IN;
  assign n9893 = ~n9976 | ~n16148;
  assign n9883 = ~n9894 | ~P2_DATAO_REG_1__SCAN_IN;
  assign n9885 = ~n8887 | ~P1_DATAO_REG_0__SCAN_IN;
  assign n9884 = ~n9894 | ~P2_DATAO_REG_0__SCAN_IN;
  assign n9887 = ~n9886 | ~n9939;
  assign n9888 = SI_1_ & SI_0_;
  assign n9994 = ~n9939 | ~n9888;
  assign n9889 = ~n9894 | ~P2_DATAO_REG_2__SCAN_IN;
  assign n9891 = ~SI_2_;
  assign n12056 = ~n9973 ^ n9972;
  assign n9892 = n10128 | n12056;
  assign n11909 = n9892 & n9893;
  assign n10164 = ~n10482;
  assign n9895 = ~P2_DATAO_REG_2__SCAN_IN;
  assign n11908 = n10482 | n9895;
  assign n16193 = ~n11909 | ~n11908;
  assign n9916 = ~n10189 | ~n16193;
  assign n9897 = ~P1_IR_REG_31__SCAN_IN;
  assign n15236 = ~n9899;
  assign n9900 = P1_IR_REG_29__SCAN_IN & n9897;
  assign n9904 = ~n9901 & ~n9900;
  assign n9903 = ~n9902 | ~P1_IR_REG_31__SCAN_IN;
  assign n9905 = ~n9904 | ~n9903;
  assign n9909 = ~n8891 | ~P1_REG1_REG_2__SCAN_IN;
  assign n9910 = ~n9906;
  assign n9908 = ~n10054 | ~P1_REG3_REG_2__SCAN_IN;
  assign n9912 = ~n10085 | ~P1_REG2_REG_2__SCAN_IN;
  assign n9911 = ~n10007 | ~P1_REG0_REG_2__SCAN_IN;
  assign n10118 = n9914 & n11296;
  assign n10093 = ~n10545;
  assign n9915 = ~n11910 | ~n10093;
  assign n9917 = ~n9916 | ~n9915;
  assign n9967 = ~n9917 ^ n10861;
  assign n9919 = ~n10864 | ~n11910;
  assign n10013 = ~n10545;
  assign n9918 = ~n16193 | ~n10013;
  assign n9968 = ~n9919 | ~n9918;
  assign n15345 = n9967 | n9968;
  assign n15423 = ~P1_IR_REG_0__SCAN_IN;
  assign n9924 = ~n8894 | ~P1_IR_REG_0__SCAN_IN;
  assign n9922 = ~n11800 | ~SI_0_;
  assign n11316 = ~n9922 ^ P2_DATAO_REG_0__SCAN_IN;
  assign n9923 = ~n9921 | ~n11316;
  assign n9926 = ~n8893 | ~P1_REG1_REG_0__SCAN_IN;
  assign n9925 = ~n10007 | ~P1_REG0_REG_0__SCAN_IN;
  assign n9928 = ~n10085 | ~P1_REG2_REG_0__SCAN_IN;
  assign n9927 = ~n10054 | ~P1_REG3_REG_0__SCAN_IN;
  assign n9929 = ~n9928 | ~n9927;
  assign n15980 = n9930 | n9929;
  assign n9931 = ~n15980 | ~n10118;
  assign n11604 = ~P1_REG1_REG_0__SCAN_IN;
  assign n9935 = ~n10864 | ~n15980;
  assign n9933 = ~n10013 | ~n16173;
  assign n9932 = n11296 | n15423;
  assign n9934 = n9933 & n9932;
  assign n11720 = ~n9935 | ~n9934;
  assign n9937 = ~n11721 | ~n11720;
  assign n9941 = ~n9938 ^ SI_1_;
  assign n9940 = n9939 & SI_0_;
  assign n12043 = ~n9941 ^ n9940;
  assign n17342 = ~n12043;
  assign n9949 = n10128 | n17342;
  assign n9947 = ~n9876;
  assign n9942 = ~P1_IR_REG_1__SCAN_IN;
  assign n9945 = ~n9942 | ~P1_IR_REG_31__SCAN_IN;
  assign n9943 = ~P1_IR_REG_31__SCAN_IN | ~P1_IR_REG_0__SCAN_IN;
  assign n9944 = ~n9943 | ~P1_IR_REG_1__SCAN_IN;
  assign n9946 = ~n9945 | ~n9944;
  assign n16155 = n9947 & n9946;
  assign n9948 = ~n8894 | ~n16155;
  assign n9952 = n9949 & n9948;
  assign n9950 = ~P2_DATAO_REG_1__SCAN_IN;
  assign n9951 = n10482 | n9950;
  assign n9959 = ~n10824 | ~n16182;
  assign n9954 = ~n8897 | ~P1_REG3_REG_1__SCAN_IN;
  assign n9955 = ~n9954 | ~n9953;
  assign n9958 = ~n11906 | ~n10013;
  assign n9960 = ~n9959 | ~n9958;
  assign n9961 = ~n9960 ^ n10803;
  assign n9964 = ~n9961;
  assign n9963 = ~n9962;
  assign n9966 = ~n8876 | ~n9310;
  assign n9965 = ~n16182 | ~n10013;
  assign n11300 = n9966 & n9965;
  assign n9970 = ~n9967;
  assign n9969 = ~n9968;
  assign n9971 = ~n9894 | ~P2_DATAO_REG_3__SCAN_IN;
  assign n9997 = ~n10001 ^ SI_3_;
  assign n9974 = ~P2_DATAO_REG_3__SCAN_IN;
  assign n9975 = ~n9990 | ~P1_IR_REG_31__SCAN_IN;
  assign n16142 = ~n9975 ^ P1_IR_REG_3__SCAN_IN;
  assign n9977 = ~n9976 | ~n16142;
  assign n9985 = ~n10824 | ~n9323;
  assign n9980 = ~n10007 | ~P1_REG0_REG_3__SCAN_IN;
  assign n9978 = ~P1_REG3_REG_3__SCAN_IN;
  assign n9979 = ~n10054 | ~n9978;
  assign n9982 = ~n10085 | ~P1_REG2_REG_3__SCAN_IN;
  assign n9981 = ~n8893 | ~P1_REG1_REG_3__SCAN_IN;
  assign n9984 = ~n11905 | ~n10013;
  assign n9986 = ~n9985 | ~n9984;
  assign n10019 = ~n9986 ^ n10803;
  assign n9988 = ~n8876 | ~n11905;
  assign n9987 = ~n9323 | ~n10013;
  assign n10020 = n9988 & n9987;
  assign n15266 = n10019 | n10020;
  assign n15307 = ~n15268 | ~n15266;
  assign n9989 = ~P2_DATAO_REG_4__SCAN_IN;
  assign n9993 = n8873 | n9989;
  assign n9991 = ~n10030 | ~P1_IR_REG_31__SCAN_IN;
  assign n16136 = ~n9991 ^ P1_IR_REG_4__SCAN_IN;
  assign n9992 = ~n8894 | ~n16136;
  assign n10000 = ~n9996 | ~n9995;
  assign n9999 = ~n9998 & ~n9997;
  assign n10035 = ~n10001 | ~SI_3_;
  assign n10003 = ~n10286 | ~P1_DATAO_REG_4__SCAN_IN;
  assign n10002 = ~n9894 | ~P2_DATAO_REG_4__SCAN_IN;
  assign n10071 = ~n10039 ^ SI_4_;
  assign n10004 = ~n16135;
  assign n10005 = n10004 | n10128;
  assign n10015 = ~n10824 | ~n16216;
  assign n10008 = ~n10007 | ~P1_REG0_REG_4__SCAN_IN;
  assign n10009 = ~P1_REG3_REG_4__SCAN_IN;
  assign n15865 = ~n10009 ^ P1_REG3_REG_3__SCAN_IN;
  assign n10011 = ~n8897 | ~n15865;
  assign n10010 = ~n10085 | ~P1_REG2_REG_4__SCAN_IN;
  assign n10012 = ~n10011 | ~n10010;
  assign n10014 = ~n11903 | ~n10013;
  assign n10016 = ~n10015 | ~n10014;
  assign n10024 = ~n10016 ^ n10803;
  assign n10018 = ~n8876 | ~n11903;
  assign n10017 = ~n16216 | ~n10093;
  assign n10025 = ~n10018 | ~n10017;
  assign n15308 = ~n10024 ^ n10025;
  assign n10022 = ~n10019;
  assign n10021 = ~n10020;
  assign n15306 = n10022 | n10021;
  assign n10023 = n15308 & n15306;
  assign n10028 = ~n15307 | ~n10023;
  assign n10026 = ~n10024;
  assign n10027 = ~n10026 | ~n10025;
  assign n10029 = ~P2_DATAO_REG_6__SCAN_IN;
  assign n10034 = n8873 | n10029;
  assign n10067 = ~n10030 & ~P1_IR_REG_4__SCAN_IN;
  assign n10031 = ~P1_IR_REG_5__SCAN_IN;
  assign n10032 = n10167 | n9897;
  assign n15477 = ~n10032 ^ P1_IR_REG_6__SCAN_IN;
  assign n10033 = ~n9976 | ~n15477;
  assign n10052 = n10034 & n10033;
  assign n10074 = ~n10039 | ~SI_4_;
  assign n10038 = ~n10286 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n10037 = ~n9894 | ~P2_DATAO_REG_5__SCAN_IN;
  assign n10046 = ~n10038 | ~n10037;
  assign n10076 = ~n10046 ^ SI_5_;
  assign n10043 = ~n10076;
  assign n10041 = ~n10039;
  assign n10040 = ~SI_4_;
  assign n10042 = ~n10041 | ~n10040;
  assign n10044 = n10043 & n10042;
  assign n10048 = ~n10045 | ~n10044;
  assign n10047 = ~n10046 | ~SI_5_;
  assign n10050 = ~n10438 | ~P1_DATAO_REG_6__SCAN_IN;
  assign n10051 = ~n10720 | ~n12090;
  assign n10062 = ~n10824 | ~n9550;
  assign n10056 = ~n10007 | ~P1_REG0_REG_6__SCAN_IN;
  assign n15380 = ~n10108 ^ P1_REG3_REG_6__SCAN_IN;
  assign n10055 = ~n10054 | ~n15380;
  assign n10060 = ~n10056 | ~n10055;
  assign n10058 = ~n13264 | ~P1_REG2_REG_6__SCAN_IN;
  assign n10057 = ~n8891 | ~P1_REG1_REG_6__SCAN_IN;
  assign n10059 = ~n10058 | ~n10057;
  assign n10061 = ~n15844 | ~n10093;
  assign n10063 = ~n10062 | ~n10061;
  assign n10099 = ~n10063 ^ n10861;
  assign n10065 = ~n8876 | ~n15844;
  assign n10064 = ~n9550 | ~n10093;
  assign n10100 = ~n10065 | ~n10064;
  assign n15373 = n10099 | n10100;
  assign n10066 = ~P2_DATAO_REG_5__SCAN_IN;
  assign n10070 = n8873 | n10066;
  assign n10068 = n10067 | n9897;
  assign n16128 = ~n10068 ^ P1_IR_REG_5__SCAN_IN;
  assign n10069 = ~n9976 | ~n16128;
  assign n10079 = n10070 & n10069;
  assign n10072 = ~n10071;
  assign n10075 = ~n10073 | ~n10072;
  assign n10077 = ~n10075 | ~n10074;
  assign n16127 = ~n10077 ^ n10076;
  assign n10078 = ~n10720 | ~n16127;
  assign n10091 = ~n10824 | ~n16227;
  assign n10080 = ~n10007 | ~P1_REG0_REG_5__SCAN_IN;
  assign n10089 = ~n10081 | ~n10080;
  assign n10083 = ~P1_REG3_REG_5__SCAN_IN;
  assign n10082 = ~P1_REG3_REG_3__SCAN_IN | ~P1_REG3_REG_4__SCAN_IN;
  assign n10084 = ~n10083 | ~n10082;
  assign n15858 = n10108 & n10084;
  assign n10087 = ~n10054 | ~n15858;
  assign n10086 = ~n10085 | ~P1_REG2_REG_5__SCAN_IN;
  assign n10088 = ~n10087 | ~n10086;
  assign n10090 = ~n15876 | ~n10093;
  assign n10092 = ~n10091 | ~n10090;
  assign n15368 = ~n10092 ^ n10861;
  assign n10095 = ~n8876 | ~n15876;
  assign n10094 = ~n16227 | ~n10093;
  assign n15366 = ~n10095 | ~n10094;
  assign n10096 = n15368 | n15366;
  assign n10097 = n15373 & n10096;
  assign n10098 = n15368 & n15366;
  assign n10103 = ~n10098 | ~n15373;
  assign n10102 = ~n10099;
  assign n10101 = ~n10100;
  assign n15372 = n10102 | n10101;
  assign n10104 = n10103 & n15372;
  assign n10105 = ~n10007 | ~P1_REG0_REG_7__SCAN_IN;
  assign n10117 = n10106 & n10105;
  assign n10107 = ~P1_REG3_REG_6__SCAN_IN | ~P1_REG3_REG_7__SCAN_IN;
  assign n10113 = ~n10200;
  assign n10109 = ~n10108;
  assign n10111 = ~n10109 | ~P1_REG3_REG_6__SCAN_IN;
  assign n10110 = ~P1_REG3_REG_7__SCAN_IN;
  assign n10112 = ~n10111 | ~n10110;
  assign n15781 = n10113 & n10112;
  assign n10115 = ~n10054 | ~n15781;
  assign n10114 = ~n13264 | ~P1_REG2_REG_7__SCAN_IN;
  assign n10116 = n10115 & n10114;
  assign n10138 = n11964 | n10863;
  assign n10122 = ~n10121 | ~SI_6_;
  assign n10147 = ~n10123 | ~n10122;
  assign n10126 = ~n13271 | ~P1_DATAO_REG_7__SCAN_IN;
  assign n10127 = ~SI_7_;
  assign n17312 = ~n10147 ^ n10146;
  assign n10136 = n17312 | n8880;
  assign n10129 = ~P2_DATAO_REG_7__SCAN_IN;
  assign n10134 = n8873 | n10129;
  assign n10130 = ~P1_IR_REG_6__SCAN_IN;
  assign n10131 = ~n10167 | ~n10130;
  assign n10132 = ~n10131 | ~P1_IR_REG_31__SCAN_IN;
  assign n11672 = ~n10132 ^ P1_IR_REG_7__SCAN_IN;
  assign n10133 = ~n9976 | ~n11672;
  assign n10135 = n10134 & n10133;
  assign n10137 = ~n10824 | ~n11963;
  assign n10139 = ~n10138 | ~n10137;
  assign n10144 = ~n10139 ^ n10861;
  assign n10141 = n10500 | n11964;
  assign n10140 = ~n11963 | ~n10118;
  assign n10143 = ~n10141 | ~n10140;
  assign n15251 = n10144 & n10143;
  assign n10142 = ~n15251;
  assign n15250 = n10144 | n10143;
  assign n15284 = ~n10145 | ~n15250;
  assign n10149 = ~n10148 | ~SI_7_;
  assign n10151 = ~n13271 | ~P1_DATAO_REG_8__SCAN_IN;
  assign n10152 = ~SI_8_;
  assign n10154 = ~n10153;
  assign n10155 = ~n10154 | ~SI_8_;
  assign n10159 = ~n13271 | ~P1_DATAO_REG_9__SCAN_IN;
  assign n10158 = ~n12871 | ~P2_DATAO_REG_9__SCAN_IN;
  assign n10160 = ~SI_9_;
  assign n10162 = ~n10161;
  assign n10163 = ~n10162 | ~SI_9_;
  assign n17300 = ~n10226 ^ n10224;
  assign n10173 = n17300 | n8880;
  assign n10193 = ~n10164;
  assign n10165 = ~P2_DATAO_REG_9__SCAN_IN;
  assign n10171 = n8873 | n10165;
  assign n10166 = ~P1_IR_REG_7__SCAN_IN & ~P1_IR_REG_6__SCAN_IN;
  assign n10236 = ~n10194 | ~n10168;
  assign n10169 = ~n10236 | ~P1_IR_REG_31__SCAN_IN;
  assign n11717 = ~n10169 ^ P1_IR_REG_9__SCAN_IN;
  assign n10170 = ~n9976 | ~n11717;
  assign n10172 = n10171 & n10170;
  assign n10185 = ~n15737 | ~n10824;
  assign n10179 = ~n13263 | ~P1_REG0_REG_9__SCAN_IN;
  assign n10174 = ~n10200 | ~P1_REG3_REG_8__SCAN_IN;
  assign n11711 = ~P1_REG3_REG_9__SCAN_IN;
  assign n10176 = n10174 & n11711;
  assign n10175 = P1_REG3_REG_9__SCAN_IN & P1_REG3_REG_8__SCAN_IN;
  assign n15741 = n10176 | n10268;
  assign n10177 = ~n15741;
  assign n10178 = ~n10054 | ~n10177;
  assign n10183 = ~n10179 | ~n10178;
  assign n10181 = ~n13264 | ~P1_REG2_REG_9__SCAN_IN;
  assign n10180 = ~n8892 | ~P1_REG1_REG_9__SCAN_IN;
  assign n10182 = ~n10181 | ~n10180;
  assign n15771 = n10183 | n10182;
  assign n10184 = ~n15771 | ~n10118;
  assign n10186 = ~n10185 | ~n10184;
  assign n15328 = ~n10186 ^ n10803;
  assign n10188 = ~n15737 | ~n10118;
  assign n10187 = ~n8876 | ~n15771;
  assign n10216 = n10188 & n10187;
  assign n10214 = n15328 | n10216;
  assign n17306 = ~n10191 ^ n10190;
  assign n10192 = ~P2_DATAO_REG_8__SCAN_IN;
  assign n10197 = n8873 | n10192;
  assign n10195 = n10194 | n9897;
  assign n11699 = ~n10195 ^ P1_IR_REG_8__SCAN_IN;
  assign n10196 = ~n9976 | ~n11699;
  assign n10198 = n10197 & n10196;
  assign n10209 = ~n10824 | ~n16258;
  assign n10203 = ~n10007 | ~P1_REG0_REG_8__SCAN_IN;
  assign n15754 = ~n10200 ^ P1_REG3_REG_8__SCAN_IN;
  assign n10201 = ~n15754;
  assign n10202 = ~n10054 | ~n10201;
  assign n10207 = ~n10203 | ~n10202;
  assign n10205 = ~n13264 | ~P1_REG2_REG_8__SCAN_IN;
  assign n10206 = ~n10205 | ~n10204;
  assign n10208 = ~n15729 | ~n10013;
  assign n10210 = ~n10209 | ~n10208;
  assign n15324 = ~n10210 ^ n10803;
  assign n10212 = ~n8876 | ~n15729;
  assign n10211 = ~n16258 | ~n10118;
  assign n15322 = n10212 & n10211;
  assign n10213 = n15324 | n15322;
  assign n10215 = n10214 & n10213;
  assign n10223 = ~n15284 | ~n10215;
  assign n15285 = ~n15324;
  assign n15286 = ~n15322;
  assign n10217 = n15285 | n15286;
  assign n15327 = ~n10216;
  assign n10218 = ~n10217 | ~n15327;
  assign n10221 = ~n15328 | ~n10218;
  assign n10219 = ~n15327 & ~n15286;
  assign n10220 = ~n10219 | ~n15324;
  assign n10222 = n10221 & n10220;
  assign n14395 = n10223 & n10222;
  assign n10229 = ~n13271 | ~P1_DATAO_REG_10__SCAN_IN;
  assign n10228 = ~n12871 | ~P2_DATAO_REG_10__SCAN_IN;
  assign n10320 = ~n10230 | ~SI_10_;
  assign n10232 = ~n13271 | ~P1_DATAO_REG_11__SCAN_IN;
  assign n10231 = ~n11800 | ~P2_DATAO_REG_11__SCAN_IN;
  assign n10233 = ~SI_11_;
  assign n10323 = ~n10234 | ~n10233;
  assign n10235 = ~n10234;
  assign n10321 = ~n10235 | ~SI_11_;
  assign n10284 = ~n10323 | ~n10321;
  assign n10245 = ~n16094 | ~n10720;
  assign n10264 = ~n10237 | ~P1_IR_REG_31__SCAN_IN;
  assign n10238 = ~P1_IR_REG_10__SCAN_IN;
  assign n10239 = ~n10264 | ~n10238;
  assign n10240 = ~n10239 | ~P1_IR_REG_31__SCAN_IN;
  assign n16095 = ~n10240 ^ P1_IR_REG_11__SCAN_IN;
  assign n10243 = ~n16095 | ~n9976;
  assign n10241 = ~P2_DATAO_REG_11__SCAN_IN;
  assign n10242 = n10193 | n10241;
  assign n10244 = n10243 & n10242;
  assign n10850 = ~n10824;
  assign n10251 = ~n10007 | ~P1_REG0_REG_11__SCAN_IN;
  assign n10246 = ~n10268 | ~P1_REG3_REG_10__SCAN_IN;
  assign n14597 = ~P1_REG3_REG_11__SCAN_IN;
  assign n10248 = n10246 & n14597;
  assign n10247 = P1_REG3_REG_11__SCAN_IN & P1_REG3_REG_10__SCAN_IN;
  assign n15691 = n10248 | n10341;
  assign n10249 = ~n15691;
  assign n10250 = ~n10054 | ~n10249;
  assign n10255 = n10251 & n10250;
  assign n10253 = ~n13264 | ~P1_REG2_REG_11__SCAN_IN;
  assign n10252 = ~n8891 | ~P1_REG1_REG_11__SCAN_IN;
  assign n10254 = n10253 & n10252;
  assign n10256 = n14457 | n10863;
  assign n10258 = ~n10257 | ~n10256;
  assign n10309 = ~n10258 ^ n10803;
  assign n10260 = n16292 | n10863;
  assign n10259 = n10500 | n14457;
  assign n10310 = n10260 & n10259;
  assign n14591 = ~n10309 | ~n10310;
  assign n10263 = ~P2_DATAO_REG_10__SCAN_IN;
  assign n10266 = n10193 | n10263;
  assign n16101 = ~n10264 ^ P1_IR_REG_10__SCAN_IN;
  assign n10265 = ~n9976 | ~n16101;
  assign n10267 = n10266 & n10265;
  assign n10271 = ~n13263 | ~P1_REG0_REG_10__SCAN_IN;
  assign n15705 = ~n10268 ^ P1_REG3_REG_10__SCAN_IN;
  assign n10269 = ~n15705;
  assign n10270 = ~n10054 | ~n10269;
  assign n10275 = ~n10271 | ~n10270;
  assign n10273 = ~n13264 | ~P1_REG2_REG_10__SCAN_IN;
  assign n10272 = ~n8891 | ~P1_REG1_REG_10__SCAN_IN;
  assign n10274 = ~n10273 | ~n10272;
  assign n10276 = ~n15734 | ~n10093;
  assign n10278 = ~n10277 | ~n10276;
  assign n10280 = ~n13105 & ~n10863;
  assign n10279 = n8876 & n15734;
  assign n14585 = n10280 | n10279;
  assign n10281 = n14587 | n14585;
  assign n10282 = n14591 & n10281;
  assign n10290 = ~n10285 | ~n10323;
  assign n10288 = ~n13271 | ~P1_DATAO_REG_12__SCAN_IN;
  assign n10287 = ~n11800 | ~P2_DATAO_REG_12__SCAN_IN;
  assign n10327 = ~n10288 | ~n10287;
  assign n10289 = ~SI_12_;
  assign n10324 = ~n10327 ^ n10289;
  assign n10297 = ~n16087 | ~n10720;
  assign n10291 = ~P2_DATAO_REG_12__SCAN_IN;
  assign n10295 = n10193 | n10291;
  assign n10293 = ~n10292 | ~P1_IR_REG_31__SCAN_IN;
  assign n16088 = ~n10293 ^ P1_IR_REG_12__SCAN_IN;
  assign n10294 = ~n9976 | ~n16088;
  assign n10296 = n10295 & n10294;
  assign n10299 = ~n13263 | ~P1_REG0_REG_12__SCAN_IN;
  assign n15656 = ~n10341 ^ P1_REG3_REG_12__SCAN_IN;
  assign n14454 = ~n15656;
  assign n10298 = ~n10054 | ~n14454;
  assign n10303 = n10299 & n10298;
  assign n10301 = ~n13264 | ~P1_REG2_REG_12__SCAN_IN;
  assign n10300 = ~n8893 | ~P1_REG1_REG_12__SCAN_IN;
  assign n10302 = n10301 & n10300;
  assign n10304 = n14559 | n10863;
  assign n10316 = ~n10305 ^ n10861;
  assign n10307 = n15659 | n10863;
  assign n10306 = n10500 | n14559;
  assign n10317 = ~n10307 | ~n10306;
  assign n10314 = ~n14449;
  assign n10308 = n14587 & n14585;
  assign n10313 = ~n14591 | ~n10308;
  assign n10312 = ~n10309;
  assign n10311 = ~n10310;
  assign n14590 = ~n10312 | ~n10311;
  assign n10319 = ~n10316;
  assign n10318 = ~n10317;
  assign n14448 = ~n10319 | ~n10318;
  assign n10419 = ~n10327 | ~SI_12_;
  assign n10329 = ~n13271 | ~P1_DATAO_REG_13__SCAN_IN;
  assign n10328 = ~n12871 | ~P2_DATAO_REG_13__SCAN_IN;
  assign n10362 = ~n10329 | ~n10328;
  assign n10359 = ~SI_13_;
  assign n10330 = ~n10362 ^ n10359;
  assign n17276 = ~n10361 ^ n10330;
  assign n10331 = ~P2_DATAO_REG_13__SCAN_IN;
  assign n10335 = n10482 | n10331;
  assign n10333 = ~n10332 | ~P1_IR_REG_31__SCAN_IN;
  assign n16081 = ~n10333 ^ P1_IR_REG_13__SCAN_IN;
  assign n10334 = ~n9976 | ~n16081;
  assign n10336 = n10335 & n10334;
  assign n10350 = ~n16315 | ~n10824;
  assign n10344 = ~n13263 | ~P1_REG0_REG_13__SCAN_IN;
  assign n10339 = ~n10341 | ~P1_REG3_REG_12__SCAN_IN;
  assign n10338 = ~P1_REG3_REG_13__SCAN_IN;
  assign n10342 = ~n10339 | ~n10338;
  assign n10340 = P1_REG3_REG_13__SCAN_IN & P1_REG3_REG_12__SCAN_IN;
  assign n15634 = ~n10342 | ~n10408;
  assign n14558 = ~n15634;
  assign n10343 = ~n10054 | ~n14558;
  assign n10348 = n10344 & n10343;
  assign n10346 = ~n13264 | ~P1_REG2_REG_13__SCAN_IN;
  assign n10345 = ~n8892 | ~P1_REG1_REG_13__SCAN_IN;
  assign n10347 = n10346 & n10345;
  assign n10349 = n14455 | n10863;
  assign n10351 = ~n10350 | ~n10349;
  assign n10354 = ~n10351 ^ n10803;
  assign n10353 = ~n16315 | ~n10118;
  assign n10352 = n10500 | n14455;
  assign n10355 = n10353 & n10352;
  assign n14554 = n10354 | n10355;
  assign n10357 = ~n10354;
  assign n10356 = ~n10355;
  assign n10360 = ~n10362;
  assign n10426 = ~n10360 | ~n10359;
  assign n10420 = ~n10362 | ~SI_13_;
  assign n10364 = ~n13271 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n10363 = ~n12871 | ~P2_DATAO_REG_14__SCAN_IN;
  assign n10430 = ~n10364 | ~n10363;
  assign n10423 = ~SI_14_;
  assign n10365 = ~n10430 ^ n10423;
  assign n12157 = ~n10387 ^ n10365;
  assign n10366 = ~P2_DATAO_REG_14__SCAN_IN;
  assign n10368 = n10482 | n10366;
  assign n10395 = n8905 | n9897;
  assign n16075 = ~n10395 ^ P1_IR_REG_14__SCAN_IN;
  assign n10367 = ~n9976 | ~n16075;
  assign n10369 = n10368 & n10367;
  assign n10378 = ~n9555 | ~n10189;
  assign n10372 = ~n13263 | ~P1_REG0_REG_14__SCAN_IN;
  assign n10404 = ~P1_REG3_REG_14__SCAN_IN;
  assign n15610 = ~n10408 ^ n10404;
  assign n14372 = ~n15610;
  assign n10371 = ~n10054 | ~n14372;
  assign n10376 = n10372 & n10371;
  assign n10374 = ~n13264 | ~P1_REG2_REG_14__SCAN_IN;
  assign n10373 = ~n8891 | ~P1_REG1_REG_14__SCAN_IN;
  assign n10375 = n10374 & n10373;
  assign n10377 = n15012 | n10863;
  assign n10379 = ~n10378 | ~n10377;
  assign n10383 = ~n10379 ^ n10803;
  assign n14367 = ~n10382 | ~n10383;
  assign n10381 = ~n11997 & ~n10863;
  assign n10380 = ~n15012 & ~n10500;
  assign n14370 = n10381 | n10380;
  assign n10386 = ~n14367 | ~n14370;
  assign n10385 = ~n10382;
  assign n10384 = ~n10383;
  assign n14368 = ~n10385 | ~n10384;
  assign n10388 = ~n10387 | ~SI_14_;
  assign n10391 = ~n13271 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n10390 = ~n11800 | ~P2_DATAO_REG_15__SCAN_IN;
  assign n10392 = ~n10433 ^ SI_15_;
  assign n10401 = ~n16068 | ~n10720;
  assign n10393 = ~P2_DATAO_REG_15__SCAN_IN;
  assign n10399 = n10193 | n10393;
  assign n10394 = ~P1_IR_REG_14__SCAN_IN;
  assign n10396 = ~n10395 | ~n10394;
  assign n10397 = ~n10396 | ~P1_IR_REG_31__SCAN_IN;
  assign n16069 = ~n10397 ^ P1_IR_REG_15__SCAN_IN;
  assign n10398 = ~n9976 | ~n16069;
  assign n10400 = n10399 & n10398;
  assign n10415 = n15024 | n10850;
  assign n10403 = ~n8892 | ~P1_REG1_REG_15__SCAN_IN;
  assign n10402 = ~n13263 | ~P1_REG0_REG_15__SCAN_IN;
  assign n10413 = n10403 & n10402;
  assign n10406 = n10408 | n10404;
  assign n10405 = ~P1_REG3_REG_15__SCAN_IN;
  assign n10409 = ~n10406 | ~n10405;
  assign n10407 = ~P1_REG3_REG_15__SCAN_IN | ~P1_REG3_REG_14__SCAN_IN;
  assign n15025 = n10409 & n10455;
  assign n10411 = ~n10054 | ~n15025;
  assign n10410 = ~n13264 | ~P1_REG2_REG_15__SCAN_IN;
  assign n10412 = n10411 & n10410;
  assign n10414 = n14997 | n10863;
  assign n10416 = ~n10415 | ~n10414;
  assign n14481 = ~n10416 ^ n10861;
  assign n10418 = n15024 | n10863;
  assign n10417 = n10500 | n14997;
  assign n10507 = ~n10418 | ~n10417;
  assign n10466 = ~n14481 | ~n10507;
  assign n10424 = ~n10430;
  assign n10425 = ~n10424 | ~n10423;
  assign n10427 = ~n10426 | ~n10425;
  assign n10428 = ~n10427 & ~n10429;
  assign n10432 = ~n10429;
  assign n10431 = n10430 & SI_14_;
  assign n10435 = ~n10432 | ~n10431;
  assign n10434 = ~n10433 | ~SI_15_;
  assign n10440 = ~n13271 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n10439 = ~n12871 | ~P2_DATAO_REG_16__SCAN_IN;
  assign n10441 = ~SI_16_;
  assign n10477 = ~n10442 | ~n10441;
  assign n10443 = ~n10442;
  assign n10444 = ~n10443 | ~SI_16_;
  assign n10445 = ~P2_DATAO_REG_16__SCAN_IN;
  assign n10449 = n10482 | n10445;
  assign n10447 = ~n10446 | ~P1_IR_REG_31__SCAN_IN;
  assign n16062 = ~n10447 ^ P1_IR_REG_16__SCAN_IN;
  assign n10448 = ~n9976 | ~n16062;
  assign n10450 = n10449 & n10448;
  assign n10462 = ~n15167 | ~n10824;
  assign n10453 = ~n8893 | ~P1_REG1_REG_16__SCAN_IN;
  assign n10452 = ~n13263 | ~P1_REG0_REG_16__SCAN_IN;
  assign n10460 = ~n10453 | ~n10452;
  assign n10454 = ~P1_REG3_REG_16__SCAN_IN;
  assign n10456 = n10455 & n10454;
  assign n14987 = ~n10540 & ~n10456;
  assign n10458 = ~n10054 | ~n14987;
  assign n10457 = ~n13264 | ~P1_REG2_REG_16__SCAN_IN;
  assign n10459 = ~n10458 | ~n10457;
  assign n10461 = ~n13151 | ~n10118;
  assign n10463 = ~n10462 | ~n10461;
  assign n10503 = ~n10463 ^ n10803;
  assign n10465 = ~n15167 | ~n10118;
  assign n10464 = ~n8876 | ~n13151;
  assign n10504 = n10465 & n10464;
  assign n14486 = n10503 | n10504;
  assign n10467 = n10466 & n14486;
  assign n10512 = ~n14484 | ~n10467;
  assign n10469 = ~n13271 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n10468 = ~n12871 | ~P2_DATAO_REG_17__SCAN_IN;
  assign n10470 = ~SI_17_;
  assign n10519 = ~n10471 | ~n10470;
  assign n10472 = ~n10471;
  assign n10473 = ~n10472 | ~SI_17_;
  assign n10474 = ~n10479;
  assign n10480 = n10552 & n10520;
  assign n10478 = ~n10476 | ~n10475;
  assign n10489 = ~n16054 | ~n10720;
  assign n10481 = ~P2_DATAO_REG_17__SCAN_IN;
  assign n10487 = n10193 | n10481;
  assign n10484 = ~n10483;
  assign n10485 = ~n10484 | ~P1_IR_REG_31__SCAN_IN;
  assign n16056 = ~n10485 ^ P1_IR_REG_17__SCAN_IN;
  assign n10486 = ~n9976 | ~n16056;
  assign n10488 = n10487 & n10486;
  assign n10498 = ~n15157 | ~n10824;
  assign n10490 = ~P1_REG3_REG_17__SCAN_IN;
  assign n14962 = ~n10540 ^ n10490;
  assign n10492 = ~n10054 | ~n14962;
  assign n10491 = ~n13263 | ~P1_REG0_REG_17__SCAN_IN;
  assign n10496 = n10492 & n10491;
  assign n10494 = ~n13264 | ~P1_REG2_REG_17__SCAN_IN;
  assign n10493 = ~n8893 | ~P1_REG1_REG_17__SCAN_IN;
  assign n10495 = n10494 & n10493;
  assign n10497 = n14998 | n10863;
  assign n10499 = ~n10498 | ~n10497;
  assign n10513 = ~n10499 ^ n10861;
  assign n10502 = ~n14961 & ~n10863;
  assign n10501 = ~n14998 & ~n10500;
  assign n10514 = n10502 | n10501;
  assign n14503 = n10513 | n10514;
  assign n10506 = ~n10503;
  assign n10505 = ~n10504;
  assign n14501 = n10506 | n10505;
  assign n10510 = n14503 & n14501;
  assign n14483 = ~n14481;
  assign n14636 = ~n10507;
  assign n10508 = n14486 & n14636;
  assign n10509 = ~n14483 | ~n10508;
  assign n10511 = n10510 & n10509;
  assign n10516 = ~n10513;
  assign n10515 = ~n10514;
  assign n14504 = n10516 | n10515;
  assign n10518 = ~n10438 | ~P1_DATAO_REG_18__SCAN_IN;
  assign n10517 = ~n11800 | ~P2_DATAO_REG_18__SCAN_IN;
  assign n10523 = ~n10518 | ~n10517;
  assign n10553 = ~n10523 ^ SI_18_;
  assign n10521 = ~n10553;
  assign n10524 = ~n10523 | ~SI_18_;
  assign n10526 = ~n13271 | ~P1_DATAO_REG_19__SCAN_IN;
  assign n10525 = ~n12871 | ~P2_DATAO_REG_19__SCAN_IN;
  assign n10527 = ~SI_19_;
  assign n10615 = ~n10528 | ~n10527;
  assign n10529 = ~n10528;
  assign n10530 = ~n10529 | ~SI_19_;
  assign n17248 = ~n10611 ^ n10612;
  assign n10535 = ~n10531 | ~n9976;
  assign n10532 = ~P2_DATAO_REG_19__SCAN_IN;
  assign n10534 = n10193 | n10532;
  assign n10536 = n10535 & n10534;
  assign n10547 = ~n15135 | ~n10824;
  assign n10539 = ~n8892 | ~P1_REG1_REG_19__SCAN_IN;
  assign n10538 = ~n10007 | ~P1_REG0_REG_19__SCAN_IN;
  assign n10544 = ~n10539 | ~n10538;
  assign n14925 = ~P1_REG3_REG_19__SCAN_IN ^ n10600;
  assign n10542 = ~n10054 | ~n14925;
  assign n10541 = ~n13264 | ~P1_REG2_REG_19__SCAN_IN;
  assign n10543 = ~n10542 | ~n10541;
  assign n10546 = ~n16391 | ~n10118;
  assign n10548 = ~n10547 | ~n10546;
  assign n14413 = ~n10548 ^ n10861;
  assign n10550 = ~n15135 | ~n10013;
  assign n10549 = ~n8876 | ~n16391;
  assign n14412 = ~n10550 | ~n10549;
  assign n14415 = n14413 | n14412;
  assign n10554 = ~n10552 | ~n10551;
  assign n17253 = ~n10554 ^ n10553;
  assign n10555 = ~P2_DATAO_REG_18__SCAN_IN;
  assign n10559 = n10193 | n10555;
  assign n16049 = ~n10557 ^ n10556;
  assign n10558 = n16049 | n9921;
  assign n10560 = n10559 & n10558;
  assign n10571 = n14610 | n10850;
  assign n10563 = ~n8891 | ~P1_REG1_REG_18__SCAN_IN;
  assign n10562 = ~n13263 | ~P1_REG0_REG_18__SCAN_IN;
  assign n10569 = ~n10563 | ~n10562;
  assign n10565 = ~n10564;
  assign n14939 = ~P1_REG3_REG_18__SCAN_IN ^ n10565;
  assign n10567 = ~n10054 | ~n14939;
  assign n10566 = ~n13264 | ~P1_REG2_REG_18__SCAN_IN;
  assign n10568 = ~n10567 | ~n10566;
  assign n10570 = ~n16388 | ~n10118;
  assign n10572 = ~n10571 | ~n10570;
  assign n10577 = ~n10572 ^ n10803;
  assign n10574 = n14610 | n10863;
  assign n10573 = ~n8876 | ~n16388;
  assign n10578 = n10574 & n10573;
  assign n10575 = ~n10577 | ~n10578;
  assign n10576 = n14415 & n10575;
  assign n14408 = ~n10577;
  assign n14607 = ~n10578;
  assign n10580 = ~n14408 | ~n14607;
  assign n10579 = ~n14412;
  assign n10581 = ~n10580 | ~n10579;
  assign n10584 = ~n14413 | ~n10581;
  assign n10582 = n14412 & n14607;
  assign n10583 = ~n10582 | ~n14408;
  assign n10585 = n10584 & n10583;
  assign n10586 = ~n10682 | ~n10612;
  assign n10593 = ~n10586 | ~n10615;
  assign n10588 = ~n10438 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n10587 = ~n12871 | ~P2_DATAO_REG_20__SCAN_IN;
  assign n10589 = ~SI_20_;
  assign n10614 = ~n10590 | ~n10589;
  assign n10591 = ~n10590;
  assign n10613 = ~n10591 | ~SI_20_;
  assign n10592 = ~n10614 | ~n10613;
  assign n10594 = ~P2_DATAO_REG_20__SCAN_IN;
  assign n10595 = n10193 | n10594;
  assign n10607 = ~n15124 | ~n10824;
  assign n10598 = ~n8891 | ~P1_REG1_REG_20__SCAN_IN;
  assign n10597 = ~n13263 | ~P1_REG0_REG_20__SCAN_IN;
  assign n10605 = ~n10598 | ~n10597;
  assign n10599 = ~P1_REG3_REG_19__SCAN_IN;
  assign n10601 = ~n10627;
  assign n14898 = ~P1_REG3_REG_20__SCAN_IN ^ n10601;
  assign n10603 = ~n8897 | ~n14898;
  assign n10602 = ~n13264 | ~P1_REG2_REG_20__SCAN_IN;
  assign n10604 = ~n10603 | ~n10602;
  assign n10606 = ~n16394 | ~n10118;
  assign n10608 = ~n10607 | ~n10606;
  assign n10641 = ~n10608 ^ n10861;
  assign n10610 = ~n15124 | ~n10013;
  assign n10609 = ~n8876 | ~n16394;
  assign n10640 = ~n10610 | ~n10609;
  assign n14428 = n10641 & n10640;
  assign n10618 = ~n10682 | ~n10648;
  assign n10617 = ~n10613;
  assign n10616 = n10615 & n10614;
  assign n10621 = ~n10618 | ~n10652;
  assign n10620 = ~n10438 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n10619 = ~n11800 | ~P2_DATAO_REG_21__SCAN_IN;
  assign n10647 = ~n10620 | ~n10619;
  assign n10650 = ~n10647 ^ SI_21_;
  assign n10622 = ~P2_DATAO_REG_21__SCAN_IN;
  assign n10623 = n10193 | n10622;
  assign n15113 = ~n14876;
  assign n10634 = ~n15113 | ~n10824;
  assign n10626 = ~n8893 | ~P1_REG1_REG_21__SCAN_IN;
  assign n10625 = ~n13263 | ~P1_REG0_REG_21__SCAN_IN;
  assign n10632 = ~n10626 | ~n10625;
  assign n10628 = ~n10666;
  assign n14877 = ~P1_REG3_REG_21__SCAN_IN ^ n10628;
  assign n10630 = ~n8897 | ~n14877;
  assign n10629 = ~n13264 | ~P1_REG2_REG_21__SCAN_IN;
  assign n10631 = ~n10630 | ~n10629;
  assign n10633 = ~n16397 | ~n10118;
  assign n10635 = ~n10634 | ~n10633;
  assign n14432 = ~n10635 ^ n10861;
  assign n10638 = ~n14432;
  assign n10637 = ~n14876 & ~n10863;
  assign n10636 = n8876 & n16397;
  assign n10639 = n10637 | n10636;
  assign n14431 = ~n10639;
  assign n10644 = ~n10638 & ~n14431;
  assign n10642 = n14432 | n10639;
  assign n14430 = n10641 | n10640;
  assign n10643 = n10642 & n14430;
  assign n10645 = n10644 | n10643;
  assign n10649 = ~n10647 | ~SI_21_;
  assign n10654 = ~n10682 | ~n10681;
  assign n10653 = ~n10649;
  assign n10651 = ~n10650;
  assign n10656 = ~n13271 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n10655 = ~n11800 | ~P2_DATAO_REG_22__SCAN_IN;
  assign n10657 = ~SI_22_;
  assign n10686 = ~n10658 | ~n10657;
  assign n10659 = ~n10658;
  assign n10660 = ~n10659 | ~SI_22_;
  assign n10684 = ~n10686 | ~n10660;
  assign n10663 = ~n16028 | ~n10720;
  assign n10661 = ~P2_DATAO_REG_22__SCAN_IN;
  assign n10662 = n10193 | n10661;
  assign n10673 = n9570 | n10850;
  assign n10665 = ~n8892 | ~P1_REG1_REG_22__SCAN_IN;
  assign n10664 = ~n13263 | ~P1_REG0_REG_22__SCAN_IN;
  assign n10671 = ~n10665 | ~n10664;
  assign n10667 = ~n10705;
  assign n14851 = ~P1_REG3_REG_22__SCAN_IN ^ n10667;
  assign n10669 = ~n10054 | ~n14851;
  assign n10668 = ~n13264 | ~P1_REG2_REG_22__SCAN_IN;
  assign n10670 = ~n10669 | ~n10668;
  assign n10672 = ~n16400 | ~n10093;
  assign n10674 = ~n10673 | ~n10672;
  assign n10678 = ~n10674 ^ n10803;
  assign n10676 = n9570 | n10863;
  assign n10675 = ~n8876 | ~n16400;
  assign n14572 = ~n10676 | ~n10675;
  assign n10679 = ~n10678;
  assign n10680 = ~n10684;
  assign n10688 = ~n10438 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n10687 = ~n11800 | ~P2_DATAO_REG_23__SCAN_IN;
  assign n10690 = n10688 & n10687;
  assign n10689 = ~SI_23_;
  assign n10693 = ~n10690 | ~n10689;
  assign n10691 = ~n10690;
  assign n10692 = ~n10691 | ~SI_23_;
  assign n10695 = ~n13271 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n10694 = ~n11800 | ~P2_DATAO_REG_24__SCAN_IN;
  assign n10697 = n10695 & n10694;
  assign n10696 = ~SI_24_;
  assign n10751 = ~n10697 | ~n10696;
  assign n10698 = ~n10697;
  assign n10699 = ~n10698 | ~SI_24_;
  assign n10748 = ~n10751 | ~n10699;
  assign n10700 = ~P2_DATAO_REG_24__SCAN_IN;
  assign n10701 = n10193 | n10700;
  assign n10712 = ~n15082 | ~n10824;
  assign n10704 = ~n8891 | ~P1_REG1_REG_24__SCAN_IN;
  assign n10703 = ~n13263 | ~P1_REG0_REG_24__SCAN_IN;
  assign n10710 = ~n10704 | ~n10703;
  assign n10706 = ~n10764;
  assign n14803 = ~P1_REG3_REG_24__SCAN_IN ^ n10706;
  assign n10708 = ~n10054 | ~n14803;
  assign n10707 = ~n13264 | ~P1_REG2_REG_24__SCAN_IN;
  assign n10709 = ~n10708 | ~n10707;
  assign n10711 = ~n16406 | ~n10013;
  assign n10713 = ~n10712 | ~n10711;
  assign n10741 = ~n10713 ^ n10803;
  assign n10715 = ~n15082 | ~n10118;
  assign n10714 = ~n8876 | ~n16406;
  assign n10742 = n10715 & n10714;
  assign n14524 = n10741 | n10742;
  assign n10719 = ~n9051 | ~n9049;
  assign n16021 = ~n10719 | ~n10718;
  assign n10722 = ~n16021 | ~n10720;
  assign n16022 = ~P2_DATAO_REG_23__SCAN_IN;
  assign n10721 = n10193 | n16022;
  assign n10732 = n14822 | n10850;
  assign n10724 = ~n8893 | ~P1_REG1_REG_23__SCAN_IN;
  assign n10723 = ~n13263 | ~P1_REG0_REG_23__SCAN_IN;
  assign n10730 = ~n10724 | ~n10723;
  assign n10726 = ~n10725;
  assign n14824 = ~P1_REG3_REG_23__SCAN_IN ^ n10726;
  assign n10728 = ~n10054 | ~n14824;
  assign n10727 = ~n13264 | ~P1_REG2_REG_23__SCAN_IN;
  assign n10729 = ~n10728 | ~n10727;
  assign n10731 = ~n16403 | ~n10118;
  assign n10733 = ~n10732 | ~n10731;
  assign n14520 = ~n10733 ^ n10861;
  assign n10735 = n14822 | n10863;
  assign n10734 = ~n8876 | ~n16403;
  assign n14518 = ~n10735 | ~n10734;
  assign n10736 = ~n14520 | ~n14518;
  assign n10737 = n14524 & n10736;
  assign n14517 = ~n14520;
  assign n10739 = ~n14518;
  assign n10740 = n14517 & n10739;
  assign n10745 = ~n14524 | ~n10740;
  assign n10744 = ~n10741;
  assign n10743 = ~n10742;
  assign n14523 = n10744 | n10743;
  assign n10746 = n10745 & n14523;
  assign n10749 = ~n10748;
  assign n10754 = ~n13271 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n10753 = ~n11800 | ~P2_DATAO_REG_25__SCAN_IN;
  assign n10756 = n10754 & n10753;
  assign n10755 = ~SI_25_;
  assign n10784 = ~n10756 | ~n10755;
  assign n10757 = ~n10756;
  assign n10758 = ~n10757 | ~SI_25_;
  assign n10781 = ~n10784 | ~n10758;
  assign n17213 = ~n10783 ^ n10781;
  assign n10759 = ~P2_DATAO_REG_25__SCAN_IN;
  assign n10760 = n10193 | n10759;
  assign n10771 = n14778 | n10850;
  assign n10763 = ~n8892 | ~P1_REG1_REG_25__SCAN_IN;
  assign n10762 = ~n13263 | ~P1_REG0_REG_25__SCAN_IN;
  assign n10769 = ~n10763 | ~n10762;
  assign n10765 = ~n10795;
  assign n14781 = ~P1_REG3_REG_25__SCAN_IN ^ n10765;
  assign n10767 = ~n10054 | ~n14781;
  assign n10766 = ~n13264 | ~P1_REG2_REG_25__SCAN_IN;
  assign n10768 = ~n10767 | ~n10766;
  assign n10770 = ~n16409 | ~n10118;
  assign n10772 = ~n10771 | ~n10770;
  assign n10776 = ~n10772 ^ n10803;
  assign n10774 = n14778 | n10863;
  assign n10773 = ~n8876 | ~n16409;
  assign n10777 = ~n10774 | ~n10773;
  assign n10775 = ~n10777;
  assign n10780 = ~n10776 | ~n10775;
  assign n10778 = ~n10776;
  assign n10779 = ~n10778 | ~n10777;
  assign n14466 = n10780 & n10779;
  assign n10782 = ~n10781;
  assign n10786 = ~n13271 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n10785 = ~n11800 | ~P2_DATAO_REG_26__SCAN_IN;
  assign n10788 = n10786 & n10785;
  assign n10787 = ~SI_26_;
  assign n10814 = ~n10788 | ~n10787;
  assign n10789 = ~n10788;
  assign n10790 = ~n10789 | ~SI_26_;
  assign n10811 = ~n10814 | ~n10790;
  assign n11804 = ~P2_DATAO_REG_26__SCAN_IN;
  assign n10791 = n10193 | n11804;
  assign n10802 = n14756 | n10850;
  assign n10794 = ~n8893 | ~P1_REG1_REG_26__SCAN_IN;
  assign n10793 = ~n13263 | ~P1_REG0_REG_26__SCAN_IN;
  assign n10800 = ~n10794 | ~n10793;
  assign n10796 = ~n10827;
  assign n14757 = ~P1_REG3_REG_26__SCAN_IN ^ n10796;
  assign n10798 = ~n10054 | ~n14757;
  assign n10797 = ~n13264 | ~P1_REG2_REG_26__SCAN_IN;
  assign n10799 = ~n10798 | ~n10797;
  assign n10801 = ~n16412 | ~n10118;
  assign n10804 = ~n10802 | ~n10801;
  assign n10807 = ~n10804 ^ n10803;
  assign n10806 = n14756 | n10863;
  assign n10805 = ~n8876 | ~n16412;
  assign n10808 = ~n10806 | ~n10805;
  assign n14621 = ~n10807 ^ n10808;
  assign n10809 = ~n10807;
  assign n10810 = ~n10809 | ~n10808;
  assign n10812 = ~n10811;
  assign n10817 = ~n10438 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n10816 = ~n11800 | ~P2_DATAO_REG_27__SCAN_IN;
  assign n10819 = n10817 & n10816;
  assign n10818 = ~SI_27_;
  assign n10843 = ~n10819 | ~n10818;
  assign n10820 = ~n10819;
  assign n10821 = ~n10820 | ~SI_27_;
  assign n10840 = ~n10843 | ~n10821;
  assign n11814 = ~P2_DATAO_REG_27__SCAN_IN;
  assign n10822 = n10193 | n11814;
  assign n10833 = ~n15052 | ~n10824;
  assign n10826 = ~n8891 | ~P1_REG1_REG_27__SCAN_IN;
  assign n10825 = ~n13263 | ~P1_REG0_REG_27__SCAN_IN;
  assign n10831 = ~n10826 | ~n10825;
  assign n10853 = ~n10827 | ~P1_REG3_REG_26__SCAN_IN;
  assign n14722 = ~P1_REG3_REG_27__SCAN_IN ^ n10853;
  assign n10829 = ~n10054 | ~n14722;
  assign n10828 = ~n13264 | ~P1_REG2_REG_27__SCAN_IN;
  assign n10830 = ~n10829 | ~n10828;
  assign n10832 = ~n16415 | ~n10118;
  assign n10834 = ~n10833 | ~n10832;
  assign n10838 = ~n10834 ^ n10861;
  assign n10836 = ~n15052 | ~n10118;
  assign n10835 = ~n8876 | ~n16415;
  assign n10837 = ~n10836 | ~n10835;
  assign n10839 = ~n10838 | ~n10837;
  assign n12019 = ~n10918 | ~n10839;
  assign n10841 = ~n10840;
  assign n10845 = ~n13271 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n10844 = ~n11800 | ~P2_DATAO_REG_28__SCAN_IN;
  assign n10846 = ~n10845 | ~n10844;
  assign n11869 = n10846 | SI_28_;
  assign n10847 = ~n10846 | ~SI_28_;
  assign n11866 = ~n11869 | ~n10847;
  assign n11825 = ~P2_DATAO_REG_28__SCAN_IN;
  assign n10848 = n10193 | n11825;
  assign n10860 = n12399 | n10850;
  assign n10852 = ~n8892 | ~P1_REG1_REG_28__SCAN_IN;
  assign n10851 = ~n13263 | ~P1_REG0_REG_28__SCAN_IN;
  assign n10858 = ~n10852 | ~n10851;
  assign n12023 = ~P1_REG3_REG_27__SCAN_IN;
  assign n10936 = ~n10853 & ~n12023;
  assign n10854 = ~n10936;
  assign n12001 = ~P1_REG3_REG_28__SCAN_IN ^ n10854;
  assign n10856 = ~n10054 | ~n12001;
  assign n10855 = ~n13264 | ~P1_REG2_REG_28__SCAN_IN;
  assign n10857 = ~n10856 | ~n10855;
  assign n10859 = ~n16418 | ~n10118;
  assign n10862 = ~n10860 | ~n10859;
  assign n10868 = ~n10862 ^ n10861;
  assign n10866 = n12399 | n10863;
  assign n10865 = ~n8876 | ~n16418;
  assign n10867 = ~n10866 | ~n10865;
  assign n10915 = ~n10868 ^ n10867;
  assign n10920 = ~n10915;
  assign n16174 = ~n13008;
  assign n16329 = n13009 & n16174;
  assign n10927 = n16329 | n13367;
  assign n10912 = ~n10927;
  assign n10869 = n16015 | n16009;
  assign n10871 = ~n10869 | ~P1_B_REG_SCAN_IN;
  assign n10870 = n16015 | P1_B_REG_SCAN_IN;
  assign n10872 = ~n10871 | ~n10870;
  assign n16007 = ~n10872 | ~n11802;
  assign n10878 = ~P1_D_REG_6__SCAN_IN & ~P1_D_REG_7__SCAN_IN;
  assign n10876 = P1_D_REG_8__SCAN_IN | P1_D_REG_9__SCAN_IN;
  assign n10874 = ~P1_D_REG_10__SCAN_IN & ~P1_D_REG_11__SCAN_IN;
  assign n10873 = ~P1_D_REG_12__SCAN_IN & ~P1_D_REG_13__SCAN_IN;
  assign n10875 = ~n10874 | ~n10873;
  assign n10877 = ~n10876 & ~n10875;
  assign n10894 = ~n10878 | ~n10877;
  assign n10880 = ~P1_D_REG_18__SCAN_IN & ~P1_D_REG_19__SCAN_IN;
  assign n10879 = ~P1_D_REG_20__SCAN_IN & ~P1_D_REG_21__SCAN_IN;
  assign n10884 = ~n10880 | ~n10879;
  assign n10882 = ~P1_D_REG_16__SCAN_IN & ~P1_D_REG_14__SCAN_IN;
  assign n10881 = ~P1_D_REG_15__SCAN_IN & ~P1_D_REG_17__SCAN_IN;
  assign n10883 = ~n10882 | ~n10881;
  assign n10892 = ~n10884 & ~n10883;
  assign n10886 = ~P1_D_REG_26__SCAN_IN & ~P1_D_REG_27__SCAN_IN;
  assign n10885 = ~P1_D_REG_28__SCAN_IN & ~P1_D_REG_31__SCAN_IN;
  assign n10890 = ~n10886 | ~n10885;
  assign n10888 = ~P1_D_REG_22__SCAN_IN & ~P1_D_REG_23__SCAN_IN;
  assign n10887 = ~P1_D_REG_24__SCAN_IN & ~P1_D_REG_25__SCAN_IN;
  assign n10889 = ~n10888 | ~n10887;
  assign n10891 = ~n10890 & ~n10889;
  assign n10893 = ~n10892 | ~n10891;
  assign n10899 = ~n10894 & ~n10893;
  assign n10896 = ~P1_D_REG_2__SCAN_IN & ~P1_D_REG_3__SCAN_IN;
  assign n10895 = ~P1_D_REG_4__SCAN_IN & ~P1_D_REG_5__SCAN_IN;
  assign n10897 = ~n10896 | ~n10895;
  assign n10898 = ~P1_D_REG_30__SCAN_IN & ~n10897;
  assign n10900 = ~n10899 | ~n10898;
  assign n10901 = ~P1_D_REG_29__SCAN_IN & ~n10900;
  assign n12010 = ~n16007 & ~n10901;
  assign n10902 = n16007 | P1_D_REG_1__SCAN_IN;
  assign n16166 = n11802 | n16009;
  assign n10903 = n16007 | P1_D_REG_0__SCAN_IN;
  assign n16162 = n16015 | n11802;
  assign n10904 = ~n12012 | ~n12392;
  assign n10934 = n12010 | n10904;
  assign n10907 = ~n10906 | ~n10905;
  assign n10909 = ~n10907 | ~P1_IR_REG_31__SCAN_IN;
  assign n10908 = ~P1_IR_REG_23__SCAN_IN;
  assign n13383 = ~n10909 ^ n10908;
  assign n11600 = n11296 & P1_STATE_REG_SCAN_IN;
  assign n10910 = ~n16008;
  assign n10921 = n10934 | n10910;
  assign n10911 = ~n10921;
  assign n15293 = ~n10912 | ~n10911;
  assign n10913 = ~n10918 | ~n15376;
  assign n10914 = ~n10920 & ~n10913;
  assign n10957 = ~n12021 | ~n10914;
  assign n10916 = ~n10915 & ~n15293;
  assign n10955 = ~n10917 | ~n10916;
  assign n10919 = ~n10918 & ~n15293;
  assign n10954 = ~n10920 | ~n10919;
  assign n15902 = n13008 | n13382;
  assign n10923 = n10921 | n15902;
  assign n10922 = ~n16008 | ~n16034;
  assign n10952 = ~n12399 & ~n15333;
  assign n13479 = ~n13383;
  assign n10924 = ~n11296;
  assign n10926 = ~n13479 & ~n10924;
  assign n10925 = ~n13009 | ~n13367;
  assign n12009 = ~n10926 | ~n10925;
  assign n10928 = ~n10934;
  assign n10929 = ~n10928 & ~n10927;
  assign n11304 = ~n12009 & ~n10929;
  assign n10933 = ~n11304 & ~P1_U3086;
  assign n11958 = n13009 | n11991;
  assign n10930 = ~n11958;
  assign n13483 = ~n10930 | ~n16008;
  assign n10931 = n15902 | P1_U3086;
  assign n10932 = ~n13483 | ~n10931;
  assign n11302 = n10932 & n10934;
  assign n10950 = ~n15311 | ~n12001;
  assign n10946 = ~n13483 & ~n10934;
  assign n15319 = ~n10946 | ~n15431;
  assign n10939 = ~n13263 | ~P1_REG0_REG_29__SCAN_IN;
  assign n13013 = ~n10936 | ~P1_REG3_REG_28__SCAN_IN;
  assign n10937 = ~n13013;
  assign n10938 = ~n8897 | ~n10937;
  assign n10943 = ~n10939 | ~n10938;
  assign n10941 = ~n13264 | ~P1_REG2_REG_29__SCAN_IN;
  assign n10940 = ~n8893 | ~P1_REG1_REG_29__SCAN_IN;
  assign n10942 = ~n10941 | ~n10940;
  assign n16421 = n10943 | n10942;
  assign n10945 = n15319 | n9756;
  assign n10944 = ~P1_REG3_REG_28__SCAN_IN | ~P1_U3086;
  assign n10948 = ~n10945 | ~n10944;
  assign n15426 = ~n15431;
  assign n15332 = ~n10946 | ~n15426;
  assign n10947 = ~n15332 & ~n14625;
  assign n10949 = ~n10948 & ~n10947;
  assign n10951 = ~n10950 | ~n10949;
  assign n10953 = ~n10952 & ~n10951;
  assign P1_U3220 = ~n10957 | ~n10956;
  assign n10958 = ~P2_IR_REG_16__SCAN_IN;
  assign n10959 = ~P2_IR_REG_21__SCAN_IN & ~P2_IR_REG_18__SCAN_IN;
  assign n10960 = ~P2_IR_REG_19__SCAN_IN & ~P2_IR_REG_15__SCAN_IN;
  assign n10972 = ~n10995 | ~n10960;
  assign n11765 = ~P2_IR_REG_20__SCAN_IN;
  assign n11102 = ~P2_IR_REG_14__SCAN_IN;
  assign n10961 = ~n11765 | ~n11102;
  assign n10962 = ~n10972 & ~n10961;
  assign n11007 = ~n10980 | ~n10962;
  assign n10992 = ~n11005 | ~n11004;
  assign n10963 = ~n10992;
  assign n11009 = ~P2_IR_REG_22__SCAN_IN;
  assign n10969 = ~P2_IR_REG_24__SCAN_IN;
  assign n10970 = ~P2_IR_REG_2__SCAN_IN & ~P2_IR_REG_25__SCAN_IN;
  assign n10971 = ~n11023 | ~n10970;
  assign n10974 = ~P2_IR_REG_14__SCAN_IN & ~P2_IR_REG_24__SCAN_IN;
  assign n10975 = ~n10974 | ~n10973;
  assign n10977 = ~n10976 & ~n10975;
  assign n10982 = ~n10981 | ~P2_IR_REG_31__SCAN_IN;
  assign n10984 = ~n10982 | ~P2_IR_REG_26__SCAN_IN;
  assign n10983 = ~n11013 | ~P2_IR_REG_31__SCAN_IN;
  assign n10985 = ~n10984 | ~n10983;
  assign n10989 = n11323 | n11809;
  assign n10986 = ~P2_IR_REG_31__SCAN_IN | ~P2_IR_REG_24__SCAN_IN;
  assign n10988 = ~n10987 | ~n10986;
  assign n10991 = ~n10990 | ~P2_IR_REG_31__SCAN_IN;
  assign n12999 = ~n10991 ^ P2_IR_REG_23__SCAN_IN;
  assign n11289 = ~n11772 & ~n12999;
  assign n10994 = ~n10992 & ~P2_IR_REG_15__SCAN_IN;
  assign n10993 = ~P2_IR_REG_16__SCAN_IN & ~P2_IR_REG_14__SCAN_IN;
  assign n10998 = ~n10994 | ~n10993;
  assign n10997 = ~n10996 | ~n10995;
  assign n10999 = ~n10998 & ~n10997;
  assign n11020 = ~n11072 | ~n10999;
  assign n11000 = ~P2_IR_REG_19__SCAN_IN;
  assign n11002 = ~P2_IR_REG_21__SCAN_IN;
  assign n11074 = ~n11072 | ~n11004;
  assign n11006 = ~n11074;
  assign n11089 = ~n11006 | ~n11005;
  assign n11008 = n11089 | n11007;
  assign n11010 = ~n11008 | ~P2_IR_REG_31__SCAN_IN;
  assign n12892 = n9800;
  assign n11011 = ~n12865 | ~n11772;
  assign n12993 = ~n12999;
  assign n11292 = ~n11011 | ~n12993;
  assign n11012 = ~P2_IR_REG_27__SCAN_IN;
  assign n11015 = ~n11012 | ~P2_IR_REG_31__SCAN_IN;
  assign n11016 = ~n11015;
  assign n12179 = n12051 | n11282;
  assign n11019 = ~n11292 | ~n12179;
  assign P2_U3150 = ~n11019 | ~P2_STATE_REG_SCAN_IN;
  assign n11021 = ~n11020 | ~P2_IR_REG_31__SCAN_IN;
  assign n17254 = ~n11021 ^ n9158;
  assign n11115 = ~n17254 | ~P2_REG2_REG_18__SCAN_IN;
  assign n11265 = ~P2_REG2_REG_17__SCAN_IN;
  assign n11251 = ~P2_REG2_REG_15__SCAN_IN;
  assign n11234 = ~P2_REG2_REG_13__SCAN_IN;
  assign n11022 = ~n11089 | ~P2_IR_REG_31__SCAN_IN;
  assign n11225 = ~n11022 ^ P2_IR_REG_11__SCAN_IN;
  assign n16984 = ~P2_REG2_REG_9__SCAN_IN;
  assign n11027 = ~n11024 | ~P2_IR_REG_2__SCAN_IN;
  assign n11026 = ~n11025 | ~P2_IR_REG_31__SCAN_IN;
  assign n11029 = ~P2_REG2_REG_2__SCAN_IN;
  assign n11030 = ~n11165 | ~n11029;
  assign n11034 = ~n11031 | ~P2_IR_REG_1__SCAN_IN;
  assign n11032 = ~P2_IR_REG_1__SCAN_IN;
  assign n11033 = ~n11032 | ~P2_IR_REG_31__SCAN_IN;
  assign n11036 = ~n11034 | ~n11033;
  assign n11035 = ~n11023;
  assign n16625 = ~n9288;
  assign n11037 = n16625 & P2_REG2_REG_0__SCAN_IN;
  assign n11039 = ~n11023 | ~P2_REG2_REG_0__SCAN_IN;
  assign n11041 = ~n16666 | ~n16665;
  assign n11044 = ~n11041 | ~n11040;
  assign n11042 = ~n11045 | ~P2_IR_REG_31__SCAN_IN;
  assign n12064 = ~n11042 ^ P2_IR_REG_3__SCAN_IN;
  assign n11047 = ~n11051 | ~P2_IR_REG_31__SCAN_IN;
  assign n11046 = ~P2_IR_REG_4__SCAN_IN;
  assign n11049 = ~n12072 | ~P2_REG2_REG_4__SCAN_IN;
  assign n11048 = n12072 | P2_REG2_REG_4__SCAN_IN;
  assign n16694 = n11049 & n11048;
  assign n11054 = ~n11050 | ~n11049;
  assign n11053 = ~n11054;
  assign n11052 = ~n9356 | ~P2_IR_REG_31__SCAN_IN;
  assign n11056 = ~n11054 | ~n17325;
  assign n17070 = ~P2_REG2_REG_5__SCAN_IN;
  assign n11057 = ~P2_IR_REG_5__SCAN_IN;
  assign n11063 = ~n11058 | ~n11057;
  assign n11059 = ~n11063 | ~P2_IR_REG_31__SCAN_IN;
  assign n11062 = ~n11059 | ~P2_IR_REG_6__SCAN_IN;
  assign n11060 = ~P2_IR_REG_6__SCAN_IN;
  assign n11061 = ~n11060 | ~P2_IR_REG_31__SCAN_IN;
  assign n11064 = ~n11062 | ~n11061;
  assign n16731 = ~n17319;
  assign n11186 = ~P2_REG2_REG_6__SCAN_IN;
  assign n11065 = ~n16731 | ~n11186;
  assign n11066 = ~n17319 | ~P2_REG2_REG_6__SCAN_IN;
  assign n16740 = ~n11065 | ~n11066;
  assign n11067 = ~n11068 | ~P2_IR_REG_31__SCAN_IN;
  assign n11197 = ~n11067 ^ P2_IR_REG_7__SCAN_IN;
  assign n11193 = ~P2_REG2_REG_7__SCAN_IN;
  assign n17022 = ~P2_REG2_REG_8__SCAN_IN;
  assign n11070 = ~n11069 | ~P2_IR_REG_31__SCAN_IN;
  assign n16777 = n17022 ^ n17307;
  assign n11073 = n11072 | n11071;
  assign n11211 = ~n11073 ^ P2_IR_REG_9__SCAN_IN;
  assign n11078 = ~P2_REG2_REG_10__SCAN_IN;
  assign n11075 = ~n11074 | ~P2_IR_REG_31__SCAN_IN;
  assign n11217 = ~n11075 ^ P2_IR_REG_10__SCAN_IN;
  assign n17295 = ~n11217;
  assign n16822 = n11078 ^ n17295;
  assign n11076 = ~n16822;
  assign n11079 = ~n11077 | ~n11076;
  assign n11080 = ~n11081;
  assign n11082 = ~n11225 & ~n11080;
  assign n11221 = ~P2_REG2_REG_11__SCAN_IN;
  assign n17289 = ~n11225;
  assign n11085 = ~P2_REG2_REG_12__SCAN_IN;
  assign n11083 = n11089 | P2_IR_REG_11__SCAN_IN;
  assign n11084 = ~n11083 | ~P2_IR_REG_31__SCAN_IN;
  assign n11231 = ~n11084 ^ P2_IR_REG_12__SCAN_IN;
  assign n17283 = ~n11231;
  assign n11087 = ~P2_IR_REG_11__SCAN_IN;
  assign n11086 = ~P2_IR_REG_12__SCAN_IN;
  assign n11088 = ~n11087 | ~n11086;
  assign n11093 = n11089 | n11088;
  assign n11090 = ~n11093 | ~P2_IR_REG_31__SCAN_IN;
  assign n11238 = ~n11090 ^ P2_IR_REG_13__SCAN_IN;
  assign n17277 = ~n11238;
  assign n11092 = ~n11238 & ~n11091;
  assign n11243 = ~P2_REG2_REG_14__SCAN_IN;
  assign n11095 = ~n11093;
  assign n11094 = ~P2_IR_REG_13__SCAN_IN;
  assign n11096 = ~n11095 | ~n11094;
  assign n11105 = ~n11096 | ~P2_IR_REG_31__SCAN_IN;
  assign n16888 = ~n11105 ^ P2_IR_REG_14__SCAN_IN;
  assign n17271 = ~n16888;
  assign n16883 = n11243 ^ n17271;
  assign n11097 = ~n11105 | ~n11102;
  assign n11098 = ~n11097 | ~P2_IR_REG_31__SCAN_IN;
  assign n12165 = ~n11098 ^ P2_IR_REG_15__SCAN_IN;
  assign n17266 = ~n12165;
  assign n11100 = ~n12165 & ~n11099;
  assign n11259 = ~P2_REG2_REG_16__SCAN_IN;
  assign n11101 = ~P2_IR_REG_15__SCAN_IN;
  assign n11103 = ~n11102 | ~n11101;
  assign n11104 = ~n11103 | ~P2_IR_REG_31__SCAN_IN;
  assign n11108 = ~n11105 | ~n11104;
  assign n17260 = ~n11108 ^ P2_IR_REG_16__SCAN_IN;
  assign n16919 = n11259 ^ n17260;
  assign n16925 = ~n17260;
  assign n11106 = ~n16925 & ~n11259;
  assign n11109 = n11108 | P2_IR_REG_16__SCAN_IN;
  assign n11110 = ~n11109 | ~P2_IR_REG_31__SCAN_IN;
  assign n12185 = ~n11110 ^ P2_IR_REG_17__SCAN_IN;
  assign n16948 = ~n12185;
  assign n11888 = ~n17254;
  assign n13958 = ~P2_REG2_REG_18__SCAN_IN;
  assign n11114 = ~n11888 | ~n13958;
  assign n11898 = ~n11115 | ~n11114;
  assign n11116 = ~n8990 | ~P2_IR_REG_31__SCAN_IN;
  assign n11117 = ~n11116 ^ n11000;
  assign n11281 = P2_REG2_REG_19__SCAN_IN ^ n11117;
  assign n11833 = n12051 & P2_STATE_REG_SCAN_IN;
  assign n16628 = ~n11292 | ~n11833;
  assign n16939 = n16628 | n8884;
  assign n16862 = ~n16939;
  assign n11154 = ~n11118 | ~n16862;
  assign n11252 = ~n8884;
  assign n16865 = n16628 | n11252;
  assign n16937 = ~n16865;
  assign n11283 = P2_REG1_REG_19__SCAN_IN ^ n11117;
  assign n11152 = ~n17254 | ~P2_REG1_REG_18__SCAN_IN;
  assign n11897 = P2_REG1_REG_18__SCAN_IN ^ n17254;
  assign n11148 = ~P2_REG1_REG_16__SCAN_IN | ~n17260;
  assign n16916 = ~P2_REG1_REG_16__SCAN_IN ^ n16925;
  assign n11144 = ~P2_REG1_REG_14__SCAN_IN | ~n17271;
  assign n16880 = ~P2_REG1_REG_14__SCAN_IN ^ n16888;
  assign n11141 = ~P2_REG1_REG_12__SCAN_IN | ~n17283;
  assign n16843 = ~P2_REG1_REG_12__SCAN_IN ^ n11231;
  assign n11138 = ~P2_REG1_REG_10__SCAN_IN | ~n17295;
  assign n16804 = ~P2_REG1_REG_10__SCAN_IN ^ n11217;
  assign n17301 = ~n11211;
  assign n11135 = ~P2_REG1_REG_8__SCAN_IN | ~n17307;
  assign n16775 = ~P2_REG1_REG_8__SCAN_IN ^ n16768;
  assign n17313 = ~n11197;
  assign n11119 = n16625 & P2_REG1_REG_0__SCAN_IN;
  assign n11121 = ~n11023 | ~P2_REG1_REG_0__SCAN_IN;
  assign n11122 = ~n16634 | ~P2_REG1_REG_1__SCAN_IN;
  assign n16663 = ~n11122 | ~n11121;
  assign n11123 = ~n9360 | ~P2_REG1_REG_2__SCAN_IN;
  assign n11125 = ~n11124 | ~n11123;
  assign n11126 = ~n11125 | ~n17330;
  assign n11173 = ~P2_REG1_REG_4__SCAN_IN;
  assign n11127 = ~n12072 | ~P2_REG1_REG_4__SCAN_IN;
  assign n16737 = ~n17319 ^ P2_REG1_REG_6__SCAN_IN;
  assign n11130 = ~n16737;
  assign n11131 = ~n17319 | ~P2_REG1_REG_6__SCAN_IN;
  assign n11134 = ~n17313 | ~n11133;
  assign n11137 = ~n17301 | ~n11136;
  assign n11140 = ~n17289 | ~n11139;
  assign n11143 = ~n17277 | ~n11142;
  assign n11147 = ~n17266 | ~n11145;
  assign n11146 = ~P2_REG1_REG_15__SCAN_IN | ~n16899;
  assign n11151 = ~n16948 | ~n11149;
  assign n11156 = ~n11282 | ~P2_REG2_REG_1__SCAN_IN;
  assign n11155 = ~n8884 | ~P2_REG1_REG_1__SCAN_IN;
  assign n11157 = ~n11156 | ~n11155;
  assign n11158 = n11157 | n9342;
  assign n11161 = ~n11157 | ~n9342;
  assign n11160 = ~n12994 | ~P2_REG2_REG_0__SCAN_IN;
  assign n11159 = ~n8884 | ~P2_REG1_REG_0__SCAN_IN;
  assign n16629 = ~n11160 | ~n11159;
  assign n16644 = n16629 | n16625;
  assign n16643 = ~n16645 | ~n16644;
  assign n16658 = n16643 & n11161;
  assign n11163 = ~n11252 | ~P2_REG2_REG_2__SCAN_IN;
  assign n11162 = ~n8884 | ~P2_REG1_REG_2__SCAN_IN;
  assign n11164 = ~n11163 | ~n11162;
  assign n16657 = ~n11164 ^ n9360;
  assign n11166 = ~n11164;
  assign n11167 = ~n11166 & ~n11165;
  assign n16681 = ~n16660 & ~n11167;
  assign n11169 = ~n11252 | ~n9608;
  assign n11168 = ~n11273 | ~n9602;
  assign n11170 = ~n11169 | ~n11168;
  assign n16680 = n12064 ^ n11170;
  assign n11171 = ~n11170 | ~n12064;
  assign n12994 = ~n8884;
  assign n17115 = ~P2_REG2_REG_4__SCAN_IN;
  assign n11175 = ~n12994 | ~n17115;
  assign n11174 = ~n11273 | ~n11173;
  assign n11176 = n11175 & n11174;
  assign n11179 = ~n11176 | ~n12072;
  assign n11177 = ~n11176;
  assign n16701 = ~n12072;
  assign n11178 = ~n11177 | ~n16701;
  assign n16704 = ~n11179 | ~n11178;
  assign n11181 = ~n12994 | ~n17070;
  assign n16713 = ~P2_REG1_REG_5__SCAN_IN;
  assign n11180 = ~n8884 | ~n16713;
  assign n11182 = ~n11181 | ~n11180;
  assign n11184 = n11182 | n12077;
  assign n11183 = ~n11182 | ~n12077;
  assign n16723 = ~n11184 | ~n11183;
  assign n11189 = ~n12994 | ~n11186;
  assign n11187 = ~P2_REG1_REG_6__SCAN_IN;
  assign n11188 = ~n11273 | ~n11187;
  assign n11190 = ~n11189 | ~n11188;
  assign n16734 = n17319 ^ n11190;
  assign n11191 = ~n11190;
  assign n11192 = ~n11191 & ~n17319;
  assign n11196 = ~n12994 | ~n11193;
  assign n11194 = ~P2_REG1_REG_7__SCAN_IN;
  assign n11195 = ~n11273 | ~n11194;
  assign n11198 = ~n11196 | ~n11195;
  assign n16755 = ~n11198 ^ n11197;
  assign n11199 = ~n11198;
  assign n11200 = ~n17313 & ~n11199;
  assign n11204 = ~n12994 | ~n17022;
  assign n11202 = ~P2_REG1_REG_8__SCAN_IN;
  assign n11203 = ~n11273 | ~n11202;
  assign n11205 = ~n11204 | ~n11203;
  assign n16771 = ~n16768 ^ n11205;
  assign n11206 = ~n11205;
  assign n11207 = ~n17307 & ~n11206;
  assign n11210 = ~n11252 | ~n16984;
  assign n11208 = ~P2_REG1_REG_9__SCAN_IN;
  assign n11209 = ~n11273 | ~n11208;
  assign n11212 = ~n11210 | ~n11209;
  assign n16791 = ~n11212 ^ n11211;
  assign n11213 = ~n11212;
  assign n11214 = ~n11213 & ~n17301;
  assign n11216 = ~n11252 | ~P2_REG2_REG_10__SCAN_IN;
  assign n11215 = ~n11273 | ~P2_REG1_REG_10__SCAN_IN;
  assign n11218 = n11216 & n11215;
  assign n16814 = ~n11218 & ~n11217;
  assign n11220 = ~n16816 & ~n16814;
  assign n11219 = ~n11218;
  assign n16813 = ~n11219 & ~n17295;
  assign n11224 = ~n11252 | ~n11221;
  assign n11222 = ~P2_REG1_REG_11__SCAN_IN;
  assign n11223 = ~n11273 | ~n11222;
  assign n11226 = ~n11224 | ~n11223;
  assign n16830 = ~n11226 ^ n11225;
  assign n11227 = ~n11226;
  assign n11228 = ~n11227 & ~n17289;
  assign n11230 = ~n11252 | ~P2_REG2_REG_12__SCAN_IN;
  assign n11229 = ~n11273 | ~P2_REG1_REG_12__SCAN_IN;
  assign n11232 = ~n11230 | ~n11229;
  assign n16848 = n11231 ^ n11232;
  assign n11233 = ~n17283 & ~n11232;
  assign n11237 = ~n11252 | ~n11234;
  assign n11235 = ~P2_REG1_REG_13__SCAN_IN;
  assign n11236 = ~n11273 | ~n11235;
  assign n11239 = ~n11237 | ~n11236;
  assign n16867 = ~n11239 ^ n11238;
  assign n11242 = ~n16868 & ~n16867;
  assign n11240 = ~n11239;
  assign n11241 = ~n17277 & ~n11240;
  assign n16886 = ~n11242 & ~n11241;
  assign n11246 = ~n11252 | ~n11243;
  assign n11244 = ~P2_REG1_REG_14__SCAN_IN;
  assign n11245 = ~n11273 | ~n11244;
  assign n11247 = ~n11246 | ~n11245;
  assign n16885 = ~n16888 ^ n11247;
  assign n11250 = ~n16886 & ~n16885;
  assign n11248 = ~n11247;
  assign n11249 = ~n17271 & ~n11248;
  assign n11255 = ~n11252 | ~n11251;
  assign n11253 = ~P2_REG1_REG_15__SCAN_IN;
  assign n11254 = ~n11273 | ~n11253;
  assign n11256 = ~n11255 | ~n11254;
  assign n16903 = ~n12165 ^ n11256;
  assign n11257 = ~n11256;
  assign n11258 = ~n17266 & ~n11257;
  assign n11262 = ~n11252 | ~n11259;
  assign n11260 = ~P2_REG1_REG_16__SCAN_IN;
  assign n11261 = ~n11273 | ~n11260;
  assign n11263 = ~n11262 | ~n11261;
  assign n16921 = n11263 ^ n17260;
  assign n11264 = ~n11263;
  assign n11268 = ~n11252 | ~n11265;
  assign n11266 = ~P2_REG1_REG_17__SCAN_IN;
  assign n11267 = ~n8884 | ~n11266;
  assign n11269 = ~n11268 | ~n11267;
  assign n16941 = ~n12185 ^ n11269;
  assign n11272 = ~n16942 & ~n16941;
  assign n11270 = ~n11269;
  assign n11271 = ~n16948 & ~n11270;
  assign n11276 = ~n11272 & ~n11271;
  assign n11275 = ~n11252 | ~P2_REG2_REG_18__SCAN_IN;
  assign n11274 = ~n11273 | ~P2_REG1_REG_18__SCAN_IN;
  assign n11277 = ~n11275 | ~n11274;
  assign n11884 = ~n11276 & ~n11277;
  assign n11279 = ~n11276;
  assign n11278 = ~n11277;
  assign n11883 = ~n11279 & ~n11278;
  assign n11280 = ~n11883 & ~n17254;
  assign n11287 = ~n11884 & ~n11280;
  assign n11285 = ~n11281 & ~n11273;
  assign n11284 = ~n11283 & ~n11282;
  assign n11286 = ~n11285 & ~n11284;
  assign n11288 = ~n11287 ^ n11286;
  assign n12995 = ~n12051;
  assign n16817 = ~P2_U3893 | ~n12995;
  assign n16945 = ~n11289 & ~P2_U3150;
  assign n11290 = ~P2_ADDR_REG_19__SCAN_IN | ~n16945;
  assign n11294 = ~P2_U3893 | ~n12051;
  assign n11822 = ~n8884 & ~P2_U3151;
  assign n11291 = n11822 & n12995;
  assign n11293 = ~n11292 | ~n11291;
  assign n16924 = ~n16949;
  assign n11770 = ~n11117;
  assign n11295 = ~n16924 | ~n11770;
  assign n13535 = ~P2_REG3_REG_19__SCAN_IN | ~P2_U3151;
  assign n11297 = ~n11296 & ~P1_U3086;
  assign P1_U3973 = ~n11337;
  assign n11299 = ~n15346 | ~n11298;
  assign n11301 = n11300 ^ n11299;
  assign n11306 = ~n11301 | ~n15376;
  assign n11303 = ~n11302 & ~P1_U3086;
  assign n15355 = ~n11304 | ~n11303;
  assign n11305 = ~P1_REG3_REG_1__SCAN_IN | ~n15355;
  assign n11312 = ~n11306 | ~n11305;
  assign n11308 = ~n15319 & ~n9307;
  assign n13035 = ~n16182;
  assign n11307 = ~n15333 & ~n13035;
  assign n11310 = ~n11308 & ~n11307;
  assign n15360 = ~n15332;
  assign n11309 = ~n15360 | ~n15980;
  assign n11311 = ~n11310 | ~n11309;
  assign P1_U3222 = n11312 | n11311;
  assign n11313 = ~n13271 | ~SI_0_;
  assign n11787 = ~n11313 ^ P1_DATAO_REG_0__SCAN_IN;
  assign n11315 = ~n11787 | ~P2_U3151;
  assign n11314 = ~n9288 | ~P2_STATE_REG_SCAN_IN;
  assign P2_U3295 = ~n11315 | ~n11314;
  assign n11318 = ~n11316 | ~P1_U3086;
  assign n11317 = ~P1_IR_REG_0__SCAN_IN | ~P1_STATE_REG_SCAN_IN;
  assign P1_U3355 = ~n11318 | ~n11317;
  assign n11830 = ~n17341;
  assign n11322 = ~n16135 | ~n11830;
  assign n11320 = ~n12072 & ~P2_U3151;
  assign n17226 = ~n17338;
  assign n12071 = ~P1_DATAO_REG_4__SCAN_IN;
  assign n11319 = ~n17226 & ~n12071;
  assign n11321 = ~n11320 & ~n11319;
  assign P2_U3291 = ~n11322 | ~n11321;
  assign n11368 = ~n11809;
  assign n11326 = ~n11728;
  assign n11325 = ~n12999 & ~P2_U3151;
  assign n17348 = ~n17350;
  assign n11374 = ~n11326 & ~n17348;
  assign n11327 = ~P2_D_REG_2__SCAN_IN;
  assign P2_U3263 = ~n11397 & ~n11327;
  assign n11328 = ~P2_D_REG_3__SCAN_IN;
  assign P2_U3262 = ~n11397 & ~n11328;
  assign n11329 = ~P2_D_REG_4__SCAN_IN;
  assign P2_U3261 = ~n11374 & ~n11329;
  assign n11330 = ~P2_D_REG_5__SCAN_IN;
  assign P2_U3260 = ~n11374 & ~n11330;
  assign n11331 = ~P2_D_REG_6__SCAN_IN;
  assign P2_U3259 = ~n11374 & ~n11331;
  assign n11332 = ~P2_D_REG_7__SCAN_IN;
  assign P2_U3258 = ~n11374 & ~n11332;
  assign n11334 = ~n11905 | ~P1_U3973;
  assign n11333 = ~n11337 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P1_U3557 = ~n11334 | ~n11333;
  assign n11336 = ~n15980 | ~P1_U3973;
  assign n11335 = ~n11337 | ~P1_DATAO_REG_0__SCAN_IN;
  assign P1_U3554 = ~n11336 | ~n11335;
  assign n11339 = ~n9310 | ~P1_U3973;
  assign n11338 = ~n11337 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P1_U3555 = ~n11339 | ~n11338;
  assign n11341 = ~n15640 | ~P1_U3973;
  assign n11340 = ~n11337 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P1_U3568 = ~n11341 | ~n11340;
  assign n11343 = ~n15729 | ~P1_U3973;
  assign n11342 = ~n11337 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P1_U3562 = ~n11343 | ~n11342;
  assign n11977 = ~n14998;
  assign n11345 = ~n11977 | ~P1_U3973;
  assign n11344 = ~n11337 | ~P1_DATAO_REG_17__SCAN_IN;
  assign P1_U3571 = ~n11345 | ~n11344;
  assign n11347 = ~n15844 | ~P1_U3973;
  assign n11346 = ~n11337 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P1_U3560 = ~n11347 | ~n11346;
  assign n11349 = ~n15823 | ~P1_U3973;
  assign n11348 = ~n11337 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P1_U3561 = ~n11349 | ~n11348;
  assign n11351 = ~n13151 | ~P1_U3973;
  assign n11350 = ~n11337 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P1_U3570 = ~n11351 | ~n11350;
  assign n11353 = ~n15711 | ~P1_U3973;
  assign n11352 = ~n11337 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P1_U3565 = ~n11353 | ~n11352;
  assign n11355 = ~n9305 | ~P1_U3973;
  assign n11354 = ~n11337 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P1_U3566 = ~n11355 | ~n11354;
  assign n11357 = ~n15661 | ~P1_U3973;
  assign n11356 = ~n11337 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P1_U3567 = ~n11357 | ~n11356;
  assign n15618 = ~n14997;
  assign n11359 = ~n15618 | ~P1_U3973;
  assign n11358 = ~n11337 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P1_U3569 = ~n11359 | ~n11358;
  assign n11361 = ~n11903 | ~P1_U3973;
  assign n11360 = ~n11337 | ~P1_DATAO_REG_4__SCAN_IN;
  assign P1_U3558 = ~n11361 | ~n11360;
  assign n11363 = ~n15876 | ~P1_U3973;
  assign n11362 = ~n11337 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P1_U3559 = ~n11363 | ~n11362;
  assign n11365 = ~n15734 | ~P1_U3973;
  assign n11364 = ~n11337 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P1_U3564 = ~n11365 | ~n11364;
  assign n11367 = ~n15771 | ~P1_U3973;
  assign n11366 = ~n11337 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P1_U3563 = ~n11367 | ~n11366;
  assign n11373 = ~n11374 & ~P2_D_REG_0__SCAN_IN;
  assign n11371 = ~n11323;
  assign n11369 = ~n11368 & ~P2_U3151;
  assign n11370 = ~n12993 | ~n11369;
  assign n11372 = ~n11371 & ~n11370;
  assign P2_U3376 = ~n11373 & ~n11372;
  assign n11397 = n11374;
  assign n11375 = ~P2_D_REG_19__SCAN_IN;
  assign P2_U3246 = ~n11397 & ~n11375;
  assign n11376 = ~P2_D_REG_20__SCAN_IN;
  assign P2_U3245 = ~n11397 & ~n11376;
  assign n11377 = ~P2_D_REG_10__SCAN_IN;
  assign P2_U3255 = ~n11397 & ~n11377;
  assign n11378 = ~P2_D_REG_11__SCAN_IN;
  assign P2_U3254 = ~n11397 & ~n11378;
  assign n11732 = ~P2_D_REG_8__SCAN_IN;
  assign P2_U3257 = ~n11397 & ~n11732;
  assign n11379 = ~P2_D_REG_21__SCAN_IN;
  assign P2_U3244 = ~n11397 & ~n11379;
  assign n11380 = ~P2_D_REG_13__SCAN_IN;
  assign P2_U3252 = ~n11397 & ~n11380;
  assign n11381 = ~P2_D_REG_14__SCAN_IN;
  assign P2_U3251 = ~n11397 & ~n11381;
  assign n11382 = ~P2_D_REG_15__SCAN_IN;
  assign P2_U3250 = ~n11397 & ~n11382;
  assign n11383 = ~P2_D_REG_18__SCAN_IN;
  assign P2_U3247 = ~n11397 & ~n11383;
  assign n11384 = ~P2_D_REG_17__SCAN_IN;
  assign P2_U3248 = ~n11397 & ~n11384;
  assign n11731 = ~P2_D_REG_9__SCAN_IN;
  assign P2_U3256 = ~n11397 & ~n11731;
  assign n11385 = ~P2_D_REG_23__SCAN_IN;
  assign P2_U3242 = ~n11397 & ~n11385;
  assign n11386 = ~P2_D_REG_24__SCAN_IN;
  assign P2_U3241 = ~n11397 & ~n11386;
  assign n11387 = ~P2_D_REG_25__SCAN_IN;
  assign P2_U3240 = ~n11397 & ~n11387;
  assign n11388 = ~P2_D_REG_12__SCAN_IN;
  assign P2_U3253 = ~n11397 & ~n11388;
  assign n11389 = ~P2_D_REG_26__SCAN_IN;
  assign P2_U3239 = ~n11397 & ~n11389;
  assign n11390 = ~P2_D_REG_27__SCAN_IN;
  assign P2_U3238 = ~n11397 & ~n11390;
  assign n11391 = ~P2_D_REG_28__SCAN_IN;
  assign P2_U3237 = ~n11397 & ~n11391;
  assign n11392 = ~P2_D_REG_16__SCAN_IN;
  assign P2_U3249 = ~n11397 & ~n11392;
  assign n11393 = ~P2_D_REG_31__SCAN_IN;
  assign P2_U3234 = ~n11397 & ~n11393;
  assign n11394 = ~P2_D_REG_22__SCAN_IN;
  assign P2_U3243 = ~n11397 & ~n11394;
  assign n11395 = ~P2_D_REG_30__SCAN_IN;
  assign P2_U3235 = ~n11397 & ~n11395;
  assign n11396 = ~P2_D_REG_29__SCAN_IN;
  assign P2_U3236 = ~n11397 & ~n11396;
  assign n11402 = ~n16054 | ~n11830;
  assign n11398 = ~P1_DATAO_REG_17__SCAN_IN;
  assign n11400 = ~n17226 & ~n11398;
  assign n11399 = ~P2_U3151 & ~n16948;
  assign n11401 = ~n11400 & ~n11399;
  assign P2_U3278 = ~n11402 | ~n11401;
  assign n11404 = ~P2_IR_REG_29__SCAN_IN;
  assign n14354 = ~n11406 | ~n11404;
  assign n12327 = n11486;
  assign n11409 = ~n12327 | ~P2_REG2_REG_11__SCAN_IN;
  assign n12216 = n11531;
  assign n11408 = ~n12216 | ~P2_REG1_REG_11__SCAN_IN;
  assign n11418 = n11409 & n11408;
  assign n12219 = n14362 & n11878;
  assign n11412 = n11495 & P2_REG3_REG_11__SCAN_IN;
  assign n16958 = n11412 | n11581;
  assign n11416 = ~n8889 | ~n16958;
  assign n11415 = ~n12881 | ~P2_REG0_REG_11__SCAN_IN;
  assign n11417 = n11416 & n11415;
  assign n14116 = ~n16507;
  assign n11420 = ~n14116 | ~P2_U3893;
  assign n17550 = ~P2_U3893;
  assign n11419 = ~n17550 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P2_U3502 = ~n11420 | ~n11419;
  assign n11422 = ~n11531 | ~P2_REG1_REG_2__SCAN_IN;
  assign n11421 = ~n12881 | ~P2_REG0_REG_2__SCAN_IN;
  assign n11426 = ~n11422 | ~n11421;
  assign n11424 = ~n12290 | ~P2_REG2_REG_2__SCAN_IN;
  assign n11423 = ~n8889 | ~P2_REG3_REG_2__SCAN_IN;
  assign n11425 = ~n11424 | ~n11423;
  assign n11428 = ~n17168 | ~P2_U3893;
  assign n11427 = ~n17550 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P2_U3493 = ~n11428 | ~n11427;
  assign n11430 = ~n12216 | ~P2_REG1_REG_5__SCAN_IN;
  assign n11429 = ~n12881 | ~P2_REG0_REG_5__SCAN_IN;
  assign n11435 = ~n11430 | ~n11429;
  assign n11433 = ~n11486 | ~P2_REG2_REG_5__SCAN_IN;
  assign n11563 = n12219;
  assign n17071 = ~n11458 ^ P2_REG3_REG_5__SCAN_IN;
  assign n11431 = ~n17071;
  assign n11432 = ~n11563 | ~n11431;
  assign n11434 = ~n11433 | ~n11432;
  assign n11437 = ~n17102 | ~P2_U3893;
  assign n11436 = ~n17550 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P2_U3496 = ~n11437 | ~n11436;
  assign n11580 = ~P2_REG3_REG_12__SCAN_IN;
  assign n11470 = ~P2_REG3_REG_13__SCAN_IN;
  assign n13574 = ~P2_REG3_REG_16__SCAN_IN;
  assign n11448 = ~n11438 | ~n13574;
  assign n11439 = n11438 | n13574;
  assign n14009 = ~n11448 | ~n11439;
  assign n11441 = ~n14009 | ~n12219;
  assign n11440 = ~n12303 | ~P2_REG1_REG_16__SCAN_IN;
  assign n11445 = ~n11441 | ~n11440;
  assign n11443 = ~n12327 | ~P2_REG2_REG_16__SCAN_IN;
  assign n11442 = ~n12881 | ~P2_REG0_REG_16__SCAN_IN;
  assign n11444 = ~n11443 | ~n11442;
  assign n11447 = ~n14270 | ~P2_U3893;
  assign n11446 = ~n17550 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P2_U3507 = ~n11447 | ~n11446;
  assign n11449 = ~n11448 | ~P2_REG3_REG_17__SCAN_IN;
  assign n13984 = ~n11590 | ~n11449;
  assign n11455 = ~n13984 | ~n8889;
  assign n11451 = ~n12303 | ~P2_REG1_REG_17__SCAN_IN;
  assign n11450 = ~n12881 | ~P2_REG0_REG_17__SCAN_IN;
  assign n11453 = ~n11451 | ~n11450;
  assign n11452 = n12327 & P2_REG2_REG_17__SCAN_IN;
  assign n11454 = ~n11453 & ~n11452;
  assign n14259 = ~n11455 | ~n11454;
  assign n11457 = ~n14259 | ~P2_U3893;
  assign n11456 = ~n17550 | ~P2_DATAO_REG_17__SCAN_IN;
  assign P2_U3508 = ~n11457 | ~n11456;
  assign n11459 = P2_REG3_REG_4__SCAN_IN & P2_REG3_REG_3__SCAN_IN;
  assign n17112 = n11459 | n11458;
  assign n11461 = ~n12219 | ~n17112;
  assign n11460 = ~n12881 | ~P2_REG0_REG_4__SCAN_IN;
  assign n11465 = ~n11461 | ~n11460;
  assign n11463 = ~n12327 | ~P2_REG2_REG_4__SCAN_IN;
  assign n11462 = ~n11531 | ~P2_REG1_REG_4__SCAN_IN;
  assign n11464 = ~n11463 | ~n11462;
  assign n17132 = n11465 | n11464;
  assign n11467 = ~n17132 | ~P2_U3893;
  assign n11466 = ~n17550 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P2_U3495 = ~n11467 | ~n11466;
  assign n11469 = ~n11486 | ~P2_REG2_REG_13__SCAN_IN;
  assign n11468 = ~n12881 | ~P2_REG0_REG_13__SCAN_IN;
  assign n11476 = n11469 & n11468;
  assign n11472 = n11471 | n11470;
  assign n14076 = ~n11534 | ~n11472;
  assign n11474 = ~n12219 | ~n14076;
  assign n11473 = ~n12216 | ~P2_REG1_REG_13__SCAN_IN;
  assign n11475 = n11474 & n11473;
  assign n11478 = ~n17465 | ~P2_U3893;
  assign n11477 = ~n17550 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P2_U3504 = ~n11478 | ~n11477;
  assign n11480 = ~n12290 | ~P2_REG2_REG_0__SCAN_IN;
  assign n11479 = ~n12881 | ~P2_REG0_REG_0__SCAN_IN;
  assign n11482 = ~n12219 | ~P2_REG3_REG_0__SCAN_IN;
  assign n11481 = ~n11531 | ~P2_REG1_REG_0__SCAN_IN;
  assign n11484 = ~n17167 | ~P2_U3893;
  assign n11483 = ~n17550 | ~P2_DATAO_REG_0__SCAN_IN;
  assign P2_U3491 = ~n11484 | ~n11483;
  assign n11485 = ~n11531 | ~P2_REG1_REG_1__SCAN_IN;
  assign n11488 = ~n11486 | ~P2_REG2_REG_1__SCAN_IN;
  assign n11487 = ~n12219 | ~P2_REG3_REG_1__SCAN_IN;
  assign n11490 = ~n17151 | ~P2_U3893;
  assign n11489 = ~n17550 | ~P2_DATAO_REG_1__SCAN_IN;
  assign P2_U3492 = ~n11490 | ~n11489;
  assign n11492 = ~n11531 | ~P2_REG1_REG_10__SCAN_IN;
  assign n11491 = ~n12881 | ~P2_REG0_REG_10__SCAN_IN;
  assign n11499 = ~n11492 | ~n11491;
  assign n11497 = ~n12327 | ~P2_REG2_REG_10__SCAN_IN;
  assign n11494 = ~n11493 | ~P2_REG3_REG_10__SCAN_IN;
  assign n16449 = ~n11495 | ~n11494;
  assign n11496 = ~n8889 | ~n16449;
  assign n11498 = ~n11497 | ~n11496;
  assign n16989 = n11499 | n11498;
  assign n11501 = ~n16989 | ~P2_U3893;
  assign n11500 = ~n17550 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P2_U3501 = ~n11501 | ~n11500;
  assign n11503 = ~n11531 | ~P2_REG1_REG_7__SCAN_IN;
  assign n11502 = ~n12881 | ~P2_REG0_REG_7__SCAN_IN;
  assign n11509 = ~n11503 | ~n11502;
  assign n11507 = ~n12327 | ~P2_REG2_REG_7__SCAN_IN;
  assign n17046 = ~n11504 ^ n9501;
  assign n11505 = ~n17046;
  assign n11506 = ~n8889 | ~n11505;
  assign n11508 = ~n11507 | ~n11506;
  assign n11511 = ~n17053 | ~P2_U3893;
  assign n11510 = ~n17550 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P2_U3498 = ~n11511 | ~n11510;
  assign n11516 = ~n12290 | ~P2_REG2_REG_8__SCAN_IN;
  assign n11514 = ~n11513 & ~n11512;
  assign n17019 = n11572 | n11514;
  assign n11515 = ~n8889 | ~n17019;
  assign n11520 = ~n11516 | ~n11515;
  assign n11518 = ~n11531 | ~P2_REG1_REG_8__SCAN_IN;
  assign n11517 = ~n12881 | ~P2_REG0_REG_8__SCAN_IN;
  assign n11519 = ~n11518 | ~n11517;
  assign n11522 = ~n17036 | ~P2_U3893;
  assign n11521 = ~n17550 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P2_U3499 = ~n11522 | ~n11521;
  assign n11524 = ~n12216 | ~P2_REG1_REG_15__SCAN_IN;
  assign n11523 = ~n12881 | ~P2_REG0_REG_15__SCAN_IN;
  assign n11526 = ~n11524 | ~n11523;
  assign n11525 = n12327 & P2_REG2_REG_15__SCAN_IN;
  assign n11528 = ~n11526 & ~n11525;
  assign n14033 = ~n11536 ^ P2_REG3_REG_15__SCAN_IN;
  assign n11527 = ~n14033 | ~n12219;
  assign n14280 = ~n14061;
  assign n11530 = ~n14280 | ~P2_U3893;
  assign n11529 = ~n17550 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P2_U3506 = ~n11530 | ~n11529;
  assign n11533 = ~n12327 | ~P2_REG2_REG_14__SCAN_IN;
  assign n11532 = ~n12303 | ~P2_REG1_REG_14__SCAN_IN;
  assign n11540 = ~n11533 | ~n11532;
  assign n11535 = ~n11534 | ~P2_REG3_REG_14__SCAN_IN;
  assign n14053 = ~n11536 | ~n11535;
  assign n11538 = ~n12219 | ~n14053;
  assign n11537 = ~n12881 | ~P2_REG0_REG_14__SCAN_IN;
  assign n11539 = ~n11538 | ~n11537;
  assign n11542 = ~n14291 | ~P2_U3893;
  assign n11541 = ~n17550 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P2_U3505 = ~n11542 | ~n11541;
  assign n11544 = ~n11531 | ~P2_REG1_REG_3__SCAN_IN;
  assign n11543 = ~n12881 | ~P2_REG0_REG_3__SCAN_IN;
  assign n11548 = n11544 & n11543;
  assign n11546 = ~n12290 | ~P2_REG2_REG_3__SCAN_IN;
  assign n11545 = ~n11563 | ~n9497;
  assign n11547 = n11546 & n11545;
  assign n17150 = ~n16543;
  assign n11550 = ~n17150 | ~P2_U3893;
  assign n11549 = ~n17550 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P2_U3494 = ~n11550 | ~n11549;
  assign n13677 = ~n11590 ^ n9494;
  assign n12256 = ~n12219;
  assign n11556 = n13677 | n12256;
  assign n11552 = ~n12303 | ~P2_REG1_REG_18__SCAN_IN;
  assign n11551 = ~n12881 | ~P2_REG0_REG_18__SCAN_IN;
  assign n11554 = ~n11552 | ~n11551;
  assign n11553 = n11486 & P2_REG2_REG_18__SCAN_IN;
  assign n11555 = ~n11554 & ~n11553;
  assign n13926 = ~n11556 | ~n11555;
  assign n11558 = ~n13926 | ~P2_U3893;
  assign n11557 = ~n17550 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P2_U3509 = ~n11558 | ~n11557;
  assign n11560 = ~n11531 | ~P2_REG1_REG_6__SCAN_IN;
  assign n11559 = ~n12881 | ~P2_REG0_REG_6__SCAN_IN;
  assign n11567 = n11560 & n11559;
  assign n11565 = ~n12327 | ~P2_REG2_REG_6__SCAN_IN;
  assign n17065 = ~n11561 ^ n9502;
  assign n11562 = ~n17065;
  assign n11564 = ~n11563 | ~n11562;
  assign n11566 = n11565 & n11564;
  assign n17078 = ~n12644;
  assign n11569 = ~n17078 | ~P2_U3893;
  assign n11568 = ~n17550 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P2_U3497 = ~n11569 | ~n11568;
  assign n11571 = ~n11531 | ~P2_REG1_REG_9__SCAN_IN;
  assign n11570 = ~n12881 | ~P2_REG0_REG_9__SCAN_IN;
  assign n11577 = ~n11571 | ~n11570;
  assign n11575 = ~n12327 | ~P2_REG2_REG_9__SCAN_IN;
  assign n16983 = ~n11572 ^ P2_REG3_REG_9__SCAN_IN;
  assign n11573 = ~n16983;
  assign n11574 = ~n8889 | ~n11573;
  assign n11576 = ~n11575 | ~n11574;
  assign n11579 = ~n17009 | ~P2_U3893;
  assign n11578 = ~n17550 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P2_U3500 = ~n11579 | ~n11578;
  assign n16510 = ~n11581 ^ n11580;
  assign n11583 = ~n11563 | ~n16510;
  assign n11582 = ~n12303 | ~P2_REG1_REG_12__SCAN_IN;
  assign n11587 = n11583 & n11582;
  assign n11585 = ~n12327 | ~P2_REG2_REG_12__SCAN_IN;
  assign n11584 = ~n12881 | ~P2_REG0_REG_12__SCAN_IN;
  assign n11586 = n11585 & n11584;
  assign n16974 = ~n13644;
  assign n11589 = ~n16974 | ~P2_U3893;
  assign n11588 = ~n17550 | ~P2_DATAO_REG_12__SCAN_IN;
  assign P2_U3503 = ~n11589 | ~n11588;
  assign n13933 = ~n12220 ^ P2_REG3_REG_19__SCAN_IN;
  assign n11596 = ~n13933 | ~n12219;
  assign n11592 = ~n12303 | ~P2_REG1_REG_19__SCAN_IN;
  assign n11591 = ~n12881 | ~P2_REG0_REG_19__SCAN_IN;
  assign n11594 = ~n11592 | ~n11591;
  assign n11593 = n12290 & P2_REG2_REG_19__SCAN_IN;
  assign n11595 = ~n11594 & ~n11593;
  assign n11598 = ~n13904 | ~P2_U3893;
  assign n11597 = ~n17550 | ~P2_DATAO_REG_19__SCAN_IN;
  assign P2_U3510 = ~n11598 | ~n11597;
  assign n14397 = ~P1_REG3_REG_10__SCAN_IN | ~P1_U3086;
  assign n11599 = ~n13367 | ~n13383;
  assign n11631 = n11599 & n9921;
  assign n16026 = n13383 | P1_U3086;
  assign n11601 = ~n11600;
  assign n11630 = ~n16026 | ~n11601;
  assign n11602 = ~n11630;
  assign n15607 = ~n11631 & ~n11602;
  assign n11603 = ~n15607 | ~P1_ADDR_REG_10__SCAN_IN;
  assign n11658 = ~n14397 | ~n11603;
  assign n14650 = P1_REG1_REG_10__SCAN_IN ^ n16101;
  assign n15408 = P1_REG1_REG_1__SCAN_IN ^ n16155;
  assign n15407 = ~n11604 & ~n15423;
  assign n15406 = ~n15408 | ~n15407;
  assign n11605 = ~n16155 | ~P1_REG1_REG_1__SCAN_IN;
  assign n15416 = ~n15406 | ~n11605;
  assign n15417 = P1_REG1_REG_2__SCAN_IN ^ n16148;
  assign n11607 = ~n15416 | ~n15417;
  assign n11606 = ~n16148 | ~P1_REG1_REG_2__SCAN_IN;
  assign n11676 = ~n11607 | ~n11606;
  assign n11608 = ~P1_REG1_REG_3__SCAN_IN;
  assign n11677 = ~n16142 ^ n11608;
  assign n11610 = ~n11676 | ~n11677;
  assign n11609 = ~n16142 | ~P1_REG1_REG_3__SCAN_IN;
  assign n15445 = ~n11610 | ~n11609;
  assign n11611 = ~P1_REG1_REG_4__SCAN_IN;
  assign n15446 = ~n16136 ^ n11611;
  assign n11613 = ~n15445 | ~n15446;
  assign n11612 = ~n16136 | ~P1_REG1_REG_4__SCAN_IN;
  assign n15470 = ~n11613 | ~n11612;
  assign n11614 = ~P1_REG1_REG_5__SCAN_IN;
  assign n15471 = ~n16128 ^ n11614;
  assign n11616 = ~n15470 | ~n15471;
  assign n11615 = ~n16128 | ~P1_REG1_REG_5__SCAN_IN;
  assign n15478 = ~n11616 | ~n11615;
  assign n11617 = ~P1_REG1_REG_6__SCAN_IN;
  assign n15479 = ~n15477 ^ n11617;
  assign n11619 = ~n15478 | ~n15479;
  assign n11618 = ~n15477 | ~P1_REG1_REG_6__SCAN_IN;
  assign n11662 = ~n11619 | ~n11618;
  assign n11620 = ~P1_REG1_REG_7__SCAN_IN;
  assign n11663 = ~n11672 ^ n11620;
  assign n11622 = ~n11662 | ~n11663;
  assign n11621 = ~n11672 | ~P1_REG1_REG_7__SCAN_IN;
  assign n11689 = ~n11622 | ~n11621;
  assign n11623 = ~P1_REG1_REG_8__SCAN_IN;
  assign n11690 = ~n11699 ^ n11623;
  assign n11625 = ~n11689 | ~n11690;
  assign n11624 = ~n11699 | ~P1_REG1_REG_8__SCAN_IN;
  assign n11707 = ~n11625 | ~n11624;
  assign n16107 = ~n11717;
  assign n11626 = ~P1_REG1_REG_9__SCAN_IN;
  assign n11628 = ~n16107 | ~n11626;
  assign n11627 = ~n11717 | ~P1_REG1_REG_9__SCAN_IN;
  assign n11706 = ~n11628 | ~n11627;
  assign n11705 = ~n11707 & ~n11706;
  assign n11629 = ~n11628;
  assign n14651 = ~n11705 & ~n11629;
  assign n11632 = n14650 ^ n14651;
  assign n15392 = ~n11631 | ~n11630;
  assign n15432 = ~n15386;
  assign n15591 = ~n15392 & ~n15432;
  assign n11656 = ~n11632 | ~n15591;
  assign n14676 = ~n16101 ^ P1_REG2_REG_10__SCAN_IN;
  assign n15399 = P1_REG2_REG_1__SCAN_IN ^ n16155;
  assign n15995 = ~P1_REG2_REG_0__SCAN_IN;
  assign n15400 = ~n15423 & ~n15995;
  assign n11634 = ~n15399 | ~n15400;
  assign n11633 = ~n16155 | ~P1_REG2_REG_1__SCAN_IN;
  assign n15438 = ~n11634 | ~n11633;
  assign n15437 = P1_REG2_REG_2__SCAN_IN ^ n16148;
  assign n11636 = ~n15438 | ~n15437;
  assign n11635 = ~n16148 | ~P1_REG2_REG_2__SCAN_IN;
  assign n11679 = ~n11636 | ~n11635;
  assign n11637 = ~P1_REG2_REG_3__SCAN_IN;
  assign n11680 = ~n16142 ^ n11637;
  assign n11639 = ~n11679 | ~n11680;
  assign n11638 = ~n16142 | ~P1_REG2_REG_3__SCAN_IN;
  assign n15453 = ~n11639 | ~n11638;
  assign n15452 = P1_REG2_REG_4__SCAN_IN ^ n16136;
  assign n11641 = ~n15453 | ~n15452;
  assign n11640 = ~n16136 | ~P1_REG2_REG_4__SCAN_IN;
  assign n15460 = ~n11641 | ~n11640;
  assign n15459 = P1_REG2_REG_5__SCAN_IN ^ n16128;
  assign n11643 = ~n15460 | ~n15459;
  assign n11642 = ~n16128 | ~P1_REG2_REG_5__SCAN_IN;
  assign n15485 = n11643 & n11642;
  assign n15486 = ~n15477 ^ P1_REG2_REG_6__SCAN_IN;
  assign n11645 = ~n15485 & ~n15486;
  assign n16122 = ~n15477;
  assign n15825 = ~P1_REG2_REG_6__SCAN_IN;
  assign n11644 = ~n16122 & ~n15825;
  assign n11665 = ~n11645 & ~n11644;
  assign n11666 = ~n11672 ^ P1_REG2_REG_7__SCAN_IN;
  assign n11647 = ~n11665 & ~n11666;
  assign n16117 = ~n11672;
  assign n15780 = ~P1_REG2_REG_7__SCAN_IN;
  assign n11646 = ~n16117 & ~n15780;
  assign n11692 = ~n11647 & ~n11646;
  assign n11693 = ~n11699 ^ P1_REG2_REG_8__SCAN_IN;
  assign n11650 = ~n11692 & ~n11693;
  assign n16112 = ~n11699;
  assign n11648 = ~P1_REG2_REG_8__SCAN_IN;
  assign n11649 = ~n16112 & ~n11648;
  assign n11702 = ~n11650 & ~n11649;
  assign n11652 = n11717 | P1_REG2_REG_9__SCAN_IN;
  assign n11651 = ~n11717 | ~P1_REG2_REG_9__SCAN_IN;
  assign n11703 = n11652 & n11651;
  assign n11653 = ~n11702 | ~n11703;
  assign n14677 = ~n11653 | ~n11652;
  assign n11654 = n14676 ^ n14677;
  assign n13482 = n15431 | n15386;
  assign n15596 = n15392 | n13482;
  assign n15574 = ~n15596;
  assign n11655 = ~n11654 | ~n15574;
  assign n11657 = ~n11656 | ~n11655;
  assign n11660 = ~n11658 & ~n11657;
  assign n15604 = ~n15392 & ~n15426;
  assign n11659 = ~n15604 | ~n16101;
  assign P1_U3253 = ~n11660 | ~n11659;
  assign n15258 = ~P1_REG3_REG_7__SCAN_IN | ~P1_U3086;
  assign n11661 = ~n15607 | ~P1_ADDR_REG_7__SCAN_IN;
  assign n11671 = ~n15258 | ~n11661;
  assign n11664 = n11663 ^ n11662;
  assign n11669 = ~n15591 | ~n11664;
  assign n11667 = n11666 ^ n11665;
  assign n11668 = ~n11667 | ~n15574;
  assign n11670 = ~n11669 | ~n11668;
  assign n11674 = ~n11671 & ~n11670;
  assign n11673 = ~n15604 | ~n11672;
  assign P1_U3250 = ~n11674 | ~n11673;
  assign n15272 = ~P1_REG3_REG_3__SCAN_IN | ~P1_U3086;
  assign n11675 = ~n15607 | ~P1_ADDR_REG_3__SCAN_IN;
  assign n11685 = ~n15272 | ~n11675;
  assign n11678 = n11677 ^ n11676;
  assign n11683 = ~n15591 | ~n11678;
  assign n11681 = n11680 ^ n11679;
  assign n11682 = ~n11681 | ~n15574;
  assign n11684 = ~n11683 | ~n11682;
  assign n11687 = ~n11685 & ~n11684;
  assign n11686 = ~n15604 | ~n16142;
  assign P1_U3246 = ~n11687 | ~n11686;
  assign n15278 = ~P1_REG3_REG_8__SCAN_IN | ~P1_U3086;
  assign n11688 = ~n15607 | ~P1_ADDR_REG_8__SCAN_IN;
  assign n11698 = ~n15278 | ~n11688;
  assign n11691 = n11690 ^ n11689;
  assign n11696 = ~n11691 | ~n15591;
  assign n11694 = n11693 ^ n11692;
  assign n11695 = ~n11694 | ~n15574;
  assign n11697 = ~n11696 | ~n11695;
  assign n11701 = ~n11698 & ~n11697;
  assign n11700 = ~n15604 | ~n11699;
  assign P1_U3251 = ~n11701 | ~n11700;
  assign n11704 = n11703 ^ n11702;
  assign n11716 = ~n15596 & ~n11704;
  assign n11709 = ~n11705;
  assign n11708 = ~n11707 | ~n11706;
  assign n11710 = ~n11709 | ~n11708;
  assign n11714 = ~n11710 | ~n15591;
  assign n15320 = ~P1_STATE_REG_SCAN_IN & ~n11711;
  assign n11712 = n15607 & P1_ADDR_REG_9__SCAN_IN;
  assign n11713 = ~n15320 & ~n11712;
  assign n11715 = ~n11714 | ~n11713;
  assign n11719 = ~n11716 & ~n11715;
  assign n11718 = ~n15604 | ~n11717;
  assign P1_U3252 = ~n11719 | ~n11718;
  assign n11727 = ~P1_REG3_REG_0__SCAN_IN | ~n15355;
  assign n15434 = ~n11721 ^ n11720;
  assign n11725 = ~n15434 & ~n15293;
  assign n15358 = ~n15319;
  assign n11723 = ~n15358 | ~n9310;
  assign n11722 = ~n15361 | ~n16173;
  assign n11724 = ~n11723 | ~n11722;
  assign n11726 = ~n11725 & ~n11724;
  assign P1_U3232 = ~n11727 | ~n11726;
  assign n11729 = ~n11323 | ~n11809;
  assign n12034 = ~n11730 | ~n11729;
  assign n11738 = ~P2_D_REG_6__SCAN_IN & ~P2_D_REG_7__SCAN_IN;
  assign n11736 = ~n11732 | ~n11731;
  assign n11734 = ~P2_D_REG_10__SCAN_IN & ~P2_D_REG_11__SCAN_IN;
  assign n11733 = ~P2_D_REG_12__SCAN_IN & ~P2_D_REG_13__SCAN_IN;
  assign n11735 = ~n11734 | ~n11733;
  assign n11737 = ~n11736 & ~n11735;
  assign n11754 = ~n11738 | ~n11737;
  assign n11740 = ~P2_D_REG_18__SCAN_IN & ~P2_D_REG_19__SCAN_IN;
  assign n11739 = ~P2_D_REG_20__SCAN_IN & ~P2_D_REG_21__SCAN_IN;
  assign n11744 = ~n11740 | ~n11739;
  assign n11742 = ~P2_D_REG_16__SCAN_IN & ~P2_D_REG_14__SCAN_IN;
  assign n11741 = ~P2_D_REG_15__SCAN_IN & ~P2_D_REG_17__SCAN_IN;
  assign n11743 = ~n11742 | ~n11741;
  assign n11752 = ~n11744 & ~n11743;
  assign n11746 = ~P2_D_REG_26__SCAN_IN & ~P2_D_REG_27__SCAN_IN;
  assign n11745 = ~P2_D_REG_28__SCAN_IN & ~P2_D_REG_31__SCAN_IN;
  assign n11750 = ~n11746 | ~n11745;
  assign n11748 = ~P2_D_REG_22__SCAN_IN & ~P2_D_REG_23__SCAN_IN;
  assign n11747 = ~P2_D_REG_24__SCAN_IN & ~P2_D_REG_25__SCAN_IN;
  assign n11749 = ~n11748 | ~n11747;
  assign n11751 = ~n11750 & ~n11749;
  assign n11753 = ~n11752 | ~n11751;
  assign n11759 = ~n11754 & ~n11753;
  assign n11756 = ~P2_D_REG_2__SCAN_IN & ~P2_D_REG_3__SCAN_IN;
  assign n11755 = ~P2_D_REG_4__SCAN_IN & ~P2_D_REG_5__SCAN_IN;
  assign n11757 = ~n11756 | ~n11755;
  assign n11758 = ~P2_D_REG_30__SCAN_IN & ~n11757;
  assign n11760 = ~n11759 | ~n11758;
  assign n11761 = ~P2_D_REG_29__SCAN_IN & ~n11760;
  assign n12552 = n11728 | n11761;
  assign n11764 = ~n12034 | ~n12552;
  assign n11763 = n11728 | P2_D_REG_1__SCAN_IN;
  assign n11762 = ~n17214 | ~n11809;
  assign n12585 = ~n11781;
  assign n12488 = n17232 | n11117;
  assign n11767 = ~n12488 & ~n17243;
  assign n11782 = ~n11767 | ~n17238;
  assign n11777 = ~n12585 & ~n11782;
  assign n12896 = ~n17243 | ~n11117;
  assign n12557 = ~n12887 | ~n12896;
  assign n11775 = n12557 & n12993;
  assign n11768 = ~n12552;
  assign n11769 = ~n11768 & ~n12034;
  assign n12583 = ~n11769 | ~n17349;
  assign n12575 = ~n17243 | ~n11770;
  assign n12895 = ~n12575;
  assign n11771 = n17452 & n12865;
  assign n11783 = n11771 & n11782;
  assign n11773 = ~n12583 | ~n12584;
  assign n11774 = n11773 & n11772;
  assign n11776 = ~n11775 | ~n11774;
  assign n11778 = ~n11777 & ~n11776;
  assign n11780 = ~P2_U3151 & ~n11778;
  assign n12997 = n17205 & n17350;
  assign n11779 = n11781 & n12997;
  assign n16601 = ~P2_STATE_REG_SCAN_IN | ~n16618;
  assign n11799 = ~P2_REG3_REG_0__SCAN_IN | ~n16601;
  assign n11795 = ~n11781 & ~n17348;
  assign n12581 = ~n11782;
  assign n11786 = ~n11795 | ~n12581;
  assign n11784 = ~n11783 | ~n17350;
  assign n11785 = n12583 | n11784;
  assign n11789 = ~n12184 | ~n9288;
  assign n11788 = ~n12179 | ~n11787;
  assign n17195 = ~n11789 | ~n11788;
  assign n17171 = ~n17167 | ~n17195;
  assign n11790 = n17167 | n17195;
  assign n17358 = n17171 & n11790;
  assign n11794 = ~n16595 | ~n17358;
  assign n11791 = ~n17185 | ~n17350;
  assign n11792 = n12583 | n11791;
  assign n13492 = ~n17452 & ~n12575;
  assign n11793 = ~n16616 | ~n17195;
  assign n11797 = ~n11794 | ~n11793;
  assign n12335 = ~n11795 | ~n17205;
  assign n12544 = ~n12051 ^ n11273;
  assign n17204 = ~n17151;
  assign n11796 = ~n16542 & ~n17204;
  assign n11798 = ~n11797 & ~n11796;
  assign P2_U3172 = ~n11799 | ~n11798;
  assign n11801 = ~n12296;
  assign n16134 = ~n16154;
  assign n11808 = ~n11801 | ~n16134;
  assign n11803 = ~n11802;
  assign n11806 = ~n11803 & ~P1_U3086;
  assign n16023 = n11800 | P1_STATE_REG_SCAN_IN;
  assign n11805 = ~n16023 & ~n11804;
  assign n11807 = ~n11806 & ~n11805;
  assign P1_U3329 = ~n11808 | ~n11807;
  assign n11813 = ~n12296 & ~n17341;
  assign n11811 = n11809 | P2_U3151;
  assign n11810 = ~n17338 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n11812 = ~n11811 | ~n11810;
  assign P2_U3269 = n11813 | n11812;
  assign n11819 = ~n12311;
  assign n11818 = ~n11819 | ~n16134;
  assign n11816 = ~n15386 & ~P1_U3086;
  assign n11815 = ~n16023 & ~n11814;
  assign n11817 = ~n11816 & ~n11815;
  assign P1_U3328 = ~n11818 | ~n11817;
  assign n11824 = ~n11819 | ~n11830;
  assign n11820 = ~P1_DATAO_REG_27__SCAN_IN;
  assign n11821 = ~n17226 & ~n11820;
  assign n11823 = ~n11822 & ~n11821;
  assign P2_U3268 = ~n11824 | ~n11823;
  assign n11831 = ~n12345;
  assign n11829 = ~n11831 | ~n16134;
  assign n11827 = ~n15431 & ~P1_U3086;
  assign n11826 = ~n16023 & ~n11825;
  assign n11828 = ~n11827 & ~n11826;
  assign P1_U3327 = ~n11829 | ~n11828;
  assign n11835 = ~n11831 | ~n11830;
  assign n11832 = n17338 & P1_DATAO_REG_28__SCAN_IN;
  assign n11834 = ~n11833 & ~n11832;
  assign P2_U3267 = ~n11835 | ~n11834;
  assign n17573 = ~P2_ADDR_REG_18__SCAN_IN | ~P1_ADDR_REG_18__SCAN_IN;
  assign n17578 = ~P2_ADDR_REG_17__SCAN_IN & ~P1_ADDR_REG_17__SCAN_IN;
  assign n17577 = P2_ADDR_REG_17__SCAN_IN & P1_ADDR_REG_17__SCAN_IN;
  assign n17582 = ~P2_ADDR_REG_16__SCAN_IN & ~P1_ADDR_REG_16__SCAN_IN;
  assign n17581 = P2_ADDR_REG_16__SCAN_IN & P1_ADDR_REG_16__SCAN_IN;
  assign n17586 = ~P2_ADDR_REG_15__SCAN_IN & ~P1_ADDR_REG_15__SCAN_IN;
  assign n17585 = P2_ADDR_REG_15__SCAN_IN & P1_ADDR_REG_15__SCAN_IN;
  assign n17590 = ~P2_ADDR_REG_14__SCAN_IN & ~P1_ADDR_REG_14__SCAN_IN;
  assign n17589 = P2_ADDR_REG_14__SCAN_IN & P1_ADDR_REG_14__SCAN_IN;
  assign n17594 = ~P2_ADDR_REG_13__SCAN_IN & ~P1_ADDR_REG_13__SCAN_IN;
  assign n17593 = P2_ADDR_REG_13__SCAN_IN & P1_ADDR_REG_13__SCAN_IN;
  assign n17598 = ~P2_ADDR_REG_12__SCAN_IN & ~P1_ADDR_REG_12__SCAN_IN;
  assign n17597 = P2_ADDR_REG_12__SCAN_IN & P1_ADDR_REG_12__SCAN_IN;
  assign n17602 = ~P2_ADDR_REG_11__SCAN_IN & ~P1_ADDR_REG_11__SCAN_IN;
  assign n17601 = P2_ADDR_REG_11__SCAN_IN & P1_ADDR_REG_11__SCAN_IN;
  assign n17606 = ~P2_ADDR_REG_10__SCAN_IN & ~P1_ADDR_REG_10__SCAN_IN;
  assign n17605 = P2_ADDR_REG_10__SCAN_IN & P1_ADDR_REG_10__SCAN_IN;
  assign n11854 = ~P2_ADDR_REG_9__SCAN_IN & ~P1_ADDR_REG_9__SCAN_IN;
  assign n11852 = ~P2_ADDR_REG_8__SCAN_IN & ~P1_ADDR_REG_8__SCAN_IN;
  assign n11850 = ~P2_ADDR_REG_7__SCAN_IN & ~P1_ADDR_REG_7__SCAN_IN;
  assign n11848 = ~P2_ADDR_REG_6__SCAN_IN & ~P1_ADDR_REG_6__SCAN_IN;
  assign n11846 = ~P2_ADDR_REG_5__SCAN_IN & ~P1_ADDR_REG_5__SCAN_IN;
  assign n11844 = ~P2_ADDR_REG_4__SCAN_IN & ~P1_ADDR_REG_4__SCAN_IN;
  assign n11842 = ~P1_ADDR_REG_3__SCAN_IN | ~P2_ADDR_REG_3__SCAN_IN;
  assign n17570 = P1_ADDR_REG_3__SCAN_IN ^ P2_ADDR_REG_3__SCAN_IN;
  assign n11840 = ~P1_ADDR_REG_2__SCAN_IN | ~P2_ADDR_REG_2__SCAN_IN;
  assign n11836 = ~P1_ADDR_REG_0__SCAN_IN | ~P2_ADDR_REG_0__SCAN_IN;
  assign n17555 = n11837 & n11836;
  assign n17554 = ~n11837 & ~n11836;
  assign n11838 = ~P2_ADDR_REG_1__SCAN_IN & ~n17554;
  assign n17572 = ~n17555 & ~n11838;
  assign n17571 = P1_ADDR_REG_2__SCAN_IN ^ P2_ADDR_REG_2__SCAN_IN;
  assign n11839 = ~n17572 | ~n17571;
  assign n17569 = ~n11840 | ~n11839;
  assign n11841 = ~n17570 | ~n17569;
  assign n17568 = ~n11842 | ~n11841;
  assign n17567 = ~P2_ADDR_REG_4__SCAN_IN ^ P1_ADDR_REG_4__SCAN_IN;
  assign n11843 = ~n17568 & ~n17567;
  assign n17566 = ~n11844 & ~n11843;
  assign n17565 = ~P2_ADDR_REG_5__SCAN_IN ^ P1_ADDR_REG_5__SCAN_IN;
  assign n11845 = ~n17566 & ~n17565;
  assign n17563 = ~P2_ADDR_REG_6__SCAN_IN ^ P1_ADDR_REG_6__SCAN_IN;
  assign n17561 = ~P2_ADDR_REG_7__SCAN_IN ^ P1_ADDR_REG_7__SCAN_IN;
  assign n17559 = ~P2_ADDR_REG_8__SCAN_IN ^ P1_ADDR_REG_8__SCAN_IN;
  assign n17557 = ~P2_ADDR_REG_9__SCAN_IN ^ P1_ADDR_REG_9__SCAN_IN;
  assign n11855 = ~n17605 & ~n17608;
  assign n11856 = ~n17601 & ~n17604;
  assign n11857 = ~n17597 & ~n17600;
  assign n11858 = ~n17593 & ~n17596;
  assign n17592 = ~n17594 & ~n11858;
  assign n11859 = ~n17589 & ~n17592;
  assign n17588 = ~n17590 & ~n11859;
  assign n11860 = ~n17585 & ~n17588;
  assign n17584 = ~n17586 & ~n11860;
  assign n11861 = ~n17581 & ~n17584;
  assign n17580 = ~n17582 & ~n11861;
  assign n11862 = ~n17577 & ~n17580;
  assign n17575 = ~n17578 & ~n11862;
  assign n17574 = P2_ADDR_REG_18__SCAN_IN | P1_ADDR_REG_18__SCAN_IN;
  assign n11863 = ~n17575 | ~n17574;
  assign n11865 = ~n17573 | ~n11863;
  assign n11864 = ~P2_ADDR_REG_19__SCAN_IN ^ P1_ADDR_REG_19__SCAN_IN;
  assign ADD_1068_U4 = ~n11865 ^ n11864;
  assign n11867 = ~n11866;
  assign n11871 = ~n13271 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n11870 = ~n11800 | ~P2_DATAO_REG_29__SCAN_IN;
  assign n12839 = ~n11871 | ~n11870;
  assign n11872 = ~n12484;
  assign n11877 = ~n11872 | ~n16134;
  assign n11875 = ~n11873 & ~P1_U3086;
  assign n12405 = ~P2_DATAO_REG_29__SCAN_IN;
  assign n11874 = ~n16023 & ~n12405;
  assign n11876 = ~n11875 & ~n11874;
  assign P1_U3326 = ~n11877 | ~n11876;
  assign n11882 = ~n12484 & ~n17341;
  assign n11880 = ~n11878 | ~P2_STATE_REG_SCAN_IN;
  assign n11879 = ~n17338 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n11881 = ~n11880 | ~n11879;
  assign P2_U3266 = n11882 | n11881;
  assign n11886 = ~n11884 & ~n11883;
  assign n11885 = ~n11886 & ~n16817;
  assign n11892 = ~n11885 & ~n11888;
  assign n11887 = ~n11886;
  assign n11890 = ~n11887 & ~n17550;
  assign n11889 = ~n16949 | ~n11888;
  assign n11891 = ~n11890 & ~n11889;
  assign n11895 = ~n11892 & ~n11891;
  assign n13678 = ~P2_REG3_REG_18__SCAN_IN | ~P2_U3151;
  assign n11893 = ~n16945 | ~P2_ADDR_REG_18__SCAN_IN;
  assign n11894 = ~n13678 | ~n11893;
  assign n11900 = ~n11899 ^ n11898;
  assign n11902 = ~n11910 | ~P1_U3973;
  assign n11901 = ~n11337 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P1_U3556 = ~n11902 | ~n11901;
  assign n13352 = ~n12402 | ~n12398;
  assign n13319 = ~n13354 | ~n13352;
  assign n11904 = n11903 | n16216;
  assign n15908 = ~n11910 & ~n16193;
  assign n15890 = ~n13286 | ~n15908;
  assign n15966 = ~n15980 | ~n16173;
  assign n15907 = ~n15969 | ~n11907;
  assign n13393 = ~n11910 | ~n15930;
  assign n11911 = ~n11903 | ~n16216;
  assign n15723 = ~n15844 | ~n13065;
  assign n11912 = ~n15842 | ~n15819;
  assign n15814 = ~n15876 & ~n16227;
  assign n11914 = ~n15819 | ~n15814;
  assign n15801 = ~n15844;
  assign n11913 = ~n15801 | ~n13065;
  assign n11915 = ~n11914 | ~n11913;
  assign n11917 = ~n11964 | ~n15785;
  assign n11963 = ~n15785;
  assign n11916 = ~n15823 | ~n11963;
  assign n15795 = ~n11917 | ~n11916;
  assign n11918 = ~n11917;
  assign n13075 = ~n16258 | ~n15729;
  assign n11968 = ~n16271 | ~n15771;
  assign n14399 = ~n15771;
  assign n13294 = ~n15737 | ~n14399;
  assign n11919 = ~n15737 & ~n15771;
  assign n15318 = ~n15734;
  assign n15677 = ~n16279 | ~n15318;
  assign n11922 = ~n9297 | ~n15711;
  assign n11924 = ~n9563 | ~n9305;
  assign n11925 = ~n15637 | ~n14455;
  assign n11926 = ~n16315 | ~n15661;
  assign n11927 = ~n11997 | ~n15012;
  assign n11928 = ~n9555 | ~n15640;
  assign n11930 = ~n15178 | ~n15618;
  assign n11932 = ~n15167 | ~n13151;
  assign n11934 = ~n15157 | ~n11977;
  assign n14937 = ~n11935 | ~n11934;
  assign n11936 = ~n14610 | ~n14972;
  assign n15146 = ~n14610;
  assign n11937 = ~n15146 | ~n16388;
  assign n14951 = ~n16391;
  assign n11938 = ~n14924 | ~n14951;
  assign n11939 = ~n15135 | ~n16391;
  assign n14866 = ~n16394;
  assign n11941 = ~n9573 | ~n14866;
  assign n11942 = ~n15124 | ~n16394;
  assign n11944 = ~n15113 | ~n16397;
  assign n11945 = ~n9570 | ~n14865;
  assign n11946 = ~n15102 | ~n16400;
  assign n14813 = ~n11947 | ~n11946;
  assign n11950 = ~n14813 | ~n11948;
  assign n11949 = ~n15092 | ~n16403;
  assign n14792 = ~n11950 | ~n11949;
  assign n11951 = ~n14802 | ~n14817;
  assign n11952 = ~n15082 | ~n16406;
  assign n11954 = ~n15071 | ~n16409;
  assign n11956 = ~n15061 | ~n16412;
  assign n11957 = ~n15052 & ~n16415;
  assign n12379 = n13319 ^ n12401;
  assign n15998 = n11958 & n13008;
  assign n11960 = n16029 & n13477;
  assign n11961 = ~n10531 & ~n11960;
  assign n15983 = ~n15998 | ~n11961;
  assign n15853 = ~n15983 | ~n14848;
  assign n12008 = ~n12379 | ~n15853;
  assign n15993 = ~n16173;
  assign n15904 = ~n13285;
  assign n13402 = ~n13047;
  assign n15790 = ~n15729;
  assign n15759 = ~n15790 | ~n16258;
  assign n11966 = ~n15725 | ~n13294;
  assign n11965 = ~n15722;
  assign n11967 = ~n11966 & ~n11965;
  assign n15757 = ~n16258;
  assign n15760 = ~n15757 | ~n15729;
  assign n11969 = ~n11971 | ~n13292;
  assign n13076 = ~n15823 | ~n15785;
  assign n11970 = n15723 & n13076;
  assign n13409 = ~n11971 | ~n11970;
  assign n11972 = ~n13412 | ~n13409;
  assign n13298 = ~n9297 | ~n14457;
  assign n13416 = n13298 & n15677;
  assign n13426 = ~n15637 | ~n15661;
  assign n13427 = ~n11997 | ~n15640;
  assign n15009 = ~n11974 | ~n13136;
  assign n13432 = ~n15024 | ~n15618;
  assign n11975 = ~n15009 | ~n13432;
  assign n14946 = ~n14961 | ~n11977;
  assign n13310 = ~n14924 | ~n16391;
  assign n11978 = n14909 & n13310;
  assign n13438 = ~n13310;
  assign n14935 = ~n15146 | ~n14972;
  assign n11979 = n13438 | n14935;
  assign n13446 = ~n15135 | ~n14951;
  assign n13325 = ~n14889 | ~n13448;
  assign n13326 = ~n15113 | ~n14891;
  assign n14861 = ~n13327 | ~n13326;
  assign n13330 = ~n15102 | ~n14865;
  assign n13338 = n15092 | n14839;
  assign n14814 = ~n13338 | ~n13336;
  assign n11980 = ~n14814;
  assign n14768 = ~n14802 | ~n16406;
  assign n13341 = ~n15082 | ~n14817;
  assign n14793 = ~n14768 | ~n13341;
  assign n13455 = ~n15071 | ~n14622;
  assign n11983 = ~n13455;
  assign n14743 = n14793 | n11983;
  assign n13346 = ~n15061 | ~n14773;
  assign n11982 = n13343 & n14768;
  assign n11984 = ~n13349;
  assign n13460 = ~n13236;
  assign n11986 = ~n14730 | ~n13460;
  assign n13351 = ~n13242;
  assign n11989 = n13319 ^ n12409;
  assign n11988 = ~n10531 | ~n13484;
  assign n11987 = ~n13376 | ~n13477;
  assign n11995 = ~n11989 | ~n15977;
  assign n15933 = ~n11990;
  assign n11993 = ~n9756 & ~n15933;
  assign n15979 = ~n11991 & ~n15431;
  assign n15875 = ~n15979;
  assign n11992 = ~n14625 & ~n15875;
  assign n11994 = ~n11993 & ~n11992;
  assign n12383 = ~n11995 | ~n11994;
  assign n15931 = ~n16182 & ~n16173;
  assign n15924 = ~n15931 | ~n15930;
  assign n11996 = ~n15882 | ~n16202;
  assign n14921 = ~n14938 | ~n14610;
  assign n11999 = ~n11998 | ~n12402;
  assign n16327 = n16174 & n13382;
  assign n12000 = ~n11999 | ~n16327;
  assign n12381 = n14703 | n12000;
  assign n12005 = ~n12381 & ~n10531;
  assign n15927 = ~n15902;
  assign n12003 = ~n12402 | ~n15927;
  assign n16000 = ~n15917;
  assign n12002 = ~n16000 | ~n12001;
  assign n12004 = ~n12003 | ~n12002;
  assign n12007 = ~n12383 & ~n12006;
  assign n12016 = ~n12008 | ~n12007;
  assign n12011 = ~n12010 & ~n12009;
  assign n12389 = ~P1_STATE_REG_SCAN_IN | ~n12011;
  assign n12014 = ~n12389;
  assign n12386 = ~n12012;
  assign n12013 = ~n12386 & ~n12392;
  assign n12015 = ~n12014 | ~n12013;
  assign n12018 = ~n12016 | ~n16004;
  assign n15961 = ~n16004;
  assign n12017 = ~n15961 | ~P1_REG2_REG_28__SCAN_IN;
  assign P1_U3265 = ~n12018 | ~n12017;
  assign n12022 = ~n12021 | ~n12020;
  assign n12033 = ~n12022 | ~n15376;
  assign n12031 = ~n14721 & ~n15333;
  assign n12029 = ~n15311 | ~n14722;
  assign n12025 = n15319 | n12398;
  assign n12024 = P1_STATE_REG_SCAN_IN | n12023;
  assign n12027 = ~n12025 | ~n12024;
  assign n12026 = ~n15332 & ~n14773;
  assign n12028 = ~n12027 & ~n12026;
  assign n12030 = ~n12029 | ~n12028;
  assign n12032 = ~n12031 & ~n12030;
  assign P1_U3214 = ~n12033 | ~n12032;
  assign n12035 = ~n12034;
  assign n12036 = ~n12035 | ~n17238;
  assign n12536 = ~n17243;
  assign n12038 = ~n12036 | ~n12536;
  assign n12037 = ~n17238 | ~n17243;
  assign n12039 = ~n9342;
  assign n12040 = ~n8884 | ~n12039;
  assign n12047 = n12051 | n12040;
  assign n12041 = ~P1_DATAO_REG_1__SCAN_IN;
  assign n12042 = n11800 & n12041;
  assign n12045 = ~n11273 & ~n12042;
  assign n12044 = n11800 | n12043;
  assign n12046 = ~n12045 | ~n12044;
  assign n12049 = n17342 | n11800;
  assign n12048 = ~n11800 | ~P1_DATAO_REG_1__SCAN_IN;
  assign n12050 = ~n12049 | ~n12048;
  assign n12052 = n12348 | n17195;
  assign n17353 = ~n17195;
  assign n16495 = n17174 & n12052;
  assign n12054 = n12053 | n17151;
  assign n16594 = ~n12055 | ~n12054;
  assign n12060 = ~n12848 | ~P1_DATAO_REG_2__SCAN_IN;
  assign n12058 = ~n12847 & ~n12056;
  assign n12057 = ~n12179 & ~n9360;
  assign n12059 = ~n12058 & ~n12057;
  assign n12061 = ~n12348 ^ n16590;
  assign n16593 = ~n12061 ^ n17168;
  assign n12062 = ~n12061;
  assign n12063 = n12062 | n17168;
  assign n12065 = ~n12184 | ~n12064;
  assign n16141 = ~n12066;
  assign n12067 = ~n12348 ^ n16466;
  assign n12070 = n12067 | n16543;
  assign n12068 = ~n12067;
  assign n12069 = n12068 | n17150;
  assign n16460 = ~n12070 | ~n12069;
  assign n12074 = ~n12205 & ~n12071;
  assign n12073 = ~n12179 & ~n12072;
  assign n12076 = ~n12074 & ~n12073;
  assign n12075 = ~n8882 | ~n16135;
  assign n17389 = n12076 & n12075;
  assign n12082 = ~n12348 ^ n17389;
  assign n16538 = ~n12082 ^ n17132;
  assign n12079 = ~n12848 | ~P1_DATAO_REG_5__SCAN_IN;
  assign n12078 = ~n12184 | ~n12077;
  assign n12081 = n12079 & n12078;
  assign n12080 = ~n16127 | ~n12263;
  assign n12084 = ~n12348 ^ n16522;
  assign n16531 = ~n12084 ^ n17102;
  assign n12083 = ~n16531;
  assign n16528 = n12082 | n17132;
  assign n12085 = ~n12084;
  assign n12087 = ~P1_DATAO_REG_6__SCAN_IN;
  assign n12089 = ~n12205 & ~n12087;
  assign n12088 = ~n12179 & ~n17319;
  assign n12092 = ~n12089 & ~n12088;
  assign n17318 = ~n12090;
  assign n12091 = ~n12090 | ~n12263;
  assign n17062 = ~n12092 | ~n12091;
  assign n12093 = ~n12348 ^ n17062;
  assign n12096 = n12093 | n12644;
  assign n12094 = ~n12093;
  assign n12095 = n12094 | n17078;
  assign n16608 = n12096 & n12095;
  assign n12101 = n17312 | n12847;
  assign n12097 = ~P1_DATAO_REG_7__SCAN_IN;
  assign n12099 = ~n12205 & ~n12097;
  assign n12098 = ~n12179 & ~n17313;
  assign n12100 = ~n12099 & ~n12098;
  assign n12119 = ~n12348 ^ n17414;
  assign n16477 = ~n12119 ^ n17053;
  assign n12106 = n17306 | n12847;
  assign n12102 = ~P1_DATAO_REG_8__SCAN_IN;
  assign n12104 = ~n12205 & ~n12102;
  assign n12103 = ~n17307 & ~n12179;
  assign n12105 = ~n12104 & ~n12103;
  assign n12118 = ~n12348 ^ n17422;
  assign n12107 = ~n12118;
  assign n12447 = ~n17036;
  assign n16485 = n12107 | n12447;
  assign n12120 = ~n16485;
  assign n16554 = n16477 | n12120;
  assign n12112 = n17300 | n12847;
  assign n12108 = ~P1_DATAO_REG_9__SCAN_IN;
  assign n12110 = ~n12205 & ~n12108;
  assign n12109 = ~n12179 & ~n17301;
  assign n12111 = ~n12110 & ~n12109;
  assign n16566 = ~n12112 | ~n12111;
  assign n12114 = ~n16566 ^ n12266;
  assign n12117 = ~n12114 | ~n17009;
  assign n12121 = ~n12117;
  assign n12113 = n16554 | n12121;
  assign n12115 = ~n12114;
  assign n16472 = ~n17009;
  assign n12116 = ~n12115 | ~n16472;
  assign n16557 = n12117 & n12116;
  assign n16479 = n12118 | n17036;
  assign n16478 = n12119 | n17053;
  assign n16483 = n16479 & n16478;
  assign n16556 = n12120 | n16483;
  assign n16560 = n16557 & n16556;
  assign n16444 = ~n12123 | ~n12122;
  assign n12132 = ~n16444 | ~n16573;
  assign n12124 = n16989 & n12122;
  assign n12130 = ~n12124 | ~n12123;
  assign n12125 = ~P1_DATAO_REG_10__SCAN_IN;
  assign n12127 = ~n12205 & ~n12125;
  assign n12126 = ~n12179 & ~n17295;
  assign n12128 = ~n12127 & ~n12126;
  assign n16445 = ~n16442 ^ n12348;
  assign n12131 = ~n12130 | ~n16445;
  assign n12137 = ~n16094 | ~n12263;
  assign n12133 = ~P1_DATAO_REG_11__SCAN_IN;
  assign n12135 = ~n12205 & ~n12133;
  assign n12134 = ~n12179 & ~n17289;
  assign n12136 = ~n12135 & ~n12134;
  assign n12138 = ~n17451 ^ n12348;
  assign n12139 = ~n12138;
  assign n12140 = n12139 | n14116;
  assign n16582 = ~n13638 | ~n12140;
  assign n12145 = ~n16087 | ~n12263;
  assign n12141 = ~P1_DATAO_REG_12__SCAN_IN;
  assign n12143 = ~n12205 & ~n12141;
  assign n12142 = ~n17283 & ~n12179;
  assign n12144 = ~n12143 & ~n12142;
  assign n12147 = ~n17463 ^ n12348;
  assign n13640 = n12147 | n13644;
  assign n12146 = n13640 & n13638;
  assign n12148 = ~n12147;
  assign n13639 = n12148 | n16974;
  assign n12153 = n17276 | n12847;
  assign n12149 = ~P1_DATAO_REG_13__SCAN_IN;
  assign n12151 = ~n12205 & ~n12149;
  assign n12150 = ~n17277 & ~n12179;
  assign n12152 = ~n12151 & ~n12150;
  assign n12155 = ~n14290 ^ n12348;
  assign n13636 = ~n12155 | ~n14050;
  assign n12154 = n13639 & n13636;
  assign n12156 = ~n12155;
  assign n13637 = ~n12156 | ~n17465;
  assign n12159 = ~n12848 | ~P1_DATAO_REG_14__SCAN_IN;
  assign n12158 = ~n16888 | ~n12184;
  assign n12160 = n12159 & n12158;
  assign n12162 = ~n12430 ^ n12348;
  assign n13504 = ~n12162 ^ n14291;
  assign n12164 = ~n13505 | ~n13504;
  assign n12163 = ~n12162;
  assign n12169 = ~n16068 | ~n8882;
  assign n12167 = ~n12165 | ~n12184;
  assign n12166 = ~n12848 | ~P1_DATAO_REG_15__SCAN_IN;
  assign n12168 = n12167 & n12166;
  assign n12170 = ~n14269 ^ n12348;
  assign n12171 = ~n12170;
  assign n12172 = n12171 | n14280;
  assign n13706 = n12173 & n12172;
  assign n12177 = n17259 | n12847;
  assign n12175 = n12179 | n17260;
  assign n12174 = ~n12848 | ~P1_DATAO_REG_16__SCAN_IN;
  assign n12176 = n12175 & n12174;
  assign n12196 = ~n14258 ^ n12266;
  assign n13585 = n12196 | n14270;
  assign n12183 = n17253 | n12847;
  assign n12178 = ~P1_DATAO_REG_18__SCAN_IN;
  assign n12181 = ~n12205 & ~n12178;
  assign n12180 = ~n12179 & ~n17254;
  assign n12182 = ~n12181 & ~n12180;
  assign n12190 = ~n13961 ^ n12348;
  assign n13674 = ~n12190 ^ n13926;
  assign n12195 = ~n13674;
  assign n12189 = ~n16054 | ~n12263;
  assign n12187 = ~n12185 | ~n12184;
  assign n12186 = ~n12848 | ~P1_DATAO_REG_17__SCAN_IN;
  assign n12188 = n12187 & n12186;
  assign n13589 = ~n14249 ^ n12266;
  assign n13672 = n13589 | n14259;
  assign n12194 = n12195 | n13672;
  assign n12192 = n13585 & n12194;
  assign n12191 = ~n12190;
  assign n12193 = n12191 | n13926;
  assign n12202 = ~n12193;
  assign n12200 = ~n12194;
  assign n13670 = n13589 & n14259;
  assign n12198 = ~n13670 & ~n12195;
  assign n12197 = ~n12196;
  assign n13587 = n12197 | n14032;
  assign n12199 = n12198 & n13587;
  assign n12201 = n12200 | n12199;
  assign n12209 = n17248 | n12847;
  assign n12204 = ~P1_DATAO_REG_19__SCAN_IN;
  assign n12207 = ~n12205 & ~n12204;
  assign n12206 = ~n12179 & ~n11117;
  assign n12208 = ~n12207 & ~n12206;
  assign n12210 = ~n14231 ^ n12348;
  assign n13530 = ~n12210 | ~n13951;
  assign n12212 = ~n13533 | ~n13530;
  assign n12211 = ~n12210;
  assign n13531 = ~n12211 | ~n13904;
  assign n12214 = ~n12848 | ~P1_DATAO_REG_20__SCAN_IN;
  assign n13621 = ~n14221 ^ n12266;
  assign n12218 = ~n12216 | ~P2_REG1_REG_20__SCAN_IN;
  assign n12217 = ~n12881 | ~P2_REG0_REG_20__SCAN_IN;
  assign n12225 = ~n12218 | ~n12217;
  assign n13910 = ~P2_REG3_REG_20__SCAN_IN ^ n12221;
  assign n12223 = ~n12219 | ~n13910;
  assign n12222 = ~n12327 | ~P2_REG2_REG_20__SCAN_IN;
  assign n12224 = ~n12223 | ~n12222;
  assign n12227 = ~n13621;
  assign n12228 = ~n12227 | ~n13932;
  assign n12230 = n17237 | n12847;
  assign n12229 = ~n12848 | ~P1_DATAO_REG_21__SCAN_IN;
  assign n13545 = ~n13895 ^ n12348;
  assign n12232 = ~n12303 | ~P2_REG1_REG_21__SCAN_IN;
  assign n12231 = ~n12881 | ~P2_REG0_REG_21__SCAN_IN;
  assign n12238 = ~n12232 | ~n12231;
  assign n13896 = ~P2_REG3_REG_21__SCAN_IN ^ n12244;
  assign n12236 = ~n11563 | ~n13896;
  assign n12235 = ~n12327 | ~P2_REG2_REG_21__SCAN_IN;
  assign n12237 = ~n12236 | ~n12235;
  assign n12239 = n13545 | n13909;
  assign n12241 = ~n16028 | ~n8882;
  assign n12240 = ~n12848 | ~P1_DATAO_REG_22__SCAN_IN;
  assign n13656 = ~n13871 ^ n12266;
  assign n12243 = ~n12303 | ~P2_REG1_REG_22__SCAN_IN;
  assign n12242 = ~n12881 | ~P2_REG0_REG_22__SCAN_IN;
  assign n12248 = ~n12243 | ~n12242;
  assign n13872 = ~P2_REG3_REG_22__SCAN_IN ^ n12255;
  assign n12246 = ~n11563 | ~n13872;
  assign n12245 = ~n12327 | ~P2_REG2_REG_22__SCAN_IN;
  assign n12247 = ~n12246 | ~n12245;
  assign n12250 = n13656 | n17522;
  assign n12249 = ~n13545;
  assign n13654 = n12249 | n17519;
  assign n12251 = ~n13656;
  assign n12252 = n12251 | n13886;
  assign n12254 = n17219 | n12847;
  assign n12253 = ~n12848 | ~P1_DATAO_REG_24__SCAN_IN;
  assign n13605 = n12348 ^ n14186;
  assign n13817 = ~n12289 ^ P2_REG3_REG_24__SCAN_IN;
  assign n12258 = ~n12303 | ~P2_REG1_REG_24__SCAN_IN;
  assign n12257 = ~n12881 | ~P2_REG0_REG_24__SCAN_IN;
  assign n12260 = ~n12258 | ~n12257;
  assign n12259 = n12327 & P2_REG2_REG_24__SCAN_IN;
  assign n12261 = ~n12260 & ~n12259;
  assign n12275 = ~n13605 | ~n17529;
  assign n12265 = ~n16021 | ~n12263;
  assign n12264 = ~n12848 | ~P1_DATAO_REG_23__SCAN_IN;
  assign n13602 = ~n14196 ^ n12266;
  assign n12273 = ~n13846 | ~n8889;
  assign n12269 = ~n12881 | ~P2_REG0_REG_23__SCAN_IN;
  assign n12268 = ~n12290 | ~P2_REG2_REG_23__SCAN_IN;
  assign n12271 = ~n12269 | ~n12268;
  assign n12270 = n12303 & P2_REG1_REG_23__SCAN_IN;
  assign n12272 = ~n12271 & ~n12270;
  assign n17525 = ~n12273 | ~n12272;
  assign n12274 = ~n13602 | ~n17525;
  assign n12276 = ~n12275 | ~n12274;
  assign n12279 = ~n13605;
  assign n12281 = ~n13602;
  assign n12277 = ~n12281 | ~n13862;
  assign n12278 = ~n12277 | ~n17529;
  assign n12283 = ~n12279 | ~n12278;
  assign n12280 = ~n17529 & ~n17525;
  assign n12282 = ~n12281 | ~n12280;
  assign n12284 = ~n12283 | ~n12282;
  assign n12286 = n17213 | n12847;
  assign n12285 = ~n12848 | ~P1_DATAO_REG_25__SCAN_IN;
  assign n12295 = n12348 ^ n14175;
  assign n12288 = ~n11531 | ~P2_REG1_REG_25__SCAN_IN;
  assign n12287 = ~n12881 | ~P2_REG0_REG_25__SCAN_IN;
  assign n12294 = ~n12288 | ~n12287;
  assign n13610 = ~P2_REG3_REG_24__SCAN_IN;
  assign n13792 = ~P2_REG3_REG_25__SCAN_IN ^ n12299;
  assign n12292 = ~n12219 | ~n13792;
  assign n12291 = ~n12290 | ~P2_REG2_REG_25__SCAN_IN;
  assign n12293 = ~n12292 | ~n12291;
  assign n13559 = ~n12295 ^ n17532;
  assign n12297 = ~n12848 | ~P1_DATAO_REG_26__SCAN_IN;
  assign n12308 = ~n14165 ^ n12348;
  assign n12300 = ~n12314;
  assign n13777 = ~P2_REG3_REG_26__SCAN_IN ^ n12300;
  assign n12302 = ~n13777 | ~n8889;
  assign n12301 = ~n12290 | ~P2_REG2_REG_26__SCAN_IN;
  assign n12307 = ~n12302 | ~n12301;
  assign n12305 = ~n12303 | ~P2_REG1_REG_26__SCAN_IN;
  assign n12304 = ~n12881 | ~P2_REG0_REG_26__SCAN_IN;
  assign n12306 = ~n12305 | ~n12304;
  assign n13688 = ~n12308 | ~n13801;
  assign n12310 = ~n13691 | ~n13688;
  assign n12309 = ~n12308;
  assign n13689 = ~n12309 | ~n17535;
  assign n12312 = ~n12848 | ~P1_DATAO_REG_27__SCAN_IN;
  assign n12353 = ~n14155 ^ n12348;
  assign n13695 = ~P2_REG3_REG_26__SCAN_IN;
  assign n12326 = ~n12314 | ~n13695;
  assign n13756 = ~P2_REG3_REG_27__SCAN_IN ^ n12326;
  assign n12315 = ~n12219 | ~n13756;
  assign n12317 = ~n12303 | ~P2_REG1_REG_27__SCAN_IN;
  assign n12316 = ~n12881 | ~P2_REG0_REG_27__SCAN_IN;
  assign n12318 = ~n12317 | ~n12316;
  assign n12349 = ~n12353 & ~n13776;
  assign n12319 = ~n12353;
  assign n12320 = ~n12319 & ~n17538;
  assign n12322 = ~n12349 & ~n12320;
  assign n12323 = ~n12321 & ~n16610;
  assign n12343 = ~n12323 | ~n12344;
  assign n12341 = ~n9510 & ~n13693;
  assign n12339 = ~n16577 | ~n13756;
  assign n12325 = ~n12303 | ~P2_REG1_REG_28__SCAN_IN;
  assign n12324 = ~n12881 | ~P2_REG0_REG_28__SCAN_IN;
  assign n12331 = ~n12325 | ~n12324;
  assign n13741 = ~P2_REG3_REG_28__SCAN_IN ^ n12358;
  assign n12329 = ~n12219 | ~n13741;
  assign n12328 = ~n12327 | ~P2_REG2_REG_28__SCAN_IN;
  assign n12330 = ~n12329 | ~n12328;
  assign n12931 = ~n17541;
  assign n12333 = n16542 | n12931;
  assign n12332 = ~P2_REG3_REG_27__SCAN_IN | ~P2_U3151;
  assign n12337 = ~n12333 | ~n12332;
  assign n12334 = ~n12544;
  assign n12336 = ~n16574 & ~n13801;
  assign n12338 = ~n12337 & ~n12336;
  assign n12340 = ~n12339 | ~n12338;
  assign n12342 = ~n12341 & ~n12340;
  assign P2_U3154 = ~n12343 | ~n12342;
  assign n12376 = ~n12344;
  assign n12347 = n12345 | n12847;
  assign n12346 = ~n12848 | ~P1_DATAO_REG_28__SCAN_IN;
  assign n12482 = ~n14146 | ~n17541;
  assign n12374 = ~n13739 ^ n12348;
  assign n12350 = ~n12349 & ~n16610;
  assign n12351 = ~n12374 | ~n12350;
  assign n12373 = ~n12376 & ~n12351;
  assign n12355 = ~n12374;
  assign n12352 = ~n16595 | ~n17538;
  assign n12354 = ~n12353 & ~n12352;
  assign n12371 = ~n12355 | ~n12354;
  assign n12854 = ~n14146;
  assign n12369 = ~n12854 & ~n13693;
  assign n12367 = ~n16577 | ~n13741;
  assign n12357 = n16574 | n13776;
  assign n12356 = ~P2_REG3_REG_28__SCAN_IN | ~P2_U3151;
  assign n12365 = ~n12357 | ~n12356;
  assign n12880 = ~n12219 | ~n12566;
  assign n12359 = ~n12290 | ~P2_REG2_REG_29__SCAN_IN;
  assign n12363 = ~n12880 | ~n12359;
  assign n12361 = ~n12303 | ~P2_REG1_REG_29__SCAN_IN;
  assign n12360 = ~n12881 | ~P2_REG0_REG_29__SCAN_IN;
  assign n12362 = ~n12361 | ~n12360;
  assign n12364 = ~n16542 & ~n13740;
  assign n12366 = ~n12365 & ~n12364;
  assign n12368 = ~n12367 | ~n12366;
  assign n12370 = ~n12369 & ~n12368;
  assign n12372 = ~n12371 | ~n12370;
  assign n12378 = ~n12373 & ~n12372;
  assign n12375 = ~n12374 & ~n16610;
  assign n12377 = ~n12376 | ~n12375;
  assign P2_U3160 = ~n12378 | ~n12377;
  assign n12385 = ~n12379 | ~n16225;
  assign n12380 = ~n12402 | ~n16329;
  assign n12382 = ~n12381 | ~n12380;
  assign n12384 = ~n12383 & ~n12382;
  assign n12395 = ~n12385 | ~n12384;
  assign n12387 = n16295 | n13376;
  assign n12388 = ~n12387 | ~n12386;
  assign n16383 = ~n12394 | ~n12392;
  assign n12391 = ~n12395 | ~n16385;
  assign n12390 = ~n16383 | ~P1_REG1_REG_28__SCAN_IN;
  assign P1_U3550 = ~n12391 | ~n12390;
  assign n12393 = ~n12392;
  assign n16326 = ~n12394 | ~n12393;
  assign n12397 = ~n12395 | ~n16338;
  assign n12396 = ~n16326 | ~P1_REG0_REG_28__SCAN_IN;
  assign P1_U3518 = ~n12397 | ~n12396;
  assign n12400 = ~n12399 | ~n12398;
  assign n12404 = ~n12401 | ~n12400;
  assign n12403 = ~n12402 | ~n16418;
  assign n12408 = ~n12404 | ~n12403;
  assign n12407 = ~n11872 | ~n10720;
  assign n12406 = n10193 | n12405;
  assign n13322 = ~n13012 ^ n16421;
  assign n13004 = ~n12408 ^ n13322;
  assign n12426 = ~n13004 | ~n16225;
  assign n12410 = ~n12409 | ~n13354;
  assign n12411 = ~n12410 | ~n13352;
  assign n12412 = ~n12411 ^ n13322;
  assign n12421 = ~n12412 | ~n15977;
  assign n12414 = ~n13264 | ~P1_REG2_REG_30__SCAN_IN;
  assign n12413 = ~n8891 | ~P1_REG1_REG_30__SCAN_IN;
  assign n12416 = n12414 & n12413;
  assign n12415 = ~n13263 | ~P1_REG0_REG_30__SCAN_IN;
  assign n16424 = n12416 & n12415;
  assign n12417 = ~n15432 | ~P1_B_REG_SCAN_IN;
  assign n14707 = ~n11990 | ~n12417;
  assign n12419 = n16424 | n14707;
  assign n12418 = ~n16418 | ~n15979;
  assign n12420 = n12419 & n12418;
  assign n13005 = ~n12421 | ~n12420;
  assign n13011 = ~n14703 ^ n13012;
  assign n12423 = ~n13011 | ~n16327;
  assign n12422 = ~n13012 | ~n16329;
  assign n12424 = ~n12423 | ~n12422;
  assign n12425 = ~n13005 & ~n12424;
  assign n12572 = ~n12426 | ~n12425;
  assign n12428 = ~n12572 | ~n16385;
  assign n12427 = ~n16383 | ~P1_REG1_REG_29__SCAN_IN;
  assign P1_U3551 = ~n12428 | ~n12427;
  assign n12492 = ~n14258;
  assign n12429 = ~n12492 | ~n14032;
  assign n12462 = ~n14258 | ~n14270;
  assign n12491 = ~n12430;
  assign n14084 = ~n14291;
  assign n14022 = ~n12491 | ~n14084;
  assign n12460 = ~n12431 & ~n14022;
  assign n14045 = ~n14290 | ~n17465;
  assign n12968 = ~n12430 | ~n14291;
  assign n14021 = n14045 & n12968;
  assign n12432 = ~n12431;
  assign n12433 = n12432 & n14021;
  assign n12461 = ~n13998 | ~n12435;
  assign n12437 = ~n17175 | ~n17171;
  assign n17184 = ~n17365;
  assign n12436 = n17151 | n17184;
  assign n12607 = ~n17168 | ~n17373;
  assign n17381 = ~n16466;
  assign n17098 = ~n16543 | ~n17381;
  assign n17095 = n17168 | n16590;
  assign n12439 = n17098 & n17095;
  assign n17111 = ~n17389;
  assign n17074 = n17132 | n17111;
  assign n12441 = n17102 | n16522;
  assign n12440 = n17074 & n12441;
  assign n12442 = ~n12441;
  assign n17082 = ~n12634 | ~n12636;
  assign n17406 = ~n17062;
  assign n12445 = n12644 & n17406;
  assign n17028 = n12644 | n17406;
  assign n17043 = ~n17414;
  assign n12499 = ~n17043 | ~n17053;
  assign n17004 = n17028 & n12499;
  assign n12959 = n17422 | n12447;
  assign n12446 = n17004 & n12959;
  assign n12449 = ~n12959;
  assign n12958 = ~n17422 | ~n12447;
  assign n17005 = ~n16473 | ~n17414;
  assign n12448 = n12958 & n17005;
  assign n12452 = n16566 & n17009;
  assign n16969 = n16442 | n16989;
  assign n17429 = ~n16566;
  assign n14124 = ~n17429 | ~n16472;
  assign n12453 = n16969 & n14124;
  assign n12454 = ~n17451 | ~n14116;
  assign n16967 = ~n16442 | ~n16989;
  assign n12455 = n12454 & n16967;
  assign n12456 = n17451 | n14116;
  assign n12457 = ~n17463 | ~n16974;
  assign n12459 = ~n14099 | ~n12457;
  assign n12458 = n17463 | n16974;
  assign n14020 = ~n14290 & ~n17465;
  assign n12901 = n14249 | n14008;
  assign n12903 = ~n14249 | ~n14008;
  assign n13969 = ~n12901 | ~n12903;
  assign n12463 = ~n14249 | ~n14259;
  assign n13945 = n13961 & n13926;
  assign n13944 = n13961 | n13926;
  assign n13923 = ~n13931 | ~n13951;
  assign n13922 = ~n14231 | ~n13904;
  assign n12909 = ~n14221 | ~n13932;
  assign n13918 = ~n12911 | ~n12909;
  assign n12915 = ~n13895 | ~n13909;
  assign n13883 = ~n12912 | ~n12915;
  assign n13856 = n13918 & n13883;
  assign n12799 = n13871 | n17522;
  assign n12465 = ~n12799;
  assign n12916 = ~n13871 | ~n13886;
  assign n13859 = ~n12919 | ~n12916;
  assign n12467 = n12465 | n13859;
  assign n12466 = n13856 & n12467;
  assign n12470 = ~n12467;
  assign n13881 = ~n13625 | ~n13932;
  assign n12468 = n13879 | n13881;
  assign n12763 = n13895 | n17519;
  assign n13857 = n12468 & n12763;
  assign n12469 = n13857 & n12799;
  assign n13810 = ~n14196 & ~n17525;
  assign n12779 = ~n13609 | ~n13837;
  assign n12474 = ~n12779;
  assign n12473 = n13810 | n12474;
  assign n13827 = ~n14196 | ~n13862;
  assign n13811 = ~n13835 | ~n14196;
  assign n12475 = n12474 | n13811;
  assign n12781 = ~n14186 | ~n17529;
  assign n12948 = ~n14175 | ~n17532;
  assign n12949 = n14175 | n17532;
  assign n13694 = ~n14165;
  assign n12477 = ~n13694 | ~n13801;
  assign n13751 = ~n14165 | ~n17535;
  assign n12478 = ~n14155 | ~n17538;
  assign n12479 = ~n12478;
  assign n12832 = ~n14155 | ~n13776;
  assign n13768 = ~n12831 | ~n12832;
  assign n12480 = n12479 | n13768;
  assign n12487 = ~n12483 | ~n12482;
  assign n12486 = n12484 | n12847;
  assign n12485 = ~n12848 | ~P1_DATAO_REG_29__SCAN_IN;
  assign n12490 = ~n12487 ^ n12985;
  assign n12489 = n17238 | n17243;
  assign n12551 = ~n12490 & ~n17356;
  assign n12733 = ~n14258 | ~n14032;
  assign n12493 = ~n12733;
  assign n12720 = n14269 | n14061;
  assign n14017 = ~n12491 | ~n14291;
  assign n12725 = ~n14269 | ~n14061;
  assign n13992 = ~n9809 | ~n12725;
  assign n12732 = ~n12492 | ~n14270;
  assign n13971 = ~n13969;
  assign n17142 = ~n17154;
  assign n12495 = ~n17175;
  assign n17177 = ~n12495 | ~n12494;
  assign n12615 = n16543 | n16466;
  assign n12496 = ~n17132 | ~n17389;
  assign n12498 = ~n17081 | ~n12634;
  assign n12642 = ~n12644 | ~n17062;
  assign n12643 = n12644 | n17062;
  assign n17030 = ~n17005 | ~n12499;
  assign n12667 = ~n17053 | ~n17414;
  assign n14090 = n17422 | n17036;
  assign n16992 = ~n16566 ^ n17009;
  assign n12960 = ~n16442 | ~n16573;
  assign n16961 = n16992 & n12960;
  assign n12684 = ~n17451 | ~n16507;
  assign n14093 = n16961 & n12684;
  assign n12500 = n14090 & n12506;
  assign n12505 = n14290 | n14050;
  assign n12962 = ~n12684;
  assign n12963 = ~n17451 & ~n16507;
  assign n12502 = ~n12963;
  assign n12501 = ~n12960;
  assign n14119 = ~n17429 | ~n17009;
  assign n12503 = n12502 & n16962;
  assign n12964 = n17463 | n13644;
  assign n12508 = n12505 & n14068;
  assign n12507 = ~n12506;
  assign n14091 = ~n17422 | ~n17036;
  assign n14066 = n12507 | n14091;
  assign n14042 = ~n14290 | ~n14050;
  assign n12708 = ~n12430 | ~n14084;
  assign n14016 = n14042 & n12708;
  assign n13991 = n14016 & n12725;
  assign n12510 = n13991 & n12733;
  assign n12512 = ~n12511 | ~n12898;
  assign n13947 = ~n12512 | ~n12903;
  assign n13974 = ~n13926;
  assign n12899 = n13961 | n13974;
  assign n12904 = ~n13961 | ~n13974;
  assign n12906 = n14231 & n13951;
  assign n12513 = ~n12906;
  assign n12900 = ~n13931 | ~n13904;
  assign n12975 = ~n13918;
  assign n13853 = ~n13859;
  assign n12515 = ~n12920;
  assign n12950 = ~n14186 | ~n13837;
  assign n12923 = n12950 & n13827;
  assign n12791 = n14175 | n13824;
  assign n13804 = ~n13609 | ~n17529;
  assign n12925 = n12791 & n13804;
  assign n12926 = ~n14175 | ~n13824;
  assign n13765 = ~n14165 | ~n13801;
  assign n12518 = n12832 & n13765;
  assign n12516 = ~n13739 | ~n12518;
  assign n12517 = n12985 | n12516;
  assign n12929 = ~n14146 & ~n12931;
  assign n12521 = n13739 | n12929;
  assign n13735 = ~n12518;
  assign n12519 = n13735 & n12831;
  assign n12531 = ~n12929;
  assign n12520 = ~n12519 | ~n12531;
  assign n12522 = ~n12521 | ~n12520;
  assign n12527 = n9417 | n12522;
  assign n13764 = n14165 | n13801;
  assign n12523 = n13735 | n13764;
  assign n13736 = ~n12523 | ~n12831;
  assign n12524 = ~n13736 | ~n13739;
  assign n12525 = ~n12524 | ~n12531;
  assign n12526 = n12985 | n12525;
  assign n12528 = ~n12527 | ~n12526;
  assign n12535 = ~n12529 | ~n12528;
  assign n12530 = n12831 & n13764;
  assign n12532 = n12531 & n12530;
  assign n12533 = n12985 & n12532;
  assign n12564 = ~n12535 & ~n12534;
  assign n12537 = ~n12536 | ~n17232;
  assign n12538 = n12537 & n11117;
  assign n12555 = ~n12538 | ~n17452;
  assign n17178 = ~n17083;
  assign n12549 = ~n12564 | ~n17178;
  assign n14049 = ~n12544 | ~n12887;
  assign n12547 = ~n12931 & ~n14049;
  assign n12539 = ~n12290 | ~P2_REG2_REG_30__SCAN_IN;
  assign n12543 = n12880 & n12539;
  assign n12541 = ~n12881 | ~P2_REG0_REG_30__SCAN_IN;
  assign n12540 = ~n12303 | ~P2_REG1_REG_30__SCAN_IN;
  assign n12542 = n12541 & n12540;
  assign n17203 = n12865 | n12544;
  assign n12545 = ~n12179 | ~P2_B_REG_SCAN_IN;
  assign n13718 = ~n17464 | ~n12545;
  assign n12546 = ~n17547 & ~n13718;
  assign n12548 = ~n12547 & ~n12546;
  assign n12550 = ~n12549 | ~n12548;
  assign n12554 = ~n12034 ^ n17349;
  assign n12553 = n12552 & n17350;
  assign n13495 = ~n17349;
  assign n12556 = n12555 | n17243;
  assign n13493 = ~n12556 | ~n8890;
  assign n13496 = n13493 & n12557;
  assign n12560 = ~n13495 | ~n13496;
  assign n12558 = ~n13493;
  assign n12559 = ~n12558 | ~n17349;
  assign n12561 = ~n12560 | ~n12559;
  assign n12565 = ~n13500 | ~n12561;
  assign n17209 = ~n17200;
  assign n12563 = ~n12580 | ~n17209;
  assign n12562 = n17209 | P2_REG2_REG_29__SCAN_IN;
  assign n12571 = ~n12563 | ~n12562;
  assign n17088 = n17238 | n12575;
  assign n17183 = ~n17088;
  assign n13983 = ~n17209 | ~n17183;
  assign n12569 = ~n12576 & ~n13983;
  assign n17123 = n12565 | n17147;
  assign n12567 = ~n12936 | ~n17196;
  assign n13720 = ~n17197 | ~n12566;
  assign n12568 = ~n12567 | ~n13720;
  assign n12570 = ~n12569 & ~n12568;
  assign P2_U3204 = ~n12571 | ~n12570;
  assign n12574 = ~n12572 | ~n16338;
  assign n12573 = ~n16326 | ~P1_REG0_REG_29__SCAN_IN;
  assign P1_U3519 = ~n12574 | ~n12573;
  assign n13000 = ~n17232;
  assign n17440 = n12575 | n13000;
  assign n12578 = ~n12576 & ~n17440;
  assign n12933 = ~n12936;
  assign n12577 = ~n12933 & ~n17452;
  assign n12579 = ~n12578 & ~n12577;
  assign n12582 = ~n17205 & ~n12581;
  assign n12587 = n12583 | n12582;
  assign n12586 = ~n12585 | ~n12584;
  assign n12588 = ~n12587 | ~n12586;
  assign n17460 = ~n12588 | ~n17350;
  assign n17472 = ~n17460;
  assign n12590 = ~n13501 | ~n17472;
  assign n12589 = ~n17460 | ~P2_REG0_REG_29__SCAN_IN;
  assign P2_U3456 = ~n12590 | ~n12589;
  assign n12592 = ~n12595 | ~n9800;
  assign n12591 = ~n12594 | ~n8890;
  assign n12593 = n12592 & n12591;
  assign n12604 = ~n17154 & ~n12593;
  assign n12597 = ~n17167 | ~n17353;
  assign n12596 = ~n12595 | ~n8890;
  assign n12598 = ~n12597 | ~n17232;
  assign n12989 = ~n17238;
  assign n12600 = ~n12598 | ~n12989;
  assign n12599 = ~n17174 | ~n17238;
  assign n12601 = ~n12600 | ~n12599;
  assign n12603 = ~n12602 | ~n12601;
  assign n12612 = ~n12604 | ~n12603;
  assign n12605 = n12623 & n8890;
  assign n12610 = ~n12606 | ~n12605;
  assign n12608 = n12607 & n9800;
  assign n12609 = ~n12608 | ~n12615;
  assign n12611 = ~n12610 | ~n12609;
  assign n12626 = ~n12612 | ~n12611;
  assign n12614 = n17132 | n8890;
  assign n12613 = ~n17389 | ~n8890;
  assign n12617 = ~n12614 | ~n12613;
  assign n12624 = ~n12617 | ~n17074;
  assign n12616 = n12624 & n12615;
  assign n12621 = ~n12626 | ~n12616;
  assign n12627 = ~n12617;
  assign n12618 = ~n17132;
  assign n12619 = ~n12627 | ~n12618;
  assign n12620 = n12619 & n12634;
  assign n12622 = ~n12621 | ~n12620;
  assign n12633 = ~n12622 | ~n8890;
  assign n12625 = n12624 & n12623;
  assign n12630 = ~n12626 | ~n12625;
  assign n12628 = ~n12627 | ~n17389;
  assign n12629 = n12628 & n12636;
  assign n12631 = ~n12630 | ~n12629;
  assign n12632 = ~n12631 | ~n12887;
  assign n12635 = n12642 & n12887;
  assign n12640 = ~n12635 | ~n12634;
  assign n12638 = ~n12643 | ~n8890;
  assign n12637 = ~n12636;
  assign n12639 = n12638 | n12637;
  assign n12641 = ~n12640 | ~n12639;
  assign n17059 = ~n12643 | ~n12642;
  assign n12646 = ~n12644 | ~n8890;
  assign n12645 = n17062 | n8890;
  assign n12647 = ~n12646 | ~n12645;
  assign n12648 = ~n17059 | ~n12647;
  assign n12649 = n12648 & n17030;
  assign n12651 = ~n17429 | ~n12887;
  assign n12650 = n17009 | n9800;
  assign n12663 = ~n12651 | ~n12650;
  assign n12655 = ~n12663 | ~n14124;
  assign n12653 = ~n14090 | ~n8890;
  assign n12652 = ~n14091 | ~n12887;
  assign n12654 = ~n12653 | ~n12652;
  assign n12669 = ~n12655 | ~n12654;
  assign n12656 = ~n12669;
  assign n12657 = n12663 | n17009;
  assign n12658 = ~n12657 | ~n12887;
  assign n12662 = ~n12658 & ~n12501;
  assign n12659 = ~n17005 | ~n16473;
  assign n12660 = ~n14090 | ~n12659;
  assign n12661 = ~n12656 | ~n12660;
  assign n12673 = ~n12662 | ~n12661;
  assign n12664 = n12663 | n16566;
  assign n12666 = ~n12664 | ~n8890;
  assign n12665 = ~n12961;
  assign n12671 = ~n12666 & ~n12665;
  assign n12668 = n12667 & n14091;
  assign n12670 = n12669 | n12668;
  assign n12672 = ~n12671 | ~n12670;
  assign n12674 = ~n12673 | ~n12672;
  assign n12679 = ~n12675 | ~n12674;
  assign n17442 = ~n16442;
  assign n12676 = ~n17442 | ~n12887;
  assign n12678 = ~n12676 | ~n12960;
  assign n12677 = n16989 | n8890;
  assign n12681 = n12963 | n9800;
  assign n12680 = ~n12684 | ~n12887;
  assign n12683 = n17451 | n8890;
  assign n12686 = ~n12684 | ~n12683;
  assign n12685 = ~n16507 | ~n12887;
  assign n12687 = ~n12686 | ~n12685;
  assign n12689 = n12692 | n12865;
  assign n12688 = ~n12964 | ~n8890;
  assign n12690 = ~n12689 | ~n12688;
  assign n12691 = ~n12964;
  assign n12694 = ~n12691 | ~n12887;
  assign n12693 = ~n12692 | ~n8890;
  assign n12703 = n12694 & n12693;
  assign n12698 = ~n12707 | ~n12703;
  assign n12695 = ~n14290;
  assign n12697 = ~n12695 | ~n8890;
  assign n12696 = ~n14050 | ~n12887;
  assign n12704 = n12697 & n12696;
  assign n12702 = ~n12698 | ~n12704;
  assign n12700 = ~n14290 | ~n9800;
  assign n12699 = n14050 | n9800;
  assign n12701 = ~n12700 | ~n12699;
  assign n12714 = ~n12702 | ~n12701;
  assign n12705 = ~n12703;
  assign n12706 = ~n12705 & ~n12704;
  assign n12712 = ~n12707 | ~n12706;
  assign n12710 = ~n14017 | ~n12865;
  assign n12709 = ~n12708 | ~n12892;
  assign n12711 = ~n12710 | ~n12709;
  assign n12713 = n12712 & n12711;
  assign n12719 = ~n12714 | ~n12713;
  assign n12716 = ~n12430 | ~n12865;
  assign n12715 = ~n14291 | ~n12892;
  assign n12717 = ~n12716 | ~n12715;
  assign n12718 = ~n12717 | ~n12968;
  assign n12723 = ~n12719 | ~n12718;
  assign n12722 = ~n12720 | ~n12865;
  assign n12721 = ~n12725 | ~n12892;
  assign n12727 = ~n12725 | ~n12724;
  assign n12726 = ~n14061 | ~n12892;
  assign n12728 = ~n12727 | ~n12726;
  assign n12730 = ~n12732 | ~n12865;
  assign n12729 = ~n12733 | ~n12892;
  assign n12731 = ~n12730 | ~n12729;
  assign n12735 = ~n12732 | ~n12892;
  assign n12734 = ~n12733 | ~n12865;
  assign n12736 = ~n12735 | ~n12734;
  assign n12738 = ~n14249 & ~n12865;
  assign n12737 = ~n14259 & ~n12892;
  assign n12739 = n12738 | n12737;
  assign n12742 = ~n14249 & ~n12892;
  assign n12741 = ~n14259 & ~n12865;
  assign n12743 = n12742 | n12741;
  assign n12745 = ~n12899 | ~n8890;
  assign n12744 = ~n12904 | ~n12892;
  assign n12746 = ~n12745 | ~n12744;
  assign n12748 = n13961 | n8890;
  assign n12747 = n13926 | n12887;
  assign n12749 = ~n12748 | ~n12747;
  assign n12750 = ~n12749 | ~n13944;
  assign n12752 = ~n12513 | ~n12892;
  assign n12751 = ~n12900 | ~n8890;
  assign n12755 = ~n14231 | ~n8890;
  assign n12754 = n13951 | n12865;
  assign n12756 = ~n12755 | ~n12754;
  assign n12757 = ~n12756 | ~n13922;
  assign n12759 = ~n12911 | ~n8890;
  assign n12758 = ~n12909 | ~n12887;
  assign n12760 = ~n12759 | ~n12758;
  assign n12762 = n13895 | n12865;
  assign n12761 = n17519 | n12887;
  assign n12772 = ~n12762 | ~n12761;
  assign n12767 = ~n12772 | ~n12763;
  assign n12765 = ~n12911 | ~n12887;
  assign n12764 = ~n12909 | ~n12865;
  assign n12766 = ~n12765 | ~n12764;
  assign n12768 = n12767 & n12766;
  assign n12770 = n13871 | n12865;
  assign n12769 = n17522 | n12887;
  assign n12798 = n12770 & n12769;
  assign n12771 = ~n13871 | ~n17522;
  assign n12776 = ~n12798 | ~n12771;
  assign n12774 = ~n12772;
  assign n12773 = ~n13895 | ~n17519;
  assign n12775 = ~n12774 | ~n12773;
  assign n12825 = n12776 & n12775;
  assign n12778 = ~n13609 | ~n12892;
  assign n12777 = ~n13837 | ~n12865;
  assign n12782 = n12778 & n12777;
  assign n12780 = ~n12782;
  assign n12803 = ~n12780 | ~n12779;
  assign n12787 = ~n12782 | ~n12781;
  assign n12783 = ~n14196 | ~n12892;
  assign n12785 = ~n12920 | ~n12783;
  assign n12784 = ~n17525 | ~n12892;
  assign n12786 = ~n12785 | ~n12784;
  assign n12788 = ~n12787 | ~n12786;
  assign n12818 = n12803 & n12788;
  assign n12789 = ~n12818;
  assign n12790 = n12825 & n12789;
  assign n12793 = ~n12791 | ~n12892;
  assign n12792 = ~n12926 | ~n12865;
  assign n12817 = ~n12793 | ~n12792;
  assign n12795 = ~n12831 | ~n12892;
  assign n12794 = ~n12832 | ~n8890;
  assign n12807 = ~n12795 | ~n12794;
  assign n12806 = n12817 & n12807;
  assign n12797 = ~n12920 | ~n12892;
  assign n12796 = ~n13827 | ~n12865;
  assign n12802 = ~n12797 | ~n12796;
  assign n12800 = ~n12798;
  assign n12801 = ~n12800 | ~n12799;
  assign n12804 = n12802 & n12801;
  assign n12828 = n12804 & n12803;
  assign n12814 = ~n12807;
  assign n12809 = n17535 | n12887;
  assign n12816 = n12809 & n12808;
  assign n12820 = ~n12816;
  assign n12811 = n14175 | n12887;
  assign n12810 = n17532 | n12865;
  assign n12812 = ~n12811 | ~n12810;
  assign n12819 = ~n12812 | ~n12949;
  assign n12813 = n12820 & n12819;
  assign n12815 = n12814 | n12813;
  assign n12827 = n12817 & n12816;
  assign n12821 = n12827 & n12818;
  assign n12823 = ~n14165 | ~n12865;
  assign n12822 = ~n17535 | ~n12892;
  assign n12824 = n12823 & n12822;
  assign n12830 = ~n12826 | ~n12825;
  assign n12829 = n12828 & n12827;
  assign n12834 = ~n12831 | ~n12865;
  assign n12833 = ~n12832 | ~n12892;
  assign n12835 = ~n12834 | ~n12833;
  assign n12837 = n14146 | n12887;
  assign n12836 = n17541 | n12865;
  assign n12859 = ~n12837 | ~n12836;
  assign n12840 = ~n12839;
  assign n12844 = ~n10438 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n12843 = ~n11800 | ~P2_DATAO_REG_30__SCAN_IN;
  assign n12845 = ~n12844 | ~n12843;
  assign n12870 = n12845 | SI_30_;
  assign n12846 = ~n12845 | ~SI_30_;
  assign n12868 = n12870 & n12846;
  assign n12850 = n15241 | n12847;
  assign n12849 = ~n12848 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n14141 = ~n12850 | ~n12849;
  assign n12939 = n14141 & n17547;
  assign n12851 = ~n12855 | ~n12936;
  assign n12852 = ~n12851 | ~n8890;
  assign n12853 = ~n12939 & ~n12852;
  assign n12856 = ~n12855 | ~n17544;
  assign n12857 = n12856 & n12887;
  assign n12947 = n14141 | n17547;
  assign n12858 = n12857 & n12947;
  assign n12861 = ~n12860 & ~n12859;
  assign n12984 = ~n12939;
  assign n12864 = n14141 | n12887;
  assign n12867 = ~n12984 | ~n12864;
  assign n12866 = ~n17547 | ~n12865;
  assign n12873 = ~n13271 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n12872 = ~n11800 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n12874 = ~n12873 | ~n12872;
  assign n12875 = ~n12874 ^ SI_31_;
  assign n12877 = n15232 | n11800;
  assign n12876 = ~n11800 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n12878 = ~n12877 | ~n12876;
  assign n12879 = ~n12327 | ~P2_REG2_REG_31__SCAN_IN;
  assign n12885 = ~n12880 | ~n12879;
  assign n12883 = ~n12303 | ~P2_REG1_REG_31__SCAN_IN;
  assign n12882 = ~n12881 | ~P2_REG0_REG_31__SCAN_IN;
  assign n12884 = ~n12883 | ~n12882;
  assign n12890 = ~n12944;
  assign n12886 = ~n14136 | ~n17551;
  assign n12986 = n12890 & n12886;
  assign n12888 = n17551 & n12887;
  assign n12889 = ~n14136 | ~n12888;
  assign n12891 = ~n12893;
  assign n12907 = ~n12900 | ~n12899;
  assign n12902 = ~n12901;
  assign n12972 = ~n12907 & ~n12902;
  assign n12905 = ~n12904 | ~n12903;
  assign n12970 = ~n12906 & ~n12905;
  assign n12908 = ~n12907 | ~n12513;
  assign n12913 = ~n12912 | ~n12911;
  assign n12917 = ~n12916 | ~n12915;
  assign n12922 = ~n12918 & ~n12917;
  assign n12921 = ~n12920 | ~n12919;
  assign n12927 = ~n12926;
  assign n12928 = ~n13735 & ~n12927;
  assign n12930 = ~n12929 & ~n13736;
  assign n12932 = ~n14146 | ~n12931;
  assign n12934 = ~n12933 | ~n17544;
  assign n12938 = ~n12935 | ~n12934;
  assign n12937 = ~n12936 | ~n13740;
  assign n12940 = ~n14141;
  assign n12941 = ~n12940 | ~n13719;
  assign n12942 = ~n14136 | ~n12941;
  assign n12943 = ~n14136 & ~n12947;
  assign n12945 = ~n12944 & ~n12943;
  assign n12983 = ~n12947;
  assign n12980 = ~n13768;
  assign n13806 = n12949 & n12948;
  assign n13829 = n13804 & n12950;
  assign n12952 = ~n17126 & ~n17175;
  assign n12951 = ~n17358 & ~n17154;
  assign n12953 = ~n12952 | ~n12951;
  assign n17107 = ~n17132 ^ n17389;
  assign n12955 = ~n12953 & ~n17107;
  assign n12954 = ~n17059 & ~n17082;
  assign n12957 = ~n12955 | ~n12954;
  assign n12956 = ~n17030;
  assign n17014 = ~n12959 | ~n12958;
  assign n14126 = ~n12961 | ~n12960;
  assign n16972 = n12963 | n12962;
  assign n12965 = n8986 | n16972;
  assign n14098 = ~n9344 | ~n12964;
  assign n12967 = ~n12965 & ~n14098;
  assign n12966 = ~n14020;
  assign n14071 = ~n12966 | ~n14045;
  assign n14024 = ~n14269 ^ n14061;
  assign n12974 = ~n12971 | ~n12970;
  assign n12973 = ~n12972;
  assign n12976 = ~n12974 & ~n12973;
  assign n12977 = ~n12976 | ~n12975;
  assign n12978 = ~n12977 & ~n13883;
  assign n12981 = ~n12980 | ~n12979;
  assign n13786 = ~n14165 ^ n13801;
  assign n12982 = ~n12981 & ~n13786;
  assign n12988 = ~n12987 | ~n12986;
  assign n12990 = ~n12988 ^ n11117;
  assign n12991 = ~n12990 & ~n12989;
  assign n12996 = ~n12995 & ~n12994;
  assign n12998 = ~n12997 | ~n12996;
  assign n13002 = ~n12998 | ~P2_B_REG_SCAN_IN;
  assign n17229 = ~n12999 | ~P2_STATE_REG_SCAN_IN;
  assign n13001 = ~n13000 & ~n17229;
  assign n13003 = ~n13002;
  assign n13021 = ~n13004 | ~n15896;
  assign n13006 = ~n16004 & ~P1_REG2_REG_29__SCAN_IN;
  assign n13019 = ~n13007 & ~n13006;
  assign n13010 = ~n13009 & ~n13008;
  assign n13017 = ~n13011 | ~n15991;
  assign n15023 = ~n16004 | ~n15927;
  assign n13015 = ~n14704 & ~n15023;
  assign n13014 = ~n15917 & ~n13013;
  assign n13016 = ~n13015 & ~n13014;
  assign n13018 = ~n13017 | ~n13016;
  assign n13020 = ~n13019 & ~n13018;
  assign P1_U3356 = ~n13021 | ~n13020;
  assign n13022 = ~n15930 | ~n13256;
  assign n13038 = ~n13023 | ~n13022;
  assign n13024 = ~n15930 | ~n13085;
  assign n13027 = n11905 | n13085;
  assign n13026 = ~n16202 | ~n13085;
  assign n13044 = ~n13027 | ~n13026;
  assign n13028 = ~n13044 | ~n15889;
  assign n13030 = ~n13401 | ~n8881;
  assign n13029 = ~n13398 | ~n13256;
  assign n13033 = ~n13031 | ~n13040;
  assign n13032 = n13398 | n9301;
  assign n13388 = ~n11906 | ~n13035;
  assign n13037 = ~n13036 | ~n13388;
  assign n13041 = ~n13039 | ~n13038;
  assign n15934 = ~n11905;
  assign n13043 = ~n13398 | ~n15934;
  assign n13046 = ~n13043 | ~n9323;
  assign n13045 = ~n13044;
  assign n13050 = ~n13046 | ~n13045;
  assign n13049 = ~n13047 | ~n13085;
  assign n13048 = ~n13406 | ~n9301;
  assign n13062 = ~n13052 | ~n13051;
  assign n13053 = ~n13401 & ~n13085;
  assign n13060 = ~n13054 | ~n13053;
  assign n13055 = n15876 | n13085;
  assign n13058 = ~n13406 | ~n13055;
  assign n13057 = ~n13056 | ~n9301;
  assign n13059 = ~n13058 | ~n13057;
  assign n13061 = n13060 & n13059;
  assign n13064 = ~n15722 | ~n13085;
  assign n13063 = ~n15723 | ~n9301;
  assign n13066 = ~n13065 | ~n13122;
  assign n13068 = ~n15722 | ~n13066;
  assign n13067 = n15844 | n9301;
  assign n13069 = ~n13068 | ~n13067;
  assign n13071 = ~n15763 | ~n8881;
  assign n13070 = ~n13076 | ~n9301;
  assign n13072 = ~n13071 | ~n13070;
  assign n13074 = n16258 | n13085;
  assign n13073 = n15729 | n13256;
  assign n13090 = n13074 & n13073;
  assign n13080 = ~n13090 | ~n13075;
  assign n13078 = ~n15763 | ~n9301;
  assign n13077 = ~n13076 | ~n13122;
  assign n13079 = ~n13078 | ~n13077;
  assign n13081 = n13080 & n13079;
  assign n13097 = ~n13082 | ~n13081;
  assign n13083 = ~n15677 | ~n13122;
  assign n13103 = ~n13084 | ~n13083;
  assign n13087 = ~n16271 | ~n13122;
  assign n13086 = n15771 | n13085;
  assign n13089 = ~n16271 | ~n9301;
  assign n13088 = n15771 | n13256;
  assign n13098 = ~n13089 | ~n13088;
  assign n13094 = ~n13099 | ~n13098;
  assign n13092 = ~n13090;
  assign n13093 = ~n13092 | ~n13091;
  assign n13095 = n13094 & n13093;
  assign n13096 = n13103 & n13095;
  assign n13101 = ~n13098;
  assign n13100 = ~n13099;
  assign n13102 = n13101 & n13100;
  assign n13109 = ~n13103 | ~n13102;
  assign n13104 = n15734 | n8881;
  assign n13107 = ~n13414 | ~n13104;
  assign n13106 = ~n13105 | ~n9301;
  assign n13108 = ~n13107 | ~n13106;
  assign n13114 = n13109 & n13108;
  assign n13110 = ~n16292 | ~n13122;
  assign n13112 = ~n13110 | ~n13298;
  assign n13111 = ~n14457 | ~n13122;
  assign n13113 = ~n13112 | ~n13111;
  assign n13115 = n13114 & n13113;
  assign n13117 = ~n13418 | ~n9301;
  assign n13116 = ~n13298 | ~n13122;
  assign n13118 = ~n13117 | ~n13116;
  assign n13120 = ~n13419 | ~n9301;
  assign n13119 = ~n13423 | ~n13122;
  assign n13121 = ~n15659 | ~n13122;
  assign n13124 = ~n13121 | ~n13423;
  assign n13123 = ~n14559 | ~n13122;
  assign n13125 = ~n13124 | ~n13123;
  assign n13130 = ~n13126 | ~n13125;
  assign n13128 = ~n13426 | ~n9301;
  assign n13127 = ~n13422 | ~n13122;
  assign n13129 = ~n13128 | ~n13127;
  assign n13135 = ~n13130 | ~n13129;
  assign n13132 = ~n13426 | ~n13122;
  assign n13131 = ~n13422 | ~n13256;
  assign n13133 = n13132 & n13131;
  assign n13141 = ~n13135 | ~n13134;
  assign n13430 = ~n13307 | ~n13136;
  assign n13139 = n13430 | n9301;
  assign n13137 = n13427 & n9301;
  assign n13138 = ~n13432 | ~n13137;
  assign n13140 = ~n13139 | ~n13138;
  assign n13145 = ~n13141 | ~n13140;
  assign n13144 = ~n13142 | ~n13307;
  assign n13143 = ~n14997 | ~n13122;
  assign n13147 = ~n13440 | ~n9301;
  assign n13146 = ~n13278 | ~n13122;
  assign n13150 = ~n9553 | ~n13122;
  assign n13153 = ~n13150 | ~n13278;
  assign n13152 = n13151 | n9301;
  assign n13154 = ~n13153 | ~n13152;
  assign n13156 = ~n8915 | ~n13122;
  assign n13155 = ~n14946 | ~n13256;
  assign n13157 = ~n14998 & ~n13256;
  assign n13158 = ~n15157 | ~n13122;
  assign n13160 = ~n13159 | ~n13158;
  assign n13165 = ~n13161 | ~n13160;
  assign n13163 = ~n14936 | ~n13256;
  assign n13162 = ~n14935 | ~n13122;
  assign n13164 = ~n13163 | ~n13162;
  assign n13170 = ~n13165 | ~n13164;
  assign n13166 = n14610 | n13122;
  assign n13168 = ~n13166 | ~n14936;
  assign n13167 = ~n16388 | ~n8896;
  assign n13169 = ~n13168 | ~n13167;
  assign n13178 = ~n13170 | ~n13169;
  assign n13172 = ~n13310 | ~n8896;
  assign n13171 = ~n13446 | ~n13122;
  assign n13176 = ~n13172 | ~n13171;
  assign n13175 = ~n13173 | ~n13122;
  assign n13174 = ~n13448 | ~n13256;
  assign n13177 = n13176 & n13179;
  assign n13186 = ~n13178 | ~n13177;
  assign n13180 = ~n15135 | ~n13256;
  assign n13182 = ~n13180 | ~n13310;
  assign n13181 = ~n16391 | ~n13256;
  assign n13185 = ~n13182 | ~n13181;
  assign n13183 = ~n15124 | ~n8896;
  assign n13184 = ~n16394 | ~n9301;
  assign n13188 = ~n13327 | ~n9301;
  assign n13187 = ~n13326 | ~n13122;
  assign n13189 = ~n13188 | ~n13187;
  assign n13195 = ~n13190 | ~n13189;
  assign n13191 = ~n15113 | ~n13256;
  assign n13193 = ~n13191 | ~n13327;
  assign n13192 = ~n16397 | ~n9301;
  assign n13194 = ~n13193 | ~n13192;
  assign n13197 = ~n13335 | ~n9301;
  assign n13196 = ~n13330 | ~n13122;
  assign n13199 = ~n14822 | ~n13256;
  assign n13198 = n16403 | n13256;
  assign n13201 = ~n13199 | ~n13198;
  assign n13206 = ~n16403 & ~n13122;
  assign n13200 = ~n14822 & ~n13206;
  assign n13204 = n13201 | n13200;
  assign n13203 = ~n13335 | ~n13122;
  assign n13202 = ~n13330 | ~n13256;
  assign n13208 = n14822 | n13122;
  assign n13207 = ~n13206;
  assign n13210 = n13208 & n13207;
  assign n13209 = ~n13336 | ~n13122;
  assign n13211 = ~n13210 | ~n13209;
  assign n13212 = n13341 & n13211;
  assign n13214 = ~n15082 | ~n13256;
  assign n13216 = ~n13214 | ~n14768;
  assign n13215 = ~n16406 | ~n9301;
  assign n13217 = ~n13216 | ~n13215;
  assign n13219 = ~n13343 | ~n9301;
  assign n13218 = ~n13455 | ~n13122;
  assign n13220 = ~n13219 | ~n13218;
  assign n13226 = ~n13221 | ~n13220;
  assign n13222 = n14778 | n13122;
  assign n13224 = ~n13222 | ~n13343;
  assign n13223 = ~n16409 | ~n9301;
  assign n13225 = ~n13224 | ~n13223;
  assign n13230 = ~n13226 | ~n13225;
  assign n13228 = ~n13349 | ~n8896;
  assign n13227 = ~n13346 | ~n13122;
  assign n13229 = ~n13228 | ~n13227;
  assign n13235 = ~n13230 | ~n13229;
  assign n13231 = n14756 | n13122;
  assign n13233 = ~n13231 | ~n13349;
  assign n13232 = ~n16412 | ~n9301;
  assign n13234 = ~n13233 | ~n13232;
  assign n13240 = ~n13235 | ~n13234;
  assign n13238 = n13236 | n13122;
  assign n13237 = n13242 | n13256;
  assign n13239 = ~n13238 | ~n13237;
  assign n13246 = ~n13240 | ~n13239;
  assign n13241 = ~n15052 & ~n13256;
  assign n13244 = n13242 | n13241;
  assign n13243 = n16415 | n9301;
  assign n13245 = ~n13244 | ~n13243;
  assign n13250 = ~n13246 | ~n13245;
  assign n13248 = ~n13354 | ~n13256;
  assign n13247 = ~n13352 | ~n13122;
  assign n13249 = ~n13248 | ~n13247;
  assign n13252 = ~n13354 | ~n13122;
  assign n13251 = ~n13352 | ~n9301;
  assign n13253 = ~n13252 | ~n13251;
  assign n13255 = ~n13254;
  assign n13257 = ~n8900 & ~n8939;
  assign n15243 = ~P2_DATAO_REG_30__SCAN_IN;
  assign n13260 = n10193 | n15243;
  assign n13262 = ~n15043 | ~n13256;
  assign n13266 = ~n13263 | ~P1_REG0_REG_31__SCAN_IN;
  assign n13265 = ~n13264 | ~P1_REG2_REG_31__SCAN_IN;
  assign n13268 = ~n13266 | ~n13265;
  assign n13267 = n8892 & P1_REG1_REG_31__SCAN_IN;
  assign n16427 = n13268 | n13267;
  assign n13275 = ~n16427;
  assign n13363 = ~n13275 & ~n16424;
  assign n13270 = ~n13363;
  assign n13272 = ~n10438 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n13274 = ~n13273 | ~n13272;
  assign n13324 = ~n15036 & ~n16427;
  assign n13276 = ~n13323 & ~n13324;
  assign n13277 = ~n13324 | ~n13256;
  assign n14746 = ~n13349 | ~n13346;
  assign n14770 = n13343 & n13455;
  assign n14862 = ~n14861;
  assign n13280 = ~n14935;
  assign n13279 = ~n8915 | ~n13278;
  assign n13435 = ~n13280 & ~n13279;
  assign n13281 = ~n13423;
  assign n15664 = ~n9678 & ~n13281;
  assign n13387 = n15980 & n15993;
  assign n16171 = n13282 | n13387;
  assign n13284 = ~n16171 & ~n13283;
  assign n15850 = ~n15842;
  assign n13291 = ~n13284 | ~n15850;
  assign n15893 = ~n13401 | ~n13398;
  assign n13289 = ~n15893 & ~n13285;
  assign n13287 = ~n15722 | ~n16034;
  assign n13288 = ~n13286 & ~n13287;
  assign n13290 = ~n13289 | ~n13288;
  assign n13293 = n13291 | n13290;
  assign n13295 = ~n13293 & ~n13292;
  assign n13296 = ~n13295 | ~n13294;
  assign n13297 = ~n13296 & ~n13409;
  assign n13299 = ~n13297 | ~n15709;
  assign n15680 = ~n13418 | ~n13298;
  assign n13300 = ~n13299 & ~n15680;
  assign n13304 = ~n15664 | ~n13300;
  assign n13302 = ~n13426;
  assign n13301 = ~n13422;
  assign n13303 = ~n15643 | ~n13440;
  assign n13306 = ~n13304 & ~n13303;
  assign n13305 = ~n15615;
  assign n15008 = ~n13432 | ~n13307;
  assign n13308 = ~n14909;
  assign n13311 = ~n13309 & ~n13308;
  assign n14911 = n13310 & n13446;
  assign n13312 = ~n13311 | ~n14911;
  assign n14888 = ~n13448 | ~n13173;
  assign n14836 = n13335 & n13330;
  assign n13315 = ~n13314 | ~n14836;
  assign n13316 = ~n14793 & ~n13315;
  assign n13317 = ~n14770 | ~n13316;
  assign n13318 = ~n14746 & ~n13317;
  assign n13320 = ~n14731 | ~n13318;
  assign n13321 = ~n13320 & ~n13319;
  assign n13474 = ~n13323;
  assign n13472 = ~n13324;
  assign n13334 = ~n13325 & ~n9665;
  assign n13328 = ~n13326 | ~n13173;
  assign n13329 = ~n13328 | ~n13327;
  assign n13332 = ~n13336 | ~n13329;
  assign n13331 = ~n13330;
  assign n13333 = ~n13332 & ~n13331;
  assign n13452 = ~n13341 | ~n13333;
  assign n13345 = ~n13334 & ~n13452;
  assign n13337 = ~n13335;
  assign n13339 = ~n13337 | ~n13336;
  assign n13340 = ~n13339 | ~n13338;
  assign n13342 = ~n13341 | ~n13340;
  assign n13344 = n13342 & n14768;
  assign n13386 = ~n13344 | ~n13343;
  assign n13348 = ~n13345 & ~n13386;
  assign n13347 = ~n13346 | ~n13455;
  assign n13350 = ~n13348 & ~n13347;
  assign n13385 = ~n13460 | ~n13349;
  assign n13353 = ~n13350 & ~n13385;
  assign n13463 = ~n13352 | ~n13351;
  assign n13356 = ~n13353 & ~n13463;
  assign n13355 = ~n14704 | ~n16421;
  assign n13466 = ~n13355 | ~n13354;
  assign n13358 = ~n13356 & ~n13466;
  assign n13357 = ~n15043 & ~n16427;
  assign n13362 = ~n13358 & ~n13357;
  assign n13359 = ~n16424;
  assign n13361 = ~n15043 & ~n13359;
  assign n13360 = ~n14704 & ~n16421;
  assign n13467 = ~n13361 & ~n13360;
  assign n13365 = ~n13362 | ~n13467;
  assign n13364 = ~n15043 | ~n13363;
  assign n13366 = ~n13365 | ~n13364;
  assign n13368 = ~n13366 | ~n13474;
  assign n13371 = ~n13368 | ~n13367;
  assign n13370 = ~n13369;
  assign n13372 = ~n13371 | ~n13370;
  assign n13373 = ~n13372 | ~n13472;
  assign n16044 = ~n10531;
  assign n13374 = ~n13373 | ~n16044;
  assign n13380 = ~n13375;
  assign n13378 = ~n13474 & ~n16044;
  assign n13377 = ~n16029 | ~n13376;
  assign n13379 = ~n13378 & ~n13377;
  assign n13381 = ~n13380 | ~n13379;
  assign n16039 = n13382 | P1_U3086;
  assign n13384 = ~n13383 & ~n16039;
  assign n13458 = ~n13385;
  assign n13454 = ~n13386;
  assign n13389 = ~n13387 & ~n16034;
  assign n13391 = ~n13389 | ~n13388;
  assign n13392 = ~n13391 | ~n13390;
  assign n13394 = n13392 | n15935;
  assign n13396 = ~n13394 | ~n13393;
  assign n13400 = ~n13396 | ~n13395;
  assign n13399 = n13398 & n13397;
  assign n13405 = ~n13400 | ~n13399;
  assign n13403 = ~n13401;
  assign n13404 = ~n13403 & ~n13402;
  assign n13407 = ~n13405 | ~n13404;
  assign n13408 = ~n13407 | ~n13406;
  assign n13411 = ~n13408 | ~n15722;
  assign n13410 = ~n13409;
  assign n13413 = ~n13411 | ~n13410;
  assign n13415 = ~n13413 | ~n13412;
  assign n13417 = ~n13415 | ~n13414;
  assign n13421 = n13417 & n13416;
  assign n13420 = ~n13419 | ~n13418;
  assign n13425 = ~n13421 & ~n13420;
  assign n13424 = ~n13423 | ~n13422;
  assign n13429 = ~n13425 & ~n13424;
  assign n13428 = ~n13427 | ~n13426;
  assign n13431 = ~n13429 & ~n13428;
  assign n13434 = ~n13431 & ~n13430;
  assign n13433 = ~n13432;
  assign n13437 = ~n13434 & ~n13433;
  assign n13436 = ~n13435;
  assign n13439 = ~n13437 & ~n13436;
  assign n13445 = ~n13439 & ~n13438;
  assign n13443 = ~n14909 | ~n13440;
  assign n13441 = ~n14935 | ~n8915;
  assign n13442 = ~n13441 | ~n14936;
  assign n13444 = ~n13443 | ~n13442;
  assign n13447 = ~n13445 | ~n13444;
  assign n13449 = ~n13447 | ~n13446;
  assign n13450 = ~n13449 | ~n13448;
  assign n13451 = ~n13450 & ~n9665;
  assign n13453 = n13452 | n13451;
  assign n13456 = ~n13454 | ~n13453;
  assign n13457 = ~n13456 | ~n13455;
  assign n13462 = ~n13458 | ~n13457;
  assign n13461 = ~n13460 | ~n13459;
  assign n13464 = ~n13462 | ~n13461;
  assign n13465 = ~n13464 & ~n13463;
  assign n13469 = ~n13466 & ~n13465;
  assign n13468 = ~n13467;
  assign n13471 = ~n13469 & ~n13468;
  assign n13470 = ~n14705 & ~n16424;
  assign n13473 = ~n13471 & ~n13470;
  assign n13475 = ~n13473 | ~n13472;
  assign n13476 = ~n13475 | ~n13474;
  assign n13481 = ~n13476 ^ n10531;
  assign n13478 = ~n13477 & ~P1_U3086;
  assign n13480 = ~n13479 | ~n13478;
  assign n13489 = ~n13481 & ~n13480;
  assign n13487 = ~n13483 & ~n13482;
  assign n13485 = n16026 | n13484;
  assign n13486 = ~n13485 | ~P1_B_REG_SCAN_IN;
  assign n13488 = ~n13487 & ~n13486;
  assign n13490 = ~n13489 & ~n13488;
  assign P1_U3242 = ~n13491 | ~n13490;
  assign n13494 = ~n13493 & ~n13492;
  assign n13498 = ~n13495 | ~n13494;
  assign n13497 = ~n13496 | ~n17349;
  assign n13499 = ~n13498 | ~n13497;
  assign n17511 = ~n13500 | ~n13499;
  assign n17512 = ~n17511;
  assign n13503 = ~n13501 | ~n17512;
  assign n13502 = ~n17511 | ~P2_REG1_REG_29__SCAN_IN;
  assign P2_U3488 = ~n13503 | ~n13502;
  assign n13506 = n13505 ^ n13504;
  assign n13517 = ~n13506 & ~n16610;
  assign n13515 = ~n16577 | ~n14053;
  assign n13513 = ~n12430 | ~n16616;
  assign n13509 = n16542 | n14061;
  assign n13507 = ~P2_REG3_REG_14__SCAN_IN;
  assign n16892 = ~P2_STATE_REG_SCAN_IN & ~n13507;
  assign n13508 = ~n16892;
  assign n13511 = ~n13509 | ~n13508;
  assign n13510 = ~n16574 & ~n14050;
  assign n13512 = ~n13511 & ~n13510;
  assign n13514 = n13513 & n13512;
  assign n13516 = ~n13515 | ~n13514;
  assign P2_U3155 = n13517 | n13516;
  assign n13519 = ~n13601 ^ n17525;
  assign n13529 = ~n13519 | ~n16595;
  assign n13525 = ~n13837 & ~n16542;
  assign n13523 = ~n16577 | ~n13846;
  assign n13521 = n16574 | n13886;
  assign n13520 = ~P2_REG3_REG_23__SCAN_IN | ~P2_U3151;
  assign n13522 = n13521 & n13520;
  assign n13524 = ~n13523 | ~n13522;
  assign n13527 = ~n13525 & ~n13524;
  assign n13526 = ~n14196 | ~n16616;
  assign n13528 = n13527 & n13526;
  assign P2_U3156 = ~n13529 | ~n13528;
  assign n13532 = ~n13531 | ~n13530;
  assign n13534 = ~n13533 ^ n13532;
  assign n13544 = ~n13534 | ~n16595;
  assign n13542 = ~n13931 & ~n13693;
  assign n13540 = ~n16577 | ~n13933;
  assign n13536 = ~n16605 | ~n17516;
  assign n13538 = ~n13536 | ~n13535;
  assign n13537 = ~n13974 & ~n16574;
  assign n13539 = ~n13538 & ~n13537;
  assign n13541 = ~n13540 | ~n13539;
  assign n13543 = ~n13542 & ~n13541;
  assign P2_U3159 = ~n13544 | ~n13543;
  assign n13546 = ~n13545 ^ n17519;
  assign n13548 = ~n13547 ^ n13546;
  assign n13558 = ~n13548 | ~n16595;
  assign n14213 = ~n13895;
  assign n13556 = ~n14213 & ~n13693;
  assign n13554 = ~n16577 | ~n13896;
  assign n13550 = n16574 | n13932;
  assign n13549 = ~P2_REG3_REG_21__SCAN_IN | ~P2_U3151;
  assign n13552 = ~n13550 | ~n13549;
  assign n13551 = ~n16542 & ~n13886;
  assign n13553 = ~n13552 & ~n13551;
  assign n13555 = ~n13554 | ~n13553;
  assign n13557 = ~n13556 & ~n13555;
  assign P2_U3163 = ~n13558 | ~n13557;
  assign n13561 = ~n13560 ^ n13559;
  assign n13571 = ~n13561 | ~n16595;
  assign n13569 = ~n14175 | ~n16616;
  assign n13567 = ~n13837 & ~n16574;
  assign n13565 = ~n16577 | ~n13792;
  assign n13563 = n16542 | n13801;
  assign n13562 = ~P2_REG3_REG_25__SCAN_IN | ~P2_U3151;
  assign n13564 = n13563 & n13562;
  assign n13566 = ~n13565 | ~n13564;
  assign n13568 = ~n13567 & ~n13566;
  assign n13570 = n13569 & n13568;
  assign P2_U3165 = ~n13571 | ~n13570;
  assign n13572 = ~n13587 | ~n13585;
  assign n13573 = n13572 ^ n13586;
  assign n13584 = ~n13573 & ~n16610;
  assign n13582 = ~n16577 | ~n14009;
  assign n13580 = ~n14258 | ~n16616;
  assign n13576 = n16542 | n14008;
  assign n16929 = ~P2_STATE_REG_SCAN_IN & ~n13574;
  assign n13575 = ~n16929;
  assign n13578 = ~n13576 | ~n13575;
  assign n13577 = ~n16574 & ~n14061;
  assign n13579 = ~n13578 & ~n13577;
  assign n13581 = n13580 & n13579;
  assign n13583 = ~n13582 | ~n13581;
  assign P2_U3166 = n13584 | n13583;
  assign n13588 = ~n13586 | ~n13585;
  assign n13671 = ~n13588 | ~n13587;
  assign n13590 = ~n13589 ^ n14008;
  assign n13591 = ~n13671 ^ n13590;
  assign n13600 = ~n13591 & ~n16610;
  assign n13598 = ~n16577 | ~n13984;
  assign n13596 = ~n14249 | ~n16616;
  assign n13592 = n13974 | n16542;
  assign n16947 = ~P2_REG3_REG_17__SCAN_IN | ~P2_U3151;
  assign n13594 = ~n13592 | ~n16947;
  assign n13593 = ~n16574 & ~n14032;
  assign n13595 = ~n13594 & ~n13593;
  assign n13597 = n13596 & n13595;
  assign n13599 = ~n13598 | ~n13597;
  assign P2_U3168 = n13600 | n13599;
  assign n13603 = ~n13518 & ~n13602;
  assign n13606 = ~n13605 ^ n17529;
  assign n13608 = ~n13607 ^ n13606;
  assign n13620 = ~n13608 | ~n16595;
  assign n13618 = ~n13609 & ~n13693;
  assign n13616 = n13817 | n16618;
  assign n16604 = ~n16574;
  assign n13614 = ~n17525 | ~n16604;
  assign n13612 = ~n16542 & ~n13824;
  assign n13611 = ~P2_STATE_REG_SCAN_IN & ~n13610;
  assign n13613 = ~n13612 & ~n13611;
  assign n13615 = n13614 & n13613;
  assign n13617 = ~n13616 | ~n13615;
  assign n13619 = ~n13618 & ~n13617;
  assign P2_U3169 = ~n13620 | ~n13619;
  assign n13622 = ~n13621 ^ n17516;
  assign n13624 = ~n13623 ^ n13622;
  assign n13635 = ~n13624 | ~n16595;
  assign n13633 = ~n13625 & ~n13693;
  assign n13631 = ~n16577 | ~n13910;
  assign n13629 = ~n13951 & ~n16574;
  assign n13627 = n16542 | n13909;
  assign n13626 = ~P2_REG3_REG_20__SCAN_IN | ~P2_U3151;
  assign n13628 = ~n13627 | ~n13626;
  assign n13630 = ~n13629 & ~n13628;
  assign n13632 = ~n13631 | ~n13630;
  assign n13634 = ~n13633 & ~n13632;
  assign P2_U3173 = ~n13635 | ~n13634;
  assign n13642 = ~n13637 | ~n13636;
  assign n16514 = ~n16580 | ~n13638;
  assign n16513 = n13640 & n13639;
  assign n16516 = ~n16514 | ~n16513;
  assign n13641 = ~n16516 | ~n13640;
  assign n13643 = n13642 ^ n13641;
  assign n13653 = ~n13643 & ~n16610;
  assign n13651 = ~n16577 | ~n14076;
  assign n13649 = ~n14290 | ~n16616;
  assign n13645 = n16574 | n13644;
  assign n16871 = ~P2_REG3_REG_13__SCAN_IN | ~P2_U3151;
  assign n13647 = ~n13645 | ~n16871;
  assign n13646 = ~n16542 & ~n14084;
  assign n13648 = ~n13647 & ~n13646;
  assign n13650 = n13649 & n13648;
  assign n13652 = ~n13651 | ~n13650;
  assign P2_U3174 = n13653 | n13652;
  assign n13658 = ~n13655 | ~n13654;
  assign n13657 = ~n13656 ^ n13886;
  assign n13659 = ~n13658 ^ n13657;
  assign n13669 = ~n13659 | ~n16595;
  assign n14205 = ~n13871;
  assign n13667 = ~n14205 & ~n13693;
  assign n13663 = ~n13862 & ~n16542;
  assign n13661 = ~n16604 | ~n17519;
  assign n13660 = ~P2_REG3_REG_22__SCAN_IN | ~P2_U3151;
  assign n13662 = ~n13661 | ~n13660;
  assign n13665 = ~n13663 & ~n13662;
  assign n13664 = ~n16577 | ~n13872;
  assign n13666 = ~n13665 | ~n13664;
  assign n13668 = ~n13667 & ~n13666;
  assign P2_U3175 = ~n13669 | ~n13668;
  assign n13673 = n13671 | n13670;
  assign n13675 = ~n13673 | ~n13672;
  assign n13676 = ~n13675 ^ n13674;
  assign n13687 = ~n13676 | ~n16595;
  assign n13962 = ~n13677;
  assign n13683 = ~n16577 | ~n13962;
  assign n13679 = ~n13904 | ~n16605;
  assign n13681 = ~n13679 | ~n13678;
  assign n13680 = ~n16574 & ~n14008;
  assign n13682 = ~n13681 & ~n13680;
  assign n13685 = ~n13683 | ~n13682;
  assign n14241 = ~n13961;
  assign n13684 = ~n14241 & ~n13693;
  assign n13686 = ~n13685 & ~n13684;
  assign P2_U3178 = ~n13687 | ~n13686;
  assign n13690 = ~n13689 | ~n13688;
  assign n13692 = ~n13691 ^ n13690;
  assign n13705 = ~n13692 | ~n16595;
  assign n13703 = ~n13694 & ~n13693;
  assign n13701 = ~n16577 | ~n13777;
  assign n13697 = n16574 | n13824;
  assign n13696 = P2_STATE_REG_SCAN_IN | n13695;
  assign n13699 = ~n13697 | ~n13696;
  assign n13698 = ~n16542 & ~n13776;
  assign n13700 = ~n13699 & ~n13698;
  assign n13702 = ~n13701 | ~n13700;
  assign n13704 = ~n13703 & ~n13702;
  assign P2_U3180 = ~n13705 | ~n13704;
  assign n13708 = ~n13707 ^ n13706;
  assign n13717 = ~n13708 & ~n16610;
  assign n13715 = ~n16577 | ~n14033;
  assign n13713 = ~n14269 | ~n16616;
  assign n13709 = n16542 | n14032;
  assign n16907 = ~P2_REG3_REG_15__SCAN_IN | ~P2_U3151;
  assign n13711 = ~n13709 | ~n16907;
  assign n13710 = ~n16574 & ~n14084;
  assign n13712 = ~n13711 & ~n13710;
  assign n13714 = n13713 & n13712;
  assign n13716 = ~n13715 | ~n13714;
  assign P2_U3181 = n13717 | n13716;
  assign n13724 = ~n14136 & ~n17123;
  assign n13722 = ~n17209 & ~P2_REG2_REG_31__SCAN_IN;
  assign n13721 = ~n14142 | ~n13720;
  assign n13725 = ~n17200 & ~n13721;
  assign n13723 = ~n13722 & ~n13725;
  assign P2_U3202 = n13724 | n13723;
  assign n13728 = ~n14141 | ~n17196;
  assign n13726 = ~n17209 & ~P2_REG2_REG_30__SCAN_IN;
  assign n13727 = n13726 | n13725;
  assign P2_U3203 = ~n13728 | ~n13727;
  assign n13730 = n13739 ^ n13729;
  assign n13732 = ~n13730 & ~n17356;
  assign n13731 = ~n13776 & ~n14049;
  assign n14151 = ~n13732 & ~n13731;
  assign n13734 = ~n14151 | ~n17209;
  assign n13733 = n17209 | P2_REG2_REG_28__SCAN_IN;
  assign n13750 = ~n13734 | ~n13733;
  assign n13737 = ~n13785 & ~n13735;
  assign n13738 = ~n13737 & ~n13736;
  assign n17108 = n17083 & n17088;
  assign n17128 = n17200 | n17108;
  assign n13746 = ~n14146 | ~n17196;
  assign n14085 = n17200 | n17203;
  assign n13744 = ~n14085 & ~n13740;
  assign n13742 = ~n13741;
  assign n13743 = ~n17120 & ~n13742;
  assign n13745 = ~n13744 & ~n13743;
  assign n13747 = ~n13746 | ~n13745;
  assign n13749 = ~n13748 & ~n13747;
  assign P2_U3205 = ~n13750 | ~n13749;
  assign n13754 = ~n17535 | ~n17166;
  assign n14159 = ~n13755 | ~n13754;
  assign n13757 = ~n17197 | ~n13756;
  assign n13758 = ~n17209 | ~n13757;
  assign n13759 = ~n17209 & ~P2_REG2_REG_27__SCAN_IN;
  assign n13763 = ~n13760 & ~n13759;
  assign n13762 = ~n14155 | ~n17196;
  assign n14107 = ~n14085;
  assign n13761 = ~n14107 | ~n17541;
  assign n13766 = ~n13785 | ~n13764;
  assign n13767 = ~n13766 | ~n13765;
  assign n14160 = n13768 ^ n13767;
  assign n13769 = ~n14160 | ~n14097;
  assign n13772 = ~n13770 | ~n17172;
  assign n13771 = ~n17532 | ~n17166;
  assign n14169 = ~n13772 | ~n13771;
  assign n13775 = n14169 | n17200;
  assign n13773 = ~P2_REG2_REG_26__SCAN_IN;
  assign n13774 = ~n17200 | ~n13773;
  assign n13784 = ~n13775 | ~n13774;
  assign n13782 = ~n14165 | ~n17196;
  assign n13780 = ~n14085 & ~n13776;
  assign n13778 = ~n13777;
  assign n13779 = ~n17120 & ~n13778;
  assign n13781 = ~n13780 & ~n13779;
  assign n13783 = n13782 & n13781;
  assign n13788 = n13784 & n13783;
  assign n14170 = n13786 ^ n13785;
  assign n13787 = ~n14170 | ~n14097;
  assign P2_U3207 = ~n13788 | ~n13787;
  assign n13789 = ~n9001 ^ n13806;
  assign n13791 = ~n13789 | ~n17172;
  assign n13790 = ~n17529 | ~n17166;
  assign n14179 = ~n13791 | ~n13790;
  assign n13796 = ~n14175 | ~n17185;
  assign n13793 = ~n13792;
  assign n13794 = ~n17120 & ~n13793;
  assign n13795 = ~n17200 & ~n13794;
  assign n13797 = ~n13796 | ~n13795;
  assign n13800 = n14179 | n13797;
  assign n13798 = ~P2_REG2_REG_25__SCAN_IN;
  assign n13799 = ~n17200 | ~n13798;
  assign n13803 = ~n13800 | ~n13799;
  assign n13802 = n14085 | n13801;
  assign n13809 = n13803 & n13802;
  assign n13807 = ~n13805 | ~n13804;
  assign n14180 = ~n13807 ^ n13806;
  assign n13808 = ~n14180 | ~n14097;
  assign P2_U3208 = ~n13809 | ~n13808;
  assign n13812 = n13834 | n13810;
  assign n13813 = ~n13812 | ~n13811;
  assign n13814 = ~n13813 ^ n13829;
  assign n13816 = ~n13814 | ~n17172;
  assign n13815 = ~n17525 | ~n17166;
  assign n14190 = ~n13816 | ~n13815;
  assign n13820 = ~n14186 | ~n17185;
  assign n13818 = ~n13817 & ~n17120;
  assign n13819 = ~n13818 & ~n17200;
  assign n13821 = ~n13820 | ~n13819;
  assign n13823 = ~n14190 & ~n13821;
  assign n13822 = ~n17209 & ~P2_REG2_REG_24__SCAN_IN;
  assign n13826 = ~n13823 & ~n13822;
  assign n13825 = ~n14085 & ~n13824;
  assign n13832 = ~n13826 & ~n13825;
  assign n13830 = ~n13828 | ~n13827;
  assign n14185 = ~n13830 ^ n13829;
  assign n13831 = ~n14185 | ~n14097;
  assign P2_U3209 = ~n13832 | ~n13831;
  assign n14195 = ~n13833 ^ n13835;
  assign n13843 = ~n14195 & ~n17083;
  assign n13836 = n13835 ^ n13834;
  assign n13841 = ~n13836 | ~n17172;
  assign n13839 = ~n13837 & ~n17203;
  assign n13838 = ~n13886 & ~n14049;
  assign n13840 = ~n13839 & ~n13838;
  assign n13842 = ~n13841 | ~n13840;
  assign n14201 = ~n13843 & ~n13842;
  assign n13845 = ~n14201 | ~n17209;
  assign n13844 = n17209 | P2_REG2_REG_23__SCAN_IN;
  assign n13852 = ~n13845 | ~n13844;
  assign n13850 = ~n14195 & ~n13983;
  assign n13848 = ~n14196 | ~n17196;
  assign n13847 = ~n13846 | ~n17197;
  assign n13849 = ~n13848 | ~n13847;
  assign n13851 = ~n13850 & ~n13849;
  assign P2_U3210 = ~n13852 | ~n13851;
  assign n14204 = ~n13854 ^ n13853;
  assign n13868 = ~n14204 & ~n17083;
  assign n13858 = ~n13855 | ~n13856;
  assign n13860 = ~n13858 | ~n13857;
  assign n13861 = ~n13860 ^ n13859;
  assign n13866 = ~n13861 | ~n17172;
  assign n13864 = ~n13862 & ~n17203;
  assign n13863 = ~n13909 & ~n14049;
  assign n13865 = ~n13864 & ~n13863;
  assign n13867 = ~n13866 | ~n13865;
  assign n14209 = ~n13868 & ~n13867;
  assign n13870 = ~n14209 | ~n17209;
  assign n13869 = n17209 | P2_REG2_REG_22__SCAN_IN;
  assign n13878 = ~n13870 | ~n13869;
  assign n13876 = ~n14204 & ~n13983;
  assign n13874 = ~n13871 | ~n17196;
  assign n13873 = ~n17197 | ~n13872;
  assign n13875 = ~n13874 | ~n13873;
  assign n13877 = ~n13876 & ~n13875;
  assign P2_U3211 = ~n13878 | ~n13877;
  assign n14212 = ~n13880 ^ n13879;
  assign n13892 = ~n14212 & ~n17083;
  assign n13882 = ~n13855 | ~n13918;
  assign n13884 = ~n13882 | ~n13881;
  assign n13885 = ~n13884 ^ n13883;
  assign n13890 = ~n13885 | ~n17172;
  assign n13888 = ~n13886 & ~n17203;
  assign n13887 = ~n13932 & ~n14049;
  assign n13889 = ~n13888 & ~n13887;
  assign n13891 = ~n13890 | ~n13889;
  assign n14217 = ~n13892 & ~n13891;
  assign n13894 = ~n14217 | ~n17209;
  assign n13893 = n17209 | P2_REG2_REG_21__SCAN_IN;
  assign n13902 = ~n13894 | ~n13893;
  assign n13900 = ~n14212 & ~n13983;
  assign n13898 = ~n13895 | ~n17196;
  assign n13897 = ~n17197 | ~n13896;
  assign n13899 = ~n13898 | ~n13897;
  assign n13901 = ~n13900 & ~n13899;
  assign P2_U3212 = ~n13902 | ~n13901;
  assign n13903 = ~n13855 ^ n13918;
  assign n13906 = ~n13903 | ~n17172;
  assign n13905 = ~n13904 | ~n17166;
  assign n14225 = ~n13906 | ~n13905;
  assign n13908 = ~n14225 & ~n17200;
  assign n13907 = ~n17209 & ~P2_REG2_REG_20__SCAN_IN;
  assign n13917 = ~n13908 & ~n13907;
  assign n13915 = ~n14221 | ~n17196;
  assign n13913 = ~n14085 & ~n13909;
  assign n13911 = ~n13910;
  assign n13912 = ~n17120 & ~n13911;
  assign n13914 = ~n13913 & ~n13912;
  assign n13916 = ~n13915 | ~n13914;
  assign n13921 = ~n13917 & ~n13916;
  assign n14220 = ~n13919 ^ n13918;
  assign n13920 = ~n14220 | ~n14097;
  assign P2_U3213 = ~n13921 | ~n13920;
  assign n13940 = ~n13923 | ~n13922;
  assign n13925 = ~n13924 ^ n13940;
  assign n13928 = ~n13925 | ~n17172;
  assign n13927 = ~n13926 | ~n17166;
  assign n14235 = ~n13928 | ~n13927;
  assign n13930 = ~n14235 & ~n17200;
  assign n13929 = ~n17209 & ~P2_REG2_REG_19__SCAN_IN;
  assign n13939 = ~n13930 & ~n13929;
  assign n13937 = ~n13931 & ~n17123;
  assign n13935 = n14085 | n13932;
  assign n13934 = ~n13933 | ~n17197;
  assign n13936 = ~n13935 | ~n13934;
  assign n13938 = n13937 | n13936;
  assign n13943 = ~n13939 & ~n13938;
  assign n14230 = ~n13941 ^ n13940;
  assign n13942 = ~n14230 | ~n14097;
  assign P2_U3214 = ~n13943 | ~n13942;
  assign n13946 = ~n13944;
  assign n13949 = ~n13946 & ~n13945;
  assign n14240 = ~n13947 ^ n13949;
  assign n13957 = ~n14240 & ~n17083;
  assign n13950 = n13949 ^ n13948;
  assign n13955 = ~n13950 | ~n17172;
  assign n13953 = ~n13951 & ~n17203;
  assign n13952 = ~n14008 & ~n14049;
  assign n13954 = ~n13953 & ~n13952;
  assign n13956 = ~n13955 | ~n13954;
  assign n14245 = ~n13957 & ~n13956;
  assign n13960 = ~n14245 | ~n17209;
  assign n13959 = ~n17200 | ~n13958;
  assign n13968 = ~n13960 | ~n13959;
  assign n13966 = ~n14240 & ~n13983;
  assign n13964 = ~n13961 | ~n17196;
  assign n13963 = ~n13962 | ~n17197;
  assign n13965 = ~n13964 | ~n13963;
  assign n13967 = ~n13966 & ~n13965;
  assign P2_U3215 = ~n13968 | ~n13967;
  assign n14248 = ~n13970 ^ n13969;
  assign n13980 = ~n14248 & ~n17083;
  assign n13973 = ~n13972 ^ n13971;
  assign n13978 = ~n13973 | ~n17172;
  assign n13976 = ~n13974 & ~n17203;
  assign n13975 = ~n14032 & ~n14049;
  assign n13977 = ~n13976 & ~n13975;
  assign n13979 = ~n13978 | ~n13977;
  assign n14254 = ~n13980 & ~n13979;
  assign n13982 = ~n14254 | ~n17209;
  assign n13981 = ~n17200 | ~n11265;
  assign n13990 = ~n13982 | ~n13981;
  assign n13988 = ~n14248 & ~n13983;
  assign n13986 = ~n14249 | ~n17196;
  assign n13985 = ~n13984 | ~n17197;
  assign n13987 = ~n13986 | ~n13985;
  assign n13989 = ~n13988 & ~n13987;
  assign P2_U3216 = ~n13990 | ~n13989;
  assign n13993 = ~n14043 | ~n13991;
  assign n13994 = n13993 & n13992;
  assign n14257 = n13998 ^ n13994;
  assign n14015 = ~n14257 | ~n14097;
  assign n13997 = n14072 | n13995;
  assign n13999 = ~n13997 | ~n13996;
  assign n14000 = ~n13999 & ~n13998;
  assign n14001 = ~n14000 & ~n17356;
  assign n14003 = ~n14001 | ~n8922;
  assign n14002 = n14061 | n14049;
  assign n14263 = ~n14003 | ~n14002;
  assign n14004 = ~n14258 | ~n17185;
  assign n14005 = ~n14004 | ~n17209;
  assign n14007 = n14263 | n14005;
  assign n14006 = ~n17200 | ~n11259;
  assign n14013 = ~n14007 | ~n14006;
  assign n14011 = n14085 | n14008;
  assign n14010 = ~n17197 | ~n14009;
  assign n14012 = n14011 & n14010;
  assign n14014 = n14013 & n14012;
  assign P2_U3217 = ~n14015 | ~n14014;
  assign n14018 = ~n14043 | ~n14016;
  assign n14019 = n14018 & n14017;
  assign n14268 = n14024 ^ n14019;
  assign n14041 = ~n14268 | ~n14097;
  assign n14046 = n14072 | n14020;
  assign n14023 = ~n14046 | ~n14021;
  assign n14025 = n14023 & n14022;
  assign n14026 = n14025 ^ n14024;
  assign n14028 = ~n14026 | ~n17172;
  assign n14027 = ~n14291 | ~n17166;
  assign n14274 = ~n14028 | ~n14027;
  assign n14030 = ~n14274 & ~n17200;
  assign n14029 = ~n17209 & ~P2_REG2_REG_15__SCAN_IN;
  assign n14039 = ~n14030 & ~n14029;
  assign n14031 = ~n14269;
  assign n14037 = ~n14031 & ~n17123;
  assign n14035 = n14085 | n14032;
  assign n14034 = ~n17197 | ~n14033;
  assign n14036 = ~n14035 | ~n14034;
  assign n14038 = n14037 | n14036;
  assign n14040 = ~n14039 & ~n14038;
  assign P2_U3218 = ~n14041 | ~n14040;
  assign n14044 = ~n14043 | ~n14042;
  assign n14279 = ~n14044 ^ n12969;
  assign n14065 = ~n14279 | ~n14097;
  assign n14047 = ~n14046 | ~n14045;
  assign n14048 = ~n14047 ^ n12969;
  assign n14052 = ~n14048 | ~n17172;
  assign n14051 = n14050 | n14049;
  assign n14284 = ~n14052 | ~n14051;
  assign n14057 = ~n12430 | ~n17185;
  assign n14054 = ~n14053;
  assign n14055 = ~n17120 & ~n14054;
  assign n14056 = ~n17200 & ~n14055;
  assign n14058 = ~n14057 | ~n14056;
  assign n14060 = n14284 | n14058;
  assign n14059 = ~n17200 | ~n11243;
  assign n14063 = ~n14060 | ~n14059;
  assign n14062 = n14085 | n14061;
  assign n14064 = n14063 & n14062;
  assign P2_U3219 = ~n14065 | ~n14064;
  assign n14069 = n14067 & n14066;
  assign n14070 = ~n14069 | ~n14068;
  assign n14289 = n14071 ^ n14070;
  assign n14089 = ~n14289 | ~n14097;
  assign n14073 = n14072 ^ n14071;
  assign n14075 = ~n14073 | ~n17172;
  assign n14074 = ~n16974 | ~n17166;
  assign n14295 = ~n14075 | ~n14074;
  assign n14080 = ~n14290 | ~n17185;
  assign n14077 = ~n14076;
  assign n14078 = ~n17120 & ~n14077;
  assign n14079 = ~n17200 & ~n14078;
  assign n14081 = ~n14080 | ~n14079;
  assign n14083 = ~n14295 & ~n14081;
  assign n14082 = ~n17209 & ~P2_REG2_REG_13__SCAN_IN;
  assign n14087 = ~n14083 & ~n14082;
  assign n14086 = ~n14085 & ~n14084;
  assign n14088 = ~n14087 & ~n14086;
  assign P2_U3220 = ~n14089 | ~n14088;
  assign n14092 = ~n17015 | ~n14090;
  assign n14095 = ~n16993 | ~n14093;
  assign n14096 = n14095 & n14094;
  assign n17461 = n14098 ^ n14096;
  assign n14113 = ~n17461 | ~n14097;
  assign n14100 = ~n14099 ^ n14098;
  assign n14102 = ~n14100 | ~n17172;
  assign n14101 = ~n14116 | ~n17166;
  assign n17469 = ~n14102 | ~n14101;
  assign n14103 = ~n17197 | ~n16510;
  assign n14104 = ~n17209 | ~n14103;
  assign n14106 = ~n17469 & ~n14104;
  assign n14105 = ~n17209 & ~P2_REG2_REG_12__SCAN_IN;
  assign n14111 = ~n14106 & ~n14105;
  assign n14109 = ~n17463 | ~n17196;
  assign n14108 = ~n14107 | ~n17465;
  assign n14110 = ~n14109 | ~n14108;
  assign n14112 = ~n14111 & ~n14110;
  assign P2_U3221 = ~n14113 | ~n14112;
  assign n14115 = ~n17200 | ~P2_REG2_REG_10__SCAN_IN;
  assign n14114 = ~n17197 | ~n16449;
  assign n14133 = ~n14115 | ~n14114;
  assign n14118 = ~n14116 | ~n17464;
  assign n14117 = ~n17009 | ~n17166;
  assign n14123 = ~n14118 | ~n14117;
  assign n14120 = ~n16993 | ~n16992;
  assign n14121 = ~n14120 | ~n14119;
  assign n17441 = n14126 ^ n14121;
  assign n14122 = ~n17441 & ~n17083;
  assign n14129 = ~n14123 & ~n14122;
  assign n16968 = ~n14125 | ~n14124;
  assign n14127 = ~n16968 ^ n14126;
  assign n14128 = ~n14127 | ~n17172;
  assign n17439 = ~n14129 | ~n14128;
  assign n14130 = ~n17441 & ~n17088;
  assign n14131 = ~n17439 & ~n14130;
  assign n14132 = ~n17200 & ~n14131;
  assign n14135 = ~n14133 & ~n14132;
  assign n14134 = ~n17196 | ~n16442;
  assign P2_U3223 = ~n14135 | ~n14134;
  assign n14137 = ~n14136;
  assign n17462 = ~n17452;
  assign n14138 = ~n14137 | ~n17462;
  assign n14300 = ~n14138 | ~n14142;
  assign n14140 = ~n14300 | ~n17512;
  assign n14139 = ~n17511 | ~P2_REG1_REG_31__SCAN_IN;
  assign P2_U3490 = ~n14140 | ~n14139;
  assign n14143 = ~n14141 | ~n17462;
  assign n14303 = ~n14143 | ~n14142;
  assign n14145 = ~n14303 | ~n17512;
  assign n14144 = ~n17511 | ~P2_REG1_REG_30__SCAN_IN;
  assign P2_U3489 = ~n14145 | ~n14144;
  assign n14148 = ~n14146 | ~n17462;
  assign n14147 = ~n17544 | ~n17464;
  assign n14149 = ~n14148 | ~n14147;
  assign n14152 = ~n14150 & ~n14149;
  assign n14306 = ~n14152 | ~n14151;
  assign n14154 = ~n14306 | ~n17512;
  assign n14153 = ~n17511 | ~P2_REG1_REG_28__SCAN_IN;
  assign P2_U3487 = ~n14154 | ~n14153;
  assign n14157 = ~n14155 | ~n17462;
  assign n14156 = ~n17541 | ~n17464;
  assign n14158 = ~n14157 | ~n14156;
  assign n14162 = ~n14159 & ~n14158;
  assign n14161 = ~n14160 | ~n9107;
  assign n14309 = ~n14162 | ~n14161;
  assign n14164 = ~n14309 | ~n17512;
  assign n14163 = ~n17511 | ~P2_REG1_REG_27__SCAN_IN;
  assign P2_U3486 = ~n14164 | ~n14163;
  assign n14167 = ~n14165 | ~n17462;
  assign n14166 = ~n17538 | ~n17464;
  assign n14168 = ~n14167 | ~n14166;
  assign n14172 = ~n14169 & ~n14168;
  assign n14171 = ~n14170 | ~n9107;
  assign n14312 = ~n14172 | ~n14171;
  assign n14174 = ~n14312 | ~n17512;
  assign n14173 = ~n17511 | ~P2_REG1_REG_26__SCAN_IN;
  assign P2_U3485 = ~n14174 | ~n14173;
  assign n14177 = ~n14175 | ~n17462;
  assign n14176 = ~n17535 | ~n17464;
  assign n14178 = ~n14177 | ~n14176;
  assign n14182 = ~n14179 & ~n14178;
  assign n14181 = ~n14180 | ~n9107;
  assign n14315 = ~n14182 | ~n14181;
  assign n14184 = ~n14315 | ~n17512;
  assign n14183 = ~n17511 | ~P2_REG1_REG_25__SCAN_IN;
  assign P2_U3484 = ~n14184 | ~n14183;
  assign n14192 = ~n14185 | ~n9107;
  assign n14188 = ~n14186 | ~n17462;
  assign n14187 = ~n17532 | ~n17464;
  assign n14189 = ~n14188 | ~n14187;
  assign n14191 = ~n14190 & ~n14189;
  assign n14318 = ~n14192 | ~n14191;
  assign n14194 = ~n14318 | ~n17512;
  assign n14193 = ~n17511 | ~P2_REG1_REG_24__SCAN_IN;
  assign P2_U3483 = ~n14194 | ~n14193;
  assign n14199 = ~n14195 & ~n17440;
  assign n14197 = ~n14196;
  assign n14198 = ~n14197 & ~n17452;
  assign n14200 = ~n14199 & ~n14198;
  assign n14321 = ~n14201 | ~n14200;
  assign n14203 = ~n14321 | ~n17512;
  assign n14202 = ~n17511 | ~P2_REG1_REG_23__SCAN_IN;
  assign P2_U3482 = ~n14203 | ~n14202;
  assign n14207 = ~n14204 & ~n17440;
  assign n14206 = ~n14205 & ~n17452;
  assign n14208 = ~n14207 & ~n14206;
  assign n14324 = ~n14209 | ~n14208;
  assign n14211 = ~n14324 | ~n17512;
  assign n14210 = ~n17511 | ~P2_REG1_REG_22__SCAN_IN;
  assign P2_U3481 = ~n14211 | ~n14210;
  assign n14215 = ~n14212 & ~n17440;
  assign n14214 = ~n14213 & ~n17452;
  assign n14216 = ~n14215 & ~n14214;
  assign n14327 = ~n14217 | ~n14216;
  assign n14219 = ~n14327 | ~n17512;
  assign n14218 = ~n17511 | ~P2_REG1_REG_21__SCAN_IN;
  assign P2_U3480 = ~n14219 | ~n14218;
  assign n14227 = ~n14220 | ~n9107;
  assign n14223 = ~n14221 | ~n17462;
  assign n14222 = ~n17519 | ~n17464;
  assign n14224 = ~n14223 | ~n14222;
  assign n14226 = ~n14225 & ~n14224;
  assign n14330 = ~n14227 | ~n14226;
  assign n14229 = ~n14330 | ~n17512;
  assign n14228 = ~n17511 | ~P2_REG1_REG_20__SCAN_IN;
  assign P2_U3479 = ~n14229 | ~n14228;
  assign n14237 = ~n14230 | ~n9107;
  assign n14233 = ~n14231 | ~n17462;
  assign n14232 = ~n17516 | ~n17464;
  assign n14234 = ~n14233 | ~n14232;
  assign n14236 = ~n14235 & ~n14234;
  assign n14333 = ~n14237 | ~n14236;
  assign n14239 = ~n14333 | ~n17512;
  assign n14238 = ~n17511 | ~P2_REG1_REG_19__SCAN_IN;
  assign P2_U3478 = ~n14239 | ~n14238;
  assign n14243 = ~n14240 & ~n17440;
  assign n14242 = ~n14241 & ~n17452;
  assign n14244 = ~n14243 & ~n14242;
  assign n14336 = ~n14245 | ~n14244;
  assign n14247 = ~n14336 | ~n17512;
  assign n14246 = ~n17511 | ~P2_REG1_REG_18__SCAN_IN;
  assign P2_U3477 = ~n14247 | ~n14246;
  assign n14252 = ~n14248 & ~n17440;
  assign n14250 = ~n14249;
  assign n14251 = ~n14250 & ~n17452;
  assign n14253 = ~n14252 & ~n14251;
  assign n14339 = ~n14254 | ~n14253;
  assign n14256 = ~n14339 | ~n17512;
  assign n14255 = ~n17511 | ~P2_REG1_REG_17__SCAN_IN;
  assign P2_U3476 = ~n14256 | ~n14255;
  assign n14265 = ~n14257 | ~n9107;
  assign n14261 = ~n14258 | ~n17462;
  assign n14260 = ~n14259 | ~n17464;
  assign n14262 = ~n14261 | ~n14260;
  assign n14264 = ~n14263 & ~n14262;
  assign n14342 = ~n14265 | ~n14264;
  assign n14267 = ~n14342 | ~n17512;
  assign n14266 = ~n17511 | ~P2_REG1_REG_16__SCAN_IN;
  assign P2_U3475 = ~n14267 | ~n14266;
  assign n14276 = ~n14268 | ~n9107;
  assign n14272 = ~n14269 | ~n17462;
  assign n14271 = ~n14270 | ~n17464;
  assign n14273 = ~n14272 | ~n14271;
  assign n14275 = ~n14274 & ~n14273;
  assign n14345 = ~n14276 | ~n14275;
  assign n14278 = ~n14345 | ~n17512;
  assign n14277 = ~n17511 | ~P2_REG1_REG_15__SCAN_IN;
  assign P2_U3474 = ~n14278 | ~n14277;
  assign n14286 = ~n14279 | ~n9107;
  assign n14282 = ~n12430 | ~n17462;
  assign n14281 = ~n14280 | ~n17464;
  assign n14283 = ~n14282 | ~n14281;
  assign n14285 = ~n14284 & ~n14283;
  assign n14348 = ~n14286 | ~n14285;
  assign n14288 = ~n14348 | ~n17512;
  assign n14287 = ~n17511 | ~P2_REG1_REG_14__SCAN_IN;
  assign P2_U3473 = ~n14288 | ~n14287;
  assign n14297 = ~n14289 | ~n9107;
  assign n14293 = ~n14290 | ~n17462;
  assign n14292 = ~n14291 | ~n17464;
  assign n14294 = ~n14293 | ~n14292;
  assign n14296 = ~n14295 & ~n14294;
  assign n14351 = ~n14297 | ~n14296;
  assign n14299 = ~n14351 | ~n17512;
  assign n14298 = ~n17511 | ~P2_REG1_REG_13__SCAN_IN;
  assign P2_U3472 = ~n14299 | ~n14298;
  assign n14302 = ~n14300 | ~n17472;
  assign n14301 = ~n17460 | ~P2_REG0_REG_31__SCAN_IN;
  assign P2_U3458 = ~n14302 | ~n14301;
  assign n14305 = ~n14303 | ~n17472;
  assign n14304 = ~n17460 | ~P2_REG0_REG_30__SCAN_IN;
  assign P2_U3457 = ~n14305 | ~n14304;
  assign n14308 = ~n14306 | ~n17472;
  assign n14307 = ~n17460 | ~P2_REG0_REG_28__SCAN_IN;
  assign P2_U3455 = ~n14308 | ~n14307;
  assign n14311 = ~n14309 | ~n17472;
  assign n14310 = ~n17460 | ~P2_REG0_REG_27__SCAN_IN;
  assign P2_U3454 = ~n14311 | ~n14310;
  assign n14314 = ~n14312 | ~n17472;
  assign n14313 = ~n17460 | ~P2_REG0_REG_26__SCAN_IN;
  assign P2_U3453 = ~n14314 | ~n14313;
  assign n14317 = ~n14315 | ~n17472;
  assign n14316 = ~n17460 | ~P2_REG0_REG_25__SCAN_IN;
  assign P2_U3452 = ~n14317 | ~n14316;
  assign n14320 = ~n14318 | ~n17472;
  assign n14319 = ~n17460 | ~P2_REG0_REG_24__SCAN_IN;
  assign P2_U3451 = ~n14320 | ~n14319;
  assign n14323 = ~n14321 | ~n17472;
  assign n14322 = ~n17460 | ~P2_REG0_REG_23__SCAN_IN;
  assign P2_U3450 = ~n14323 | ~n14322;
  assign n14326 = ~n14324 | ~n17472;
  assign n14325 = ~n17460 | ~P2_REG0_REG_22__SCAN_IN;
  assign P2_U3449 = ~n14326 | ~n14325;
  assign n14329 = ~n14327 | ~n17472;
  assign n14328 = ~n17460 | ~P2_REG0_REG_21__SCAN_IN;
  assign P2_U3448 = ~n14329 | ~n14328;
  assign n14332 = ~n14330 | ~n17472;
  assign n14331 = ~n17460 | ~P2_REG0_REG_20__SCAN_IN;
  assign P2_U3447 = ~n14332 | ~n14331;
  assign n14335 = ~n14333 | ~n17472;
  assign n14334 = ~n17460 | ~P2_REG0_REG_19__SCAN_IN;
  assign P2_U3446 = ~n14335 | ~n14334;
  assign n14338 = ~n14336 | ~n17472;
  assign n14337 = ~n17460 | ~P2_REG0_REG_18__SCAN_IN;
  assign P2_U3444 = ~n14338 | ~n14337;
  assign n14341 = ~n14339 | ~n17472;
  assign n14340 = ~n17460 | ~P2_REG0_REG_17__SCAN_IN;
  assign P2_U3441 = ~n14341 | ~n14340;
  assign n14344 = ~n14342 | ~n17472;
  assign n14343 = ~n17460 | ~P2_REG0_REG_16__SCAN_IN;
  assign P2_U3438 = ~n14344 | ~n14343;
  assign n14347 = ~n14345 | ~n17472;
  assign n14346 = ~n17460 | ~P2_REG0_REG_15__SCAN_IN;
  assign P2_U3435 = ~n14347 | ~n14346;
  assign n14350 = ~n14348 | ~n17472;
  assign n14349 = ~n17460 | ~P2_REG0_REG_14__SCAN_IN;
  assign P2_U3432 = ~n14350 | ~n14349;
  assign n14353 = ~n14351 | ~n17472;
  assign n14352 = ~n17460 | ~P2_REG0_REG_13__SCAN_IN;
  assign P2_U3429 = ~n14353 | ~n14352;
  assign n14361 = ~n15232 & ~n17341;
  assign n14357 = ~n14354;
  assign n14355 = ~P2_IR_REG_31__SCAN_IN | ~P2_STATE_REG_SCAN_IN;
  assign n14356 = ~n14355 & ~P2_IR_REG_30__SCAN_IN;
  assign n14359 = ~n14357 | ~n14356;
  assign n14358 = ~n17338 | ~P1_DATAO_REG_31__SCAN_IN;
  assign n14360 = ~n14359 | ~n14358;
  assign P2_U3264 = n14361 | n14360;
  assign n14366 = ~n15241 & ~n17341;
  assign n14364 = ~n14362 | ~P2_STATE_REG_SCAN_IN;
  assign n14363 = ~n17338 | ~P1_DATAO_REG_30__SCAN_IN;
  assign n14365 = ~n14364 | ~n14363;
  assign P2_U3265 = n14366 | n14365;
  assign n14369 = ~n14368 | ~n14367;
  assign n14371 = n14370 ^ n14369;
  assign n14381 = ~n14371 & ~n15293;
  assign n14379 = ~n15311 | ~n14372;
  assign n14377 = ~n9555 | ~n15361;
  assign n14373 = n15332 | n14455;
  assign n15533 = ~P1_REG3_REG_14__SCAN_IN | ~P1_U3086;
  assign n14375 = ~n14373 | ~n15533;
  assign n14374 = ~n15319 & ~n14997;
  assign n14376 = ~n14375 & ~n14374;
  assign n14378 = n14377 & n14376;
  assign n14380 = ~n14379 | ~n14378;
  assign P1_U3215 = n14381 | n14380;
  assign n14383 = ~n14520 ^ n14518;
  assign n14384 = ~n14382 ^ n14383;
  assign n14394 = ~n14384 | ~n15376;
  assign n14392 = ~n14822 & ~n15333;
  assign n14390 = ~n15311 | ~n14824;
  assign n14386 = n15332 | n14865;
  assign n14385 = ~P1_REG3_REG_23__SCAN_IN | ~P1_U3086;
  assign n14388 = ~n14386 | ~n14385;
  assign n14387 = ~n15319 & ~n14817;
  assign n14389 = ~n14388 & ~n14387;
  assign n14391 = ~n14390 | ~n14389;
  assign n14393 = ~n14392 & ~n14391;
  assign P1_U3216 = ~n14394 | ~n14393;
  assign n14586 = ~n14395 ^ n14587;
  assign n14396 = ~n14586 ^ n14585;
  assign n14403 = ~n14396 | ~n15376;
  assign n14398 = ~n15358 | ~n15711;
  assign n14401 = ~n14398 | ~n14397;
  assign n14400 = ~n15332 & ~n14399;
  assign n14402 = ~n14401 & ~n14400;
  assign n14405 = ~n14403 | ~n14402;
  assign n14404 = ~n15381 & ~n15705;
  assign n14407 = ~n14405 & ~n14404;
  assign n14406 = ~n16279 | ~n15361;
  assign P1_U3217 = ~n14407 | ~n14406;
  assign n14608 = ~n14409 ^ n14408;
  assign n14411 = ~n14608 & ~n14607;
  assign n14410 = ~n14409 & ~n14408;
  assign n14417 = ~n14411 & ~n14410;
  assign n14414 = ~n14413 | ~n14412;
  assign n14416 = ~n14415 | ~n14414;
  assign n14418 = ~n14417 ^ n14416;
  assign n14427 = ~n14418 | ~n15376;
  assign n14425 = ~n14924 & ~n15333;
  assign n14423 = ~n15311 | ~n14925;
  assign n14419 = ~n15319 & ~n14866;
  assign n14649 = P1_U3086 & P1_REG3_REG_19__SCAN_IN;
  assign n14421 = n14419 | n14649;
  assign n14420 = ~n15332 & ~n14972;
  assign n14422 = ~n14421 & ~n14420;
  assign n14424 = ~n14423 | ~n14422;
  assign n14426 = ~n14425 & ~n14424;
  assign P1_U3219 = ~n14427 | ~n14426;
  assign n14429 = ~n14430;
  assign n14538 = ~n14429 & ~n14428;
  assign n14541 = ~n14539 | ~n14538;
  assign n14434 = ~n14541 | ~n14430;
  assign n14433 = ~n14432 ^ n14431;
  assign n14435 = ~n14434 ^ n14433;
  assign n14445 = ~n14435 | ~n15376;
  assign n14443 = ~n14876 & ~n15333;
  assign n14441 = ~n15311 | ~n14877;
  assign n14437 = n15332 | n14866;
  assign n14436 = ~P1_REG3_REG_21__SCAN_IN | ~P1_U3086;
  assign n14439 = ~n14437 | ~n14436;
  assign n14438 = ~n15319 & ~n14865;
  assign n14440 = ~n14439 & ~n14438;
  assign n14442 = ~n14441 | ~n14440;
  assign n14444 = ~n14443 & ~n14442;
  assign P1_U3223 = ~n14445 | ~n14444;
  assign n14452 = ~n14447 | ~n14446;
  assign n14450 = ~n14448;
  assign n14451 = ~n14450 & ~n14449;
  assign n14453 = ~n14452 ^ n14451;
  assign n14465 = ~n14453 & ~n15293;
  assign n14463 = ~n15311 | ~n14454;
  assign n14461 = n15659 | n15333;
  assign n14456 = n15319 | n14455;
  assign n15508 = ~P1_REG3_REG_12__SCAN_IN | ~P1_U3086;
  assign n14459 = ~n14456 | ~n15508;
  assign n14458 = ~n15332 & ~n14457;
  assign n14460 = ~n14459 & ~n14458;
  assign n14462 = n14461 & n14460;
  assign n14464 = ~n14463 | ~n14462;
  assign P1_U3224 = n14465 | n14464;
  assign n14469 = n14467 | n14466;
  assign n14470 = ~n14469 | ~n14468;
  assign n14480 = ~n14470 | ~n15376;
  assign n14478 = ~n14778 & ~n15333;
  assign n14476 = ~n15311 | ~n14781;
  assign n14472 = n15332 | n14817;
  assign n14471 = ~P1_REG3_REG_25__SCAN_IN | ~P1_U3086;
  assign n14474 = ~n14472 | ~n14471;
  assign n14473 = ~n15319 & ~n14773;
  assign n14475 = ~n14474 & ~n14473;
  assign n14477 = ~n14476 | ~n14475;
  assign n14479 = ~n14478 & ~n14477;
  assign P1_U3225 = ~n14480 | ~n14479;
  assign n14482 = ~n14484;
  assign n14635 = ~n14482 & ~n14481;
  assign n14485 = ~n14635 & ~n14636;
  assign n14634 = ~n14484 & ~n14483;
  assign n14488 = ~n14485 & ~n14634;
  assign n14487 = n14486 & n14501;
  assign n14502 = ~n14488 | ~n14487;
  assign n14490 = ~n14502;
  assign n14489 = ~n14488 & ~n14487;
  assign n14491 = ~n14490 & ~n14489;
  assign n14500 = ~n14491 & ~n15293;
  assign n14498 = ~n15311 | ~n14987;
  assign n14496 = ~n15167 | ~n15361;
  assign n14492 = n15332 | n14997;
  assign n15562 = ~P1_REG3_REG_16__SCAN_IN | ~P1_U3086;
  assign n14494 = ~n14492 | ~n15562;
  assign n14493 = ~n15319 & ~n14998;
  assign n14495 = ~n14494 & ~n14493;
  assign n14497 = n14496 & n14495;
  assign n14499 = ~n14498 | ~n14497;
  assign P1_U3226 = n14500 | n14499;
  assign n14506 = ~n14502 | ~n14501;
  assign n14505 = ~n14504 | ~n14503;
  assign n14507 = ~n14506 ^ n14505;
  assign n14516 = ~n14507 & ~n15293;
  assign n14512 = ~n15157 | ~n15361;
  assign n14508 = n15319 | n14972;
  assign n15577 = ~P1_REG3_REG_17__SCAN_IN | ~P1_U3086;
  assign n14510 = ~n14508 | ~n15577;
  assign n14509 = ~n15332 & ~n15011;
  assign n14511 = ~n14510 & ~n14509;
  assign n14514 = n14512 & n14511;
  assign n14513 = ~n15311 | ~n14962;
  assign n14515 = ~n14514 | ~n14513;
  assign P1_U3228 = n14516 | n14515;
  assign n14519 = ~n10738 | ~n14517;
  assign n14522 = ~n14519 | ~n14518;
  assign n14521 = ~n14382 | ~n14520;
  assign n14526 = ~n14522 | ~n14521;
  assign n14525 = ~n14524 | ~n14523;
  assign n14527 = ~n14526 ^ n14525;
  assign n14537 = ~n14527 | ~n15376;
  assign n14535 = ~n14802 & ~n15333;
  assign n14533 = ~n15311 | ~n14803;
  assign n14529 = n15332 | n14839;
  assign n14528 = ~P1_REG3_REG_24__SCAN_IN | ~P1_U3086;
  assign n14531 = ~n14529 | ~n14528;
  assign n14530 = ~n15319 & ~n14622;
  assign n14532 = ~n14531 & ~n14530;
  assign n14534 = ~n14533 | ~n14532;
  assign n14536 = ~n14535 & ~n14534;
  assign P1_U3229 = ~n14537 | ~n14536;
  assign n14540 = n14539 | n14538;
  assign n14542 = ~n14541 | ~n14540;
  assign n14552 = ~n14542 | ~n15376;
  assign n14550 = ~n9573 & ~n15333;
  assign n14548 = ~n15311 | ~n14898;
  assign n14544 = ~n15360 | ~n16391;
  assign n14543 = ~P1_REG3_REG_20__SCAN_IN | ~P1_U3086;
  assign n14546 = ~n14544 | ~n14543;
  assign n14545 = ~n15319 & ~n14891;
  assign n14547 = ~n14546 & ~n14545;
  assign n14549 = ~n14548 | ~n14547;
  assign n14551 = ~n14550 & ~n14549;
  assign P1_U3233 = ~n14552 | ~n14551;
  assign n14555 = ~n14554 | ~n14553;
  assign n14557 = ~n14556 ^ n14555;
  assign n14569 = ~n14557 & ~n15293;
  assign n14567 = ~n15311 | ~n14558;
  assign n14565 = ~n16315 | ~n15361;
  assign n14561 = n15332 | n14559;
  assign n15519 = P1_U3086 & P1_REG3_REG_13__SCAN_IN;
  assign n14560 = ~n15519;
  assign n14563 = ~n14561 | ~n14560;
  assign n14562 = ~n15319 & ~n15012;
  assign n14564 = ~n14563 & ~n14562;
  assign n14566 = n14565 & n14564;
  assign n14568 = ~n14567 | ~n14566;
  assign P1_U3234 = n14569 | n14568;
  assign n14573 = ~n14571 | ~n14570;
  assign n14574 = ~n14573 ^ n14572;
  assign n14584 = ~n14574 | ~n15376;
  assign n14582 = ~n9570 & ~n15333;
  assign n14580 = ~n15311 | ~n14851;
  assign n14576 = n15332 | n14891;
  assign n14575 = ~P1_REG3_REG_22__SCAN_IN | ~P1_U3086;
  assign n14578 = ~n14576 | ~n14575;
  assign n14577 = ~n15319 & ~n14839;
  assign n14579 = ~n14578 & ~n14577;
  assign n14581 = ~n14580 | ~n14579;
  assign n14583 = ~n14582 & ~n14581;
  assign P1_U3235 = ~n14584 | ~n14583;
  assign n14589 = ~n14586 & ~n14585;
  assign n14588 = ~n14395 & ~n14587;
  assign n14594 = n14589 | n14588;
  assign n14593 = ~n14591 | ~n14590;
  assign n14592 = ~n14594 & ~n14593;
  assign n14596 = ~n14592 & ~n15293;
  assign n14595 = ~n14594 | ~n14593;
  assign n14602 = ~n14596 | ~n14595;
  assign n15491 = ~P1_STATE_REG_SCAN_IN & ~n14597;
  assign n14599 = ~n15360 | ~n15734;
  assign n14598 = ~n15358 | ~n9305;
  assign n14600 = ~n14599 | ~n14598;
  assign n14601 = ~n15491 & ~n14600;
  assign n14604 = ~n14602 | ~n14601;
  assign n14603 = ~n15381 & ~n15691;
  assign n14606 = ~n14604 & ~n14603;
  assign n14605 = ~n9297 | ~n15361;
  assign P1_U3236 = ~n14606 | ~n14605;
  assign n14609 = ~n14608 ^ n14607;
  assign n14619 = ~n14609 | ~n15376;
  assign n14617 = ~n14610 & ~n15333;
  assign n14615 = ~n15311 | ~n14939;
  assign n14611 = ~n15358 | ~n16391;
  assign n15588 = ~P1_REG3_REG_18__SCAN_IN | ~P1_U3086;
  assign n14613 = ~n14611 | ~n15588;
  assign n14612 = ~n15332 & ~n14998;
  assign n14614 = ~n14613 & ~n14612;
  assign n14616 = ~n14615 | ~n14614;
  assign n14618 = ~n14617 & ~n14616;
  assign P1_U3238 = ~n14619 | ~n14618;
  assign n14631 = ~n14756 & ~n15333;
  assign n14629 = ~n15311 | ~n14757;
  assign n14624 = n15332 | n14622;
  assign n14623 = ~P1_REG3_REG_26__SCAN_IN | ~P1_U3086;
  assign n14627 = ~n14624 | ~n14623;
  assign n14626 = ~n15319 & ~n14625;
  assign n14628 = ~n14627 & ~n14626;
  assign n14630 = ~n14629 | ~n14628;
  assign n14632 = ~n14631 & ~n14630;
  assign P1_U3240 = ~n14633 | ~n14632;
  assign n14637 = ~n14635 & ~n14634;
  assign n14638 = ~n14637 ^ n14636;
  assign n14647 = ~n14638 | ~n15376;
  assign n14645 = ~n15024 & ~n15333;
  assign n14643 = ~n15311 | ~n15025;
  assign n14639 = ~n15332 & ~n15012;
  assign n15547 = P1_U3086 & P1_REG3_REG_15__SCAN_IN;
  assign n14641 = n14639 | n15547;
  assign n14640 = ~n15319 & ~n15011;
  assign n14642 = ~n14641 & ~n14640;
  assign n14644 = ~n14643 | ~n14642;
  assign n14646 = ~n14645 & ~n14644;
  assign P1_U3241 = ~n14647 | ~n14646;
  assign n14648 = P1_ADDR_REG_19__SCAN_IN & n15607;
  assign n14675 = ~n14649 & ~n14648;
  assign n14672 = ~n10531 ^ P1_REG1_REG_19__SCAN_IN;
  assign n15603 = ~n16049;
  assign n14670 = ~n15603 | ~P1_REG1_REG_18__SCAN_IN;
  assign n15590 = ~n16049 ^ P1_REG1_REG_18__SCAN_IN;
  assign n14668 = ~P1_REG1_REG_17__SCAN_IN & ~n16056;
  assign n14666 = ~n16062 & ~P1_REG1_REG_16__SCAN_IN;
  assign n14661 = ~n16075 | ~P1_REG1_REG_14__SCAN_IN;
  assign n15535 = P1_REG1_REG_14__SCAN_IN ^ n16075;
  assign n14659 = ~n16081 | ~P1_REG1_REG_13__SCAN_IN;
  assign n14657 = ~n16088 & ~P1_REG1_REG_12__SCAN_IN;
  assign n15510 = ~P1_REG1_REG_12__SCAN_IN ^ n16088;
  assign n14655 = ~n16095 | ~P1_REG1_REG_11__SCAN_IN;
  assign n15496 = P1_REG1_REG_11__SCAN_IN ^ n16095;
  assign n14653 = ~n14651 | ~n14650;
  assign n14652 = ~n16101 | ~P1_REG1_REG_10__SCAN_IN;
  assign n15495 = ~n14653 | ~n14652;
  assign n14654 = ~n15496 | ~n15495;
  assign n15509 = ~n14655 | ~n14654;
  assign n14656 = ~n15510 & ~n15509;
  assign n15524 = ~n14657 & ~n14656;
  assign n15523 = P1_REG1_REG_13__SCAN_IN ^ n16081;
  assign n14658 = ~n15524 | ~n15523;
  assign n15534 = ~n14659 | ~n14658;
  assign n14660 = ~n15535 | ~n15534;
  assign n14662 = ~n14661 | ~n14660;
  assign n14664 = ~n16069 | ~n14662;
  assign n15550 = n16069 ^ n14662;
  assign n14663 = ~P1_REG1_REG_15__SCAN_IN | ~n15550;
  assign n15559 = ~n14664 | ~n14663;
  assign n15558 = ~P1_REG1_REG_16__SCAN_IN ^ n16062;
  assign n14665 = ~n15559 & ~n15558;
  assign n15578 = ~n14666 & ~n14665;
  assign n15579 = ~P1_REG1_REG_17__SCAN_IN ^ n16056;
  assign n14667 = ~n15578 & ~n15579;
  assign n15589 = ~n14668 & ~n14667;
  assign n14669 = ~n15590 | ~n15589;
  assign n14671 = ~n14670 | ~n14669;
  assign n14673 = ~n14672 ^ n14671;
  assign n14674 = ~n15591 | ~n14673;
  assign n14700 = ~n14675 | ~n14674;
  assign n15594 = ~n16049 ^ P1_REG2_REG_18__SCAN_IN;
  assign n14694 = ~P1_REG2_REG_17__SCAN_IN & ~n16056;
  assign n14692 = ~n16062 | ~P1_REG2_REG_16__SCAN_IN;
  assign n15564 = P1_REG2_REG_16__SCAN_IN ^ n16062;
  assign n14687 = ~n16075 | ~P1_REG2_REG_14__SCAN_IN;
  assign n15538 = P1_REG2_REG_14__SCAN_IN ^ n16075;
  assign n14685 = ~n16081 | ~P1_REG2_REG_13__SCAN_IN;
  assign n14683 = ~n16088 & ~P1_REG2_REG_12__SCAN_IN;
  assign n14681 = ~n16095 | ~P1_REG2_REG_11__SCAN_IN;
  assign n15493 = P1_REG2_REG_11__SCAN_IN ^ n16095;
  assign n14678 = ~n16101 | ~P1_REG2_REG_10__SCAN_IN;
  assign n15492 = ~n14679 | ~n14678;
  assign n14680 = ~n15493 | ~n15492;
  assign n15505 = ~n14681 | ~n14680;
  assign n15504 = ~P1_REG2_REG_12__SCAN_IN ^ n16088;
  assign n14682 = ~n15505 & ~n15504;
  assign n15520 = ~n14683 & ~n14682;
  assign n15521 = P1_REG2_REG_13__SCAN_IN ^ n16081;
  assign n14684 = ~n15520 | ~n15521;
  assign n15537 = ~n14685 | ~n14684;
  assign n14686 = ~n15538 | ~n15537;
  assign n14688 = ~n14687 | ~n14686;
  assign n14690 = ~n16069 | ~n14688;
  assign n15548 = n16069 ^ n14688;
  assign n14689 = ~P1_REG2_REG_15__SCAN_IN | ~n15548;
  assign n15563 = ~n14690 | ~n14689;
  assign n14691 = ~n15564 | ~n15563;
  assign n15573 = ~n14692 | ~n14691;
  assign n15572 = ~P1_REG2_REG_17__SCAN_IN ^ n16056;
  assign n14693 = ~n15573 & ~n15572;
  assign n15593 = ~n14694 & ~n14693;
  assign n15597 = ~n15594 | ~n15593;
  assign n14695 = ~n15603 | ~P1_REG2_REG_18__SCAN_IN;
  assign n14697 = ~n15597 | ~n14695;
  assign n14696 = P1_REG2_REG_19__SCAN_IN ^ n10531;
  assign n14698 = ~n14697 ^ n14696;
  assign n14699 = ~n14698 & ~n15596;
  assign n14702 = ~n14700 & ~n14699;
  assign n14701 = ~n15604 | ~n10531;
  assign P1_U3262 = ~n14702 | ~n14701;
  assign n14713 = ~n15035 | ~n15991;
  assign n14711 = ~n15036 & ~n15023;
  assign n14709 = ~n15961 | ~P1_REG2_REG_31__SCAN_IN;
  assign n14708 = ~n14707;
  assign n15044 = n14708 & n16427;
  assign n14714 = ~n16004 | ~n15044;
  assign n14710 = ~n14709 | ~n14714;
  assign n14712 = ~n14711 & ~n14710;
  assign P1_U3263 = ~n14713 | ~n14712;
  assign n15042 = ~n15043 ^ n8918;
  assign n14719 = ~n15042 | ~n15991;
  assign n14717 = ~n15043 & ~n15023;
  assign n14715 = ~n15961 | ~P1_REG2_REG_30__SCAN_IN;
  assign n14716 = ~n14715 | ~n14714;
  assign n14718 = ~n14717 & ~n14716;
  assign P1_U3264 = ~n14719 | ~n14718;
  assign n15747 = ~n15896;
  assign n14729 = ~n15050 & ~n15747;
  assign n15051 = ~n14720 ^ n15052;
  assign n14727 = ~n15051 | ~n15991;
  assign n14725 = ~n14721 & ~n15023;
  assign n14723 = ~n14722;
  assign n14724 = ~n15917 & ~n14723;
  assign n14726 = ~n14725 & ~n14724;
  assign n14728 = ~n14727 | ~n14726;
  assign n14740 = ~n14729 & ~n14728;
  assign n14732 = n14731 ^ n14730;
  assign n14736 = ~n14732 & ~n16170;
  assign n14734 = ~n16412 | ~n15979;
  assign n14733 = ~n16418 | ~n11990;
  assign n14735 = ~n14734 | ~n14733;
  assign n14738 = ~n15056 | ~n16004;
  assign n14737 = n16004 | P1_REG2_REG_27__SCAN_IN;
  assign n14739 = ~n14738 | ~n14737;
  assign P1_U3266 = ~n14740 | ~n14739;
  assign n15059 = n14746 ^ n14741;
  assign n14766 = ~n15059 | ~n15896;
  assign n14745 = n14742 | n14743;
  assign n14747 = ~n14745 | ~n14744;
  assign n14748 = ~n14747 ^ n14746;
  assign n14752 = ~n14748 | ~n15977;
  assign n14750 = ~n16409 | ~n15979;
  assign n14749 = ~n16415 | ~n11990;
  assign n14751 = n14750 & n14749;
  assign n15065 = ~n14752 | ~n14751;
  assign n14754 = n15065 | n15961;
  assign n14753 = n16004 | P1_REG2_REG_26__SCAN_IN;
  assign n14764 = ~n14754 | ~n14753;
  assign n15060 = ~n14755 ^ n14756;
  assign n14762 = ~n15060 | ~n15991;
  assign n14760 = n14756 | n15023;
  assign n14758 = ~n14757;
  assign n14759 = n15917 | n14758;
  assign n14761 = n14760 & n14759;
  assign n14763 = n14762 & n14761;
  assign n14765 = n14764 & n14763;
  assign P1_U3267 = ~n14766 | ~n14765;
  assign n15070 = ~n14767 ^ n14770;
  assign n14788 = ~n15070 | ~n15853;
  assign n14769 = n14742 | n14793;
  assign n14771 = n14769 & n14768;
  assign n14772 = ~n14771 ^ n14770;
  assign n14777 = ~n14772 | ~n15977;
  assign n14775 = ~n14817 & ~n15875;
  assign n14774 = ~n14773 & ~n15933;
  assign n14776 = ~n14775 & ~n14774;
  assign n15075 = ~n14777 | ~n14776;
  assign n14780 = ~n14779 ^ n14778;
  assign n16289 = ~n16327;
  assign n15073 = n14780 | n16289;
  assign n14785 = ~n15073 & ~n10531;
  assign n14783 = ~n15071 | ~n15927;
  assign n14782 = ~n16000 | ~n14781;
  assign n14784 = ~n14783 | ~n14782;
  assign n14786 = n14785 | n14784;
  assign n14787 = ~n15075 & ~n14786;
  assign n14789 = ~n14788 | ~n14787;
  assign n14791 = ~n14789 | ~n16004;
  assign n14790 = ~n15961 | ~P1_REG2_REG_25__SCAN_IN;
  assign P1_U3268 = ~n14791 | ~n14790;
  assign n15080 = n14792 ^ n14793;
  assign n14812 = ~n15080 | ~n15896;
  assign n14794 = ~n14742 ^ n14793;
  assign n14798 = n14794 | n16170;
  assign n14796 = ~n16403 | ~n15979;
  assign n14795 = ~n16409 | ~n11990;
  assign n14797 = n14796 & n14795;
  assign n15086 = ~n14798 | ~n14797;
  assign n14800 = ~n15086 & ~n15961;
  assign n14799 = ~n16004 & ~P1_REG2_REG_24__SCAN_IN;
  assign n14810 = ~n14800 & ~n14799;
  assign n15081 = ~n14801 ^ n15082;
  assign n14808 = ~n15081 | ~n15991;
  assign n14806 = ~n14802 & ~n15023;
  assign n14804 = ~n14803;
  assign n14805 = ~n15917 & ~n14804;
  assign n14807 = ~n14806 & ~n14805;
  assign n14809 = ~n14808 | ~n14807;
  assign n14811 = ~n14810 & ~n14809;
  assign P1_U3269 = ~n14812 | ~n14811;
  assign n15091 = n14813 ^ n14814;
  assign n14831 = ~n15091 | ~n15853;
  assign n14816 = ~n14815 ^ n14814;
  assign n14821 = ~n14816 | ~n15977;
  assign n14819 = ~n14865 & ~n15875;
  assign n14818 = ~n14817 & ~n15933;
  assign n14820 = ~n14819 & ~n14818;
  assign n15096 = ~n14821 | ~n14820;
  assign n14823 = ~n8985 ^ n14822;
  assign n15094 = ~n14823 | ~n16327;
  assign n14828 = ~n15094 & ~n10531;
  assign n14826 = ~n15092 | ~n15927;
  assign n14825 = ~n16000 | ~n14824;
  assign n14827 = ~n14826 | ~n14825;
  assign n14829 = n14828 | n14827;
  assign n14830 = ~n15096 & ~n14829;
  assign n14832 = ~n14831 | ~n14830;
  assign n14834 = ~n14832 | ~n16004;
  assign n14833 = ~n15961 | ~P1_REG2_REG_23__SCAN_IN;
  assign P1_U3270 = ~n14834 | ~n14833;
  assign n15101 = n14836 ^ n14835;
  assign n14845 = ~n15101 & ~n15983;
  assign n14838 = n14837 ^ n14836;
  assign n14843 = ~n14838 | ~n15977;
  assign n14841 = ~n14839 & ~n15933;
  assign n14840 = ~n14891 & ~n15875;
  assign n14842 = ~n14841 & ~n14840;
  assign n14844 = ~n14843 | ~n14842;
  assign n15108 = ~n14845 & ~n14844;
  assign n14847 = ~n15108 | ~n16004;
  assign n14846 = n16004 | P1_REG2_REG_22__SCAN_IN;
  assign n14859 = ~n14847 | ~n14846;
  assign n15675 = ~n14848;
  assign n15954 = ~n16004 | ~n15675;
  assign n14857 = ~n15101 & ~n15954;
  assign n14849 = ~n9006 | ~n15102;
  assign n14850 = n14849 & n16327;
  assign n15104 = ~n14850 | ~n8985;
  assign n14986 = ~n16004 | ~n16044;
  assign n14855 = ~n15104 & ~n14986;
  assign n14853 = ~n15102 | ~n15992;
  assign n14852 = ~n16000 | ~n14851;
  assign n14854 = ~n14853 | ~n14852;
  assign n14856 = n14855 | n14854;
  assign n14858 = ~n14857 & ~n14856;
  assign P1_U3271 = ~n14859 | ~n14858;
  assign n15111 = ~n14860 ^ n14861;
  assign n14872 = ~n15111 & ~n15983;
  assign n14864 = ~n14863 ^ n14862;
  assign n14870 = ~n14864 | ~n15977;
  assign n14868 = ~n14865 & ~n15933;
  assign n14867 = ~n14866 & ~n15875;
  assign n14869 = ~n14868 & ~n14867;
  assign n14871 = ~n14870 | ~n14869;
  assign n15119 = ~n14872 & ~n14871;
  assign n14874 = ~n15119 | ~n16004;
  assign n14873 = n16004 | P1_REG2_REG_21__SCAN_IN;
  assign n14886 = ~n14874 | ~n14873;
  assign n14884 = ~n15111 & ~n15954;
  assign n15112 = ~n14875 ^ n15113;
  assign n14882 = ~n15112 | ~n15991;
  assign n14880 = ~n14876 & ~n15023;
  assign n14878 = ~n14877;
  assign n14879 = ~n15917 & ~n14878;
  assign n14881 = ~n14880 & ~n14879;
  assign n14883 = ~n14882 | ~n14881;
  assign n14885 = ~n14884 & ~n14883;
  assign P1_U3272 = ~n14886 | ~n14885;
  assign n15122 = n14887 ^ n14888;
  assign n14907 = ~n15122 | ~n15896;
  assign n14890 = n14889 ^ n14888;
  assign n14895 = ~n14890 | ~n15977;
  assign n14893 = ~n14951 & ~n15875;
  assign n14892 = ~n14891 & ~n15933;
  assign n14894 = ~n14893 & ~n14892;
  assign n15128 = ~n14895 | ~n14894;
  assign n14897 = ~n15128 & ~n15961;
  assign n14896 = ~n16004 & ~P1_REG2_REG_20__SCAN_IN;
  assign n14905 = ~n14897 & ~n14896;
  assign n15123 = ~n14923 ^ n9573;
  assign n14903 = ~n15123 | ~n15991;
  assign n14901 = ~n9573 & ~n15023;
  assign n14899 = ~n14898;
  assign n14900 = ~n15917 & ~n14899;
  assign n14902 = ~n14901 & ~n14900;
  assign n14904 = ~n14903 | ~n14902;
  assign n14906 = ~n14905 & ~n14904;
  assign P1_U3273 = ~n14907 | ~n14906;
  assign n15133 = ~n14908 ^ n14911;
  assign n14934 = ~n15133 | ~n15896;
  assign n14910 = ~n14947 | ~n14909;
  assign n14913 = ~n14910 | ~n14935;
  assign n14912 = ~n14911;
  assign n14914 = ~n14913 ^ n14912;
  assign n14918 = n14914 | n16170;
  assign n14916 = ~n16388 | ~n15979;
  assign n14915 = ~n16394 | ~n11990;
  assign n14917 = n14916 & n14915;
  assign n15139 = ~n14918 | ~n14917;
  assign n14920 = n15139 | n15961;
  assign n14919 = n16004 | P1_REG2_REG_19__SCAN_IN;
  assign n14932 = ~n14920 | ~n14919;
  assign n14922 = ~n14921 | ~n15135;
  assign n15134 = n14923 & n14922;
  assign n14930 = ~n15134 | ~n15991;
  assign n14928 = ~n14924 & ~n15023;
  assign n14926 = ~n14925;
  assign n14927 = ~n15917 & ~n14926;
  assign n14929 = ~n14928 & ~n14927;
  assign n14931 = n14930 & n14929;
  assign n14933 = n14932 & n14931;
  assign P1_U3274 = ~n14934 | ~n14933;
  assign n14948 = ~n14936 | ~n14935;
  assign n15144 = n14948 ^ n14937;
  assign n14945 = ~n15144 | ~n15896;
  assign n15145 = ~n14938 ^ n15146;
  assign n14943 = n15145 & n15991;
  assign n14941 = ~n15146 | ~n15992;
  assign n14940 = ~n16000 | ~n14939;
  assign n14942 = ~n14941 | ~n14940;
  assign n14944 = ~n14943 & ~n14942;
  assign n14959 = ~n14945 | ~n14944;
  assign n14949 = ~n14947 | ~n14946;
  assign n14950 = ~n14949 ^ n14948;
  assign n14955 = ~n14950 | ~n15977;
  assign n14953 = ~n14951 & ~n15933;
  assign n14952 = ~n14998 & ~n15875;
  assign n14954 = ~n14953 & ~n14952;
  assign n15150 = ~n14955 | ~n14954;
  assign n14957 = ~n15150 & ~n15961;
  assign n14956 = ~n16004 & ~P1_REG2_REG_18__SCAN_IN;
  assign n14958 = ~n14957 & ~n14956;
  assign P1_U3275 = n14959 | n14958;
  assign n14969 = ~n14961 ^ n14998;
  assign n15155 = ~n14960 ^ n14969;
  assign n14968 = ~n15155 | ~n15896;
  assign n15156 = ~n14984 ^ n14961;
  assign n14966 = n15156 & n15991;
  assign n14964 = ~n15992 | ~n15157;
  assign n14963 = ~n16000 | ~n14962;
  assign n14965 = ~n14964 | ~n14963;
  assign n14967 = ~n14966 & ~n14965;
  assign n14980 = ~n14968 | ~n14967;
  assign n14971 = ~n14970 ^ n14969;
  assign n14976 = ~n14971 | ~n15977;
  assign n14974 = ~n14972 & ~n15933;
  assign n14973 = ~n15011 & ~n15875;
  assign n14975 = ~n14974 & ~n14973;
  assign n15161 = ~n14976 | ~n14975;
  assign n14978 = ~n15161 & ~n15961;
  assign n14977 = ~n16004 & ~P1_REG2_REG_17__SCAN_IN;
  assign n14979 = ~n14978 & ~n14977;
  assign P1_U3276 = n14980 | n14979;
  assign n15166 = n14981 ^ n14994;
  assign n14993 = ~n15166 | ~n15896;
  assign n14983 = ~n14982 | ~n15167;
  assign n14985 = n14983 & n16327;
  assign n15169 = ~n14985 | ~n14984;
  assign n14991 = ~n15169 & ~n14986;
  assign n14989 = ~n15992 | ~n15167;
  assign n14988 = ~n16000 | ~n14987;
  assign n14990 = ~n14989 | ~n14988;
  assign n14992 = ~n14991 & ~n14990;
  assign n15006 = ~n14993 | ~n14992;
  assign n14996 = n14995 ^ n14994;
  assign n15002 = ~n14996 | ~n15977;
  assign n15000 = ~n14997 & ~n15875;
  assign n14999 = ~n14998 & ~n15933;
  assign n15001 = ~n15000 & ~n14999;
  assign n15171 = ~n15002 | ~n15001;
  assign n15004 = ~n15171 & ~n15961;
  assign n15003 = ~n16004 & ~P1_REG2_REG_16__SCAN_IN;
  assign n15005 = ~n15004 & ~n15003;
  assign P1_U3277 = n15006 | n15005;
  assign n15176 = ~n15007 ^ n15008;
  assign n15018 = ~n15176 & ~n15983;
  assign n15010 = n15009 ^ n15008;
  assign n15016 = ~n15010 | ~n15977;
  assign n15014 = ~n15011 & ~n15933;
  assign n15013 = ~n15012 & ~n15875;
  assign n15015 = ~n15014 & ~n15013;
  assign n15017 = ~n15016 | ~n15015;
  assign n15184 = ~n15018 & ~n15017;
  assign n15021 = ~n15184 | ~n16004;
  assign n15019 = ~P1_REG2_REG_15__SCAN_IN;
  assign n15020 = ~n15961 | ~n15019;
  assign n15034 = ~n15021 | ~n15020;
  assign n15032 = ~n15176 & ~n15954;
  assign n15177 = ~n15022 ^ n15024;
  assign n15030 = ~n15177 | ~n15991;
  assign n15028 = ~n15024 & ~n15023;
  assign n15026 = ~n15025;
  assign n15027 = ~n15917 & ~n15026;
  assign n15029 = ~n15028 & ~n15027;
  assign n15031 = ~n15030 | ~n15029;
  assign n15033 = ~n15032 & ~n15031;
  assign P1_U3278 = ~n15034 | ~n15033;
  assign n15039 = ~n15035 | ~n16327;
  assign n16291 = ~n16329;
  assign n15037 = ~n15036 & ~n16291;
  assign n15038 = ~n15037 & ~n15044;
  assign n15187 = ~n15039 | ~n15038;
  assign n15041 = ~n15187 | ~n16385;
  assign n15040 = ~n16383 | ~P1_REG1_REG_31__SCAN_IN;
  assign P1_U3553 = ~n15041 | ~n15040;
  assign n15047 = ~n15042 | ~n16327;
  assign n15045 = ~n15043 & ~n16291;
  assign n15046 = ~n15045 & ~n15044;
  assign n15190 = ~n15047 | ~n15046;
  assign n15049 = ~n15190 | ~n16385;
  assign n15048 = ~n16383 | ~P1_REG1_REG_30__SCAN_IN;
  assign P1_U3552 = ~n15049 | ~n15048;
  assign n16318 = ~n16225;
  assign n15054 = ~n15051 | ~n16327;
  assign n15053 = ~n15052 | ~n16329;
  assign n15055 = ~n15054 | ~n15053;
  assign n15058 = ~n15193 | ~n16385;
  assign n15057 = ~n16383 | ~P1_REG1_REG_27__SCAN_IN;
  assign P1_U3549 = ~n15058 | ~n15057;
  assign n15067 = ~n15059 | ~n16225;
  assign n15063 = ~n15060 | ~n16327;
  assign n15062 = ~n15061 | ~n16329;
  assign n15064 = ~n15063 | ~n15062;
  assign n15066 = ~n15065 & ~n15064;
  assign n15196 = ~n15067 | ~n15066;
  assign n15069 = ~n15196 | ~n16385;
  assign n15068 = ~n16383 | ~P1_REG1_REG_26__SCAN_IN;
  assign P1_U3548 = ~n15069 | ~n15068;
  assign n15077 = ~n15070 | ~n16225;
  assign n15072 = ~n15071 | ~n16329;
  assign n15074 = ~n15073 | ~n15072;
  assign n15199 = ~n15077 | ~n15076;
  assign n15079 = ~n15199 | ~n16385;
  assign n15078 = ~n16383 | ~P1_REG1_REG_25__SCAN_IN;
  assign P1_U3547 = ~n15079 | ~n15078;
  assign n15088 = ~n15080 | ~n16225;
  assign n15084 = ~n15081 | ~n16327;
  assign n15083 = ~n15082 | ~n16329;
  assign n15085 = ~n15084 | ~n15083;
  assign n15087 = ~n15086 & ~n15085;
  assign n15202 = ~n15088 | ~n15087;
  assign n15090 = ~n15202 | ~n16385;
  assign n15089 = ~n16383 | ~P1_REG1_REG_24__SCAN_IN;
  assign P1_U3546 = ~n15090 | ~n15089;
  assign n15098 = ~n15091 | ~n16225;
  assign n15093 = ~n15092 | ~n16329;
  assign n15095 = ~n15094 | ~n15093;
  assign n15097 = ~n15096 & ~n15095;
  assign n15205 = ~n15098 | ~n15097;
  assign n15100 = ~n15205 | ~n16385;
  assign n15099 = ~n16383 | ~P1_REG1_REG_23__SCAN_IN;
  assign P1_U3545 = ~n15100 | ~n15099;
  assign n15106 = ~n15101 & ~n16295;
  assign n15103 = ~n15102 | ~n16329;
  assign n15105 = ~n15104 | ~n15103;
  assign n15107 = ~n15106 & ~n15105;
  assign n15208 = ~n15108 | ~n15107;
  assign n15110 = ~n15208 | ~n16385;
  assign n15109 = ~n16383 | ~P1_REG1_REG_22__SCAN_IN;
  assign P1_U3544 = ~n15110 | ~n15109;
  assign n15117 = ~n15111 & ~n16295;
  assign n15115 = ~n15112 | ~n16327;
  assign n15114 = ~n15113 | ~n16329;
  assign n15116 = ~n15115 | ~n15114;
  assign n15118 = ~n15117 & ~n15116;
  assign n15211 = ~n15119 | ~n15118;
  assign n15121 = ~n15211 | ~n16385;
  assign n15120 = ~n16383 | ~P1_REG1_REG_21__SCAN_IN;
  assign P1_U3543 = ~n15121 | ~n15120;
  assign n15130 = ~n15122 | ~n16225;
  assign n15126 = ~n15123 | ~n16327;
  assign n15125 = ~n15124 | ~n16329;
  assign n15127 = ~n15126 | ~n15125;
  assign n15129 = ~n15128 & ~n15127;
  assign n15214 = ~n15130 | ~n15129;
  assign n15132 = ~n15214 | ~n16385;
  assign n15131 = ~n16383 | ~P1_REG1_REG_20__SCAN_IN;
  assign P1_U3542 = ~n15132 | ~n15131;
  assign n15141 = ~n15133 | ~n16225;
  assign n15137 = ~n15134 | ~n16327;
  assign n15136 = ~n15135 | ~n16329;
  assign n15138 = ~n15137 | ~n15136;
  assign n15140 = ~n15139 & ~n15138;
  assign n15217 = ~n15141 | ~n15140;
  assign n15143 = ~n15217 | ~n16385;
  assign n15142 = ~n16383 | ~P1_REG1_REG_19__SCAN_IN;
  assign P1_U3541 = ~n15143 | ~n15142;
  assign n15152 = ~n15144 | ~n16225;
  assign n15148 = ~n15145 | ~n16327;
  assign n15147 = ~n15146 | ~n16329;
  assign n15149 = ~n15148 | ~n15147;
  assign n15151 = ~n15150 & ~n15149;
  assign n15220 = ~n15152 | ~n15151;
  assign n15154 = ~n15220 | ~n16385;
  assign n15153 = ~n16383 | ~P1_REG1_REG_18__SCAN_IN;
  assign P1_U3540 = ~n15154 | ~n15153;
  assign n15163 = ~n15155 | ~n16225;
  assign n15159 = ~n15156 | ~n16327;
  assign n15158 = ~n15157 | ~n16329;
  assign n15160 = ~n15159 | ~n15158;
  assign n15162 = ~n15161 & ~n15160;
  assign n15223 = ~n15163 | ~n15162;
  assign n15165 = ~n15223 | ~n16385;
  assign n15164 = ~n16383 | ~P1_REG1_REG_17__SCAN_IN;
  assign P1_U3539 = ~n15165 | ~n15164;
  assign n15173 = ~n15166 | ~n16225;
  assign n15168 = ~n15167 | ~n16329;
  assign n15170 = ~n15169 | ~n15168;
  assign n15172 = ~n15171 & ~n15170;
  assign n15226 = ~n15173 | ~n15172;
  assign n15175 = ~n15226 | ~n16385;
  assign n15174 = ~n16383 | ~P1_REG1_REG_16__SCAN_IN;
  assign P1_U3538 = ~n15175 | ~n15174;
  assign n15182 = ~n15176 & ~n16295;
  assign n15180 = ~n15177 | ~n16327;
  assign n15179 = ~n15178 | ~n16329;
  assign n15181 = ~n15180 | ~n15179;
  assign n15183 = ~n15182 & ~n15181;
  assign n15229 = ~n15184 | ~n15183;
  assign n15186 = ~n15229 | ~n16385;
  assign n15185 = ~n16383 | ~P1_REG1_REG_15__SCAN_IN;
  assign P1_U3537 = ~n15186 | ~n15185;
  assign n15189 = ~n15187 | ~n16338;
  assign n15188 = ~n16326 | ~P1_REG0_REG_31__SCAN_IN;
  assign P1_U3521 = ~n15189 | ~n15188;
  assign n15192 = ~n15190 | ~n16338;
  assign n15191 = ~n16326 | ~P1_REG0_REG_30__SCAN_IN;
  assign P1_U3520 = ~n15192 | ~n15191;
  assign n15194 = ~n16326 | ~P1_REG0_REG_27__SCAN_IN;
  assign P1_U3517 = ~n15195 | ~n15194;
  assign n15198 = ~n15196 | ~n16338;
  assign n15197 = ~n16326 | ~P1_REG0_REG_26__SCAN_IN;
  assign P1_U3516 = ~n15198 | ~n15197;
  assign n15201 = ~n15199 | ~n16338;
  assign n15200 = ~n16326 | ~P1_REG0_REG_25__SCAN_IN;
  assign P1_U3515 = ~n15201 | ~n15200;
  assign n15204 = ~n15202 | ~n16338;
  assign n15203 = ~n16326 | ~P1_REG0_REG_24__SCAN_IN;
  assign P1_U3514 = ~n15204 | ~n15203;
  assign n15207 = ~n15205 | ~n16338;
  assign n15206 = ~n16326 | ~P1_REG0_REG_23__SCAN_IN;
  assign P1_U3513 = ~n15207 | ~n15206;
  assign n15210 = ~n15208 | ~n16338;
  assign n15209 = ~n16326 | ~P1_REG0_REG_22__SCAN_IN;
  assign P1_U3512 = ~n15210 | ~n15209;
  assign n15213 = ~n15211 | ~n16338;
  assign n15212 = ~n16326 | ~P1_REG0_REG_21__SCAN_IN;
  assign P1_U3511 = ~n15213 | ~n15212;
  assign n15216 = ~n15214 | ~n16338;
  assign n15215 = ~n16326 | ~P1_REG0_REG_20__SCAN_IN;
  assign P1_U3510 = ~n15216 | ~n15215;
  assign n15219 = ~n15217 | ~n16338;
  assign n15218 = ~n16326 | ~P1_REG0_REG_19__SCAN_IN;
  assign P1_U3509 = ~n15219 | ~n15218;
  assign n15222 = ~n15220 | ~n16338;
  assign n15221 = ~n16326 | ~P1_REG0_REG_18__SCAN_IN;
  assign P1_U3507 = ~n15222 | ~n15221;
  assign n15225 = ~n15223 | ~n16338;
  assign n15224 = ~n16326 | ~P1_REG0_REG_17__SCAN_IN;
  assign P1_U3504 = ~n15225 | ~n15224;
  assign n15228 = ~n15226 | ~n16338;
  assign n15227 = ~n16326 | ~P1_REG0_REG_16__SCAN_IN;
  assign P1_U3501 = ~n15228 | ~n15227;
  assign n15231 = ~n15229 | ~n16338;
  assign n15230 = ~n16326 | ~P1_REG0_REG_15__SCAN_IN;
  assign P1_U3498 = ~n15231 | ~n15230;
  assign n15240 = ~n15232 & ~n16154;
  assign n15234 = n15233 & P1_IR_REG_31__SCAN_IN;
  assign n15235 = ~n15234 | ~P1_STATE_REG_SCAN_IN;
  assign n15238 = n15236 | n15235;
  assign n16159 = ~n16023;
  assign n15237 = ~n16159 | ~P2_DATAO_REG_31__SCAN_IN;
  assign n15239 = ~n15238 | ~n15237;
  assign P1_U3324 = n15240 | n15239;
  assign n15242 = ~n15241;
  assign n15247 = ~n15242 | ~n16134;
  assign n15245 = ~n9906 & ~P1_U3086;
  assign n15244 = ~n16023 & ~n15243;
  assign n15246 = ~n15245 & ~n15244;
  assign P1_U3325 = ~n15247 | ~n15246;
  assign U123 = ~P1_WR_REG_SCAN_IN ^ P2_WR_REG_SCAN_IN;
  assign U126 = ~P2_RD_REG_SCAN_IN ^ P1_RD_REG_SCAN_IN;
  assign n15249 = ~n15360 | ~n15844;
  assign n15248 = ~n15361 | ~n11963;
  assign n15257 = ~n15249 | ~n15248;
  assign n15252 = ~n15250;
  assign n15253 = ~n15252 & ~n15251;
  assign n15255 = ~n15254 ^ n15253;
  assign n15256 = ~n15255 & ~n15293;
  assign n15263 = ~n15257 & ~n15256;
  assign n15261 = ~n15311 | ~n15781;
  assign n15259 = n15319 | n15790;
  assign n15260 = n15259 & n15258;
  assign n15262 = n15261 & n15260;
  assign P1_U3213 = ~n15263 | ~n15262;
  assign n15265 = ~n15360 | ~n11910;
  assign n15264 = ~n15361 | ~n9323;
  assign n15271 = ~n15265 | ~n15264;
  assign n15267 = ~n15306 | ~n15266;
  assign n15269 = ~n15268 ^ n15267;
  assign n15270 = ~n15269 & ~n15293;
  assign n15277 = ~n15271 & ~n15270;
  assign n15273 = ~n15358 | ~n11903;
  assign n15275 = ~n15273 | ~n15272;
  assign n15274 = ~P1_REG3_REG_3__SCAN_IN & ~n15381;
  assign n15276 = ~n15275 & ~n15274;
  assign P1_U3218 = ~n15277 | ~n15276;
  assign n15279 = ~n15358 | ~n15771;
  assign n15283 = ~n15279 | ~n15278;
  assign n15281 = ~n15360 | ~n15823;
  assign n15280 = ~n15361 | ~n16258;
  assign n15282 = ~n15281 | ~n15280;
  assign n15291 = ~n15283 & ~n15282;
  assign n15323 = ~n15284 ^ n15285;
  assign n15287 = ~n15323 ^ n15286;
  assign n15289 = ~n15287 & ~n15293;
  assign n15288 = ~n15381 & ~n15754;
  assign n15290 = ~n15289 & ~n15288;
  assign P1_U3221 = ~n15291 | ~n15290;
  assign n15292 = ~n15319 & ~n15801;
  assign n15464 = P1_U3086 & P1_REG3_REG_5__SCAN_IN;
  assign n15302 = ~n15292 & ~n15464;
  assign n15367 = ~n15369 ^ n15368;
  assign n15294 = n15366 ^ n15367;
  assign n15300 = ~n15294 & ~n15293;
  assign n15298 = ~n15311 | ~n15858;
  assign n15901 = ~n11903;
  assign n15296 = n15332 | n15901;
  assign n15295 = ~n15361 | ~n16227;
  assign n15297 = n15296 & n15295;
  assign n15299 = ~n15298 | ~n15297;
  assign n15301 = ~n15300 & ~n15299;
  assign P1_U3227 = ~n15302 | ~n15301;
  assign n15304 = ~n15332 & ~n15934;
  assign n15303 = ~n15333 & ~n15882;
  assign n15317 = ~n15304 & ~n15303;
  assign n15305 = ~n15358 | ~n15876;
  assign n15444 = ~P1_REG3_REG_4__SCAN_IN | ~P1_U3086;
  assign n15315 = ~n15305 | ~n15444;
  assign n15309 = ~n15307 | ~n15306;
  assign n15310 = ~n15308 ^ n15309;
  assign n15313 = ~n15310 | ~n15376;
  assign n15312 = ~n15311 | ~n15865;
  assign n15314 = ~n15313 | ~n15312;
  assign n15316 = ~n15315 & ~n15314;
  assign P1_U3230 = ~n15317 | ~n15316;
  assign n15321 = ~n15319 & ~n15318;
  assign n15341 = ~n15321 & ~n15320;
  assign n15326 = ~n15323 | ~n15322;
  assign n15325 = ~n15284 | ~n15324;
  assign n15330 = ~n15326 | ~n15325;
  assign n15329 = ~n15328 ^ n15327;
  assign n15331 = ~n15330 ^ n15329;
  assign n15337 = ~n15331 | ~n15376;
  assign n15335 = ~n15332 & ~n15790;
  assign n15334 = ~n16271 & ~n15333;
  assign n15336 = ~n15335 & ~n15334;
  assign n15339 = ~n15337 | ~n15336;
  assign n15338 = ~n15381 & ~n15741;
  assign n15340 = ~n15339 & ~n15338;
  assign P1_U3231 = ~n15341 | ~n15340;
  assign n15343 = ~n15360 | ~n9310;
  assign n15342 = ~n15361 | ~n16193;
  assign n15354 = ~n15343 | ~n15342;
  assign n15349 = ~n15345 | ~n15344;
  assign n15348 = ~n15347 | ~n15346;
  assign n15350 = n15349 ^ n15348;
  assign n15352 = ~n15350 | ~n15376;
  assign n15351 = ~n15358 | ~n11905;
  assign n15353 = ~n15352 | ~n15351;
  assign n15357 = ~n15354 & ~n15353;
  assign n15356 = ~P1_REG3_REG_2__SCAN_IN | ~n15355;
  assign P1_U3237 = ~n15357 | ~n15356;
  assign n15359 = ~n15358 | ~n15823;
  assign n15476 = ~P1_REG3_REG_6__SCAN_IN | ~P1_U3086;
  assign n15365 = ~n15359 | ~n15476;
  assign n15363 = ~n15360 | ~n15876;
  assign n15362 = ~n15361 | ~n9550;
  assign n15364 = ~n15363 | ~n15362;
  assign n15385 = ~n15365 & ~n15364;
  assign n15371 = ~n15367 & ~n15366;
  assign n15370 = ~n15369 & ~n15368;
  assign n15375 = ~n15371 & ~n15370;
  assign n15374 = n15373 & n15372;
  assign n15379 = ~n15375 & ~n15374;
  assign n15377 = ~n15375 | ~n15374;
  assign n15378 = ~n15377 | ~n15376;
  assign n15383 = ~n15379 & ~n15378;
  assign n15826 = ~n15380;
  assign n15382 = ~n15381 & ~n15826;
  assign n15384 = ~n15383 & ~n15382;
  assign P1_U3239 = ~n15385 | ~n15384;
  assign n15388 = ~n15432 | ~P1_REG2_REG_0__SCAN_IN;
  assign n15387 = ~n15386 | ~P1_REG1_REG_0__SCAN_IN;
  assign n15389 = ~n15388 | ~n15387;
  assign n15390 = ~n15389 | ~n15426;
  assign n15391 = ~n15423 ^ n15390;
  assign n15394 = ~n15392 & ~n15391;
  assign n15393 = P1_U3086 & P1_REG3_REG_0__SCAN_IN;
  assign n15396 = ~n15394 & ~n15393;
  assign n15395 = ~n15607 | ~P1_ADDR_REG_0__SCAN_IN;
  assign P1_U3243 = ~n15396 | ~n15395;
  assign n15398 = ~P1_ADDR_REG_1__SCAN_IN | ~n15607;
  assign n15397 = ~P1_REG3_REG_1__SCAN_IN | ~P1_U3086;
  assign n15405 = ~n15398 | ~n15397;
  assign n15401 = n15400 ^ n15399;
  assign n15403 = ~n15574 | ~n15401;
  assign n15402 = ~n15604 | ~n16155;
  assign n15404 = ~n15403 | ~n15402;
  assign n15413 = ~n15405 & ~n15404;
  assign n15410 = ~n15406;
  assign n15409 = ~n15408 & ~n15407;
  assign n15411 = ~n15410 & ~n15409;
  assign n15412 = ~n15591 | ~n15411;
  assign P1_U3244 = ~n15413 | ~n15412;
  assign n15415 = ~P1_ADDR_REG_2__SCAN_IN | ~n15607;
  assign n15414 = ~P1_REG3_REG_2__SCAN_IN | ~P1_U3086;
  assign n15422 = ~n15415 | ~n15414;
  assign n15420 = ~n15604 | ~n16148;
  assign n15418 = n15417 ^ n15416;
  assign n15419 = ~n15591 | ~n15418;
  assign n15421 = ~n15420 | ~n15419;
  assign n15442 = ~n15422 & ~n15421;
  assign n15424 = ~n15423 | ~P1_REG2_REG_0__SCAN_IN;
  assign n15425 = ~n15432 | ~n15424;
  assign n15429 = ~n15425 | ~n15426;
  assign n15427 = ~n15426 | ~P1_REG2_REG_0__SCAN_IN;
  assign n15428 = ~n15427 | ~P1_IR_REG_0__SCAN_IN;
  assign n15430 = ~n15429 | ~n15428;
  assign n15436 = ~n15430 | ~P1_U3973;
  assign n15433 = ~n15432 & ~n15431;
  assign n15435 = n15434 & n15433;
  assign n15456 = ~n15436 & ~n15435;
  assign n15439 = ~n15438 ^ n15437;
  assign n15440 = ~n15596 & ~n15439;
  assign n15441 = ~n15456 & ~n15440;
  assign P1_U3245 = ~n15442 | ~n15441;
  assign n15443 = ~n15607 | ~P1_ADDR_REG_4__SCAN_IN;
  assign n15451 = ~n15444 | ~n15443;
  assign n15449 = ~n15604 | ~n16136;
  assign n15447 = n15446 ^ n15445;
  assign n15448 = ~n15591 | ~n15447;
  assign n15450 = ~n15449 | ~n15448;
  assign n15458 = ~n15451 & ~n15450;
  assign n15454 = ~n15453 ^ n15452;
  assign n15455 = ~n15596 & ~n15454;
  assign n15457 = ~n15456 & ~n15455;
  assign P1_U3247 = ~n15458 | ~n15457;
  assign n15461 = ~n15460 ^ n15459;
  assign n15469 = ~n15596 & ~n15461;
  assign n15463 = ~n15607;
  assign n15462 = ~P1_ADDR_REG_5__SCAN_IN;
  assign n15465 = ~n15463 & ~n15462;
  assign n15467 = ~n15465 & ~n15464;
  assign n15466 = ~n15604 | ~n16128;
  assign n15468 = ~n15467 | ~n15466;
  assign n15474 = ~n15469 & ~n15468;
  assign n15472 = n15471 ^ n15470;
  assign n15473 = ~n15591 | ~n15472;
  assign P1_U3248 = ~n15474 | ~n15473;
  assign n15475 = ~n15607 | ~P1_ADDR_REG_6__SCAN_IN;
  assign n15484 = ~n15476 | ~n15475;
  assign n15482 = ~n15604 | ~n15477;
  assign n15480 = n15479 ^ n15478;
  assign n15481 = ~n15591 | ~n15480;
  assign n15483 = ~n15482 | ~n15481;
  assign n15489 = ~n15484 & ~n15483;
  assign n15487 = n15486 ^ n15485;
  assign n15488 = ~n15574 | ~n15487;
  assign P1_U3249 = ~n15489 | ~n15488;
  assign n15490 = n15607 & P1_ADDR_REG_11__SCAN_IN;
  assign n15503 = ~n15491 & ~n15490;
  assign n15494 = ~n15493 ^ n15492;
  assign n15501 = ~n15596 & ~n15494;
  assign n15497 = n15496 ^ n15495;
  assign n15499 = ~n15497 | ~n15591;
  assign n15498 = ~n15604 | ~n16095;
  assign n15500 = ~n15499 | ~n15498;
  assign n15502 = ~n15501 & ~n15500;
  assign P1_U3254 = ~n15503 | ~n15502;
  assign n15506 = ~n15505 ^ n15504;
  assign n15517 = ~n15506 | ~n15574;
  assign n15507 = ~n15607 | ~P1_ADDR_REG_12__SCAN_IN;
  assign n15515 = ~n15508 | ~n15507;
  assign n15513 = ~n15604 | ~n16088;
  assign n15511 = ~n15510 ^ n15509;
  assign n15512 = ~n15511 | ~n15591;
  assign n15514 = ~n15513 | ~n15512;
  assign n15516 = ~n15515 & ~n15514;
  assign P1_U3255 = ~n15517 | ~n15516;
  assign n15518 = n15607 & P1_ADDR_REG_13__SCAN_IN;
  assign n15531 = ~n15519 & ~n15518;
  assign n15522 = ~n15521 ^ n15520;
  assign n15529 = ~n15596 & ~n15522;
  assign n15525 = n15524 ^ n15523;
  assign n15527 = ~n15525 | ~n15591;
  assign n15526 = ~n15604 | ~n16081;
  assign n15528 = ~n15527 | ~n15526;
  assign n15530 = ~n15529 & ~n15528;
  assign P1_U3256 = ~n15531 | ~n15530;
  assign n15532 = ~n15607 | ~P1_ADDR_REG_14__SCAN_IN;
  assign n15543 = ~n15533 | ~n15532;
  assign n15536 = n15535 ^ n15534;
  assign n15541 = ~n15536 | ~n15591;
  assign n15539 = n15538 ^ n15537;
  assign n15540 = ~n15539 | ~n15574;
  assign n15542 = ~n15541 | ~n15540;
  assign n15545 = ~n15543 & ~n15542;
  assign n15544 = ~n15604 | ~n16075;
  assign P1_U3257 = ~n15545 | ~n15544;
  assign n15546 = n15607 & P1_ADDR_REG_15__SCAN_IN;
  assign n15557 = ~n15547 & ~n15546;
  assign n15549 = ~n15548 ^ P1_REG2_REG_15__SCAN_IN;
  assign n15555 = ~n15596 & ~n15549;
  assign n15551 = P1_REG1_REG_15__SCAN_IN ^ n15550;
  assign n15553 = ~n15551 | ~n15591;
  assign n15552 = ~n15604 | ~n16069;
  assign n15554 = ~n15553 | ~n15552;
  assign n15556 = ~n15555 & ~n15554;
  assign P1_U3258 = ~n15557 | ~n15556;
  assign n15560 = ~n15559 ^ n15558;
  assign n15571 = ~n15560 | ~n15591;
  assign n15561 = ~n15607 | ~P1_ADDR_REG_16__SCAN_IN;
  assign n15569 = ~n15562 | ~n15561;
  assign n15565 = n15564 ^ n15563;
  assign n15567 = ~n15565 | ~n15574;
  assign n15566 = ~n15604 | ~n16062;
  assign n15568 = ~n15567 | ~n15566;
  assign n15570 = ~n15569 & ~n15568;
  assign P1_U3259 = ~n15571 | ~n15570;
  assign n15575 = ~n15573 ^ n15572;
  assign n15586 = ~n15575 | ~n15574;
  assign n15576 = ~n15607 | ~P1_ADDR_REG_17__SCAN_IN;
  assign n15584 = ~n15577 | ~n15576;
  assign n15580 = ~n15579 ^ n15578;
  assign n15582 = ~n15580 | ~n15591;
  assign n15581 = ~n15604 | ~n16056;
  assign n15583 = ~n15582 | ~n15581;
  assign n15585 = ~n15584 & ~n15583;
  assign P1_U3260 = ~n15586 | ~n15585;
  assign n15587 = ~n15607 | ~P1_ADDR_REG_18__SCAN_IN;
  assign n15602 = ~n15588 | ~n15587;
  assign n15592 = n15590 ^ n15589;
  assign n15600 = ~n15592 | ~n15591;
  assign n15595 = ~n15594 & ~n15593;
  assign n15598 = ~n15596 & ~n15595;
  assign n15599 = ~n15598 | ~n15597;
  assign n15601 = ~n15600 | ~n15599;
  assign n15606 = ~n15602 & ~n15601;
  assign n15605 = ~n15604 | ~n15603;
  assign P1_U3261 = ~n15606 | ~n15605;
  assign P1_U3085 = ~n15607 & ~P1_U3973;
  assign n15609 = ~n15992 | ~n9555;
  assign n15608 = ~n15961 | ~P1_REG2_REG_14__SCAN_IN;
  assign n15612 = ~n15609 | ~n15608;
  assign n15611 = ~n15917 & ~n15610;
  assign n15631 = ~n15612 & ~n15611;
  assign n16328 = ~n15613 ^ n9555;
  assign n15626 = ~n16328 | ~n15991;
  assign n15627 = ~n15615 ^ n15614;
  assign n16335 = ~n15627;
  assign n15942 = ~n15983;
  assign n15624 = ~n16335 | ~n15942;
  assign n15617 = ~n15616 ^ n15615;
  assign n15622 = ~n15617 & ~n16170;
  assign n15620 = ~n15661 | ~n15979;
  assign n15619 = ~n15618 | ~n11990;
  assign n15621 = ~n15620 | ~n15619;
  assign n15623 = ~n15622 & ~n15621;
  assign n16333 = ~n15624 | ~n15623;
  assign n15625 = ~n16333 | ~n16004;
  assign n15629 = ~n15626 | ~n15625;
  assign n15628 = ~n15627 & ~n15954;
  assign n15630 = ~n15629 & ~n15628;
  assign P1_U3279 = ~n15631 | ~n15630;
  assign n15633 = ~n15992 | ~n16315;
  assign n15632 = ~n15961 | ~P1_REG2_REG_13__SCAN_IN;
  assign n15636 = ~n15633 | ~n15632;
  assign n15635 = ~n15917 & ~n15634;
  assign n15653 = ~n15636 & ~n15635;
  assign n16314 = ~n15637 ^ n15638;
  assign n15651 = ~n16314 | ~n15991;
  assign n16319 = n15639 ^ n15643;
  assign n15649 = ~n16319 & ~n15747;
  assign n15642 = ~n9305 | ~n15979;
  assign n15641 = ~n15640 | ~n11990;
  assign n15647 = ~n15642 | ~n15641;
  assign n15645 = n15644 ^ n15643;
  assign n15646 = ~n15645 & ~n16170;
  assign n16323 = ~n15647 & ~n15646;
  assign n15648 = ~n15961 & ~n16323;
  assign n15650 = ~n15649 & ~n15648;
  assign n15652 = n15651 & n15650;
  assign P1_U3280 = ~n15653 | ~n15652;
  assign n15655 = ~n15992 | ~n9563;
  assign n15654 = ~n15961 | ~P1_REG2_REG_12__SCAN_IN;
  assign n15658 = ~n15655 | ~n15654;
  assign n15657 = ~n15917 & ~n15656;
  assign n15673 = ~n15658 & ~n15657;
  assign n16303 = ~n15697 ^ n15659;
  assign n15671 = ~n16303 | ~n15991;
  assign n16307 = n15660 ^ n15664;
  assign n15669 = ~n16307 & ~n15747;
  assign n15663 = ~n15711 | ~n15979;
  assign n15662 = ~n15661 | ~n11990;
  assign n15667 = ~n15663 | ~n15662;
  assign n15665 = n9025 ^ n15664;
  assign n15666 = ~n15665 & ~n16170;
  assign n16311 = ~n15667 & ~n15666;
  assign n15668 = ~n15961 & ~n16311;
  assign n15670 = ~n15669 & ~n15668;
  assign n15672 = n15671 & n15670;
  assign P1_U3281 = ~n15673 | ~n15672;
  assign n16296 = ~n15674 ^ n15680;
  assign n15676 = ~n16296;
  assign n15690 = ~n15676 | ~n15675;
  assign n15679 = ~n15678 | ~n15677;
  assign n15681 = n15680 ^ n15679;
  assign n15687 = ~n15681 | ~n15977;
  assign n15683 = ~n15979 | ~n15734;
  assign n15682 = ~n11990 | ~n9305;
  assign n15685 = ~n15683 | ~n15682;
  assign n15684 = ~n16296 & ~n15983;
  assign n15686 = ~n15685 & ~n15684;
  assign n16298 = ~n15687 | ~n15686;
  assign n15688 = ~n16292 & ~n15902;
  assign n15689 = ~n16298 & ~n15688;
  assign n15693 = ~n15690 | ~n15689;
  assign n15692 = ~n15917 & ~n15691;
  assign n15694 = ~n15693 & ~n15692;
  assign n15700 = ~n15961 & ~n15694;
  assign n15696 = n15695 | n16292;
  assign n16290 = ~n15697 | ~n15696;
  assign n15698 = ~n15991;
  assign n15699 = ~n16290 & ~n15698;
  assign n15702 = ~n15700 & ~n15699;
  assign n15701 = ~P1_REG2_REG_11__SCAN_IN | ~n15961;
  assign P1_U3282 = ~n15702 | ~n15701;
  assign n15704 = ~n15992 | ~n16279;
  assign n15703 = ~n15961 | ~P1_REG2_REG_10__SCAN_IN;
  assign n15707 = ~n15704 | ~n15703;
  assign n15706 = ~n15917 & ~n15705;
  assign n15721 = ~n15707 & ~n15706;
  assign n16278 = ~n15708 ^ n16279;
  assign n15719 = ~n16278 | ~n15991;
  assign n16282 = n9026 ^ n15709;
  assign n15717 = ~n16282 & ~n15747;
  assign n15715 = ~n15710 & ~n16170;
  assign n15713 = ~n15711 | ~n11990;
  assign n15712 = ~n15771 | ~n15979;
  assign n15714 = ~n15713 | ~n15712;
  assign n16286 = ~n15715 & ~n15714;
  assign n15716 = ~n15961 & ~n16286;
  assign n15718 = ~n15717 & ~n15716;
  assign n15720 = n15719 & n15718;
  assign P1_U3283 = ~n15721 | ~n15720;
  assign n15724 = ~n15818 | ~n15722;
  assign n15791 = n15724 & n15723;
  assign n15764 = ~n15791 | ~n15795;
  assign n15726 = ~n15764 | ~n15725;
  assign n15727 = ~n15726 | ~n15760;
  assign n15728 = n15727 ^ n15746;
  assign n15731 = ~n15728 | ~n15977;
  assign n15730 = ~n15729 | ~n15979;
  assign n16270 = ~n15731 | ~n15730;
  assign n15733 = ~n15732 ^ n16271;
  assign n15736 = ~n15733 | ~n16327;
  assign n15735 = ~n15734 | ~n11990;
  assign n16273 = ~n15736 | ~n15735;
  assign n15739 = ~n16273 | ~n16044;
  assign n15738 = ~n15737 | ~n15927;
  assign n15740 = ~n15739 | ~n15738;
  assign n15743 = n16270 | n15740;
  assign n15742 = ~n15917 & ~n15741;
  assign n15744 = ~n15743 & ~n15742;
  assign n15749 = ~n15961 & ~n15744;
  assign n16268 = n15745 ^ n15746;
  assign n15748 = ~n16268 & ~n15747;
  assign n15751 = ~n15749 & ~n15748;
  assign n15750 = ~P1_REG2_REG_9__SCAN_IN | ~n15961;
  assign P1_U3284 = ~n15751 | ~n15750;
  assign n15753 = ~n15992 | ~n16258;
  assign n15752 = ~n15961 | ~P1_REG2_REG_8__SCAN_IN;
  assign n15756 = ~n15753 | ~n15752;
  assign n15755 = ~n15917 & ~n15754;
  assign n15779 = ~n15756 & ~n15755;
  assign n16257 = ~n15788 ^ n15757;
  assign n15762 = ~n15991 | ~n16257;
  assign n15766 = ~n15760 | ~n15759;
  assign n16261 = ~n15758 ^ n15766;
  assign n15768 = ~n16261;
  assign n15971 = ~n15954;
  assign n15761 = ~n15768 | ~n15971;
  assign n15777 = ~n15762 | ~n15761;
  assign n15765 = ~n15764 | ~n15763;
  assign n15767 = n15766 ^ n15765;
  assign n15770 = ~n15767 | ~n15977;
  assign n15769 = ~n15768 | ~n15942;
  assign n15775 = ~n15770 | ~n15769;
  assign n15773 = ~n15823 | ~n15979;
  assign n15772 = ~n15771 | ~n11990;
  assign n15774 = ~n15773 | ~n15772;
  assign n16265 = ~n15775 & ~n15774;
  assign n15776 = ~n15961 & ~n16265;
  assign n15778 = ~n15777 & ~n15776;
  assign P1_U3285 = ~n15779 | ~n15778;
  assign n15784 = ~n16004 & ~n15780;
  assign n15782 = ~n15781;
  assign n15783 = ~n15917 & ~n15782;
  assign n15812 = ~n15784 & ~n15783;
  assign n15787 = ~n15786 & ~n15785;
  assign n15789 = ~n15787 & ~n16289;
  assign n16252 = n15789 & n15788;
  assign n15806 = n16252 & n16044;
  assign n15800 = ~n15790 & ~n15933;
  assign n15792 = ~n15791 ^ n15795;
  assign n15798 = ~n15792 | ~n15977;
  assign n15796 = ~n15794 | ~n15795;
  assign n16248 = ~n9785 | ~n15796;
  assign n15797 = ~n15942 | ~n16248;
  assign n15799 = ~n15798 | ~n15797;
  assign n15803 = n15800 | n15799;
  assign n15802 = ~n15801 & ~n15875;
  assign n16254 = ~n15803 & ~n15802;
  assign n15804 = ~n11963 | ~n15927;
  assign n15805 = ~n16254 | ~n15804;
  assign n15807 = ~n15806 & ~n15805;
  assign n15810 = ~n15961 & ~n15807;
  assign n15808 = ~n16248;
  assign n15809 = ~n15808 & ~n15954;
  assign n15811 = ~n15810 & ~n15809;
  assign P1_U3286 = ~n15812 | ~n15811;
  assign n15849 = ~n15813 & ~n15850;
  assign n15815 = ~n15849 & ~n15814;
  assign n15833 = n15819 ^ n15815;
  assign n15817 = ~n15833 | ~n15942;
  assign n15816 = ~n15876 | ~n15979;
  assign n15822 = ~n15817 | ~n15816;
  assign n15820 = n15818 ^ n15819;
  assign n15821 = ~n15820 & ~n16170;
  assign n16245 = ~n15822 & ~n15821;
  assign n16237 = ~n15823 | ~n11990;
  assign n15824 = ~n16245 | ~n16237;
  assign n15832 = ~n15824 | ~n16004;
  assign n15828 = ~n16004 & ~n15825;
  assign n15827 = ~n15917 & ~n15826;
  assign n15830 = ~n15828 & ~n15827;
  assign n15829 = ~n15992 | ~n9550;
  assign n15831 = n15830 & n15829;
  assign n15835 = ~n15832 | ~n15831;
  assign n16241 = ~n15833;
  assign n15834 = ~n16241 & ~n15954;
  assign n15837 = ~n15835 & ~n15834;
  assign n16238 = ~n9032 ^ n9550;
  assign n15836 = ~n15991 | ~n16238;
  assign P1_U3287 = ~n15837 | ~n15836;
  assign n15838 = ~n15884 | ~n16227;
  assign n15839 = ~n15838 | ~n16327;
  assign n16231 = ~n9032 & ~n15839;
  assign n15841 = ~n16231 | ~n16044;
  assign n15840 = ~n16227 | ~n15927;
  assign n15856 = ~n15841 | ~n15840;
  assign n15843 = ~n15842 ^ n9021;
  assign n15848 = ~n15843 & ~n16170;
  assign n15846 = ~n11903 | ~n15979;
  assign n15845 = ~n15844 | ~n11990;
  assign n15847 = ~n15846 | ~n15845;
  assign n16233 = ~n15848 & ~n15847;
  assign n15852 = ~n15849;
  assign n15851 = ~n15813 | ~n15850;
  assign n16226 = ~n15852 | ~n15851;
  assign n15854 = ~n16226 | ~n15853;
  assign n15855 = ~n16233 | ~n15854;
  assign n15857 = ~n15856 & ~n15855;
  assign n15861 = n15857 | n15961;
  assign n15859 = ~n15858;
  assign n15860 = n15917 | n15859;
  assign n15863 = n15861 & n15860;
  assign n15862 = ~P1_REG2_REG_5__SCAN_IN | ~n15961;
  assign P1_U3288 = ~n15863 | ~n15862;
  assign n15864 = ~P1_REG2_REG_4__SCAN_IN;
  assign n15868 = ~n16004 & ~n15864;
  assign n15866 = ~n15865;
  assign n15867 = ~n15917 & ~n15866;
  assign n15870 = ~n15868 & ~n15867;
  assign n15869 = ~n15992 | ~n16216;
  assign n15900 = n15870 & n15869;
  assign n15873 = ~n15872 | ~n15871;
  assign n15874 = n15893 ^ n15873;
  assign n15881 = ~n15874 | ~n15977;
  assign n15879 = ~n15934 & ~n15875;
  assign n15877 = ~n15876;
  assign n15878 = ~n15877 & ~n15933;
  assign n15880 = ~n15879 & ~n15878;
  assign n16220 = ~n15881 | ~n15880;
  assign n15883 = ~n15924 & ~n9323;
  assign n15886 = ~n15883 & ~n15882;
  assign n15885 = ~n15884 | ~n16327;
  assign n16221 = n15886 | n15885;
  assign n15887 = ~n16221 & ~n10531;
  assign n15888 = ~n16220 & ~n15887;
  assign n15898 = ~n15961 & ~n15888;
  assign n15891 = n15890 & n15889;
  assign n15895 = n15892 & n15891;
  assign n15894 = ~n15893;
  assign n16215 = ~n15895 ^ n15894;
  assign n15897 = n15896 & n16215;
  assign n15899 = ~n15898 & ~n15897;
  assign P1_U3289 = ~n15900 | ~n15899;
  assign n16204 = ~n15901 & ~n15933;
  assign n15903 = ~n16202 & ~n15902;
  assign n15915 = ~n16204 & ~n15903;
  assign n15938 = ~n15935 | ~n15904;
  assign n15905 = ~n15938 | ~n13390;
  assign n15906 = ~n15905 ^ n13286;
  assign n15914 = ~n15906 & ~n16170;
  assign n15941 = n15907 & n13285;
  assign n15909 = ~n15941 & ~n15908;
  assign n16208 = ~n15909 ^ n13286;
  assign n15910 = ~n16208;
  assign n15912 = ~n15910 | ~n15942;
  assign n15911 = ~n11910 | ~n15979;
  assign n15913 = ~n15912 | ~n15911;
  assign n16212 = ~n15914 & ~n15913;
  assign n15916 = ~n15915 | ~n16212;
  assign n15921 = ~n15916 | ~n16004;
  assign n15919 = P1_REG2_REG_3__SCAN_IN & n15961;
  assign n15918 = ~P1_REG3_REG_3__SCAN_IN & ~n15917;
  assign n15920 = ~n15919 & ~n15918;
  assign n15923 = ~n15921 | ~n15920;
  assign n15922 = ~n15954 & ~n16208;
  assign n15926 = ~n15923 & ~n15922;
  assign n16205 = ~n15924 ^ n16202;
  assign n15925 = ~n15991 | ~n16205;
  assign P1_U3290 = ~n15926 | ~n15925;
  assign n15929 = ~n16000 | ~P1_REG3_REG_2__SCAN_IN;
  assign n15928 = ~n16193 | ~n15927;
  assign n15951 = ~n15929 | ~n15928;
  assign n15932 = ~n15931 ^ n15930;
  assign n16197 = ~n15932 & ~n16289;
  assign n15949 = ~n16197 | ~n16044;
  assign n15946 = ~n15934 & ~n15933;
  assign n15936 = ~n15935;
  assign n15937 = ~n15936 | ~n13285;
  assign n15939 = ~n15938 | ~n15937;
  assign n15944 = ~n15977 | ~n15939;
  assign n15940 = ~n15907 & ~n13285;
  assign n15953 = ~n15941 & ~n15940;
  assign n16192 = ~n15953;
  assign n15943 = ~n15942 | ~n16192;
  assign n15945 = ~n15944 | ~n15943;
  assign n15948 = ~n15946 & ~n15945;
  assign n15947 = ~n9310 | ~n15979;
  assign n16199 = n15948 & n15947;
  assign n15950 = ~n15949 | ~n16199;
  assign n15952 = ~n15951 & ~n15950;
  assign n15956 = ~n15961 & ~n15952;
  assign n15955 = ~n15954 & ~n15953;
  assign n15958 = ~n15956 & ~n15955;
  assign n15957 = ~P1_REG2_REG_2__SCAN_IN | ~n15961;
  assign P1_U3291 = ~n15958 | ~n15957;
  assign n15960 = ~n15992 | ~n16182;
  assign n16181 = ~n16182 ^ n15993;
  assign n15959 = ~n15991 | ~n16181;
  assign n15965 = ~n15960 | ~n15959;
  assign n15963 = ~n15961 | ~P1_REG2_REG_1__SCAN_IN;
  assign n15962 = ~P1_REG3_REG_1__SCAN_IN | ~n16000;
  assign n15964 = ~n15963 | ~n15962;
  assign n15973 = ~n15965 & ~n15964;
  assign n15967 = ~n15966;
  assign n15970 = ~n15968 | ~n15967;
  assign n16187 = ~n15970 | ~n15969;
  assign n15972 = ~n15971 | ~n16187;
  assign n15990 = n15973 & n15972;
  assign n15976 = ~n13283 | ~n15974;
  assign n15978 = ~n15976 | ~n15975;
  assign n15988 = ~n15978 | ~n15977;
  assign n15982 = ~n15980 | ~n15979;
  assign n15981 = ~n11910 | ~n11990;
  assign n15986 = ~n15982 | ~n15981;
  assign n15984 = ~n16187;
  assign n15985 = ~n15984 & ~n15983;
  assign n15987 = ~n15986 & ~n15985;
  assign n16186 = ~n15988 | ~n15987;
  assign n15989 = ~n16004 | ~n16186;
  assign P1_U3292 = ~n15990 | ~n15989;
  assign n15994 = ~n15992 & ~n15991;
  assign n15997 = ~n15994 & ~n15993;
  assign n15996 = ~n16004 & ~n15995;
  assign n16006 = ~n15997 & ~n15996;
  assign n15999 = ~n16171 | ~n15998;
  assign n16176 = ~n9310 | ~n11990;
  assign n16002 = n15999 & n16176;
  assign n16001 = ~n16000 | ~P1_REG3_REG_0__SCAN_IN;
  assign n16003 = ~n16002 | ~n16001;
  assign n16005 = ~n16004 | ~n16003;
  assign P1_U3293 = ~n16006 | ~n16005;
  assign P1_U3294 = P1_D_REG_31__SCAN_IN & n16165;
  assign P1_U3295 = P1_D_REG_30__SCAN_IN & n16165;
  assign P1_U3296 = P1_D_REG_29__SCAN_IN & n16165;
  assign P1_U3297 = P1_D_REG_28__SCAN_IN & n16165;
  assign P1_U3298 = P1_D_REG_27__SCAN_IN & n16165;
  assign P1_U3299 = P1_D_REG_26__SCAN_IN & n16165;
  assign P1_U3300 = P1_D_REG_25__SCAN_IN & n16165;
  assign P1_U3301 = P1_D_REG_24__SCAN_IN & n16165;
  assign P1_U3302 = P1_D_REG_23__SCAN_IN & n16165;
  assign P1_U3303 = P1_D_REG_22__SCAN_IN & n16165;
  assign P1_U3304 = P1_D_REG_21__SCAN_IN & n16165;
  assign P1_U3305 = P1_D_REG_20__SCAN_IN & n16165;
  assign P1_U3306 = P1_D_REG_19__SCAN_IN & n16165;
  assign P1_U3307 = P1_D_REG_18__SCAN_IN & n16165;
  assign P1_U3308 = P1_D_REG_17__SCAN_IN & n16165;
  assign P1_U3309 = P1_D_REG_16__SCAN_IN & n16165;
  assign P1_U3310 = P1_D_REG_15__SCAN_IN & n16165;
  assign P1_U3311 = P1_D_REG_14__SCAN_IN & n16165;
  assign P1_U3312 = P1_D_REG_13__SCAN_IN & n16165;
  assign P1_U3313 = P1_D_REG_12__SCAN_IN & n16165;
  assign P1_U3314 = P1_D_REG_11__SCAN_IN & n16165;
  assign P1_U3315 = P1_D_REG_10__SCAN_IN & n16165;
  assign P1_U3316 = P1_D_REG_9__SCAN_IN & n16165;
  assign P1_U3317 = P1_D_REG_8__SCAN_IN & n16165;
  assign P1_U3318 = P1_D_REG_7__SCAN_IN & n16165;
  assign P1_U3319 = P1_D_REG_6__SCAN_IN & n16165;
  assign P1_U3320 = P1_D_REG_5__SCAN_IN & n16165;
  assign P1_U3321 = P1_D_REG_4__SCAN_IN & n16165;
  assign P1_U3322 = P1_D_REG_3__SCAN_IN & n16165;
  assign P1_U3323 = P1_D_REG_2__SCAN_IN & n16165;
  assign n16012 = ~n17213 & ~n16154;
  assign n16010 = ~n16009;
  assign n16011 = ~n16010 & ~P1_U3086;
  assign n16014 = ~n16012 & ~n16011;
  assign n16013 = ~n16159 | ~P2_DATAO_REG_25__SCAN_IN;
  assign P1_U3330 = ~n16014 | ~n16013;
  assign n16018 = ~n17219 & ~n16154;
  assign n16016 = ~n16015;
  assign n16017 = ~n16016 & ~P1_U3086;
  assign n16020 = ~n16018 & ~n16017;
  assign n16019 = ~n16159 | ~P2_DATAO_REG_24__SCAN_IN;
  assign P1_U3331 = ~n16020 | ~n16019;
  assign n17224 = ~n16021;
  assign n16025 = ~n17224 & ~n16154;
  assign n16024 = ~n16023 & ~n16022;
  assign n16027 = ~n16025 & ~n16024;
  assign P1_U3332 = ~n16027 | ~n16026;
  assign n17231 = ~n16028;
  assign n16031 = ~n17231 & ~n16154;
  assign n16030 = ~n16029 & ~P1_U3086;
  assign n16033 = ~n16031 & ~n16030;
  assign n16032 = ~n16159 | ~P2_DATAO_REG_22__SCAN_IN;
  assign P1_U3333 = ~n16033 | ~n16032;
  assign n16036 = ~n17237 & ~n16154;
  assign n16035 = ~n16034 & ~P1_U3086;
  assign n16038 = ~n16036 & ~n16035;
  assign n16037 = ~n16159 | ~P2_DATAO_REG_21__SCAN_IN;
  assign P1_U3334 = ~n16038 | ~n16037;
  assign n16041 = ~n12213 & ~n16154;
  assign n16040 = ~n16039;
  assign n16043 = ~n16041 & ~n16040;
  assign n16042 = ~n16159 | ~P2_DATAO_REG_20__SCAN_IN;
  assign P1_U3335 = ~n16043 | ~n16042;
  assign n16046 = ~n17248 & ~n16154;
  assign n16045 = ~n16044 & ~P1_U3086;
  assign n16048 = ~n16046 & ~n16045;
  assign n16047 = ~n16159 | ~P2_DATAO_REG_19__SCAN_IN;
  assign P1_U3336 = ~n16048 | ~n16047;
  assign n16051 = ~n17253 & ~n16154;
  assign n16050 = ~n16049 & ~P1_U3086;
  assign n16053 = ~n16051 & ~n16050;
  assign n16052 = ~n16159 | ~P2_DATAO_REG_18__SCAN_IN;
  assign P1_U3337 = ~n16053 | ~n16052;
  assign n16055 = ~n16054;
  assign n16059 = ~n16055 & ~n16154;
  assign n16057 = ~n16056;
  assign n16058 = ~n16057 & ~P1_U3086;
  assign n16061 = ~n16059 & ~n16058;
  assign n16060 = ~n16159 | ~P2_DATAO_REG_17__SCAN_IN;
  assign P1_U3338 = ~n16061 | ~n16060;
  assign n16065 = ~n17259 & ~n16154;
  assign n16063 = ~n16062;
  assign n16064 = ~n16063 & ~P1_U3086;
  assign n16067 = ~n16065 & ~n16064;
  assign n16066 = ~n16159 | ~P2_DATAO_REG_16__SCAN_IN;
  assign P1_U3339 = ~n16067 | ~n16066;
  assign n17265 = ~n16068;
  assign n16072 = ~n17265 & ~n16154;
  assign n16070 = ~n16069;
  assign n16071 = ~n16070 & ~P1_U3086;
  assign n16074 = ~n16072 & ~n16071;
  assign n16073 = ~n16159 | ~P2_DATAO_REG_15__SCAN_IN;
  assign P1_U3340 = ~n16074 | ~n16073;
  assign n16078 = ~n12157 & ~n16154;
  assign n16076 = ~n16075;
  assign n16077 = ~n16076 & ~P1_U3086;
  assign n16080 = ~n16078 & ~n16077;
  assign n16079 = ~n16159 | ~P2_DATAO_REG_14__SCAN_IN;
  assign P1_U3341 = ~n16080 | ~n16079;
  assign n16084 = ~n17276 & ~n16154;
  assign n16082 = ~n16081;
  assign n16083 = ~n16082 & ~P1_U3086;
  assign n16086 = ~n16084 & ~n16083;
  assign n16085 = ~n16159 | ~P2_DATAO_REG_13__SCAN_IN;
  assign P1_U3342 = ~n16086 | ~n16085;
  assign n17282 = ~n16087;
  assign n16091 = ~n17282 & ~n16154;
  assign n16089 = ~n16088;
  assign n16090 = ~n16089 & ~P1_U3086;
  assign n16093 = ~n16091 & ~n16090;
  assign n16092 = ~n16159 | ~P2_DATAO_REG_12__SCAN_IN;
  assign P1_U3343 = ~n16093 | ~n16092;
  assign n17288 = ~n16094;
  assign n16098 = ~n17288 & ~n16154;
  assign n16096 = ~n16095;
  assign n16097 = ~n16096 & ~P1_U3086;
  assign n16100 = ~n16098 & ~n16097;
  assign n16099 = ~n16159 | ~P2_DATAO_REG_11__SCAN_IN;
  assign P1_U3344 = ~n16100 | ~n16099;
  assign n16104 = ~n17294 & ~n16154;
  assign n16102 = ~n16101;
  assign n16103 = ~n16102 & ~P1_U3086;
  assign n16106 = ~n16104 & ~n16103;
  assign n16105 = ~n16159 | ~P2_DATAO_REG_10__SCAN_IN;
  assign P1_U3345 = ~n16106 | ~n16105;
  assign n16109 = ~n17300 & ~n16154;
  assign n16108 = ~n16107 & ~P1_U3086;
  assign n16111 = ~n16109 & ~n16108;
  assign n16110 = ~n16159 | ~P2_DATAO_REG_9__SCAN_IN;
  assign P1_U3346 = ~n16111 | ~n16110;
  assign n16114 = ~n17306 & ~n16154;
  assign n16113 = ~n16112 & ~P1_U3086;
  assign n16116 = ~n16114 & ~n16113;
  assign n16115 = ~n16159 | ~P2_DATAO_REG_8__SCAN_IN;
  assign P1_U3347 = ~n16116 | ~n16115;
  assign n16119 = ~n17312 & ~n16154;
  assign n16118 = ~n16117 & ~P1_U3086;
  assign n16121 = ~n16119 & ~n16118;
  assign n16120 = ~n16159 | ~P2_DATAO_REG_7__SCAN_IN;
  assign P1_U3348 = ~n16121 | ~n16120;
  assign n16124 = ~n17318 & ~n16154;
  assign n16123 = ~n16122 & ~P1_U3086;
  assign n16126 = ~n16124 & ~n16123;
  assign n16125 = ~n16159 | ~P2_DATAO_REG_6__SCAN_IN;
  assign P1_U3349 = ~n16126 | ~n16125;
  assign n17324 = ~n16127;
  assign n16131 = ~n17324 & ~n16154;
  assign n16129 = ~n16128;
  assign n16130 = ~n16129 & ~P1_U3086;
  assign n16133 = ~n16131 & ~n16130;
  assign n16132 = ~n16159 | ~P2_DATAO_REG_5__SCAN_IN;
  assign P1_U3350 = ~n16133 | ~n16132;
  assign n16138 = ~n16135 | ~n16134;
  assign n16137 = ~n16136 | ~P1_STATE_REG_SCAN_IN;
  assign n16140 = n16138 & n16137;
  assign n16139 = ~n16159 | ~P2_DATAO_REG_4__SCAN_IN;
  assign P1_U3351 = ~n16140 | ~n16139;
  assign n16145 = ~n12066 & ~n16154;
  assign n16143 = ~n16142;
  assign n16144 = ~n16143 & ~P1_U3086;
  assign n16147 = ~n16145 & ~n16144;
  assign n16146 = ~n16159 | ~P2_DATAO_REG_3__SCAN_IN;
  assign P1_U3352 = ~n16147 | ~n16146;
  assign n16151 = ~n12056 & ~n16154;
  assign n16149 = ~n16148;
  assign n16150 = ~n16149 & ~P1_U3086;
  assign n16153 = ~n16151 & ~n16150;
  assign n16152 = ~n16159 | ~P2_DATAO_REG_2__SCAN_IN;
  assign P1_U3353 = ~n16153 | ~n16152;
  assign n16158 = ~n17342 & ~n16154;
  assign n16156 = ~n16155;
  assign n16157 = ~n16156 & ~P1_U3086;
  assign n16161 = ~n16158 & ~n16157;
  assign n16160 = ~n16159 | ~P2_DATAO_REG_1__SCAN_IN;
  assign P1_U3354 = ~n16161 | ~n16160;
  assign n16164 = ~P1_D_REG_0__SCAN_IN | ~n16165;
  assign n16167 = ~n16165;
  assign n16163 = ~n16167 | ~n16162;
  assign P1_U3439 = ~n16164 | ~n16163;
  assign n16169 = ~P1_D_REG_1__SCAN_IN | ~n16165;
  assign n16168 = ~n16167 | ~n16166;
  assign P1_U3440 = ~n16169 | ~n16168;
  assign n16180 = ~P1_REG0_REG_0__SCAN_IN | ~n16326;
  assign n16172 = ~n16318 | ~n16170;
  assign n16178 = ~n16172 | ~n16171;
  assign n16175 = ~n16174 | ~n16173;
  assign n16177 = n16176 & n16175;
  assign n16341 = ~n16178 | ~n16177;
  assign n16179 = ~n16338 | ~n16341;
  assign P1_U3453 = ~n16180 | ~n16179;
  assign n16191 = ~P1_REG0_REG_1__SCAN_IN | ~n16326;
  assign n16184 = ~n16181 | ~n16327;
  assign n16183 = ~n16329 | ~n16182;
  assign n16185 = ~n16184 | ~n16183;
  assign n16189 = ~n16186 & ~n16185;
  assign n16334 = ~n16295;
  assign n16188 = ~n16187 | ~n16334;
  assign n16344 = ~n16189 | ~n16188;
  assign n16190 = ~n16338 | ~n16344;
  assign P1_U3456 = ~n16191 | ~n16190;
  assign n16201 = ~P1_REG0_REG_2__SCAN_IN | ~n16326;
  assign n16195 = ~n16192 | ~n16334;
  assign n16194 = ~n16193 | ~n16329;
  assign n16196 = ~n16195 | ~n16194;
  assign n16198 = ~n16197 & ~n16196;
  assign n16347 = ~n16199 | ~n16198;
  assign n16200 = ~n16338 | ~n16347;
  assign P1_U3459 = ~n16201 | ~n16200;
  assign n16214 = ~P1_REG0_REG_3__SCAN_IN | ~n16326;
  assign n16203 = ~n16291 & ~n16202;
  assign n16207 = ~n16204 & ~n16203;
  assign n16206 = ~n16205 | ~n16327;
  assign n16210 = ~n16207 | ~n16206;
  assign n16209 = ~n16208 & ~n16295;
  assign n16211 = ~n16210 & ~n16209;
  assign n16350 = ~n16212 | ~n16211;
  assign n16213 = ~n16338 | ~n16350;
  assign P1_U3462 = ~n16214 | ~n16213;
  assign n16224 = ~P1_REG0_REG_4__SCAN_IN | ~n16326;
  assign n16218 = ~n16215 | ~n16225;
  assign n16217 = ~n16329 | ~n16216;
  assign n16219 = ~n16218 | ~n16217;
  assign n16222 = ~n16220 & ~n16219;
  assign n16353 = ~n16222 | ~n16221;
  assign n16223 = ~n16338 | ~n16353;
  assign P1_U3465 = ~n16224 | ~n16223;
  assign n16235 = ~P1_REG0_REG_5__SCAN_IN | ~n16326;
  assign n16229 = ~n16226 | ~n16225;
  assign n16228 = ~n16227 | ~n16329;
  assign n16230 = ~n16229 | ~n16228;
  assign n16232 = ~n16231 & ~n16230;
  assign n16356 = ~n16233 | ~n16232;
  assign n16234 = ~n16338 | ~n16356;
  assign P1_U3468 = ~n16235 | ~n16234;
  assign n16247 = ~P1_REG0_REG_6__SCAN_IN | ~n16326;
  assign n16236 = ~n9550 | ~n16329;
  assign n16240 = n16237 & n16236;
  assign n16239 = ~n16238 | ~n16327;
  assign n16243 = ~n16240 | ~n16239;
  assign n16242 = ~n16241 & ~n16295;
  assign n16244 = ~n16243 & ~n16242;
  assign n16359 = ~n16245 | ~n16244;
  assign n16246 = ~n16338 | ~n16359;
  assign P1_U3471 = ~n16247 | ~n16246;
  assign n16256 = ~P1_REG0_REG_7__SCAN_IN | ~n16326;
  assign n16250 = ~n16248 | ~n16334;
  assign n16249 = ~n11963 | ~n16329;
  assign n16251 = ~n16250 | ~n16249;
  assign n16253 = ~n16252 & ~n16251;
  assign n16362 = ~n16254 | ~n16253;
  assign n16255 = ~n16338 | ~n16362;
  assign P1_U3474 = ~n16256 | ~n16255;
  assign n16267 = ~P1_REG0_REG_8__SCAN_IN | ~n16326;
  assign n16260 = ~n16257 | ~n16327;
  assign n16259 = ~n16258 | ~n16329;
  assign n16263 = ~n16260 | ~n16259;
  assign n16262 = ~n16261 & ~n16295;
  assign n16264 = ~n16263 & ~n16262;
  assign n16365 = ~n16265 | ~n16264;
  assign n16266 = ~n16338 | ~n16365;
  assign P1_U3477 = ~n16267 | ~n16266;
  assign n16277 = ~P1_REG0_REG_9__SCAN_IN | ~n16326;
  assign n16269 = ~n16268 & ~n16318;
  assign n16275 = ~n16270 & ~n16269;
  assign n16272 = ~n16271 & ~n16291;
  assign n16274 = ~n16273 & ~n16272;
  assign n16368 = ~n16275 | ~n16274;
  assign n16276 = ~n16338 | ~n16368;
  assign P1_U3480 = ~n16277 | ~n16276;
  assign n16288 = ~P1_REG0_REG_10__SCAN_IN | ~n16326;
  assign n16281 = ~n16278 | ~n16327;
  assign n16280 = ~n16279 | ~n16329;
  assign n16284 = ~n16281 | ~n16280;
  assign n16283 = ~n16282 & ~n16318;
  assign n16285 = ~n16284 & ~n16283;
  assign n16371 = ~n16286 | ~n16285;
  assign n16287 = ~n16338 | ~n16371;
  assign P1_U3483 = ~n16288 | ~n16287;
  assign n16302 = ~P1_REG0_REG_11__SCAN_IN | ~n16326;
  assign n16294 = ~n16290 & ~n16289;
  assign n16293 = ~n16292 & ~n16291;
  assign n16300 = ~n16294 & ~n16293;
  assign n16297 = ~n16296 & ~n16295;
  assign n16299 = ~n16298 & ~n16297;
  assign n16374 = ~n16300 | ~n16299;
  assign n16301 = ~n16338 | ~n16374;
  assign P1_U3486 = ~n16302 | ~n16301;
  assign n16313 = ~P1_REG0_REG_12__SCAN_IN | ~n16326;
  assign n16306 = ~n16303 | ~n16327;
  assign n16305 = ~n9563 | ~n16329;
  assign n16309 = ~n16306 | ~n16305;
  assign n16308 = ~n16307 & ~n16318;
  assign n16310 = ~n16309 & ~n16308;
  assign n16377 = ~n16311 | ~n16310;
  assign n16312 = ~n16338 | ~n16377;
  assign P1_U3489 = ~n16313 | ~n16312;
  assign n16325 = ~P1_REG0_REG_13__SCAN_IN | ~n16326;
  assign n16317 = ~n16314 | ~n16327;
  assign n16316 = ~n16315 | ~n16329;
  assign n16321 = ~n16317 | ~n16316;
  assign n16320 = ~n16319 & ~n16318;
  assign n16322 = ~n16321 & ~n16320;
  assign n16380 = ~n16323 | ~n16322;
  assign n16324 = ~n16338 | ~n16380;
  assign P1_U3492 = ~n16325 | ~n16324;
  assign n16340 = ~P1_REG0_REG_14__SCAN_IN | ~n16326;
  assign n16331 = ~n16328 | ~n16327;
  assign n16330 = ~n9555 | ~n16329;
  assign n16332 = ~n16331 | ~n16330;
  assign n16337 = ~n16333 & ~n16332;
  assign n16336 = ~n16335 | ~n16334;
  assign n16384 = ~n16337 | ~n16336;
  assign n16339 = ~n16338 | ~n16384;
  assign P1_U3495 = ~n16340 | ~n16339;
  assign n16343 = ~P1_REG1_REG_0__SCAN_IN | ~n16383;
  assign n16342 = ~n16385 | ~n16341;
  assign P1_U3522 = ~n16343 | ~n16342;
  assign n16346 = ~P1_REG1_REG_1__SCAN_IN | ~n16383;
  assign n16345 = ~n16385 | ~n16344;
  assign P1_U3523 = ~n16346 | ~n16345;
  assign n16349 = ~P1_REG1_REG_2__SCAN_IN | ~n16383;
  assign n16348 = ~n16385 | ~n16347;
  assign P1_U3524 = ~n16349 | ~n16348;
  assign n16352 = ~P1_REG1_REG_3__SCAN_IN | ~n16383;
  assign n16351 = ~n16385 | ~n16350;
  assign P1_U3525 = ~n16352 | ~n16351;
  assign n16355 = ~P1_REG1_REG_4__SCAN_IN | ~n16383;
  assign n16354 = ~n16385 | ~n16353;
  assign P1_U3526 = ~n16355 | ~n16354;
  assign n16358 = ~P1_REG1_REG_5__SCAN_IN | ~n16383;
  assign n16357 = ~n16385 | ~n16356;
  assign P1_U3527 = ~n16358 | ~n16357;
  assign n16361 = ~P1_REG1_REG_6__SCAN_IN | ~n16383;
  assign n16360 = ~n16385 | ~n16359;
  assign P1_U3528 = ~n16361 | ~n16360;
  assign n16364 = ~P1_REG1_REG_7__SCAN_IN | ~n16383;
  assign n16363 = ~n16385 | ~n16362;
  assign P1_U3529 = ~n16364 | ~n16363;
  assign n16367 = ~P1_REG1_REG_8__SCAN_IN | ~n16383;
  assign n16366 = ~n16385 | ~n16365;
  assign P1_U3530 = ~n16367 | ~n16366;
  assign n16370 = ~P1_REG1_REG_9__SCAN_IN | ~n16383;
  assign n16369 = ~n16385 | ~n16368;
  assign P1_U3531 = ~n16370 | ~n16369;
  assign n16373 = ~P1_REG1_REG_10__SCAN_IN | ~n16383;
  assign n16372 = ~n16385 | ~n16371;
  assign P1_U3532 = ~n16373 | ~n16372;
  assign n16376 = ~P1_REG1_REG_11__SCAN_IN | ~n16383;
  assign n16375 = ~n16385 | ~n16374;
  assign P1_U3533 = ~n16376 | ~n16375;
  assign n16379 = ~P1_REG1_REG_12__SCAN_IN | ~n16383;
  assign n16378 = ~n16385 | ~n16377;
  assign P1_U3534 = ~n16379 | ~n16378;
  assign n16382 = ~P1_REG1_REG_13__SCAN_IN | ~n16383;
  assign n16381 = ~n16385 | ~n16380;
  assign P1_U3535 = ~n16382 | ~n16381;
  assign n16387 = ~P1_REG1_REG_14__SCAN_IN | ~n16383;
  assign n16386 = ~n16385 | ~n16384;
  assign P1_U3536 = ~n16387 | ~n16386;
  assign n16390 = ~P1_DATAO_REG_18__SCAN_IN | ~n11337;
  assign n16389 = ~P1_U3973 | ~n16388;
  assign P1_U3572 = ~n16390 | ~n16389;
  assign n16393 = ~P1_DATAO_REG_19__SCAN_IN | ~n11337;
  assign n16392 = ~P1_U3973 | ~n16391;
  assign P1_U3573 = ~n16393 | ~n16392;
  assign n16396 = ~P1_DATAO_REG_20__SCAN_IN | ~n11337;
  assign n16395 = ~P1_U3973 | ~n16394;
  assign P1_U3574 = ~n16396 | ~n16395;
  assign n16399 = ~P1_DATAO_REG_21__SCAN_IN | ~n11337;
  assign n16398 = ~P1_U3973 | ~n16397;
  assign P1_U3575 = ~n16399 | ~n16398;
  assign n16402 = ~P1_DATAO_REG_22__SCAN_IN | ~n11337;
  assign n16401 = ~P1_U3973 | ~n16400;
  assign P1_U3576 = ~n16402 | ~n16401;
  assign n16405 = ~P1_DATAO_REG_23__SCAN_IN | ~n11337;
  assign n16404 = ~P1_U3973 | ~n16403;
  assign P1_U3577 = ~n16405 | ~n16404;
  assign n16408 = ~P1_DATAO_REG_24__SCAN_IN | ~n11337;
  assign n16407 = ~P1_U3973 | ~n16406;
  assign P1_U3578 = ~n16408 | ~n16407;
  assign n16411 = ~P1_DATAO_REG_25__SCAN_IN | ~n11337;
  assign n16410 = ~P1_U3973 | ~n16409;
  assign P1_U3579 = ~n16411 | ~n16410;
  assign n16414 = ~P1_DATAO_REG_26__SCAN_IN | ~n11337;
  assign n16413 = ~P1_U3973 | ~n16412;
  assign P1_U3580 = ~n16414 | ~n16413;
  assign n16417 = ~P1_DATAO_REG_27__SCAN_IN | ~n11337;
  assign n16416 = ~P1_U3973 | ~n16415;
  assign P1_U3581 = ~n16417 | ~n16416;
  assign n16420 = ~P1_DATAO_REG_28__SCAN_IN | ~n11337;
  assign n16419 = ~P1_U3973 | ~n16418;
  assign P1_U3582 = ~n16420 | ~n16419;
  assign n16423 = ~P1_DATAO_REG_29__SCAN_IN | ~n11337;
  assign n16422 = ~P1_U3973 | ~n16421;
  assign P1_U3583 = ~n16423 | ~n16422;
  assign n16426 = ~P1_DATAO_REG_30__SCAN_IN | ~n11337;
  assign n16425 = n11337 | n16424;
  assign P1_U3584 = ~n16426 | ~n16425;
  assign n16429 = ~P1_DATAO_REG_31__SCAN_IN | ~n11337;
  assign n16428 = ~P1_U3973 | ~n16427;
  assign P1_U3585 = ~n16429 | ~n16428;
  assign n16430 = ~n16616 | ~n17043;
  assign n16753 = ~P2_REG3_REG_7__SCAN_IN | ~P2_U3151;
  assign n16434 = ~n16430 | ~n16753;
  assign n16432 = ~n16604 | ~n17078;
  assign n16431 = ~n16605 | ~n17036;
  assign n16433 = ~n16432 | ~n16431;
  assign n16439 = ~n16434 & ~n16433;
  assign n16435 = n16477 ^ n16555;
  assign n16437 = ~n16435 & ~n16610;
  assign n16436 = ~n17046 & ~n16618;
  assign n16438 = ~n16437 & ~n16436;
  assign P2_U3153 = ~n16439 | ~n16438;
  assign n16441 = ~n16542 & ~n16507;
  assign n16440 = ~n16574 & ~n16472;
  assign n16455 = ~n16441 & ~n16440;
  assign n16443 = ~n16616 | ~n16442;
  assign n16808 = ~P2_REG3_REG_10__SCAN_IN | ~P2_U3151;
  assign n16453 = ~n16443 | ~n16808;
  assign n16447 = ~n16444;
  assign n16446 = ~n16445 ^ n16573;
  assign n16448 = ~n16447 ^ n16446;
  assign n16451 = ~n16448 | ~n16595;
  assign n16450 = ~n16577 | ~n16449;
  assign n16452 = ~n16451 | ~n16450;
  assign n16454 = ~n16453 & ~n16452;
  assign P2_U3157 = ~n16455 | ~n16454;
  assign n16457 = ~n16605 | ~n17132;
  assign n16456 = ~n16604 | ~n17168;
  assign n16465 = ~n16457 | ~n16456;
  assign n16463 = ~n16458;
  assign n16461 = ~n16459 | ~n16460;
  assign n16462 = ~n16461 | ~n16595;
  assign n16464 = ~n16463 & ~n16462;
  assign n16471 = ~n16465 & ~n16464;
  assign n16467 = ~n16616 | ~n16466;
  assign n16678 = ~P2_REG3_REG_3__SCAN_IN | ~P2_U3151;
  assign n16469 = ~n16467 | ~n16678;
  assign n16468 = ~P2_REG3_REG_3__SCAN_IN & ~n16618;
  assign n16470 = ~n16469 & ~n16468;
  assign P2_U3158 = ~n16471 | ~n16470;
  assign n16475 = ~n16542 & ~n16472;
  assign n16474 = ~n16574 & ~n16473;
  assign n16494 = ~n16475 & ~n16474;
  assign n17018 = ~n17422;
  assign n16476 = ~n16616 | ~n17018;
  assign n16770 = ~P2_REG3_REG_8__SCAN_IN | ~P2_U3151;
  assign n16492 = ~n16476 | ~n16770;
  assign n16484 = n16555 | n16477;
  assign n16481 = n16484 & n16478;
  assign n16480 = n16485 & n16479;
  assign n16482 = ~n16481 & ~n16480;
  assign n16488 = ~n16482 & ~n16610;
  assign n16486 = n16484 & n16483;
  assign n16487 = ~n16486 | ~n16485;
  assign n16490 = ~n16488 | ~n16487;
  assign n16489 = ~n16577 | ~n17019;
  assign n16491 = ~n16490 | ~n16489;
  assign n16493 = ~n16492 & ~n16491;
  assign P2_U3161 = ~n16494 | ~n16493;
  assign n16497 = ~n16496 ^ n16495;
  assign n16505 = ~n16497 | ~n16595;
  assign n16499 = ~n16604 | ~n17167;
  assign n16498 = ~n16616 | ~n17184;
  assign n16503 = ~n16499 | ~n16498;
  assign n16501 = ~P2_REG3_REG_1__SCAN_IN | ~n16601;
  assign n16500 = ~n16605 | ~n17168;
  assign n16502 = ~n16501 | ~n16500;
  assign n16504 = ~n16503 & ~n16502;
  assign P2_U3162 = ~n16505 | ~n16504;
  assign n16506 = ~n16605 | ~n17465;
  assign n16852 = ~P2_REG3_REG_12__SCAN_IN | ~P2_U3151;
  assign n16509 = ~n16506 | ~n16852;
  assign n16508 = ~n16574 & ~n16507;
  assign n16521 = ~n16509 & ~n16508;
  assign n16512 = ~n16577 | ~n16510;
  assign n16511 = ~n17463 | ~n16616;
  assign n16519 = ~n16512 | ~n16511;
  assign n16515 = ~n16514 & ~n16513;
  assign n16517 = ~n16515 & ~n16610;
  assign n16518 = n16517 & n16516;
  assign n16520 = ~n16519 & ~n16518;
  assign P2_U3164 = ~n16521 | ~n16520;
  assign n16523 = ~n16616 | ~n16522;
  assign n16720 = ~P2_REG3_REG_5__SCAN_IN | ~P2_U3151;
  assign n16527 = ~n16523 | ~n16720;
  assign n16525 = ~n16605 | ~n17078;
  assign n16524 = ~n16604 | ~n17132;
  assign n16526 = ~n16525 | ~n16524;
  assign n16536 = ~n16527 & ~n16526;
  assign n16529 = n16539 | n16538;
  assign n16530 = ~n16529 | ~n16528;
  assign n16532 = n16531 ^ n16530;
  assign n16534 = ~n16532 & ~n16610;
  assign n16533 = ~n17071 & ~n16618;
  assign n16535 = ~n16534 & ~n16533;
  assign P2_U3167 = ~n16536 | ~n16535;
  assign n16537 = ~n16616 | ~n17111;
  assign n16702 = ~P2_REG3_REG_4__SCAN_IN | ~P2_U3151;
  assign n16549 = ~n16537 | ~n16702;
  assign n16540 = ~n16539 ^ n16538;
  assign n16547 = ~n16540 | ~n16595;
  assign n16541 = ~n17102;
  assign n16545 = ~n16542 & ~n16541;
  assign n16544 = ~n16574 & ~n16543;
  assign n16546 = ~n16545 & ~n16544;
  assign n16548 = ~n16547 | ~n16546;
  assign n16551 = ~n16549 & ~n16548;
  assign n16550 = ~n17112 | ~n16577;
  assign P2_U3170 = ~n16551 | ~n16550;
  assign n16553 = ~n16604 | ~n17036;
  assign n16552 = ~n16605 | ~n16989;
  assign n16565 = ~n16553 | ~n16552;
  assign n16561 = n16555 | n16554;
  assign n16558 = n16561 & n16556;
  assign n16559 = ~n16558 & ~n16557;
  assign n16563 = ~n16559 & ~n16610;
  assign n16562 = ~n16561 | ~n16560;
  assign n16564 = n16563 & n16562;
  assign n16571 = ~n16565 & ~n16564;
  assign n16567 = ~n16616 | ~n16566;
  assign n16795 = ~P2_REG3_REG_9__SCAN_IN | ~P2_U3151;
  assign n16569 = ~n16567 | ~n16795;
  assign n16568 = ~n16983 & ~n16618;
  assign n16570 = ~n16569 & ~n16568;
  assign P2_U3171 = ~n16571 | ~n16570;
  assign n16572 = ~n16605 | ~n16974;
  assign n16834 = ~P2_REG3_REG_11__SCAN_IN | ~P2_U3151;
  assign n16576 = ~n16572 | ~n16834;
  assign n16575 = ~n16574 & ~n16573;
  assign n16589 = ~n16576 & ~n16575;
  assign n16579 = ~n16577 | ~n16958;
  assign n16578 = ~n17451 | ~n16616;
  assign n16587 = ~n16579 | ~n16578;
  assign n16585 = ~n16580;
  assign n16583 = ~n16581 | ~n16582;
  assign n16584 = ~n16583 | ~n16595;
  assign n16586 = ~n16585 & ~n16584;
  assign n16588 = ~n16587 & ~n16586;
  assign P2_U3176 = ~n16589 | ~n16588;
  assign n16592 = ~n16604 | ~n17151;
  assign n16591 = ~n16616 | ~n16590;
  assign n16600 = ~n16592 | ~n16591;
  assign n16596 = ~n16594 ^ n16593;
  assign n16598 = ~n16596 | ~n16595;
  assign n16597 = ~n16605 | ~n17150;
  assign n16599 = ~n16598 | ~n16597;
  assign n16603 = ~n16600 & ~n16599;
  assign n16602 = ~P2_REG3_REG_2__SCAN_IN | ~n16601;
  assign P2_U3177 = ~n16603 | ~n16602;
  assign n16607 = ~n16604 | ~n17102;
  assign n16606 = ~n16605 | ~n17053;
  assign n16615 = ~n16607 | ~n16606;
  assign n16611 = ~n16609 & ~n16608;
  assign n16613 = ~n16611 & ~n16610;
  assign n16614 = n16613 & n16612;
  assign n16622 = ~n16615 & ~n16614;
  assign n16617 = ~n16616 | ~n17062;
  assign n16732 = ~P2_REG3_REG_6__SCAN_IN | ~P2_U3151;
  assign n16620 = ~n16617 | ~n16732;
  assign n16619 = ~n17065 & ~n16618;
  assign n16621 = ~n16620 & ~n16619;
  assign P2_U3179 = ~n16622 | ~n16621;
  assign n16624 = ~P2_ADDR_REG_0__SCAN_IN | ~n16945;
  assign n16623 = ~P2_REG3_REG_0__SCAN_IN | ~P2_U3151;
  assign n16627 = ~n16624 | ~n16623;
  assign n16626 = ~n16949 & ~n16625;
  assign n16633 = ~n16627 & ~n16626;
  assign n16631 = ~n16817 | ~n16628;
  assign n16630 = n9288 ^ n16629;
  assign n16632 = ~n16631 | ~n16630;
  assign P2_U3182 = ~n16633 | ~n16632;
  assign n16637 = ~n16949 & ~n9342;
  assign n16635 = P2_REG1_REG_1__SCAN_IN ^ n16634;
  assign n16636 = ~n16865 & ~n16635;
  assign n16654 = ~n16637 & ~n16636;
  assign n16640 = ~n16639 | ~n16638;
  assign n16642 = ~n16862 | ~n16640;
  assign n16641 = ~P2_REG3_REG_1__SCAN_IN | ~P2_U3151;
  assign n16652 = ~n16642 | ~n16641;
  assign n16650 = ~P2_ADDR_REG_1__SCAN_IN | ~n16945;
  assign n16647 = ~n16643;
  assign n16646 = ~n16645 & ~n16644;
  assign n16648 = ~n16647 & ~n16646;
  assign n16649 = ~n16943 | ~n16648;
  assign n16651 = ~n16650 | ~n16649;
  assign n16653 = ~n16652 & ~n16651;
  assign P2_U3183 = ~n16654 | ~n16653;
  assign n16656 = ~n16924 | ~n11165;
  assign n16655 = ~P2_REG3_REG_2__SCAN_IN | ~P2_U3151;
  assign n16673 = ~n16656 | ~n16655;
  assign n16659 = n16658 & n16657;
  assign n16661 = ~n16660 & ~n16659;
  assign n16671 = ~n16661 | ~n16943;
  assign n16664 = n16663 ^ n16662;
  assign n16669 = ~n16865 & ~n16664;
  assign n16667 = n16666 ^ n16665;
  assign n16668 = ~n16939 & ~n16667;
  assign n16670 = ~n16669 & ~n16668;
  assign n16672 = ~n16671 | ~n16670;
  assign n16675 = ~n16673 & ~n16672;
  assign n16674 = ~n16945 | ~P2_ADDR_REG_2__SCAN_IN;
  assign P2_U3184 = ~n16675 | ~n16674;
  assign n16677 = ~n16676 ^ P2_REG1_REG_3__SCAN_IN;
  assign n16679 = ~n16937 | ~n16677;
  assign n16690 = ~n16679 | ~n16678;
  assign n16682 = ~n16681 ^ n16680;
  assign n16688 = ~n16682 | ~n16943;
  assign n16686 = ~n16949 & ~n17330;
  assign n16684 = n16683 ^ P2_REG2_REG_3__SCAN_IN;
  assign n16685 = ~n16939 & ~n16684;
  assign n16687 = ~n16686 & ~n16685;
  assign n16689 = ~n16688 | ~n16687;
  assign n16692 = ~n16690 & ~n16689;
  assign n16691 = ~n16945 | ~P2_ADDR_REG_3__SCAN_IN;
  assign P2_U3185 = ~n16692 | ~n16691;
  assign n16695 = n16693 ^ n16694;
  assign n16700 = ~n16939 & ~n16695;
  assign n16698 = n16697 ^ n16696;
  assign n16699 = ~n16698 & ~n16865;
  assign n16712 = ~n16700 & ~n16699;
  assign n16703 = ~n16924 | ~n16701;
  assign n16710 = ~n16703 | ~n16702;
  assign n16708 = ~P2_ADDR_REG_4__SCAN_IN | ~n16945;
  assign n16706 = n16705 ^ n16704;
  assign n16707 = ~n16706 | ~n16943;
  assign n16709 = ~n16708 | ~n16707;
  assign n16711 = ~n16710 & ~n16709;
  assign P2_U3186 = ~n16712 | ~n16711;
  assign n16715 = ~n16714 ^ n16713;
  assign n16717 = ~n16715 & ~n16865;
  assign n16716 = ~n16949 & ~n17325;
  assign n16730 = ~n16717 & ~n16716;
  assign n16719 = n16718 ^ P2_REG2_REG_5__SCAN_IN;
  assign n16721 = ~n16719 | ~n16862;
  assign n16728 = ~n16721 | ~n16720;
  assign n16726 = ~P2_ADDR_REG_5__SCAN_IN | ~n16945;
  assign n16724 = n16723 ^ n16722;
  assign n16725 = ~n16724 | ~n16943;
  assign n16727 = ~n16726 | ~n16725;
  assign n16729 = ~n16728 & ~n16727;
  assign P2_U3187 = ~n16730 | ~n16729;
  assign n16733 = ~n16924 | ~n16731;
  assign n16748 = ~n16733 | ~n16732;
  assign n16736 = ~n16735 ^ n16734;
  assign n16746 = ~n16736 | ~n16943;
  assign n16739 = ~n16738 ^ n16737;
  assign n16744 = ~n16739 & ~n16865;
  assign n16742 = n16740 ^ n16741;
  assign n16743 = ~n16742 & ~n16939;
  assign n16745 = ~n16744 & ~n16743;
  assign n16747 = ~n16746 | ~n16745;
  assign n16750 = ~n16748 & ~n16747;
  assign n16749 = ~n16945 | ~P2_ADDR_REG_6__SCAN_IN;
  assign P2_U3188 = ~n16750 | ~n16749;
  assign n16752 = n16751 ^ P2_REG2_REG_7__SCAN_IN;
  assign n16754 = ~n16752 | ~n16862;
  assign n16765 = ~n16754 | ~n16753;
  assign n16757 = ~n16756 ^ n16755;
  assign n16763 = ~n16757 | ~n16943;
  assign n16759 = n16758 ^ P2_REG1_REG_7__SCAN_IN;
  assign n16761 = ~n16759 & ~n16865;
  assign n16760 = ~n16949 & ~n17313;
  assign n16762 = ~n16761 & ~n16760;
  assign n16764 = ~n16763 | ~n16762;
  assign n16767 = ~n16765 & ~n16764;
  assign n16766 = ~n16945 | ~P2_ADDR_REG_7__SCAN_IN;
  assign P2_U3189 = ~n16767 | ~n16766;
  assign n16769 = ~n16768 | ~n16924;
  assign n16784 = ~n16770 | ~n16769;
  assign n16773 = ~n16772 ^ n16771;
  assign n16782 = ~n16773 | ~n16943;
  assign n16776 = n16774 ^ n16775;
  assign n16780 = ~n16776 & ~n16865;
  assign n16778 = n9029 ^ n16777;
  assign n16779 = ~n16778 & ~n16939;
  assign n16781 = ~n16780 & ~n16779;
  assign n16783 = ~n16782 | ~n16781;
  assign n16786 = ~n16784 & ~n16783;
  assign n16785 = ~n16945 | ~P2_ADDR_REG_8__SCAN_IN;
  assign P2_U3190 = ~n16786 | ~n16785;
  assign n16788 = ~P2_REG1_REG_9__SCAN_IN ^ n16787;
  assign n16803 = ~n16788 | ~n16937;
  assign n16790 = ~n16789 ^ P2_REG2_REG_9__SCAN_IN;
  assign n16801 = ~n16790 & ~n16939;
  assign n16793 = ~n16792 ^ n16791;
  assign n16799 = ~n16793 | ~n16943;
  assign n16794 = ~n16945 | ~P2_ADDR_REG_9__SCAN_IN;
  assign n16797 = ~n16795 | ~n16794;
  assign n16796 = ~n16949 & ~n17301;
  assign n16798 = ~n16797 & ~n16796;
  assign n16800 = ~n16799 | ~n16798;
  assign n16802 = ~n16801 & ~n16800;
  assign P2_U3191 = ~n16803 | ~n16802;
  assign n16806 = ~n16805 ^ n16804;
  assign n16812 = ~n16806 | ~n16937;
  assign n16807 = ~n16945 | ~P2_ADDR_REG_10__SCAN_IN;
  assign n16810 = ~n16808 | ~n16807;
  assign n16809 = ~n16949 & ~n17295;
  assign n16811 = ~n16810 & ~n16809;
  assign n16820 = ~n16812 | ~n16811;
  assign n16815 = ~n16814 & ~n16813;
  assign n16818 = ~n16816 ^ n16815;
  assign n16819 = ~n16818 & ~n16817;
  assign n16825 = ~n16820 & ~n16819;
  assign n16823 = ~n16821 ^ n16822;
  assign n16824 = ~n16823 | ~n16862;
  assign P2_U3192 = ~n16825 | ~n16824;
  assign n16827 = ~P2_REG1_REG_11__SCAN_IN ^ n16826;
  assign n16842 = ~n16827 | ~n16937;
  assign n16829 = ~n16828 ^ P2_REG2_REG_11__SCAN_IN;
  assign n16840 = ~n16829 & ~n16939;
  assign n16832 = ~n16831 ^ n16830;
  assign n16838 = ~n16832 | ~n16943;
  assign n16833 = ~n16945 | ~P2_ADDR_REG_11__SCAN_IN;
  assign n16836 = ~n16834 | ~n16833;
  assign n16835 = ~n16949 & ~n17289;
  assign n16837 = ~n16836 & ~n16835;
  assign n16839 = ~n16838 | ~n16837;
  assign n16841 = ~n16840 & ~n16839;
  assign P2_U3193 = ~n16842 | ~n16841;
  assign n16845 = ~n16844 ^ n16843;
  assign n16860 = ~n16845 | ~n16937;
  assign n16847 = n9020 ^ n16846;
  assign n16858 = ~n16847 & ~n16939;
  assign n16850 = ~n16849 ^ n16848;
  assign n16856 = ~n16850 | ~n16943;
  assign n16851 = ~n16945 | ~P2_ADDR_REG_12__SCAN_IN;
  assign n16854 = ~n16852 | ~n16851;
  assign n16853 = ~n16949 & ~n17283;
  assign n16855 = ~n16854 & ~n16853;
  assign n16857 = ~n16856 | ~n16855;
  assign n16859 = ~n16858 & ~n16857;
  assign P2_U3194 = ~n16860 | ~n16859;
  assign n16863 = P2_REG2_REG_13__SCAN_IN ^ n16861;
  assign n16879 = ~n16863 | ~n16862;
  assign n16866 = n16864 ^ P2_REG1_REG_13__SCAN_IN;
  assign n16877 = ~n16866 & ~n16865;
  assign n16869 = ~n16868 ^ n16867;
  assign n16875 = ~n16869 | ~n16943;
  assign n16870 = ~n16945 | ~P2_ADDR_REG_13__SCAN_IN;
  assign n16873 = ~n16871 | ~n16870;
  assign n16872 = ~n16949 & ~n17277;
  assign n16874 = ~n16873 & ~n16872;
  assign n16876 = ~n16875 | ~n16874;
  assign n16878 = ~n16877 & ~n16876;
  assign P2_U3195 = ~n16879 | ~n16878;
  assign n16882 = ~n16881 ^ n16880;
  assign n16898 = ~n16882 | ~n16937;
  assign n16884 = n8901 ^ n16883;
  assign n16896 = ~n16884 & ~n16939;
  assign n16887 = ~n16886 ^ n16885;
  assign n16894 = ~n16887 | ~n16943;
  assign n16890 = ~n16945 | ~P2_ADDR_REG_14__SCAN_IN;
  assign n16889 = ~n16888 | ~n16924;
  assign n16891 = ~n16890 | ~n16889;
  assign n16893 = ~n16892 & ~n16891;
  assign n16895 = ~n16894 | ~n16893;
  assign n16897 = ~n16896 & ~n16895;
  assign P2_U3196 = ~n16898 | ~n16897;
  assign n16900 = ~P2_REG1_REG_15__SCAN_IN ^ n16899;
  assign n16915 = ~n16900 | ~n16937;
  assign n16902 = ~P2_REG2_REG_15__SCAN_IN ^ n16901;
  assign n16913 = ~n16902 & ~n16939;
  assign n16905 = ~n16904 ^ n16903;
  assign n16911 = ~n16905 | ~n16943;
  assign n16906 = ~n16945 | ~P2_ADDR_REG_15__SCAN_IN;
  assign n16909 = ~n16907 | ~n16906;
  assign n16908 = ~n16949 & ~n17266;
  assign n16910 = ~n16909 & ~n16908;
  assign n16912 = ~n16911 | ~n16910;
  assign n16914 = ~n16913 & ~n16912;
  assign P2_U3197 = ~n16915 | ~n16914;
  assign n16918 = ~n16917 ^ n16916;
  assign n16935 = ~n16918 | ~n16937;
  assign n16920 = n8987 ^ n16919;
  assign n16933 = ~n16920 & ~n16939;
  assign n16923 = ~n16922 ^ n16921;
  assign n16931 = ~n16923 | ~n16943;
  assign n16927 = ~n16945 | ~P2_ADDR_REG_16__SCAN_IN;
  assign n16926 = ~n16925 | ~n16924;
  assign n16928 = ~n16927 | ~n16926;
  assign n16930 = ~n16929 & ~n16928;
  assign n16932 = ~n16931 | ~n16930;
  assign n16934 = ~n16933 & ~n16932;
  assign P2_U3198 = ~n16935 | ~n16934;
  assign n16938 = ~P2_REG1_REG_17__SCAN_IN ^ n16936;
  assign n16957 = ~n16938 | ~n16937;
  assign n16955 = ~n16940 & ~n16939;
  assign n16944 = ~n16942 ^ n16941;
  assign n16953 = ~n16944 | ~n16943;
  assign n16946 = ~n16945 | ~P2_ADDR_REG_17__SCAN_IN;
  assign n16951 = ~n16947 | ~n16946;
  assign n16950 = ~n16949 & ~n16948;
  assign n16952 = ~n16951 & ~n16950;
  assign n16954 = ~n16953 | ~n16952;
  assign n16956 = ~n16955 & ~n16954;
  assign P2_U3199 = ~n16957 | ~n16956;
  assign n16960 = ~P2_REG2_REG_11__SCAN_IN | ~n17200;
  assign n16959 = ~n17197 | ~n16958;
  assign n16966 = ~n16960 | ~n16959;
  assign n16963 = ~n16993 | ~n16961;
  assign n16964 = ~n16963 | ~n16962;
  assign n17450 = n16972 ^ n16964;
  assign n16965 = ~n17450 & ~n17128;
  assign n16982 = ~n16966 & ~n16965;
  assign n16970 = ~n16968 | ~n16967;
  assign n16971 = ~n16970 | ~n16969;
  assign n16973 = n16972 ^ n16971;
  assign n16978 = ~n16973 & ~n17356;
  assign n16976 = ~n16974 | ~n17464;
  assign n16975 = ~n16989 | ~n17166;
  assign n16977 = ~n16976 | ~n16975;
  assign n17457 = ~n16978 & ~n16977;
  assign n16979 = ~n17451 | ~n17185;
  assign n16980 = ~n17457 | ~n16979;
  assign n16981 = ~n17209 | ~n16980;
  assign P2_U3222 = ~n16982 | ~n16981;
  assign n16986 = ~n16983 & ~n17120;
  assign n16985 = ~n17209 & ~n16984;
  assign n17003 = ~n16986 & ~n16985;
  assign n16988 = ~n16987 ^ n16992;
  assign n16997 = ~n16988 | ~n17172;
  assign n16991 = ~n17166 | ~n17036;
  assign n16990 = ~n17464 | ~n16989;
  assign n16995 = ~n16991 | ~n16990;
  assign n17432 = ~n16993 ^ n16992;
  assign n16994 = ~n17083 & ~n17432;
  assign n16996 = ~n16995 & ~n16994;
  assign n17431 = ~n16997 | ~n16996;
  assign n16998 = ~n17088 & ~n17432;
  assign n16999 = ~n17431 & ~n16998;
  assign n17001 = ~n17200 & ~n16999;
  assign n17000 = ~n17123 & ~n17429;
  assign n17002 = ~n17001 & ~n17000;
  assign P2_U3224 = ~n17003 | ~n17002;
  assign n17006 = ~n17029 | ~n17004;
  assign n17007 = n17006 & n17005;
  assign n17008 = n17014 ^ n17007;
  assign n17013 = ~n17008 & ~n17356;
  assign n17011 = ~n17009 | ~n17464;
  assign n17010 = ~n17053 | ~n17166;
  assign n17012 = ~n17011 | ~n17010;
  assign n17426 = ~n17013 & ~n17012;
  assign n17421 = ~n17015 ^ n17014;
  assign n17016 = n17421 | n17108;
  assign n17017 = ~n17426 | ~n17016;
  assign n17026 = ~n17017 | ~n17209;
  assign n17021 = ~n17196 | ~n17018;
  assign n17020 = ~n17197 | ~n17019;
  assign n17024 = ~n17021 | ~n17020;
  assign n17023 = ~n17022 & ~n17209;
  assign n17025 = ~n17024 & ~n17023;
  assign P2_U3225 = ~n17026 | ~n17025;
  assign n17413 = ~n17027 ^ n17030;
  assign n17033 = ~n17413;
  assign n17041 = ~n17033 | ~n17183;
  assign n17031 = ~n17029 | ~n17028;
  assign n17032 = ~n17031 ^ n17030;
  assign n17035 = ~n17032 | ~n17172;
  assign n17034 = ~n17033 | ~n17178;
  assign n17040 = ~n17035 | ~n17034;
  assign n17038 = ~n17078 | ~n17166;
  assign n17037 = ~n17036 | ~n17464;
  assign n17039 = ~n17038 | ~n17037;
  assign n17418 = ~n17040 & ~n17039;
  assign n17042 = ~n17041 | ~n17418;
  assign n17050 = ~n17042 | ~n17209;
  assign n17045 = ~n17196 | ~n17043;
  assign n17044 = ~n17200 | ~P2_REG2_REG_7__SCAN_IN;
  assign n17048 = ~n17045 | ~n17044;
  assign n17047 = ~n17046 & ~n17120;
  assign n17049 = ~n17048 & ~n17047;
  assign P2_U3226 = ~n17050 | ~n17049;
  assign n17052 = n17059 ^ n17051;
  assign n17057 = ~n17052 & ~n17356;
  assign n17055 = ~n17053 | ~n17464;
  assign n17054 = ~n17102 | ~n17166;
  assign n17056 = ~n17055 | ~n17054;
  assign n17410 = ~n17057 & ~n17056;
  assign n17405 = n17058 ^ n17059;
  assign n17060 = n17405 | n17108;
  assign n17061 = ~n17410 | ~n17060;
  assign n17069 = ~n17061 | ~n17209;
  assign n17064 = ~n17196 | ~n17062;
  assign n17063 = ~n17200 | ~P2_REG2_REG_6__SCAN_IN;
  assign n17067 = ~n17064 | ~n17063;
  assign n17066 = ~n17065 & ~n17120;
  assign n17068 = ~n17067 & ~n17066;
  assign P2_U3227 = ~n17069 | ~n17068;
  assign n17073 = ~n17070 & ~n17209;
  assign n17072 = ~n17071 & ~n17120;
  assign n17094 = ~n17073 & ~n17072;
  assign n17076 = ~n17075 | ~n17074;
  assign n17077 = ~n17076 ^ n17082;
  assign n17087 = ~n17077 | ~n17172;
  assign n17080 = ~n17166 | ~n17132;
  assign n17079 = ~n17464 | ~n17078;
  assign n17085 = ~n17080 | ~n17079;
  assign n17399 = n17081 ^ n17082;
  assign n17084 = ~n17399 & ~n17083;
  assign n17086 = ~n17085 & ~n17084;
  assign n17398 = ~n17087 | ~n17086;
  assign n17089 = ~n17399 & ~n17088;
  assign n17090 = ~n17398 & ~n17089;
  assign n17092 = ~n17200 & ~n17090;
  assign n17091 = ~n17123 & ~n17396;
  assign n17093 = ~n17092 & ~n17091;
  assign P2_U3228 = ~n17094 | ~n17093;
  assign n17130 = ~n17096 | ~n17095;
  assign n17099 = ~n17130 | ~n17097;
  assign n17100 = ~n17099 | ~n17098;
  assign n17101 = n17107 ^ n17100;
  assign n17106 = ~n17101 & ~n17356;
  assign n17104 = ~n17150 | ~n17166;
  assign n17103 = ~n17102 | ~n17464;
  assign n17105 = ~n17104 | ~n17103;
  assign n17393 = ~n17106 & ~n17105;
  assign n17109 = n17388 | n17108;
  assign n17110 = ~n17393 | ~n17109;
  assign n17119 = ~n17110 | ~n17209;
  assign n17114 = ~n17196 | ~n17111;
  assign n17113 = ~n17197 | ~n17112;
  assign n17117 = ~n17114 | ~n17113;
  assign n17116 = ~n17115 & ~n17209;
  assign n17118 = ~n17117 & ~n17116;
  assign P2_U3229 = ~n17119 | ~n17118;
  assign n17122 = ~P2_REG2_REG_3__SCAN_IN | ~n17200;
  assign n17121 = n17120 | P2_REG3_REG_3__SCAN_IN;
  assign n17125 = ~n17122 | ~n17121;
  assign n17124 = ~n17123 & ~n17381;
  assign n17140 = ~n17125 & ~n17124;
  assign n17380 = ~n17127 ^ n17126;
  assign n17138 = ~n17380 & ~n17128;
  assign n17131 = ~n17130 ^ n17129;
  assign n17136 = ~n17131 & ~n17356;
  assign n17134 = ~n17132 | ~n17464;
  assign n17133 = ~n17168 | ~n17166;
  assign n17135 = ~n17134 | ~n17133;
  assign n17385 = ~n17136 & ~n17135;
  assign n17137 = ~n17200 & ~n17385;
  assign n17139 = ~n17138 & ~n17137;
  assign P2_U3230 = ~n17140 | ~n17139;
  assign n17144 = ~n17141;
  assign n17372 = ~n17144 & ~n17143;
  assign n17157 = ~n17372;
  assign n17146 = ~n17157 | ~n17183;
  assign n17145 = ~P2_REG3_REG_2__SCAN_IN | ~n17197;
  assign n17149 = ~n17146 | ~n17145;
  assign n17148 = ~n17373 & ~n17147;
  assign n17162 = ~n17149 & ~n17148;
  assign n17153 = ~n17150 | ~n17464;
  assign n17152 = ~n17151 | ~n17166;
  assign n17161 = ~n17153 | ~n17152;
  assign n17156 = ~n17155 ^ n17154;
  assign n17159 = ~n17156 | ~n17172;
  assign n17158 = ~n17157 | ~n17178;
  assign n17160 = ~n17159 | ~n17158;
  assign n17377 = ~n17161 & ~n17160;
  assign n17163 = ~n17162 | ~n17377;
  assign n17165 = ~n17209 | ~n17163;
  assign n17164 = ~n17200 | ~P2_REG2_REG_2__SCAN_IN;
  assign P2_U3231 = ~n17165 | ~n17164;
  assign n17170 = ~n17167 | ~n17166;
  assign n17169 = ~n17168 | ~n17464;
  assign n17182 = ~n17170 | ~n17169;
  assign n17173 = ~n17175 ^ n17171;
  assign n17180 = ~n17173 | ~n17172;
  assign n17176 = ~n17175 | ~n17174;
  assign n17363 = ~n17177 | ~n17176;
  assign n17179 = ~n17363 | ~n17178;
  assign n17181 = ~n17180 | ~n17179;
  assign n17369 = ~n17182 & ~n17181;
  assign n17189 = ~n17369;
  assign n17187 = ~n17363 | ~n17183;
  assign n17186 = ~n17185 | ~n17184;
  assign n17188 = ~n17187 | ~n17186;
  assign n17190 = ~n17189 & ~n17188;
  assign n17192 = ~n17200 & ~n17190;
  assign n17191 = ~n17209 & ~n9632;
  assign n17194 = ~n17192 & ~n17191;
  assign n17193 = ~P2_REG3_REG_1__SCAN_IN | ~n17197;
  assign P2_U3232 = ~n17194 | ~n17193;
  assign n17199 = ~n17196 | ~n17195;
  assign n17198 = ~n17197 | ~P2_REG3_REG_0__SCAN_IN;
  assign n17202 = ~n17199 | ~n17198;
  assign n17201 = P2_REG2_REG_0__SCAN_IN & n17200;
  assign n17212 = ~n17202 & ~n17201;
  assign n17355 = ~n17204 & ~n17203;
  assign n17208 = ~n17355;
  assign n17206 = ~n17205 & ~n17462;
  assign n17207 = ~n17358 | ~n17206;
  assign n17210 = ~n17208 | ~n17207;
  assign n17211 = ~n17210 | ~n17209;
  assign P2_U3233 = ~n17212 | ~n17211;
  assign n17216 = ~n17213 & ~n17341;
  assign n17215 = ~n17214 & ~P2_U3151;
  assign n17218 = ~n17216 & ~n17215;
  assign n17217 = ~n17338 | ~P1_DATAO_REG_25__SCAN_IN;
  assign P2_U3270 = ~n17218 | ~n17217;
  assign n17221 = ~n17219 & ~n17341;
  assign n17220 = ~n11323 & ~P2_U3151;
  assign n17223 = ~n17221 & ~n17220;
  assign n17222 = ~n17338 | ~P1_DATAO_REG_24__SCAN_IN;
  assign P2_U3271 = ~n17223 | ~n17222;
  assign n17228 = ~n17224 & ~n17341;
  assign n17225 = ~P1_DATAO_REG_23__SCAN_IN;
  assign n17227 = ~n17226 & ~n17225;
  assign n17230 = ~n17228 & ~n17227;
  assign P2_U3272 = ~n17230 | ~n17229;
  assign n17234 = ~n17231 & ~n17341;
  assign n17233 = ~n17232 & ~P2_U3151;
  assign n17236 = ~n17234 & ~n17233;
  assign n17235 = ~n17338 | ~P1_DATAO_REG_22__SCAN_IN;
  assign P2_U3273 = ~n17236 | ~n17235;
  assign n17240 = ~n17237 & ~n17341;
  assign n17239 = ~n17238 & ~P2_U3151;
  assign n17242 = ~n17240 & ~n17239;
  assign n17241 = ~n17338 | ~P1_DATAO_REG_21__SCAN_IN;
  assign P2_U3274 = ~n17242 | ~n17241;
  assign n17245 = ~n12213 & ~n17341;
  assign n17244 = ~n17243 & ~P2_U3151;
  assign n17247 = ~n17245 & ~n17244;
  assign n17246 = ~n17338 | ~P1_DATAO_REG_20__SCAN_IN;
  assign P2_U3275 = ~n17247 | ~n17246;
  assign n17250 = ~n17248 & ~n17341;
  assign n17249 = ~n11117 & ~P2_U3151;
  assign n17252 = ~n17250 & ~n17249;
  assign n17251 = ~n17338 | ~P1_DATAO_REG_19__SCAN_IN;
  assign P2_U3276 = ~n17252 | ~n17251;
  assign n17256 = ~n17253 & ~n17341;
  assign n17255 = ~n17254 & ~P2_U3151;
  assign n17258 = ~n17256 & ~n17255;
  assign n17257 = ~n17338 | ~P1_DATAO_REG_18__SCAN_IN;
  assign P2_U3277 = ~n17258 | ~n17257;
  assign n17262 = ~n17259 & ~n17341;
  assign n17261 = ~n17260 & ~P2_U3151;
  assign n17264 = ~n17262 & ~n17261;
  assign n17263 = ~n17338 | ~P1_DATAO_REG_16__SCAN_IN;
  assign P2_U3279 = ~n17264 | ~n17263;
  assign n17268 = ~n17265 & ~n17341;
  assign n17267 = ~n17266 & ~P2_U3151;
  assign n17270 = ~n17268 & ~n17267;
  assign n17269 = ~n17338 | ~P1_DATAO_REG_15__SCAN_IN;
  assign P2_U3280 = ~n17270 | ~n17269;
  assign n17273 = ~n12157 & ~n17341;
  assign n17272 = ~n17271 & ~P2_U3151;
  assign n17275 = ~n17273 & ~n17272;
  assign n17274 = ~n17338 | ~P1_DATAO_REG_14__SCAN_IN;
  assign P2_U3281 = ~n17275 | ~n17274;
  assign n17279 = ~n17276 & ~n17341;
  assign n17278 = ~n17277 & ~P2_U3151;
  assign n17281 = ~n17279 & ~n17278;
  assign n17280 = ~n17338 | ~P1_DATAO_REG_13__SCAN_IN;
  assign P2_U3282 = ~n17281 | ~n17280;
  assign n17285 = ~n17282 & ~n17341;
  assign n17284 = ~n17283 & ~P2_U3151;
  assign n17287 = ~n17285 & ~n17284;
  assign n17286 = ~n17338 | ~P1_DATAO_REG_12__SCAN_IN;
  assign P2_U3283 = ~n17287 | ~n17286;
  assign n17291 = ~n17288 & ~n17341;
  assign n17290 = ~n17289 & ~P2_U3151;
  assign n17293 = ~n17291 & ~n17290;
  assign n17292 = ~n17338 | ~P1_DATAO_REG_11__SCAN_IN;
  assign P2_U3284 = ~n17293 | ~n17292;
  assign n17297 = ~n17294 & ~n17341;
  assign n17296 = ~n17295 & ~P2_U3151;
  assign n17299 = ~n17297 & ~n17296;
  assign n17298 = ~n17338 | ~P1_DATAO_REG_10__SCAN_IN;
  assign P2_U3285 = ~n17299 | ~n17298;
  assign n17303 = ~n17300 & ~n17341;
  assign n17302 = ~n17301 & ~P2_U3151;
  assign n17305 = ~n17303 & ~n17302;
  assign n17304 = ~n17338 | ~P1_DATAO_REG_9__SCAN_IN;
  assign P2_U3286 = ~n17305 | ~n17304;
  assign n17309 = ~n17306 & ~n17341;
  assign n17308 = ~n17307 & ~P2_U3151;
  assign n17311 = ~n17309 & ~n17308;
  assign n17310 = ~n17338 | ~P1_DATAO_REG_8__SCAN_IN;
  assign P2_U3287 = ~n17311 | ~n17310;
  assign n17315 = ~n17312 & ~n17341;
  assign n17314 = ~n17313 & ~P2_U3151;
  assign n17317 = ~n17315 & ~n17314;
  assign n17316 = ~n17338 | ~P1_DATAO_REG_7__SCAN_IN;
  assign P2_U3288 = ~n17317 | ~n17316;
  assign n17321 = ~n17318 & ~n17341;
  assign n17320 = ~n17319 & ~P2_U3151;
  assign n17323 = ~n17321 & ~n17320;
  assign n17322 = ~n17338 | ~P1_DATAO_REG_6__SCAN_IN;
  assign P2_U3289 = ~n17323 | ~n17322;
  assign n17327 = ~n17324 & ~n17341;
  assign n17326 = ~n17325 & ~P2_U3151;
  assign n17329 = ~n17327 & ~n17326;
  assign n17328 = ~n17338 | ~P1_DATAO_REG_5__SCAN_IN;
  assign P2_U3290 = ~n17329 | ~n17328;
  assign n17332 = ~n12066 & ~n17341;
  assign n17331 = ~n17330 & ~P2_U3151;
  assign n17334 = ~n17332 & ~n17331;
  assign n17333 = ~n17338 | ~P1_DATAO_REG_3__SCAN_IN;
  assign P2_U3292 = ~n17334 | ~n17333;
  assign n17337 = ~n12056 & ~n17341;
  assign n17336 = ~n9360 & ~P2_U3151;
  assign n17340 = ~n17337 & ~n17336;
  assign n17339 = ~n17338 | ~P1_DATAO_REG_2__SCAN_IN;
  assign P2_U3293 = ~n17340 | ~n17339;
  assign n17345 = ~n17342 & ~n17341;
  assign n17344 = ~n9342 & ~P2_U3151;
  assign n17347 = ~n17345 & ~n17344;
  assign n17346 = ~n17338 | ~P1_DATAO_REG_1__SCAN_IN;
  assign P2_U3294 = ~n17347 | ~n17346;
  assign n17352 = ~P2_D_REG_1__SCAN_IN | ~n17348;
  assign n17351 = ~n17350 | ~n17349;
  assign P2_U3377 = ~n17352 | ~n17351;
  assign n17362 = ~P2_REG0_REG_0__SCAN_IN | ~n17460;
  assign n17354 = ~n17353 & ~n17452;
  assign n17360 = ~n17355 & ~n17354;
  assign n17357 = ~n17449 | ~n17356;
  assign n17359 = ~n17358 | ~n17357;
  assign n17475 = ~n17360 | ~n17359;
  assign n17361 = ~n17472 | ~n17475;
  assign P2_U3390 = ~n17362 | ~n17361;
  assign n17371 = ~P2_REG0_REG_1__SCAN_IN | ~n17460;
  assign n17364 = ~n17363;
  assign n17367 = ~n17364 & ~n17440;
  assign n17366 = ~n17365 & ~n17452;
  assign n17368 = ~n17367 & ~n17366;
  assign n17478 = ~n17369 | ~n17368;
  assign n17370 = ~n17472 | ~n17478;
  assign P2_U3393 = ~n17371 | ~n17370;
  assign n17379 = ~P2_REG0_REG_2__SCAN_IN | ~n17460;
  assign n17375 = ~n17372 & ~n17440;
  assign n17374 = ~n17373 & ~n17452;
  assign n17376 = ~n17375 & ~n17374;
  assign n17481 = ~n17377 | ~n17376;
  assign n17378 = ~n17472 | ~n17481;
  assign P2_U3396 = ~n17379 | ~n17378;
  assign n17387 = ~P2_REG0_REG_3__SCAN_IN | ~n17460;
  assign n17383 = ~n17380 & ~n17449;
  assign n17382 = ~n17381 & ~n17452;
  assign n17384 = ~n17383 & ~n17382;
  assign n17484 = ~n17385 | ~n17384;
  assign n17386 = ~n17472 | ~n17484;
  assign P2_U3399 = ~n17387 | ~n17386;
  assign n17395 = ~P2_REG0_REG_4__SCAN_IN | ~n17460;
  assign n17391 = ~n17388 & ~n17449;
  assign n17390 = ~n17389 & ~n17452;
  assign n17392 = ~n17391 & ~n17390;
  assign n17487 = ~n17393 | ~n17392;
  assign n17394 = ~n17472 | ~n17487;
  assign P2_U3402 = ~n17395 | ~n17394;
  assign n17404 = ~P2_REG0_REG_5__SCAN_IN | ~n17460;
  assign n17397 = ~n17396 & ~n17452;
  assign n17402 = ~n17398 & ~n17397;
  assign n17400 = ~n17399;
  assign n17433 = ~n17440;
  assign n17401 = ~n17400 | ~n17433;
  assign n17490 = ~n17402 | ~n17401;
  assign n17403 = ~n17472 | ~n17490;
  assign P2_U3405 = ~n17404 | ~n17403;
  assign n17412 = ~P2_REG0_REG_6__SCAN_IN | ~n17460;
  assign n17408 = ~n17405 & ~n17449;
  assign n17407 = ~n17406 & ~n17452;
  assign n17409 = ~n17408 & ~n17407;
  assign n17493 = ~n17410 | ~n17409;
  assign n17411 = ~n17472 | ~n17493;
  assign P2_U3408 = ~n17412 | ~n17411;
  assign n17420 = ~P2_REG0_REG_7__SCAN_IN | ~n17460;
  assign n17416 = ~n17413 & ~n17440;
  assign n17415 = ~n17414 & ~n17452;
  assign n17417 = ~n17416 & ~n17415;
  assign n17496 = ~n17418 | ~n17417;
  assign n17419 = ~n17472 | ~n17496;
  assign P2_U3411 = ~n17420 | ~n17419;
  assign n17428 = ~P2_REG0_REG_8__SCAN_IN | ~n17460;
  assign n17424 = ~n17421 & ~n17449;
  assign n17423 = ~n17422 & ~n17452;
  assign n17425 = ~n17424 & ~n17423;
  assign n17499 = ~n17426 | ~n17425;
  assign n17427 = ~n17472 | ~n17499;
  assign P2_U3414 = ~n17428 | ~n17427;
  assign n17438 = ~P2_REG0_REG_9__SCAN_IN | ~n17460;
  assign n17430 = ~n17429 & ~n17452;
  assign n17436 = ~n17431 & ~n17430;
  assign n17434 = ~n17432;
  assign n17435 = ~n17434 | ~n17433;
  assign n17502 = ~n17436 | ~n17435;
  assign n17437 = ~n17472 | ~n17502;
  assign P2_U3417 = ~n17438 | ~n17437;
  assign n17448 = ~P2_REG0_REG_10__SCAN_IN | ~n17460;
  assign n17446 = ~n17439;
  assign n17444 = ~n17441 & ~n17440;
  assign n17443 = ~n17442 & ~n17452;
  assign n17445 = ~n17444 & ~n17443;
  assign n17505 = ~n17446 | ~n17445;
  assign n17447 = ~n17472 | ~n17505;
  assign P2_U3420 = ~n17448 | ~n17447;
  assign n17459 = ~P2_REG0_REG_11__SCAN_IN | ~n17460;
  assign n17455 = ~n17450 & ~n17449;
  assign n17453 = ~n17451;
  assign n17454 = ~n17453 & ~n17452;
  assign n17456 = ~n17455 & ~n17454;
  assign n17508 = ~n17457 | ~n17456;
  assign n17458 = ~n17472 | ~n17508;
  assign P2_U3423 = ~n17459 | ~n17458;
  assign n17474 = ~P2_REG0_REG_12__SCAN_IN | ~n17460;
  assign n17471 = ~n17461 | ~n9107;
  assign n17467 = ~n17463 | ~n17462;
  assign n17466 = ~n17465 | ~n17464;
  assign n17468 = ~n17467 | ~n17466;
  assign n17470 = ~n17469 & ~n17468;
  assign n17513 = ~n17471 | ~n17470;
  assign n17473 = ~n17513 | ~n17472;
  assign P2_U3426 = ~n17474 | ~n17473;
  assign n17477 = ~P2_REG1_REG_0__SCAN_IN | ~n17511;
  assign n17476 = ~n17512 | ~n17475;
  assign P2_U3459 = ~n17477 | ~n17476;
  assign n17480 = ~P2_REG1_REG_1__SCAN_IN | ~n17511;
  assign n17479 = ~n17512 | ~n17478;
  assign P2_U3460 = ~n17480 | ~n17479;
  assign n17483 = ~P2_REG1_REG_2__SCAN_IN | ~n17511;
  assign n17482 = ~n17512 | ~n17481;
  assign P2_U3461 = ~n17483 | ~n17482;
  assign n17486 = ~P2_REG1_REG_3__SCAN_IN | ~n17511;
  assign n17485 = ~n17512 | ~n17484;
  assign P2_U3462 = ~n17486 | ~n17485;
  assign n17489 = ~P2_REG1_REG_4__SCAN_IN | ~n17511;
  assign n17488 = ~n17512 | ~n17487;
  assign P2_U3463 = ~n17489 | ~n17488;
  assign n17492 = ~P2_REG1_REG_5__SCAN_IN | ~n17511;
  assign n17491 = ~n17512 | ~n17490;
  assign P2_U3464 = ~n17492 | ~n17491;
  assign n17495 = ~P2_REG1_REG_6__SCAN_IN | ~n17511;
  assign n17494 = ~n17512 | ~n17493;
  assign P2_U3465 = ~n17495 | ~n17494;
  assign n17498 = ~P2_REG1_REG_7__SCAN_IN | ~n17511;
  assign n17497 = ~n17512 | ~n17496;
  assign P2_U3466 = ~n17498 | ~n17497;
  assign n17501 = ~P2_REG1_REG_8__SCAN_IN | ~n17511;
  assign n17500 = ~n17512 | ~n17499;
  assign P2_U3467 = ~n17501 | ~n17500;
  assign n17504 = ~P2_REG1_REG_9__SCAN_IN | ~n17511;
  assign n17503 = ~n17512 | ~n17502;
  assign P2_U3468 = ~n17504 | ~n17503;
  assign n17507 = ~P2_REG1_REG_10__SCAN_IN | ~n17511;
  assign n17506 = ~n17512 | ~n17505;
  assign P2_U3469 = ~n17507 | ~n17506;
  assign n17510 = ~P2_REG1_REG_11__SCAN_IN | ~n17511;
  assign n17509 = ~n17512 | ~n17508;
  assign P2_U3470 = ~n17510 | ~n17509;
  assign n17515 = ~P2_REG1_REG_12__SCAN_IN | ~n17511;
  assign n17514 = ~n17513 | ~n17512;
  assign P2_U3471 = ~n17515 | ~n17514;
  assign n17518 = ~P2_DATAO_REG_20__SCAN_IN | ~n17550;
  assign n17517 = ~P2_U3893 | ~n17516;
  assign P2_U3511 = ~n17518 | ~n17517;
  assign n17521 = ~P2_DATAO_REG_21__SCAN_IN | ~n17550;
  assign n17520 = ~P2_U3893 | ~n17519;
  assign P2_U3512 = ~n17521 | ~n17520;
  assign n17524 = ~P2_DATAO_REG_22__SCAN_IN | ~n17550;
  assign n17523 = ~P2_U3893 | ~n17522;
  assign P2_U3513 = ~n17524 | ~n17523;
  assign n17528 = ~P2_DATAO_REG_23__SCAN_IN | ~n17550;
  assign n17527 = ~P2_U3893 | ~n17525;
  assign P2_U3514 = ~n17528 | ~n17527;
  assign n17531 = ~P2_DATAO_REG_24__SCAN_IN | ~n17550;
  assign n17530 = ~P2_U3893 | ~n17529;
  assign P2_U3515 = ~n17531 | ~n17530;
  assign n17534 = ~P2_DATAO_REG_25__SCAN_IN | ~n17550;
  assign n17533 = ~P2_U3893 | ~n17532;
  assign P2_U3516 = ~n17534 | ~n17533;
  assign n17537 = ~P2_DATAO_REG_26__SCAN_IN | ~n17550;
  assign n17536 = ~P2_U3893 | ~n17535;
  assign P2_U3517 = ~n17537 | ~n17536;
  assign n17540 = ~P2_DATAO_REG_27__SCAN_IN | ~n17550;
  assign n17539 = ~P2_U3893 | ~n17538;
  assign P2_U3518 = ~n17540 | ~n17539;
  assign n17543 = ~P2_DATAO_REG_28__SCAN_IN | ~n17550;
  assign n17542 = ~P2_U3893 | ~n17541;
  assign P2_U3519 = ~n17543 | ~n17542;
  assign n17546 = ~P2_DATAO_REG_29__SCAN_IN | ~n17550;
  assign n17545 = ~P2_U3893 | ~n17544;
  assign P2_U3520 = ~n17546 | ~n17545;
  assign n17549 = ~P2_DATAO_REG_30__SCAN_IN | ~n17550;
  assign n17548 = n17550 | n17547;
  assign P2_U3521 = ~n17549 | ~n17548;
  assign n17553 = ~P2_DATAO_REG_31__SCAN_IN | ~n17550;
  assign n17552 = ~P2_U3893 | ~n17551;
  assign P2_U3522 = ~n17553 | ~n17552;
  assign n17556 = ~n17555 & ~n17554;
  assign ADD_1068_U5 = P2_ADDR_REG_1__SCAN_IN ^ n17556;
  assign ADD_1068_U46 = P1_ADDR_REG_0__SCAN_IN ^ P2_ADDR_REG_0__SCAN_IN;
  assign ADD_1068_U47 = ~n17558 ^ n17557;
  assign ADD_1068_U48 = ~n17560 ^ n17559;
  assign ADD_1068_U49 = ~n17562 ^ n17561;
  assign ADD_1068_U50 = ~n17564 ^ n17563;
  assign ADD_1068_U51 = ~n17566 ^ n17565;
  assign ADD_1068_U52 = ~n17568 ^ n17567;
  assign ADD_1068_U53 = n17570 ^ n17569;
  assign ADD_1068_U54 = n17572 ^ n17571;
  assign n17576 = ~n17574 | ~n17573;
  assign ADD_1068_U55 = ~n17576 ^ n17575;
  assign n17579 = ~n17578 & ~n17577;
  assign ADD_1068_U56 = n17580 ^ n17579;
  assign n17583 = ~n17582 & ~n17581;
  assign ADD_1068_U57 = n17584 ^ n17583;
  assign n17587 = ~n17586 & ~n17585;
  assign ADD_1068_U58 = n17588 ^ n17587;
  assign n17591 = ~n17590 & ~n17589;
  assign ADD_1068_U59 = n17592 ^ n17591;
  assign n17595 = ~n17594 & ~n17593;
  assign ADD_1068_U60 = n17596 ^ n17595;
  assign n17599 = ~n17598 & ~n17597;
  assign ADD_1068_U61 = n17600 ^ n17599;
  assign n17603 = ~n17602 & ~n17601;
  assign ADD_1068_U62 = n17604 ^ n17603;
  assign n17607 = ~n17606 & ~n17605;
  assign ADD_1068_U63 = n17608 ^ n17607;
  assign n13271 = n10286;
  assign n9976 = ~n9920;
  assign n11273 = ~n11282;
  assign n13056 = n10079 & n10078;
  assign n13065 = n10052 & n10051;
  assign n17237 = ~n10621 ^ n10650;
endmodule


