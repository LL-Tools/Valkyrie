

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput127, keyinput126, keyinput125, keyinput124, keyinput123, 
        keyinput122, keyinput121, keyinput120, keyinput119, keyinput118, 
        keyinput117, keyinput116, keyinput115, keyinput114, keyinput113, 
        keyinput112, keyinput111, keyinput110, keyinput109, keyinput108, 
        keyinput107, keyinput106, keyinput105, keyinput104, keyinput103, 
        keyinput102, keyinput101, keyinput100, keyinput99, keyinput98, 
        keyinput97, keyinput96, keyinput95, keyinput94, keyinput93, keyinput92, 
        keyinput91, keyinput90, keyinput89, keyinput88, keyinput87, keyinput86, 
        keyinput85, keyinput84, keyinput83, keyinput82, keyinput81, keyinput80, 
        keyinput79, keyinput78, keyinput77, keyinput76, keyinput75, keyinput74, 
        keyinput73, keyinput72, keyinput71, keyinput70, keyinput69, keyinput68, 
        keyinput67, keyinput66, keyinput65, keyinput64, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4409, n4410, n4411, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433;

  MUX2_X1 U4915 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9357), .S(n4525), .Z(n9359) );
  NAND2_X1 U4916 ( .A1(n5322), .A2(n5202), .ZN(n5169) );
  NAND2_X2 U4917 ( .A1(n5851), .A2(n7300), .ZN(n9613) );
  INV_X2 U4919 ( .A(n5129), .ZN(n5171) );
  NAND2_X1 U4920 ( .A1(n5057), .A2(n5089), .ZN(n5092) );
  INV_X1 U4921 ( .A(n5600), .ZN(n5220) );
  INV_X1 U4923 ( .A(n5946), .ZN(n6165) );
  INV_X1 U4925 ( .A(n5322), .ZN(n5745) );
  INV_X2 U4926 ( .A(n5345), .ZN(n5445) );
  AND3_X1 U4927 ( .A1(n5961), .A2(n5960), .A3(n5031), .ZN(n7232) );
  NAND2_X1 U4928 ( .A1(n5946), .A2(n5212), .ZN(n6004) );
  INV_X1 U4930 ( .A(n6332), .ZN(n8285) );
  AND2_X1 U4931 ( .A1(n8197), .A2(n8186), .ZN(n8345) );
  OR2_X1 U4932 ( .A1(n5088), .A2(n5089), .ZN(n5091) );
  NOR2_X2 U4933 ( .A1(n9886), .A2(n9878), .ZN(n9858) );
  INV_X1 U4934 ( .A(n7140), .ZN(n6383) );
  XNOR2_X1 U4935 ( .A(n8296), .B(n8297), .ZN(n6267) );
  NAND2_X1 U4936 ( .A1(n4744), .A2(n4748), .ZN(n8041) );
  NAND2_X1 U4937 ( .A1(n4944), .A2(n4945), .ZN(n8552) );
  OR2_X1 U4938 ( .A1(n6267), .A2(SI_29_), .ZN(n6268) );
  XNOR2_X1 U4939 ( .A(n5672), .B(n5671), .ZN(n7646) );
  AND4_X1 U4941 ( .A1(n5068), .A2(n5054), .A3(n5053), .A4(n5052), .ZN(n4409)
         );
  INV_X1 U4942 ( .A(n5951), .ZN(n4410) );
  OAI21_X2 U4943 ( .B1(n5133), .B2(n5134), .A(n5132), .ZN(n4877) );
  NOR2_X2 U4945 ( .A1(n7859), .A2(n10011), .ZN(n7858) );
  NOR2_X4 U4946 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5934) );
  INV_X4 U4948 ( .A(n4410), .ZN(n4411) );
  AOI21_X1 U4950 ( .B1(n4428), .B2(n6487), .A(n4510), .ZN(n4674) );
  NOR2_X1 U4951 ( .A1(n4538), .A2(n4462), .ZN(n8314) );
  INV_X1 U4952 ( .A(n10028), .ZN(n9720) );
  NAND2_X1 U4953 ( .A1(n9817), .A2(n4616), .ZN(n9799) );
  NAND2_X1 U4954 ( .A1(n8300), .A2(n8299), .ZN(n8323) );
  NAND2_X1 U4955 ( .A1(n9277), .A2(n5625), .ZN(n9215) );
  NAND2_X1 U4956 ( .A1(n6267), .A2(SI_29_), .ZN(n8300) );
  NAND2_X1 U4957 ( .A1(n6243), .A2(n6242), .ZN(n9103) );
  NAND2_X1 U4958 ( .A1(n4758), .A2(n7961), .ZN(n7948) );
  AOI21_X1 U4959 ( .B1(n4733), .B2(n4731), .A(n4477), .ZN(n4730) );
  INV_X1 U4960 ( .A(n4733), .ZN(n4732) );
  NAND2_X1 U4961 ( .A1(n5755), .A2(n5754), .ZN(n9781) );
  NAND2_X1 U4962 ( .A1(n5734), .A2(n5733), .ZN(n9792) );
  NAND2_X1 U4963 ( .A1(n6204), .A2(n6203), .ZN(n9119) );
  OAI21_X1 U4964 ( .B1(n7342), .B2(n4628), .A(n4629), .ZN(n7630) );
  NAND2_X1 U4965 ( .A1(n7758), .A2(n4931), .ZN(n7805) );
  NAND2_X1 U4966 ( .A1(n4841), .A2(n4840), .ZN(n7342) );
  OR2_X1 U4967 ( .A1(n5630), .A2(n5631), .ZN(n5650) );
  AND2_X1 U4968 ( .A1(n7610), .A2(n4448), .ZN(n4765) );
  OAI21_X1 U4969 ( .B1(n5400), .B2(n5399), .A(n5398), .ZN(n5427) );
  INV_X2 U4970 ( .A(n9916), .ZN(n4415) );
  NAND3_X1 U4971 ( .A1(n5118), .A2(n5117), .A3(n5116), .ZN(n9647) );
  INV_X1 U4972 ( .A(n8398), .ZN(n6284) );
  NAND3_X1 U4973 ( .A1(n4613), .A2(n5130), .A3(n5131), .ZN(n9645) );
  NAND4_X2 U4974 ( .A1(n5975), .A2(n5974), .A3(n5973), .A4(n5972), .ZN(n8398)
         );
  CLKBUF_X1 U4975 ( .A(n5322), .Z(n5817) );
  AND4_X1 U4976 ( .A1(n5944), .A2(n5943), .A3(n5942), .A4(n5941), .ZN(n6280)
         );
  AND2_X1 U4977 ( .A1(n5196), .A2(n5195), .ZN(n7331) );
  AND3_X1 U4978 ( .A1(n5969), .A2(n5968), .A3(n5967), .ZN(n10331) );
  AND3_X1 U4980 ( .A1(n5939), .A2(n4641), .A3(n5938), .ZN(n7137) );
  AOI21_X1 U4981 ( .B1(n4881), .B2(n4886), .A(n4472), .ZN(n4879) );
  NAND2_X1 U4982 ( .A1(n4999), .A2(n4997), .ZN(n10079) );
  INV_X2 U4983 ( .A(n6004), .ZN(n5962) );
  NAND2_X2 U4984 ( .A1(n5920), .A2(n8022), .ZN(n5971) );
  AND2_X1 U4985 ( .A1(n4883), .A2(n4500), .ZN(n4881) );
  NAND2_X1 U4986 ( .A1(n10075), .A2(n4998), .ZN(n4997) );
  XNOR2_X1 U4987 ( .A(n6323), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8165) );
  XNOR2_X1 U4988 ( .A(n5060), .B(P1_IR_REG_29__SCAN_IN), .ZN(n10083) );
  INV_X1 U4989 ( .A(n8509), .ZN(n8533) );
  NAND2_X1 U4990 ( .A1(n9164), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5918) );
  XNOR2_X1 U4991 ( .A(n6164), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8509) );
  NAND2_X1 U4992 ( .A1(n5092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5060) );
  XNOR2_X1 U4993 ( .A(n6321), .B(n6320), .ZN(n8329) );
  XNOR2_X1 U4994 ( .A(n5094), .B(n5056), .ZN(n6554) );
  AND3_X1 U4995 ( .A1(n4694), .A2(n4950), .A3(n4693), .ZN(n5911) );
  AND2_X1 U4996 ( .A1(n4422), .A2(n5909), .ZN(n4950) );
  NOR2_X1 U4997 ( .A1(n5049), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4800) );
  AND2_X1 U4998 ( .A1(n5141), .A2(n5051), .ZN(n5184) );
  AND4_X1 U4999 ( .A1(n5896), .A2(n5895), .A3(n8937), .A4(n5982), .ZN(n5898)
         );
  INV_X1 U5000 ( .A(n5965), .ZN(n4416) );
  NAND2_X1 U5001 ( .A1(n4905), .A2(n4908), .ZN(n4910) );
  AND2_X1 U5002 ( .A1(n5906), .A2(n5907), .ZN(n4951) );
  NAND2_X1 U5003 ( .A1(n4906), .A2(n4907), .ZN(n4911) );
  INV_X1 U5004 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5540) );
  NOR2_X1 U5005 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5896) );
  NOR2_X1 U5006 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5895) );
  INV_X1 U5007 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n8937) );
  INV_X4 U5008 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X4 U5009 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U5010 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5051) );
  INV_X1 U5011 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5561) );
  INV_X1 U5012 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5074) );
  NOR2_X1 U5013 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5141) );
  INV_X1 U5014 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6128) );
  NOR2_X1 U5015 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5900) );
  NOR2_X1 U5016 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5901) );
  NOR2_X2 U5017 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_RD_REG_SCAN_IN), .ZN(
        n4906) );
  INV_X1 U5018 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4907) );
  AND2_X1 U5019 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n4905) );
  INV_X1 U5020 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4908) );
  INV_X1 U5021 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6320) );
  XNOR2_X2 U5022 ( .A(n5846), .B(P1_IR_REG_22__SCAN_IN), .ZN(n5851) );
  OAI21_X2 U5023 ( .B1(n8033), .B2(n8386), .A(n7999), .ZN(n8078) );
  BUF_X4 U5024 ( .A(n5963), .Z(n6241) );
  NAND2_X1 U5025 ( .A1(n6897), .A2(n6896), .ZN(n4417) );
  BUF_X4 U5026 ( .A(n6902), .Z(n8011) );
  OAI21_X2 U5027 ( .B1(n6346), .B2(n6352), .A(n6369), .ZN(n6351) );
  AOI22_X4 U5028 ( .A1(n8041), .A2(n8040), .B1(n8677), .B2(n7991), .ZN(n8087)
         );
  NAND2_X2 U5029 ( .A1(n9858), .A2(n4423), .ZN(n9808) );
  INV_X1 U5030 ( .A(n6004), .ZN(n4418) );
  NAND2_X1 U5032 ( .A1(n4768), .A2(n9424), .ZN(n9427) );
  NOR2_X1 U5033 ( .A1(n5483), .A2(n4901), .ZN(n4900) );
  AND2_X1 U5034 ( .A1(n5904), .A2(n6128), .ZN(n5905) );
  INV_X1 U5035 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5904) );
  OR2_X1 U5036 ( .A1(n9911), .A2(n9259), .ZN(n9497) );
  NAND2_X1 U5037 ( .A1(n5301), .A2(n5300), .ZN(n5326) );
  AND2_X1 U5038 ( .A1(n6240), .A2(n6239), .ZN(n8590) );
  AOI21_X1 U5039 ( .B1(n9793), .B2(n5171), .A(n5740), .ZN(n9269) );
  NAND2_X1 U5040 ( .A1(n9919), .A2(n6403), .ZN(n5025) );
  NAND2_X1 U5041 ( .A1(n4790), .A2(n4792), .ZN(n4788) );
  NAND2_X1 U5042 ( .A1(n9467), .A2(n9466), .ZN(n4777) );
  OAI21_X1 U5043 ( .B1(n4547), .B2(n4546), .A(n8234), .ZN(n8237) );
  OAI21_X1 U5044 ( .B1(n8229), .B2(n8285), .A(n8231), .ZN(n4546) );
  NOR2_X1 U5045 ( .A1(n8230), .A2(n8312), .ZN(n4547) );
  AOI21_X1 U5046 ( .B1(n9493), .B2(n4802), .A(n4478), .ZN(n4803) );
  NOR2_X1 U5047 ( .A1(n4804), .A2(n4806), .ZN(n4802) );
  AND2_X1 U5048 ( .A1(n4834), .A2(n4832), .ZN(n4831) );
  NAND2_X1 U5049 ( .A1(n9527), .A2(n9526), .ZN(n4832) );
  AND2_X1 U5050 ( .A1(n4494), .A2(n4835), .ZN(n4834) );
  INV_X1 U5051 ( .A(n4837), .ZN(n4828) );
  INV_X1 U5052 ( .A(n4494), .ZN(n4827) );
  AOI21_X1 U5053 ( .B1(n4826), .B2(n4829), .A(n9534), .ZN(n4825) );
  INV_X1 U5054 ( .A(n4830), .ZN(n4829) );
  NAND2_X1 U5055 ( .A1(n4786), .A2(n4782), .ZN(n9516) );
  OAI21_X1 U5056 ( .B1(n4787), .B2(n9511), .A(n9533), .ZN(n4786) );
  NOR2_X1 U5057 ( .A1(n6222), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6233) );
  INV_X1 U5058 ( .A(n4914), .ZN(n4913) );
  OAI21_X1 U5059 ( .B1(n4921), .B2(n4915), .A(n4919), .ZN(n4914) );
  AND2_X1 U5060 ( .A1(n4888), .A2(n5033), .ZN(n4887) );
  NAND2_X1 U5061 ( .A1(n7987), .A2(n8675), .ZN(n4757) );
  INV_X1 U5062 ( .A(n7983), .ZN(n4756) );
  NOR2_X1 U5063 ( .A1(n4683), .A2(n8587), .ZN(n4682) );
  INV_X1 U5064 ( .A(n4684), .ZN(n4683) );
  OR2_X1 U5065 ( .A1(n8052), .A2(n8624), .ZN(n8155) );
  OR2_X1 U5066 ( .A1(n8683), .A2(n8663), .ZN(n8263) );
  OR2_X1 U5067 ( .A1(n9152), .A2(n8074), .ZN(n8254) );
  NAND2_X1 U5068 ( .A1(n8177), .A2(n8178), .ZN(n8171) );
  AND2_X1 U5069 ( .A1(n9168), .A2(n5921), .ZN(n5970) );
  OR2_X1 U5070 ( .A1(n9103), .A2(n8577), .ZN(n8149) );
  OR2_X1 U5071 ( .A1(n8761), .A2(n8604), .ZN(n8289) );
  INV_X1 U5072 ( .A(n6308), .ZN(n4672) );
  NAND2_X1 U5073 ( .A1(n5928), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6345) );
  AND2_X1 U5074 ( .A1(n5910), .A2(n5905), .ZN(n4696) );
  INV_X1 U5075 ( .A(n5903), .ZN(n4695) );
  NAND2_X1 U5076 ( .A1(n4603), .A2(n6421), .ZN(n5202) );
  AND2_X1 U5077 ( .A1(n6500), .A2(n9613), .ZN(n4603) );
  INV_X1 U5078 ( .A(n5531), .ZN(n4599) );
  INV_X1 U5079 ( .A(n6411), .ZN(n5013) );
  AND2_X1 U5080 ( .A1(n5019), .A2(n4482), .ZN(n5017) );
  NOR2_X1 U5081 ( .A1(n9827), .A2(n4726), .ZN(n4725) );
  INV_X1 U5082 ( .A(n4727), .ZN(n4726) );
  OR2_X1 U5083 ( .A1(n10003), .A2(n7854), .ZN(n9495) );
  INV_X1 U5084 ( .A(n4632), .ZN(n4631) );
  INV_X1 U5085 ( .A(n6390), .ZN(n5003) );
  AND2_X1 U5086 ( .A1(n9595), .A2(n9608), .ZN(n6460) );
  INV_X1 U5087 ( .A(n5050), .ZN(n4799) );
  NAND2_X1 U5088 ( .A1(n4799), .A2(n4800), .ZN(n4556) );
  AND2_X1 U5089 ( .A1(n5673), .A2(n5656), .ZN(n5671) );
  NAND2_X1 U5090 ( .A1(n4893), .A2(n4891), .ZN(n5558) );
  AOI21_X1 U5091 ( .B1(n4899), .B2(n4894), .A(n4892), .ZN(n4891) );
  INV_X1 U5092 ( .A(n5533), .ZN(n4892) );
  INV_X1 U5093 ( .A(SI_14_), .ZN(n5453) );
  AOI21_X1 U5094 ( .B1(n4887), .B2(n4885), .A(n4884), .ZN(n4883) );
  INV_X1 U5095 ( .A(n5324), .ZN(n4885) );
  INV_X1 U5096 ( .A(n5352), .ZN(n4884) );
  NAND2_X1 U5097 ( .A1(n4838), .A2(n5270), .ZN(n5297) );
  INV_X1 U5098 ( .A(n5190), .ZN(n5191) );
  NAND2_X1 U5099 ( .A1(n7992), .A2(n8662), .ZN(n4740) );
  NAND2_X1 U5100 ( .A1(n4938), .A2(n4937), .ZN(n4936) );
  AND2_X1 U5101 ( .A1(n5921), .A2(n5920), .ZN(n5994) );
  AND2_X1 U5102 ( .A1(n8022), .A2(n9168), .ZN(n5951) );
  NOR2_X1 U5103 ( .A1(n5984), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U5104 ( .A(n7048), .B(n6799), .ZN(n6786) );
  OR2_X1 U5105 ( .A1(n8402), .A2(n4867), .ZN(n4526) );
  NAND2_X1 U5106 ( .A1(n4870), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4867) );
  NAND2_X1 U5107 ( .A1(n8426), .A2(n4870), .ZN(n4866) );
  OR2_X1 U5108 ( .A1(n8456), .A2(n8455), .ZN(n8491) );
  XNOR2_X1 U5109 ( .A(n8506), .B(n8527), .ZN(n10291) );
  AOI21_X1 U5110 ( .B1(n4647), .B2(n4645), .A(n4461), .ZN(n4644) );
  AOI21_X1 U5111 ( .B1(n7686), .B2(n8209), .A(n6039), .ZN(n7759) );
  AND2_X1 U5112 ( .A1(n8208), .A2(n8214), .ZN(n8353) );
  NAND2_X1 U5113 ( .A1(n7759), .A2(n8353), .ZN(n7758) );
  NAND2_X1 U5114 ( .A1(n7473), .A2(n8344), .ZN(n4927) );
  NAND2_X1 U5115 ( .A1(n7022), .A2(n10324), .ZN(n8177) );
  OAI22_X1 U5116 ( .A1(n8575), .A2(n6315), .B1(n8590), .B2(n9110), .ZN(n8567)
         );
  OR2_X1 U5117 ( .A1(n8129), .A2(n8590), .ZN(n8293) );
  OAI22_X1 U5118 ( .A1(n8621), .A2(n8626), .B1(n8614), .B2(n8627), .ZN(n8612)
         );
  OR2_X1 U5119 ( .A1(n8627), .A2(n8635), .ZN(n8156) );
  NAND2_X1 U5120 ( .A1(n5238), .A2(n5264), .ZN(n4985) );
  NOR2_X1 U5121 ( .A1(n9328), .A2(n4983), .ZN(n4982) );
  NAND2_X1 U5122 ( .A1(n4967), .A2(n4421), .ZN(n4586) );
  NAND2_X1 U5123 ( .A1(n7300), .A2(n9605), .ZN(n9608) );
  NAND2_X1 U5124 ( .A1(n5081), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5846) );
  AND2_X1 U5125 ( .A1(n5641), .A2(n5640), .ZN(n9370) );
  AND3_X1 U5126 ( .A1(n5571), .A2(n5570), .A3(n5569), .ZN(n9259) );
  NAND2_X1 U5127 ( .A1(n5086), .A2(n5824), .ZN(n6500) );
  AND2_X1 U5128 ( .A1(n5080), .A2(n4430), .ZN(n5086) );
  AND2_X1 U5129 ( .A1(n7725), .A2(n7868), .ZN(n5080) );
  NAND2_X1 U5130 ( .A1(n4615), .A2(n9517), .ZN(n9767) );
  NAND2_X1 U5131 ( .A1(n9799), .A2(n4454), .ZN(n4615) );
  NAND2_X1 U5132 ( .A1(n9827), .A2(n9512), .ZN(n9801) );
  OAI21_X1 U5133 ( .B1(n4568), .B2(n4571), .A(n4569), .ZN(n9807) );
  NAND2_X1 U5134 ( .A1(n4572), .A2(n4432), .ZN(n4571) );
  AOI21_X1 U5135 ( .B1(n4572), .B2(n4455), .A(n4570), .ZN(n4569) );
  NOR2_X1 U5136 ( .A1(n9827), .A2(n9625), .ZN(n4570) );
  AOI21_X1 U5137 ( .B1(n4561), .B2(n4559), .A(n4508), .ZN(n4558) );
  INV_X1 U5138 ( .A(n4561), .ZN(n4560) );
  NAND2_X1 U5139 ( .A1(n6960), .A2(n6425), .ZN(n9425) );
  AND2_X1 U5140 ( .A1(n9529), .A2(n9588), .ZN(n9576) );
  NAND2_X1 U5141 ( .A1(n9767), .A2(n9768), .ZN(n9766) );
  NAND2_X1 U5142 ( .A1(n5612), .A2(n5611), .ZN(n9878) );
  NAND2_X1 U5143 ( .A1(n4995), .A2(P1_IR_REG_30__SCAN_IN), .ZN(n4999) );
  NAND2_X1 U5144 ( .A1(n10075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4995) );
  INV_X1 U5145 ( .A(n5087), .ZN(n5057) );
  NAND2_X1 U5146 ( .A1(n5541), .A2(n5540), .ZN(n5073) );
  NAND2_X1 U5147 ( .A1(n6418), .A2(n6417), .ZN(n6452) );
  INV_X1 U5148 ( .A(n9444), .ZN(n4796) );
  AOI21_X1 U5149 ( .B1(n4791), .B2(n4793), .A(n9441), .ZN(n4790) );
  NAND2_X1 U5150 ( .A1(n4541), .A2(n8223), .ZN(n8224) );
  NAND2_X1 U5151 ( .A1(n8228), .A2(n8222), .ZN(n4541) );
  NAND2_X1 U5152 ( .A1(n9468), .A2(n9534), .ZN(n4775) );
  NAND2_X1 U5153 ( .A1(n4777), .A2(n9533), .ZN(n4776) );
  OAI21_X1 U5154 ( .B1(n8237), .B2(n8713), .A(n8236), .ZN(n8238) );
  NAND2_X1 U5155 ( .A1(n4774), .A2(n4772), .ZN(n9491) );
  NOR2_X1 U5156 ( .A1(n6436), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U5157 ( .A1(n9485), .A2(n9396), .ZN(n4774) );
  INV_X1 U5158 ( .A(n9487), .ZN(n4773) );
  INV_X1 U5159 ( .A(n4804), .ZN(n4801) );
  NOR2_X1 U5160 ( .A1(n9500), .A2(n4803), .ZN(n9501) );
  INV_X1 U5161 ( .A(n9506), .ZN(n4785) );
  OAI21_X1 U5162 ( .B1(n4545), .B2(n8278), .A(n4544), .ZN(n8284) );
  AOI22_X1 U5163 ( .A1(n8273), .A2(n8274), .B1(n8275), .B2(n6332), .ZN(n4545)
         );
  NAND2_X1 U5164 ( .A1(n4831), .A2(n4833), .ZN(n4824) );
  OR2_X1 U5165 ( .A1(n4836), .A2(n9524), .ZN(n4833) );
  AND2_X1 U5166 ( .A1(n9455), .A2(n9443), .ZN(n9447) );
  NAND2_X1 U5167 ( .A1(n8566), .A2(n8295), .ZN(n4539) );
  NAND2_X1 U5168 ( .A1(n5940), .A2(n10319), .ZN(n8176) );
  AOI21_X1 U5169 ( .B1(n4817), .B2(n4424), .A(n10024), .ZN(n4813) );
  NOR2_X1 U5170 ( .A1(n9536), .A2(n4816), .ZN(n4815) );
  OAI21_X1 U5171 ( .B1(n10028), .B2(n9533), .A(n9591), .ZN(n4816) );
  AOI21_X1 U5172 ( .B1(n5626), .B2(n4920), .A(n4511), .ZN(n4919) );
  INV_X1 U5173 ( .A(n5607), .ZN(n4920) );
  INV_X1 U5174 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5044) );
  NAND2_X1 U5175 ( .A1(n7561), .A2(n5038), .ZN(n7831) );
  INV_X1 U5176 ( .A(n7714), .ZN(n4980) );
  NAND2_X1 U5177 ( .A1(n4813), .A2(n4814), .ZN(n4812) );
  INV_X1 U5178 ( .A(n4817), .ZN(n4814) );
  OAI211_X1 U5179 ( .C1(n4819), .C2(n9523), .A(n4820), .B(n4475), .ZN(n9531)
         );
  INV_X1 U5180 ( .A(n4825), .ZN(n4819) );
  NOR2_X1 U5181 ( .A1(n4809), .A2(n10028), .ZN(n4808) );
  INV_X1 U5182 ( .A(n4815), .ZN(n4809) );
  AND2_X1 U5183 ( .A1(n9875), .A2(n9475), .ZN(n4640) );
  NAND2_X1 U5184 ( .A1(n7268), .A2(n6429), .ZN(n9390) );
  OAI211_X1 U5185 ( .C1(n4910), .C2(P2_DATAO_REG_2__SCAN_IN), .A(n4548), .B(
        n4549), .ZN(n5137) );
  NAND2_X1 U5186 ( .A1(n8370), .A2(n9088), .ZN(n4938) );
  XNOR2_X1 U5187 ( .A(n6711), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n10226) );
  NAND2_X1 U5188 ( .A1(n6785), .A2(n6784), .ZN(n7048) );
  NOR2_X1 U5189 ( .A1(n10243), .A2(n4875), .ZN(n7031) );
  NOR2_X1 U5190 ( .A1(n10254), .A2(n10376), .ZN(n4875) );
  NAND2_X1 U5191 ( .A1(n7194), .A2(n5041), .ZN(n7195) );
  XNOR2_X1 U5192 ( .A(n7831), .B(n7562), .ZN(n7563) );
  NOR2_X1 U5193 ( .A1(n8405), .A2(n8404), .ZN(n8437) );
  NOR2_X1 U5194 ( .A1(n7834), .A2(n9037), .ZN(n8404) );
  AND2_X1 U5195 ( .A1(n8512), .A2(n8511), .ZN(n8513) );
  AND2_X1 U5196 ( .A1(n6245), .A2(n6244), .ZN(n6254) );
  OAI21_X1 U5197 ( .B1(n8587), .B2(n4435), .A(n4687), .ZN(n4686) );
  OR2_X1 U5198 ( .A1(n8761), .A2(n8385), .ZN(n4687) );
  AND2_X1 U5199 ( .A1(n6143), .A2(n6142), .ZN(n6155) );
  NOR2_X1 U5200 ( .A1(n6119), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6143) );
  NOR2_X1 U5201 ( .A1(n6290), .A2(n4652), .ZN(n4660) );
  INV_X1 U5202 ( .A(n8329), .ZN(n6478) );
  AND2_X1 U5203 ( .A1(n6353), .A2(n6588), .ZN(n6477) );
  CLKBUF_X1 U5204 ( .A(n6893), .Z(n6349) );
  INV_X1 U5205 ( .A(n4948), .ZN(n4947) );
  OAI21_X1 U5206 ( .B1(n8578), .B2(n4949), .A(n8147), .ZN(n4948) );
  OR2_X1 U5207 ( .A1(n8083), .A2(n8591), .ZN(n8364) );
  AND2_X1 U5208 ( .A1(n8669), .A2(n8649), .ZN(n4673) );
  OR2_X1 U5209 ( .A1(n9133), .A2(n8662), .ZN(n8154) );
  INV_X1 U5210 ( .A(n6310), .ZN(n4668) );
  NAND2_X1 U5211 ( .A1(n6309), .A2(n4670), .ZN(n4669) );
  OR2_X1 U5212 ( .A1(n7980), .A2(n7981), .ZN(n8248) );
  NAND2_X1 U5213 ( .A1(n4651), .A2(n4649), .ZN(n7930) );
  NOR2_X1 U5214 ( .A1(n4450), .A2(n4650), .ZN(n4649) );
  INV_X1 U5215 ( .A(n6303), .ZN(n4650) );
  OR2_X1 U5216 ( .A1(n8112), .A2(n7922), .ZN(n8225) );
  OR2_X1 U5217 ( .A1(n7969), .A2(n8104), .ZN(n8232) );
  INV_X1 U5218 ( .A(n5905), .ZN(n4692) );
  NOR3_X1 U5219 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U5220 ( .A1(n6339), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  INV_X1 U5221 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5982) );
  NAND2_X1 U5222 ( .A1(n6099), .A2(n5897), .ZN(n5956) );
  OAI211_X1 U5223 ( .C1(n5169), .C2(n4956), .A(n4955), .B(n4953), .ZN(n5108)
         );
  NAND2_X1 U5224 ( .A1(n5169), .A2(n4954), .ZN(n4953) );
  OR2_X1 U5225 ( .A1(n9759), .A2(n6413), .ZN(n9528) );
  NOR2_X1 U5226 ( .A1(n9759), .A2(n9781), .ZN(n4721) );
  NAND2_X1 U5227 ( .A1(n9781), .A2(n9236), .ZN(n9518) );
  INV_X1 U5228 ( .A(n5017), .ZN(n5016) );
  INV_X1 U5229 ( .A(n4640), .ZN(n4635) );
  NOR2_X1 U5230 ( .A1(n9842), .A2(n9861), .ZN(n4727) );
  NOR2_X1 U5231 ( .A1(n6440), .A2(n4638), .ZN(n4637) );
  INV_X1 U5232 ( .A(n9856), .ZN(n4638) );
  INV_X1 U5233 ( .A(n9632), .ZN(n9258) );
  NOR2_X1 U5234 ( .A1(n6401), .A2(n4567), .ZN(n4566) );
  INV_X1 U5235 ( .A(n6399), .ZN(n4567) );
  NOR2_X1 U5236 ( .A1(n9229), .A2(n10187), .ZN(n4722) );
  NAND2_X1 U5237 ( .A1(n9390), .A2(n9388), .ZN(n7340) );
  OR2_X1 U5238 ( .A1(n7459), .A2(n7344), .ZN(n9455) );
  AND2_X1 U5239 ( .A1(n7264), .A2(n9442), .ZN(n7268) );
  INV_X1 U5240 ( .A(n9425), .ZN(n4770) );
  NAND2_X1 U5241 ( .A1(n7148), .A2(n6392), .ZN(n7261) );
  INV_X1 U5242 ( .A(n4993), .ZN(n4992) );
  OAI21_X1 U5243 ( .B1(n9444), .B2(n4994), .A(n7283), .ZN(n4993) );
  INV_X1 U5244 ( .A(n6393), .ZN(n4994) );
  NAND2_X1 U5245 ( .A1(n7261), .A2(n9444), .ZN(n7260) );
  AND2_X1 U5246 ( .A1(n4797), .A2(n9442), .ZN(n9548) );
  NAND2_X1 U5247 ( .A1(n6266), .A2(n6265), .ZN(n8296) );
  INV_X1 U5248 ( .A(n5723), .ZN(n5724) );
  AND2_X1 U5249 ( .A1(n5748), .A2(n5732), .ZN(n5746) );
  AND3_X1 U5250 ( .A1(n5561), .A2(n5540), .A3(n5074), .ZN(n5068) );
  OR2_X1 U5251 ( .A1(n5486), .A2(n9019), .ZN(n4896) );
  NOR2_X1 U5252 ( .A1(n5050), .A2(n5049), .ZN(n5027) );
  NAND2_X2 U5253 ( .A1(n4911), .A2(n4910), .ZN(n5153) );
  NAND2_X1 U5254 ( .A1(n8122), .A2(n8123), .ZN(n4743) );
  INV_X1 U5255 ( .A(n8109), .ZN(n4762) );
  NAND2_X1 U5256 ( .A1(n7917), .A2(n8391), .ZN(n4761) );
  OR2_X1 U5257 ( .A1(n4737), .A2(n7994), .ZN(n4736) );
  AOI21_X1 U5258 ( .B1(n8086), .B2(n4740), .A(n4738), .ZN(n4737) );
  INV_X1 U5259 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5906) );
  OR2_X1 U5260 ( .A1(n6711), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U5261 ( .A1(n6793), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7029) );
  NAND2_X1 U5262 ( .A1(n6786), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7050) );
  AND2_X1 U5263 ( .A1(n7030), .A2(n4876), .ZN(n10243) );
  INV_X1 U5264 ( .A(n10244), .ZN(n4876) );
  XNOR2_X1 U5265 ( .A(n7031), .B(n10269), .ZN(n10266) );
  AND2_X1 U5266 ( .A1(n6347), .A2(n6369), .ZN(n6370) );
  AND3_X1 U5267 ( .A1(n4526), .A2(n4521), .A3(n4866), .ZN(n8472) );
  NAND2_X1 U5268 ( .A1(n8491), .A2(n5037), .ZN(n8495) );
  NAND2_X1 U5269 ( .A1(n8477), .A2(n8476), .ZN(n8505) );
  OAI21_X1 U5270 ( .B1(n10288), .B2(n4701), .A(n4700), .ZN(n10097) );
  NAND2_X1 U5271 ( .A1(n4702), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U5272 ( .A1(n8514), .A2(n4702), .ZN(n4700) );
  INV_X1 U5273 ( .A(n10098), .ZN(n4702) );
  AOI21_X1 U5274 ( .B1(n8535), .B2(n10298), .A(n8534), .ZN(n8536) );
  AOI21_X1 U5275 ( .B1(n10096), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n4523), .ZN(
        n4714) );
  AOI21_X1 U5276 ( .B1(n8552), .B2(n8553), .A(n6262), .ZN(n8335) );
  AND2_X1 U5277 ( .A1(n8293), .A2(n8294), .ZN(n8578) );
  NOR2_X1 U5278 ( .A1(n4690), .A2(n4426), .ZN(n4684) );
  AND2_X1 U5279 ( .A1(n6228), .A2(n6227), .ZN(n8604) );
  AND3_X1 U5280 ( .A1(n6192), .A2(n6191), .A3(n6190), .ZN(n8624) );
  AND2_X1 U5281 ( .A1(n8156), .A2(n8276), .ZN(n8626) );
  AND3_X1 U5282 ( .A1(n6202), .A2(n6201), .A3(n6200), .ZN(n8635) );
  AOI21_X1 U5283 ( .B1(n6163), .B2(n8696), .A(n4929), .ZN(n4928) );
  INV_X1 U5284 ( .A(n8263), .ZN(n4929) );
  INV_X1 U5285 ( .A(n8361), .ZN(n8657) );
  OR2_X1 U5286 ( .A1(n6057), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6067) );
  NAND2_X1 U5287 ( .A1(n6047), .A2(n6046), .ZN(n6057) );
  INV_X1 U5288 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6046) );
  OAI21_X1 U5289 ( .B1(n4661), .B2(n4657), .A(n4654), .ZN(n7592) );
  INV_X1 U5290 ( .A(n4658), .ZN(n4657) );
  AOI21_X1 U5291 ( .B1(n4658), .B2(n4656), .A(n4655), .ZN(n4654) );
  NOR2_X1 U5292 ( .A1(n6291), .A2(n4659), .ZN(n4658) );
  NAND2_X1 U5293 ( .A1(n6003), .A2(n8198), .ZN(n7473) );
  AND2_X1 U5294 ( .A1(n8203), .A2(n8193), .ZN(n8344) );
  NAND2_X1 U5295 ( .A1(n4653), .A2(n6289), .ZN(n7477) );
  NAND2_X1 U5296 ( .A1(n4661), .A2(n4660), .ZN(n4653) );
  AND4_X1 U5297 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n7614)
         );
  NAND2_X1 U5298 ( .A1(n6284), .A2(n7257), .ZN(n8186) );
  INV_X1 U5299 ( .A(n8184), .ZN(n8341) );
  OR2_X1 U5300 ( .A1(n5946), .A2(n5959), .ZN(n5031) );
  AOI22_X1 U5301 ( .A1(n8567), .A2(n6316), .B1(n8557), .B2(n9103), .ZN(n8555)
         );
  INV_X1 U5302 ( .A(n8553), .ZN(n8554) );
  XNOR2_X1 U5303 ( .A(n9097), .B(n8569), .ZN(n8553) );
  AND2_X1 U5304 ( .A1(n8149), .A2(n8147), .ZN(n8566) );
  NAND2_X1 U5305 ( .A1(n8625), .A2(n8626), .ZN(n4926) );
  OR2_X1 U5306 ( .A1(n6888), .A2(n8312), .ZN(n8676) );
  INV_X1 U5307 ( .A(n8717), .ZN(n8678) );
  AND2_X1 U5308 ( .A1(n6888), .A2(n8285), .ZN(n8717) );
  NAND2_X1 U5309 ( .A1(n8336), .A2(n6479), .ZN(n8722) );
  NOR2_X1 U5310 ( .A1(n4932), .A2(n8195), .ZN(n4931) );
  AND3_X1 U5311 ( .A1(n5989), .A2(n5988), .A3(n5987), .ZN(n10337) );
  OR2_X1 U5312 ( .A1(n8165), .A2(n8379), .ZN(n10359) );
  INV_X1 U5313 ( .A(n8722), .ZN(n8673) );
  AND2_X1 U5314 ( .A1(n5368), .A2(n5369), .ZN(n9196) );
  NAND2_X1 U5315 ( .A1(n7434), .A2(n5295), .ZN(n5323) );
  NAND2_X1 U5316 ( .A1(n4611), .A2(n9309), .ZN(n4610) );
  INV_X1 U5317 ( .A(n9307), .ZN(n4611) );
  OR2_X1 U5318 ( .A1(n5516), .A2(n5497), .ZN(n5545) );
  AND2_X1 U5319 ( .A1(n4599), .A2(n5481), .ZN(n4597) );
  NAND2_X1 U5320 ( .A1(n4479), .A2(n4599), .ZN(n4596) );
  OAI21_X1 U5321 ( .B1(n9186), .B2(n9266), .A(n9265), .ZN(n9264) );
  AND2_X1 U5322 ( .A1(n5323), .A2(n4498), .ZN(n7783) );
  OR2_X1 U5323 ( .A1(n5412), .A2(n5411), .ZN(n5436) );
  INV_X1 U5324 ( .A(n4610), .ZN(n4608) );
  NAND2_X1 U5325 ( .A1(n5369), .A2(n9309), .ZN(n4605) );
  NAND2_X1 U5326 ( .A1(n9196), .A2(n9197), .ZN(n9195) );
  NAND2_X1 U5327 ( .A1(n5668), .A2(n4582), .ZN(n4957) );
  AND2_X1 U5328 ( .A1(n5687), .A2(n5686), .ZN(n9512) );
  AND4_X1 U5329 ( .A1(n5318), .A2(n5317), .A3(n5316), .A4(n5315), .ZN(n7452)
         );
  AND4_X1 U5330 ( .A1(n5230), .A2(n5229), .A3(n5228), .A4(n5227), .ZN(n7153)
         );
  NAND2_X1 U5331 ( .A1(n5005), .A2(n4458), .ZN(n9739) );
  AOI21_X1 U5332 ( .B1(n5007), .B2(n5012), .A(n4459), .ZN(n5006) );
  AOI21_X1 U5333 ( .B1(n5011), .B2(n4420), .A(n4464), .ZN(n5010) );
  AND2_X1 U5334 ( .A1(n9784), .A2(n9514), .ZN(n9800) );
  OR2_X1 U5335 ( .A1(n5016), .A2(n4576), .ZN(n4575) );
  INV_X1 U5336 ( .A(n6407), .ZN(n4576) );
  INV_X1 U5337 ( .A(n4573), .ZN(n4572) );
  OAI21_X1 U5338 ( .B1(n5016), .B2(n4574), .A(n5014), .ZN(n4573) );
  NAND2_X1 U5339 ( .A1(n4436), .A2(n6407), .ZN(n4574) );
  AOI21_X1 U5340 ( .B1(n5017), .B2(n5015), .A(n4469), .ZN(n5014) );
  NAND2_X1 U5341 ( .A1(n9858), .A2(n4725), .ZN(n9825) );
  AND2_X1 U5342 ( .A1(n5020), .A2(n6410), .ZN(n5019) );
  OR2_X1 U5343 ( .A1(n6409), .A2(n5021), .ZN(n5020) );
  NAND2_X1 U5344 ( .A1(n4437), .A2(n6408), .ZN(n5021) );
  INV_X1 U5345 ( .A(n6408), .ZN(n5022) );
  AND2_X1 U5346 ( .A1(n9365), .A2(n9372), .ZN(n9840) );
  OAI21_X1 U5347 ( .B1(n4568), .B2(n4436), .A(n6407), .ZN(n9874) );
  NAND2_X1 U5348 ( .A1(n6439), .A2(n9497), .ZN(n9893) );
  NOR2_X1 U5349 ( .A1(n9920), .A2(n9911), .ZN(n9910) );
  NAND2_X1 U5350 ( .A1(n9910), .A2(n9892), .ZN(n9886) );
  NAND2_X1 U5351 ( .A1(n5025), .A2(n5023), .ZN(n6406) );
  NOR2_X1 U5352 ( .A1(n5024), .A2(n4512), .ZN(n5023) );
  AND2_X1 U5353 ( .A1(n9497), .A2(n9481), .ZN(n9904) );
  NAND2_X1 U5354 ( .A1(n6400), .A2(n6399), .ZN(n4565) );
  NAND2_X1 U5355 ( .A1(n7696), .A2(n4566), .ZN(n4562) );
  NAND2_X1 U5356 ( .A1(n7852), .A2(n9563), .ZN(n7851) );
  AOI21_X1 U5357 ( .B1(n6434), .B2(n4631), .A(n4630), .ZN(n4629) );
  NAND2_X1 U5358 ( .A1(n7342), .A2(n4632), .ZN(n7669) );
  AND2_X1 U5359 ( .A1(n9601), .A2(n9605), .ZN(n9611) );
  OAI211_X1 U5360 ( .C1(n7066), .C2(n5003), .A(n4552), .B(n7265), .ZN(n7148)
         );
  NAND2_X1 U5361 ( .A1(n6945), .A2(n5001), .ZN(n4552) );
  NOR2_X1 U5362 ( .A1(n5002), .A2(n5003), .ZN(n5001) );
  INV_X1 U5363 ( .A(n6388), .ZN(n5002) );
  NAND2_X1 U5364 ( .A1(n7067), .A2(n7066), .ZN(n7065) );
  AND2_X1 U5365 ( .A1(n9440), .A2(n9438), .ZN(n9547) );
  NAND2_X1 U5366 ( .A1(n10205), .A2(n7088), .ZN(n6462) );
  INV_X1 U5367 ( .A(n9777), .ZN(n9922) );
  NAND2_X1 U5368 ( .A1(n7657), .A2(n5214), .ZN(n4878) );
  INV_X1 U5369 ( .A(n9352), .ZN(n7845) );
  INV_X1 U5370 ( .A(n6489), .ZN(n7081) );
  AOI21_X1 U5371 ( .B1(n10202), .B2(n6461), .A(n6460), .ZN(n7080) );
  NAND2_X1 U5372 ( .A1(n4409), .A2(n5215), .ZN(n4555) );
  AOI21_X1 U5373 ( .B1(n5085), .B2(P1_IR_REG_24__SCAN_IN), .A(n5084), .ZN(
        n5824) );
  AND2_X1 U5374 ( .A1(n10074), .A2(n5083), .ZN(n5084) );
  XNOR2_X1 U5375 ( .A(n5705), .B(n5704), .ZN(n7679) );
  XNOR2_X1 U5376 ( .A(n5849), .B(n5848), .ZN(n6533) );
  INV_X1 U5377 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5848) );
  XNOR2_X1 U5378 ( .A(n5632), .B(SI_21_), .ZN(n7602) );
  OAI21_X1 U5379 ( .B1(n5609), .B2(n5608), .A(n5607), .ZN(n5627) );
  NAND2_X1 U5380 ( .A1(n4890), .A2(n5482), .ZN(n5505) );
  NAND2_X1 U5381 ( .A1(n4882), .A2(n4883), .ZN(n5371) );
  OR2_X1 U5382 ( .A1(n5326), .A2(n4886), .ZN(n4882) );
  XNOR2_X1 U5383 ( .A(n5326), .B(n5325), .ZN(n6527) );
  INV_X1 U5384 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U5385 ( .A1(n4839), .A2(n5243), .ZN(n5267) );
  NOR2_X1 U5386 ( .A1(n7952), .A2(n7953), .ZN(n7979) );
  XNOR2_X1 U5387 ( .A(n7998), .B(n7997), .ZN(n8033) );
  INV_X1 U5388 ( .A(n4749), .ZN(n4748) );
  OAI22_X1 U5389 ( .A1(n4754), .A2(n4750), .B1(n8692), .B2(n7989), .ZN(n4749)
         );
  AND2_X1 U5390 ( .A1(n6997), .A2(n6275), .ZN(n8384) );
  AND3_X1 U5391 ( .A1(n6209), .A2(n6208), .A3(n6207), .ZN(n8623) );
  NAND2_X1 U5392 ( .A1(n7749), .A2(n7748), .ZN(n7893) );
  INV_X1 U5393 ( .A(n8649), .ZN(n8677) );
  NAND2_X1 U5394 ( .A1(n6196), .A2(n6195), .ZN(n8627) );
  NAND2_X1 U5395 ( .A1(n6231), .A2(n6230), .ZN(n8129) );
  NOR2_X1 U5396 ( .A1(n4935), .A2(n8373), .ZN(n4934) );
  INV_X1 U5397 ( .A(n8577), .ZN(n8557) );
  XNOR2_X1 U5398 ( .A(n5990), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6799) );
  OR2_X1 U5399 ( .A1(n6727), .A2(n8376), .ZN(n10302) );
  XNOR2_X1 U5400 ( .A(n8472), .B(n8490), .ZN(n8450) );
  NOR2_X1 U5401 ( .A1(n8450), .A2(n8808), .ZN(n8474) );
  NAND2_X1 U5402 ( .A1(n4529), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4528) );
  NAND2_X1 U5403 ( .A1(n8507), .A2(n4529), .ZN(n4527) );
  NOR2_X1 U5404 ( .A1(n4468), .A2(n4529), .ZN(n4865) );
  INV_X1 U5405 ( .A(n4861), .ZN(n4860) );
  OAI211_X1 U5406 ( .C1(n10102), .C2(n10101), .A(n4438), .B(n4862), .ZN(n4861)
         );
  AOI21_X1 U5407 ( .B1(n10096), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n4524), .ZN(
        n4862) );
  OR2_X1 U5408 ( .A1(n5946), .A2(n5937), .ZN(n5938) );
  NAND2_X1 U5409 ( .A1(n6131), .A2(n6130), .ZN(n9152) );
  INV_X1 U5410 ( .A(n9147), .ZN(n9158) );
  AND2_X1 U5411 ( .A1(n6466), .A2(n9329), .ZN(n4973) );
  NOR2_X1 U5412 ( .A1(n4975), .A2(n9354), .ZN(n4974) );
  INV_X1 U5413 ( .A(n4441), .ZN(n4975) );
  NAND2_X1 U5414 ( .A1(n5882), .A2(n5770), .ZN(n6465) );
  INV_X1 U5415 ( .A(n9892), .ZN(n9992) );
  XNOR2_X1 U5416 ( .A(n5323), .B(n4498), .ZN(n7715) );
  NAND2_X1 U5417 ( .A1(n5495), .A2(n5494), .ZN(n10011) );
  NAND2_X1 U5418 ( .A1(n5544), .A2(n5543), .ZN(n10003) );
  NAND2_X1 U5419 ( .A1(n4587), .A2(n4585), .ZN(n9277) );
  AND2_X1 U5420 ( .A1(n4964), .A2(n4586), .ZN(n4585) );
  INV_X1 U5421 ( .A(n4965), .ZN(n4964) );
  AND2_X1 U5422 ( .A1(n4716), .A2(n5142), .ZN(n4715) );
  OR2_X1 U5423 ( .A1(n5587), .A2(n4550), .ZN(n5143) );
  INV_X1 U5424 ( .A(n7336), .ZN(n9334) );
  NAND2_X1 U5425 ( .A1(n9606), .A2(n9605), .ZN(n9607) );
  NAND2_X1 U5426 ( .A1(n5089), .A2(n10074), .ZN(n5090) );
  NAND2_X1 U5427 ( .A1(n6500), .A2(n6498), .ZN(n9614) );
  INV_X1 U5428 ( .A(n9371), .ZN(n9628) );
  INV_X1 U5429 ( .A(n7854), .ZN(n9631) );
  NAND4_X1 U5430 ( .A1(n5175), .A2(n5174), .A3(n5173), .A4(n5172), .ZN(n6385)
         );
  NAND2_X1 U5431 ( .A1(n5387), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5064) );
  NAND2_X1 U5432 ( .A1(n5221), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5063) );
  AND2_X1 U5433 ( .A1(n5115), .A2(n5114), .ZN(n5116) );
  INV_X1 U5434 ( .A(n6450), .ZN(n4856) );
  OR2_X1 U5435 ( .A1(n4415), .A2(n9705), .ZN(n9778) );
  NOR2_X2 U5436 ( .A1(n9614), .A2(n6462), .ZN(n10184) );
  INV_X1 U5437 ( .A(n9927), .ZN(n10186) );
  AOI21_X1 U5438 ( .B1(n9766), .B2(n4844), .A(n4843), .ZN(n4842) );
  INV_X1 U5439 ( .A(n4855), .ZN(n4854) );
  INV_X1 U5440 ( .A(n6495), .ZN(n4852) );
  AOI21_X1 U5441 ( .B1(n6452), .B2(n6494), .A(n6493), .ZN(n6495) );
  INV_X1 U5442 ( .A(n9759), .ZN(n10035) );
  AOI21_X1 U5443 ( .B1(n9725), .B2(n10217), .A(n4557), .ZN(n4855) );
  NAND2_X1 U5444 ( .A1(n9729), .A2(n4856), .ZN(n4557) );
  NAND2_X1 U5445 ( .A1(n10220), .A2(n10205), .ZN(n10067) );
  NAND2_X1 U5446 ( .A1(n4578), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4577) );
  NAND2_X1 U5447 ( .A1(n5562), .A2(n5561), .ZN(n4578) );
  NAND2_X1 U5448 ( .A1(n9422), .A2(n9421), .ZN(n4768) );
  OAI21_X1 U5449 ( .B1(n9439), .B2(n4789), .A(n4474), .ZN(n4795) );
  INV_X1 U5450 ( .A(n4790), .ZN(n4789) );
  AND2_X1 U5451 ( .A1(n9443), .A2(n9546), .ZN(n4794) );
  OAI211_X1 U5452 ( .C1(n8219), .C2(n8312), .A(n8221), .B(n4542), .ZN(n8228)
         );
  OR2_X1 U5453 ( .A1(n8220), .A2(n8285), .ZN(n4542) );
  AND2_X1 U5454 ( .A1(n9497), .A2(n9498), .ZN(n4805) );
  NOR2_X1 U5455 ( .A1(n9894), .A2(n9499), .ZN(n4804) );
  AND2_X1 U5456 ( .A1(n9528), .A2(n9534), .ZN(n4835) );
  AOI21_X1 U5457 ( .B1(n9510), .B2(n9840), .A(n4473), .ZN(n4787) );
  INV_X1 U5458 ( .A(n9801), .ZN(n9511) );
  NAND2_X1 U5459 ( .A1(n9800), .A2(n9513), .ZN(n4783) );
  AOI211_X1 U5460 ( .C1(n9505), .C2(n9840), .A(n9533), .B(n4785), .ZN(n4784)
         );
  NAND2_X1 U5461 ( .A1(n4444), .A2(n9542), .ZN(n9545) );
  INV_X1 U5462 ( .A(n9577), .ZN(n4818) );
  INV_X1 U5463 ( .A(n4831), .ZN(n4822) );
  AOI21_X1 U5464 ( .B1(n4825), .B2(n4821), .A(n4823), .ZN(n4820) );
  INV_X1 U5465 ( .A(n4826), .ZN(n4821) );
  NAND2_X1 U5466 ( .A1(n4859), .A2(n9447), .ZN(n6428) );
  INV_X1 U5467 ( .A(n9432), .ZN(n4859) );
  INV_X1 U5468 ( .A(n9447), .ZN(n9552) );
  NAND2_X1 U5469 ( .A1(n4922), .A2(n5626), .ZN(n4921) );
  INV_X1 U5470 ( .A(n5608), .ZN(n4922) );
  NAND2_X1 U5471 ( .A1(n4918), .A2(n5581), .ZN(n4915) );
  NOR2_X1 U5472 ( .A1(n4921), .A2(n4917), .ZN(n4916) );
  INV_X1 U5473 ( .A(n5581), .ZN(n4917) );
  AND2_X1 U5474 ( .A1(n8578), .A2(n8291), .ZN(n4540) );
  NOR2_X1 U5475 ( .A1(n6023), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6032) );
  INV_X1 U5476 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8776) );
  INV_X1 U5477 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n8893) );
  OAI21_X1 U5478 ( .B1(n6977), .B2(n5202), .A(n5107), .ZN(n4952) );
  INV_X1 U5479 ( .A(n4502), .ZN(n4918) );
  INV_X1 U5480 ( .A(n4896), .ZN(n4895) );
  INV_X1 U5481 ( .A(SI_17_), .ZN(n5536) );
  INV_X1 U5482 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5048) );
  NOR2_X1 U5483 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n5046) );
  NOR2_X1 U5484 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5045) );
  AND2_X1 U5485 ( .A1(n4736), .A2(n4734), .ZN(n4733) );
  INV_X1 U5486 ( .A(n4434), .ZN(n4731) );
  INV_X1 U5487 ( .A(n8336), .ZN(n4937) );
  OR2_X1 U5488 ( .A1(n6662), .A2(n10368), .ZN(n6710) );
  NAND2_X1 U5489 ( .A1(n6710), .A2(n6709), .ZN(n10225) );
  NAND2_X1 U5490 ( .A1(n10225), .A2(n10226), .ZN(n10224) );
  NAND2_X1 U5491 ( .A1(n4698), .A2(n4449), .ZN(n6785) );
  AOI21_X1 U5492 ( .B1(n4466), .B2(n6786), .A(n4706), .ZN(n7053) );
  INV_X1 U5493 ( .A(n7306), .ZN(n4874) );
  INV_X1 U5494 ( .A(n8427), .ZN(n4870) );
  NOR2_X1 U5495 ( .A1(n8453), .A2(n8452), .ZN(n8489) );
  AND2_X1 U5496 ( .A1(n8451), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8452) );
  AND2_X1 U5497 ( .A1(n8505), .A2(n8504), .ZN(n8506) );
  AND2_X1 U5498 ( .A1(n6233), .A2(n6232), .ZN(n6245) );
  OR2_X1 U5499 ( .A1(n6212), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6222) );
  NOR2_X1 U5500 ( .A1(n6176), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6185) );
  INV_X1 U5501 ( .A(n4647), .ZN(n4646) );
  AND2_X1 U5502 ( .A1(n4648), .A2(n8252), .ZN(n4647) );
  NAND2_X1 U5503 ( .A1(n8339), .A2(n6307), .ZN(n4648) );
  INV_X1 U5504 ( .A(n6307), .ZN(n4645) );
  AND2_X1 U5505 ( .A1(n6032), .A2(n8776), .ZN(n6047) );
  INV_X1 U5506 ( .A(n6289), .ZN(n4659) );
  INV_X1 U5507 ( .A(n4660), .ZN(n4656) );
  NOR2_X1 U5508 ( .A1(n10342), .A2(n7614), .ZN(n4655) );
  CLKBUF_X1 U5509 ( .A(n6279), .Z(n8342) );
  INV_X1 U5510 ( .A(n8167), .ZN(n5947) );
  OR2_X1 U5511 ( .A1(n6376), .A2(n8384), .ZN(n8334) );
  INV_X1 U5512 ( .A(n5911), .ZN(n6338) );
  INV_X1 U5513 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6372) );
  INV_X1 U5514 ( .A(n7178), .ZN(n4983) );
  NAND2_X1 U5515 ( .A1(n4499), .A2(n4980), .ZN(n4979) );
  NAND2_X1 U5516 ( .A1(n7782), .A2(n4499), .ZN(n4978) );
  NAND2_X1 U5517 ( .A1(n7783), .A2(n4499), .ZN(n4976) );
  NAND2_X1 U5518 ( .A1(n5235), .A2(n5234), .ZN(n4600) );
  NAND2_X1 U5519 ( .A1(n4960), .A2(n5207), .ZN(n5235) );
  NOR2_X1 U5520 ( .A1(n5339), .A2(n7786), .ZN(n5357) );
  NOR2_X1 U5521 ( .A1(n5635), .A2(n9035), .ZN(n5659) );
  AND2_X1 U5522 ( .A1(n4596), .A2(n4594), .ZN(n4593) );
  INV_X1 U5523 ( .A(n9256), .ZN(n4594) );
  NOR2_X1 U5524 ( .A1(n5545), .A2(n7582), .ZN(n5566) );
  AND2_X1 U5525 ( .A1(n5844), .A2(n6489), .ZN(n5865) );
  NAND2_X1 U5526 ( .A1(n4602), .A2(n6500), .ZN(n5322) );
  NAND2_X1 U5527 ( .A1(n4812), .A2(n9594), .ZN(n4811) );
  INV_X1 U5528 ( .A(n4433), .ZN(n5015) );
  NAND2_X1 U5529 ( .A1(n9895), .A2(n4640), .ZN(n4639) );
  INV_X1 U5530 ( .A(n6404), .ZN(n5024) );
  OR2_X1 U5531 ( .A1(n9992), .A2(n9280), .ZN(n9496) );
  INV_X1 U5532 ( .A(n4566), .ZN(n4559) );
  NOR2_X1 U5533 ( .A1(n5466), .A2(n5465), .ZN(n5496) );
  AND2_X1 U5534 ( .A1(n9396), .A2(n9487), .ZN(n9558) );
  INV_X1 U5535 ( .A(n9463), .ZN(n4630) );
  AND2_X1 U5536 ( .A1(n5357), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5383) );
  AND2_X1 U5537 ( .A1(n6432), .A2(n9457), .ZN(n4632) );
  INV_X1 U5538 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5248) );
  NOR2_X1 U5539 ( .A1(n7150), .A2(n9334), .ZN(n7151) );
  OR2_X1 U5540 ( .A1(n6452), .A2(n6885), .ZN(n9529) );
  OAI211_X1 U5541 ( .C1(n4617), .C2(n4770), .A(n9429), .B(n4619), .ZN(n6427)
         );
  OR2_X1 U5542 ( .A1(n4617), .A2(n4769), .ZN(n4619) );
  AND2_X1 U5543 ( .A1(n6265), .A2(n5811), .ZN(n6263) );
  AND2_X1 U5544 ( .A1(n5185), .A2(n5055), .ZN(n4798) );
  AND2_X1 U5545 ( .A1(n5806), .A2(n5780), .ZN(n5804) );
  INV_X1 U5546 ( .A(SI_19_), .ZN(n5583) );
  NAND2_X1 U5547 ( .A1(n4880), .A2(n4879), .ZN(n5400) );
  INV_X1 U5548 ( .A(n4887), .ZN(n4886) );
  NAND2_X1 U5549 ( .A1(n5303), .A2(n5302), .ZN(n5324) );
  AND2_X1 U5550 ( .A1(n5138), .A2(n5189), .ZN(n5139) );
  XNOR2_X1 U5551 ( .A(n5930), .B(P2_IR_REG_27__SCAN_IN), .ZN(n6331) );
  NAND2_X1 U5552 ( .A1(n4751), .A2(n4752), .ZN(n4750) );
  INV_X1 U5553 ( .A(n8114), .ZN(n4751) );
  AND2_X1 U5554 ( .A1(n4440), .A2(n4746), .ZN(n4745) );
  INV_X1 U5555 ( .A(n4750), .ZN(n4746) );
  XNOR2_X1 U5556 ( .A(n7137), .B(n4417), .ZN(n6900) );
  INV_X1 U5557 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n8799) );
  AND2_X1 U5558 ( .A1(n8225), .A2(n8223), .ZN(n8352) );
  XNOR2_X1 U5559 ( .A(n4417), .B(n7232), .ZN(n7014) );
  OR2_X1 U5560 ( .A1(n4753), .A2(n8070), .ZN(n4752) );
  INV_X1 U5561 ( .A(n4757), .ZN(n4753) );
  AND2_X1 U5562 ( .A1(n7985), .A2(n4757), .ZN(n4754) );
  INV_X1 U5563 ( .A(n7484), .ZN(n4767) );
  AND4_X1 U5564 ( .A1(n6124), .A2(n6123), .A3(n6122), .A4(n6121), .ZN(n7981)
         );
  AND4_X1 U5565 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n7750)
         );
  OR2_X1 U5566 ( .A1(n6713), .A2(n6721), .ZN(n6714) );
  NAND2_X1 U5567 ( .A1(n4699), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6768) );
  INV_X1 U5568 ( .A(n6706), .ZN(n4699) );
  NAND3_X1 U5569 ( .A1(n6714), .A2(n6761), .A3(P2_REG1_REG_3__SCAN_IN), .ZN(
        n6763) );
  NOR2_X1 U5570 ( .A1(n10266), .A2(n10378), .ZN(n10265) );
  NAND2_X1 U5571 ( .A1(n7201), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7316) );
  OAI21_X1 U5572 ( .B1(n7201), .B2(n4705), .A(n4703), .ZN(n7561) );
  AOI21_X1 U5573 ( .B1(n7315), .B2(n4704), .A(n7320), .ZN(n4703) );
  INV_X1 U5574 ( .A(n7315), .ZN(n4705) );
  AND2_X1 U5575 ( .A1(n7316), .A2(n7315), .ZN(n7321) );
  OR2_X1 U5576 ( .A1(n7196), .A2(n4873), .ZN(n4871) );
  NAND2_X1 U5577 ( .A1(n4874), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U5578 ( .A1(n7304), .A2(n4874), .ZN(n4872) );
  NOR2_X1 U5579 ( .A1(n7196), .A2(n7762), .ZN(n7305) );
  AND2_X1 U5580 ( .A1(n7563), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7833) );
  NAND2_X1 U5581 ( .A1(n4712), .A2(n4711), .ZN(n8405) );
  NAND2_X1 U5582 ( .A1(n7832), .A2(n4713), .ZN(n4711) );
  NOR2_X1 U5583 ( .A1(n8442), .A2(n8441), .ZN(n8453) );
  NAND2_X1 U5584 ( .A1(n8495), .A2(n8494), .ZN(n8512) );
  NOR2_X1 U5585 ( .A1(n10291), .A2(n10292), .ZN(n10290) );
  NOR2_X1 U5586 ( .A1(n10288), .A2(n10289), .ZN(n10287) );
  NAND2_X1 U5587 ( .A1(n4681), .A2(n4679), .ZN(n8575) );
  AND2_X1 U5588 ( .A1(n4685), .A2(n4680), .ZN(n4679) );
  INV_X1 U5589 ( .A(n4686), .ZN(n4685) );
  NOR2_X1 U5590 ( .A1(n8338), .A2(n4925), .ZN(n4924) );
  INV_X1 U5591 ( .A(n8156), .ZN(n4925) );
  OR2_X1 U5592 ( .A1(n6205), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6212) );
  NAND2_X1 U5593 ( .A1(n6197), .A2(n8799), .ZN(n6205) );
  AOI22_X1 U5594 ( .A1(n8633), .A2(n6312), .B1(n8624), .B2(n9130), .ZN(n8621)
         );
  AND2_X1 U5595 ( .A1(n8155), .A2(n8152), .ZN(n8638) );
  NAND2_X1 U5596 ( .A1(n6155), .A2(n6154), .ZN(n6168) );
  OR2_X1 U5597 ( .A1(n6168), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6176) );
  OR2_X1 U5598 ( .A1(n6108), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6119) );
  AND4_X1 U5599 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n7773)
         );
  NAND2_X1 U5600 ( .A1(n4662), .A2(n6286), .ZN(n4661) );
  NOR2_X1 U5601 ( .A1(n6288), .A2(n4663), .ZN(n4662) );
  INV_X1 U5602 ( .A(n6285), .ZN(n4663) );
  NAND2_X1 U5603 ( .A1(n7253), .A2(n4923), .ZN(n7372) );
  AND2_X1 U5604 ( .A1(n8199), .A2(n8186), .ZN(n4923) );
  NOR2_X1 U5605 ( .A1(n5932), .A2(n9356), .ZN(n4642) );
  AND2_X1 U5606 ( .A1(n6357), .A2(n6356), .ZN(n6915) );
  AND2_X1 U5607 ( .A1(n8334), .A2(n8306), .ZN(n8368) );
  AOI21_X1 U5608 ( .B1(n4947), .B2(n4949), .A(n4946), .ZN(n4945) );
  INV_X1 U5609 ( .A(n8149), .ZN(n4946) );
  AOI21_X1 U5610 ( .B1(n4665), .B2(n4667), .A(n4664), .ZN(n8648) );
  INV_X1 U5611 ( .A(n4666), .ZN(n4664) );
  AOI21_X1 U5612 ( .B1(n4667), .B2(n4671), .A(n4673), .ZN(n4666) );
  NAND2_X1 U5613 ( .A1(n4669), .A2(n6310), .ZN(n8658) );
  AND2_X1 U5614 ( .A1(n4669), .A2(n4667), .ZN(n8661) );
  AND2_X1 U5615 ( .A1(n6167), .A2(n6166), .ZN(n9139) );
  INV_X1 U5616 ( .A(n8252), .ZN(n8706) );
  OR2_X1 U5617 ( .A1(n7940), .A2(n8339), .ZN(n7942) );
  AND2_X1 U5618 ( .A1(n8248), .A2(n8247), .ZN(n8339) );
  OR2_X1 U5619 ( .A1(n7936), .A2(n8720), .ZN(n8713) );
  AND2_X1 U5620 ( .A1(n6088), .A2(n6087), .ZN(n8732) );
  INV_X1 U5621 ( .A(n8352), .ZN(n7894) );
  OR2_X1 U5622 ( .A1(n8312), .A2(n6894), .ZN(n6887) );
  INV_X1 U5623 ( .A(n9071), .ZN(n10353) );
  NAND2_X1 U5624 ( .A1(n6866), .A2(n6875), .ZN(n6925) );
  XNOR2_X1 U5625 ( .A(n6371), .B(n6372), .ZN(n6658) );
  AND2_X1 U5626 ( .A1(n4496), .A2(n5910), .ZN(n4933) );
  NAND2_X1 U5627 ( .A1(n5915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5927) );
  CLKBUF_X1 U5628 ( .A(n6329), .Z(n6330) );
  XNOR2_X1 U5629 ( .A(n6345), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U5630 ( .A1(n6149), .A2(n4951), .ZN(n6276) );
  AND2_X1 U5631 ( .A1(n5986), .A2(n5985), .ZN(n6783) );
  NOR2_X1 U5632 ( .A1(n5958), .A2(n4416), .ZN(n6711) );
  NAND2_X1 U5633 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5957) );
  AND2_X1 U5634 ( .A1(n5801), .A2(n5800), .ZN(n6467) );
  INV_X1 U5635 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5465) );
  XNOR2_X1 U5636 ( .A(n5178), .B(n5820), .ZN(n5180) );
  OR2_X1 U5637 ( .A1(n7365), .A2(n5600), .ZN(n5177) );
  NAND2_X1 U5638 ( .A1(n5169), .A2(n6975), .ZN(n5126) );
  INV_X1 U5639 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9035) );
  INV_X1 U5640 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5411) );
  INV_X1 U5641 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5497) );
  INV_X1 U5642 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7786) );
  OAI21_X1 U5643 ( .B1(n4968), .B2(n4966), .A(n9279), .ZN(n4965) );
  NOR2_X1 U5644 ( .A1(n4589), .A2(n4966), .ZN(n4588) );
  INV_X1 U5645 ( .A(n4590), .ZN(n4589) );
  NAND2_X1 U5646 ( .A1(n9316), .A2(n9317), .ZN(n4969) );
  AND2_X1 U5647 ( .A1(n4419), .A2(n9317), .ZN(n4968) );
  NAND2_X1 U5648 ( .A1(n9195), .A2(n5369), .ZN(n9306) );
  NAND2_X1 U5649 ( .A1(n5955), .A2(n4717), .ZN(n4716) );
  INV_X1 U5650 ( .A(n6416), .ZN(n4717) );
  INV_X1 U5651 ( .A(n5108), .ZN(n5111) );
  AOI21_X1 U5652 ( .B1(n4593), .B2(n4591), .A(n4517), .ZN(n4590) );
  INV_X1 U5653 ( .A(n4597), .ZN(n4591) );
  INV_X1 U5654 ( .A(n4593), .ZN(n4592) );
  INV_X1 U5655 ( .A(n9321), .ZN(n9301) );
  NOR2_X1 U5656 ( .A1(n5234), .A2(n4959), .ZN(n4958) );
  INV_X1 U5657 ( .A(n5207), .ZN(n4959) );
  AND2_X1 U5658 ( .A1(n5865), .A2(n6458), .ZN(n5864) );
  NAND2_X1 U5659 ( .A1(n9175), .A2(n5481), .ZN(n4598) );
  NAND2_X1 U5660 ( .A1(n4889), .A2(n6444), .ZN(n4780) );
  NAND2_X1 U5661 ( .A1(n9604), .A2(n7300), .ZN(n4889) );
  INV_X1 U5662 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5089) );
  NAND2_X1 U5663 ( .A1(n4554), .A2(n4553), .ZN(n5087) );
  INV_X1 U5664 ( .A(n4556), .ZN(n4553) );
  NOR2_X1 U5665 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5026) );
  AND2_X1 U5666 ( .A1(n5762), .A2(n5761), .ZN(n9236) );
  AND2_X1 U5667 ( .A1(n5712), .A2(n5711), .ZN(n9235) );
  AND2_X1 U5668 ( .A1(n5666), .A2(n5665), .ZN(n9217) );
  AND2_X1 U5669 ( .A1(n5620), .A2(n5619), .ZN(n9371) );
  AND4_X1 U5670 ( .A1(n5520), .A2(n5519), .A3(n5518), .A4(n5517), .ZN(n7853)
         );
  AND4_X1 U5671 ( .A1(n5471), .A2(n5470), .A3(n5469), .A4(n5468), .ZN(n7795)
         );
  AND4_X1 U5672 ( .A1(n5441), .A2(n5440), .A3(n5439), .A4(n5438), .ZN(n7703)
         );
  AND4_X1 U5673 ( .A1(n5417), .A2(n5416), .A3(n5415), .A4(n5414), .ZN(n7666)
         );
  AND4_X1 U5674 ( .A1(n5391), .A2(n5390), .A3(n5389), .A4(n5388), .ZN(n7506)
         );
  AND4_X1 U5675 ( .A1(n5364), .A2(n5363), .A3(n5362), .A4(n5361), .ZN(n7665)
         );
  AND4_X1 U5676 ( .A1(n5344), .A2(n5343), .A3(n5342), .A4(n5341), .ZN(n7344)
         );
  AND4_X1 U5677 ( .A1(n5287), .A2(n5286), .A3(n5285), .A4(n5284), .ZN(n7280)
         );
  INV_X1 U5678 ( .A(n5251), .ZN(n5221) );
  NAND2_X1 U5679 ( .A1(n5171), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5114) );
  AND2_X1 U5680 ( .A1(n9358), .A2(n6534), .ZN(n6536) );
  NOR2_X1 U5681 ( .A1(n6452), .A2(n4720), .ZN(n4718) );
  NAND2_X1 U5682 ( .A1(n7909), .A2(n9595), .ZN(n9300) );
  INV_X1 U5683 ( .A(n9574), .ZN(n9738) );
  NAND2_X1 U5684 ( .A1(n9791), .A2(n10039), .ZN(n9776) );
  AND2_X1 U5685 ( .A1(n5737), .A2(n5756), .ZN(n9793) );
  AND2_X1 U5686 ( .A1(n9800), .A2(n9801), .ZN(n4616) );
  AOI21_X1 U5687 ( .B1(n4637), .B2(n4635), .A(n4634), .ZN(n4633) );
  INV_X1 U5688 ( .A(n4637), .ZN(n4636) );
  INV_X1 U5689 ( .A(n9503), .ZN(n4634) );
  AND2_X1 U5690 ( .A1(n4639), .A2(n9416), .ZN(n9851) );
  NAND2_X1 U5691 ( .A1(n4639), .A2(n4637), .ZN(n9850) );
  NAND2_X1 U5692 ( .A1(n9858), .A2(n10058), .ZN(n9859) );
  NOR2_X1 U5693 ( .A1(n4425), .A2(n4849), .ZN(n4847) );
  NAND2_X1 U5694 ( .A1(n7858), .A2(n6455), .ZN(n9920) );
  NOR2_X1 U5695 ( .A1(n9563), .A2(n4564), .ZN(n4561) );
  NOR2_X1 U5696 ( .A1(n4723), .A2(n10015), .ZN(n7800) );
  INV_X1 U5697 ( .A(n9558), .ZN(n7636) );
  OR2_X1 U5698 ( .A1(n10187), .A2(n7506), .ZN(n9460) );
  AND2_X1 U5699 ( .A1(n9466), .A2(n9463), .ZN(n9557) );
  NAND2_X1 U5700 ( .A1(n7661), .A2(n4722), .ZN(n7638) );
  NAND2_X1 U5701 ( .A1(n5383), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5412) );
  NAND2_X1 U5702 ( .A1(n7661), .A2(n6454), .ZN(n7662) );
  INV_X1 U5703 ( .A(n9551), .ZN(n4840) );
  AND2_X1 U5704 ( .A1(n7351), .A2(n9205), .ZN(n7661) );
  NAND2_X1 U5705 ( .A1(n4991), .A2(n4990), .ZN(n7448) );
  AOI21_X1 U5706 ( .B1(n4992), .B2(n4994), .A(n4463), .ZN(n4990) );
  NOR2_X1 U5707 ( .A1(n7291), .A2(n7502), .ZN(n7455) );
  NAND2_X1 U5708 ( .A1(n7151), .A2(n6453), .ZN(n7291) );
  NAND2_X1 U5709 ( .A1(n6945), .A2(n6388), .ZN(n7067) );
  NAND2_X1 U5710 ( .A1(n7073), .A2(n7380), .ZN(n7150) );
  NOR2_X1 U5711 ( .A1(n6986), .A2(n6947), .ZN(n7073) );
  NAND2_X1 U5712 ( .A1(n6987), .A2(n7365), .ZN(n6986) );
  AND2_X1 U5713 ( .A1(n6974), .A2(n6383), .ZN(n6987) );
  NOR2_X1 U5714 ( .A1(n6975), .A2(n6977), .ZN(n6974) );
  AND2_X1 U5715 ( .A1(n5850), .A2(n9535), .ZN(n6456) );
  OAI21_X1 U5716 ( .B1(n6457), .B2(P1_D_REG_1__SCAN_IN), .A(n10072), .ZN(n7078) );
  OAI21_X1 U5717 ( .B1(n4845), .B2(n9755), .A(n9738), .ZN(n4843) );
  NAND2_X1 U5718 ( .A1(n5782), .A2(n5781), .ZN(n9759) );
  NAND2_X1 U5719 ( .A1(n7260), .A2(n6393), .ZN(n7279) );
  OAI21_X1 U5720 ( .B1(n7261), .B2(n4994), .A(n4992), .ZN(n7278) );
  NAND2_X1 U5721 ( .A1(n7290), .A2(n10208), .ZN(n10217) );
  INV_X1 U5722 ( .A(n9614), .ZN(n6458) );
  AND2_X1 U5723 ( .A1(n5000), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4998) );
  XNOR2_X1 U5724 ( .A(n8323), .B(n8322), .ZN(n9408) );
  AND2_X1 U5725 ( .A1(n5722), .A2(n5679), .ZN(n5698) );
  XNOR2_X1 U5726 ( .A(n5069), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U5727 ( .A1(n5075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U5728 ( .A1(n4987), .A2(n4986), .ZN(n5070) );
  AND2_X1 U5729 ( .A1(n5068), .A2(n5067), .ZN(n4986) );
  INV_X1 U5730 ( .A(n5491), .ZN(n4987) );
  OAI21_X1 U5731 ( .B1(n5491), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U5732 ( .A1(n4897), .A2(n4896), .ZN(n5535) );
  NAND2_X1 U5733 ( .A1(n4890), .A2(n4898), .ZN(n4897) );
  XNOR2_X1 U5734 ( .A(n4858), .B(n5033), .ZN(n6531) );
  OAI21_X1 U5735 ( .B1(n5326), .B2(n5325), .A(n5324), .ZN(n4858) );
  INV_X1 U5736 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5330) );
  INV_X1 U5737 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5331) );
  INV_X1 U5738 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5185) );
  OAI21_X1 U5739 ( .B1(n5153), .B2(n5100), .A(n5099), .ZN(n5101) );
  INV_X1 U5740 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5100) );
  NAND2_X1 U5741 ( .A1(n5153), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5099) );
  AND2_X1 U5742 ( .A1(n4764), .A2(n4448), .ZN(n7611) );
  NOR2_X1 U5743 ( .A1(n8024), .A2(n4742), .ZN(n4741) );
  INV_X1 U5744 ( .A(n8007), .ZN(n4742) );
  AND4_X1 U5745 ( .A1(n6072), .A2(n6071), .A3(n6070), .A4(n6069), .ZN(n7922)
         );
  AND4_X1 U5746 ( .A1(n6161), .A2(n6160), .A3(n6159), .A4(n6158), .ZN(n8663)
         );
  OAI21_X1 U5747 ( .B1(n8011), .B2(n6911), .A(n8167), .ZN(n6904) );
  NAND2_X1 U5748 ( .A1(n6183), .A2(n6182), .ZN(n8052) );
  AND4_X1 U5749 ( .A1(n6096), .A2(n6095), .A3(n6094), .A4(n6093), .ZN(n8235)
         );
  NAND2_X1 U5750 ( .A1(n6221), .A2(n6220), .ZN(n8761) );
  NAND2_X1 U5751 ( .A1(n8134), .A2(n7983), .ZN(n8064) );
  AND4_X1 U5752 ( .A1(n6135), .A2(n6134), .A3(n6133), .A4(n6132), .ZN(n8074)
         );
  NAND2_X1 U5753 ( .A1(n4755), .A2(n7985), .ZN(n8071) );
  NAND2_X1 U5754 ( .A1(n6140), .A2(n6139), .ZN(n9076) );
  NAND2_X1 U5755 ( .A1(n7998), .A2(n7997), .ZN(n7999) );
  NAND2_X1 U5756 ( .A1(n6211), .A2(n6210), .ZN(n8083) );
  AND4_X1 U5757 ( .A1(n6062), .A2(n6061), .A3(n6060), .A4(n6059), .ZN(n7754)
         );
  OAI21_X1 U5758 ( .B1(n7915), .B2(n4760), .A(n4759), .ZN(n4758) );
  NAND2_X1 U5759 ( .A1(n4762), .A2(n4761), .ZN(n4760) );
  INV_X1 U5760 ( .A(n7901), .ZN(n4759) );
  NAND2_X1 U5761 ( .A1(n8087), .A2(n4434), .ZN(n4735) );
  AND4_X1 U5762 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n8104)
         );
  AND4_X1 U5763 ( .A1(n6148), .A2(n6147), .A3(n6146), .A4(n6145), .ZN(n8675)
         );
  NAND2_X1 U5764 ( .A1(n4747), .A2(n4752), .ZN(n8115) );
  NAND2_X1 U5765 ( .A1(n4755), .A2(n4754), .ZN(n4747) );
  NAND2_X1 U5766 ( .A1(n6153), .A2(n6152), .ZN(n8683) );
  INV_X1 U5767 ( .A(n8396), .ZN(n7490) );
  NAND2_X1 U5768 ( .A1(n7485), .A2(n7484), .ZN(n7487) );
  NAND2_X1 U5769 ( .A1(n7013), .A2(n8381), .ZN(n8141) );
  XNOR2_X1 U5770 ( .A(n6277), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8379) );
  AND2_X1 U5771 ( .A1(n6997), .A2(n6996), .ZN(n8539) );
  INV_X1 U5772 ( .A(n8590), .ZN(n8568) );
  INV_X1 U5773 ( .A(n8604), .ZN(n8385) );
  INV_X1 U5774 ( .A(n8635), .ZN(n8614) );
  INV_X1 U5775 ( .A(n8675), .ZN(n8707) );
  INV_X1 U5776 ( .A(n8074), .ZN(n8691) );
  INV_X1 U5777 ( .A(n7981), .ZN(n8718) );
  INV_X1 U5778 ( .A(n8104), .ZN(n8389) );
  INV_X1 U5779 ( .A(n7754), .ZN(n8391) );
  INV_X1 U5780 ( .A(n7773), .ZN(n8392) );
  INV_X1 U5781 ( .A(n7750), .ZN(n8393) );
  AND2_X1 U5782 ( .A1(n5950), .A2(n5949), .ZN(n5953) );
  OR2_X1 U5783 ( .A1(n6866), .A2(n6501), .ZN(n8399) );
  INV_X1 U5784 ( .A(n10283), .ZN(n10096) );
  AND2_X1 U5785 ( .A1(n7050), .A2(n7049), .ZN(n5042) );
  INV_X1 U5786 ( .A(n7030), .ZN(n10245) );
  OAI21_X1 U5787 ( .B1(n10266), .B2(n4536), .A(n4535), .ZN(n7192) );
  NAND2_X1 U5788 ( .A1(n4537), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4536) );
  INV_X1 U5789 ( .A(n4869), .ZN(n8425) );
  OR2_X1 U5790 ( .A1(n8402), .A2(n8403), .ZN(n4869) );
  INV_X1 U5791 ( .A(n8426), .ZN(n4868) );
  NAND2_X1 U5792 ( .A1(n4526), .A2(n4866), .ZN(n8449) );
  OR2_X1 U5793 ( .A1(n8474), .A2(n8473), .ZN(n8477) );
  OAI21_X1 U5794 ( .B1(n8518), .B2(n10302), .A(n4465), .ZN(n4531) );
  NOR2_X1 U5795 ( .A1(n10097), .A2(n8516), .ZN(n8517) );
  INV_X1 U5796 ( .A(n8508), .ZN(n4534) );
  INV_X1 U5797 ( .A(n6336), .ZN(n4676) );
  NAND2_X1 U5798 ( .A1(n4691), .A2(n4684), .ZN(n4688) );
  OR2_X1 U5799 ( .A1(n10359), .A2(n7125), .ZN(n8731) );
  NAND2_X1 U5800 ( .A1(n4691), .A2(n4689), .ZN(n8602) );
  INV_X1 U5801 ( .A(n9139), .ZN(n8669) );
  NAND2_X1 U5802 ( .A1(n6118), .A2(n6117), .ZN(n7980) );
  NAND2_X1 U5803 ( .A1(n7758), .A2(n8208), .ZN(n7772) );
  NAND2_X1 U5804 ( .A1(n4543), .A2(n6031), .ZN(n7743) );
  NAND2_X1 U5805 ( .A1(n6527), .A2(n5962), .ZN(n4543) );
  AND3_X1 U5806 ( .A1(n6022), .A2(n6021), .A3(n6020), .ZN(n10348) );
  NAND2_X1 U5807 ( .A1(n4927), .A2(n8193), .ZN(n7593) );
  NAND2_X1 U5808 ( .A1(n7253), .A2(n8186), .ZN(n7241) );
  INV_X1 U5809 ( .A(n10337), .ZN(n7248) );
  NAND2_X1 U5810 ( .A1(n10317), .A2(n10308), .ZN(n8728) );
  INV_X1 U5811 ( .A(n8699), .ZN(n10312) );
  AND2_X1 U5812 ( .A1(n10384), .A2(n10325), .ZN(n9084) );
  NAND2_X1 U5813 ( .A1(n8328), .A2(n8327), .ZN(n9088) );
  INV_X1 U5814 ( .A(n8744), .ZN(n9094) );
  NAND2_X1 U5815 ( .A1(n6253), .A2(n6252), .ZN(n9097) );
  AOI21_X1 U5816 ( .B1(n8561), .B2(n8722), .A(n8560), .ZN(n9095) );
  NAND2_X1 U5817 ( .A1(n8559), .A2(n8558), .ZN(n8560) );
  XNOR2_X1 U5818 ( .A(n8555), .B(n8554), .ZN(n8561) );
  NAND2_X1 U5819 ( .A1(n8756), .A2(n8293), .ZN(n8565) );
  NAND2_X1 U5820 ( .A1(n4926), .A2(n8156), .ZN(n8611) );
  INV_X1 U5821 ( .A(n8052), .ZN(n9130) );
  NAND2_X1 U5822 ( .A1(n6175), .A2(n6174), .ZN(n9133) );
  NAND2_X1 U5823 ( .A1(n6107), .A2(n6106), .ZN(n9159) );
  INV_X1 U5824 ( .A(n8732), .ZN(n7936) );
  NAND2_X1 U5825 ( .A1(n6077), .A2(n6076), .ZN(n7969) );
  AND3_X1 U5826 ( .A1(n5993), .A2(n5992), .A3(n5991), .ZN(n7467) );
  AND2_X1 U5827 ( .A1(n6658), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6875) );
  NAND2_X1 U5828 ( .A1(n6343), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6344) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7710) );
  INV_X1 U5830 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7647) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7379) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7302) );
  INV_X1 U5833 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9018) );
  NOR2_X1 U5834 ( .A1(n6129), .A2(n6137), .ZN(n8523) );
  INV_X1 U5835 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6832) );
  INV_X1 U5836 ( .A(n8463), .ZN(n8451) );
  INV_X1 U5837 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6562) );
  INV_X1 U5838 ( .A(n7562), .ZN(n7830) );
  INV_X1 U5839 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U5840 ( .A1(n5936), .A2(n5935), .ZN(n6689) );
  NOR2_X1 U5841 ( .A1(n9188), .A2(n4582), .ZN(n4581) );
  NAND2_X1 U5842 ( .A1(n9195), .A2(n4612), .ZN(n4609) );
  INV_X1 U5843 ( .A(n4605), .ZN(n4612) );
  NAND2_X1 U5844 ( .A1(n9175), .A2(n4597), .ZN(n4595) );
  INV_X1 U5845 ( .A(n7459), .ZN(n10213) );
  NAND2_X1 U5846 ( .A1(n4981), .A2(n5349), .ZN(n4977) );
  INV_X1 U5847 ( .A(n7783), .ZN(n4981) );
  NAND2_X1 U5848 ( .A1(n4963), .A2(n4967), .ZN(n9278) );
  NAND2_X1 U5849 ( .A1(n9315), .A2(n4968), .ZN(n4963) );
  INV_X1 U5850 ( .A(n4607), .ZN(n4606) );
  AOI21_X1 U5851 ( .B1(n4605), .B2(n4607), .A(n4515), .ZN(n4604) );
  NOR2_X1 U5852 ( .A1(n9224), .A2(n4608), .ZN(n4607) );
  NAND2_X1 U5853 ( .A1(n4957), .A2(n9189), .ZN(n9299) );
  NAND2_X1 U5854 ( .A1(n5658), .A2(n5657), .ZN(n9842) );
  AND2_X1 U5855 ( .A1(n5151), .A2(n5152), .ZN(n6820) );
  NAND2_X1 U5856 ( .A1(n5565), .A2(n5564), .ZN(n9911) );
  OR2_X1 U5857 ( .A1(n5872), .A2(n5871), .ZN(n9337) );
  INV_X1 U5858 ( .A(n9283), .ZN(n9351) );
  INV_X1 U5859 ( .A(n9236), .ZN(n9622) );
  INV_X1 U5860 ( .A(n9512), .ZN(n9625) );
  INV_X1 U5861 ( .A(n9217), .ZN(n9626) );
  OR2_X1 U5862 ( .A1(n5501), .A2(n5500), .ZN(n9632) );
  OR2_X1 U5863 ( .A1(n5129), .A2(n6830), .ZN(n5131) );
  AOI22_X1 U5864 ( .A1(n4614), .A2(P1_REG0_REG_2__SCAN_IN), .B1(
        P1_REG2_REG_2__SCAN_IN), .B2(n5387), .ZN(n4613) );
  OR2_X1 U5865 ( .A1(n6500), .A2(n6499), .ZN(n9646) );
  AND2_X1 U5866 ( .A1(n6556), .A2(n5856), .ZN(n10173) );
  NAND2_X1 U5867 ( .A1(n9754), .A2(n9753), .ZN(n9950) );
  OAI21_X1 U5868 ( .B1(n9807), .B2(n5008), .A(n5006), .ZN(n9756) );
  NAND2_X1 U5869 ( .A1(n5009), .A2(n5010), .ZN(n9772) );
  NAND2_X1 U5870 ( .A1(n9807), .A2(n5011), .ZN(n5009) );
  OAI21_X1 U5871 ( .B1(n9807), .B2(n4420), .A(n6411), .ZN(n9790) );
  OAI21_X1 U5872 ( .B1(n9885), .B2(n4575), .A(n4572), .ZN(n9824) );
  AOI211_X1 U5873 ( .C1(n9827), .C2(n4728), .A(n9922), .B(n9826), .ZN(n9972)
         );
  NAND2_X1 U5874 ( .A1(n5018), .A2(n5019), .ZN(n9839) );
  NAND2_X1 U5875 ( .A1(n9874), .A2(n4433), .ZN(n5018) );
  OAI21_X1 U5876 ( .B1(n9874), .B2(n4437), .A(n6408), .ZN(n9857) );
  AND2_X1 U5877 ( .A1(n5590), .A2(n5589), .ZN(n9892) );
  NAND2_X1 U5878 ( .A1(n5025), .A2(n6404), .ZN(n9903) );
  NAND2_X1 U5879 ( .A1(n7851), .A2(n9484), .ZN(n9928) );
  NAND2_X1 U5880 ( .A1(n4562), .A2(n4563), .ZN(n7857) );
  NAND2_X1 U5881 ( .A1(n4562), .A2(n4561), .ZN(n10008) );
  NAND2_X1 U5882 ( .A1(n5511), .A2(n5510), .ZN(n9352) );
  OAI21_X1 U5883 ( .B1(n7696), .B2(n6400), .A(n6399), .ZN(n7799) );
  INV_X1 U5884 ( .A(n10184), .ZN(n9774) );
  NAND2_X1 U5885 ( .A1(n7065), .A2(n6390), .ZN(n7149) );
  NAND2_X1 U5886 ( .A1(n9422), .A2(n4620), .ZN(n7068) );
  NAND2_X1 U5887 ( .A1(n9422), .A2(n9428), .ZN(n6948) );
  NOR2_X1 U5888 ( .A1(n6969), .A2(n4771), .ZN(n7171) );
  INV_X1 U5889 ( .A(n9778), .ZN(n10189) );
  AND2_X1 U5890 ( .A1(n6456), .A2(n9605), .ZN(n9777) );
  NAND2_X1 U5891 ( .A1(n5356), .A2(n5355), .ZN(n7426) );
  NOR2_X1 U5892 ( .A1(n9950), .A2(n4625), .ZN(n10033) );
  NAND2_X1 U5893 ( .A1(n4627), .A2(n4626), .ZN(n4625) );
  INV_X1 U5894 ( .A(n9951), .ZN(n4626) );
  NAND2_X1 U5895 ( .A1(n9952), .A2(n10217), .ZN(n4627) );
  NOR2_X1 U5896 ( .A1(n10035), .A2(n10067), .ZN(n4623) );
  INV_X1 U5897 ( .A(n9878), .ZN(n10062) );
  NAND2_X1 U5898 ( .A1(n5409), .A2(n5408), .ZN(n9229) );
  INV_X1 U5899 ( .A(n7426), .ZN(n9205) );
  AND2_X1 U5900 ( .A1(n5247), .A2(n5246), .ZN(n7336) );
  INV_X1 U5901 ( .A(n6389), .ZN(n7380) );
  NAND2_X1 U5902 ( .A1(n6458), .A2(n6457), .ZN(n10202) );
  XNOR2_X1 U5903 ( .A(n5079), .B(P1_IR_REG_26__SCAN_IN), .ZN(n7868) );
  INV_X1 U5904 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8783) );
  INV_X1 U5905 ( .A(n9601), .ZN(n9535) );
  INV_X1 U5906 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8952) );
  INV_X1 U5907 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8976) );
  INV_X1 U5908 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8975) );
  INV_X1 U5909 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6943) );
  INV_X1 U5910 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9016) );
  INV_X1 U5911 ( .A(n10133), .ZN(n7411) );
  INV_X1 U5912 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6778) );
  INV_X1 U5913 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6563) );
  INV_X1 U5914 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6542) );
  INV_X1 U5915 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6528) );
  INV_X1 U5916 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7548) );
  NAND2_X1 U5917 ( .A1(n4863), .A2(n4460), .ZN(P2_U3200) );
  NAND2_X1 U5918 ( .A1(n4864), .A2(n10228), .ZN(n4863) );
  OR2_X1 U5919 ( .A1(n4865), .A2(n10094), .ZN(n4864) );
  OAI21_X1 U5920 ( .B1(n4532), .B2(n10293), .A(n4530), .ZN(P2_U3201) );
  XNOR2_X1 U5921 ( .A(n4534), .B(n4533), .ZN(n4532) );
  INV_X1 U5922 ( .A(n4531), .ZN(n4530) );
  INV_X1 U5923 ( .A(n8519), .ZN(n4533) );
  OAI21_X1 U5924 ( .B1(n4678), .B2(n4675), .A(n4674), .ZN(P2_U3456) );
  INV_X1 U5925 ( .A(n6487), .ZN(n4675) );
  AOI21_X1 U5926 ( .B1(n6465), .B2(n4974), .A(n4972), .ZN(n4970) );
  OR2_X1 U5927 ( .A1(n4429), .A2(n6476), .ZN(n4972) );
  OAI21_X1 U5928 ( .B1(n10039), .B2(n9283), .A(n5891), .ZN(n5892) );
  AOI21_X1 U5929 ( .B1(n4778), .B2(n9607), .A(n4476), .ZN(n9618) );
  AND2_X1 U5930 ( .A1(n4857), .A2(n4856), .ZN(n9734) );
  AOI21_X1 U5931 ( .B1(n4853), .B2(n4854), .A(n4852), .ZN(n4851) );
  AOI21_X1 U5932 ( .B1(n4855), .B2(n9906), .A(n6496), .ZN(n4853) );
  AND2_X1 U5933 ( .A1(n4855), .A2(n4857), .ZN(n6497) );
  NAND2_X1 U5934 ( .A1(n4624), .A2(n4621), .ZN(P1_U3517) );
  NOR2_X1 U5935 ( .A1(n4623), .A2(n4622), .ZN(n4621) );
  OR2_X1 U5936 ( .A1(n10033), .A2(n10218), .ZN(n4624) );
  NOR2_X1 U5937 ( .A1(n10220), .A2(n10034), .ZN(n4622) );
  INV_X2 U5938 ( .A(n5153), .ZN(n5212) );
  OR2_X1 U5939 ( .A1(n9878), .A2(n9371), .ZN(n9416) );
  AND2_X1 U5940 ( .A1(n4598), .A2(n4447), .ZN(n9242) );
  NAND2_X1 U5941 ( .A1(n5605), .A2(n9207), .ZN(n4419) );
  NOR2_X1 U5942 ( .A1(n9810), .A2(n9624), .ZN(n4420) );
  INV_X2 U5943 ( .A(n5170), .ZN(n4614) );
  NAND2_X1 U5944 ( .A1(n4456), .A2(n4957), .ZN(n9187) );
  INV_X1 U5945 ( .A(n5851), .ZN(n5850) );
  AND2_X1 U5946 ( .A1(n4590), .A2(n4592), .ZN(n4421) );
  AND2_X1 U5947 ( .A1(n4951), .A2(n4457), .ZN(n4422) );
  AND2_X1 U5948 ( .A1(n4725), .A2(n4724), .ZN(n4423) );
  NAND2_X1 U5949 ( .A1(n9720), .A2(n9619), .ZN(n4424) );
  AND2_X1 U5950 ( .A1(n4848), .A2(n9929), .ZN(n4425) );
  AND2_X1 U5951 ( .A1(n8083), .A2(n8615), .ZN(n4426) );
  INV_X1 U5952 ( .A(n5012), .ZN(n5011) );
  OR2_X1 U5953 ( .A1(n5013), .A2(n6412), .ZN(n5012) );
  INV_X1 U5954 ( .A(n6452), .ZN(n6491) );
  AND2_X1 U5955 ( .A1(n9484), .A2(n9492), .ZN(n9563) );
  AND2_X1 U5956 ( .A1(n8277), .A2(n6332), .ZN(n4427) );
  NAND2_X1 U5957 ( .A1(n4677), .A2(n10367), .ZN(n4428) );
  AND2_X1 U5958 ( .A1(n6466), .A2(n4442), .ZN(n4429) );
  NAND2_X1 U5959 ( .A1(n5813), .A2(n5812), .ZN(n9742) );
  INV_X1 U5960 ( .A(n9742), .ZN(n10032) );
  INV_X1 U5961 ( .A(n8591), .ZN(n8615) );
  AND2_X1 U5962 ( .A1(n6218), .A2(n6217), .ZN(n8591) );
  NAND2_X1 U5963 ( .A1(n4516), .A2(n7178), .ZN(n7177) );
  INV_X1 U5964 ( .A(n10095), .ZN(n4529) );
  AND2_X1 U5965 ( .A1(n6500), .A2(n9611), .ZN(n5236) );
  INV_X1 U5966 ( .A(n5236), .ZN(n5345) );
  NAND2_X1 U5967 ( .A1(n6897), .A2(n6896), .ZN(n6902) );
  AND2_X1 U5968 ( .A1(n5184), .A2(n5185), .ZN(n5215) );
  NAND3_X1 U5969 ( .A1(n5027), .A2(n4409), .A3(n5215), .ZN(n4430) );
  OR2_X1 U5970 ( .A1(n4555), .A2(n4556), .ZN(n4431) );
  NAND2_X1 U5971 ( .A1(n9827), .A2(n9625), .ZN(n4432) );
  NOR2_X1 U5972 ( .A1(n6409), .A2(n5022), .ZN(n4433) );
  AND2_X1 U5973 ( .A1(n4740), .A2(n4739), .ZN(n4434) );
  NAND2_X1 U5974 ( .A1(n8764), .A2(n8591), .ZN(n4435) );
  NAND2_X1 U5975 ( .A1(n5463), .A2(n5462), .ZN(n10015) );
  NOR2_X1 U5976 ( .A1(n9892), .A2(n9280), .ZN(n4436) );
  NOR2_X1 U5977 ( .A1(n9878), .A2(n9628), .ZN(n4437) );
  INV_X1 U5978 ( .A(n9436), .ZN(n4769) );
  INV_X1 U5979 ( .A(n10254), .ZN(n7052) );
  INV_X1 U5980 ( .A(n8206), .ZN(n8347) );
  AND2_X1 U5981 ( .A1(n7685), .A2(n8212), .ZN(n8206) );
  OR3_X1 U5982 ( .A1(n10093), .A2(n10092), .A3(n10091), .ZN(n4438) );
  AND2_X1 U5983 ( .A1(n9791), .A2(n4719), .ZN(n4439) );
  NOR2_X1 U5984 ( .A1(n7986), .A2(n4756), .ZN(n4440) );
  NAND2_X2 U5985 ( .A1(n4996), .A2(n4999), .ZN(n5251) );
  AND2_X1 U5986 ( .A1(n5803), .A2(n5802), .ZN(n4441) );
  INV_X1 U5987 ( .A(n5008), .ZN(n5007) );
  NAND2_X1 U5988 ( .A1(n5010), .A2(n4453), .ZN(n5008) );
  NAND2_X1 U5989 ( .A1(n5143), .A2(n4715), .ZN(n7140) );
  AND2_X1 U5990 ( .A1(n6467), .A2(n9329), .ZN(n4442) );
  AND2_X1 U5991 ( .A1(n8393), .A2(n7743), .ZN(n4443) );
  AND3_X1 U5992 ( .A1(n9543), .A2(n6423), .A3(n9541), .ZN(n4444) );
  INV_X1 U5993 ( .A(n9428), .ZN(n4618) );
  NAND2_X1 U5994 ( .A1(n5634), .A2(n5633), .ZN(n9861) );
  NAND2_X1 U5995 ( .A1(n5434), .A2(n5433), .ZN(n9294) );
  AND2_X1 U5996 ( .A1(n9895), .A2(n9475), .ZN(n4445) );
  AND2_X1 U5997 ( .A1(n6342), .A2(n6343), .ZN(n6347) );
  AND2_X1 U5998 ( .A1(n8549), .A2(n6278), .ZN(n4446) );
  NAND2_X1 U5999 ( .A1(n5480), .A2(n5479), .ZN(n4447) );
  OR2_X1 U6000 ( .A1(n9119), .A2(n8623), .ZN(n8279) );
  NAND2_X1 U6001 ( .A1(n7607), .A2(n8395), .ZN(n4448) );
  NAND2_X1 U6002 ( .A1(n4743), .A2(n4741), .ZN(n8025) );
  AND2_X1 U6003 ( .A1(n6765), .A2(n4697), .ZN(n4449) );
  NAND2_X1 U6004 ( .A1(n4878), .A2(n5680), .ZN(n9827) );
  INV_X1 U6005 ( .A(n5169), .ZN(n5600) );
  NOR2_X1 U6006 ( .A1(n8657), .A2(n4668), .ZN(n4667) );
  NOR2_X1 U6007 ( .A1(n7969), .A2(n8389), .ZN(n4450) );
  AND2_X1 U6008 ( .A1(n4722), .A2(n7639), .ZN(n4451) );
  NOR2_X1 U6009 ( .A1(n10287), .A2(n8514), .ZN(n4452) );
  NAND2_X1 U6010 ( .A1(n5382), .A2(n5381), .ZN(n10187) );
  OR2_X1 U6011 ( .A1(n9781), .A2(n9622), .ZN(n4453) );
  AND2_X1 U6012 ( .A1(n9789), .A2(n9784), .ZN(n4454) );
  INV_X1 U6013 ( .A(n9781), .ZN(n10039) );
  INV_X1 U6014 ( .A(n9526), .ZN(n4836) );
  AND2_X1 U6015 ( .A1(n4575), .A2(n4432), .ZN(n4455) );
  AND2_X1 U6016 ( .A1(n9189), .A2(n9297), .ZN(n4456) );
  AND2_X1 U6017 ( .A1(n6320), .A2(n5908), .ZN(n4457) );
  INV_X1 U6018 ( .A(n4792), .ZN(n4791) );
  OAI21_X1 U6019 ( .B1(n4793), .B2(n9438), .A(n9442), .ZN(n4792) );
  INV_X1 U6020 ( .A(n4988), .ZN(n5081) );
  NOR2_X1 U6021 ( .A1(n5075), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4988) );
  AND2_X1 U6022 ( .A1(n5004), .A2(n6414), .ZN(n4458) );
  INV_X1 U6023 ( .A(n4671), .ZN(n4670) );
  OR2_X1 U6024 ( .A1(n6311), .A2(n4672), .ZN(n4671) );
  AND2_X1 U6025 ( .A1(n9781), .A2(n9622), .ZN(n4459) );
  AND2_X1 U6026 ( .A1(n10100), .A2(n4860), .ZN(n4460) );
  INV_X1 U6027 ( .A(n4690), .ZN(n4689) );
  NOR2_X1 U6028 ( .A1(n6313), .A2(n8623), .ZN(n4690) );
  OR2_X1 U6029 ( .A1(n10011), .A2(n9258), .ZN(n9484) );
  INV_X1 U6030 ( .A(n9484), .ZN(n4848) );
  INV_X1 U6031 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10074) );
  AND2_X1 U6032 ( .A1(n9152), .A2(n8691), .ZN(n4461) );
  NAND2_X1 U6033 ( .A1(n6406), .A2(n6405), .ZN(n9885) );
  INV_X1 U6034 ( .A(n9885), .ZN(n4568) );
  AND2_X1 U6035 ( .A1(n8151), .A2(n8150), .ZN(n4462) );
  NOR2_X1 U6036 ( .A1(n7502), .A2(n9640), .ZN(n4463) );
  INV_X1 U6037 ( .A(n4564), .ZN(n4563) );
  OAI21_X1 U6038 ( .B1(n6401), .B2(n4565), .A(n6402), .ZN(n4564) );
  NOR2_X1 U6039 ( .A1(n9792), .A2(n9623), .ZN(n4464) );
  AND2_X1 U6040 ( .A1(n8536), .A2(n4714), .ZN(n4465) );
  AND2_X1 U6041 ( .A1(n9516), .A2(n9515), .ZN(n9523) );
  NOR2_X1 U6042 ( .A1(n10248), .A2(n4709), .ZN(n4466) );
  NAND2_X1 U6043 ( .A1(n9496), .A2(n4805), .ZN(n4467) );
  OAI21_X1 U6044 ( .B1(n4848), .B2(n9494), .A(n9492), .ZN(n4806) );
  OR2_X1 U6045 ( .A1(n10290), .A2(n8507), .ZN(n4468) );
  INV_X1 U6046 ( .A(n8195), .ZN(n8208) );
  AND2_X1 U6047 ( .A1(n7766), .A2(n8392), .ZN(n8195) );
  AND2_X1 U6048 ( .A1(n9842), .A2(n9626), .ZN(n4469) );
  NAND2_X1 U6049 ( .A1(n6149), .A2(n5906), .ZN(n4470) );
  NAND2_X1 U6050 ( .A1(n6149), .A2(n4422), .ZN(n4471) );
  INV_X1 U6051 ( .A(n4720), .ZN(n4719) );
  NAND2_X1 U6052 ( .A1(n10032), .A2(n4721), .ZN(n4720) );
  AND2_X1 U6053 ( .A1(n5370), .A2(SI_10_), .ZN(n4472) );
  INV_X1 U6054 ( .A(n4845), .ZN(n4844) );
  OAI21_X1 U6055 ( .B1(n9571), .B2(n9518), .A(n9526), .ZN(n4845) );
  NAND2_X1 U6056 ( .A1(n9366), .A2(n9365), .ZN(n4473) );
  AND2_X1 U6057 ( .A1(n4788), .A2(n4796), .ZN(n4474) );
  INV_X1 U6058 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5056) );
  INV_X1 U6059 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5067) );
  INV_X1 U6060 ( .A(n9441), .ZN(n4797) );
  NOR2_X1 U6061 ( .A1(n5534), .A2(n4895), .ZN(n4894) );
  OR2_X1 U6062 ( .A1(n9523), .A2(n4822), .ZN(n4475) );
  INV_X1 U6063 ( .A(n4899), .ZN(n4898) );
  NAND2_X1 U6064 ( .A1(n4501), .A2(n5482), .ZN(n4899) );
  NOR2_X1 U6065 ( .A1(n9609), .A2(n9608), .ZN(n4476) );
  NOR2_X1 U6066 ( .A1(n7996), .A2(n8614), .ZN(n4477) );
  AND2_X1 U6067 ( .A1(n4801), .A2(n4467), .ZN(n4478) );
  INV_X1 U6068 ( .A(n4967), .ZN(n4966) );
  NAND2_X1 U6069 ( .A1(n4481), .A2(n4419), .ZN(n4967) );
  OR2_X1 U6070 ( .A1(n6426), .A2(n4618), .ZN(n4617) );
  NAND2_X1 U6071 ( .A1(n5532), .A2(n4447), .ZN(n4479) );
  OR2_X1 U6072 ( .A1(n9522), .A2(n9533), .ZN(n4480) );
  NAND2_X1 U6073 ( .A1(n5606), .A2(n4969), .ZN(n4481) );
  INV_X1 U6074 ( .A(n8690), .ZN(n8696) );
  AND2_X1 U6075 ( .A1(n8260), .A2(n8680), .ZN(n8690) );
  OR2_X1 U6076 ( .A1(n9842), .A2(n9626), .ZN(n4482) );
  AND2_X1 U6077 ( .A1(n5006), .A2(n9571), .ZN(n4483) );
  AND2_X1 U6078 ( .A1(n8158), .A2(n8285), .ZN(n4484) );
  AND2_X1 U6079 ( .A1(n4688), .A2(n4435), .ZN(n4485) );
  AND2_X1 U6080 ( .A1(n8289), .A2(n8290), .ZN(n8587) );
  NOR2_X1 U6081 ( .A1(n8332), .A2(n8333), .ZN(n4486) );
  AND2_X1 U6082 ( .A1(n9088), .A2(n8539), .ZN(n4487) );
  OR2_X1 U6083 ( .A1(n4815), .A2(n4813), .ZN(n4488) );
  AND2_X1 U6084 ( .A1(n8334), .A2(n9097), .ZN(n4489) );
  AND2_X1 U6085 ( .A1(n8206), .A2(n8193), .ZN(n4490) );
  NAND2_X1 U6086 ( .A1(n9522), .A2(n9526), .ZN(n4491) );
  AND2_X1 U6087 ( .A1(n5184), .A2(n4798), .ZN(n4492) );
  AND2_X1 U6088 ( .A1(n4894), .A2(n4900), .ZN(n4493) );
  NAND2_X1 U6089 ( .A1(n10032), .A2(n9620), .ZN(n4494) );
  INV_X1 U6090 ( .A(n7994), .ZN(n4739) );
  AND2_X1 U6091 ( .A1(n7993), .A2(n8624), .ZN(n7994) );
  NAND2_X1 U6092 ( .A1(n9563), .A2(n9929), .ZN(n4495) );
  AND2_X1 U6093 ( .A1(n5913), .A2(n5912), .ZN(n4496) );
  NAND2_X1 U6094 ( .A1(n7052), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4497) );
  XOR2_X1 U6095 ( .A(n5321), .B(n5743), .Z(n4498) );
  NAND2_X1 U6096 ( .A1(n8134), .A2(n4440), .ZN(n4755) );
  INV_X1 U6097 ( .A(n5587), .ZN(n5610) );
  NAND2_X1 U6098 ( .A1(n5351), .A2(n5350), .ZN(n4499) );
  NAND2_X1 U6099 ( .A1(n7893), .A2(n7892), .ZN(n7915) );
  NAND2_X1 U6100 ( .A1(n5707), .A2(n5706), .ZN(n9810) );
  INV_X1 U6101 ( .A(n9810), .ZN(n4724) );
  INV_X1 U6102 ( .A(n9297), .ZN(n4584) );
  OR2_X1 U6103 ( .A1(n8695), .A2(n8696), .ZN(n8679) );
  NOR2_X1 U6104 ( .A1(n7715), .A2(n7714), .ZN(n7713) );
  INV_X1 U6105 ( .A(n5669), .ZN(n4582) );
  NOR2_X1 U6106 ( .A1(n6040), .A2(n5903), .ZN(n6126) );
  INV_X1 U6107 ( .A(n8285), .ZN(n8312) );
  XOR2_X1 U6108 ( .A(n5370), .B(SI_10_), .Z(n4500) );
  XOR2_X1 U6109 ( .A(n5485), .B(SI_15_), .Z(n4501) );
  OAI21_X1 U6110 ( .B1(n9175), .B2(n4592), .A(n4590), .ZN(n9315) );
  NAND2_X1 U6111 ( .A1(n4651), .A2(n6303), .ZN(n7874) );
  NAND2_X1 U6112 ( .A1(n7942), .A2(n6307), .ZN(n8705) );
  NAND2_X1 U6113 ( .A1(n6309), .A2(n6308), .ZN(n8672) );
  NAND2_X1 U6114 ( .A1(n4595), .A2(n4596), .ZN(n9255) );
  NAND2_X1 U6115 ( .A1(n4609), .A2(n4610), .ZN(n9223) );
  NOR2_X1 U6116 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5402) );
  XOR2_X1 U6117 ( .A(n5580), .B(SI_18_), .Z(n4502) );
  INV_X1 U6118 ( .A(n10269), .ZN(n7038) );
  AND2_X1 U6119 ( .A1(n6029), .A2(n6019), .ZN(n10269) );
  INV_X1 U6120 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5845) );
  OR2_X1 U6121 ( .A1(n7551), .A2(n10382), .ZN(n4503) );
  NAND2_X1 U6122 ( .A1(n9858), .A2(n4727), .ZN(n4728) );
  NOR2_X1 U6123 ( .A1(n7833), .A2(n7832), .ZN(n4504) );
  AND4_X1 U6124 ( .A1(n6181), .A2(n6180), .A3(n6179), .A4(n6178), .ZN(n8662)
         );
  AND2_X1 U6125 ( .A1(n8679), .A2(n6163), .ZN(n4505) );
  INV_X1 U6126 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4909) );
  INV_X1 U6127 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4550) );
  NAND2_X1 U6128 ( .A1(n7342), .A2(n9457), .ZN(n4506) );
  AND2_X1 U6129 ( .A1(n9306), .A2(n9307), .ZN(n4507) );
  AND2_X1 U6130 ( .A1(n7639), .A2(n9635), .ZN(n9488) );
  INV_X1 U6131 ( .A(n9488), .ZN(n9396) );
  AND2_X1 U6132 ( .A1(n10011), .A2(n9632), .ZN(n4508) );
  AND2_X1 U6133 ( .A1(n4869), .A2(n4868), .ZN(n4509) );
  INV_X1 U6134 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5000) );
  AND2_X1 U6135 ( .A1(n6376), .A2(n9158), .ZN(n4510) );
  AND2_X1 U6136 ( .A1(n6126), .A2(n5905), .ZN(n6149) );
  AND2_X1 U6137 ( .A1(n5629), .A2(n5628), .ZN(n4511) );
  AND2_X1 U6138 ( .A1(n9911), .A2(n9630), .ZN(n4512) );
  OR2_X1 U6139 ( .A1(n4977), .A2(n7713), .ZN(n4513) );
  AND2_X1 U6140 ( .A1(n4713), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4514) );
  NOR2_X1 U6141 ( .A1(n5423), .A2(n5422), .ZN(n4515) );
  AND3_X2 U6142 ( .A1(n6490), .A2(n7080), .A3(n6489), .ZN(n10223) );
  NAND2_X1 U6143 ( .A1(n7082), .A2(n9774), .ZN(n9916) );
  INV_X1 U6144 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6099) );
  NAND2_X1 U6145 ( .A1(n4661), .A2(n6287), .ZN(n7369) );
  AND2_X1 U6146 ( .A1(n4600), .A2(n5237), .ZN(n4516) );
  XNOR2_X1 U6147 ( .A(n6344), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U6148 ( .A1(n7216), .A2(n7215), .ZN(n7388) );
  AND2_X1 U6149 ( .A1(n5556), .A2(n5555), .ZN(n4517) );
  NOR2_X1 U6150 ( .A1(n7006), .A2(n7007), .ZN(n4518) );
  NAND2_X1 U6151 ( .A1(n7661), .A2(n4451), .ZN(n4723) );
  NOR2_X1 U6152 ( .A1(n7305), .A2(n7304), .ZN(n4519) );
  AND2_X1 U6153 ( .A1(n4984), .A2(n5264), .ZN(n4520) );
  NAND2_X1 U6154 ( .A1(n6338), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6371) );
  NAND2_X1 U6155 ( .A1(n8451), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4521) );
  NAND2_X1 U6156 ( .A1(n4960), .A2(n4958), .ZN(n5237) );
  AND2_X1 U6157 ( .A1(n5850), .A2(n9705), .ZN(n9533) );
  AND2_X1 U6158 ( .A1(n6901), .A2(n6932), .ZN(n6903) );
  NOR2_X1 U6159 ( .A1(n10265), .A2(n7032), .ZN(n4522) );
  OR2_X1 U6160 ( .A1(n6727), .A2(n6664), .ZN(n10293) );
  INV_X1 U6161 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n4704) );
  AND2_X1 U6162 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n4523) );
  AND2_X1 U6163 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_U3151), .ZN(n4524) );
  INV_X1 U6164 ( .A(n7300), .ZN(n9705) );
  XNOR2_X1 U6165 ( .A(n4577), .B(n5074), .ZN(n7300) );
  NAND2_X1 U6166 ( .A1(n5072), .A2(n5075), .ZN(n9605) );
  INV_X1 U6167 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n4709) );
  INV_X1 U6168 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n4551) );
  NOR2_X1 U6169 ( .A1(n4811), .A2(n4808), .ZN(n4807) );
  NAND2_X1 U6170 ( .A1(n9603), .A2(n9705), .ZN(n4781) );
  NAND2_X1 U6171 ( .A1(n4781), .A2(n4779), .ZN(n4778) );
  AOI21_X1 U6172 ( .B1(n4830), .B2(n4828), .A(n4827), .ZN(n4826) );
  NAND2_X1 U6173 ( .A1(n4810), .A2(n4807), .ZN(n9599) );
  NAND2_X1 U6174 ( .A1(n5139), .A2(n4877), .ZN(n5193) );
  AOI21_X1 U6175 ( .B1(n9538), .B2(n9537), .A(n4780), .ZN(n4779) );
  NOR2_X1 U6176 ( .A1(n4427), .A2(n4484), .ZN(n4544) );
  NOR2_X1 U6177 ( .A1(n8316), .A2(n8315), .ZN(n8320) );
  NOR2_X1 U6178 ( .A1(n8314), .A2(n4489), .ZN(n8308) );
  AOI21_X1 U6179 ( .B1(n8292), .B2(n4540), .A(n4539), .ZN(n4538) );
  NOR2_X1 U6180 ( .A1(n8314), .A2(n5034), .ZN(n8304) );
  AOI21_X1 U6181 ( .B1(n8318), .B2(n8317), .A(n6332), .ZN(n4943) );
  AOI21_X1 U6182 ( .B1(n4940), .B2(n4934), .A(n4487), .ZN(n8374) );
  OAI21_X1 U6183 ( .B1(n10291), .B2(n4528), .A(n4527), .ZN(n10094) );
  NAND2_X1 U6184 ( .A1(n7032), .A2(n4537), .ZN(n4535) );
  INV_X1 U6185 ( .A(n7033), .ZN(n4537) );
  NAND2_X1 U6186 ( .A1(n6714), .A2(n6761), .ZN(n6715) );
  NAND2_X1 U6187 ( .A1(n6763), .A2(n6761), .ZN(n6759) );
  NAND2_X1 U6188 ( .A1(n5934), .A2(n5897), .ZN(n5965) );
  AOI21_X2 U6189 ( .B1(n5193), .B2(n5192), .A(n5191), .ZN(n5209) );
  NAND3_X1 U6190 ( .A1(n4906), .A2(n4550), .A3(n4907), .ZN(n4549) );
  INV_X1 U6191 ( .A(n5137), .ZN(n5135) );
  NAND3_X1 U6192 ( .A1(n4911), .A2(n4910), .A3(n4551), .ZN(n4548) );
  NAND2_X1 U6193 ( .A1(n6946), .A2(n9544), .ZN(n6945) );
  AND3_X2 U6194 ( .A1(n4409), .A2(n5215), .A3(n5026), .ZN(n4554) );
  OAI21_X1 U6195 ( .B1(n7696), .B2(n4560), .A(n4558), .ZN(n9919) );
  NAND2_X1 U6196 ( .A1(n4957), .A2(n4583), .ZN(n4579) );
  NAND2_X1 U6197 ( .A1(n4579), .A2(n4580), .ZN(n9186) );
  NAND2_X1 U6198 ( .A1(n5670), .A2(n5669), .ZN(n9189) );
  NAND2_X1 U6199 ( .A1(n5670), .A2(n4581), .ZN(n4580) );
  NOR2_X1 U6200 ( .A1(n9188), .A2(n4584), .ZN(n4583) );
  NAND2_X1 U6201 ( .A1(n9175), .A2(n4588), .ZN(n4587) );
  NAND3_X1 U6202 ( .A1(n4600), .A2(n4982), .A3(n5237), .ZN(n4601) );
  NAND3_X1 U6203 ( .A1(n4985), .A2(n5265), .A3(n4601), .ZN(n7433) );
  NAND2_X1 U6204 ( .A1(n5076), .A2(n9613), .ZN(n4602) );
  OAI21_X1 U6205 ( .B1(n9195), .B2(n4606), .A(n4604), .ZN(n9287) );
  INV_X1 U6206 ( .A(n7340), .ZN(n4841) );
  INV_X1 U6207 ( .A(n4617), .ZN(n4620) );
  NAND2_X1 U6208 ( .A1(n4770), .A2(n4769), .ZN(n9422) );
  INV_X1 U6209 ( .A(n6434), .ZN(n4628) );
  OAI21_X2 U6210 ( .B1(n9895), .B2(n4636), .A(n4633), .ZN(n9835) );
  NAND2_X1 U6211 ( .A1(n5946), .A2(n4642), .ZN(n4641) );
  NAND2_X2 U6212 ( .A1(n6331), .A2(n6329), .ZN(n5946) );
  OR2_X1 U6213 ( .A1(n7940), .A2(n4646), .ZN(n4643) );
  NAND2_X1 U6214 ( .A1(n4643), .A2(n4644), .ZN(n8689) );
  NAND2_X1 U6215 ( .A1(n7807), .A2(n7894), .ZN(n4651) );
  INV_X1 U6216 ( .A(n6287), .ZN(n4652) );
  NAND2_X1 U6217 ( .A1(n6286), .A2(n6285), .ZN(n7242) );
  INV_X1 U6218 ( .A(n6309), .ZN(n4665) );
  NAND2_X1 U6219 ( .A1(n6337), .A2(n8722), .ZN(n4678) );
  NAND2_X1 U6220 ( .A1(n4678), .A2(n4677), .ZN(n6488) );
  AND2_X1 U6221 ( .A1(n4678), .A2(n4676), .ZN(n8551) );
  NOR2_X2 U6222 ( .A1(n6336), .A2(n4446), .ZN(n4677) );
  NAND2_X1 U6223 ( .A1(n8612), .A2(n4682), .ZN(n4681) );
  OR2_X1 U6224 ( .A1(n8612), .A2(n6314), .ZN(n4691) );
  NAND3_X1 U6225 ( .A1(n4684), .A2(n6314), .A3(n8588), .ZN(n4680) );
  INV_X1 U6226 ( .A(n6040), .ZN(n4693) );
  NOR2_X1 U6227 ( .A1(n4692), .A2(n5903), .ZN(n4694) );
  NAND4_X1 U6228 ( .A1(n4950), .A2(n4696), .A3(n4695), .A4(n4693), .ZN(n5928)
         );
  NAND2_X1 U6229 ( .A1(n6766), .A2(n9025), .ZN(n4697) );
  NAND2_X1 U6230 ( .A1(n6706), .A2(n6766), .ZN(n4698) );
  OAI21_X1 U6231 ( .B1(n7049), .B2(n10248), .A(n4497), .ZN(n4706) );
  OAI21_X1 U6232 ( .B1(n6786), .B2(n4708), .A(n4707), .ZN(n4710) );
  AOI21_X1 U6233 ( .B1(n4709), .B2(n7049), .A(n10248), .ZN(n4707) );
  INV_X1 U6234 ( .A(n7049), .ZN(n4708) );
  INV_X1 U6235 ( .A(n4710), .ZN(n10247) );
  NAND2_X1 U6236 ( .A1(n7563), .A2(n4514), .ZN(n4712) );
  INV_X1 U6237 ( .A(n7835), .ZN(n4713) );
  NAND2_X2 U6238 ( .A1(n5106), .A2(n5105), .ZN(n6977) );
  NAND2_X1 U6239 ( .A1(n9791), .A2(n4718), .ZN(n9719) );
  NAND2_X1 U6240 ( .A1(n9791), .A2(n4721), .ZN(n9757) );
  INV_X1 U6241 ( .A(n4723), .ZN(n7697) );
  INV_X1 U6242 ( .A(n4728), .ZN(n9841) );
  NAND2_X1 U6243 ( .A1(n4729), .A2(n7015), .ZN(n7016) );
  OAI21_X1 U6244 ( .B1(n6934), .B2(n6935), .A(n4729), .ZN(n6936) );
  NAND2_X1 U6245 ( .A1(n6934), .A2(n6935), .ZN(n4729) );
  OAI21_X2 U6246 ( .B1(n8087), .B2(n4732), .A(n4730), .ZN(n7998) );
  NAND2_X1 U6247 ( .A1(n4735), .A2(n4736), .ZN(n8093) );
  INV_X1 U6248 ( .A(n8094), .ZN(n4734) );
  OAI21_X1 U6249 ( .B1(n8087), .B2(n8086), .A(n4740), .ZN(n8047) );
  INV_X1 U6250 ( .A(n8048), .ZN(n4738) );
  NAND2_X1 U6251 ( .A1(n4743), .A2(n8007), .ZN(n8023) );
  NAND2_X1 U6252 ( .A1(n8134), .A2(n4745), .ZN(n4744) );
  NAND2_X2 U6253 ( .A1(n4766), .A2(n4765), .ZN(n7739) );
  NAND2_X1 U6254 ( .A1(n7485), .A2(n4763), .ZN(n4766) );
  NOR2_X1 U6255 ( .A1(n4767), .A2(n7486), .ZN(n4763) );
  CLKBUF_X1 U6256 ( .A(n4766), .Z(n4764) );
  NAND2_X1 U6257 ( .A1(n6933), .A2(n6932), .ZN(n6934) );
  NAND2_X4 U6258 ( .A1(n9358), .A2(n5212), .ZN(n5587) );
  NAND2_X4 U6259 ( .A1(n5856), .A2(n6554), .ZN(n9358) );
  OR2_X1 U6260 ( .A1(n5587), .A2(n4909), .ZN(n5106) );
  OAI21_X1 U6261 ( .B1(n6999), .B2(n6423), .A(n6971), .ZN(n6973) );
  NAND2_X1 U6262 ( .A1(n6999), .A2(n6423), .ZN(n6971) );
  AND2_X1 U6263 ( .A1(n6970), .A2(n6423), .ZN(n4771) );
  NAND2_X1 U6264 ( .A1(n4776), .A2(n4775), .ZN(n9485) );
  NOR2_X1 U6265 ( .A1(n4784), .A2(n4783), .ZN(n4782) );
  INV_X1 U6266 ( .A(n9440), .ZN(n4793) );
  NAND2_X1 U6267 ( .A1(n4795), .A2(n4794), .ZN(n9445) );
  NAND4_X1 U6268 ( .A1(n4409), .A2(n4799), .A3(n4800), .A4(n4492), .ZN(n5093)
         );
  NAND2_X1 U6269 ( .A1(n9532), .A2(n4488), .ZN(n4810) );
  NAND2_X1 U6270 ( .A1(n4818), .A2(n9534), .ZN(n4817) );
  NAND3_X1 U6271 ( .A1(n9576), .A2(n4480), .A3(n4824), .ZN(n4823) );
  AOI21_X1 U6272 ( .B1(n4837), .B2(n9524), .A(n4491), .ZN(n4830) );
  AND2_X1 U6273 ( .A1(n9525), .A2(n9528), .ZN(n4837) );
  NAND2_X1 U6274 ( .A1(n5267), .A2(n5266), .ZN(n4838) );
  NAND2_X1 U6275 ( .A1(n5240), .A2(n5239), .ZN(n4839) );
  NAND2_X1 U6276 ( .A1(n5209), .A2(SI_4_), .ZN(n5210) );
  OR2_X2 U6277 ( .A1(n9893), .A2(n9894), .ZN(n9895) );
  OAI21_X1 U6278 ( .B1(n9766), .B2(n9571), .A(n4844), .ZN(n9735) );
  NAND2_X1 U6279 ( .A1(n9766), .A2(n9518), .ZN(n9750) );
  INV_X1 U6280 ( .A(n4842), .ZN(n6442) );
  INV_X1 U6281 ( .A(n7852), .ZN(n4846) );
  OAI21_X1 U6282 ( .B1(n4846), .B2(n4495), .A(n4847), .ZN(n9905) );
  INV_X1 U6283 ( .A(n9495), .ZN(n4849) );
  NAND2_X1 U6284 ( .A1(n6451), .A2(n4853), .ZN(n4850) );
  NAND2_X1 U6285 ( .A1(n4850), .A2(n4851), .ZN(P1_U3551) );
  NAND2_X1 U6286 ( .A1(n6451), .A2(n9931), .ZN(n4857) );
  XNOR2_X1 U6287 ( .A(n8424), .B(n8438), .ZN(n8402) );
  NAND2_X1 U6288 ( .A1(n4871), .A2(n4872), .ZN(n7552) );
  NAND3_X1 U6289 ( .A1(n4871), .A2(n4872), .A3(n4503), .ZN(n7553) );
  NAND2_X1 U6290 ( .A1(n10224), .A2(n6712), .ZN(n6713) );
  OR2_X1 U6291 ( .A1(n5139), .A2(n4877), .ZN(n5140) );
  NAND2_X1 U6292 ( .A1(n5326), .A2(n4881), .ZN(n4880) );
  NAND2_X1 U6293 ( .A1(n5325), .A2(n5324), .ZN(n4888) );
  NAND2_X1 U6294 ( .A1(n5452), .A2(n4493), .ZN(n4893) );
  NAND2_X1 U6295 ( .A1(n5452), .A2(n4900), .ZN(n4890) );
  NAND2_X1 U6296 ( .A1(n5452), .A2(n5451), .ZN(n5484) );
  INV_X1 U6297 ( .A(n5451), .ZN(n4901) );
  NAND3_X1 U6298 ( .A1(n4904), .A2(n4903), .A3(n4902), .ZN(n5097) );
  NAND3_X1 U6299 ( .A1(n4905), .A2(n4908), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4902) );
  NAND3_X1 U6300 ( .A1(n4906), .A2(n4907), .A3(P2_DATAO_REG_1__SCAN_IN), .ZN(
        n4903) );
  NAND3_X1 U6301 ( .A1(n4911), .A2(P1_DATAO_REG_1__SCAN_IN), .A3(n4910), .ZN(
        n4904) );
  NAND2_X1 U6302 ( .A1(n5582), .A2(n4916), .ZN(n4912) );
  OAI21_X1 U6303 ( .B1(n5582), .B2(n4918), .A(n5581), .ZN(n5609) );
  NAND2_X1 U6304 ( .A1(n4912), .A2(n4913), .ZN(n5630) );
  NAND2_X1 U6305 ( .A1(n5976), .A2(n8345), .ZN(n7253) );
  NAND2_X1 U6306 ( .A1(n4926), .A2(n4924), .ZN(n8599) );
  NAND2_X1 U6307 ( .A1(n4927), .A2(n4490), .ZN(n7686) );
  NAND2_X1 U6308 ( .A1(n8695), .A2(n6163), .ZN(n4930) );
  INV_X1 U6309 ( .A(n8222), .ZN(n4932) );
  NAND2_X1 U6310 ( .A1(n5911), .A2(n4933), .ZN(n5915) );
  AOI21_X1 U6311 ( .B1(n4939), .B2(n4486), .A(n4936), .ZN(n4935) );
  NAND2_X1 U6312 ( .A1(n8335), .A2(n8334), .ZN(n4939) );
  OAI21_X1 U6313 ( .B1(n4943), .B2(n4941), .A(n8329), .ZN(n4940) );
  OAI21_X1 U6314 ( .B1(n8320), .B2(n4942), .A(n8331), .ZN(n4941) );
  NAND2_X1 U6315 ( .A1(n8319), .A2(n6332), .ZN(n4942) );
  NAND2_X1 U6316 ( .A1(n8579), .A2(n4947), .ZN(n4944) );
  INV_X1 U6317 ( .A(n8293), .ZN(n4949) );
  NAND2_X1 U6318 ( .A1(n8579), .A2(n8578), .ZN(n8756) );
  AND2_X1 U6319 ( .A1(n5202), .A2(n6977), .ZN(n4954) );
  OAI21_X1 U6320 ( .B1(n5107), .B2(n5202), .A(n4952), .ZN(n4955) );
  NAND2_X1 U6321 ( .A1(n5107), .A2(n5820), .ZN(n4956) );
  INV_X2 U6322 ( .A(n5202), .ZN(n5820) );
  NAND2_X1 U6323 ( .A1(n6847), .A2(n4961), .ZN(n4960) );
  NAND2_X1 U6324 ( .A1(n6847), .A2(n5183), .ZN(n7006) );
  NOR2_X1 U6325 ( .A1(n7007), .A2(n4962), .ZN(n4961) );
  INV_X1 U6326 ( .A(n5183), .ZN(n4962) );
  OAI21_X1 U6327 ( .B1(n9315), .B2(n9316), .A(n9317), .ZN(n9206) );
  NAND2_X1 U6328 ( .A1(n6468), .A2(n4973), .ZN(n4971) );
  NAND2_X1 U6329 ( .A1(n4971), .A2(n4970), .ZN(P1_U3214) );
  NAND2_X1 U6330 ( .A1(n6465), .A2(n4441), .ZN(n6469) );
  OAI211_X1 U6331 ( .C1(n7715), .C2(n4979), .A(n4978), .B(n4976), .ZN(n5367)
         );
  NAND2_X1 U6332 ( .A1(n7177), .A2(n5237), .ZN(n4984) );
  NAND3_X1 U6333 ( .A1(n5112), .A2(n5127), .A3(n6837), .ZN(n6819) );
  NAND2_X1 U6334 ( .A1(n4989), .A2(n6820), .ZN(n6823) );
  NAND2_X1 U6335 ( .A1(n6819), .A2(n5127), .ZN(n4989) );
  AND2_X1 U6336 ( .A1(n5112), .A2(n5127), .ZN(n6836) );
  NAND2_X1 U6337 ( .A1(n7261), .A2(n4992), .ZN(n4991) );
  AND2_X1 U6338 ( .A1(n10083), .A2(n4997), .ZN(n4996) );
  INV_X1 U6339 ( .A(n10083), .ZN(n5062) );
  NAND2_X1 U6340 ( .A1(n9807), .A2(n4483), .ZN(n5005) );
  NAND3_X1 U6341 ( .A1(n5006), .A2(n5008), .A3(n9571), .ZN(n5004) );
  NAND2_X1 U6342 ( .A1(n5215), .A2(n5027), .ZN(n5491) );
  NAND2_X1 U6343 ( .A1(n8148), .A2(n8285), .ZN(n8151) );
  OR2_X1 U6344 ( .A1(n6415), .A2(n6416), .ZN(n6418) );
  AND2_X1 U6345 ( .A1(n9502), .A2(n9501), .ZN(n9509) );
  INV_X1 U6346 ( .A(n9827), .ZN(n10050) );
  XNOR2_X1 U6347 ( .A(n5927), .B(n5926), .ZN(n6329) );
  XNOR2_X1 U6348 ( .A(n6264), .B(n6263), .ZN(n7908) );
  NAND2_X1 U6349 ( .A1(n5970), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5924) );
  OAI21_X2 U6350 ( .B1(n6415), .B2(n6004), .A(n6269), .ZN(n6376) );
  NAND2_X1 U6351 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  INV_X1 U6352 ( .A(n5237), .ZN(n5238) );
  INV_X1 U6353 ( .A(n6423), .ZN(n6381) );
  XNOR2_X1 U6354 ( .A(n6380), .B(n6977), .ZN(n6423) );
  AOI22_X1 U6355 ( .A1(n6380), .A2(n5745), .B1(n5236), .B2(n6977), .ZN(n5110)
         );
  BUF_X4 U6356 ( .A(n5970), .Z(n6271) );
  AND2_X1 U6357 ( .A1(n5032), .A2(n6464), .ZN(n5028) );
  AND2_X1 U6358 ( .A1(n6377), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5029) );
  INV_X1 U6359 ( .A(n10384), .ZN(n6377) );
  NAND2_X2 U6360 ( .A1(n6926), .A2(n8606), .ZN(n10317) );
  AND2_X1 U6361 ( .A1(n6486), .A2(n6485), .ZN(n10365) );
  AND2_X1 U6362 ( .A1(n6376), .A2(n9084), .ZN(n5030) );
  OR2_X1 U6363 ( .A1(n6491), .A2(n10067), .ZN(n5032) );
  AND2_X1 U6364 ( .A1(n5352), .A2(n5329), .ZN(n5033) );
  INV_X1 U6365 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5897) );
  INV_X1 U6366 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5083) );
  AND2_X1 U6367 ( .A1(n8306), .A2(n8569), .ZN(n5034) );
  AND2_X1 U6368 ( .A1(n8149), .A2(n6332), .ZN(n5035) );
  AND2_X1 U6369 ( .A1(n5875), .A2(n9329), .ZN(n5036) );
  NAND2_X1 U6370 ( .A1(n9232), .A2(n9233), .ZN(n5882) );
  INV_X1 U6371 ( .A(n8279), .ZN(n8338) );
  OR2_X1 U6372 ( .A1(n8490), .A2(n8489), .ZN(n5037) );
  OR2_X1 U6373 ( .A1(n7551), .A2(n7317), .ZN(n5038) );
  INV_X1 U6374 ( .A(n7834), .ZN(n8414) );
  INV_X1 U6375 ( .A(n10361), .ZN(n6278) );
  AND2_X1 U6376 ( .A1(n7978), .A2(n8242), .ZN(n5039) );
  INV_X1 U6377 ( .A(n10003), .ZN(n6455) );
  NAND2_X1 U6378 ( .A1(n8645), .A2(n8154), .ZN(n8636) );
  NAND2_X1 U6379 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), 
        .ZN(n5040) );
  OR2_X1 U6380 ( .A1(n7193), .A2(n10380), .ZN(n5041) );
  AND2_X1 U6381 ( .A1(n6465), .A2(n9329), .ZN(n5043) );
  INV_X1 U6382 ( .A(n10001), .ZN(n6494) );
  NAND2_X1 U6383 ( .A1(n5864), .A2(n5852), .ZN(n9354) );
  INV_X1 U6384 ( .A(n9354), .ZN(n9329) );
  NAND2_X1 U6385 ( .A1(n8334), .A2(n5035), .ZN(n8150) );
  INV_X1 U6386 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5908) );
  INV_X1 U6387 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5899) );
  NAND2_X1 U6388 ( .A1(n6711), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6698) );
  NAND2_X1 U6389 ( .A1(n5294), .A2(n5293), .ZN(n5295) );
  INV_X1 U6390 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5312) );
  INV_X1 U6391 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6392 ( .A1(n8000), .A2(n8591), .ZN(n8001) );
  OR2_X1 U6393 ( .A1(n6703), .A2(n6721), .ZN(n6704) );
  NAND2_X1 U6394 ( .A1(n7029), .A2(n7028), .ZN(n7030) );
  NAND2_X1 U6395 ( .A1(n8176), .A2(n8170), .ZN(n6279) );
  INV_X1 U6396 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6340) );
  OR2_X1 U6397 ( .A1(n5647), .A2(n5646), .ZN(n5648) );
  OR2_X1 U6398 ( .A1(n5313), .A2(n5312), .ZN(n5339) );
  INV_X1 U6399 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n7582) );
  OR2_X1 U6400 ( .A1(n5614), .A2(n5613), .ZN(n5635) );
  INV_X1 U6401 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8999) );
  AND2_X1 U6402 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5223) );
  NAND2_X1 U6403 ( .A1(n9647), .A2(n6975), .ZN(n6967) );
  INV_X1 U6404 ( .A(SI_26_), .ZN(n8930) );
  INV_X1 U6405 ( .A(SI_16_), .ZN(n9021) );
  INV_X1 U6406 ( .A(SI_9_), .ZN(n8774) );
  AND2_X1 U6407 ( .A1(n6185), .A2(n6184), .ZN(n6197) );
  NAND2_X1 U6408 ( .A1(n6903), .A2(n6904), .ZN(n6933) );
  INV_X1 U6409 ( .A(n7561), .ZN(n7319) );
  INV_X1 U6410 ( .A(n8491), .ZN(n8454) );
  NAND2_X1 U6411 ( .A1(n6345), .A2(n5929), .ZN(n5930) );
  NOR2_X1 U6412 ( .A1(n6078), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6090) );
  OR2_X1 U6413 ( .A1(n6351), .A2(n6368), .ZN(n6481) );
  NAND2_X1 U6414 ( .A1(n8557), .A2(n8719), .ZN(n8558) );
  AND2_X1 U6415 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  OR2_X1 U6416 ( .A1(n6483), .A2(n6482), .ZN(n6872) );
  INV_X1 U6417 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5907) );
  OR2_X1 U6418 ( .A1(n6074), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n6085) );
  OR2_X1 U6419 ( .A1(n5681), .A2(n9191), .ZN(n5736) );
  OAI21_X1 U6420 ( .B1(n6416), .B2(n6511), .A(n5103), .ZN(n5104) );
  AND2_X1 U6421 ( .A1(n5566), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5591) );
  OR2_X1 U6422 ( .A1(n5736), .A2(n5735), .ZN(n5756) );
  NAND2_X1 U6423 ( .A1(n5591), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5614) );
  NOR2_X1 U6424 ( .A1(n5756), .A2(n5889), .ZN(n5783) );
  INV_X1 U6425 ( .A(n9629), .ZN(n9280) );
  OR2_X1 U6426 ( .A1(n5436), .A2(n8999), .ZN(n5466) );
  INV_X1 U6427 ( .A(n6958), .ZN(n9541) );
  INV_X1 U6428 ( .A(n10204), .ZN(n6453) );
  INV_X1 U6429 ( .A(n6967), .ZN(n6970) );
  INV_X1 U6430 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5058) );
  INV_X1 U6431 ( .A(SI_15_), .ZN(n9019) );
  OR2_X1 U6432 ( .A1(n8062), .A2(n8691), .ZN(n7985) );
  OR2_X1 U6433 ( .A1(n6010), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6023) );
  OR2_X1 U6434 ( .A1(n6067), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6078) );
  OR2_X1 U6435 ( .A1(n10359), .A2(n6878), .ZN(n6924) );
  AND3_X1 U6436 ( .A1(n6887), .A2(n6324), .A3(n10359), .ZN(n7775) );
  NOR2_X1 U6437 ( .A1(n6872), .A2(n6925), .ZN(n6890) );
  OAI21_X1 U6438 ( .B1(n5934), .B2(n5957), .A(n5956), .ZN(n5958) );
  INV_X1 U6439 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9191) );
  INV_X1 U6440 ( .A(n9337), .ZN(n9349) );
  AND2_X1 U6441 ( .A1(n6533), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6498) );
  NOR2_X1 U6442 ( .A1(n9720), .A2(n9719), .ZN(n9718) );
  INV_X1 U6443 ( .A(n9571), .ZN(n9755) );
  INV_X1 U6444 ( .A(n9568), .ZN(n9823) );
  INV_X1 U6445 ( .A(n9858), .ZN(n9877) );
  INV_X1 U6446 ( .A(n7858), .ZN(n9923) );
  NAND2_X1 U6447 ( .A1(n4769), .A2(n9428), .ZN(n6983) );
  AND2_X1 U6448 ( .A1(n5856), .A2(n9595), .ZN(n9321) );
  INV_X1 U6449 ( .A(n9557), .ZN(n7512) );
  INV_X1 U6450 ( .A(n7151), .ZN(n7273) );
  INV_X1 U6451 ( .A(n9931), .ZN(n9906) );
  INV_X1 U6452 ( .A(n7674), .ZN(n10208) );
  AND2_X1 U6453 ( .A1(n5773), .A2(n5753), .ZN(n5771) );
  AND2_X1 U6454 ( .A1(n5559), .A2(n5539), .ZN(n5557) );
  OR2_X1 U6455 ( .A1(n5405), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5430) );
  INV_X1 U6456 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n9036) );
  INV_X1 U6457 ( .A(n8127), .ZN(n8137) );
  NOR2_X1 U6458 ( .A1(n7979), .A2(n5039), .ZN(n8136) );
  NAND2_X1 U6459 ( .A1(n6352), .A2(n6370), .ZN(n6866) );
  INV_X1 U6460 ( .A(n8477), .ZN(n8480) );
  OR2_X1 U6461 ( .A1(n6925), .A2(n6924), .ZN(n8606) );
  INV_X1 U6462 ( .A(n8676), .ZN(n8719) );
  AND2_X1 U6463 ( .A1(n7686), .A2(n7594), .ZN(n10347) );
  INV_X1 U6464 ( .A(n10331), .ZN(n7257) );
  INV_X1 U6465 ( .A(n8606), .ZN(n10314) );
  INV_X1 U6466 ( .A(n7467), .ZN(n7470) );
  AND3_X1 U6467 ( .A1(n6483), .A2(n6916), .A3(n6924), .ZN(n6375) );
  OAI21_X1 U6468 ( .B1(n8656), .B2(n8159), .A(n8267), .ZN(n8645) );
  AND2_X1 U6469 ( .A1(n8232), .A2(n8233), .ZN(n8231) );
  OR2_X1 U6470 ( .A1(n7775), .A2(n6278), .ZN(n9071) );
  AND2_X1 U6471 ( .A1(n6105), .A2(n6115), .ZN(n8463) );
  AND2_X1 U6472 ( .A1(n4525), .A2(P2_U3151), .ZN(n9166) );
  AND2_X1 U6473 ( .A1(n5791), .A2(n5790), .ZN(n6413) );
  AND3_X1 U6474 ( .A1(n5550), .A2(n5549), .A3(n5548), .ZN(n7854) );
  AND2_X1 U6475 ( .A1(n6537), .A2(n6536), .ZN(n6556) );
  INV_X1 U6476 ( .A(n9701), .ZN(n10175) );
  AND2_X1 U6477 ( .A1(n6556), .A2(n6555), .ZN(n10158) );
  AND2_X1 U6478 ( .A1(n9495), .A2(n9478), .ZN(n9929) );
  INV_X1 U6479 ( .A(n9469), .ZN(n9559) );
  NAND2_X1 U6480 ( .A1(n7297), .A2(n7086), .ZN(n9876) );
  NOR2_X1 U6481 ( .A1(n10223), .A2(n6492), .ZN(n6493) );
  AND2_X1 U6482 ( .A1(n5843), .A2(n10073), .ZN(n6489) );
  AND2_X1 U6483 ( .A1(n6456), .A2(n9608), .ZN(n10205) );
  AND2_X1 U6484 ( .A1(n9533), .A2(n9605), .ZN(n7674) );
  AND2_X1 U6485 ( .A1(n7078), .A2(n6462), .ZN(n6490) );
  NAND2_X1 U6486 ( .A1(n5826), .A2(n7868), .ZN(n6457) );
  INV_X1 U6487 ( .A(n7680), .ZN(n5842) );
  AND2_X1 U6488 ( .A1(n5824), .A2(n4430), .ZN(n7680) );
  AND2_X1 U6489 ( .A1(n5430), .A2(n5406), .ZN(n7408) );
  INV_X4 U6490 ( .A(n5212), .ZN(n9356) );
  NOR2_X1 U6491 ( .A1(n4525), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10082) );
  INV_X1 U6492 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9651) );
  OAI21_X1 U6493 ( .B1(n10281), .B2(n8770), .A(n7539), .ZN(n7540) );
  INV_X1 U6494 ( .A(n8141), .ZN(n7495) );
  AND2_X1 U6495 ( .A1(n6863), .A2(n6862), .ZN(n8131) );
  NAND2_X1 U6496 ( .A1(n6261), .A2(n6260), .ZN(n8569) );
  INV_X1 U6497 ( .A(n8663), .ZN(n8692) );
  INV_X1 U6498 ( .A(n8235), .ZN(n8720) );
  INV_X1 U6499 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10281) );
  INV_X2 U6500 ( .A(n10317), .ZN(n8741) );
  OR2_X1 U6501 ( .A1(n6926), .A2(n8731), .ZN(n8699) );
  NOR2_X1 U6502 ( .A1(n5030), .A2(n5029), .ZN(n6378) );
  INV_X1 U6503 ( .A(n9084), .ZN(n9075) );
  NAND2_X1 U6504 ( .A1(n10384), .A2(n9071), .ZN(n9087) );
  AND2_X2 U6505 ( .A1(n6915), .A2(n6375), .ZN(n10384) );
  INV_X1 U6506 ( .A(n8129), .ZN(n9110) );
  OR2_X1 U6507 ( .A1(n10365), .A2(n10359), .ZN(n9147) );
  OR2_X1 U6508 ( .A1(n10365), .A2(n10353), .ZN(n9162) );
  AND3_X1 U6509 ( .A1(n10340), .A2(n10339), .A3(n10338), .ZN(n10375) );
  INV_X2 U6510 ( .A(n10365), .ZN(n10367) );
  AND2_X1 U6511 ( .A1(n6544), .A2(n6351), .ZN(n6587) );
  INV_X1 U6512 ( .A(n6587), .ZN(n6565) );
  INV_X1 U6513 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7604) );
  INV_X1 U6514 ( .A(n6783), .ZN(n6790) );
  AND2_X1 U6515 ( .A1(n6537), .A2(n6535), .ZN(n10155) );
  NAND2_X1 U6516 ( .A1(n6469), .A2(n5854), .ZN(n5880) );
  INV_X1 U6517 ( .A(n5892), .ZN(n5893) );
  AND2_X1 U6518 ( .A1(n5862), .A2(n5861), .ZN(n6885) );
  INV_X1 U6519 ( .A(n9370), .ZN(n9627) );
  INV_X1 U6520 ( .A(n10173), .ZN(n9674) );
  OR2_X1 U6521 ( .A1(n6550), .A2(n9610), .ZN(n9701) );
  INV_X1 U6522 ( .A(n10158), .ZN(n10182) );
  OR2_X1 U6523 ( .A1(n4415), .A2(n7085), .ZN(n7297) );
  NAND2_X1 U6524 ( .A1(n10223), .A2(n10205), .ZN(n10001) );
  INV_X1 U6525 ( .A(n9792), .ZN(n10043) );
  NAND3_X1 U6526 ( .A1(n7081), .A2(n7080), .A3(n6490), .ZN(n10218) );
  INV_X2 U6527 ( .A(n10218), .ZN(n10220) );
  INV_X1 U6528 ( .A(n10202), .ZN(n10201) );
  INV_X1 U6529 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8977) );
  INV_X1 U6530 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7094) );
  INV_X1 U6531 ( .A(n7408), .ZN(n6809) );
  INV_X1 U6532 ( .A(n7656), .ZN(n10085) );
  OAI21_X1 U6533 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n10403), .ZN(n10401) );
  INV_X2 U6534 ( .A(n8399), .ZN(P2_U3893) );
  NAND2_X1 U6535 ( .A1(n6379), .A2(n6378), .ZN(P2_U3488) );
  INV_X2 U6536 ( .A(n9646), .ZN(P1_U3973) );
  NOR2_X1 U6537 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5047) );
  NAND4_X1 U6538 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5050)
         );
  NAND3_X1 U6539 ( .A1(n5402), .A2(n5048), .A3(n5330), .ZN(n5049) );
  NOR2_X1 U6540 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5054) );
  NOR2_X1 U6541 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5053) );
  NOR2_X1 U6542 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5052) );
  INV_X1 U6543 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5055) );
  INV_X1 U6544 ( .A(n5092), .ZN(n5059) );
  NAND2_X1 U6545 ( .A1(n5059), .A2(n5058), .ZN(n10075) );
  NAND2_X1 U6546 ( .A1(n5171), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5066) );
  OR2_X2 U6547 ( .A1(n10079), .A2(n10083), .ZN(n5170) );
  INV_X1 U6548 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5061) );
  OR2_X1 U6549 ( .A1(n5170), .A2(n5061), .ZN(n5065) );
  AND2_X2 U6550 ( .A1(n10079), .A2(n5062), .ZN(n5387) );
  NAND4_X2 U6551 ( .A1(n5066), .A2(n5065), .A3(n5064), .A4(n5063), .ZN(n6380)
         );
  OR2_X2 U6552 ( .A1(n5070), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n5075) );
  NAND2_X1 U6553 ( .A1(n5070), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5071) );
  MUX2_X1 U6554 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5071), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5072) );
  INV_X1 U6555 ( .A(n9611), .ZN(n6421) );
  NAND2_X1 U6556 ( .A1(n5073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U6557 ( .A1(n6421), .A2(n9608), .ZN(n5076) );
  NAND2_X1 U6558 ( .A1(n4430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5077) );
  MUX2_X1 U6559 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5077), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5078) );
  NAND2_X1 U6560 ( .A1(n5078), .A2(n4431), .ZN(n5827) );
  INV_X1 U6561 ( .A(n5827), .ZN(n7725) );
  NAND2_X1 U6562 ( .A1(n4431), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5079) );
  NOR2_X1 U6563 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5082) );
  AOI21_X1 U6564 ( .B1(n4988), .B2(n5082), .A(n10074), .ZN(n5085) );
  NAND2_X1 U6565 ( .A1(n5087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5088) );
  NAND3_X2 U6566 ( .A1(n5092), .A2(n5091), .A3(n5090), .ZN(n5856) );
  NAND2_X1 U6567 ( .A1(n5093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5094) );
  NAND2_X2 U6568 ( .A1(n9358), .A2(n9356), .ZN(n6416) );
  INV_X1 U6569 ( .A(n5097), .ZN(n5096) );
  INV_X1 U6570 ( .A(SI_1_), .ZN(n5095) );
  NAND2_X1 U6571 ( .A1(n5096), .A2(n5095), .ZN(n5098) );
  NAND2_X1 U6572 ( .A1(n5097), .A2(SI_1_), .ZN(n5132) );
  NAND2_X1 U6573 ( .A1(n5098), .A2(n5132), .ZN(n5134) );
  NAND2_X1 U6574 ( .A1(n5101), .A2(SI_0_), .ZN(n5133) );
  XNOR2_X1 U6575 ( .A(n5134), .B(n5133), .ZN(n6511) );
  INV_X1 U6576 ( .A(n9358), .ZN(n5165) );
  NAND2_X1 U6577 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5102) );
  XNOR2_X1 U6578 ( .A(n5102), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6574) );
  NAND2_X1 U6579 ( .A1(n5165), .A2(n6574), .ZN(n5103) );
  INV_X1 U6580 ( .A(n5104), .ZN(n5105) );
  INV_X1 U6581 ( .A(n5110), .ZN(n5109) );
  NAND2_X1 U6582 ( .A1(n6380), .A2(n5236), .ZN(n5107) );
  NAND2_X1 U6583 ( .A1(n5109), .A2(n5108), .ZN(n5112) );
  NAND2_X1 U6584 ( .A1(n5111), .A2(n5110), .ZN(n5127) );
  INV_X1 U6585 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8996) );
  NAND2_X1 U6586 ( .A1(n5387), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5118) );
  OR2_X1 U6587 ( .A1(n5251), .A2(n8996), .ZN(n5117) );
  INV_X1 U6588 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5113) );
  OR2_X1 U6589 ( .A1(n5170), .A2(n5113), .ZN(n5115) );
  NAND2_X1 U6590 ( .A1(n9647), .A2(n5236), .ZN(n5122) );
  INV_X1 U6591 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5121) );
  NAND2_X1 U6592 ( .A1(n9356), .A2(SI_0_), .ZN(n5120) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5119) );
  XNOR2_X1 U6594 ( .A(n5120), .B(n5119), .ZN(n10086) );
  MUX2_X1 U6595 ( .A(n5121), .B(n10086), .S(n9358), .Z(n7104) );
  INV_X1 U6596 ( .A(n7104), .ZN(n6975) );
  OAI211_X1 U6597 ( .C1(n8996), .C2(n6500), .A(n5122), .B(n5126), .ZN(n6735)
         );
  NAND2_X1 U6598 ( .A1(n9647), .A2(n5745), .ZN(n5125) );
  INV_X1 U6599 ( .A(n6500), .ZN(n5123) );
  AOI22_X1 U6600 ( .A1(n6975), .A2(n5236), .B1(n5123), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n5124) );
  NAND2_X1 U6601 ( .A1(n5125), .A2(n5124), .ZN(n6734) );
  AOI22_X1 U6602 ( .A1(n6735), .A2(n6734), .B1(n5820), .B2(n5126), .ZN(n6837)
         );
  INV_X1 U6603 ( .A(n5127), .ZN(n6821) );
  INV_X1 U6604 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5128) );
  INV_X1 U6605 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6830) );
  INV_X1 U6606 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6571) );
  OR2_X1 U6607 ( .A1(n5251), .A2(n6571), .ZN(n5130) );
  NAND2_X1 U6608 ( .A1(n9645), .A2(n5236), .ZN(n5145) );
  NAND2_X1 U6609 ( .A1(n5135), .A2(SI_2_), .ZN(n5189) );
  INV_X1 U6610 ( .A(SI_2_), .ZN(n5136) );
  NAND2_X1 U6611 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  AND2_X1 U6612 ( .A1(n5140), .A2(n5193), .ZN(n5955) );
  INV_X1 U6613 ( .A(n5955), .ZN(n6509) );
  OR2_X1 U6614 ( .A1(n5141), .A2(n10074), .ZN(n5162) );
  XNOR2_X1 U6615 ( .A(n5162), .B(P1_IR_REG_2__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U6616 ( .A1(n5165), .A2(n6740), .ZN(n5142) );
  NAND2_X1 U6617 ( .A1(n5169), .A2(n7140), .ZN(n5144) );
  NAND2_X1 U6618 ( .A1(n5145), .A2(n5144), .ZN(n5146) );
  XNOR2_X1 U6619 ( .A(n5146), .B(n5820), .ZN(n5150) );
  INV_X1 U6620 ( .A(n5150), .ZN(n5148) );
  AOI22_X1 U6621 ( .A1(n9645), .A2(n5745), .B1(n5236), .B2(n7140), .ZN(n5149)
         );
  INV_X1 U6622 ( .A(n5149), .ZN(n5147) );
  NAND2_X1 U6623 ( .A1(n5148), .A2(n5147), .ZN(n5151) );
  NAND2_X1 U6624 ( .A1(n5150), .A2(n5149), .ZN(n5152) );
  NAND2_X1 U6625 ( .A1(n6823), .A2(n5152), .ZN(n6848) );
  INV_X2 U6626 ( .A(n6416), .ZN(n5214) );
  NAND2_X1 U6627 ( .A1(n5193), .A2(n5189), .ZN(n5158) );
  MUX2_X1 U6628 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n5153), .Z(n5154) );
  NAND2_X1 U6629 ( .A1(n5154), .A2(SI_3_), .ZN(n5188) );
  INV_X1 U6630 ( .A(n5154), .ZN(n5156) );
  INV_X1 U6631 ( .A(SI_3_), .ZN(n5155) );
  NAND2_X1 U6632 ( .A1(n5156), .A2(n5155), .ZN(n5190) );
  AND2_X1 U6633 ( .A1(n5188), .A2(n5190), .ZN(n5157) );
  NAND2_X1 U6634 ( .A1(n5158), .A2(n5157), .ZN(n5160) );
  OR2_X1 U6635 ( .A1(n5158), .A2(n5157), .ZN(n5159) );
  AND2_X1 U6636 ( .A1(n5160), .A2(n5159), .ZN(n6504) );
  NAND2_X1 U6637 ( .A1(n5214), .A2(n6504), .ZN(n5168) );
  NAND2_X1 U6638 ( .A1(n5610), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5167) );
  INV_X1 U6639 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6640 ( .A1(n5162), .A2(n5161), .ZN(n5163) );
  NAND2_X1 U6641 ( .A1(n5163), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5164) );
  XNOR2_X1 U6642 ( .A(n5164), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U6643 ( .A1(n5165), .A2(n6604), .ZN(n5166) );
  AND3_X2 U6644 ( .A1(n5168), .A2(n5167), .A3(n5166), .ZN(n7365) );
  NAND2_X1 U6645 ( .A1(n4614), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5175) );
  OR2_X1 U6646 ( .A1(n5129), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5174) );
  INV_X1 U6647 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6594) );
  OR2_X1 U6648 ( .A1(n9364), .A2(n6594), .ZN(n5173) );
  INV_X1 U6649 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6577) );
  OR2_X1 U6650 ( .A1(n5251), .A2(n6577), .ZN(n5172) );
  NAND2_X1 U6651 ( .A1(n6385), .A2(n5236), .ZN(n5176) );
  NAND2_X1 U6652 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6653 ( .A1(n6385), .A2(n5745), .ZN(n5179) );
  OAI21_X1 U6654 ( .B1(n7365), .B2(n5345), .A(n5179), .ZN(n5181) );
  XNOR2_X1 U6655 ( .A(n5180), .B(n5181), .ZN(n6849) );
  NAND2_X1 U6656 ( .A1(n6848), .A2(n6849), .ZN(n6847) );
  INV_X1 U6657 ( .A(n5180), .ZN(n5182) );
  OR2_X1 U6658 ( .A1(n5182), .A2(n5181), .ZN(n5183) );
  INV_X1 U6659 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6516) );
  OR2_X1 U6660 ( .A1(n5184), .A2(n10074), .ZN(n5186) );
  XNOR2_X1 U6661 ( .A(n5186), .B(n5185), .ZN(n9659) );
  OAI22_X1 U6662 ( .A1(n5587), .A2(n6516), .B1(n9358), .B2(n9659), .ZN(n5187)
         );
  INV_X1 U6663 ( .A(n5187), .ZN(n5196) );
  AND2_X1 U6664 ( .A1(n5189), .A2(n5188), .ZN(n5192) );
  MUX2_X1 U6665 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n9356), .Z(n5208) );
  XNOR2_X1 U6666 ( .A(n5208), .B(SI_4_), .ZN(n5194) );
  XNOR2_X1 U6667 ( .A(n5209), .B(n5194), .ZN(n6515) );
  NAND2_X1 U6668 ( .A1(n6515), .A2(n5214), .ZN(n5195) );
  NAND2_X1 U6669 ( .A1(n4614), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5200) );
  INV_X1 U6670 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6596) );
  OR2_X1 U6671 ( .A1(n9364), .A2(n6596), .ZN(n5199) );
  INV_X1 U6672 ( .A(n5223), .ZN(n5225) );
  OAI21_X1 U6673 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(n5225), .ZN(n7108) );
  OR2_X1 U6674 ( .A1(n5129), .A2(n7108), .ZN(n5198) );
  INV_X1 U6675 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6605) );
  OR2_X1 U6676 ( .A1(n5251), .A2(n6605), .ZN(n5197) );
  NAND4_X1 U6677 ( .A1(n5200), .A2(n5199), .A3(n5198), .A4(n5197), .ZN(n9644)
         );
  NAND2_X1 U6678 ( .A1(n9644), .A2(n5236), .ZN(n5201) );
  OAI21_X1 U6679 ( .B1(n7331), .B2(n5600), .A(n5201), .ZN(n5203) );
  XNOR2_X1 U6680 ( .A(n5203), .B(n5743), .ZN(n5206) );
  NAND2_X1 U6681 ( .A1(n9644), .A2(n5745), .ZN(n5204) );
  OAI21_X1 U6682 ( .B1(n7331), .B2(n5345), .A(n5204), .ZN(n5205) );
  XNOR2_X1 U6683 ( .A(n5206), .B(n5205), .ZN(n7007) );
  NAND2_X1 U6684 ( .A1(n5206), .A2(n5205), .ZN(n5207) );
  OAI21_X1 U6685 ( .B1(n5209), .B2(SI_4_), .A(n5208), .ZN(n5211) );
  NAND2_X1 U6686 ( .A1(n5211), .A2(n5210), .ZN(n5240) );
  INV_X1 U6687 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6522) );
  INV_X1 U6688 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6514) );
  MUX2_X1 U6689 ( .A(n6522), .B(n6514), .S(n9356), .Z(n5241) );
  XNOR2_X1 U6690 ( .A(n5241), .B(SI_5_), .ZN(n5239) );
  INV_X1 U6691 ( .A(n5239), .ZN(n5213) );
  XNOR2_X1 U6692 ( .A(n5240), .B(n5213), .ZN(n6513) );
  NAND2_X1 U6693 ( .A1(n6513), .A2(n5214), .ZN(n5219) );
  OR2_X1 U6694 ( .A1(n5215), .A2(n10074), .ZN(n5216) );
  XNOR2_X1 U6695 ( .A(n5216), .B(n5331), .ZN(n6616) );
  OAI22_X1 U6696 ( .A1(n5587), .A2(n6514), .B1(n9358), .B2(n6616), .ZN(n5217)
         );
  INV_X1 U6697 ( .A(n5217), .ZN(n5218) );
  NAND2_X1 U6698 ( .A1(n5219), .A2(n5218), .ZN(n6389) );
  NAND2_X1 U6699 ( .A1(n6389), .A2(n5220), .ZN(n5232) );
  NAND2_X1 U6700 ( .A1(n9360), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5230) );
  INV_X1 U6701 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5222) );
  OR2_X1 U6702 ( .A1(n5170), .A2(n5222), .ZN(n5229) );
  NAND2_X1 U6703 ( .A1(n5223), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5249) );
  INV_X1 U6704 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5224) );
  NAND2_X1 U6705 ( .A1(n5225), .A2(n5224), .ZN(n5226) );
  NAND2_X1 U6706 ( .A1(n5249), .A2(n5226), .ZN(n7179) );
  OR2_X1 U6707 ( .A1(n5129), .A2(n7179), .ZN(n5228) );
  INV_X1 U6708 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7083) );
  OR2_X1 U6709 ( .A1(n9364), .A2(n7083), .ZN(n5227) );
  OR2_X1 U6710 ( .A1(n7153), .A2(n5345), .ZN(n5231) );
  NAND2_X1 U6711 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  XNOR2_X1 U6712 ( .A(n5233), .B(n5743), .ZN(n5234) );
  INV_X1 U6713 ( .A(n7153), .ZN(n9643) );
  AOI22_X1 U6714 ( .A1(n9643), .A2(n5745), .B1(n6389), .B2(n5445), .ZN(n7178)
         );
  INV_X1 U6715 ( .A(n5241), .ZN(n5242) );
  NAND2_X1 U6716 ( .A1(n5242), .A2(SI_5_), .ZN(n5243) );
  INV_X1 U6717 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6526) );
  INV_X1 U6718 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6512) );
  MUX2_X1 U6719 ( .A(n6526), .B(n6512), .S(n9356), .Z(n5268) );
  XNOR2_X1 U6720 ( .A(n5268), .B(SI_6_), .ZN(n5266) );
  XNOR2_X1 U6721 ( .A(n5267), .B(n5266), .ZN(n6525) );
  OR2_X1 U6722 ( .A1(n6525), .A2(n6416), .ZN(n5247) );
  NAND2_X1 U6723 ( .A1(n5215), .A2(n5331), .ZN(n5244) );
  NAND2_X1 U6724 ( .A1(n5244), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5272) );
  XNOR2_X1 U6725 ( .A(n5272), .B(n5332), .ZN(n6649) );
  OAI22_X1 U6726 ( .A1(n5587), .A2(n6512), .B1(n9358), .B2(n6649), .ZN(n5245)
         );
  INV_X1 U6727 ( .A(n5245), .ZN(n5246) );
  NAND2_X1 U6728 ( .A1(n4614), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5255) );
  INV_X1 U6729 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7163) );
  OR2_X1 U6730 ( .A1(n9364), .A2(n7163), .ZN(n5254) );
  NOR2_X1 U6731 ( .A1(n5249), .A2(n5248), .ZN(n5280) );
  INV_X1 U6732 ( .A(n5280), .ZN(n5282) );
  NAND2_X1 U6733 ( .A1(n5249), .A2(n5248), .ZN(n5250) );
  NAND2_X1 U6734 ( .A1(n5282), .A2(n5250), .ZN(n9335) );
  OR2_X1 U6735 ( .A1(n5129), .A2(n9335), .ZN(n5253) );
  INV_X1 U6736 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6627) );
  OR2_X1 U6737 ( .A1(n5251), .A2(n6627), .ZN(n5252) );
  NAND4_X1 U6738 ( .A1(n5255), .A2(n5254), .A3(n5253), .A4(n5252), .ZN(n9642)
         );
  INV_X1 U6739 ( .A(n9642), .ZN(n6391) );
  OAI22_X1 U6740 ( .A1(n7336), .A2(n5600), .B1(n6391), .B2(n5345), .ZN(n5256)
         );
  XNOR2_X1 U6741 ( .A(n5256), .B(n5820), .ZN(n5259) );
  OR2_X1 U6742 ( .A1(n7336), .A2(n5345), .ZN(n5258) );
  NAND2_X1 U6743 ( .A1(n9642), .A2(n5745), .ZN(n5257) );
  AND2_X1 U6744 ( .A1(n5258), .A2(n5257), .ZN(n5260) );
  NAND2_X1 U6745 ( .A1(n5259), .A2(n5260), .ZN(n5265) );
  INV_X1 U6746 ( .A(n5259), .ZN(n5262) );
  INV_X1 U6747 ( .A(n5260), .ZN(n5261) );
  NAND2_X1 U6748 ( .A1(n5262), .A2(n5261), .ZN(n5263) );
  NAND2_X1 U6749 ( .A1(n5265), .A2(n5263), .ZN(n9328) );
  INV_X1 U6750 ( .A(n9328), .ZN(n5264) );
  INV_X1 U6751 ( .A(n5268), .ZN(n5269) );
  NAND2_X1 U6752 ( .A1(n5269), .A2(SI_6_), .ZN(n5270) );
  INV_X1 U6753 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6524) );
  INV_X1 U6754 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6507) );
  MUX2_X1 U6755 ( .A(n6524), .B(n6507), .S(n9356), .Z(n5298) );
  XNOR2_X1 U6756 ( .A(n5298), .B(SI_7_), .ZN(n5296) );
  INV_X1 U6757 ( .A(n5296), .ZN(n5271) );
  XNOR2_X1 U6758 ( .A(n5297), .B(n5271), .ZN(n6506) );
  NAND2_X1 U6759 ( .A1(n6506), .A2(n5214), .ZN(n5278) );
  NAND2_X1 U6760 ( .A1(n5272), .A2(n5332), .ZN(n5273) );
  NAND2_X1 U6761 ( .A1(n5273), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5274) );
  NAND2_X1 U6762 ( .A1(n5274), .A2(n9036), .ZN(n5306) );
  OR2_X1 U6763 ( .A1(n5274), .A2(n9036), .ZN(n5275) );
  NAND2_X1 U6764 ( .A1(n5306), .A2(n5275), .ZN(n6679) );
  OAI22_X1 U6765 ( .A1(n5587), .A2(n6507), .B1(n9358), .B2(n6679), .ZN(n5276)
         );
  INV_X1 U6766 ( .A(n5276), .ZN(n5277) );
  NAND2_X1 U6767 ( .A1(n5278), .A2(n5277), .ZN(n10204) );
  NAND2_X1 U6768 ( .A1(n9360), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5287) );
  INV_X1 U6769 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5279) );
  OR2_X1 U6770 ( .A1(n5170), .A2(n5279), .ZN(n5286) );
  NAND2_X1 U6771 ( .A1(n5280), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5313) );
  INV_X1 U6772 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6773 ( .A1(n5282), .A2(n5281), .ZN(n5283) );
  NAND2_X1 U6774 ( .A1(n5313), .A2(n5283), .ZN(n7439) );
  OR2_X1 U6775 ( .A1(n5129), .A2(n7439), .ZN(n5285) );
  INV_X1 U6776 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7272) );
  OR2_X1 U6777 ( .A1(n9364), .A2(n7272), .ZN(n5284) );
  INV_X1 U6778 ( .A(n7280), .ZN(n9641) );
  AOI22_X1 U6779 ( .A1(n10204), .A2(n5445), .B1(n5745), .B2(n9641), .ZN(n5293)
         );
  NAND2_X1 U6780 ( .A1(n10204), .A2(n5220), .ZN(n5289) );
  OR2_X1 U6781 ( .A1(n7280), .A2(n5345), .ZN(n5288) );
  NAND2_X1 U6782 ( .A1(n5289), .A2(n5288), .ZN(n5290) );
  XNOR2_X1 U6783 ( .A(n5290), .B(n5743), .ZN(n5292) );
  XOR2_X1 U6784 ( .A(n5293), .B(n5292), .Z(n7436) );
  INV_X1 U6785 ( .A(n7436), .ZN(n5291) );
  NAND2_X1 U6786 ( .A1(n7433), .A2(n5291), .ZN(n7434) );
  INV_X1 U6787 ( .A(n5292), .ZN(n5294) );
  NAND2_X1 U6788 ( .A1(n5297), .A2(n5296), .ZN(n5301) );
  INV_X1 U6789 ( .A(n5298), .ZN(n5299) );
  NAND2_X1 U6790 ( .A1(n5299), .A2(SI_7_), .ZN(n5300) );
  INV_X1 U6791 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6530) );
  MUX2_X1 U6792 ( .A(n6530), .B(n6528), .S(n5153), .Z(n5303) );
  INV_X1 U6793 ( .A(SI_8_), .ZN(n5302) );
  INV_X1 U6794 ( .A(n5303), .ZN(n5304) );
  NAND2_X1 U6795 ( .A1(n5304), .A2(SI_8_), .ZN(n5305) );
  NAND2_X1 U6796 ( .A1(n5324), .A2(n5305), .ZN(n5325) );
  NAND2_X1 U6797 ( .A1(n6527), .A2(n5214), .ZN(n5310) );
  NAND2_X1 U6798 ( .A1(n5306), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5307) );
  XNOR2_X1 U6799 ( .A(n5307), .B(n5330), .ZN(n9677) );
  OAI22_X1 U6800 ( .A1(n5587), .A2(n6528), .B1(n9358), .B2(n9677), .ZN(n5308)
         );
  INV_X1 U6801 ( .A(n5308), .ZN(n5309) );
  NAND2_X1 U6802 ( .A1(n5310), .A2(n5309), .ZN(n7502) );
  NAND2_X1 U6803 ( .A1(n7502), .A2(n5220), .ZN(n5320) );
  NAND2_X1 U6804 ( .A1(n9360), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5318) );
  INV_X1 U6805 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5311) );
  OR2_X1 U6806 ( .A1(n5170), .A2(n5311), .ZN(n5317) );
  NAND2_X1 U6807 ( .A1(n5313), .A2(n5312), .ZN(n5314) );
  NAND2_X1 U6808 ( .A1(n5339), .A2(n5314), .ZN(n7292) );
  OR2_X1 U6809 ( .A1(n5129), .A2(n7292), .ZN(n5316) );
  INV_X1 U6810 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6673) );
  OR2_X1 U6811 ( .A1(n9364), .A2(n6673), .ZN(n5315) );
  OR2_X1 U6812 ( .A1(n7452), .A2(n5345), .ZN(n5319) );
  NAND2_X1 U6813 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  INV_X1 U6814 ( .A(n7502), .ZN(n7720) );
  OAI22_X1 U6815 ( .A1(n7720), .A2(n5345), .B1(n7452), .B2(n5817), .ZN(n7714)
         );
  MUX2_X1 U6816 ( .A(n6532), .B(n6542), .S(n9356), .Z(n5327) );
  NAND2_X1 U6817 ( .A1(n5327), .A2(n8774), .ZN(n5352) );
  INV_X1 U6818 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6819 ( .A1(n5328), .A2(SI_9_), .ZN(n5329) );
  NAND2_X1 U6820 ( .A1(n6531), .A2(n5214), .ZN(n5338) );
  AND4_X1 U6821 ( .A1(n5332), .A2(n5331), .A3(n9036), .A4(n5330), .ZN(n5333)
         );
  NAND2_X1 U6822 ( .A1(n5215), .A2(n5333), .ZN(n5353) );
  NAND2_X1 U6823 ( .A1(n5353), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5335) );
  INV_X1 U6824 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n5334) );
  XNOR2_X1 U6825 ( .A(n5335), .B(n5334), .ZN(n10111) );
  OAI22_X1 U6826 ( .A1(n5587), .A2(n6542), .B1(n9358), .B2(n10111), .ZN(n5336)
         );
  INV_X1 U6827 ( .A(n5336), .ZN(n5337) );
  NAND2_X1 U6828 ( .A1(n5338), .A2(n5337), .ZN(n7459) );
  NAND2_X1 U6829 ( .A1(n7459), .A2(n5220), .ZN(n5347) );
  NAND2_X1 U6830 ( .A1(n4614), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5344) );
  INV_X1 U6831 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n8990) );
  OR2_X1 U6832 ( .A1(n5251), .A2(n8990), .ZN(n5343) );
  INV_X1 U6833 ( .A(n5357), .ZN(n5359) );
  NAND2_X1 U6834 ( .A1(n5339), .A2(n7786), .ZN(n5340) );
  NAND2_X1 U6835 ( .A1(n5359), .A2(n5340), .ZN(n7785) );
  OR2_X1 U6836 ( .A1(n5129), .A2(n7785), .ZN(n5342) );
  INV_X1 U6837 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7457) );
  OR2_X1 U6838 ( .A1(n9364), .A2(n7457), .ZN(n5341) );
  OR2_X1 U6839 ( .A1(n7344), .A2(n5345), .ZN(n5346) );
  NAND2_X1 U6840 ( .A1(n5347), .A2(n5346), .ZN(n5348) );
  XNOR2_X1 U6841 ( .A(n5348), .B(n5743), .ZN(n5351) );
  OAI22_X1 U6842 ( .A1(n10213), .A2(n5345), .B1(n7344), .B2(n5817), .ZN(n5350)
         );
  XNOR2_X1 U6843 ( .A(n5351), .B(n5350), .ZN(n7782) );
  INV_X1 U6844 ( .A(n7782), .ZN(n5349) );
  MUX2_X1 U6845 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n9356), .Z(n5370) );
  XNOR2_X1 U6846 ( .A(n5371), .B(n4500), .ZN(n6546) );
  NAND2_X1 U6847 ( .A1(n6546), .A2(n5214), .ZN(n5356) );
  INV_X1 U6848 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U6849 ( .A1(n5353), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5459) );
  OR2_X1 U6850 ( .A1(n5459), .A2(n10074), .ZN(n5404) );
  INV_X1 U6851 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5376) );
  XNOR2_X1 U6852 ( .A(n5404), .B(n5376), .ZN(n6807) );
  OAI22_X1 U6853 ( .A1(n5587), .A2(n6548), .B1(n9358), .B2(n6807), .ZN(n5354)
         );
  INV_X1 U6854 ( .A(n5354), .ZN(n5355) );
  NAND2_X1 U6855 ( .A1(n4614), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5364) );
  INV_X1 U6856 ( .A(n5383), .ZN(n5385) );
  INV_X1 U6857 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U6858 ( .A1(n5359), .A2(n5358), .ZN(n5360) );
  NAND2_X1 U6859 ( .A1(n5385), .A2(n5360), .ZN(n9199) );
  OR2_X1 U6860 ( .A1(n5129), .A2(n9199), .ZN(n5363) );
  INV_X1 U6861 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7352) );
  OR2_X1 U6862 ( .A1(n9364), .A2(n7352), .ZN(n5362) );
  INV_X1 U6863 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8991) );
  OR2_X1 U6864 ( .A1(n5251), .A2(n8991), .ZN(n5361) );
  INV_X1 U6865 ( .A(n7665), .ZN(n9638) );
  AOI22_X1 U6866 ( .A1(n7426), .A2(n5220), .B1(n5445), .B2(n9638), .ZN(n5365)
         );
  XNOR2_X1 U6867 ( .A(n5365), .B(n5743), .ZN(n5366) );
  OR2_X1 U6868 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  NAND2_X1 U6869 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  AOI22_X1 U6870 ( .A1(n7426), .A2(n5445), .B1(n5745), .B2(n9638), .ZN(n9197)
         );
  MUX2_X1 U6871 ( .A(n6562), .B(n6563), .S(n9356), .Z(n5373) );
  INV_X1 U6872 ( .A(SI_11_), .ZN(n5372) );
  NAND2_X1 U6873 ( .A1(n5373), .A2(n5372), .ZN(n5398) );
  INV_X1 U6874 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6875 ( .A1(n5374), .A2(SI_11_), .ZN(n5375) );
  NAND2_X1 U6876 ( .A1(n5398), .A2(n5375), .ZN(n5399) );
  XNOR2_X1 U6877 ( .A(n5400), .B(n5399), .ZN(n6561) );
  NAND2_X1 U6878 ( .A1(n6561), .A2(n5214), .ZN(n5382) );
  NAND2_X1 U6879 ( .A1(n5404), .A2(n5376), .ZN(n5377) );
  NAND2_X1 U6880 ( .A1(n5377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5379) );
  INV_X1 U6881 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U6882 ( .A(n5379), .B(n5378), .ZN(n10118) );
  OAI22_X1 U6883 ( .A1(n5587), .A2(n6563), .B1(n9358), .B2(n10118), .ZN(n5380)
         );
  INV_X1 U6884 ( .A(n5380), .ZN(n5381) );
  NAND2_X1 U6885 ( .A1(n10187), .A2(n5220), .ZN(n5393) );
  NAND2_X1 U6886 ( .A1(n4614), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5391) );
  INV_X1 U6887 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6808) );
  OR2_X1 U6888 ( .A1(n5251), .A2(n6808), .ZN(n5390) );
  INV_X1 U6889 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5384) );
  NAND2_X1 U6890 ( .A1(n5385), .A2(n5384), .ZN(n5386) );
  NAND2_X1 U6891 ( .A1(n5412), .A2(n5386), .ZN(n10183) );
  OR2_X1 U6892 ( .A1(n5129), .A2(n10183), .ZN(n5389) );
  INV_X1 U6893 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6803) );
  OR2_X1 U6894 ( .A1(n9364), .A2(n6803), .ZN(n5388) );
  OR2_X1 U6895 ( .A1(n7506), .A2(n5345), .ZN(n5392) );
  NAND2_X1 U6896 ( .A1(n5393), .A2(n5392), .ZN(n5394) );
  XNOR2_X1 U6897 ( .A(n5394), .B(n5820), .ZN(n5397) );
  NOR2_X1 U6898 ( .A1(n7506), .A2(n5817), .ZN(n5395) );
  AOI21_X1 U6899 ( .B1(n10187), .B2(n5445), .A(n5395), .ZN(n5396) );
  OR2_X1 U6900 ( .A1(n5397), .A2(n5396), .ZN(n9307) );
  NAND2_X1 U6901 ( .A1(n5397), .A2(n5396), .ZN(n9309) );
  MUX2_X1 U6902 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n4525), .Z(n5424) );
  XNOR2_X1 U6903 ( .A(n5424), .B(SI_12_), .ZN(n5426) );
  INV_X1 U6904 ( .A(n5426), .ZN(n5401) );
  XNOR2_X1 U6905 ( .A(n5427), .B(n5401), .ZN(n6592) );
  NAND2_X1 U6906 ( .A1(n6592), .A2(n5214), .ZN(n5409) );
  INV_X1 U6907 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6650) );
  OR2_X1 U6908 ( .A1(n5402), .A2(n10074), .ZN(n5403) );
  NAND2_X1 U6909 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U6910 ( .A1(n5405), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5406) );
  OAI22_X1 U6911 ( .A1(n5587), .A2(n6650), .B1(n9358), .B2(n6809), .ZN(n5407)
         );
  INV_X1 U6912 ( .A(n5407), .ZN(n5408) );
  NAND2_X1 U6913 ( .A1(n4614), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5417) );
  INV_X1 U6914 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5410) );
  OR2_X1 U6915 ( .A1(n5251), .A2(n5410), .ZN(n5416) );
  NAND2_X1 U6916 ( .A1(n5412), .A2(n5411), .ZN(n5413) );
  NAND2_X1 U6917 ( .A1(n5436), .A2(n5413), .ZN(n9227) );
  OR2_X1 U6918 ( .A1(n5129), .A2(n9227), .ZN(n5415) );
  INV_X1 U6919 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7516) );
  OR2_X1 U6920 ( .A1(n9364), .A2(n7516), .ZN(n5414) );
  INV_X1 U6921 ( .A(n7666), .ZN(n9636) );
  AOI22_X1 U6922 ( .A1(n9229), .A2(n5445), .B1(n5745), .B2(n9636), .ZN(n5421)
         );
  NAND2_X1 U6923 ( .A1(n9229), .A2(n5220), .ZN(n5419) );
  OR2_X1 U6924 ( .A1(n7666), .A2(n5345), .ZN(n5418) );
  NAND2_X1 U6925 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  XNOR2_X1 U6926 ( .A(n5420), .B(n5743), .ZN(n5423) );
  XOR2_X1 U6927 ( .A(n5421), .B(n5423), .Z(n9224) );
  INV_X1 U6928 ( .A(n5421), .ZN(n5422) );
  NAND2_X1 U6929 ( .A1(n5424), .A2(SI_12_), .ZN(n5425) );
  OAI21_X1 U6930 ( .B1(n5427), .B2(n5426), .A(n5425), .ZN(n5448) );
  INV_X1 U6931 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n5428) );
  MUX2_X1 U6932 ( .A(n5428), .B(n6778), .S(n9356), .Z(n5449) );
  XNOR2_X1 U6933 ( .A(n5449), .B(SI_13_), .ZN(n5447) );
  INV_X1 U6934 ( .A(n5447), .ZN(n5429) );
  XNOR2_X1 U6935 ( .A(n5448), .B(n5429), .ZN(n6732) );
  NAND2_X1 U6936 ( .A1(n6732), .A2(n5214), .ZN(n5434) );
  NAND2_X1 U6937 ( .A1(n5430), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5431) );
  XNOR2_X1 U6938 ( .A(n5431), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10133) );
  OAI22_X1 U6939 ( .A1(n5587), .A2(n6778), .B1(n9358), .B2(n7411), .ZN(n5432)
         );
  INV_X1 U6940 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U6941 ( .A1(n9294), .A2(n5220), .ZN(n5443) );
  NAND2_X1 U6942 ( .A1(n9360), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5441) );
  INV_X1 U6943 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5435) );
  OR2_X1 U6944 ( .A1(n5170), .A2(n5435), .ZN(n5440) );
  NAND2_X1 U6945 ( .A1(n5436), .A2(n8999), .ZN(n5437) );
  NAND2_X1 U6946 ( .A1(n5466), .A2(n5437), .ZN(n9292) );
  OR2_X1 U6947 ( .A1(n5129), .A2(n9292), .ZN(n5439) );
  INV_X1 U6948 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7640) );
  OR2_X1 U6949 ( .A1(n9364), .A2(n7640), .ZN(n5438) );
  OR2_X1 U6950 ( .A1(n7703), .A2(n5345), .ZN(n5442) );
  NAND2_X1 U6951 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  XNOR2_X1 U6952 ( .A(n5444), .B(n5743), .ZN(n5476) );
  NOR2_X1 U6953 ( .A1(n7703), .A2(n5817), .ZN(n5446) );
  AOI21_X1 U6954 ( .B1(n9294), .B2(n5445), .A(n5446), .ZN(n5477) );
  XNOR2_X1 U6955 ( .A(n5476), .B(n5477), .ZN(n9288) );
  NAND2_X1 U6956 ( .A1(n9287), .A2(n9288), .ZN(n9175) );
  NAND2_X1 U6957 ( .A1(n5448), .A2(n5447), .ZN(n5452) );
  INV_X1 U6958 ( .A(n5449), .ZN(n5450) );
  NAND2_X1 U6959 ( .A1(n5450), .A2(SI_13_), .ZN(n5451) );
  MUX2_X1 U6960 ( .A(n6832), .B(n9016), .S(n9356), .Z(n5454) );
  NAND2_X1 U6961 ( .A1(n5454), .A2(n5453), .ZN(n5482) );
  INV_X1 U6962 ( .A(n5454), .ZN(n5455) );
  NAND2_X1 U6963 ( .A1(n5455), .A2(SI_14_), .ZN(n5456) );
  NAND2_X1 U6964 ( .A1(n5482), .A2(n5456), .ZN(n5483) );
  XNOR2_X1 U6965 ( .A(n5484), .B(n5483), .ZN(n6831) );
  NAND2_X1 U6966 ( .A1(n6831), .A2(n5214), .ZN(n5463) );
  NOR2_X1 U6967 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5457) );
  AND2_X1 U6968 ( .A1(n5402), .A2(n5457), .ZN(n5458) );
  NAND2_X1 U6969 ( .A1(n5459), .A2(n5458), .ZN(n5506) );
  NAND2_X1 U6970 ( .A1(n5506), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U6971 ( .A(n5460), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10145) );
  INV_X1 U6972 ( .A(n10145), .ZN(n7407) );
  OAI22_X1 U6973 ( .A1(n5587), .A2(n9016), .B1(n9358), .B2(n7407), .ZN(n5461)
         );
  INV_X1 U6974 ( .A(n5461), .ZN(n5462) );
  NAND2_X1 U6975 ( .A1(n10015), .A2(n5220), .ZN(n5473) );
  NAND2_X1 U6976 ( .A1(n4614), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5471) );
  INV_X1 U6977 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5464) );
  OR2_X1 U6978 ( .A1(n9364), .A2(n5464), .ZN(n5470) );
  INV_X1 U6979 ( .A(n5496), .ZN(n5514) );
  NAND2_X1 U6980 ( .A1(n5466), .A2(n5465), .ZN(n5467) );
  NAND2_X1 U6981 ( .A1(n5514), .A2(n5467), .ZN(n9182) );
  OR2_X1 U6982 ( .A1(n5129), .A2(n9182), .ZN(n5469) );
  INV_X1 U6983 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7402) );
  OR2_X1 U6984 ( .A1(n5251), .A2(n7402), .ZN(n5468) );
  OR2_X1 U6985 ( .A1(n7795), .A2(n5345), .ZN(n5472) );
  NAND2_X1 U6986 ( .A1(n5473), .A2(n5472), .ZN(n5474) );
  XNOR2_X1 U6987 ( .A(n5474), .B(n5820), .ZN(n9177) );
  NOR2_X1 U6988 ( .A1(n7795), .A2(n5817), .ZN(n5475) );
  AOI21_X1 U6989 ( .B1(n10015), .B2(n5445), .A(n5475), .ZN(n9176) );
  INV_X1 U6990 ( .A(n5476), .ZN(n5478) );
  AND2_X1 U6991 ( .A1(n5478), .A2(n5477), .ZN(n9173) );
  AOI21_X1 U6992 ( .B1(n9177), .B2(n9176), .A(n9173), .ZN(n5481) );
  INV_X1 U6993 ( .A(n9177), .ZN(n5480) );
  INV_X1 U6994 ( .A(n9176), .ZN(n5479) );
  MUX2_X1 U6995 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n9356), .Z(n5485) );
  INV_X1 U6996 ( .A(n5485), .ZN(n5486) );
  MUX2_X1 U6997 ( .A(n5487), .B(n6943), .S(n9356), .Z(n5488) );
  NAND2_X1 U6998 ( .A1(n5488), .A2(n9021), .ZN(n5533) );
  INV_X1 U6999 ( .A(n5488), .ZN(n5489) );
  NAND2_X1 U7000 ( .A1(n5489), .A2(SI_16_), .ZN(n5490) );
  NAND2_X1 U7001 ( .A1(n5533), .A2(n5490), .ZN(n5534) );
  XNOR2_X1 U7002 ( .A(n5535), .B(n5534), .ZN(n6913) );
  NAND2_X1 U7003 ( .A1(n6913), .A2(n5214), .ZN(n5495) );
  NAND2_X1 U7004 ( .A1(n5491), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5492) );
  XNOR2_X1 U7005 ( .A(n5492), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7576) );
  INV_X1 U7006 ( .A(n7576), .ZN(n7574) );
  OAI22_X1 U7007 ( .A1(n5587), .A2(n6943), .B1(n9358), .B2(n7574), .ZN(n5493)
         );
  INV_X1 U7008 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7009 ( .A1(n5496), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U7010 ( .A1(n5516), .A2(n5497), .ZN(n5498) );
  NAND2_X1 U7011 ( .A1(n5545), .A2(n5498), .ZN(n9251) );
  INV_X1 U7012 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n7575) );
  OAI22_X1 U7013 ( .A1(n9251), .A2(n5129), .B1(n5251), .B2(n7575), .ZN(n5501)
         );
  INV_X1 U7014 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U7015 ( .A1(n4614), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5499) );
  OAI21_X1 U7016 ( .B1(n9364), .B2(n7861), .A(n5499), .ZN(n5500) );
  AOI22_X1 U7017 ( .A1(n10011), .A2(n5220), .B1(n5445), .B2(n9632), .ZN(n5502)
         );
  XOR2_X1 U7018 ( .A(n5743), .B(n5502), .Z(n9245) );
  NAND2_X1 U7019 ( .A1(n10011), .A2(n5445), .ZN(n5504) );
  NAND2_X1 U7020 ( .A1(n9632), .A2(n5745), .ZN(n5503) );
  NAND2_X1 U7021 ( .A1(n5504), .A2(n5503), .ZN(n5526) );
  XNOR2_X1 U7022 ( .A(n5505), .B(n4501), .ZN(n6886) );
  NAND2_X1 U7023 ( .A1(n6886), .A2(n5214), .ZN(n5511) );
  INV_X1 U7024 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6908) );
  OAI21_X1 U7025 ( .B1(n5506), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5507) );
  MUX2_X1 U7026 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5507), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n5508) );
  NAND2_X1 U7027 ( .A1(n5508), .A2(n5491), .ZN(n7413) );
  OAI22_X1 U7028 ( .A1(n5587), .A2(n6908), .B1(n9358), .B2(n7413), .ZN(n5509)
         );
  INV_X1 U7029 ( .A(n5509), .ZN(n5510) );
  NAND2_X1 U7030 ( .A1(n9352), .A2(n5220), .ZN(n5522) );
  NAND2_X1 U7031 ( .A1(n9360), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5520) );
  INV_X1 U7032 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5512) );
  OR2_X1 U7033 ( .A1(n5170), .A2(n5512), .ZN(n5519) );
  INV_X1 U7034 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U7035 ( .A1(n5514), .A2(n5513), .ZN(n5515) );
  NAND2_X1 U7036 ( .A1(n5516), .A2(n5515), .ZN(n9348) );
  OR2_X1 U7037 ( .A1(n5129), .A2(n9348), .ZN(n5518) );
  INV_X1 U7038 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8994) );
  OR2_X1 U7039 ( .A1(n9364), .A2(n8994), .ZN(n5517) );
  OR2_X1 U7040 ( .A1(n7853), .A2(n5345), .ZN(n5521) );
  NAND2_X1 U7041 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  XNOR2_X1 U7042 ( .A(n5523), .B(n5743), .ZN(n5529) );
  NAND2_X1 U7043 ( .A1(n9352), .A2(n5445), .ZN(n5525) );
  OR2_X1 U7044 ( .A1(n7853), .A2(n5817), .ZN(n5524) );
  NAND2_X1 U7045 ( .A1(n5525), .A2(n5524), .ZN(n9344) );
  AOI22_X1 U7046 ( .A1(n9245), .A2(n5526), .B1(n5529), .B2(n9344), .ZN(n5532)
         );
  INV_X1 U7047 ( .A(n5529), .ZN(n9243) );
  INV_X1 U7048 ( .A(n9344), .ZN(n5527) );
  INV_X1 U7049 ( .A(n5526), .ZN(n9244) );
  AOI21_X1 U7050 ( .B1(n9243), .B2(n5527), .A(n9244), .ZN(n5530) );
  NAND2_X1 U7051 ( .A1(n9244), .A2(n5527), .ZN(n5528) );
  OAI22_X1 U7052 ( .A1(n9245), .A2(n5530), .B1(n5529), .B2(n5528), .ZN(n5531)
         );
  MUX2_X1 U7053 ( .A(n9018), .B(n7094), .S(n4525), .Z(n5537) );
  NAND2_X1 U7054 ( .A1(n5537), .A2(n5536), .ZN(n5559) );
  INV_X1 U7055 ( .A(n5537), .ZN(n5538) );
  NAND2_X1 U7056 ( .A1(n5538), .A2(SI_17_), .ZN(n5539) );
  XNOR2_X1 U7057 ( .A(n5558), .B(n5557), .ZN(n7077) );
  NAND2_X1 U7058 ( .A1(n7077), .A2(n5214), .ZN(n5544) );
  XNOR2_X1 U7059 ( .A(n5541), .B(n5540), .ZN(n9689) );
  OAI22_X1 U7060 ( .A1(n5587), .A2(n7094), .B1(n9358), .B2(n9689), .ZN(n5542)
         );
  INV_X1 U7061 ( .A(n5542), .ZN(n5543) );
  NAND2_X1 U7062 ( .A1(n10003), .A2(n5220), .ZN(n5552) );
  INV_X1 U7063 ( .A(n5566), .ZN(n5567) );
  NAND2_X1 U7064 ( .A1(n5545), .A2(n7582), .ZN(n5546) );
  NAND2_X1 U7065 ( .A1(n5567), .A2(n5546), .ZN(n9924) );
  OR2_X1 U7066 ( .A1(n9924), .A2(n5129), .ZN(n5550) );
  AOI22_X1 U7067 ( .A1(n9360), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n4614), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5549) );
  INV_X1 U7068 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5547) );
  OR2_X1 U7069 ( .A1(n9364), .A2(n5547), .ZN(n5548) );
  NAND2_X1 U7070 ( .A1(n9631), .A2(n5445), .ZN(n5551) );
  NAND2_X1 U7071 ( .A1(n5552), .A2(n5551), .ZN(n5553) );
  XNOR2_X1 U7072 ( .A(n5553), .B(n5820), .ZN(n5556) );
  NOR2_X1 U7073 ( .A1(n7854), .A2(n5817), .ZN(n5554) );
  AOI21_X1 U7074 ( .B1(n10003), .B2(n5445), .A(n5554), .ZN(n5555) );
  NOR2_X1 U7075 ( .A1(n5556), .A2(n5555), .ZN(n9256) );
  NAND2_X1 U7076 ( .A1(n5558), .A2(n5557), .ZN(n5560) );
  NAND2_X1 U7077 ( .A1(n5560), .A2(n5559), .ZN(n5582) );
  MUX2_X1 U7078 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4525), .Z(n5580) );
  XNOR2_X1 U7079 ( .A(n5582), .B(n4502), .ZN(n7115) );
  NAND2_X1 U7080 ( .A1(n7115), .A2(n5214), .ZN(n5565) );
  INV_X1 U7081 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9017) );
  XNOR2_X1 U7082 ( .A(n5562), .B(n5561), .ZN(n10170) );
  OAI22_X1 U7083 ( .A1(n5587), .A2(n9017), .B1(n9358), .B2(n10170), .ZN(n5563)
         );
  INV_X1 U7084 ( .A(n5563), .ZN(n5564) );
  NAND2_X1 U7085 ( .A1(n9911), .A2(n5220), .ZN(n5573) );
  INV_X1 U7086 ( .A(n5591), .ZN(n5593) );
  INV_X1 U7087 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U7088 ( .A1(n5567), .A2(n9322), .ZN(n5568) );
  AND2_X1 U7089 ( .A1(n5593), .A2(n5568), .ZN(n9912) );
  NAND2_X1 U7090 ( .A1(n9912), .A2(n5171), .ZN(n5571) );
  AOI22_X1 U7091 ( .A1(n9360), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n4614), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5570) );
  INV_X1 U7092 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n10166) );
  OR2_X1 U7093 ( .A1(n9364), .A2(n10166), .ZN(n5569) );
  INV_X1 U7094 ( .A(n9259), .ZN(n9630) );
  NAND2_X1 U7095 ( .A1(n9630), .A2(n5445), .ZN(n5572) );
  NAND2_X1 U7096 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  XNOR2_X1 U7097 ( .A(n5574), .B(n5820), .ZN(n5576) );
  NOR2_X1 U7098 ( .A1(n9259), .A2(n5817), .ZN(n5575) );
  AOI21_X1 U7099 ( .B1(n9911), .B2(n5445), .A(n5575), .ZN(n5577) );
  AND2_X1 U7100 ( .A1(n5576), .A2(n5577), .ZN(n9316) );
  INV_X1 U7101 ( .A(n5576), .ZN(n5579) );
  INV_X1 U7102 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U7103 ( .A1(n5579), .A2(n5578), .ZN(n9317) );
  NAND2_X1 U7104 ( .A1(n5580), .A2(SI_18_), .ZN(n5581) );
  MUX2_X1 U7105 ( .A(n7302), .B(n8975), .S(n4525), .Z(n5584) );
  NAND2_X1 U7106 ( .A1(n5584), .A2(n5583), .ZN(n5607) );
  INV_X1 U7107 ( .A(n5584), .ZN(n5585) );
  NAND2_X1 U7108 ( .A1(n5585), .A2(SI_19_), .ZN(n5586) );
  NAND2_X1 U7109 ( .A1(n5607), .A2(n5586), .ZN(n5608) );
  XNOR2_X1 U7110 ( .A(n5609), .B(n5608), .ZN(n7299) );
  NAND2_X1 U7111 ( .A1(n7299), .A2(n5214), .ZN(n5590) );
  OAI22_X1 U7112 ( .A1(n5587), .A2(n8975), .B1(n7300), .B2(n9358), .ZN(n5588)
         );
  INV_X1 U7113 ( .A(n5588), .ZN(n5589) );
  INV_X1 U7114 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7115 ( .A1(n5593), .A2(n5592), .ZN(n5594) );
  NAND2_X1 U7116 ( .A1(n5614), .A2(n5594), .ZN(n9889) );
  OR2_X1 U7117 ( .A1(n9889), .A2(n5129), .ZN(n5599) );
  INV_X1 U7118 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9693) );
  NAND2_X1 U7119 ( .A1(n4614), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U7120 ( .A1(n5387), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5595) );
  OAI211_X1 U7121 ( .C1(n5251), .C2(n9693), .A(n5596), .B(n5595), .ZN(n5597)
         );
  INV_X1 U7122 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7123 ( .A1(n5599), .A2(n5598), .ZN(n9629) );
  OAI22_X1 U7124 ( .A1(n9892), .A2(n5600), .B1(n9280), .B2(n5345), .ZN(n5601)
         );
  XNOR2_X1 U7125 ( .A(n5601), .B(n5820), .ZN(n9208) );
  OR2_X1 U7126 ( .A1(n9892), .A2(n5345), .ZN(n5603) );
  NAND2_X1 U7127 ( .A1(n9629), .A2(n5745), .ZN(n5602) );
  AND2_X1 U7128 ( .A1(n5603), .A2(n5602), .ZN(n5604) );
  NAND2_X1 U7129 ( .A1(n9208), .A2(n5604), .ZN(n5606) );
  INV_X1 U7130 ( .A(n9208), .ZN(n5605) );
  INV_X1 U7131 ( .A(n5604), .ZN(n9207) );
  MUX2_X1 U7132 ( .A(n7379), .B(n8976), .S(n4525), .Z(n5629) );
  XNOR2_X1 U7133 ( .A(n5629), .B(SI_20_), .ZN(n5626) );
  XNOR2_X1 U7134 ( .A(n5627), .B(n5626), .ZN(n7378) );
  NAND2_X1 U7135 ( .A1(n7378), .A2(n5214), .ZN(n5612) );
  NAND2_X1 U7136 ( .A1(n5610), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5611) );
  INV_X1 U7137 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5613) );
  NAND2_X1 U7138 ( .A1(n5614), .A2(n5613), .ZN(n5615) );
  AND2_X1 U7139 ( .A1(n5635), .A2(n5615), .ZN(n9879) );
  NAND2_X1 U7140 ( .A1(n9879), .A2(n5171), .ZN(n5620) );
  INV_X1 U7141 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n8951) );
  NAND2_X1 U7142 ( .A1(n9360), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U7143 ( .A1(n4614), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5616) );
  OAI211_X1 U7144 ( .C1(n8951), .C2(n9364), .A(n5617), .B(n5616), .ZN(n5618)
         );
  INV_X1 U7145 ( .A(n5618), .ZN(n5619) );
  AOI22_X1 U7146 ( .A1(n9878), .A2(n5220), .B1(n5445), .B2(n9628), .ZN(n5621)
         );
  XOR2_X1 U7147 ( .A(n5743), .B(n5621), .Z(n5623) );
  OAI22_X1 U7148 ( .A1(n10062), .A2(n5345), .B1(n9371), .B2(n5817), .ZN(n5622)
         );
  NOR2_X1 U7149 ( .A1(n5623), .A2(n5622), .ZN(n5624) );
  AOI21_X1 U7150 ( .B1(n5623), .B2(n5622), .A(n5624), .ZN(n9279) );
  INV_X1 U7151 ( .A(n5624), .ZN(n5625) );
  INV_X1 U7152 ( .A(SI_20_), .ZN(n5628) );
  MUX2_X1 U7153 ( .A(n7604), .B(n8952), .S(n4525), .Z(n5631) );
  NAND2_X1 U7154 ( .A1(n5630), .A2(n5631), .ZN(n5651) );
  NAND2_X1 U7155 ( .A1(n5650), .A2(n5651), .ZN(n5632) );
  NAND2_X1 U7156 ( .A1(n7602), .A2(n5214), .ZN(n5634) );
  NAND2_X1 U7157 ( .A1(n5610), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5633) );
  NAND2_X1 U7158 ( .A1(n9861), .A2(n5220), .ZN(n5643) );
  INV_X1 U7159 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7160 ( .A1(n5635), .A2(n9035), .ZN(n5636) );
  NAND2_X1 U7161 ( .A1(n5660), .A2(n5636), .ZN(n9862) );
  OR2_X1 U7162 ( .A1(n9862), .A2(n5129), .ZN(n5641) );
  INV_X1 U7163 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9984) );
  NAND2_X1 U7164 ( .A1(n5387), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U7165 ( .A1(n4614), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5637) );
  OAI211_X1 U7166 ( .C1(n5251), .C2(n9984), .A(n5638), .B(n5637), .ZN(n5639)
         );
  INV_X1 U7167 ( .A(n5639), .ZN(n5640) );
  NAND2_X1 U7168 ( .A1(n9627), .A2(n5445), .ZN(n5642) );
  NAND2_X1 U7169 ( .A1(n5643), .A2(n5642), .ZN(n5644) );
  XNOR2_X1 U7170 ( .A(n5644), .B(n5743), .ZN(n5647) );
  AOI22_X1 U7171 ( .A1(n9861), .A2(n5445), .B1(n5745), .B2(n9627), .ZN(n5645)
         );
  XNOR2_X1 U7172 ( .A(n5647), .B(n5645), .ZN(n9216) );
  NAND2_X1 U7173 ( .A1(n9215), .A2(n9216), .ZN(n9214) );
  INV_X1 U7174 ( .A(n5645), .ZN(n5646) );
  NAND2_X1 U7175 ( .A1(n9214), .A2(n5648), .ZN(n5670) );
  INV_X1 U7176 ( .A(n5670), .ZN(n5668) );
  INV_X1 U7177 ( .A(SI_21_), .ZN(n5649) );
  NAND2_X1 U7178 ( .A1(n5650), .A2(n5649), .ZN(n5652) );
  NAND2_X1 U7179 ( .A1(n5652), .A2(n5651), .ZN(n5672) );
  MUX2_X1 U7180 ( .A(n7647), .B(n8977), .S(n4525), .Z(n5654) );
  INV_X1 U7181 ( .A(SI_22_), .ZN(n5653) );
  NAND2_X1 U7182 ( .A1(n5654), .A2(n5653), .ZN(n5673) );
  INV_X1 U7183 ( .A(n5654), .ZN(n5655) );
  NAND2_X1 U7184 ( .A1(n5655), .A2(SI_22_), .ZN(n5656) );
  NAND2_X1 U7185 ( .A1(n7646), .A2(n5214), .ZN(n5658) );
  NAND2_X1 U7186 ( .A1(n5610), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5657) );
  NAND2_X1 U7187 ( .A1(n5659), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5681) );
  INV_X1 U7188 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U7189 ( .A1(n5660), .A2(n8923), .ZN(n5661) );
  NAND2_X1 U7190 ( .A1(n5681), .A2(n5661), .ZN(n9843) );
  OR2_X1 U7191 ( .A1(n9843), .A2(n5129), .ZN(n5666) );
  INV_X1 U7192 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U7193 ( .A1(n5387), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U7194 ( .A1(n4614), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5662) );
  OAI211_X1 U7195 ( .C1(n5251), .C2(n9979), .A(n5663), .B(n5662), .ZN(n5664)
         );
  INV_X1 U7196 ( .A(n5664), .ZN(n5665) );
  AOI22_X1 U7197 ( .A1(n9842), .A2(n5220), .B1(n5445), .B2(n9626), .ZN(n5667)
         );
  XNOR2_X1 U7198 ( .A(n5667), .B(n5743), .ZN(n5669) );
  AOI22_X1 U7199 ( .A1(n9842), .A2(n5445), .B1(n5745), .B2(n9626), .ZN(n9297)
         );
  NAND2_X1 U7200 ( .A1(n5672), .A2(n5671), .ZN(n5674) );
  NAND2_X1 U7201 ( .A1(n5674), .A2(n5673), .ZN(n5699) );
  INV_X1 U7202 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5675) );
  MUX2_X1 U7203 ( .A(n5675), .B(n8783), .S(n4525), .Z(n5677) );
  INV_X1 U7204 ( .A(SI_23_), .ZN(n5676) );
  NAND2_X1 U7205 ( .A1(n5677), .A2(n5676), .ZN(n5722) );
  INV_X1 U7206 ( .A(n5677), .ZN(n5678) );
  NAND2_X1 U7207 ( .A1(n5678), .A2(SI_23_), .ZN(n5679) );
  XNOR2_X1 U7208 ( .A(n5699), .B(n5698), .ZN(n7657) );
  NAND2_X1 U7209 ( .A1(n5610), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5680) );
  NAND2_X1 U7210 ( .A1(n9827), .A2(n5220), .ZN(n5689) );
  NAND2_X1 U7211 ( .A1(n5681), .A2(n9191), .ZN(n5682) );
  NAND2_X1 U7212 ( .A1(n5736), .A2(n5682), .ZN(n9828) );
  OR2_X1 U7213 ( .A1(n9828), .A2(n5129), .ZN(n5687) );
  INV_X1 U7214 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9974) );
  NAND2_X1 U7215 ( .A1(n5387), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U7216 ( .A1(n4614), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5683) );
  OAI211_X1 U7217 ( .C1(n5251), .C2(n9974), .A(n5684), .B(n5683), .ZN(n5685)
         );
  INV_X1 U7218 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U7219 ( .A1(n9625), .A2(n5445), .ZN(n5688) );
  NAND2_X1 U7220 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  XNOR2_X1 U7221 ( .A(n5690), .B(n5820), .ZN(n5692) );
  NOR2_X1 U7222 ( .A1(n9512), .A2(n5817), .ZN(n5691) );
  AOI21_X1 U7223 ( .B1(n9827), .B2(n5445), .A(n5691), .ZN(n5693) );
  NAND2_X1 U7224 ( .A1(n5692), .A2(n5693), .ZN(n5697) );
  INV_X1 U7225 ( .A(n5692), .ZN(n5695) );
  INV_X1 U7226 ( .A(n5693), .ZN(n5694) );
  NAND2_X1 U7227 ( .A1(n5695), .A2(n5694), .ZN(n5696) );
  NAND2_X1 U7228 ( .A1(n5697), .A2(n5696), .ZN(n9188) );
  INV_X1 U7229 ( .A(n5697), .ZN(n9266) );
  NAND2_X1 U7230 ( .A1(n5699), .A2(n5698), .ZN(n5726) );
  NAND2_X1 U7231 ( .A1(n5726), .A2(n5722), .ZN(n5705) );
  INV_X1 U7232 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n5700) );
  MUX2_X1 U7233 ( .A(n7710), .B(n5700), .S(n4525), .Z(n5702) );
  INV_X1 U7234 ( .A(SI_24_), .ZN(n5701) );
  NAND2_X1 U7235 ( .A1(n5702), .A2(n5701), .ZN(n5721) );
  INV_X1 U7236 ( .A(n5702), .ZN(n5703) );
  NAND2_X1 U7237 ( .A1(n5703), .A2(SI_24_), .ZN(n5723) );
  AND2_X1 U7238 ( .A1(n5721), .A2(n5723), .ZN(n5704) );
  NAND2_X1 U7239 ( .A1(n7679), .A2(n5214), .ZN(n5707) );
  NAND2_X1 U7240 ( .A1(n5610), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5706) );
  NAND2_X1 U7241 ( .A1(n9810), .A2(n5220), .ZN(n5714) );
  XNOR2_X1 U7242 ( .A(n5736), .B(P1_REG3_REG_24__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U7243 ( .A1(n9811), .A2(n5171), .ZN(n5712) );
  INV_X1 U7244 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U7245 ( .A1(n5387), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5709) );
  NAND2_X1 U7246 ( .A1(n4614), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5708) );
  OAI211_X1 U7247 ( .C1(n5251), .C2(n9969), .A(n5709), .B(n5708), .ZN(n5710)
         );
  INV_X1 U7248 ( .A(n5710), .ZN(n5711) );
  OR2_X1 U7249 ( .A1(n9235), .A2(n5345), .ZN(n5713) );
  NAND2_X1 U7250 ( .A1(n5714), .A2(n5713), .ZN(n5715) );
  XNOR2_X1 U7251 ( .A(n5715), .B(n5820), .ZN(n5718) );
  NOR2_X1 U7252 ( .A1(n9235), .A2(n5817), .ZN(n5716) );
  AOI21_X1 U7253 ( .B1(n9810), .B2(n5445), .A(n5716), .ZN(n5717) );
  NAND2_X1 U7254 ( .A1(n5718), .A2(n5717), .ZN(n5720) );
  OR2_X1 U7255 ( .A1(n5718), .A2(n5717), .ZN(n5719) );
  AND2_X1 U7256 ( .A1(n5720), .A2(n5719), .ZN(n9265) );
  NAND2_X1 U7257 ( .A1(n9264), .A2(n5720), .ZN(n9232) );
  AND2_X1 U7258 ( .A1(n5722), .A2(n5721), .ZN(n5725) );
  AOI21_X2 U7259 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5747) );
  INV_X1 U7260 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5728) );
  INV_X1 U7261 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n5727) );
  MUX2_X1 U7262 ( .A(n5728), .B(n5727), .S(n4525), .Z(n5730) );
  INV_X1 U7263 ( .A(SI_25_), .ZN(n5729) );
  NAND2_X1 U7264 ( .A1(n5730), .A2(n5729), .ZN(n5748) );
  INV_X1 U7265 ( .A(n5730), .ZN(n5731) );
  NAND2_X1 U7266 ( .A1(n5731), .A2(SI_25_), .ZN(n5732) );
  XNOR2_X1 U7267 ( .A(n5747), .B(n5746), .ZN(n7724) );
  NAND2_X1 U7268 ( .A1(n7724), .A2(n5214), .ZN(n5734) );
  NAND2_X1 U7269 ( .A1(n5610), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5733) );
  NAND2_X1 U7270 ( .A1(n9792), .A2(n5169), .ZN(n5742) );
  INV_X1 U7271 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9272) );
  INV_X1 U7272 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9237) );
  OAI21_X1 U7273 ( .B1(n5736), .B2(n9272), .A(n9237), .ZN(n5737) );
  NAND2_X1 U7274 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n5735) );
  INV_X1 U7275 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10041) );
  NAND2_X1 U7276 ( .A1(n9360), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5739) );
  NAND2_X1 U7277 ( .A1(n5387), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5738) );
  OAI211_X1 U7278 ( .C1(n5170), .C2(n10041), .A(n5739), .B(n5738), .ZN(n5740)
         );
  OR2_X1 U7279 ( .A1(n9269), .A2(n5345), .ZN(n5741) );
  NAND2_X1 U7280 ( .A1(n5742), .A2(n5741), .ZN(n5744) );
  XNOR2_X1 U7281 ( .A(n5744), .B(n5743), .ZN(n5769) );
  INV_X1 U7282 ( .A(n9269), .ZN(n9623) );
  AOI22_X1 U7283 ( .A1(n9792), .A2(n5445), .B1(n5745), .B2(n9623), .ZN(n5767)
         );
  XNOR2_X1 U7284 ( .A(n5769), .B(n5767), .ZN(n9233) );
  NAND2_X1 U7285 ( .A1(n5747), .A2(n5746), .ZN(n5749) );
  NAND2_X1 U7286 ( .A1(n5749), .A2(n5748), .ZN(n5772) );
  INV_X1 U7287 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7870) );
  INV_X1 U7288 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n5750) );
  MUX2_X1 U7289 ( .A(n7870), .B(n5750), .S(n4525), .Z(n5751) );
  NAND2_X1 U7290 ( .A1(n5751), .A2(n8930), .ZN(n5773) );
  INV_X1 U7291 ( .A(n5751), .ZN(n5752) );
  NAND2_X1 U7292 ( .A1(n5752), .A2(SI_26_), .ZN(n5753) );
  XNOR2_X1 U7293 ( .A(n5772), .B(n5771), .ZN(n7867) );
  NAND2_X1 U7294 ( .A1(n7867), .A2(n5214), .ZN(n5755) );
  NAND2_X1 U7295 ( .A1(n5610), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7296 ( .A1(n9781), .A2(n5220), .ZN(n5764) );
  INV_X1 U7297 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5889) );
  INV_X1 U7298 ( .A(n5783), .ZN(n5785) );
  NAND2_X1 U7299 ( .A1(n5756), .A2(n5889), .ZN(n5757) );
  NAND2_X1 U7300 ( .A1(n5785), .A2(n5757), .ZN(n9775) );
  OR2_X1 U7301 ( .A1(n9775), .A2(n5129), .ZN(n5762) );
  INV_X1 U7302 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U7303 ( .A1(n5387), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5759) );
  NAND2_X1 U7304 ( .A1(n4614), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5758) );
  OAI211_X1 U7305 ( .C1(n5251), .C2(n9959), .A(n5759), .B(n5758), .ZN(n5760)
         );
  INV_X1 U7306 ( .A(n5760), .ZN(n5761) );
  NAND2_X1 U7307 ( .A1(n9622), .A2(n5445), .ZN(n5763) );
  NAND2_X1 U7308 ( .A1(n5764), .A2(n5763), .ZN(n5765) );
  XNOR2_X1 U7309 ( .A(n5765), .B(n5820), .ZN(n5798) );
  NOR2_X1 U7310 ( .A1(n9236), .A2(n5817), .ZN(n5766) );
  AOI21_X1 U7311 ( .B1(n9781), .B2(n5445), .A(n5766), .ZN(n5799) );
  XNOR2_X1 U7312 ( .A(n5798), .B(n5799), .ZN(n5884) );
  INV_X1 U7313 ( .A(n5767), .ZN(n5768) );
  NOR2_X1 U7314 ( .A1(n5769), .A2(n5768), .ZN(n5883) );
  NOR2_X1 U7315 ( .A1(n5884), .A2(n5883), .ZN(n5770) );
  NAND2_X1 U7316 ( .A1(n5772), .A2(n5771), .ZN(n5774) );
  NAND2_X1 U7317 ( .A1(n5774), .A2(n5773), .ZN(n5805) );
  INV_X1 U7318 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5776) );
  INV_X1 U7319 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5775) );
  MUX2_X1 U7320 ( .A(n5776), .B(n5775), .S(n4525), .Z(n5778) );
  INV_X1 U7321 ( .A(SI_27_), .ZN(n5777) );
  NAND2_X1 U7322 ( .A1(n5778), .A2(n5777), .ZN(n5806) );
  INV_X1 U7323 ( .A(n5778), .ZN(n5779) );
  NAND2_X1 U7324 ( .A1(n5779), .A2(SI_27_), .ZN(n5780) );
  XNOR2_X1 U7325 ( .A(n5805), .B(n5804), .ZN(n7885) );
  NAND2_X1 U7326 ( .A1(n7885), .A2(n5214), .ZN(n5782) );
  NAND2_X1 U7327 ( .A1(n5610), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5781) );
  NAND2_X1 U7328 ( .A1(n9759), .A2(n5169), .ZN(n5793) );
  NAND2_X1 U7329 ( .A1(n5783), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n9728) );
  INV_X1 U7330 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5784) );
  NAND2_X1 U7331 ( .A1(n5785), .A2(n5784), .ZN(n5786) );
  NAND2_X1 U7332 ( .A1(n9728), .A2(n5786), .ZN(n6470) );
  OR2_X1 U7333 ( .A1(n6470), .A2(n5129), .ZN(n5791) );
  INV_X1 U7334 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9953) );
  NAND2_X1 U7335 ( .A1(n5387), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5788) );
  NAND2_X1 U7336 ( .A1(n4614), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5787) );
  OAI211_X1 U7337 ( .C1(n5251), .C2(n9953), .A(n5788), .B(n5787), .ZN(n5789)
         );
  INV_X1 U7338 ( .A(n5789), .ZN(n5790) );
  INV_X1 U7339 ( .A(n6413), .ZN(n9621) );
  NAND2_X1 U7340 ( .A1(n9621), .A2(n5445), .ZN(n5792) );
  NAND2_X1 U7341 ( .A1(n5793), .A2(n5792), .ZN(n5794) );
  XNOR2_X1 U7342 ( .A(n5794), .B(n5820), .ZN(n5797) );
  NOR2_X1 U7343 ( .A1(n6413), .A2(n5817), .ZN(n5795) );
  AOI21_X1 U7344 ( .B1(n9759), .B2(n5445), .A(n5795), .ZN(n5796) );
  NAND2_X1 U7345 ( .A1(n5797), .A2(n5796), .ZN(n5875) );
  OAI21_X1 U7346 ( .B1(n5797), .B2(n5796), .A(n5875), .ZN(n6466) );
  INV_X1 U7347 ( .A(n6466), .ZN(n5803) );
  INV_X1 U7348 ( .A(n5798), .ZN(n5801) );
  INV_X1 U7349 ( .A(n5799), .ZN(n5800) );
  INV_X1 U7350 ( .A(n6467), .ZN(n5802) );
  NAND2_X1 U7351 ( .A1(n5805), .A2(n5804), .ZN(n5807) );
  NAND2_X1 U7352 ( .A1(n5807), .A2(n5806), .ZN(n6264) );
  INV_X1 U7353 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8782) );
  INV_X1 U7354 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n5808) );
  MUX2_X1 U7355 ( .A(n8782), .B(n5808), .S(n4525), .Z(n5809) );
  INV_X1 U7356 ( .A(SI_28_), .ZN(n8992) );
  NAND2_X1 U7357 ( .A1(n5809), .A2(n8992), .ZN(n6265) );
  INV_X1 U7358 ( .A(n5809), .ZN(n5810) );
  NAND2_X1 U7359 ( .A1(n5810), .A2(SI_28_), .ZN(n5811) );
  NAND2_X1 U7360 ( .A1(n7908), .A2(n5214), .ZN(n5813) );
  NAND2_X1 U7361 ( .A1(n5610), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5812) );
  NAND2_X1 U7362 ( .A1(n9742), .A2(n5445), .ZN(n5819) );
  XNOR2_X1 U7363 ( .A(n9728), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9744) );
  INV_X1 U7364 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U7365 ( .A1(n5387), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5815) );
  INV_X1 U7366 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n10030) );
  OR2_X1 U7367 ( .A1(n5170), .A2(n10030), .ZN(n5814) );
  OAI211_X1 U7368 ( .C1(n5251), .C2(n9948), .A(n5815), .B(n5814), .ZN(n5816)
         );
  AOI21_X1 U7369 ( .B1(n9744), .B2(n5171), .A(n5816), .ZN(n6471) );
  OR2_X1 U7370 ( .A1(n6471), .A2(n5817), .ZN(n5818) );
  NAND2_X1 U7371 ( .A1(n5819), .A2(n5818), .ZN(n5821) );
  XNOR2_X1 U7372 ( .A(n5821), .B(n5820), .ZN(n5823) );
  INV_X1 U7373 ( .A(n6471), .ZN(n9620) );
  AOI22_X1 U7374 ( .A1(n9742), .A2(n5169), .B1(n5445), .B2(n9620), .ZN(n5822)
         );
  XNOR2_X1 U7375 ( .A(n5823), .B(n5822), .ZN(n5876) );
  INV_X1 U7376 ( .A(n5876), .ZN(n5853) );
  NAND2_X1 U7377 ( .A1(n5827), .A2(P1_B_REG_SCAN_IN), .ZN(n5825) );
  MUX2_X1 U7378 ( .A(P1_B_REG_SCAN_IN), .B(n5825), .S(n5842), .Z(n5826) );
  INV_X1 U7379 ( .A(n7868), .ZN(n5841) );
  NAND2_X1 U7380 ( .A1(n5841), .A2(n5827), .ZN(n10072) );
  NOR2_X1 U7381 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .ZN(
        n8984) );
  NOR4_X1 U7382 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_27__SCAN_IN), .ZN(n5830) );
  NOR4_X1 U7383 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5829) );
  NOR4_X1 U7384 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n5828) );
  AND4_X1 U7385 ( .A1(n8984), .A2(n5830), .A3(n5829), .A4(n5828), .ZN(n5836)
         );
  NOR4_X1 U7386 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n5834) );
  NOR4_X1 U7387 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5833) );
  NOR4_X1 U7388 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n5832) );
  NOR4_X1 U7389 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n5831) );
  AND4_X1 U7390 ( .A1(n5834), .A2(n5833), .A3(n5832), .A4(n5831), .ZN(n5835)
         );
  NAND2_X1 U7391 ( .A1(n5836), .A2(n5835), .ZN(n6459) );
  INV_X1 U7392 ( .A(n6459), .ZN(n5837) );
  NOR2_X1 U7393 ( .A1(n6457), .A2(n5837), .ZN(n5838) );
  NOR2_X1 U7394 ( .A1(n7078), .A2(n5838), .ZN(n5844) );
  INV_X1 U7395 ( .A(n6457), .ZN(n5840) );
  INV_X1 U7396 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U7397 ( .A1(n5840), .A2(n5839), .ZN(n5843) );
  NAND2_X1 U7398 ( .A1(n5842), .A2(n5841), .ZN(n10073) );
  NAND2_X1 U7399 ( .A1(n5846), .A2(n5845), .ZN(n5847) );
  NAND2_X1 U7400 ( .A1(n5847), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5849) );
  AND2_X1 U7401 ( .A1(n5851), .A2(n9601), .ZN(n9595) );
  NOR2_X1 U7402 ( .A1(n10205), .A2(n9595), .ZN(n5852) );
  NAND2_X1 U7403 ( .A1(n5853), .A2(n9329), .ZN(n5881) );
  AND2_X1 U7404 ( .A1(n5876), .A2(n5036), .ZN(n5854) );
  INV_X1 U7405 ( .A(n9605), .ZN(n6444) );
  NAND2_X1 U7406 ( .A1(n6456), .A2(n6444), .ZN(n7088) );
  INV_X1 U7407 ( .A(n7088), .ZN(n5855) );
  AOI21_X2 U7408 ( .B1(n5864), .B2(n5855), .A(n10184), .ZN(n9283) );
  INV_X1 U7409 ( .A(n5856), .ZN(n7909) );
  NAND2_X1 U7410 ( .A1(n5171), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5857) );
  OR2_X1 U7411 ( .A1(n9728), .A2(n5857), .ZN(n5862) );
  INV_X1 U7412 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U7413 ( .A1(n4614), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U7414 ( .A1(n5387), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5858) );
  OAI211_X1 U7415 ( .C1(n5251), .C2(n6492), .A(n5859), .B(n5858), .ZN(n5860)
         );
  INV_X1 U7416 ( .A(n5860), .ZN(n5861) );
  OAI22_X1 U7417 ( .A1(n6413), .A2(n9300), .B1(n6885), .B2(n9301), .ZN(n9736)
         );
  INV_X1 U7418 ( .A(n9736), .ZN(n5874) );
  INV_X1 U7419 ( .A(n9608), .ZN(n5863) );
  AND2_X2 U7420 ( .A1(n5864), .A2(n5863), .ZN(n9346) );
  INV_X1 U7421 ( .A(n9346), .ZN(n9323) );
  INV_X1 U7422 ( .A(n5865), .ZN(n5866) );
  NAND2_X1 U7423 ( .A1(n5866), .A2(n6462), .ZN(n5869) );
  INV_X1 U7424 ( .A(n6460), .ZN(n5867) );
  AND2_X1 U7425 ( .A1(n5867), .A2(n6500), .ZN(n5868) );
  AOI21_X1 U7426 ( .B1(n5869), .B2(n5868), .A(P1_U3086), .ZN(n5872) );
  INV_X1 U7427 ( .A(n6533), .ZN(n5870) );
  NAND2_X1 U7428 ( .A1(n5870), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9617) );
  INV_X1 U7429 ( .A(n9617), .ZN(n5871) );
  AOI22_X1 U7430 ( .A1(n9744), .A2(n9337), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n5873) );
  OAI21_X1 U7431 ( .B1(n5874), .B2(n9323), .A(n5873), .ZN(n5878) );
  NOR3_X1 U7432 ( .A1(n5876), .A2(n9354), .A3(n5875), .ZN(n5877) );
  AOI211_X1 U7433 ( .C1(n9742), .C2(n9351), .A(n5878), .B(n5877), .ZN(n5879)
         );
  OAI211_X1 U7434 ( .C1(n6469), .C2(n5881), .A(n5880), .B(n5879), .ZN(P1_U3220) );
  INV_X1 U7435 ( .A(n5883), .ZN(n5886) );
  INV_X1 U7436 ( .A(n5884), .ZN(n5885) );
  AOI21_X1 U7437 ( .B1(n5882), .B2(n5886), .A(n5885), .ZN(n5887) );
  INV_X1 U7438 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U7439 ( .A1(n5888), .A2(n5043), .ZN(n5894) );
  OAI22_X1 U7440 ( .A1(n6413), .A2(n9301), .B1(n9269), .B2(n9300), .ZN(n9769)
         );
  OAI22_X1 U7441 ( .A1(n9775), .A2(n9349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5889), .ZN(n5890) );
  AOI21_X1 U7442 ( .B1(n9769), .B2(n9346), .A(n5890), .ZN(n5891) );
  NAND2_X1 U7443 ( .A1(n5894), .A2(n5893), .ZN(P1_U3240) );
  NAND2_X1 U7444 ( .A1(n5898), .A2(n4416), .ZN(n6040) );
  NOR2_X1 U7445 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5902) );
  NAND4_X1 U7446 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(n5903)
         );
  INV_X1 U7447 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5909) );
  INV_X1 U7448 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5913) );
  INV_X1 U7449 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7450 ( .A1(n5927), .A2(n5040), .ZN(n5914) );
  XNOR2_X2 U7451 ( .A(n5914), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8022) );
  INV_X1 U7452 ( .A(n5915), .ZN(n5917) );
  NOR2_X1 U7453 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n5916) );
  NAND2_X1 U7454 ( .A1(n5917), .A2(n5916), .ZN(n9164) );
  XNOR2_X2 U7455 ( .A(n5918), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5920) );
  INV_X1 U7456 ( .A(n5920), .ZN(n9168) );
  NAND2_X1 U7457 ( .A1(n5951), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5925) );
  INV_X1 U7458 ( .A(n8022), .ZN(n5921) );
  INV_X1 U7459 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5919) );
  OR2_X1 U7460 ( .A1(n5971), .A2(n5919), .ZN(n5923) );
  NAND2_X1 U7461 ( .A1(n5994), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5922) );
  AND4_X2 U7462 ( .A1(n5925), .A2(n5924), .A3(n5923), .A4(n5922), .ZN(n6899)
         );
  INV_X1 U7463 ( .A(n6899), .ZN(n5940) );
  INV_X1 U7464 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5926) );
  NAND2_X1 U7465 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n5929) );
  AND2_X2 U7466 ( .A1(n5946), .A2(n9356), .ZN(n5963) );
  INV_X1 U7467 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7468 ( .A1(n5963), .A2(n5931), .ZN(n5939) );
  INV_X1 U7469 ( .A(n6511), .ZN(n5932) );
  NAND2_X1 U7470 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5933) );
  MUX2_X1 U7471 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5933), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n5936) );
  INV_X1 U7472 ( .A(n5934), .ZN(n5935) );
  INV_X1 U7473 ( .A(n6689), .ZN(n5937) );
  INV_X1 U7474 ( .A(n7137), .ZN(n10319) );
  NAND2_X1 U7475 ( .A1(n7137), .A2(n6899), .ZN(n8170) );
  INV_X1 U7476 ( .A(n6279), .ZN(n5948) );
  NAND2_X1 U7477 ( .A1(n5994), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5944) );
  NAND2_X1 U7478 ( .A1(n5970), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7479 ( .A1(n6991), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7480 ( .A1(n5951), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7481 ( .A1(n5212), .A2(SI_0_), .ZN(n5945) );
  XNOR2_X1 U7482 ( .A(n5945), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9172) );
  MUX2_X1 U7483 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9172), .S(n5946), .Z(n6911) );
  NAND2_X1 U7484 ( .A1(n6280), .A2(n6911), .ZN(n8167) );
  NAND2_X1 U7485 ( .A1(n5948), .A2(n5947), .ZN(n7127) );
  NAND2_X1 U7486 ( .A1(n7127), .A2(n8170), .ZN(n7225) );
  NAND2_X1 U7487 ( .A1(n6991), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7488 ( .A1(n5994), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5950) );
  NAND2_X1 U7489 ( .A1(n5970), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7490 ( .A1(n5951), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5952) );
  NAND3_X2 U7491 ( .A1(n5954), .A2(n5953), .A3(n5952), .ZN(n8400) );
  INV_X2 U7492 ( .A(n8400), .ZN(n7022) );
  NAND2_X1 U7493 ( .A1(n4418), .A2(n5955), .ZN(n5961) );
  NAND2_X1 U7494 ( .A1(n5963), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5960) );
  INV_X1 U7495 ( .A(n6711), .ZN(n5959) );
  INV_X1 U7496 ( .A(n7232), .ZN(n10324) );
  NAND2_X1 U7497 ( .A1(n7232), .A2(n8400), .ZN(n8178) );
  INV_X1 U7498 ( .A(n8171), .ZN(n7227) );
  NAND2_X1 U7499 ( .A1(n7225), .A2(n7227), .ZN(n7224) );
  NAND2_X1 U7500 ( .A1(n7224), .A2(n8177), .ZN(n5976) );
  NAND2_X1 U7501 ( .A1(n5962), .A2(n6504), .ZN(n5969) );
  NAND2_X1 U7502 ( .A1(n6241), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7503 ( .A1(n5965), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5964) );
  MUX2_X1 U7504 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5964), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5966) );
  OR2_X1 U7505 ( .A1(n5965), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n5984) );
  AND2_X1 U7506 ( .A1(n5966), .A2(n5984), .ZN(n6754) );
  NAND2_X1 U7507 ( .A1(n6165), .A2(n6754), .ZN(n5967) );
  NAND2_X1 U7508 ( .A1(n5951), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5975) );
  INV_X1 U7509 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U7510 ( .A1(n5994), .A2(n7256), .ZN(n5974) );
  NAND2_X1 U7511 ( .A1(n6271), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5973) );
  INV_X4 U7512 ( .A(n5971), .ZN(n6991) );
  NAND2_X1 U7513 ( .A1(n6991), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7514 ( .A1(n10331), .A2(n8398), .ZN(n8197) );
  NAND2_X1 U7515 ( .A1(n5951), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5981) );
  NAND2_X1 U7516 ( .A1(n6991), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5980) );
  NOR2_X1 U7517 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5996) );
  INV_X1 U7518 ( .A(n5996), .ZN(n5997) );
  NAND2_X1 U7519 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5977) );
  NAND2_X1 U7520 ( .A1(n5997), .A2(n5977), .ZN(n7247) );
  NAND2_X1 U7521 ( .A1(n4414), .A2(n7247), .ZN(n5979) );
  NAND2_X1 U7522 ( .A1(n6271), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5978) );
  NAND4_X1 U7523 ( .A1(n5981), .A2(n5980), .A3(n5979), .A4(n5978), .ZN(n8397)
         );
  INV_X1 U7524 ( .A(n8397), .ZN(n7393) );
  NAND2_X1 U7525 ( .A1(n5962), .A2(n6515), .ZN(n5989) );
  NAND2_X1 U7526 ( .A1(n6241), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n5988) );
  NAND2_X1 U7527 ( .A1(n5984), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5983) );
  MUX2_X1 U7528 ( .A(n5983), .B(P2_IR_REG_31__SCAN_IN), .S(n5982), .Z(n5986)
         );
  INV_X1 U7529 ( .A(n6006), .ZN(n5985) );
  NAND2_X1 U7530 ( .A1(n6165), .A2(n6783), .ZN(n5987) );
  NAND2_X1 U7531 ( .A1(n7393), .A2(n7248), .ZN(n8199) );
  NAND2_X1 U7532 ( .A1(n10337), .A2(n8397), .ZN(n7371) );
  NAND2_X1 U7533 ( .A1(n5962), .A2(n6513), .ZN(n5993) );
  NAND2_X1 U7534 ( .A1(n6241), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n5992) );
  OR2_X1 U7535 ( .A1(n6006), .A2(n6099), .ZN(n5990) );
  NAND2_X1 U7536 ( .A1(n6165), .A2(n6799), .ZN(n5991) );
  NAND2_X1 U7537 ( .A1(n4411), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7538 ( .A1(n6991), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6001) );
  INV_X1 U7539 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5995) );
  NAND2_X1 U7540 ( .A1(n5996), .A2(n5995), .ZN(n6010) );
  NAND2_X1 U7541 ( .A1(n5997), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7542 ( .A1(n6010), .A2(n5998), .ZN(n7384) );
  NAND2_X1 U7543 ( .A1(n4414), .A2(n7384), .ZN(n6000) );
  NAND2_X1 U7544 ( .A1(n6271), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5999) );
  NAND4_X1 U7545 ( .A1(n6002), .A2(n6001), .A3(n6000), .A4(n5999), .ZN(n8396)
         );
  NAND2_X1 U7546 ( .A1(n7467), .A2(n8396), .ZN(n8202) );
  AND2_X1 U7547 ( .A1(n7371), .A2(n8202), .ZN(n8187) );
  NAND2_X1 U7548 ( .A1(n7372), .A2(n8187), .ZN(n6003) );
  NAND2_X1 U7549 ( .A1(n7490), .A2(n7470), .ZN(n8198) );
  NAND2_X1 U7550 ( .A1(n6241), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6009) );
  INV_X1 U7551 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7552 ( .A1(n6006), .A2(n6005), .ZN(n6016) );
  NAND2_X1 U7553 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7554 ( .A(n6007), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10254) );
  NAND2_X1 U7555 ( .A1(n6165), .A2(n10254), .ZN(n6008) );
  OAI211_X1 U7556 ( .C1(n6004), .C2(n6525), .A(n6009), .B(n6008), .ZN(n7492)
         );
  INV_X1 U7557 ( .A(n7492), .ZN(n10342) );
  NAND2_X1 U7558 ( .A1(n6991), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6015) );
  NAND2_X1 U7559 ( .A1(n4411), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7560 ( .A1(n6010), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6011) );
  NAND2_X1 U7561 ( .A1(n6023), .A2(n6011), .ZN(n7474) );
  NAND2_X1 U7562 ( .A1(n4413), .A2(n7474), .ZN(n6013) );
  NAND2_X1 U7563 ( .A1(n6271), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6012) );
  INV_X1 U7564 ( .A(n7614), .ZN(n8395) );
  AND2_X1 U7565 ( .A1(n10342), .A2(n8395), .ZN(n8189) );
  INV_X1 U7566 ( .A(n8189), .ZN(n8203) );
  NAND2_X1 U7567 ( .A1(n7614), .A2(n7492), .ZN(n8193) );
  NAND2_X1 U7568 ( .A1(n5962), .A2(n6506), .ZN(n6022) );
  NAND2_X1 U7569 ( .A1(n6241), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6021) );
  OR2_X1 U7570 ( .A1(n6016), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n6017) );
  NAND2_X1 U7571 ( .A1(n6017), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6018) );
  NAND2_X1 U7572 ( .A1(n6018), .A2(n8937), .ZN(n6029) );
  OR2_X1 U7573 ( .A1(n6018), .A2(n8937), .ZN(n6019) );
  NAND2_X1 U7574 ( .A1(n6165), .A2(n10269), .ZN(n6020) );
  NAND2_X1 U7575 ( .A1(n4411), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7576 ( .A1(n6271), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6027) );
  INV_X1 U7577 ( .A(n6032), .ZN(n6033) );
  NAND2_X1 U7578 ( .A1(n6023), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6024) );
  NAND2_X1 U7579 ( .A1(n6033), .A2(n6024), .ZN(n7612) );
  NAND2_X1 U7580 ( .A1(n4413), .A2(n7612), .ZN(n6026) );
  NAND2_X1 U7581 ( .A1(n6991), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6025) );
  NAND4_X1 U7582 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n8394)
         );
  NAND2_X1 U7583 ( .A1(n10348), .A2(n8394), .ZN(n7685) );
  INV_X1 U7584 ( .A(n8394), .ZN(n7734) );
  INV_X1 U7585 ( .A(n10348), .ZN(n7613) );
  NAND2_X1 U7586 ( .A1(n7734), .A2(n7613), .ZN(n8212) );
  NAND2_X1 U7587 ( .A1(n6029), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6030) );
  XNOR2_X1 U7588 ( .A(n6030), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7193) );
  AOI22_X1 U7589 ( .A1(n6241), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6165), .B2(
        n7193), .ZN(n6031) );
  INV_X1 U7590 ( .A(n7743), .ZN(n10352) );
  NAND2_X1 U7591 ( .A1(n6991), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6038) );
  NAND2_X1 U7592 ( .A1(n4411), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6037) );
  INV_X1 U7593 ( .A(n6047), .ZN(n6048) );
  NAND2_X1 U7594 ( .A1(n6033), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U7595 ( .A1(n6048), .A2(n6034), .ZN(n7729) );
  NAND2_X1 U7596 ( .A1(n4414), .A2(n7729), .ZN(n6036) );
  NAND2_X1 U7597 ( .A1(n6271), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6035) );
  AND2_X1 U7598 ( .A1(n10352), .A2(n8393), .ZN(n8194) );
  INV_X1 U7599 ( .A(n8194), .ZN(n7684) );
  AND2_X1 U7600 ( .A1(n7684), .A2(n7685), .ZN(n8209) );
  NAND2_X1 U7601 ( .A1(n7743), .A2(n7750), .ZN(n8213) );
  INV_X1 U7602 ( .A(n8213), .ZN(n6039) );
  NAND2_X1 U7603 ( .A1(n6531), .A2(n5962), .ZN(n6045) );
  NAND2_X1 U7604 ( .A1(n6040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6041) );
  MUX2_X1 U7605 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6041), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n6043) );
  NOR2_X1 U7606 ( .A1(n6040), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6063) );
  INV_X1 U7607 ( .A(n6063), .ZN(n6042) );
  NAND2_X1 U7608 ( .A1(n6043), .A2(n6042), .ZN(n7313) );
  INV_X1 U7609 ( .A(n7313), .ZN(n7203) );
  AOI22_X1 U7610 ( .A1(n6241), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6165), .B2(
        n7203), .ZN(n6044) );
  NAND2_X1 U7611 ( .A1(n6045), .A2(n6044), .ZN(n10313) );
  INV_X1 U7612 ( .A(n10313), .ZN(n7766) );
  NAND2_X1 U7613 ( .A1(n4411), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7614 ( .A1(n6048), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6049) );
  NAND2_X1 U7615 ( .A1(n6057), .A2(n6049), .ZN(n10315) );
  NAND2_X1 U7616 ( .A1(n4414), .A2(n10315), .ZN(n6052) );
  NAND2_X1 U7617 ( .A1(n6271), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6051) );
  NAND2_X1 U7618 ( .A1(n6991), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6050) );
  NAND2_X1 U7619 ( .A1(n10313), .A2(n7773), .ZN(n8214) );
  NAND2_X1 U7620 ( .A1(n6546), .A2(n5962), .ZN(n6056) );
  OR2_X1 U7621 ( .A1(n6063), .A2(n6099), .ZN(n6054) );
  XNOR2_X1 U7622 ( .A(n6054), .B(P2_IR_REG_10__SCAN_IN), .ZN(n7551) );
  AOI22_X1 U7623 ( .A1(n6241), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6165), .B2(
        n7551), .ZN(n6055) );
  NAND2_X1 U7624 ( .A1(n6056), .A2(n6055), .ZN(n7924) );
  NAND2_X1 U7625 ( .A1(n4411), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6062) );
  NAND2_X1 U7626 ( .A1(n6991), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7627 ( .A1(n6057), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7628 ( .A1(n6067), .A2(n6058), .ZN(n7918) );
  NAND2_X1 U7629 ( .A1(n4414), .A2(n7918), .ZN(n6060) );
  NAND2_X1 U7630 ( .A1(n6271), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6059) );
  OR2_X1 U7631 ( .A1(n7924), .A2(n7754), .ZN(n8222) );
  NAND2_X1 U7632 ( .A1(n6561), .A2(n5962), .ZN(n6066) );
  NAND2_X1 U7633 ( .A1(n6063), .A2(n8893), .ZN(n6074) );
  NAND2_X1 U7634 ( .A1(n6074), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6064) );
  XNOR2_X1 U7635 ( .A(n6064), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7562) );
  AOI22_X1 U7636 ( .A1(n6241), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6165), .B2(
        n7562), .ZN(n6065) );
  NAND2_X1 U7637 ( .A1(n6066), .A2(n6065), .ZN(n8112) );
  NAND2_X1 U7638 ( .A1(n6991), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6072) );
  NAND2_X1 U7639 ( .A1(n4411), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6071) );
  NAND2_X1 U7640 ( .A1(n6067), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6068) );
  NAND2_X1 U7641 ( .A1(n6078), .A2(n6068), .ZN(n8100) );
  NAND2_X1 U7642 ( .A1(n4413), .A2(n8100), .ZN(n6070) );
  NAND2_X1 U7643 ( .A1(n6271), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7644 ( .A1(n8112), .A2(n7922), .ZN(n8223) );
  NAND2_X1 U7645 ( .A1(n7924), .A2(n7754), .ZN(n8215) );
  AND2_X1 U7646 ( .A1(n8223), .A2(n8215), .ZN(n8227) );
  NAND2_X1 U7647 ( .A1(n7805), .A2(n8227), .ZN(n6073) );
  NAND2_X1 U7648 ( .A1(n6073), .A2(n8225), .ZN(n7873) );
  NAND2_X1 U7649 ( .A1(n6592), .A2(n5962), .ZN(n6077) );
  NAND2_X1 U7650 ( .A1(n6085), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6075) );
  XNOR2_X1 U7651 ( .A(n6075), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7834) );
  AOI22_X1 U7652 ( .A1(n6241), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6165), .B2(
        n7834), .ZN(n6076) );
  NAND2_X1 U7653 ( .A1(n6991), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U7654 ( .A1(n4411), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6082) );
  INV_X1 U7655 ( .A(n6090), .ZN(n6091) );
  NAND2_X1 U7656 ( .A1(n6078), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7657 ( .A1(n6091), .A2(n6079), .ZN(n7964) );
  NAND2_X1 U7658 ( .A1(n4413), .A2(n7964), .ZN(n6081) );
  NAND2_X1 U7659 ( .A1(n6271), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6080) );
  NAND2_X1 U7660 ( .A1(n7969), .A2(n8104), .ZN(n8233) );
  NAND2_X1 U7661 ( .A1(n7873), .A2(n8231), .ZN(n6084) );
  NAND2_X1 U7662 ( .A1(n6084), .A2(n8232), .ZN(n7927) );
  NAND2_X1 U7663 ( .A1(n6732), .A2(n5962), .ZN(n6088) );
  NOR2_X1 U7664 ( .A1(n6085), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6101) );
  OR2_X1 U7665 ( .A1(n6101), .A2(n6099), .ZN(n6086) );
  XNOR2_X1 U7666 ( .A(n6086), .B(P2_IR_REG_13__SCAN_IN), .ZN(n8438) );
  AOI22_X1 U7667 ( .A1(n6241), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6165), .B2(
        n8438), .ZN(n6087) );
  NAND2_X1 U7668 ( .A1(n4411), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7669 ( .A1(n6271), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6095) );
  INV_X1 U7670 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7671 ( .A1(n6090), .A2(n6089), .ZN(n6108) );
  NAND2_X1 U7672 ( .A1(n6091), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7673 ( .A1(n6108), .A2(n6092), .ZN(n8736) );
  NAND2_X1 U7674 ( .A1(n4413), .A2(n8736), .ZN(n6094) );
  NAND2_X1 U7675 ( .A1(n6991), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7676 ( .A1(n7936), .A2(n8720), .ZN(n8239) );
  NAND2_X1 U7677 ( .A1(n8713), .A2(n8239), .ZN(n7928) );
  NAND2_X1 U7678 ( .A1(n7927), .A2(n7928), .ZN(n6098) );
  OR2_X1 U7679 ( .A1(n7936), .A2(n8235), .ZN(n6097) );
  NAND2_X1 U7680 ( .A1(n6098), .A2(n6097), .ZN(n8726) );
  NAND2_X1 U7681 ( .A1(n6831), .A2(n5962), .ZN(n6107) );
  INV_X1 U7682 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6100) );
  AOI21_X1 U7683 ( .B1(n6101), .B2(n6100), .A(n6099), .ZN(n6102) );
  NAND2_X1 U7684 ( .A1(n6102), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n6105) );
  INV_X1 U7685 ( .A(n6102), .ZN(n6104) );
  INV_X1 U7686 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6103) );
  NAND2_X1 U7687 ( .A1(n6104), .A2(n6103), .ZN(n6115) );
  AOI22_X1 U7688 ( .A1(n6241), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6165), .B2(
        n8463), .ZN(n6106) );
  NAND2_X1 U7689 ( .A1(n6991), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7690 ( .A1(n4411), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6112) );
  NAND2_X1 U7691 ( .A1(n6108), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7692 ( .A1(n6119), .A2(n6109), .ZN(n8723) );
  NAND2_X1 U7693 ( .A1(n4414), .A2(n8723), .ZN(n6111) );
  NAND2_X1 U7694 ( .A1(n6271), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6110) );
  NAND4_X1 U7695 ( .A1(n6113), .A2(n6112), .A3(n6111), .A4(n6110), .ZN(n8388)
         );
  XNOR2_X1 U7696 ( .A(n9159), .B(n8388), .ZN(n8727) );
  NAND2_X1 U7697 ( .A1(n8726), .A2(n8727), .ZN(n6114) );
  INV_X1 U7698 ( .A(n8388), .ZN(n8242) );
  OR2_X1 U7699 ( .A1(n9159), .A2(n8242), .ZN(n8244) );
  NAND2_X1 U7700 ( .A1(n6114), .A2(n8244), .ZN(n7939) );
  NAND2_X1 U7701 ( .A1(n6886), .A2(n5962), .ZN(n6118) );
  NAND2_X1 U7702 ( .A1(n6115), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6116) );
  XNOR2_X1 U7703 ( .A(n6116), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8490) );
  AOI22_X1 U7704 ( .A1(n6241), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6165), .B2(
        n8490), .ZN(n6117) );
  NAND2_X1 U7705 ( .A1(n6991), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7706 ( .A1(n4411), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6123) );
  INV_X1 U7707 ( .A(n6143), .ZN(n6141) );
  NAND2_X1 U7708 ( .A1(n6119), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6120) );
  NAND2_X1 U7709 ( .A1(n6141), .A2(n6120), .ZN(n8142) );
  NAND2_X1 U7710 ( .A1(n4414), .A2(n8142), .ZN(n6122) );
  NAND2_X1 U7711 ( .A1(n6271), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7712 ( .A1(n7980), .A2(n7981), .ZN(n8247) );
  NAND2_X1 U7713 ( .A1(n7939), .A2(n8339), .ZN(n6125) );
  NAND2_X1 U7714 ( .A1(n6125), .A2(n8248), .ZN(n8704) );
  NAND2_X1 U7715 ( .A1(n6913), .A2(n5962), .ZN(n6131) );
  NOR2_X1 U7716 ( .A1(n6126), .A2(n6099), .ZN(n6127) );
  MUX2_X1 U7717 ( .A(n6099), .B(n6127), .S(P2_IR_REG_16__SCAN_IN), .Z(n6129)
         );
  AND2_X1 U7718 ( .A1(n6126), .A2(n6128), .ZN(n6137) );
  AOI22_X1 U7719 ( .A1(n6241), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6165), .B2(
        n8523), .ZN(n6130) );
  NAND2_X1 U7720 ( .A1(n6991), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7721 ( .A1(n4411), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6134) );
  XNOR2_X1 U7722 ( .A(n6141), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U7723 ( .A1(n4414), .A2(n8710), .ZN(n6133) );
  NAND2_X1 U7724 ( .A1(n6271), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7725 ( .A1(n9152), .A2(n8074), .ZN(n8253) );
  NAND2_X1 U7726 ( .A1(n8254), .A2(n8253), .ZN(n8252) );
  NAND2_X1 U7727 ( .A1(n8704), .A2(n8706), .ZN(n6136) );
  NAND2_X2 U7728 ( .A1(n6136), .A2(n8254), .ZN(n8695) );
  NAND2_X1 U7729 ( .A1(n7077), .A2(n5962), .ZN(n6140) );
  OR2_X1 U7730 ( .A1(n6137), .A2(n6099), .ZN(n6138) );
  XNOR2_X1 U7731 ( .A(n6138), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8527) );
  AOI22_X1 U7732 ( .A1(n6241), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6165), .B2(
        n8527), .ZN(n6139) );
  NAND2_X1 U7733 ( .A1(n6991), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6148) );
  NAND2_X1 U7734 ( .A1(n4411), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6147) );
  OAI21_X1 U7735 ( .B1(n6141), .B2(P2_REG3_REG_16__SCAN_IN), .A(
        P2_REG3_REG_17__SCAN_IN), .ZN(n6144) );
  NOR2_X1 U7736 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_REG3_REG_17__SCAN_IN), 
        .ZN(n6142) );
  INV_X1 U7737 ( .A(n6155), .ZN(n6156) );
  NAND2_X1 U7738 ( .A1(n6144), .A2(n6156), .ZN(n8697) );
  NAND2_X1 U7739 ( .A1(n4413), .A2(n8697), .ZN(n6146) );
  NAND2_X1 U7740 ( .A1(n6271), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6145) );
  OR2_X1 U7741 ( .A1(n9076), .A2(n8675), .ZN(n8260) );
  NAND2_X1 U7742 ( .A1(n9076), .A2(n8675), .ZN(n8680) );
  NAND2_X1 U7743 ( .A1(n7115), .A2(n5962), .ZN(n6153) );
  INV_X1 U7744 ( .A(n6149), .ZN(n6150) );
  NAND2_X1 U7745 ( .A1(n6150), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6151) );
  XNOR2_X1 U7746 ( .A(n6151), .B(P2_IR_REG_18__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U7747 ( .A1(n5963), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6165), .B2(
        n10092), .ZN(n6152) );
  NAND2_X1 U7748 ( .A1(n4411), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6161) );
  NAND2_X1 U7749 ( .A1(n6991), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n6160) );
  INV_X1 U7750 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7751 ( .A1(n6156), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6157) );
  NAND2_X1 U7752 ( .A1(n6168), .A2(n6157), .ZN(n8684) );
  NAND2_X1 U7753 ( .A1(n4413), .A2(n8684), .ZN(n6159) );
  NAND2_X1 U7754 ( .A1(n6271), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6158) );
  AND2_X1 U7755 ( .A1(n8683), .A2(n8663), .ZN(n8265) );
  INV_X1 U7756 ( .A(n8265), .ZN(n8259) );
  NAND2_X1 U7757 ( .A1(n8263), .A2(n8259), .ZN(n8682) );
  INV_X1 U7758 ( .A(n8680), .ZN(n6162) );
  NOR2_X1 U7759 ( .A1(n8682), .A2(n6162), .ZN(n6163) );
  NAND2_X1 U7760 ( .A1(n7299), .A2(n5962), .ZN(n6167) );
  NAND2_X1 U7761 ( .A1(n4470), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6164) );
  AOI22_X1 U7762 ( .A1(n6241), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8509), .B2(
        n6165), .ZN(n6166) );
  NAND2_X1 U7763 ( .A1(n4411), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6173) );
  NAND2_X1 U7764 ( .A1(n6991), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7765 ( .A1(n6168), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7766 ( .A1(n6176), .A2(n6169), .ZN(n8668) );
  NAND2_X1 U7767 ( .A1(n4414), .A2(n8668), .ZN(n6171) );
  NAND2_X1 U7768 ( .A1(n6271), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6170) );
  NAND4_X1 U7769 ( .A1(n6173), .A2(n6172), .A3(n6171), .A4(n6170), .ZN(n8649)
         );
  AND2_X1 U7770 ( .A1(n9139), .A2(n8649), .ZN(n8159) );
  NAND2_X1 U7771 ( .A1(n8669), .A2(n8677), .ZN(n8267) );
  NAND2_X1 U7772 ( .A1(n7378), .A2(n5962), .ZN(n6175) );
  NAND2_X1 U7773 ( .A1(n5963), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6174) );
  INV_X1 U7774 ( .A(n6185), .ZN(n6186) );
  NAND2_X1 U7775 ( .A1(n6176), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6177) );
  NAND2_X1 U7776 ( .A1(n6186), .A2(n6177), .ZN(n8653) );
  NAND2_X1 U7777 ( .A1(n8653), .A2(n4413), .ZN(n6181) );
  NAND2_X1 U7778 ( .A1(n4411), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7779 ( .A1(n6991), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7780 ( .A1(n6271), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7781 ( .A1(n7602), .A2(n5962), .ZN(n6183) );
  NAND2_X1 U7782 ( .A1(n5963), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6182) );
  INV_X1 U7783 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6184) );
  INV_X1 U7784 ( .A(n6197), .ZN(n6198) );
  NAND2_X1 U7785 ( .A1(n6186), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6187) );
  NAND2_X1 U7786 ( .A1(n6198), .A2(n6187), .ZN(n8640) );
  NAND2_X1 U7787 ( .A1(n8640), .A2(n4414), .ZN(n6192) );
  NAND2_X1 U7788 ( .A1(n4411), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6189) );
  NAND2_X1 U7789 ( .A1(n6991), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6188) );
  AND2_X1 U7790 ( .A1(n6189), .A2(n6188), .ZN(n6191) );
  NAND2_X1 U7791 ( .A1(n6271), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6190) );
  NAND2_X1 U7792 ( .A1(n8052), .A2(n8624), .ZN(n8152) );
  NAND2_X1 U7793 ( .A1(n9133), .A2(n8662), .ZN(n8637) );
  NAND2_X1 U7794 ( .A1(n8152), .A2(n8637), .ZN(n8275) );
  INV_X1 U7795 ( .A(n8275), .ZN(n6193) );
  NAND2_X1 U7796 ( .A1(n8636), .A2(n6193), .ZN(n6194) );
  NAND2_X1 U7797 ( .A1(n6194), .A2(n8155), .ZN(n8625) );
  NAND2_X1 U7798 ( .A1(n7646), .A2(n5962), .ZN(n6196) );
  NAND2_X1 U7799 ( .A1(n5963), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6195) );
  NAND2_X1 U7800 ( .A1(n6198), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6199) );
  NAND2_X1 U7801 ( .A1(n6205), .A2(n6199), .ZN(n8628) );
  NAND2_X1 U7802 ( .A1(n8628), .A2(n4413), .ZN(n6202) );
  AOI22_X1 U7803 ( .A1(n6991), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n4411), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n6201) );
  NAND2_X1 U7804 ( .A1(n6271), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7805 ( .A1(n8627), .A2(n8635), .ZN(n8276) );
  NAND2_X1 U7806 ( .A1(n7657), .A2(n5962), .ZN(n6204) );
  NAND2_X1 U7807 ( .A1(n5963), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6203) );
  NAND2_X1 U7808 ( .A1(n6205), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7809 ( .A1(n6212), .A2(n6206), .ZN(n8618) );
  NAND2_X1 U7810 ( .A1(n8618), .A2(n4413), .ZN(n6209) );
  AOI22_X1 U7811 ( .A1(n6271), .A2(P2_REG1_REG_23__SCAN_IN), .B1(n4411), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7812 ( .A1(n6991), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7813 ( .A1(n7679), .A2(n5962), .ZN(n6211) );
  NAND2_X1 U7814 ( .A1(n5963), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6210) );
  NAND2_X1 U7815 ( .A1(n6212), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6213) );
  NAND2_X1 U7816 ( .A1(n6222), .A2(n6213), .ZN(n8605) );
  NAND2_X1 U7817 ( .A1(n8605), .A2(n4414), .ZN(n6218) );
  INV_X1 U7818 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8768) );
  INV_X1 U7819 ( .A(n6271), .ZN(n6994) );
  NAND2_X1 U7820 ( .A1(n4411), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7821 ( .A1(n6991), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6214) );
  OAI211_X1 U7822 ( .C1(n8768), .C2(n6994), .A(n6215), .B(n6214), .ZN(n6216)
         );
  INV_X1 U7823 ( .A(n6216), .ZN(n6217) );
  AND2_X1 U7824 ( .A1(n8083), .A2(n8591), .ZN(n8280) );
  INV_X1 U7825 ( .A(n8280), .ZN(n8363) );
  NAND2_X1 U7826 ( .A1(n9119), .A2(n8623), .ZN(n8598) );
  AND2_X1 U7827 ( .A1(n8363), .A2(n8598), .ZN(n8283) );
  NAND2_X1 U7828 ( .A1(n8599), .A2(n8283), .ZN(n6219) );
  NAND2_X1 U7829 ( .A1(n6219), .A2(n8364), .ZN(n8586) );
  NAND2_X1 U7830 ( .A1(n7724), .A2(n4418), .ZN(n6221) );
  NAND2_X1 U7831 ( .A1(n5963), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6220) );
  INV_X1 U7832 ( .A(n6233), .ZN(n6234) );
  NAND2_X1 U7833 ( .A1(n6222), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U7834 ( .A1(n6234), .A2(n6223), .ZN(n8592) );
  NAND2_X1 U7835 ( .A1(n8592), .A2(n4414), .ZN(n6228) );
  INV_X1 U7836 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n8762) );
  NAND2_X1 U7837 ( .A1(n6991), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7838 ( .A1(n4411), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6224) );
  OAI211_X1 U7839 ( .C1(n8762), .C2(n6994), .A(n6225), .B(n6224), .ZN(n6226)
         );
  INV_X1 U7840 ( .A(n6226), .ZN(n6227) );
  NAND2_X1 U7841 ( .A1(n8761), .A2(n8604), .ZN(n8290) );
  NAND2_X1 U7842 ( .A1(n8586), .A2(n8290), .ZN(n6229) );
  NAND2_X1 U7843 ( .A1(n6229), .A2(n8289), .ZN(n8579) );
  NAND2_X1 U7844 ( .A1(n7867), .A2(n4418), .ZN(n6231) );
  NAND2_X1 U7845 ( .A1(n5963), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6230) );
  INV_X1 U7846 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6232) );
  INV_X1 U7847 ( .A(n6245), .ZN(n6246) );
  NAND2_X1 U7848 ( .A1(n6234), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6235) );
  NAND2_X1 U7849 ( .A1(n6246), .A2(n6235), .ZN(n8581) );
  NAND2_X1 U7850 ( .A1(n8581), .A2(n4413), .ZN(n6240) );
  INV_X1 U7851 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U7852 ( .A1(n6991), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7853 ( .A1(n4411), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6236) );
  OAI211_X1 U7854 ( .C1(n8758), .C2(n6994), .A(n6237), .B(n6236), .ZN(n6238)
         );
  INV_X1 U7855 ( .A(n6238), .ZN(n6239) );
  NAND2_X1 U7856 ( .A1(n8129), .A2(n8590), .ZN(n8294) );
  NAND2_X1 U7857 ( .A1(n7885), .A2(n5962), .ZN(n6243) );
  NAND2_X1 U7858 ( .A1(n6241), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6242) );
  INV_X1 U7859 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6244) );
  INV_X1 U7860 ( .A(n6254), .ZN(n6255) );
  NAND2_X1 U7861 ( .A1(n6246), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7862 ( .A1(n6255), .A2(n6247), .ZN(n8572) );
  INV_X1 U7863 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U7864 ( .A1(n6271), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7865 ( .A1(n4411), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6248) );
  OAI211_X1 U7866 ( .C1(n5971), .C2(n8571), .A(n6249), .B(n6248), .ZN(n6250)
         );
  AOI21_X1 U7867 ( .B1(n8572), .B2(n4413), .A(n6250), .ZN(n8577) );
  NAND2_X1 U7868 ( .A1(n9103), .A2(n8577), .ZN(n8147) );
  NAND2_X1 U7869 ( .A1(n7908), .A2(n5962), .ZN(n6253) );
  NAND2_X1 U7870 ( .A1(n5963), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6252) );
  INV_X1 U7871 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U7872 ( .A1(n6254), .A2(n8014), .ZN(n8540) );
  NAND2_X1 U7873 ( .A1(n6255), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U7874 ( .A1(n8540), .A2(n6256), .ZN(n8562) );
  NAND2_X1 U7875 ( .A1(n8562), .A2(n4413), .ZN(n6261) );
  INV_X1 U7876 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U7877 ( .A1(n4411), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7878 ( .A1(n6271), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6257) );
  OAI211_X1 U7879 ( .C1(n8830), .C2(n5971), .A(n6258), .B(n6257), .ZN(n6259)
         );
  INV_X1 U7880 ( .A(n6259), .ZN(n6260) );
  INV_X1 U7881 ( .A(n8569), .ZN(n8028) );
  NOR2_X1 U7882 ( .A1(n9097), .A2(n8028), .ZN(n6262) );
  NAND2_X1 U7883 ( .A1(n6264), .A2(n6263), .ZN(n6266) );
  MUX2_X1 U7884 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n4525), .Z(n8297) );
  NAND2_X2 U7885 ( .A1(n8300), .A2(n6268), .ZN(n6415) );
  NAND2_X1 U7886 ( .A1(n5963), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6269) );
  INV_X1 U7887 ( .A(n4414), .ZN(n6270) );
  OR2_X1 U7888 ( .A1(n8540), .A2(n6270), .ZN(n6997) );
  INV_X1 U7889 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U7890 ( .A1(n6271), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U7891 ( .A1(n4411), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6272) );
  OAI211_X1 U7892 ( .C1(n5971), .C2(n9039), .A(n6273), .B(n6272), .ZN(n6274)
         );
  INV_X1 U7893 ( .A(n6274), .ZN(n6275) );
  NAND2_X1 U7894 ( .A1(n6376), .A2(n8384), .ZN(n8306) );
  XNOR2_X1 U7895 ( .A(n8335), .B(n8368), .ZN(n8549) );
  NAND2_X1 U7896 ( .A1(n6276), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7897 ( .A1(n8329), .A2(n8509), .ZN(n6878) );
  NAND2_X1 U7898 ( .A1(n4471), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6277) );
  OR2_X1 U7899 ( .A1(n6878), .A2(n8379), .ZN(n10361) );
  INV_X1 U7900 ( .A(n8662), .ZN(n8387) );
  INV_X1 U7901 ( .A(n6280), .ZN(n7132) );
  NAND2_X1 U7902 ( .A1(n7132), .A2(n6911), .ZN(n7130) );
  NAND2_X1 U7903 ( .A1(n8342), .A2(n7130), .ZN(n7129) );
  NAND2_X1 U7904 ( .A1(n10319), .A2(n6899), .ZN(n7226) );
  NAND2_X1 U7905 ( .A1(n7129), .A2(n7226), .ZN(n6281) );
  NAND2_X1 U7906 ( .A1(n6281), .A2(n8171), .ZN(n7229) );
  NAND2_X1 U7907 ( .A1(n7232), .A2(n7022), .ZN(n6282) );
  NAND2_X1 U7908 ( .A1(n7229), .A2(n6282), .ZN(n7254) );
  NAND2_X1 U7909 ( .A1(n7257), .A2(n8398), .ZN(n6283) );
  NAND2_X1 U7910 ( .A1(n7254), .A2(n6283), .ZN(n6286) );
  NAND2_X1 U7911 ( .A1(n10331), .A2(n6284), .ZN(n6285) );
  AND2_X1 U7912 ( .A1(n10337), .A2(n7393), .ZN(n6288) );
  NAND2_X1 U7913 ( .A1(n7248), .A2(n8397), .ZN(n6287) );
  NOR2_X1 U7914 ( .A1(n7467), .A2(n7490), .ZN(n6290) );
  NAND2_X1 U7915 ( .A1(n7467), .A2(n7490), .ZN(n6289) );
  AND2_X1 U7916 ( .A1(n10342), .A2(n7614), .ZN(n6291) );
  OR2_X1 U7917 ( .A1(n8206), .A2(n4443), .ZN(n6292) );
  OR2_X1 U7918 ( .A1(n7592), .A2(n6292), .ZN(n6296) );
  NAND2_X1 U7919 ( .A1(n10348), .A2(n7734), .ZN(n7688) );
  NAND2_X1 U7920 ( .A1(n10352), .A2(n7750), .ZN(n6293) );
  AND2_X1 U7921 ( .A1(n7688), .A2(n6293), .ZN(n6294) );
  OR2_X1 U7922 ( .A1(n4443), .A2(n6294), .ZN(n6295) );
  NAND2_X1 U7923 ( .A1(n6296), .A2(n6295), .ZN(n7760) );
  NAND2_X1 U7924 ( .A1(n10313), .A2(n8392), .ZN(n6297) );
  NAND2_X1 U7925 ( .A1(n7760), .A2(n6297), .ZN(n6299) );
  OR2_X1 U7926 ( .A1(n10313), .A2(n8392), .ZN(n6298) );
  NAND2_X1 U7927 ( .A1(n6299), .A2(n6298), .ZN(n7770) );
  NAND2_X1 U7928 ( .A1(n7924), .A2(n8391), .ZN(n6300) );
  NAND2_X1 U7929 ( .A1(n7770), .A2(n6300), .ZN(n6302) );
  OR2_X1 U7930 ( .A1(n7924), .A2(n8391), .ZN(n6301) );
  NAND2_X1 U7931 ( .A1(n6302), .A2(n6301), .ZN(n7807) );
  INV_X1 U7932 ( .A(n7922), .ZN(n8390) );
  OR2_X1 U7933 ( .A1(n8112), .A2(n8390), .ZN(n6303) );
  INV_X1 U7934 ( .A(n8727), .ZN(n8715) );
  NAND2_X1 U7935 ( .A1(n7969), .A2(n8389), .ZN(n7929) );
  NAND4_X1 U7936 ( .A1(n7930), .A2(n8715), .A3(n8239), .A4(n7929), .ZN(n6306)
         );
  OAI22_X1 U7937 ( .A1(n8727), .A2(n8713), .B1(n8388), .B2(n9159), .ZN(n6304)
         );
  INV_X1 U7938 ( .A(n6304), .ZN(n6305) );
  NAND2_X1 U7939 ( .A1(n6306), .A2(n6305), .ZN(n7940) );
  NAND2_X1 U7940 ( .A1(n7980), .A2(n8718), .ZN(n6307) );
  NAND2_X1 U7941 ( .A1(n8689), .A2(n8696), .ZN(n6309) );
  NAND2_X1 U7942 ( .A1(n9076), .A2(n8707), .ZN(n6308) );
  AND2_X1 U7943 ( .A1(n8683), .A2(n8692), .ZN(n6311) );
  OR2_X1 U7944 ( .A1(n8683), .A2(n8692), .ZN(n6310) );
  INV_X1 U7945 ( .A(n8159), .ZN(n8264) );
  NAND2_X1 U7946 ( .A1(n8264), .A2(n8267), .ZN(n8361) );
  NAND2_X1 U7947 ( .A1(n8154), .A2(n8637), .ZN(n8647) );
  NAND2_X1 U7948 ( .A1(n8648), .A2(n8647), .ZN(n8646) );
  OAI21_X1 U7949 ( .B1(n9133), .B2(n8387), .A(n8646), .ZN(n8633) );
  INV_X1 U7950 ( .A(n8638), .ZN(n6312) );
  INV_X1 U7951 ( .A(n8623), .ZN(n8386) );
  NOR2_X1 U7952 ( .A1(n9119), .A2(n8386), .ZN(n6314) );
  INV_X1 U7953 ( .A(n9119), .ZN(n6313) );
  INV_X1 U7954 ( .A(n8083), .ZN(n8764) );
  NOR2_X1 U7955 ( .A1(n8129), .A2(n8568), .ZN(n6315) );
  INV_X1 U7956 ( .A(n8566), .ZN(n6316) );
  NAND2_X1 U7957 ( .A1(n9097), .A2(n8569), .ZN(n6318) );
  INV_X1 U7958 ( .A(n9097), .ZN(n6317) );
  AOI22_X1 U7959 ( .A1(n8555), .A2(n6318), .B1(n8028), .B2(n6317), .ZN(n6319)
         );
  XNOR2_X1 U7960 ( .A(n6319), .B(n8368), .ZN(n6337) );
  NAND2_X1 U7961 ( .A1(n6321), .A2(n6320), .ZN(n6322) );
  NAND2_X1 U7962 ( .A1(n6322), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7963 ( .A1(n8165), .A2(n6478), .ZN(n8336) );
  NAND2_X1 U7964 ( .A1(n8379), .A2(n8509), .ZN(n6479) );
  NAND2_X1 U7965 ( .A1(n8165), .A2(n8379), .ZN(n6332) );
  NAND2_X1 U7966 ( .A1(n8329), .A2(n8533), .ZN(n6894) );
  INV_X1 U7967 ( .A(n8379), .ZN(n8163) );
  AOI21_X1 U7968 ( .B1(n8163), .B2(n6478), .A(n8509), .ZN(n6324) );
  NAND2_X1 U7969 ( .A1(n8549), .A2(n7775), .ZN(n6335) );
  INV_X1 U7970 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n8747) );
  NAND2_X1 U7971 ( .A1(n4411), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7972 ( .A1(n6991), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6325) );
  OAI211_X1 U7973 ( .C1(n6994), .C2(n8747), .A(n6326), .B(n6325), .ZN(n6327)
         );
  INV_X1 U7974 ( .A(n6327), .ZN(n6328) );
  AND2_X1 U7975 ( .A1(n6997), .A2(n6328), .ZN(n8303) );
  INV_X1 U7976 ( .A(n8303), .ZN(n8383) );
  INV_X1 U7977 ( .A(n6331), .ZN(n6664) );
  INV_X2 U7978 ( .A(n6664), .ZN(n8376) );
  OAI21_X1 U7979 ( .B1(n6330), .B2(n8376), .A(n5946), .ZN(n6888) );
  NAND2_X1 U7980 ( .A1(n5946), .A2(P2_B_REG_SCAN_IN), .ZN(n6333) );
  AND2_X1 U7981 ( .A1(n8717), .A2(n6333), .ZN(n8537) );
  AOI22_X1 U7982 ( .A1(n8383), .A2(n8537), .B1(n8719), .B2(n8569), .ZN(n6334)
         );
  NAND2_X1 U7983 ( .A1(n6371), .A2(n6372), .ZN(n6339) );
  OR2_X1 U7984 ( .A1(n6341), .A2(n6340), .ZN(n6342) );
  NAND2_X1 U7985 ( .A1(n6341), .A2(n6340), .ZN(n6343) );
  XNOR2_X1 U7986 ( .A(n6347), .B(P2_B_REG_SCAN_IN), .ZN(n6346) );
  INV_X1 U7987 ( .A(n6369), .ZN(n7871) );
  INV_X1 U7988 ( .A(n6347), .ZN(n7711) );
  NAND2_X1 U7989 ( .A1(n7871), .A2(n7711), .ZN(n6590) );
  OAI21_X1 U7990 ( .B1(n6351), .B2(P2_D_REG_0__SCAN_IN), .A(n6590), .ZN(n6348)
         );
  INV_X1 U7991 ( .A(n6348), .ZN(n6893) );
  NAND3_X1 U7992 ( .A1(n6478), .A2(n8379), .A3(n8533), .ZN(n6350) );
  NAND2_X1 U7993 ( .A1(n6332), .A2(n6350), .ZN(n6354) );
  NAND2_X1 U7994 ( .A1(n6349), .A2(n6354), .ZN(n6357) );
  OR2_X1 U7995 ( .A1(n6351), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6353) );
  OR2_X1 U7996 ( .A1(n6352), .A2(n6369), .ZN(n6588) );
  INV_X1 U7997 ( .A(n6354), .ZN(n6355) );
  NAND2_X1 U7998 ( .A1(n6477), .A2(n6355), .ZN(n6356) );
  INV_X1 U7999 ( .A(n6477), .ZN(n6358) );
  NAND2_X1 U8000 ( .A1(n6348), .A2(n6358), .ZN(n6483) );
  NOR2_X1 U8001 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .ZN(
        n8985) );
  NOR4_X1 U8002 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6361) );
  NOR4_X1 U8003 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6360) );
  NOR4_X1 U8004 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6359) );
  AND4_X1 U8005 ( .A1(n8985), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n6367)
         );
  NOR4_X1 U8006 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n6365) );
  NOR4_X1 U8007 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6364) );
  NOR4_X1 U8008 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6363) );
  NOR4_X1 U8009 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6362) );
  AND4_X1 U8010 ( .A1(n6365), .A2(n6364), .A3(n6363), .A4(n6362), .ZN(n6366)
         );
  AND2_X1 U8011 ( .A1(n6367), .A2(n6366), .ZN(n6368) );
  INV_X1 U8012 ( .A(n6894), .ZN(n6373) );
  NOR2_X1 U8013 ( .A1(n6332), .A2(n6373), .ZN(n6864) );
  NOR2_X1 U8014 ( .A1(n6925), .A2(n6864), .ZN(n6374) );
  AND2_X1 U8015 ( .A1(n6481), .A2(n6374), .ZN(n6916) );
  NAND2_X1 U8016 ( .A1(n6488), .A2(n10384), .ZN(n6379) );
  INV_X1 U8017 ( .A(n10359), .ZN(n10325) );
  NAND2_X1 U8018 ( .A1(n6967), .A2(n6381), .ZN(n6968) );
  OR2_X1 U8019 ( .A1(n6380), .A2(n6977), .ZN(n6382) );
  NAND2_X1 U8020 ( .A1(n6968), .A2(n6382), .ZN(n6956) );
  XNOR2_X1 U8021 ( .A(n9645), .B(n6383), .ZN(n6958) );
  NAND2_X1 U8022 ( .A1(n6956), .A2(n6958), .ZN(n6955) );
  OR2_X1 U8023 ( .A1(n9645), .A2(n7140), .ZN(n6384) );
  NAND2_X1 U8024 ( .A1(n6955), .A2(n6384), .ZN(n6982) );
  NOR2_X1 U8025 ( .A1(n6385), .A2(n7365), .ZN(n9436) );
  NAND2_X1 U8026 ( .A1(n6385), .A2(n7365), .ZN(n9428) );
  NAND2_X1 U8027 ( .A1(n6982), .A2(n6983), .ZN(n6981) );
  INV_X1 U8028 ( .A(n6385), .ZN(n6827) );
  NAND2_X1 U8029 ( .A1(n6827), .A2(n7365), .ZN(n6386) );
  NAND2_X1 U8030 ( .A1(n6981), .A2(n6386), .ZN(n6946) );
  OR2_X1 U8031 ( .A1(n9644), .A2(n7331), .ZN(n9423) );
  NAND2_X1 U8032 ( .A1(n9644), .A2(n7331), .ZN(n9435) );
  NAND2_X1 U8033 ( .A1(n9423), .A2(n9435), .ZN(n9544) );
  INV_X1 U8034 ( .A(n9644), .ZN(n6387) );
  NAND2_X1 U8035 ( .A1(n6387), .A2(n7331), .ZN(n6388) );
  OR2_X1 U8036 ( .A1(n6389), .A2(n7153), .ZN(n9440) );
  NAND2_X1 U8037 ( .A1(n6389), .A2(n7153), .ZN(n9438) );
  INV_X1 U8038 ( .A(n9547), .ZN(n7066) );
  NAND2_X1 U8039 ( .A1(n7380), .A2(n7153), .ZN(n6390) );
  AND2_X1 U8040 ( .A1(n7336), .A2(n9642), .ZN(n9441) );
  NAND2_X1 U8041 ( .A1(n9334), .A2(n6391), .ZN(n9442) );
  INV_X1 U8042 ( .A(n9548), .ZN(n7265) );
  NAND2_X1 U8043 ( .A1(n7336), .A2(n6391), .ZN(n6392) );
  OR2_X1 U8044 ( .A1(n10204), .A2(n7280), .ZN(n9546) );
  NAND2_X1 U8045 ( .A1(n10204), .A2(n7280), .ZN(n7284) );
  NAND2_X1 U8046 ( .A1(n9546), .A2(n7284), .ZN(n9444) );
  OR2_X1 U8047 ( .A1(n10204), .A2(n9641), .ZN(n6393) );
  OR2_X1 U8048 ( .A1(n7502), .A2(n7452), .ZN(n9443) );
  NAND2_X1 U8049 ( .A1(n7502), .A2(n7452), .ZN(n9448) );
  NAND2_X1 U8050 ( .A1(n9443), .A2(n9448), .ZN(n7283) );
  INV_X1 U8051 ( .A(n7452), .ZN(n9640) );
  NAND2_X1 U8052 ( .A1(n7459), .A2(n7344), .ZN(n9458) );
  NAND2_X1 U8053 ( .A1(n9455), .A2(n9458), .ZN(n7451) );
  NAND2_X1 U8054 ( .A1(n7448), .A2(n7451), .ZN(n7447) );
  INV_X1 U8055 ( .A(n7344), .ZN(n9639) );
  OR2_X1 U8056 ( .A1(n7459), .A2(n9639), .ZN(n6394) );
  NAND2_X1 U8057 ( .A1(n7447), .A2(n6394), .ZN(n7350) );
  OR2_X1 U8058 ( .A1(n7426), .A2(n7665), .ZN(n9461) );
  NAND2_X1 U8059 ( .A1(n7426), .A2(n7665), .ZN(n9457) );
  NAND2_X1 U8060 ( .A1(n9461), .A2(n9457), .ZN(n9551) );
  NAND2_X1 U8061 ( .A1(n7350), .A2(n9551), .ZN(n7349) );
  OR2_X1 U8062 ( .A1(n7426), .A2(n9638), .ZN(n6395) );
  NAND2_X1 U8063 ( .A1(n7349), .A2(n6395), .ZN(n7660) );
  NAND2_X1 U8064 ( .A1(n10187), .A2(n7506), .ZN(n9464) );
  NAND2_X1 U8065 ( .A1(n9460), .A2(n9464), .ZN(n9555) );
  NAND2_X1 U8066 ( .A1(n7660), .A2(n9555), .ZN(n7659) );
  INV_X1 U8067 ( .A(n7506), .ZN(n9637) );
  OR2_X1 U8068 ( .A1(n10187), .A2(n9637), .ZN(n6396) );
  NAND2_X1 U8069 ( .A1(n7659), .A2(n6396), .ZN(n7513) );
  OR2_X1 U8070 ( .A1(n9229), .A2(n7666), .ZN(n9466) );
  NAND2_X1 U8071 ( .A1(n9229), .A2(n7666), .ZN(n9463) );
  NAND2_X1 U8072 ( .A1(n7513), .A2(n7512), .ZN(n7511) );
  OR2_X1 U8073 ( .A1(n9229), .A2(n9636), .ZN(n6397) );
  NAND2_X1 U8074 ( .A1(n7511), .A2(n6397), .ZN(n7637) );
  INV_X1 U8075 ( .A(n9294), .ZN(n7639) );
  INV_X1 U8076 ( .A(n7703), .ZN(n9635) );
  NAND2_X1 U8077 ( .A1(n9294), .A2(n7703), .ZN(n9487) );
  NAND2_X1 U8078 ( .A1(n7637), .A2(n7636), .ZN(n7635) );
  OR2_X1 U8079 ( .A1(n9294), .A2(n9635), .ZN(n6398) );
  NAND2_X1 U8080 ( .A1(n7635), .A2(n6398), .ZN(n7696) );
  INV_X1 U8081 ( .A(n7795), .ZN(n9634) );
  NOR2_X1 U8082 ( .A1(n10015), .A2(n9634), .ZN(n6400) );
  NAND2_X1 U8083 ( .A1(n10015), .A2(n9634), .ZN(n6399) );
  INV_X1 U8084 ( .A(n7853), .ZN(n9633) );
  AND2_X1 U8085 ( .A1(n9352), .A2(n9633), .ZN(n6401) );
  OR2_X1 U8086 ( .A1(n9352), .A2(n9633), .ZN(n6402) );
  NAND2_X1 U8087 ( .A1(n10011), .A2(n9258), .ZN(n9492) );
  OR2_X1 U8088 ( .A1(n10003), .A2(n9631), .ZN(n6403) );
  NAND2_X1 U8089 ( .A1(n10003), .A2(n9631), .ZN(n6404) );
  OR2_X1 U8090 ( .A1(n9911), .A2(n9630), .ZN(n6405) );
  NAND2_X1 U8091 ( .A1(n9892), .A2(n9280), .ZN(n6407) );
  NAND2_X1 U8092 ( .A1(n9878), .A2(n9628), .ZN(n6408) );
  AND2_X1 U8093 ( .A1(n9861), .A2(n9627), .ZN(n6409) );
  OR2_X1 U8094 ( .A1(n9861), .A2(n9627), .ZN(n6410) );
  INV_X1 U8095 ( .A(n9235), .ZN(n9624) );
  NAND2_X1 U8096 ( .A1(n9810), .A2(n9624), .ZN(n6411) );
  AND2_X1 U8097 ( .A1(n9792), .A2(n9623), .ZN(n6412) );
  NAND2_X1 U8098 ( .A1(n9759), .A2(n6413), .ZN(n9526) );
  NAND2_X1 U8099 ( .A1(n9528), .A2(n9526), .ZN(n9571) );
  OR2_X1 U8100 ( .A1(n9759), .A2(n9621), .ZN(n6414) );
  NAND2_X1 U8101 ( .A1(n9742), .A2(n6471), .ZN(n9522) );
  NAND2_X1 U8102 ( .A1(n4494), .A2(n9522), .ZN(n9574) );
  NOR2_X1 U8103 ( .A1(n9739), .A2(n9738), .ZN(n9741) );
  AOI21_X1 U8104 ( .B1(n9742), .B2(n9620), .A(n9741), .ZN(n6420) );
  NAND2_X1 U8105 ( .A1(n5610), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n6417) );
  NAND2_X1 U8106 ( .A1(n6452), .A2(n6885), .ZN(n9588) );
  INV_X1 U8107 ( .A(n9576), .ZN(n6419) );
  XNOR2_X1 U8108 ( .A(n6420), .B(n6419), .ZN(n9725) );
  INV_X1 U8109 ( .A(n6456), .ZN(n7002) );
  OAI21_X1 U8110 ( .B1(n9613), .B2(n6421), .A(n7002), .ZN(n7098) );
  AND2_X1 U8111 ( .A1(n9613), .A2(n9608), .ZN(n6422) );
  OR2_X1 U8112 ( .A1(n7098), .A2(n6422), .ZN(n7290) );
  OR2_X1 U8113 ( .A1(n9792), .A2(n9269), .ZN(n9519) );
  NAND2_X1 U8114 ( .A1(n9792), .A2(n9269), .ZN(n9517) );
  NAND2_X1 U8115 ( .A1(n9519), .A2(n9517), .ZN(n9570) );
  INV_X1 U8116 ( .A(n9570), .ZN(n9789) );
  OR2_X1 U8117 ( .A1(n9810), .A2(n9235), .ZN(n9784) );
  NOR2_X1 U8118 ( .A1(n9647), .A2(n7104), .ZN(n6999) );
  INV_X1 U8119 ( .A(n6380), .ZN(n6826) );
  NAND2_X1 U8120 ( .A1(n6826), .A2(n6977), .ZN(n6957) );
  NAND2_X1 U8121 ( .A1(n6971), .A2(n6957), .ZN(n6424) );
  NAND2_X1 U8122 ( .A1(n6424), .A2(n9541), .ZN(n6960) );
  INV_X1 U8123 ( .A(n9645), .ZN(n6835) );
  NAND2_X1 U8124 ( .A1(n6835), .A2(n7140), .ZN(n6425) );
  INV_X1 U8125 ( .A(n9435), .ZN(n6426) );
  AND2_X1 U8126 ( .A1(n9438), .A2(n9423), .ZN(n9429) );
  NAND2_X1 U8127 ( .A1(n6427), .A2(n9440), .ZN(n7264) );
  AND2_X1 U8128 ( .A1(n9448), .A2(n7284), .ZN(n9432) );
  NAND2_X1 U8129 ( .A1(n6428), .A2(n9458), .ZN(n9553) );
  INV_X1 U8130 ( .A(n9553), .ZN(n6429) );
  NAND2_X1 U8131 ( .A1(n9546), .A2(n4797), .ZN(n6430) );
  NOR2_X1 U8132 ( .A1(n9552), .A2(n6430), .ZN(n6431) );
  OR2_X1 U8133 ( .A1(n9553), .A2(n6431), .ZN(n9388) );
  INV_X1 U8134 ( .A(n9555), .ZN(n6432) );
  INV_X1 U8135 ( .A(n9460), .ZN(n6433) );
  NOR2_X1 U8136 ( .A1(n7512), .A2(n6433), .ZN(n6434) );
  NAND2_X1 U8137 ( .A1(n7630), .A2(n9396), .ZN(n7701) );
  NAND2_X1 U8138 ( .A1(n7701), .A2(n9487), .ZN(n6435) );
  OR2_X1 U8139 ( .A1(n10015), .A2(n7795), .ZN(n9489) );
  NAND2_X1 U8140 ( .A1(n10015), .A2(n7795), .ZN(n9486) );
  NAND2_X1 U8141 ( .A1(n9489), .A2(n9486), .ZN(n9469) );
  NAND2_X1 U8142 ( .A1(n6435), .A2(n9559), .ZN(n7793) );
  AND2_X1 U8143 ( .A1(n7845), .A2(n9633), .ZN(n9473) );
  INV_X1 U8144 ( .A(n9473), .ZN(n9382) );
  NAND2_X1 U8145 ( .A1(n9352), .A2(n7853), .ZN(n9494) );
  NAND2_X1 U8146 ( .A1(n9382), .A2(n9494), .ZN(n9561) );
  INV_X1 U8147 ( .A(n9486), .ZN(n6436) );
  NOR2_X1 U8148 ( .A1(n9561), .A2(n6436), .ZN(n6437) );
  NAND2_X1 U8149 ( .A1(n7793), .A2(n6437), .ZN(n6438) );
  NAND2_X1 U8150 ( .A1(n6438), .A2(n9382), .ZN(n7852) );
  NAND2_X1 U8151 ( .A1(n10003), .A2(n7854), .ZN(n9478) );
  NAND2_X1 U8152 ( .A1(n9911), .A2(n9259), .ZN(n9481) );
  NAND2_X1 U8153 ( .A1(n9905), .A2(n9904), .ZN(n6439) );
  NAND2_X1 U8154 ( .A1(n9992), .A2(n9280), .ZN(n9475) );
  NAND2_X1 U8155 ( .A1(n9496), .A2(n9475), .ZN(n9894) );
  XNOR2_X1 U8156 ( .A(n9878), .B(n9628), .ZN(n9875) );
  INV_X1 U8157 ( .A(n9416), .ZN(n6440) );
  XNOR2_X1 U8158 ( .A(n9861), .B(n9627), .ZN(n9856) );
  NAND2_X1 U8159 ( .A1(n9861), .A2(n9370), .ZN(n9503) );
  OR2_X1 U8160 ( .A1(n9842), .A2(n9217), .ZN(n9365) );
  NAND2_X1 U8161 ( .A1(n9842), .A2(n9217), .ZN(n9372) );
  NAND2_X1 U8162 ( .A1(n9835), .A2(n9840), .ZN(n6441) );
  NAND2_X1 U8163 ( .A1(n6441), .A2(n9372), .ZN(n9818) );
  OR2_X1 U8164 ( .A1(n9827), .A2(n9512), .ZN(n9366) );
  NAND2_X1 U8165 ( .A1(n9366), .A2(n9801), .ZN(n9568) );
  NAND2_X1 U8166 ( .A1(n9818), .A2(n9823), .ZN(n9817) );
  NAND2_X1 U8167 ( .A1(n9810), .A2(n9235), .ZN(n9514) );
  OR2_X1 U8168 ( .A1(n9781), .A2(n9236), .ZN(n9520) );
  NAND2_X1 U8169 ( .A1(n9520), .A2(n9518), .ZN(n9771) );
  INV_X1 U8170 ( .A(n9771), .ZN(n9768) );
  NAND2_X1 U8171 ( .A1(n6442), .A2(n9522), .ZN(n6443) );
  XNOR2_X1 U8172 ( .A(n9576), .B(n6443), .ZN(n6451) );
  NAND2_X1 U8173 ( .A1(n9601), .A2(n6444), .ZN(n6445) );
  OAI21_X2 U8174 ( .B1(n5850), .B2(n7300), .A(n6445), .ZN(n9931) );
  INV_X1 U8175 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9942) );
  NOR2_X1 U8176 ( .A1(n5251), .A2(n9942), .ZN(n6448) );
  INV_X1 U8177 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8773) );
  NOR2_X1 U8178 ( .A1(n9364), .A2(n8773), .ZN(n6447) );
  INV_X1 U8179 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10026) );
  NOR2_X1 U8180 ( .A1(n5170), .A2(n10026), .ZN(n6446) );
  OR3_X1 U8181 ( .A1(n6448), .A2(n6447), .A3(n6446), .ZN(n9619) );
  INV_X1 U8182 ( .A(n9619), .ZN(n9412) );
  INV_X1 U8183 ( .A(P1_B_REG_SCAN_IN), .ZN(n8805) );
  OR2_X1 U8184 ( .A1(n6554), .A2(n8805), .ZN(n6449) );
  NAND2_X1 U8185 ( .A1(n9321), .A2(n6449), .ZN(n9711) );
  OAI22_X1 U8186 ( .A1(n6471), .A2(n9300), .B1(n9412), .B2(n9711), .ZN(n6450)
         );
  INV_X1 U8187 ( .A(n7331), .ZN(n6947) );
  AND2_X1 U8188 ( .A1(n7455), .A2(n10213), .ZN(n7351) );
  INV_X1 U8189 ( .A(n10187), .ZN(n6454) );
  INV_X1 U8190 ( .A(n10015), .ZN(n7700) );
  NAND2_X1 U8191 ( .A1(n7845), .A2(n7800), .ZN(n7859) );
  NOR2_X2 U8192 ( .A1(n9792), .A2(n9808), .ZN(n9791) );
  OAI211_X1 U8193 ( .C1(n6491), .C2(n4439), .A(n9777), .B(n9719), .ZN(n9729)
         );
  OR2_X1 U8194 ( .A1(n9614), .A2(n6459), .ZN(n6461) );
  INV_X1 U8195 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6463) );
  OR2_X1 U8196 ( .A1(n10220), .A2(n6463), .ZN(n6464) );
  OAI21_X1 U8197 ( .B1(n6497), .B2(n10218), .A(n5028), .ZN(P1_U3519) );
  INV_X1 U8198 ( .A(n6465), .ZN(n6468) );
  INV_X1 U8199 ( .A(n6470), .ZN(n9760) );
  AOI22_X1 U8200 ( .A1(n9760), .A2(n9337), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6475) );
  OR2_X1 U8201 ( .A1(n6471), .A2(n9301), .ZN(n6473) );
  INV_X1 U8202 ( .A(n9300), .ZN(n9320) );
  NAND2_X1 U8203 ( .A1(n9622), .A2(n9320), .ZN(n6472) );
  NAND2_X1 U8204 ( .A1(n6473), .A2(n6472), .ZN(n9752) );
  NAND2_X1 U8205 ( .A1(n9752), .A2(n9346), .ZN(n6474) );
  OAI211_X1 U8206 ( .C1(n10035), .C2(n9283), .A(n6475), .B(n6474), .ZN(n6476)
         );
  AND2_X1 U8207 ( .A1(n6349), .A2(n6477), .ZN(n6918) );
  NAND2_X1 U8208 ( .A1(n6918), .A2(n6481), .ZN(n6879) );
  NOR2_X1 U8209 ( .A1(n6879), .A2(n6925), .ZN(n6860) );
  INV_X1 U8210 ( .A(n8165), .ZN(n7603) );
  NAND2_X1 U8211 ( .A1(n7603), .A2(n6478), .ZN(n8340) );
  OR2_X1 U8212 ( .A1(n8340), .A2(n6479), .ZN(n6861) );
  NAND2_X1 U8213 ( .A1(n6887), .A2(n6861), .ZN(n6480) );
  NAND2_X1 U8214 ( .A1(n6860), .A2(n6480), .ZN(n6486) );
  INV_X1 U8215 ( .A(n6481), .ZN(n6482) );
  AND2_X1 U8216 ( .A1(n10359), .A2(n8312), .ZN(n6484) );
  NAND2_X1 U8217 ( .A1(n6484), .A2(n6861), .ZN(n6858) );
  INV_X1 U8218 ( .A(n6878), .ZN(n7125) );
  NAND2_X1 U8219 ( .A1(n6858), .A2(n8731), .ZN(n6869) );
  NAND2_X1 U8220 ( .A1(n6890), .A2(n6869), .ZN(n6485) );
  OR2_X1 U8221 ( .A1(n10367), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6487) );
  INV_X1 U8222 ( .A(n10223), .ZN(n6496) );
  INV_X1 U8223 ( .A(n6498), .ZN(n6499) );
  INV_X1 U8224 ( .A(n6875), .ZN(n6501) );
  NAND2_X1 U8225 ( .A1(n6866), .A2(n6332), .ZN(n6502) );
  NAND2_X1 U8226 ( .A1(n6502), .A2(n6658), .ZN(n6663) );
  NAND2_X1 U8227 ( .A1(n6663), .A2(n5946), .ZN(n6503) );
  NAND2_X1 U8228 ( .A1(n6503), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NAND2_X2 U8229 ( .A1(n5212), .A2(P2_U3151), .ZN(n9169) );
  INV_X1 U8230 ( .A(n9166), .ZN(n9171) );
  OAI222_X1 U8231 ( .A1(n9169), .A2(n6511), .B1(n9171), .B2(n5931), .C1(
        P2_U3151), .C2(n6689), .ZN(P2_U3294) );
  INV_X1 U8232 ( .A(n6504), .ZN(n6518) );
  INV_X1 U8233 ( .A(n6754), .ZN(n6721) );
  INV_X1 U8234 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6505) );
  OAI222_X1 U8235 ( .A1(n9169), .A2(n6518), .B1(n6721), .B2(P2_U3151), .C1(
        n6505), .C2(n9171), .ZN(P2_U3292) );
  OAI222_X1 U8236 ( .A1(n9169), .A2(n6509), .B1(n5959), .B2(P2_U3151), .C1(
        n4551), .C2(n9171), .ZN(P2_U3293) );
  NAND2_X1 U8237 ( .A1(n4525), .A2(P1_U3086), .ZN(n7911) );
  INV_X1 U8238 ( .A(n6506), .ZN(n6523) );
  INV_X1 U8239 ( .A(n10082), .ZN(n7682) );
  OAI222_X1 U8240 ( .A1(n6679), .A2(P1_U3086), .B1(n7911), .B2(n6523), .C1(
        n6507), .C2(n7682), .ZN(P1_U3348) );
  INV_X1 U8241 ( .A(n7911), .ZN(n7656) );
  AOI22_X1 U8242 ( .A1(n10082), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n6740), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6508) );
  OAI21_X1 U8243 ( .B1(n6509), .B2(n10085), .A(n6508), .ZN(P1_U3353) );
  AOI22_X1 U8244 ( .A1(n10082), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        P1_STATE_REG_SCAN_IN), .B2(n6574), .ZN(n6510) );
  OAI21_X1 U8245 ( .B1(n6511), .B2(n10085), .A(n6510), .ZN(P1_U3354) );
  OAI222_X1 U8246 ( .A1(n6649), .A2(P1_U3086), .B1(n10085), .B2(n6525), .C1(
        n6512), .C2(n7682), .ZN(P1_U3349) );
  INV_X1 U8247 ( .A(n6513), .ZN(n6521) );
  OAI222_X1 U8248 ( .A1(n6616), .A2(P1_U3086), .B1(n10085), .B2(n6521), .C1(
        n6514), .C2(n7682), .ZN(P1_U3350) );
  INV_X1 U8249 ( .A(n6515), .ZN(n6519) );
  OAI222_X1 U8250 ( .A1(n9659), .A2(P1_U3086), .B1(n10085), .B2(n6519), .C1(
        n6516), .C2(n7682), .ZN(P1_U3351) );
  INV_X1 U8251 ( .A(n6604), .ZN(n6595) );
  INV_X1 U8252 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6517) );
  OAI222_X1 U8253 ( .A1(P1_U3086), .A2(n6595), .B1(n10085), .B2(n6518), .C1(
        n6517), .C2(n7682), .ZN(P1_U3352) );
  INV_X1 U8254 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6520) );
  OAI222_X1 U8255 ( .A1(n9171), .A2(n6520), .B1(n9169), .B2(n6519), .C1(
        P2_U3151), .C2(n6790), .ZN(P2_U3291) );
  INV_X1 U8256 ( .A(n6799), .ZN(n7047) );
  OAI222_X1 U8257 ( .A1(n9171), .A2(n6522), .B1(n9169), .B2(n6521), .C1(
        P2_U3151), .C2(n7047), .ZN(P2_U3290) );
  OAI222_X1 U8258 ( .A1(n9171), .A2(n6524), .B1(n9169), .B2(n6523), .C1(
        P2_U3151), .C2(n7038), .ZN(P2_U3288) );
  OAI222_X1 U8259 ( .A1(n9171), .A2(n6526), .B1(n9169), .B2(n6525), .C1(
        P2_U3151), .C2(n7052), .ZN(P2_U3289) );
  INV_X1 U8260 ( .A(n6527), .ZN(n6529) );
  OAI222_X1 U8261 ( .A1(n9677), .A2(P1_U3086), .B1(n10085), .B2(n6529), .C1(
        n6528), .C2(n7682), .ZN(P1_U3347) );
  INV_X1 U8262 ( .A(n7193), .ZN(n7056) );
  OAI222_X1 U8263 ( .A1(n9171), .A2(n6530), .B1(n9169), .B2(n6529), .C1(
        P2_U3151), .C2(n7056), .ZN(P2_U3287) );
  INV_X1 U8264 ( .A(n6531), .ZN(n6543) );
  OAI222_X1 U8265 ( .A1(n9169), .A2(n6543), .B1(n7313), .B2(P2_U3151), .C1(
        n6532), .C2(n9171), .ZN(P2_U3286) );
  NAND2_X1 U8266 ( .A1(n9614), .A2(n9617), .ZN(n6537) );
  NAND2_X1 U8267 ( .A1(n9595), .A2(n6533), .ZN(n6534) );
  INV_X1 U8268 ( .A(n6536), .ZN(n6535) );
  INV_X1 U8269 ( .A(n10155), .ZN(n10171) );
  INV_X1 U8270 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6541) );
  INV_X1 U8271 ( .A(n6554), .ZN(n9610) );
  INV_X1 U8272 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7100) );
  AOI21_X1 U8273 ( .B1(n9610), .B2(n7100), .A(n5856), .ZN(n6739) );
  OAI21_X1 U8274 ( .B1(n9610), .B2(P1_REG1_REG_0__SCAN_IN), .A(n6739), .ZN(
        n6538) );
  XNOR2_X1 U8275 ( .A(n6538), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6539) );
  AOI22_X1 U8276 ( .A1(n6556), .A2(n6539), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6540) );
  OAI21_X1 U8277 ( .B1(n10171), .B2(n6541), .A(n6540), .ZN(P1_U3243) );
  OAI222_X1 U8278 ( .A1(P1_U3086), .A2(n10111), .B1(n10085), .B2(n6543), .C1(
        n6542), .C2(n7682), .ZN(P1_U3346) );
  NOR2_X1 U8279 ( .A1(n10155), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8280 ( .A(n6925), .ZN(n6544) );
  INV_X1 U8281 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n8880) );
  NOR2_X1 U8282 ( .A1(n6587), .A2(n8880), .ZN(P2_U3238) );
  INV_X1 U8283 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n8819) );
  NOR2_X1 U8284 ( .A1(n6587), .A2(n8819), .ZN(P2_U3241) );
  INV_X1 U8285 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n8936) );
  NOR2_X1 U8286 ( .A1(n6587), .A2(n8936), .ZN(P2_U3255) );
  INV_X1 U8287 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n8821) );
  NOR2_X1 U8288 ( .A1(n6587), .A2(n8821), .ZN(P2_U3244) );
  NAND2_X1 U8289 ( .A1(n6380), .A2(P1_U3973), .ZN(n6545) );
  OAI21_X1 U8290 ( .B1(P1_U3973), .B2(n5931), .A(n6545), .ZN(P1_U3555) );
  INV_X1 U8291 ( .A(n6546), .ZN(n6549) );
  INV_X1 U8292 ( .A(n7551), .ZN(n7555) );
  INV_X1 U8293 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6547) );
  OAI222_X1 U8294 ( .A1(n9169), .A2(n6549), .B1(n7555), .B2(P2_U3151), .C1(
        n6547), .C2(n9171), .ZN(P2_U3285) );
  OAI222_X1 U8295 ( .A1(P1_U3086), .A2(n6807), .B1(n10085), .B2(n6549), .C1(
        n6548), .C2(n7682), .ZN(P1_U3345) );
  INV_X1 U8296 ( .A(n6556), .ZN(n6550) );
  INV_X1 U8297 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6978) );
  XNOR2_X1 U8298 ( .A(n6574), .B(n6978), .ZN(n6573) );
  AND2_X1 U8299 ( .A1(P1_REG1_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6572) );
  XNOR2_X1 U8300 ( .A(n6573), .B(n6572), .ZN(n6560) );
  INV_X1 U8301 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6551) );
  INV_X1 U8302 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6841) );
  OAI22_X1 U8303 ( .A1(n10171), .A2(n6551), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6841), .ZN(n6552) );
  AOI21_X1 U8304 ( .B1(n6574), .B2(n10173), .A(n6552), .ZN(n6559) );
  AND2_X1 U8305 ( .A1(P1_REG2_REG_0__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6736) );
  INV_X1 U8306 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6553) );
  MUX2_X1 U8307 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6553), .S(n6574), .Z(n6557)
         );
  NOR2_X1 U8308 ( .A1(n5856), .A2(n6554), .ZN(n6555) );
  NAND2_X1 U8309 ( .A1(n6574), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6567) );
  OAI211_X1 U8310 ( .C1(n6574), .C2(P1_REG2_REG_1__SCAN_IN), .A(n6736), .B(
        n6567), .ZN(n6568) );
  OAI211_X1 U8311 ( .C1(n6736), .C2(n6557), .A(n10158), .B(n6568), .ZN(n6558)
         );
  OAI211_X1 U8312 ( .C1(n9701), .C2(n6560), .A(n6559), .B(n6558), .ZN(P1_U3244) );
  INV_X1 U8313 ( .A(n6561), .ZN(n6564) );
  OAI222_X1 U8314 ( .A1(n9171), .A2(n6562), .B1(n9169), .B2(n6564), .C1(
        P2_U3151), .C2(n7830), .ZN(P2_U3284) );
  OAI222_X1 U8315 ( .A1(n10118), .A2(P1_U3086), .B1(n7911), .B2(n6564), .C1(
        n6563), .C2(n7682), .ZN(P1_U3344) );
  AND2_X1 U8316 ( .A1(n6565), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8317 ( .A1(n6565), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8318 ( .A1(n6565), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8319 ( .A1(n6565), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8320 ( .A1(n6565), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8321 ( .A1(n6565), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8322 ( .A1(n6565), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8323 ( .A1(n6565), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8324 ( .A1(n6565), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8325 ( .A1(n6565), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8326 ( .A1(n6565), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  INV_X1 U8327 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6566) );
  XNOR2_X1 U8328 ( .A(n6740), .B(n6566), .ZN(n6743) );
  NAND2_X1 U8329 ( .A1(n6568), .A2(n6567), .ZN(n6741) );
  AOI22_X1 U8330 ( .A1(n6743), .A2(n6741), .B1(n6740), .B2(
        P1_REG2_REG_2__SCAN_IN), .ZN(n6570) );
  MUX2_X1 U8331 ( .A(n6594), .B(P1_REG2_REG_3__SCAN_IN), .S(n6604), .Z(n6569)
         );
  NOR2_X1 U8332 ( .A1(n6570), .A2(n6569), .ZN(n9658) );
  AOI211_X1 U8333 ( .C1(n6570), .C2(n6569), .A(n9658), .B(n10182), .ZN(n6584)
         );
  MUX2_X1 U8334 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6571), .S(n6740), .Z(n6747)
         );
  NAND2_X1 U8335 ( .A1(n6573), .A2(n6572), .ZN(n6576) );
  NAND2_X1 U8336 ( .A1(n6574), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6575) );
  NAND2_X1 U8337 ( .A1(n6576), .A2(n6575), .ZN(n6746) );
  NAND2_X1 U8338 ( .A1(n6747), .A2(n6746), .ZN(n6745) );
  NAND2_X1 U8339 ( .A1(n6740), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6580) );
  NAND2_X1 U8340 ( .A1(n6745), .A2(n6580), .ZN(n6579) );
  MUX2_X1 U8341 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6577), .S(n6604), .Z(n6578)
         );
  NAND2_X1 U8342 ( .A1(n6579), .A2(n6578), .ZN(n9662) );
  MUX2_X1 U8343 ( .A(n6577), .B(P1_REG1_REG_3__SCAN_IN), .S(n6604), .Z(n6581)
         );
  NAND3_X1 U8344 ( .A1(n6581), .A2(n6745), .A3(n6580), .ZN(n6582) );
  AND3_X1 U8345 ( .A1(n10175), .A2(n9662), .A3(n6582), .ZN(n6583) );
  NOR2_X1 U8346 ( .A1(n6584), .A2(n6583), .ZN(n6586) );
  AND2_X1 U8347 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6852) );
  AOI21_X1 U8348 ( .B1(n10155), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6852), .ZN(
        n6585) );
  OAI211_X1 U8349 ( .C1(n6595), .C2(n9674), .A(n6586), .B(n6585), .ZN(P1_U3246) );
  INV_X1 U8350 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n8916) );
  INV_X1 U8351 ( .A(n6588), .ZN(n6589) );
  AOI22_X1 U8352 ( .A1(n6565), .A2(n8916), .B1(n6875), .B2(n6589), .ZN(
        P2_U3377) );
  INV_X1 U8353 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n8978) );
  INV_X1 U8354 ( .A(n6590), .ZN(n6591) );
  AOI22_X1 U8355 ( .A1(n6565), .A2(n8978), .B1(n6875), .B2(n6591), .ZN(
        P2_U3376) );
  INV_X1 U8356 ( .A(n6592), .ZN(n6651) );
  INV_X1 U8357 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6593) );
  OAI222_X1 U8358 ( .A1(n9169), .A2(n6651), .B1(n8414), .B2(P2_U3151), .C1(
        n6593), .C2(n9171), .ZN(P2_U3283) );
  NAND2_X1 U8359 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7182) );
  INV_X1 U8360 ( .A(n9659), .ZN(n9648) );
  NOR2_X1 U8361 ( .A1(n6595), .A2(n6594), .ZN(n9653) );
  MUX2_X1 U8362 ( .A(n6596), .B(P1_REG2_REG_4__SCAN_IN), .S(n9659), .Z(n6597)
         );
  OAI21_X1 U8363 ( .B1(n9658), .B2(n9653), .A(n6597), .ZN(n9656) );
  INV_X1 U8364 ( .A(n9656), .ZN(n6598) );
  AOI21_X1 U8365 ( .B1(n9648), .B2(P1_REG2_REG_4__SCAN_IN), .A(n6598), .ZN(
        n6600) );
  MUX2_X1 U8366 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7083), .S(n6616), .Z(n6599)
         );
  NOR2_X1 U8367 ( .A1(n6600), .A2(n6599), .ZN(n6617) );
  AOI211_X1 U8368 ( .C1(n6600), .C2(n6599), .A(n6617), .B(n10182), .ZN(n6601)
         );
  INV_X1 U8369 ( .A(n6601), .ZN(n6602) );
  NAND2_X1 U8370 ( .A1(n7182), .A2(n6602), .ZN(n6603) );
  AOI21_X1 U8371 ( .B1(n10155), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n6603), .ZN(
        n6615) );
  NAND2_X1 U8372 ( .A1(n6604), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9661) );
  NAND2_X1 U8373 ( .A1(n9662), .A2(n9661), .ZN(n6607) );
  MUX2_X1 U8374 ( .A(n6605), .B(P1_REG1_REG_4__SCAN_IN), .S(n9659), .Z(n6606)
         );
  NAND2_X1 U8375 ( .A1(n6607), .A2(n6606), .ZN(n9664) );
  NAND2_X1 U8376 ( .A1(n9648), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U8377 ( .A1(n9664), .A2(n6612), .ZN(n6610) );
  INV_X1 U8378 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6608) );
  MUX2_X1 U8379 ( .A(n6608), .B(P1_REG1_REG_5__SCAN_IN), .S(n6616), .Z(n6609)
         );
  NAND2_X1 U8380 ( .A1(n6610), .A2(n6609), .ZN(n6644) );
  MUX2_X1 U8381 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6608), .S(n6616), .Z(n6611)
         );
  NAND3_X1 U8382 ( .A1(n9664), .A2(n6612), .A3(n6611), .ZN(n6613) );
  NAND3_X1 U8383 ( .A1(n10175), .A2(n6644), .A3(n6613), .ZN(n6614) );
  OAI211_X1 U8384 ( .C1(n9674), .C2(n6616), .A(n6615), .B(n6614), .ZN(P1_U3248) );
  NAND2_X1 U8385 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n7442) );
  INV_X1 U8386 ( .A(n6649), .ZN(n6618) );
  INV_X1 U8387 ( .A(n6616), .ZN(n6624) );
  AOI21_X1 U8388 ( .B1(n6624), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6617), .ZN(
        n6638) );
  MUX2_X1 U8389 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7163), .S(n6649), .Z(n6637)
         );
  NOR2_X1 U8390 ( .A1(n6638), .A2(n6637), .ZN(n6636) );
  AOI21_X1 U8391 ( .B1(P1_REG2_REG_6__SCAN_IN), .B2(n6618), .A(n6636), .ZN(
        n6620) );
  MUX2_X1 U8392 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n7272), .S(n6679), .Z(n6619)
         );
  NOR2_X1 U8393 ( .A1(n6620), .A2(n6619), .ZN(n9671) );
  AOI211_X1 U8394 ( .C1(n6620), .C2(n6619), .A(n9671), .B(n10182), .ZN(n6621)
         );
  INV_X1 U8395 ( .A(n6621), .ZN(n6622) );
  NAND2_X1 U8396 ( .A1(n7442), .A2(n6622), .ZN(n6623) );
  AOI21_X1 U8397 ( .B1(n10155), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n6623), .ZN(
        n6635) );
  NAND2_X1 U8398 ( .A1(n6624), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6643) );
  NAND2_X1 U8399 ( .A1(n6644), .A2(n6643), .ZN(n6626) );
  MUX2_X1 U8400 ( .A(n6627), .B(P1_REG1_REG_6__SCAN_IN), .S(n6649), .Z(n6625)
         );
  NAND2_X1 U8401 ( .A1(n6626), .A2(n6625), .ZN(n6646) );
  OR2_X1 U8402 ( .A1(n6649), .A2(n6627), .ZN(n6632) );
  NAND2_X1 U8403 ( .A1(n6646), .A2(n6632), .ZN(n6630) );
  INV_X1 U8404 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6628) );
  MUX2_X1 U8405 ( .A(n6628), .B(P1_REG1_REG_7__SCAN_IN), .S(n6679), .Z(n6629)
         );
  NAND2_X1 U8406 ( .A1(n6630), .A2(n6629), .ZN(n9680) );
  MUX2_X1 U8407 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n6628), .S(n6679), .Z(n6631)
         );
  NAND3_X1 U8408 ( .A1(n6646), .A2(n6632), .A3(n6631), .ZN(n6633) );
  NAND3_X1 U8409 ( .A1(n10175), .A2(n9680), .A3(n6633), .ZN(n6634) );
  OAI211_X1 U8410 ( .C1(n9674), .C2(n6679), .A(n6635), .B(n6634), .ZN(P1_U3250) );
  NAND2_X1 U8411 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9331) );
  AOI211_X1 U8412 ( .C1(n6638), .C2(n6637), .A(n6636), .B(n10182), .ZN(n6639)
         );
  INV_X1 U8413 ( .A(n6639), .ZN(n6640) );
  NAND2_X1 U8414 ( .A1(n9331), .A2(n6640), .ZN(n6641) );
  AOI21_X1 U8415 ( .B1(n10155), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n6641), .ZN(
        n6648) );
  MUX2_X1 U8416 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6627), .S(n6649), .Z(n6642)
         );
  NAND3_X1 U8417 ( .A1(n6644), .A2(n6643), .A3(n6642), .ZN(n6645) );
  NAND3_X1 U8418 ( .A1(n10175), .A2(n6646), .A3(n6645), .ZN(n6647) );
  OAI211_X1 U8419 ( .C1(n9674), .C2(n6649), .A(n6648), .B(n6647), .ZN(P1_U3249) );
  OAI222_X1 U8420 ( .A1(P1_U3086), .A2(n6809), .B1(n7911), .B2(n6651), .C1(
        n6650), .C2(n7682), .ZN(P1_U3343) );
  AND2_X1 U8421 ( .A1(n6565), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8422 ( .A1(n6565), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8423 ( .A1(n6565), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8424 ( .A1(n6565), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U8425 ( .A1(n6565), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8426 ( .A1(n6565), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8427 ( .A1(n6565), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8428 ( .A1(n6565), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8429 ( .A1(n6565), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8430 ( .A1(n6565), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8431 ( .A1(n6565), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8432 ( .A1(n6565), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8433 ( .A1(n6565), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8434 ( .A1(n6565), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8435 ( .A1(n6565), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  NOR2_X1 U8436 ( .A1(n8376), .A2(P2_U3151), .ZN(n7887) );
  NAND2_X1 U8437 ( .A1(n6663), .A2(n7887), .ZN(n6652) );
  MUX2_X1 U8438 ( .A(n8399), .B(n6652), .S(n6330), .Z(n10284) );
  INV_X1 U8439 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6656) );
  INV_X1 U8440 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6928) );
  INV_X1 U8441 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6653) );
  MUX2_X1 U8442 ( .A(n6928), .B(n6653), .S(n8376), .Z(n6722) );
  AND2_X1 U8443 ( .A1(n6722), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6723) );
  MUX2_X1 U8444 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n8376), .Z(n6690) );
  XNOR2_X1 U8445 ( .A(n6690), .B(n6689), .ZN(n6692) );
  XOR2_X1 U8446 ( .A(n6723), .B(n6692), .Z(n6654) );
  INV_X1 U8447 ( .A(n6330), .ZN(n8375) );
  NOR2_X2 U8448 ( .A1(n8399), .A2(n8375), .ZN(n10298) );
  NAND2_X1 U8449 ( .A1(n6654), .A2(n10298), .ZN(n6655) );
  OAI21_X1 U8450 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n6656), .A(n6655), .ZN(n6657) );
  INV_X1 U8451 ( .A(n6657), .ZN(n6672) );
  INV_X1 U8452 ( .A(n6658), .ZN(n7012) );
  NOR2_X1 U8453 ( .A1(n6866), .A2(n7012), .ZN(n6659) );
  OR2_X1 U8454 ( .A1(P2_U3150), .A2(n6659), .ZN(n10283) );
  INV_X1 U8455 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10368) );
  INV_X1 U8456 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6725) );
  AND2_X1 U8457 ( .A1(n6725), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6660) );
  NAND2_X1 U8458 ( .A1(n5934), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8459 ( .B1(n6689), .B2(n6660), .A(n6709), .ZN(n6662) );
  INV_X1 U8460 ( .A(n6710), .ZN(n6661) );
  AOI21_X1 U8461 ( .B1(n10368), .B2(n6662), .A(n6661), .ZN(n6669) );
  NOR2_X1 U8462 ( .A1(n6330), .A2(P2_U3151), .ZN(n7912) );
  NAND2_X1 U8463 ( .A1(n7912), .A2(n6663), .ZN(n6727) );
  AND2_X1 U8464 ( .A1(n6725), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8465 ( .A1(n5934), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6700) );
  OAI21_X1 U8466 ( .B1(n6689), .B2(n6665), .A(n6700), .ZN(n6667) );
  OR2_X1 U8467 ( .A1(n6667), .A2(n5919), .ZN(n6701) );
  INV_X1 U8468 ( .A(n6701), .ZN(n6666) );
  AOI21_X1 U8469 ( .B1(n5919), .B2(n6667), .A(n6666), .ZN(n6668) );
  OAI22_X1 U8470 ( .A1(n6669), .A2(n10293), .B1(n10302), .B2(n6668), .ZN(n6670) );
  AOI21_X1 U8471 ( .B1(n10096), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n6670), .ZN(
        n6671) );
  OAI211_X1 U8472 ( .C1(n10284), .C2(n6689), .A(n6672), .B(n6671), .ZN(
        P2_U3183) );
  AND2_X1 U8473 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9201) );
  INV_X1 U8474 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U8475 ( .A1(n6679), .A2(n7272), .ZN(n9670) );
  MUX2_X1 U8476 ( .A(n6673), .B(P1_REG2_REG_8__SCAN_IN), .S(n9677), .Z(n9669)
         );
  OAI21_X1 U8477 ( .B1(n9671), .B2(n9670), .A(n9669), .ZN(n9673) );
  OAI21_X1 U8478 ( .B1(n6673), .B2(n9677), .A(n9673), .ZN(n10104) );
  MUX2_X1 U8479 ( .A(n7457), .B(P1_REG2_REG_9__SCAN_IN), .S(n10111), .Z(n6674)
         );
  INV_X1 U8480 ( .A(n6674), .ZN(n10105) );
  NOR2_X1 U8481 ( .A1(n10104), .A2(n10105), .ZN(n10103) );
  AOI21_X1 U8482 ( .B1(n7457), .B2(n10111), .A(n10103), .ZN(n6676) );
  MUX2_X1 U8483 ( .A(n7352), .B(P1_REG2_REG_10__SCAN_IN), .S(n6807), .Z(n6675)
         );
  NAND2_X1 U8484 ( .A1(n6676), .A2(n6675), .ZN(n6802) );
  OAI211_X1 U8485 ( .C1(n6676), .C2(n6675), .A(n6802), .B(n10158), .ZN(n6677)
         );
  OAI21_X1 U8486 ( .B1(n10171), .B2(n10417), .A(n6677), .ZN(n6678) );
  NOR2_X1 U8487 ( .A1(n9201), .A2(n6678), .ZN(n6687) );
  OR2_X1 U8488 ( .A1(n6679), .A2(n6628), .ZN(n9679) );
  NAND2_X1 U8489 ( .A1(n9680), .A2(n9679), .ZN(n6682) );
  INV_X1 U8490 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6680) );
  MUX2_X1 U8491 ( .A(n6680), .B(P1_REG1_REG_8__SCAN_IN), .S(n9677), .Z(n6681)
         );
  NAND2_X1 U8492 ( .A1(n6682), .A2(n6681), .ZN(n9682) );
  OR2_X1 U8493 ( .A1(n9677), .A2(n6680), .ZN(n6683) );
  NAND2_X1 U8494 ( .A1(n9682), .A2(n6683), .ZN(n10107) );
  MUX2_X1 U8495 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n8990), .S(n10111), .Z(n10106) );
  NOR2_X1 U8496 ( .A1(n10107), .A2(n10106), .ZN(n10109) );
  AOI21_X1 U8497 ( .B1(n8990), .B2(n10111), .A(n10109), .ZN(n6685) );
  MUX2_X1 U8498 ( .A(n8991), .B(P1_REG1_REG_10__SCAN_IN), .S(n6807), .Z(n6684)
         );
  NAND2_X1 U8499 ( .A1(n6685), .A2(n6684), .ZN(n6806) );
  OAI211_X1 U8500 ( .C1(n6685), .C2(n6684), .A(n6806), .B(n10175), .ZN(n6686)
         );
  OAI211_X1 U8501 ( .C1(n9674), .C2(n6807), .A(n6687), .B(n6686), .ZN(P1_U3253) );
  NAND2_X1 U8502 ( .A1(n7132), .A2(P2_U3893), .ZN(n6688) );
  OAI21_X1 U8503 ( .B1(P2_U3893), .B2(n5119), .A(n6688), .ZN(P2_U3491) );
  INV_X1 U8504 ( .A(n6690), .ZN(n6691) );
  OAI22_X1 U8505 ( .A1(n6692), .A2(n6723), .B1(n5937), .B2(n6691), .ZN(n10237)
         );
  MUX2_X1 U8506 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8376), .Z(n6693) );
  XNOR2_X1 U8507 ( .A(n6693), .B(n6711), .ZN(n10238) );
  AOI22_X1 U8508 ( .A1(n10237), .A2(n10238), .B1(n6693), .B2(n5959), .ZN(n6695) );
  MUX2_X1 U8509 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8376), .Z(n6753) );
  XNOR2_X1 U8510 ( .A(n6753), .B(n6754), .ZN(n6694) );
  NAND2_X1 U8511 ( .A1(n6695), .A2(n6694), .ZN(n6758) );
  OAI21_X1 U8512 ( .B1(n6695), .B2(n6694), .A(n6758), .ZN(n6696) );
  NAND2_X1 U8513 ( .A1(n6696), .A2(n10298), .ZN(n6720) );
  INV_X1 U8514 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9025) );
  INV_X1 U8515 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6697) );
  NAND2_X1 U8516 ( .A1(n6699), .A2(n6698), .ZN(n10231) );
  NAND2_X1 U8517 ( .A1(n6701), .A2(n6700), .ZN(n10230) );
  NAND2_X1 U8518 ( .A1(n10231), .A2(n10230), .ZN(n10229) );
  OR2_X1 U8519 ( .A1(n6711), .A2(n6697), .ZN(n6702) );
  NAND2_X1 U8520 ( .A1(n10229), .A2(n6702), .ZN(n6703) );
  NAND2_X1 U8521 ( .A1(n6703), .A2(n6721), .ZN(n6766) );
  NAND2_X1 U8522 ( .A1(n6766), .A2(n6704), .ZN(n6706) );
  INV_X1 U8523 ( .A(n6768), .ZN(n6705) );
  AOI21_X1 U8524 ( .B1(n9025), .B2(n6706), .A(n6705), .ZN(n6707) );
  NAND2_X1 U8525 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7021) );
  OAI21_X1 U8526 ( .B1(n10302), .B2(n6707), .A(n7021), .ZN(n6718) );
  INV_X1 U8527 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6708) );
  OR2_X1 U8528 ( .A1(n6711), .A2(n6708), .ZN(n6712) );
  NAND2_X1 U8529 ( .A1(n6713), .A2(n6721), .ZN(n6761) );
  INV_X1 U8530 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10372) );
  NAND2_X1 U8531 ( .A1(n6715), .A2(n10372), .ZN(n6716) );
  AOI21_X1 U8532 ( .B1(n6763), .B2(n6716), .A(n10293), .ZN(n6717) );
  AOI211_X1 U8533 ( .C1(P2_ADDR_REG_3__SCAN_IN), .C2(n10096), .A(n6718), .B(
        n6717), .ZN(n6719) );
  OAI211_X1 U8534 ( .C1(n10284), .C2(n6721), .A(n6720), .B(n6719), .ZN(
        P2_U3185) );
  INV_X1 U8535 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6731) );
  INV_X1 U8536 ( .A(n10298), .ZN(n10091) );
  INV_X1 U8537 ( .A(n6722), .ZN(n6724) );
  AOI21_X1 U8538 ( .B1(n6725), .B2(n6724), .A(n6723), .ZN(n6726) );
  AOI21_X1 U8539 ( .B1(n6727), .B2(n10091), .A(n6726), .ZN(n6728) );
  AOI21_X1 U8540 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .A(n6728), .ZN(
        n6730) );
  INV_X1 U8541 ( .A(n10284), .ZN(n10270) );
  NAND2_X1 U8542 ( .A1(n10270), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6729) );
  OAI211_X1 U8543 ( .C1(n10283), .C2(n6731), .A(n6730), .B(n6729), .ZN(
        P2_U3182) );
  INV_X1 U8544 ( .A(n6732), .ZN(n6779) );
  AOI22_X1 U8545 ( .A1(n8438), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n9166), .ZN(n6733) );
  OAI21_X1 U8546 ( .B1(n6779), .B2(n9169), .A(n6733), .ZN(P2_U3282) );
  XNOR2_X1 U8547 ( .A(n6735), .B(n6734), .ZN(n6842) );
  MUX2_X1 U8548 ( .A(n6842), .B(n6736), .S(n9610), .Z(n6737) );
  NAND2_X1 U8549 ( .A1(n6737), .A2(n7909), .ZN(n6738) );
  OAI211_X1 U8550 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n6739), .A(n6738), .B(
        P1_U3973), .ZN(n9668) );
  AOI22_X1 U8551 ( .A1(n10155), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n6751) );
  NAND2_X1 U8552 ( .A1(n10173), .A2(n6740), .ZN(n6750) );
  INV_X1 U8553 ( .A(n6741), .ZN(n6742) );
  XNOR2_X1 U8554 ( .A(n6743), .B(n6742), .ZN(n6744) );
  NAND2_X1 U8555 ( .A1(n10158), .A2(n6744), .ZN(n6749) );
  OAI211_X1 U8556 ( .C1(n6747), .C2(n6746), .A(n10175), .B(n6745), .ZN(n6748)
         );
  AND4_X1 U8557 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6752)
         );
  NAND2_X1 U8558 ( .A1(n9668), .A2(n6752), .ZN(P1_U3245) );
  INV_X1 U8559 ( .A(n6753), .ZN(n6755) );
  NAND2_X1 U8560 ( .A1(n6755), .A2(n6754), .ZN(n6757) );
  MUX2_X1 U8561 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8376), .Z(n6780) );
  XNOR2_X1 U8562 ( .A(n6780), .B(n6783), .ZN(n6756) );
  NAND3_X1 U8563 ( .A1(n6758), .A2(n6757), .A3(n6756), .ZN(n6781) );
  NAND2_X1 U8564 ( .A1(n6781), .A2(n10298), .ZN(n6777) );
  AOI21_X1 U8565 ( .B1(n6758), .B2(n6757), .A(n6756), .ZN(n6776) );
  NOR2_X1 U8566 ( .A1(n10284), .A2(n6790), .ZN(n6774) );
  INV_X1 U8567 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10374) );
  MUX2_X1 U8568 ( .A(n10374), .B(P2_REG1_REG_4__SCAN_IN), .S(n6783), .Z(n6760)
         );
  NAND2_X1 U8569 ( .A1(n6759), .A2(n6760), .ZN(n6792) );
  INV_X1 U8570 ( .A(n6760), .ZN(n6762) );
  NAND3_X1 U8571 ( .A1(n6763), .A2(n6762), .A3(n6761), .ZN(n6764) );
  AND2_X1 U8572 ( .A1(n6792), .A2(n6764), .ZN(n6772) );
  INV_X1 U8573 ( .A(n10302), .ZN(n10233) );
  XNOR2_X1 U8574 ( .A(n6783), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n6765) );
  INV_X1 U8575 ( .A(n6765), .ZN(n6767) );
  NAND3_X1 U8576 ( .A1(n6768), .A2(n6767), .A3(n6766), .ZN(n6769) );
  NAND2_X1 U8577 ( .A1(n6785), .A2(n6769), .ZN(n6770) );
  NAND2_X1 U8578 ( .A1(n10233), .A2(n6770), .ZN(n6771) );
  NAND2_X1 U8579 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7218) );
  OAI211_X1 U8580 ( .C1(n6772), .C2(n10293), .A(n6771), .B(n7218), .ZN(n6773)
         );
  AOI211_X1 U8581 ( .C1(n10096), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6774), .B(
        n6773), .ZN(n6775) );
  OAI21_X1 U8582 ( .B1(n6777), .B2(n6776), .A(n6775), .ZN(P2_U3186) );
  OAI222_X1 U8583 ( .A1(n7411), .A2(P1_U3086), .B1(n7911), .B2(n6779), .C1(
        n6778), .C2(n7682), .ZN(P1_U3342) );
  INV_X1 U8584 ( .A(n6780), .ZN(n6782) );
  OAI21_X1 U8585 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(n7036) );
  MUX2_X1 U8586 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8376), .Z(n7034) );
  XNOR2_X1 U8587 ( .A(n7034), .B(n6799), .ZN(n7035) );
  XNOR2_X1 U8588 ( .A(n7036), .B(n7035), .ZN(n6801) );
  INV_X1 U8589 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n6797) );
  NAND2_X1 U8590 ( .A1(n6790), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6784) );
  INV_X1 U8591 ( .A(n6786), .ZN(n6787) );
  NAND2_X1 U8592 ( .A1(n6787), .A2(n4709), .ZN(n6788) );
  NAND2_X1 U8593 ( .A1(n7050), .A2(n6788), .ZN(n6789) );
  AND2_X1 U8594 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7395) );
  AOI21_X1 U8595 ( .B1(n10233), .B2(n6789), .A(n7395), .ZN(n6796) );
  INV_X1 U8596 ( .A(n10293), .ZN(n10228) );
  NAND2_X1 U8597 ( .A1(n6790), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8598 ( .A1(n6792), .A2(n6791), .ZN(n7027) );
  XNOR2_X1 U8599 ( .A(n7027), .B(n6799), .ZN(n6793) );
  OAI21_X1 U8600 ( .B1(n6793), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7029), .ZN(
        n6794) );
  NAND2_X1 U8601 ( .A1(n10228), .A2(n6794), .ZN(n6795) );
  OAI211_X1 U8602 ( .C1(n6797), .C2(n10283), .A(n6796), .B(n6795), .ZN(n6798)
         );
  AOI21_X1 U8603 ( .B1(n6799), .B2(n10270), .A(n6798), .ZN(n6800) );
  OAI21_X1 U8604 ( .B1(n6801), .B2(n10091), .A(n6800), .ZN(P2_U3187) );
  AOI22_X1 U8605 ( .A1(n7408), .A2(n7516), .B1(P1_REG2_REG_12__SCAN_IN), .B2(
        n6809), .ZN(n6805) );
  OAI21_X1 U8606 ( .B1(n7352), .B2(n6807), .A(n6802), .ZN(n10125) );
  MUX2_X1 U8607 ( .A(n6803), .B(P1_REG2_REG_11__SCAN_IN), .S(n10118), .Z(
        n10124) );
  NAND2_X1 U8608 ( .A1(n10125), .A2(n10124), .ZN(n10123) );
  OAI21_X1 U8609 ( .B1(n6803), .B2(n10118), .A(n10123), .ZN(n6804) );
  NOR2_X1 U8610 ( .A1(n6805), .A2(n6804), .ZN(n7409) );
  AOI21_X1 U8611 ( .B1(n6805), .B2(n6804), .A(n7409), .ZN(n6818) );
  OAI21_X1 U8612 ( .B1(n8991), .B2(n6807), .A(n6806), .ZN(n10122) );
  MUX2_X1 U8613 ( .A(n6808), .B(P1_REG1_REG_11__SCAN_IN), .S(n10118), .Z(
        n10121) );
  NAND2_X1 U8614 ( .A1(n10122), .A2(n10121), .ZN(n10120) );
  OAI21_X1 U8615 ( .B1(n6808), .B2(n10118), .A(n10120), .ZN(n6811) );
  AOI22_X1 U8616 ( .A1(n7408), .A2(n5410), .B1(P1_REG1_REG_12__SCAN_IN), .B2(
        n6809), .ZN(n6810) );
  NOR2_X1 U8617 ( .A1(n6811), .A2(n6810), .ZN(n7400) );
  AOI21_X1 U8618 ( .B1(n6811), .B2(n6810), .A(n7400), .ZN(n6815) );
  AND2_X1 U8619 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6812) );
  AOI21_X1 U8620 ( .B1(n10155), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n6812), .ZN(
        n6814) );
  NAND2_X1 U8621 ( .A1(n10173), .A2(n7408), .ZN(n6813) );
  OAI211_X1 U8622 ( .C1(n6815), .C2(n9701), .A(n6814), .B(n6813), .ZN(n6816)
         );
  INV_X1 U8623 ( .A(n6816), .ZN(n6817) );
  OAI21_X1 U8624 ( .B1(n6818), .B2(n10182), .A(n6817), .ZN(P1_U3255) );
  NOR2_X1 U8625 ( .A1(n9337), .A2(P1_U3086), .ZN(n6846) );
  INV_X1 U8626 ( .A(n6819), .ZN(n6822) );
  NOR3_X1 U8627 ( .A1(n6822), .A2(n6821), .A3(n6820), .ZN(n6825) );
  INV_X1 U8628 ( .A(n6823), .ZN(n6824) );
  OAI21_X1 U8629 ( .B1(n6825), .B2(n6824), .A(n9329), .ZN(n6829) );
  OAI22_X1 U8630 ( .A1(n6827), .A2(n9301), .B1(n6826), .B2(n9300), .ZN(n6962)
         );
  AOI22_X1 U8631 ( .A1(n9351), .A2(n7140), .B1(n9346), .B2(n6962), .ZN(n6828)
         );
  OAI211_X1 U8632 ( .C1(n6846), .C2(n6830), .A(n6829), .B(n6828), .ZN(P1_U3237) );
  INV_X1 U8633 ( .A(n6831), .ZN(n6833) );
  OAI222_X1 U8634 ( .A1(n9171), .A2(n6832), .B1(n9169), .B2(n6833), .C1(
        P2_U3151), .C2(n8451), .ZN(P2_U3281) );
  OAI222_X1 U8635 ( .A1(n7407), .A2(P1_U3086), .B1(n7911), .B2(n6833), .C1(
        n9016), .C2(n7682), .ZN(P1_U3341) );
  INV_X1 U8636 ( .A(n9647), .ZN(n6834) );
  OAI22_X1 U8637 ( .A1(n6835), .A2(n9301), .B1(n6834), .B2(n9300), .ZN(n6972)
         );
  AOI22_X1 U8638 ( .A1(n9351), .A2(n6977), .B1(n9346), .B2(n6972), .ZN(n6840)
         );
  OAI21_X1 U8639 ( .B1(n6837), .B2(n6836), .A(n6819), .ZN(n6838) );
  NAND2_X1 U8640 ( .A1(n6838), .A2(n9329), .ZN(n6839) );
  OAI211_X1 U8641 ( .C1(n6846), .C2(n6841), .A(n6840), .B(n6839), .ZN(P1_U3222) );
  INV_X1 U8642 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6845) );
  NAND2_X1 U8643 ( .A1(n6380), .A2(n9321), .ZN(n7096) );
  OAI22_X1 U8644 ( .A1(n9323), .A2(n7096), .B1(n9354), .B2(n6842), .ZN(n6843)
         );
  AOI21_X1 U8645 ( .B1(n6975), .B2(n9351), .A(n6843), .ZN(n6844) );
  OAI21_X1 U8646 ( .B1(n6846), .B2(n6845), .A(n6844), .ZN(P1_U3232) );
  OAI21_X1 U8647 ( .B1(n6849), .B2(n6848), .A(n6847), .ZN(n6856) );
  NAND2_X1 U8648 ( .A1(n9645), .A2(n9320), .ZN(n6851) );
  NAND2_X1 U8649 ( .A1(n9644), .A2(n9321), .ZN(n6850) );
  NAND2_X1 U8650 ( .A1(n6851), .A2(n6850), .ZN(n6984) );
  AOI21_X1 U8651 ( .B1(n9346), .B2(n6984), .A(n6852), .ZN(n6854) );
  INV_X1 U8652 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n7116) );
  NAND2_X1 U8653 ( .A1(n9337), .A2(n7116), .ZN(n6853) );
  OAI211_X1 U8654 ( .C1(n9283), .C2(n7365), .A(n6854), .B(n6853), .ZN(n6855)
         );
  AOI21_X1 U8655 ( .B1(n6856), .B2(n9329), .A(n6855), .ZN(n6857) );
  INV_X1 U8656 ( .A(n6857), .ZN(P1_U3218) );
  INV_X1 U8657 ( .A(n6911), .ZN(n6931) );
  NAND2_X1 U8658 ( .A1(n7132), .A2(n6931), .ZN(n8164) );
  AND2_X1 U8659 ( .A1(n8167), .A2(n8164), .ZN(n8343) );
  INV_X1 U8660 ( .A(n6858), .ZN(n6859) );
  NAND2_X1 U8661 ( .A1(n6860), .A2(n6859), .ZN(n6863) );
  INV_X1 U8662 ( .A(n6861), .ZN(n6868) );
  NAND2_X1 U8663 ( .A1(n6890), .A2(n6868), .ZN(n6862) );
  INV_X1 U8664 ( .A(n6864), .ZN(n6865) );
  NAND2_X1 U8665 ( .A1(n6866), .A2(n6865), .ZN(n6867) );
  AOI21_X1 U8666 ( .B1(n6872), .B2(n6868), .A(n6867), .ZN(n6871) );
  NAND2_X1 U8667 ( .A1(n6879), .A2(n6869), .ZN(n6870) );
  NAND2_X1 U8668 ( .A1(n6871), .A2(n6870), .ZN(n6874) );
  NOR2_X1 U8669 ( .A1(n6925), .A2(n6887), .ZN(n8377) );
  AND2_X1 U8670 ( .A1(n6872), .A2(n8377), .ZN(n6873) );
  AOI21_X1 U8671 ( .B1(n6874), .B2(P2_STATE_REG_SCAN_IN), .A(n6873), .ZN(n7013) );
  AND2_X1 U8672 ( .A1(n7013), .A2(n6875), .ZN(n6940) );
  INV_X1 U8673 ( .A(n6940), .ZN(n6876) );
  NAND2_X1 U8674 ( .A1(n6876), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6883) );
  INV_X1 U8675 ( .A(n6887), .ZN(n6921) );
  AND2_X1 U8676 ( .A1(n6888), .A2(n6921), .ZN(n6877) );
  NAND2_X1 U8677 ( .A1(n6890), .A2(n6877), .ZN(n8127) );
  NAND2_X1 U8678 ( .A1(n6879), .A2(n6878), .ZN(n6881) );
  NOR2_X1 U8679 ( .A1(n6925), .A2(n10359), .ZN(n6880) );
  AND2_X2 U8680 ( .A1(n6881), .A2(n6880), .ZN(n8119) );
  AOI22_X1 U8681 ( .A1(n8137), .A2(n5940), .B1(n8119), .B2(n6911), .ZN(n6882)
         );
  OAI211_X1 U8682 ( .C1(n8343), .C2(n8131), .A(n6883), .B(n6882), .ZN(P2_U3172) );
  NAND2_X1 U8683 ( .A1(n9646), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6884) );
  OAI21_X1 U8684 ( .B1(n6885), .B2(n9646), .A(n6884), .ZN(P1_U3583) );
  INV_X1 U8685 ( .A(n6886), .ZN(n6909) );
  INV_X1 U8686 ( .A(n8490), .ZN(n8481) );
  INV_X1 U8687 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9020) );
  OAI222_X1 U8688 ( .A1(n9169), .A2(n6909), .B1(n8481), .B2(P2_U3151), .C1(
        n9020), .C2(n9171), .ZN(P2_U3280) );
  INV_X1 U8689 ( .A(n8119), .ZN(n8145) );
  NOR2_X1 U8690 ( .A1(n6888), .A2(n6887), .ZN(n6889) );
  NAND2_X1 U8691 ( .A1(n6890), .A2(n6889), .ZN(n8139) );
  OAI22_X1 U8692 ( .A1(n8145), .A2(n10319), .B1(n8139), .B2(n6280), .ZN(n6891)
         );
  AOI21_X1 U8693 ( .B1(n8137), .B2(n8400), .A(n6891), .ZN(n6907) );
  INV_X1 U8694 ( .A(n8340), .ZN(n6892) );
  NAND2_X1 U8695 ( .A1(n6893), .A2(n6892), .ZN(n6897) );
  NAND2_X1 U8696 ( .A1(n8165), .A2(n8329), .ZN(n6895) );
  AND2_X1 U8697 ( .A1(n6895), .A2(n6894), .ZN(n6896) );
  INV_X1 U8698 ( .A(n6900), .ZN(n6898) );
  NAND2_X1 U8699 ( .A1(n6898), .A2(n5940), .ZN(n6901) );
  NAND2_X1 U8700 ( .A1(n6900), .A2(n6899), .ZN(n6932) );
  OAI21_X1 U8701 ( .B1(n6903), .B2(n6904), .A(n6933), .ZN(n6905) );
  INV_X1 U8702 ( .A(n8131), .ZN(n8133) );
  NAND2_X1 U8703 ( .A1(n6905), .A2(n8133), .ZN(n6906) );
  OAI211_X1 U8704 ( .C1(n6940), .C2(n6656), .A(n6907), .B(n6906), .ZN(P2_U3162) );
  OAI222_X1 U8705 ( .A1(P1_U3086), .A2(n7413), .B1(n7911), .B2(n6909), .C1(
        n6908), .C2(n7682), .ZN(P1_U3340) );
  NOR2_X1 U8706 ( .A1(n6899), .A2(n8678), .ZN(n6922) );
  AOI21_X1 U8707 ( .B1(n8673), .B2(n10353), .A(n8343), .ZN(n6910) );
  AOI211_X1 U8708 ( .C1(n10325), .C2(n6911), .A(n6922), .B(n6910), .ZN(n6941)
         );
  NAND2_X1 U8709 ( .A1(n10365), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6912) );
  OAI21_X1 U8710 ( .B1(n6941), .B2(n10365), .A(n6912), .ZN(P2_U3390) );
  INV_X1 U8711 ( .A(n6913), .ZN(n6944) );
  AOI22_X1 U8712 ( .A1(n8523), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9166), .ZN(n6914) );
  OAI21_X1 U8713 ( .B1(n6944), .B2(n9169), .A(n6914), .ZN(P2_U3279) );
  INV_X1 U8714 ( .A(n6915), .ZN(n6920) );
  INV_X1 U8715 ( .A(n6916), .ZN(n6917) );
  NOR2_X1 U8716 ( .A1(n6918), .A2(n6917), .ZN(n6919) );
  NAND2_X1 U8717 ( .A1(n6920), .A2(n6919), .ZN(n6926) );
  NOR3_X1 U8718 ( .A1(n8343), .A2(n6921), .A3(n10325), .ZN(n6923) );
  NOR2_X1 U8719 ( .A1(n6923), .A2(n6922), .ZN(n6927) );
  MUX2_X1 U8720 ( .A(n6928), .B(n6927), .S(n10317), .Z(n6930) );
  NAND2_X1 U8721 ( .A1(n10314), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6929) );
  OAI211_X1 U8722 ( .C1(n8699), .C2(n6931), .A(n6930), .B(n6929), .ZN(P2_U3233) );
  INV_X1 U8723 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n9027) );
  XNOR2_X1 U8724 ( .A(n7014), .B(n7022), .ZN(n6935) );
  NAND2_X1 U8725 ( .A1(n6936), .A2(n8133), .ZN(n6939) );
  OAI22_X1 U8726 ( .A1(n8145), .A2(n7232), .B1(n8139), .B2(n6899), .ZN(n6937)
         );
  AOI21_X1 U8727 ( .B1(n8137), .B2(n8398), .A(n6937), .ZN(n6938) );
  OAI211_X1 U8728 ( .C1(n6940), .C2(n9027), .A(n6939), .B(n6938), .ZN(P2_U3177) );
  OR2_X1 U8729 ( .A1(n6941), .A2(n6377), .ZN(n6942) );
  OAI21_X1 U8730 ( .B1(n10384), .B2(n6653), .A(n6942), .ZN(P2_U3459) );
  OAI222_X1 U8731 ( .A1(n7574), .A2(P1_U3086), .B1(n7911), .B2(n6944), .C1(
        n6943), .C2(n7682), .ZN(P1_U3339) );
  OAI21_X1 U8732 ( .B1(n6946), .B2(n9544), .A(n6945), .ZN(n7106) );
  AOI211_X1 U8733 ( .C1(n6947), .C2(n6986), .A(n9922), .B(n7073), .ZN(n7111)
         );
  INV_X1 U8734 ( .A(n9544), .ZN(n9421) );
  XNOR2_X1 U8735 ( .A(n6948), .B(n9421), .ZN(n6952) );
  OR2_X1 U8736 ( .A1(n7153), .A2(n9301), .ZN(n6950) );
  NAND2_X1 U8737 ( .A1(n6385), .A2(n9320), .ZN(n6949) );
  NAND2_X1 U8738 ( .A1(n6950), .A2(n6949), .ZN(n7004) );
  INV_X1 U8739 ( .A(n7004), .ZN(n6951) );
  OAI21_X1 U8740 ( .B1(n6952), .B2(n9906), .A(n6951), .ZN(n7107) );
  AOI211_X1 U8741 ( .C1(n10217), .C2(n7106), .A(n7111), .B(n7107), .ZN(n7334)
         );
  OAI22_X1 U8742 ( .A1(n10001), .A2(n7331), .B1(n10223), .B2(n6605), .ZN(n6953) );
  INV_X1 U8743 ( .A(n6953), .ZN(n6954) );
  OAI21_X1 U8744 ( .B1(n7334), .B2(n6496), .A(n6954), .ZN(P1_U3526) );
  OAI21_X1 U8745 ( .B1(n6956), .B2(n6958), .A(n6955), .ZN(n7145) );
  INV_X1 U8746 ( .A(n7145), .ZN(n6964) );
  INV_X1 U8747 ( .A(n7290), .ZN(n7672) );
  NAND3_X1 U8748 ( .A1(n6971), .A2(n6958), .A3(n6957), .ZN(n6959) );
  AOI21_X1 U8749 ( .B1(n6960), .B2(n6959), .A(n9906), .ZN(n6961) );
  AOI211_X1 U8750 ( .C1(n7672), .C2(n7145), .A(n6962), .B(n6961), .ZN(n7147)
         );
  INV_X1 U8751 ( .A(n6987), .ZN(n6963) );
  OAI211_X1 U8752 ( .C1(n6383), .C2(n6974), .A(n6963), .B(n9777), .ZN(n7143)
         );
  OAI211_X1 U8753 ( .C1(n6964), .C2(n10208), .A(n7147), .B(n7143), .ZN(n7359)
         );
  OAI22_X1 U8754 ( .A1(n10001), .A2(n6383), .B1(n10223), .B2(n6571), .ZN(n6965) );
  AOI21_X1 U8755 ( .B1(n7359), .B2(n10223), .A(n6965), .ZN(n6966) );
  INV_X1 U8756 ( .A(n6966), .ZN(P1_U3524) );
  INV_X1 U8757 ( .A(n6968), .ZN(n6969) );
  INV_X1 U8758 ( .A(n10217), .ZN(n10018) );
  AOI21_X1 U8759 ( .B1(n6973), .B2(n9931), .A(n6972), .ZN(n7176) );
  AOI211_X1 U8760 ( .C1(n6975), .C2(n6977), .A(n9922), .B(n6974), .ZN(n7174)
         );
  INV_X1 U8761 ( .A(n7174), .ZN(n6976) );
  OAI211_X1 U8762 ( .C1(n7171), .C2(n10018), .A(n7176), .B(n6976), .ZN(n7362)
         );
  INV_X1 U8763 ( .A(n6977), .ZN(n9383) );
  OAI22_X1 U8764 ( .A1(n10001), .A2(n9383), .B1(n10223), .B2(n6978), .ZN(n6979) );
  AOI21_X1 U8765 ( .B1(n7362), .B2(n10223), .A(n6979), .ZN(n6980) );
  INV_X1 U8766 ( .A(n6980), .ZN(P1_U3523) );
  OAI21_X1 U8767 ( .B1(n6982), .B2(n6983), .A(n6981), .ZN(n7122) );
  INV_X1 U8768 ( .A(n7122), .ZN(n6988) );
  INV_X1 U8769 ( .A(n6983), .ZN(n9542) );
  XNOR2_X1 U8770 ( .A(n9542), .B(n9425), .ZN(n6985) );
  AOI21_X1 U8771 ( .B1(n6985), .B2(n9931), .A(n6984), .ZN(n7124) );
  OAI211_X1 U8772 ( .C1(n6987), .C2(n7365), .A(n9777), .B(n6986), .ZN(n7120)
         );
  OAI211_X1 U8773 ( .C1(n6988), .C2(n10018), .A(n7124), .B(n7120), .ZN(n7367)
         );
  OAI22_X1 U8774 ( .A1(n10001), .A2(n7365), .B1(n10223), .B2(n6577), .ZN(n6989) );
  AOI21_X1 U8775 ( .B1(n7367), .B2(n10223), .A(n6989), .ZN(n6990) );
  INV_X1 U8776 ( .A(n6990), .ZN(P1_U3525) );
  INV_X1 U8777 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U8778 ( .A1(n6991), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U8779 ( .A1(n4411), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6992) );
  OAI211_X1 U8780 ( .C1(n9038), .C2(n6994), .A(n6993), .B(n6992), .ZN(n6995)
         );
  INV_X1 U8781 ( .A(n6995), .ZN(n6996) );
  NAND2_X1 U8782 ( .A1(n8399), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n6998) );
  OAI21_X1 U8783 ( .B1(n8539), .B2(n8399), .A(n6998), .ZN(P2_U3522) );
  INV_X1 U8784 ( .A(n6999), .ZN(n7000) );
  NAND2_X1 U8785 ( .A1(n9647), .A2(n7104), .ZN(n9385) );
  NAND2_X1 U8786 ( .A1(n7000), .A2(n9385), .ZN(n9540) );
  OAI21_X1 U8787 ( .B1(n10217), .B2(n9931), .A(n9540), .ZN(n7001) );
  OAI211_X1 U8788 ( .C1(n7002), .C2(n7104), .A(n7001), .B(n7096), .ZN(n10020)
         );
  NAND2_X1 U8789 ( .A1(n10020), .A2(n10220), .ZN(n7003) );
  OAI21_X1 U8790 ( .B1(n10220), .B2(n5113), .A(n7003), .ZN(P1_U3453) );
  INV_X1 U8791 ( .A(n7108), .ZN(n7010) );
  NAND2_X1 U8792 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n9649) );
  NAND2_X1 U8793 ( .A1(n9346), .A2(n7004), .ZN(n7005) );
  OAI211_X1 U8794 ( .C1(n9283), .C2(n7331), .A(n9649), .B(n7005), .ZN(n7009)
         );
  AOI211_X1 U8795 ( .C1(n7007), .C2(n7006), .A(n9354), .B(n4518), .ZN(n7008)
         );
  AOI211_X1 U8796 ( .C1(n7010), .C2(n9337), .A(n7009), .B(n7008), .ZN(n7011)
         );
  INV_X1 U8797 ( .A(n7011), .ZN(P1_U3230) );
  NAND2_X1 U8798 ( .A1(n7012), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8381) );
  OR2_X1 U8799 ( .A1(n7014), .A2(n8400), .ZN(n7015) );
  XNOR2_X1 U8800 ( .A(n8011), .B(n10331), .ZN(n7210) );
  XNOR2_X1 U8801 ( .A(n7210), .B(n8398), .ZN(n7017) );
  AOI21_X1 U8802 ( .B1(n7016), .B2(n7017), .A(n8131), .ZN(n7020) );
  INV_X1 U8803 ( .A(n7016), .ZN(n7019) );
  INV_X1 U8804 ( .A(n7017), .ZN(n7018) );
  NAND2_X1 U8805 ( .A1(n7019), .A2(n7018), .ZN(n7212) );
  NAND2_X1 U8806 ( .A1(n7020), .A2(n7212), .ZN(n7026) );
  INV_X1 U8807 ( .A(n7021), .ZN(n7024) );
  OAI22_X1 U8808 ( .A1(n7022), .A2(n8139), .B1(n8127), .B2(n7393), .ZN(n7023)
         );
  AOI211_X1 U8809 ( .C1(n8119), .C2(n7257), .A(n7024), .B(n7023), .ZN(n7025)
         );
  OAI211_X1 U8810 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n7495), .A(n7026), .B(
        n7025), .ZN(P2_U3158) );
  NAND2_X1 U8811 ( .A1(n7027), .A2(n7047), .ZN(n7028) );
  INV_X1 U8812 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U8813 ( .A1(n10254), .A2(P2_REG1_REG_6__SCAN_IN), .B1(n10376), .B2(
        n7052), .ZN(n10244) );
  NOR2_X1 U8814 ( .A1(n10269), .A2(n7031), .ZN(n7032) );
  INV_X1 U8815 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10378) );
  INV_X1 U8816 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U8817 ( .A1(n7193), .A2(P2_REG1_REG_8__SCAN_IN), .B1(n10380), .B2(
        n7056), .ZN(n7033) );
  AOI21_X1 U8818 ( .B1(n4522), .B2(n7033), .A(n7192), .ZN(n7064) );
  MUX2_X1 U8819 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8376), .Z(n7037) );
  AOI22_X1 U8820 ( .A1(n7036), .A2(n7035), .B1(n7034), .B2(n7047), .ZN(n10257)
         );
  XNOR2_X1 U8821 ( .A(n7037), .B(n10254), .ZN(n10256) );
  NAND2_X1 U8822 ( .A1(n10257), .A2(n10256), .ZN(n10255) );
  OAI21_X1 U8823 ( .B1(n7037), .B2(n7052), .A(n10255), .ZN(n10276) );
  MUX2_X1 U8824 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8376), .Z(n7039) );
  NOR2_X1 U8825 ( .A1(n7039), .A2(n7038), .ZN(n7040) );
  AOI21_X1 U8826 ( .B1(n7039), .B2(n7038), .A(n7040), .ZN(n10277) );
  NAND2_X1 U8827 ( .A1(n10276), .A2(n10277), .ZN(n10275) );
  INV_X1 U8828 ( .A(n7040), .ZN(n7041) );
  NAND2_X1 U8829 ( .A1(n10275), .A2(n7041), .ZN(n7044) );
  MUX2_X1 U8830 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8376), .Z(n7042) );
  NOR2_X1 U8831 ( .A1(n7042), .A2(n7056), .ZN(n7188) );
  AOI21_X1 U8832 ( .B1(n7042), .B2(n7056), .A(n7188), .ZN(n7043) );
  AND2_X1 U8833 ( .A1(n7044), .A2(n7043), .ZN(n7187) );
  NOR2_X1 U8834 ( .A1(n7044), .A2(n7043), .ZN(n7045) );
  OAI21_X1 U8835 ( .B1(n7187), .B2(n7045), .A(n10298), .ZN(n7063) );
  INV_X1 U8836 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U8837 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7730) );
  OAI21_X1 U8838 ( .B1(n10283), .B2(n7046), .A(n7730), .ZN(n7061) );
  NAND2_X1 U8839 ( .A1(n7048), .A2(n7047), .ZN(n7049) );
  INV_X1 U8840 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7051) );
  AOI22_X1 U8841 ( .A1(n10254), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n7051), .B2(
        n7052), .ZN(n10248) );
  NOR2_X1 U8842 ( .A1(n10269), .A2(n7053), .ZN(n7054) );
  INV_X1 U8843 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10264) );
  XNOR2_X1 U8844 ( .A(n7053), .B(n10269), .ZN(n10263) );
  NOR2_X1 U8845 ( .A1(n10264), .A2(n10263), .ZN(n10262) );
  NOR2_X1 U8846 ( .A1(n7054), .A2(n10262), .ZN(n7058) );
  INV_X1 U8847 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7055) );
  OR2_X1 U8848 ( .A1(n7193), .A2(n7055), .ZN(n7200) );
  OAI21_X1 U8849 ( .B1(n7056), .B2(P2_REG2_REG_8__SCAN_IN), .A(n7200), .ZN(
        n7057) );
  NOR2_X1 U8850 ( .A1(n7058), .A2(n7057), .ZN(n7198) );
  AOI21_X1 U8851 ( .B1(n7058), .B2(n7057), .A(n7198), .ZN(n7059) );
  NOR2_X1 U8852 ( .A1(n7059), .A2(n10302), .ZN(n7060) );
  AOI211_X1 U8853 ( .C1(n10270), .C2(n7193), .A(n7061), .B(n7060), .ZN(n7062)
         );
  OAI211_X1 U8854 ( .C1(n7064), .C2(n10293), .A(n7063), .B(n7062), .ZN(
        P2_U3190) );
  OAI21_X1 U8855 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n7091) );
  INV_X1 U8856 ( .A(n7091), .ZN(n7074) );
  NAND2_X1 U8857 ( .A1(n7068), .A2(n9423), .ZN(n7069) );
  XNOR2_X1 U8858 ( .A(n7069), .B(n9547), .ZN(n7072) );
  NAND2_X1 U8859 ( .A1(n9644), .A2(n9320), .ZN(n7071) );
  NAND2_X1 U8860 ( .A1(n9642), .A2(n9321), .ZN(n7070) );
  NAND2_X1 U8861 ( .A1(n7071), .A2(n7070), .ZN(n7180) );
  AOI21_X1 U8862 ( .B1(n7072), .B2(n9931), .A(n7180), .ZN(n7084) );
  OAI211_X1 U8863 ( .C1(n7073), .C2(n7380), .A(n9777), .B(n7150), .ZN(n7087)
         );
  OAI211_X1 U8864 ( .C1(n7074), .C2(n10018), .A(n7084), .B(n7087), .ZN(n7382)
         );
  OAI22_X1 U8865 ( .A1(n10001), .A2(n7380), .B1(n10223), .B2(n6608), .ZN(n7075) );
  AOI21_X1 U8866 ( .B1(n7382), .B2(n10223), .A(n7075), .ZN(n7076) );
  INV_X1 U8867 ( .A(n7076), .ZN(P1_U3527) );
  INV_X1 U8868 ( .A(n7077), .ZN(n7095) );
  INV_X1 U8869 ( .A(n8527), .ZN(n10285) );
  OAI222_X1 U8870 ( .A1(n9169), .A2(n7095), .B1(n10285), .B2(P2_U3151), .C1(
        n9018), .C2(n9171), .ZN(P2_U3278) );
  INV_X1 U8871 ( .A(n7078), .ZN(n7079) );
  NAND3_X1 U8872 ( .A1(n7081), .A2(n7080), .A3(n7079), .ZN(n7082) );
  MUX2_X1 U8873 ( .A(n7084), .B(n7083), .S(n4415), .Z(n7093) );
  NAND2_X1 U8874 ( .A1(n9705), .A2(n9611), .ZN(n7085) );
  OR2_X1 U8875 ( .A1(n4415), .A2(n7290), .ZN(n7086) );
  NOR2_X1 U8876 ( .A1(n7087), .A2(n9778), .ZN(n7090) );
  OR2_X2 U8877 ( .A1(n4415), .A2(n7088), .ZN(n9927) );
  OAI22_X1 U8878 ( .A1(n9927), .A2(n7380), .B1(n9774), .B2(n7179), .ZN(n7089)
         );
  AOI211_X1 U8879 ( .C1(n7091), .C2(n9876), .A(n7090), .B(n7089), .ZN(n7092)
         );
  NAND2_X1 U8880 ( .A1(n7093), .A2(n7092), .ZN(P1_U3288) );
  OAI222_X1 U8881 ( .A1(P1_U3086), .A2(n9689), .B1(n7911), .B2(n7095), .C1(
        n7094), .C2(n7682), .ZN(P1_U3338) );
  AOI21_X1 U8882 ( .B1(n10189), .B2(n9777), .A(n10186), .ZN(n7105) );
  INV_X1 U8883 ( .A(n9540), .ZN(n7099) );
  NAND2_X1 U8884 ( .A1(n10184), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7097) );
  OAI211_X1 U8885 ( .C1(n7099), .C2(n7098), .A(n7097), .B(n7096), .ZN(n7102)
         );
  NOR2_X1 U8886 ( .A1(n9916), .A2(n7100), .ZN(n7101) );
  AOI21_X1 U8887 ( .B1(n9916), .B2(n7102), .A(n7101), .ZN(n7103) );
  OAI21_X1 U8888 ( .B1(n7105), .B2(n7104), .A(n7103), .ZN(P1_U3293) );
  INV_X1 U8889 ( .A(n9876), .ZN(n9936) );
  INV_X1 U8890 ( .A(n7106), .ZN(n7114) );
  NAND2_X1 U8891 ( .A1(n7107), .A2(n9916), .ZN(n7113) );
  NOR2_X1 U8892 ( .A1(n9927), .A2(n7331), .ZN(n7110) );
  OAI22_X1 U8893 ( .A1(n9916), .A2(n6596), .B1(n7108), .B2(n9774), .ZN(n7109)
         );
  AOI211_X1 U8894 ( .C1(n7111), .C2(n10189), .A(n7110), .B(n7109), .ZN(n7112)
         );
  OAI211_X1 U8895 ( .C1(n9936), .C2(n7114), .A(n7113), .B(n7112), .ZN(P1_U3289) );
  INV_X1 U8896 ( .A(n7115), .ZN(n7160) );
  INV_X1 U8897 ( .A(n10092), .ZN(n10101) );
  INV_X1 U8898 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n8974) );
  OAI222_X1 U8899 ( .A1(n9169), .A2(n7160), .B1(n10101), .B2(P2_U3151), .C1(
        n8974), .C2(n9171), .ZN(P2_U3277) );
  INV_X1 U8900 ( .A(n7365), .ZN(n7118) );
  OAI22_X1 U8901 ( .A1(n9916), .A2(n6594), .B1(n9774), .B2(
        P1_REG3_REG_3__SCAN_IN), .ZN(n7117) );
  AOI21_X1 U8902 ( .B1(n10186), .B2(n7118), .A(n7117), .ZN(n7119) );
  OAI21_X1 U8903 ( .B1(n9778), .B2(n7120), .A(n7119), .ZN(n7121) );
  AOI21_X1 U8904 ( .B1(n9876), .B2(n7122), .A(n7121), .ZN(n7123) );
  OAI21_X1 U8905 ( .B1(n4415), .B2(n7124), .A(n7123), .ZN(P1_U3290) );
  NAND2_X1 U8906 ( .A1(n7125), .A2(n8165), .ZN(n7239) );
  NOR2_X1 U8907 ( .A1(n8741), .A2(n7239), .ZN(n8548) );
  INV_X1 U8908 ( .A(n8548), .ZN(n7237) );
  NAND2_X1 U8909 ( .A1(n8342), .A2(n8167), .ZN(n7126) );
  NAND2_X1 U8910 ( .A1(n7127), .A2(n7126), .ZN(n7128) );
  INV_X1 U8911 ( .A(n7128), .ZN(n10320) );
  NAND2_X1 U8912 ( .A1(n7128), .A2(n7775), .ZN(n7135) );
  OAI21_X1 U8913 ( .B1(n7130), .B2(n8342), .A(n7129), .ZN(n7131) );
  NAND2_X1 U8914 ( .A1(n7131), .A2(n8722), .ZN(n7134) );
  AOI22_X1 U8915 ( .A1(n7132), .A2(n8719), .B1(n8717), .B2(n8400), .ZN(n7133)
         );
  NAND3_X1 U8916 ( .A1(n7135), .A2(n7134), .A3(n7133), .ZN(n10321) );
  MUX2_X1 U8917 ( .A(n10321), .B(P2_REG2_REG_1__SCAN_IN), .S(n8741), .Z(n7136)
         );
  INV_X1 U8918 ( .A(n7136), .ZN(n7139) );
  AOI22_X1 U8919 ( .A1(n10312), .A2(n7137), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10314), .ZN(n7138) );
  OAI211_X1 U8920 ( .C1(n7237), .C2(n10320), .A(n7139), .B(n7138), .ZN(
        P2_U3232) );
  INV_X1 U8921 ( .A(n7297), .ZN(n10190) );
  NAND2_X1 U8922 ( .A1(n10186), .A2(n7140), .ZN(n7142) );
  AOI22_X1 U8923 ( .A1(n4415), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n10184), .ZN(n7141) );
  OAI211_X1 U8924 ( .C1(n7143), .C2(n9778), .A(n7142), .B(n7141), .ZN(n7144)
         );
  AOI21_X1 U8925 ( .B1(n10190), .B2(n7145), .A(n7144), .ZN(n7146) );
  OAI21_X1 U8926 ( .B1(n7147), .B2(n4415), .A(n7146), .ZN(P1_U3291) );
  OAI21_X1 U8927 ( .B1(n7149), .B2(n7265), .A(n7148), .ZN(n7161) );
  AOI21_X1 U8928 ( .B1(n7150), .B2(n9334), .A(n9922), .ZN(n7152) );
  AND2_X1 U8929 ( .A1(n7152), .A2(n7273), .ZN(n7166) );
  XNOR2_X1 U8930 ( .A(n7264), .B(n9548), .ZN(n7157) );
  OR2_X1 U8931 ( .A1(n7153), .A2(n9300), .ZN(n7155) );
  OR2_X1 U8932 ( .A1(n7280), .A2(n9301), .ZN(n7154) );
  NAND2_X1 U8933 ( .A1(n7155), .A2(n7154), .ZN(n9333) );
  INV_X1 U8934 ( .A(n9333), .ZN(n7156) );
  OAI21_X1 U8935 ( .B1(n7157), .B2(n9906), .A(n7156), .ZN(n7162) );
  AOI211_X1 U8936 ( .C1(n10217), .C2(n7161), .A(n7166), .B(n7162), .ZN(n7339)
         );
  OAI22_X1 U8937 ( .A1(n10001), .A2(n7336), .B1(n10223), .B2(n6627), .ZN(n7158) );
  INV_X1 U8938 ( .A(n7158), .ZN(n7159) );
  OAI21_X1 U8939 ( .B1(n7339), .B2(n6496), .A(n7159), .ZN(P1_U3528) );
  OAI222_X1 U8940 ( .A1(P1_U3086), .A2(n10170), .B1(n7911), .B2(n7160), .C1(
        n9017), .C2(n7682), .ZN(P1_U3337) );
  INV_X1 U8941 ( .A(n7161), .ZN(n7169) );
  INV_X1 U8942 ( .A(n7162), .ZN(n7164) );
  MUX2_X1 U8943 ( .A(n7164), .B(n7163), .S(n4415), .Z(n7168) );
  OAI22_X1 U8944 ( .A1(n9927), .A2(n7336), .B1(n9774), .B2(n9335), .ZN(n7165)
         );
  AOI21_X1 U8945 ( .B1(n7166), .B2(n10189), .A(n7165), .ZN(n7167) );
  OAI211_X1 U8946 ( .C1(n9936), .C2(n7169), .A(n7168), .B(n7167), .ZN(P1_U3287) );
  AOI22_X1 U8947 ( .A1(n4415), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10184), .ZN(n7170) );
  OAI21_X1 U8948 ( .B1(n9927), .B2(n9383), .A(n7170), .ZN(n7173) );
  NOR2_X1 U8949 ( .A1(n9936), .A2(n7171), .ZN(n7172) );
  AOI211_X1 U8950 ( .C1(n7174), .C2(n10189), .A(n7173), .B(n7172), .ZN(n7175)
         );
  OAI21_X1 U8951 ( .B1(n4415), .B2(n7176), .A(n7175), .ZN(P1_U3292) );
  OAI21_X1 U8952 ( .B1(n7178), .B2(n4516), .A(n7177), .ZN(n7185) );
  NOR2_X1 U8953 ( .A1(n9349), .A2(n7179), .ZN(n7184) );
  NAND2_X1 U8954 ( .A1(n9346), .A2(n7180), .ZN(n7181) );
  OAI211_X1 U8955 ( .C1(n9283), .C2(n7380), .A(n7182), .B(n7181), .ZN(n7183)
         );
  AOI211_X1 U8956 ( .C1(n7185), .C2(n9329), .A(n7184), .B(n7183), .ZN(n7186)
         );
  INV_X1 U8957 ( .A(n7186), .ZN(P1_U3227) );
  NOR2_X1 U8958 ( .A1(n7188), .A2(n7187), .ZN(n7308) );
  MUX2_X1 U8959 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8376), .Z(n7189) );
  OR2_X1 U8960 ( .A1(n7189), .A2(n7313), .ZN(n7307) );
  AND2_X1 U8961 ( .A1(n7189), .A2(n7313), .ZN(n7309) );
  INV_X1 U8962 ( .A(n7309), .ZN(n7190) );
  NAND2_X1 U8963 ( .A1(n7307), .A2(n7190), .ZN(n7191) );
  XNOR2_X1 U8964 ( .A(n7308), .B(n7191), .ZN(n7208) );
  INV_X1 U8965 ( .A(n7192), .ZN(n7194) );
  NAND2_X1 U8966 ( .A1(n7195), .A2(n7313), .ZN(n7303) );
  OAI21_X1 U8967 ( .B1(n7195), .B2(n7313), .A(n7303), .ZN(n7196) );
  INV_X1 U8968 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7762) );
  AOI21_X1 U8969 ( .B1(n7196), .B2(n7762), .A(n7305), .ZN(n7197) );
  NOR2_X1 U8970 ( .A1(n7197), .A2(n10293), .ZN(n7207) );
  INV_X1 U8971 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8888) );
  INV_X1 U8972 ( .A(n7198), .ZN(n7199) );
  NAND2_X1 U8973 ( .A1(n7200), .A2(n7199), .ZN(n7314) );
  XNOR2_X1 U8974 ( .A(n7314), .B(n7203), .ZN(n7201) );
  OAI21_X1 U8975 ( .B1(n7201), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7316), .ZN(
        n7202) );
  AND2_X1 U8976 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7751) );
  AOI21_X1 U8977 ( .B1(n10233), .B2(n7202), .A(n7751), .ZN(n7205) );
  NAND2_X1 U8978 ( .A1(n10270), .A2(n7203), .ZN(n7204) );
  OAI211_X1 U8979 ( .C1(n8888), .C2(n10283), .A(n7205), .B(n7204), .ZN(n7206)
         );
  AOI211_X1 U8980 ( .C1(n7208), .C2(n10298), .A(n7207), .B(n7206), .ZN(n7209)
         );
  INV_X1 U8981 ( .A(n7209), .ZN(P2_U3191) );
  INV_X1 U8982 ( .A(n7247), .ZN(n7223) );
  NAND2_X1 U8983 ( .A1(n7210), .A2(n8398), .ZN(n7211) );
  AND2_X1 U8984 ( .A1(n7212), .A2(n7211), .ZN(n7216) );
  XNOR2_X1 U8985 ( .A(n8011), .B(n10337), .ZN(n7213) );
  OR2_X1 U8986 ( .A1(n7213), .A2(n8397), .ZN(n7387) );
  NAND2_X1 U8987 ( .A1(n7213), .A2(n8397), .ZN(n7214) );
  AND2_X1 U8988 ( .A1(n7387), .A2(n7214), .ZN(n7215) );
  OAI21_X1 U8989 ( .B1(n7216), .B2(n7215), .A(n7388), .ZN(n7217) );
  NAND2_X1 U8990 ( .A1(n7217), .A2(n8133), .ZN(n7222) );
  INV_X1 U8991 ( .A(n7218), .ZN(n7220) );
  OAI22_X1 U8992 ( .A1(n6284), .A2(n8139), .B1(n8127), .B2(n7490), .ZN(n7219)
         );
  AOI211_X1 U8993 ( .C1(n8119), .C2(n7248), .A(n7220), .B(n7219), .ZN(n7221)
         );
  OAI211_X1 U8994 ( .C1(n7223), .C2(n7495), .A(n7222), .B(n7221), .ZN(P2_U3170) );
  OAI21_X1 U8995 ( .B1(n7225), .B2(n7227), .A(n7224), .ZN(n10326) );
  INV_X1 U8996 ( .A(n10326), .ZN(n7238) );
  OAI22_X1 U8997 ( .A1(n6284), .A2(n8678), .B1(n6899), .B2(n8676), .ZN(n7231)
         );
  NAND3_X1 U8998 ( .A1(n7129), .A2(n7227), .A3(n7226), .ZN(n7228) );
  AOI21_X1 U8999 ( .B1(n7229), .B2(n7228), .A(n8673), .ZN(n7230) );
  AOI211_X1 U9000 ( .C1(n7775), .C2(n10326), .A(n7231), .B(n7230), .ZN(n10328)
         );
  INV_X1 U9001 ( .A(n10328), .ZN(n7234) );
  OAI22_X1 U9002 ( .A1(n7232), .A2(n8731), .B1(n9027), .B2(n8606), .ZN(n7233)
         );
  NOR2_X1 U9003 ( .A1(n7234), .A2(n7233), .ZN(n7235) );
  MUX2_X1 U9004 ( .A(n6697), .B(n7235), .S(n10317), .Z(n7236) );
  OAI21_X1 U9005 ( .B1(n7238), .B2(n7237), .A(n7236), .ZN(P2_U3231) );
  INV_X1 U9006 ( .A(n7239), .ZN(n7240) );
  OR2_X1 U9007 ( .A1(n7775), .A2(n7240), .ZN(n10308) );
  AND2_X1 U9008 ( .A1(n7371), .A2(n8199), .ZN(n8184) );
  XNOR2_X1 U9009 ( .A(n7241), .B(n8341), .ZN(n10336) );
  XNOR2_X1 U9010 ( .A(n7242), .B(n8341), .ZN(n7243) );
  NAND2_X1 U9011 ( .A1(n7243), .A2(n8722), .ZN(n7245) );
  AOI22_X1 U9012 ( .A1(n8719), .A2(n8398), .B1(n8396), .B2(n8717), .ZN(n7244)
         );
  AND2_X1 U9013 ( .A1(n7245), .A2(n7244), .ZN(n10340) );
  INV_X1 U9014 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7246) );
  MUX2_X1 U9015 ( .A(n10340), .B(n7246), .S(n8741), .Z(n7250) );
  AOI22_X1 U9016 ( .A1(n10312), .A2(n7248), .B1(n10314), .B2(n7247), .ZN(n7249) );
  OAI211_X1 U9017 ( .C1(n8728), .C2(n10336), .A(n7250), .B(n7249), .ZN(
        P2_U3229) );
  INV_X1 U9018 ( .A(n8345), .ZN(n7251) );
  NAND3_X1 U9019 ( .A1(n7224), .A2(n8177), .A3(n7251), .ZN(n7252) );
  AND2_X1 U9020 ( .A1(n7253), .A2(n7252), .ZN(n10332) );
  XOR2_X1 U9021 ( .A(n7254), .B(n8345), .Z(n7255) );
  AOI222_X1 U9022 ( .A1(n8722), .A2(n7255), .B1(n8397), .B2(n8717), .C1(n8400), 
        .C2(n8719), .ZN(n10330) );
  MUX2_X1 U9023 ( .A(n9025), .B(n10330), .S(n10317), .Z(n7259) );
  AOI22_X1 U9024 ( .A1(n10312), .A2(n7257), .B1(n10314), .B2(n7256), .ZN(n7258) );
  OAI211_X1 U9025 ( .C1(n10332), .C2(n8728), .A(n7259), .B(n7258), .ZN(
        P2_U3230) );
  OAI21_X1 U9026 ( .B1(n7261), .B2(n9444), .A(n7260), .ZN(n7271) );
  INV_X1 U9027 ( .A(n7271), .ZN(n10209) );
  OR2_X1 U9028 ( .A1(n7452), .A2(n9301), .ZN(n7263) );
  NAND2_X1 U9029 ( .A1(n9642), .A2(n9320), .ZN(n7262) );
  NAND2_X1 U9030 ( .A1(n7263), .A2(n7262), .ZN(n7438) );
  INV_X1 U9031 ( .A(n7264), .ZN(n7266) );
  OAI21_X1 U9032 ( .B1(n7266), .B2(n7265), .A(n4797), .ZN(n7267) );
  NAND2_X1 U9033 ( .A1(n7267), .A2(n9444), .ZN(n7269) );
  OR2_X1 U9034 ( .A1(n9444), .A2(n9441), .ZN(n9433) );
  OR2_X1 U9035 ( .A1(n7268), .A2(n9433), .ZN(n7285) );
  AOI21_X1 U9036 ( .B1(n7269), .B2(n7285), .A(n9906), .ZN(n7270) );
  AOI211_X1 U9037 ( .C1(n7672), .C2(n7271), .A(n7438), .B(n7270), .ZN(n10207)
         );
  MUX2_X1 U9038 ( .A(n7272), .B(n10207), .S(n9916), .Z(n7277) );
  AOI21_X1 U9039 ( .B1(n7273), .B2(n10204), .A(n9922), .ZN(n7274) );
  AND2_X1 U9040 ( .A1(n7291), .A2(n7274), .ZN(n10203) );
  OAI22_X1 U9041 ( .A1(n9927), .A2(n6453), .B1(n9774), .B2(n7439), .ZN(n7275)
         );
  AOI21_X1 U9042 ( .B1(n10203), .B2(n10189), .A(n7275), .ZN(n7276) );
  OAI211_X1 U9043 ( .C1(n10209), .C2(n7297), .A(n7277), .B(n7276), .ZN(
        P1_U3286) );
  OAI21_X1 U9044 ( .B1(n7279), .B2(n7283), .A(n7278), .ZN(n7499) );
  INV_X1 U9045 ( .A(n7499), .ZN(n7298) );
  OR2_X1 U9046 ( .A1(n7280), .A2(n9300), .ZN(n7282) );
  OR2_X1 U9047 ( .A1(n7344), .A2(n9301), .ZN(n7281) );
  NAND2_X1 U9048 ( .A1(n7282), .A2(n7281), .ZN(n7716) );
  INV_X1 U9049 ( .A(n7716), .ZN(n7289) );
  INV_X1 U9050 ( .A(n7283), .ZN(n7287) );
  AND2_X1 U9051 ( .A1(n7285), .A2(n7284), .ZN(n7286) );
  NAND3_X1 U9052 ( .A1(n7285), .A2(n7287), .A3(n7284), .ZN(n7449) );
  OAI211_X1 U9053 ( .C1(n7287), .C2(n7286), .A(n7449), .B(n9931), .ZN(n7288)
         );
  OAI211_X1 U9054 ( .C1(n7298), .C2(n7290), .A(n7289), .B(n7288), .ZN(n7497)
         );
  NAND2_X1 U9055 ( .A1(n7497), .A2(n9916), .ZN(n7296) );
  AOI211_X1 U9056 ( .C1(n7502), .C2(n7291), .A(n9922), .B(n7455), .ZN(n7498)
         );
  INV_X1 U9057 ( .A(n7292), .ZN(n7717) );
  AOI22_X1 U9058 ( .A1(n4415), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7717), .B2(
        n10184), .ZN(n7293) );
  OAI21_X1 U9059 ( .B1(n7720), .B2(n9927), .A(n7293), .ZN(n7294) );
  AOI21_X1 U9060 ( .B1(n7498), .B2(n10189), .A(n7294), .ZN(n7295) );
  OAI211_X1 U9061 ( .C1(n7298), .C2(n7297), .A(n7296), .B(n7295), .ZN(P1_U3285) );
  INV_X1 U9062 ( .A(n7299), .ZN(n7301) );
  OAI222_X1 U9063 ( .A1(n7300), .A2(P1_U3086), .B1(n7911), .B2(n7301), .C1(
        n8975), .C2(n7682), .ZN(P1_U3336) );
  OAI222_X1 U9064 ( .A1(n9171), .A2(n7302), .B1(n9169), .B2(n7301), .C1(n8533), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  INV_X1 U9065 ( .A(n7303), .ZN(n7304) );
  INV_X1 U9066 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U9067 ( .A1(n7551), .A2(P2_REG1_REG_10__SCAN_IN), .B1(n10382), .B2(
        n7555), .ZN(n7306) );
  AOI21_X1 U9068 ( .B1(n4519), .B2(n7306), .A(n7552), .ZN(n7329) );
  OAI21_X1 U9069 ( .B1(n7309), .B2(n7308), .A(n7307), .ZN(n7311) );
  MUX2_X1 U9070 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8376), .Z(n7556) );
  XNOR2_X1 U9071 ( .A(n7556), .B(n7551), .ZN(n7310) );
  NAND2_X1 U9072 ( .A1(n7310), .A2(n7311), .ZN(n7557) );
  OAI21_X1 U9073 ( .B1(n7311), .B2(n7310), .A(n7557), .ZN(n7312) );
  NAND2_X1 U9074 ( .A1(n7312), .A2(n10298), .ZN(n7328) );
  NAND2_X1 U9075 ( .A1(n7314), .A2(n7313), .ZN(n7315) );
  INV_X1 U9076 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U9077 ( .A1(n7551), .A2(n7317), .ZN(n7318) );
  NAND2_X1 U9078 ( .A1(n7318), .A2(n5038), .ZN(n7320) );
  AOI21_X1 U9079 ( .B1(n7321), .B2(n7320), .A(n7319), .ZN(n7324) );
  INV_X1 U9080 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7322) );
  NOR2_X1 U9081 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7322), .ZN(n7919) );
  INV_X1 U9082 ( .A(n7919), .ZN(n7323) );
  OAI21_X1 U9083 ( .B1(n10302), .B2(n7324), .A(n7323), .ZN(n7326) );
  INV_X1 U9084 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n10416) );
  NOR2_X1 U9085 ( .A1(n10283), .A2(n10416), .ZN(n7325) );
  AOI211_X1 U9086 ( .C1(n10270), .C2(n7551), .A(n7326), .B(n7325), .ZN(n7327)
         );
  OAI211_X1 U9087 ( .C1(n7329), .C2(n10293), .A(n7328), .B(n7327), .ZN(
        P2_U3192) );
  INV_X1 U9088 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7330) );
  OAI22_X1 U9089 ( .A1(n10067), .A2(n7331), .B1(n10220), .B2(n7330), .ZN(n7332) );
  INV_X1 U9090 ( .A(n7332), .ZN(n7333) );
  OAI21_X1 U9091 ( .B1(n7334), .B2(n10218), .A(n7333), .ZN(P1_U3465) );
  INV_X1 U9092 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7335) );
  OAI22_X1 U9093 ( .A1(n10067), .A2(n7336), .B1(n10220), .B2(n7335), .ZN(n7337) );
  INV_X1 U9094 ( .A(n7337), .ZN(n7338) );
  OAI21_X1 U9095 ( .B1(n7339), .B2(n10218), .A(n7338), .ZN(P1_U3471) );
  NAND2_X1 U9096 ( .A1(n7340), .A2(n9551), .ZN(n7341) );
  NAND2_X1 U9097 ( .A1(n7342), .A2(n7341), .ZN(n7343) );
  NAND2_X1 U9098 ( .A1(n7343), .A2(n9931), .ZN(n7348) );
  OR2_X1 U9099 ( .A1(n7344), .A2(n9300), .ZN(n7346) );
  OR2_X1 U9100 ( .A1(n7506), .A2(n9301), .ZN(n7345) );
  NAND2_X1 U9101 ( .A1(n7346), .A2(n7345), .ZN(n9202) );
  INV_X1 U9102 ( .A(n9202), .ZN(n7347) );
  NAND2_X1 U9103 ( .A1(n7348), .A2(n7347), .ZN(n7423) );
  INV_X1 U9104 ( .A(n7423), .ZN(n7357) );
  OAI21_X1 U9105 ( .B1(n7350), .B2(n9551), .A(n7349), .ZN(n7425) );
  NAND2_X1 U9106 ( .A1(n7425), .A2(n9876), .ZN(n7356) );
  INV_X1 U9107 ( .A(n7351), .ZN(n7454) );
  AOI211_X1 U9108 ( .C1(n7426), .C2(n7454), .A(n9922), .B(n7661), .ZN(n7424)
         );
  NOR2_X1 U9109 ( .A1(n9205), .A2(n9927), .ZN(n7354) );
  OAI22_X1 U9110 ( .A1(n9916), .A2(n7352), .B1(n9199), .B2(n9774), .ZN(n7353)
         );
  AOI211_X1 U9111 ( .C1(n7424), .C2(n10189), .A(n7354), .B(n7353), .ZN(n7355)
         );
  OAI211_X1 U9112 ( .C1(n4415), .C2(n7357), .A(n7356), .B(n7355), .ZN(P1_U3283) );
  OAI22_X1 U9113 ( .A1(n10067), .A2(n6383), .B1(n10220), .B2(n5128), .ZN(n7358) );
  AOI21_X1 U9114 ( .B1(n7359), .B2(n10220), .A(n7358), .ZN(n7360) );
  INV_X1 U9115 ( .A(n7360), .ZN(P1_U3459) );
  OAI22_X1 U9116 ( .A1(n10067), .A2(n9383), .B1(n10220), .B2(n5061), .ZN(n7361) );
  AOI21_X1 U9117 ( .B1(n7362), .B2(n10220), .A(n7361), .ZN(n7363) );
  INV_X1 U9118 ( .A(n7363), .ZN(P1_U3456) );
  INV_X1 U9119 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7364) );
  OAI22_X1 U9120 ( .A1(n10067), .A2(n7365), .B1(n10220), .B2(n7364), .ZN(n7366) );
  AOI21_X1 U9121 ( .B1(n7367), .B2(n10220), .A(n7366), .ZN(n7368) );
  INV_X1 U9122 ( .A(n7368), .ZN(P1_U3462) );
  XNOR2_X1 U9123 ( .A(n7490), .B(n7470), .ZN(n8349) );
  XNOR2_X1 U9124 ( .A(n7369), .B(n8349), .ZN(n7370) );
  OAI222_X1 U9125 ( .A1(n8678), .A2(n7614), .B1(n8676), .B2(n7393), .C1(n8673), 
        .C2(n7370), .ZN(n7464) );
  INV_X1 U9126 ( .A(n7464), .ZN(n7377) );
  NAND2_X1 U9127 ( .A1(n7372), .A2(n7371), .ZN(n7373) );
  XNOR2_X1 U9128 ( .A(n7373), .B(n8349), .ZN(n7465) );
  INV_X1 U9129 ( .A(n8728), .ZN(n8738) );
  AOI22_X1 U9130 ( .A1(n10312), .A2(n7470), .B1(n10314), .B2(n7384), .ZN(n7374) );
  OAI21_X1 U9131 ( .B1(n4709), .B2(n10317), .A(n7374), .ZN(n7375) );
  AOI21_X1 U9132 ( .B1(n7465), .B2(n8738), .A(n7375), .ZN(n7376) );
  OAI21_X1 U9133 ( .B1(n7377), .B2(n8741), .A(n7376), .ZN(P2_U3228) );
  INV_X1 U9134 ( .A(n7378), .ZN(n7432) );
  OAI222_X1 U9135 ( .A1(n9169), .A2(n7432), .B1(P2_U3151), .B2(n8329), .C1(
        n7379), .C2(n9171), .ZN(P2_U3275) );
  OAI22_X1 U9136 ( .A1(n10067), .A2(n7380), .B1(n10220), .B2(n5222), .ZN(n7381) );
  AOI21_X1 U9137 ( .B1(n7382), .B2(n10220), .A(n7381), .ZN(n7383) );
  INV_X1 U9138 ( .A(n7383), .ZN(P1_U3468) );
  INV_X1 U9139 ( .A(n7384), .ZN(n7398) );
  INV_X1 U9140 ( .A(n7388), .ZN(n7386) );
  INV_X1 U9141 ( .A(n7387), .ZN(n7385) );
  XNOR2_X1 U9142 ( .A(n8011), .B(n7467), .ZN(n7483) );
  XNOR2_X1 U9143 ( .A(n7483), .B(n7490), .ZN(n7389) );
  NOR3_X1 U9144 ( .A1(n7386), .A2(n7385), .A3(n7389), .ZN(n7392) );
  NAND2_X1 U9145 ( .A1(n7388), .A2(n7387), .ZN(n7390) );
  NAND2_X1 U9146 ( .A1(n7390), .A2(n7389), .ZN(n7485) );
  INV_X1 U9147 ( .A(n7485), .ZN(n7391) );
  OAI21_X1 U9148 ( .B1(n7392), .B2(n7391), .A(n8133), .ZN(n7397) );
  OAI22_X1 U9149 ( .A1(n7393), .A2(n8139), .B1(n8127), .B2(n7614), .ZN(n7394)
         );
  AOI211_X1 U9150 ( .C1(n8119), .C2(n7470), .A(n7395), .B(n7394), .ZN(n7396)
         );
  OAI211_X1 U9151 ( .C1(n7398), .C2(n7495), .A(n7397), .B(n7396), .ZN(P2_U3167) );
  AOI22_X1 U9152 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n7574), .B1(n7576), .B2(
        n7575), .ZN(n7406) );
  XNOR2_X1 U9153 ( .A(n7407), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10151) );
  INV_X1 U9154 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7401) );
  XNOR2_X1 U9155 ( .A(n10133), .B(n7401), .ZN(n10138) );
  NOR2_X1 U9156 ( .A1(n7408), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7399) );
  NOR2_X1 U9157 ( .A1(n7400), .A2(n7399), .ZN(n10139) );
  NAND2_X1 U9158 ( .A1(n10138), .A2(n10139), .ZN(n10137) );
  OAI21_X1 U9159 ( .B1(n7411), .B2(n7401), .A(n10137), .ZN(n10150) );
  NAND2_X1 U9160 ( .A1(n10151), .A2(n10150), .ZN(n10149) );
  OAI21_X1 U9161 ( .B1(n7407), .B2(n7402), .A(n10149), .ZN(n7403) );
  INV_X1 U9162 ( .A(n7413), .ZN(n10156) );
  NAND2_X1 U9163 ( .A1(n7403), .A2(n10156), .ZN(n7404) );
  XNOR2_X1 U9164 ( .A(n7403), .B(n7413), .ZN(n10161) );
  NAND2_X1 U9165 ( .A1(n10161), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n10160) );
  NAND2_X1 U9166 ( .A1(n7404), .A2(n10160), .ZN(n7405) );
  NOR2_X1 U9167 ( .A1(n7406), .A2(n7405), .ZN(n7573) );
  AOI21_X1 U9168 ( .B1(n7406), .B2(n7405), .A(n7573), .ZN(n7422) );
  NAND2_X1 U9169 ( .A1(n10145), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n7412) );
  AOI22_X1 U9170 ( .A1(n10145), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n5464), .B2(
        n7407), .ZN(n10148) );
  AOI22_X1 U9171 ( .A1(n10133), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7640), .B2(
        n7411), .ZN(n10136) );
  NOR2_X1 U9172 ( .A1(n7408), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7410) );
  NOR2_X1 U9173 ( .A1(n7410), .A2(n7409), .ZN(n10135) );
  NAND2_X1 U9174 ( .A1(n10136), .A2(n10135), .ZN(n10134) );
  OAI21_X1 U9175 ( .B1(n7640), .B2(n7411), .A(n10134), .ZN(n10147) );
  NAND2_X1 U9176 ( .A1(n10148), .A2(n10147), .ZN(n10146) );
  NAND2_X1 U9177 ( .A1(n7412), .A2(n10146), .ZN(n7414) );
  NAND2_X1 U9178 ( .A1(n7414), .A2(n10156), .ZN(n7415) );
  XNOR2_X1 U9179 ( .A(n7414), .B(n7413), .ZN(n10159) );
  NAND2_X1 U9180 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10159), .ZN(n10157) );
  NAND2_X1 U9181 ( .A1(n7415), .A2(n10157), .ZN(n7417) );
  AOI22_X1 U9182 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7576), .B1(n7574), .B2(
        n7861), .ZN(n7416) );
  NAND2_X1 U9183 ( .A1(n7416), .A2(n7417), .ZN(n7577) );
  OAI211_X1 U9184 ( .C1(n7417), .C2(n7416), .A(n10158), .B(n7577), .ZN(n7420)
         );
  NAND2_X1 U9185 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U9186 ( .A1(n10173), .A2(n7576), .ZN(n7419) );
  NAND2_X1 U9187 ( .A1(n10155), .A2(P1_ADDR_REG_16__SCAN_IN), .ZN(n7418) );
  AND4_X1 U9188 ( .A1(n7420), .A2(n9250), .A3(n7419), .A4(n7418), .ZN(n7421)
         );
  OAI21_X1 U9189 ( .B1(n7422), .B2(n9701), .A(n7421), .ZN(P1_U3259) );
  AOI211_X1 U9190 ( .C1(n7425), .C2(n10217), .A(n7424), .B(n7423), .ZN(n7431)
         );
  AOI22_X1 U9191 ( .A1(n7426), .A2(n6494), .B1(n6496), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7427) );
  OAI21_X1 U9192 ( .B1(n7431), .B2(n6496), .A(n7427), .ZN(P1_U3532) );
  INV_X1 U9193 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7428) );
  OAI22_X1 U9194 ( .A1(n9205), .A2(n10067), .B1(n10220), .B2(n7428), .ZN(n7429) );
  INV_X1 U9195 ( .A(n7429), .ZN(n7430) );
  OAI21_X1 U9196 ( .B1(n7431), .B2(n10218), .A(n7430), .ZN(P1_U3483) );
  OAI222_X1 U9197 ( .A1(P1_U3086), .A2(n9605), .B1(n7911), .B2(n7432), .C1(
        n8976), .C2(n7682), .ZN(P1_U3335) );
  INV_X1 U9198 ( .A(n7433), .ZN(n7437) );
  INV_X1 U9199 ( .A(n7434), .ZN(n7435) );
  AOI21_X1 U9200 ( .B1(n7437), .B2(n7436), .A(n7435), .ZN(n7446) );
  NAND2_X1 U9201 ( .A1(n9346), .A2(n7438), .ZN(n7443) );
  INV_X1 U9202 ( .A(n7439), .ZN(n7440) );
  NAND2_X1 U9203 ( .A1(n9337), .A2(n7440), .ZN(n7441) );
  NAND3_X1 U9204 ( .A1(n7443), .A2(n7442), .A3(n7441), .ZN(n7444) );
  AOI21_X1 U9205 ( .B1(n10204), .B2(n9351), .A(n7444), .ZN(n7445) );
  OAI21_X1 U9206 ( .B1(n7446), .B2(n9354), .A(n7445), .ZN(P1_U3213) );
  OAI21_X1 U9207 ( .B1(n7448), .B2(n7451), .A(n7447), .ZN(n10216) );
  INV_X1 U9208 ( .A(n10216), .ZN(n7463) );
  NAND2_X1 U9209 ( .A1(n7449), .A2(n9443), .ZN(n7450) );
  XOR2_X1 U9210 ( .A(n7451), .B(n7450), .Z(n7453) );
  OR2_X1 U9211 ( .A1(n7452), .A2(n9300), .ZN(n7787) );
  OAI21_X1 U9212 ( .B1(n7453), .B2(n9906), .A(n7787), .ZN(n10214) );
  OAI211_X1 U9213 ( .C1(n10213), .C2(n7455), .A(n7454), .B(n9777), .ZN(n7456)
         );
  OR2_X1 U9214 ( .A1(n7665), .A2(n9301), .ZN(n7788) );
  AND2_X1 U9215 ( .A1(n7456), .A2(n7788), .ZN(n10211) );
  OAI22_X1 U9216 ( .A1(n9916), .A2(n7457), .B1(n7785), .B2(n9774), .ZN(n7458)
         );
  AOI21_X1 U9217 ( .B1(n10186), .B2(n7459), .A(n7458), .ZN(n7460) );
  OAI21_X1 U9218 ( .B1(n10211), .B2(n9778), .A(n7460), .ZN(n7461) );
  AOI21_X1 U9219 ( .B1(n10214), .B2(n9916), .A(n7461), .ZN(n7462) );
  OAI21_X1 U9220 ( .B1(n9936), .B2(n7463), .A(n7462), .ZN(P1_U3284) );
  AOI21_X1 U9221 ( .B1(n7465), .B2(n9071), .A(n7464), .ZN(n7472) );
  INV_X1 U9222 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n7466) );
  OAI22_X1 U9223 ( .A1(n7467), .A2(n9147), .B1(n10367), .B2(n7466), .ZN(n7468)
         );
  INV_X1 U9224 ( .A(n7468), .ZN(n7469) );
  OAI21_X1 U9225 ( .B1(n7472), .B2(n10365), .A(n7469), .ZN(P2_U3405) );
  AOI22_X1 U9226 ( .A1(n9084), .A2(n7470), .B1(n6377), .B2(
        P2_REG1_REG_5__SCAN_IN), .ZN(n7471) );
  OAI21_X1 U9227 ( .B1(n7472), .B2(n6377), .A(n7471), .ZN(P2_U3464) );
  XOR2_X1 U9228 ( .A(n7473), .B(n8344), .Z(n10343) );
  INV_X1 U9229 ( .A(n7474), .ZN(n7496) );
  OAI22_X1 U9230 ( .A1(n8699), .A2(n10342), .B1(n7496), .B2(n8606), .ZN(n7475)
         );
  AOI21_X1 U9231 ( .B1(n8741), .B2(P2_REG2_REG_6__SCAN_IN), .A(n7475), .ZN(
        n7482) );
  INV_X1 U9232 ( .A(n8344), .ZN(n7476) );
  XNOR2_X1 U9233 ( .A(n7477), .B(n7476), .ZN(n7478) );
  NAND2_X1 U9234 ( .A1(n7478), .A2(n8722), .ZN(n7480) );
  AOI22_X1 U9235 ( .A1(n8719), .A2(n8396), .B1(n8394), .B2(n8717), .ZN(n7479)
         );
  NAND2_X1 U9236 ( .A1(n7480), .A2(n7479), .ZN(n10344) );
  NAND2_X1 U9237 ( .A1(n10344), .A2(n10317), .ZN(n7481) );
  OAI211_X1 U9238 ( .C1(n10343), .C2(n8728), .A(n7482), .B(n7481), .ZN(
        P2_U3227) );
  OR2_X1 U9239 ( .A1(n7483), .A2(n8396), .ZN(n7484) );
  XNOR2_X1 U9240 ( .A(n8011), .B(n7492), .ZN(n7606) );
  XNOR2_X1 U9241 ( .A(n7606), .B(n7614), .ZN(n7486) );
  AOI21_X1 U9242 ( .B1(n7487), .B2(n7486), .A(n8131), .ZN(n7488) );
  NAND2_X1 U9243 ( .A1(n7488), .A2(n4764), .ZN(n7494) );
  INV_X1 U9244 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7489) );
  NOR2_X1 U9245 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7489), .ZN(n10249) );
  OAI22_X1 U9246 ( .A1(n7490), .A2(n8139), .B1(n8127), .B2(n7734), .ZN(n7491)
         );
  AOI211_X1 U9247 ( .C1(n8119), .C2(n7492), .A(n10249), .B(n7491), .ZN(n7493)
         );
  OAI211_X1 U9248 ( .C1(n7496), .C2(n7495), .A(n7494), .B(n7493), .ZN(P2_U3179) );
  AOI211_X1 U9249 ( .C1(n7674), .C2(n7499), .A(n7498), .B(n7497), .ZN(n7504)
         );
  OAI22_X1 U9250 ( .A1(n7720), .A2(n10067), .B1(n10220), .B2(n5311), .ZN(n7500) );
  INV_X1 U9251 ( .A(n7500), .ZN(n7501) );
  OAI21_X1 U9252 ( .B1(n7504), .B2(n10218), .A(n7501), .ZN(P1_U3477) );
  AOI22_X1 U9253 ( .A1(n6494), .A2(n7502), .B1(n6496), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n7503) );
  OAI21_X1 U9254 ( .B1(n7504), .B2(n6496), .A(n7503), .ZN(P1_U3530) );
  NAND2_X1 U9255 ( .A1(n7669), .A2(n9460), .ZN(n7505) );
  XNOR2_X1 U9256 ( .A(n7505), .B(n9557), .ZN(n7510) );
  OR2_X1 U9257 ( .A1(n7703), .A2(n9301), .ZN(n7508) );
  OR2_X1 U9258 ( .A1(n7506), .A2(n9300), .ZN(n7507) );
  NAND2_X1 U9259 ( .A1(n7508), .A2(n7507), .ZN(n9225) );
  INV_X1 U9260 ( .A(n9225), .ZN(n7509) );
  OAI21_X1 U9261 ( .B1(n7510), .B2(n9906), .A(n7509), .ZN(n7622) );
  INV_X1 U9262 ( .A(n7622), .ZN(n7521) );
  OAI21_X1 U9263 ( .B1(n7513), .B2(n7512), .A(n7511), .ZN(n7624) );
  NAND2_X1 U9264 ( .A1(n7624), .A2(n9876), .ZN(n7520) );
  INV_X1 U9265 ( .A(n7638), .ZN(n7514) );
  AOI211_X1 U9266 ( .C1(n9229), .C2(n7662), .A(n9922), .B(n7514), .ZN(n7623)
         );
  INV_X1 U9267 ( .A(n9229), .ZN(n7515) );
  NOR2_X1 U9268 ( .A1(n7515), .A2(n9927), .ZN(n7518) );
  OAI22_X1 U9269 ( .A1(n9916), .A2(n7516), .B1(n9227), .B2(n9774), .ZN(n7517)
         );
  AOI211_X1 U9270 ( .C1(n7623), .C2(n10189), .A(n7518), .B(n7517), .ZN(n7519)
         );
  OAI211_X1 U9271 ( .C1(n4415), .C2(n7521), .A(n7520), .B(n7519), .ZN(P1_U3281) );
  INV_X1 U9272 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10390) );
  NOR2_X1 U9273 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7522) );
  AOI21_X1 U9274 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7522), .ZN(n10394) );
  INV_X1 U9275 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n10396) );
  INV_X1 U9276 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U9277 ( .A1(n10396), .A2(n10397), .ZN(n10395) );
  NOR2_X1 U9278 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n10400) );
  INV_X1 U9279 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7524) );
  INV_X1 U9280 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7523) );
  AOI22_X1 U9281 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_14__SCAN_IN), 
        .B1(n7524), .B2(n7523), .ZN(n10405) );
  INV_X1 U9282 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n8411) );
  INV_X1 U9283 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U9284 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(P2_ADDR_REG_13__SCAN_IN), 
        .B1(n8411), .B2(n10131), .ZN(n10408) );
  NOR2_X1 U9285 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7525) );
  AOI21_X1 U9286 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7525), .ZN(n10411) );
  NAND2_X1 U9287 ( .A1(n10416), .A2(n10417), .ZN(n10415) );
  INV_X1 U9288 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8770) );
  AOI22_X1 U9289 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_7__SCAN_IN), 
        .B1(n10281), .B2(n8770), .ZN(n10426) );
  NOR2_X1 U9290 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7533) );
  XOR2_X1 U9291 ( .A(n9651), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n10433) );
  NAND2_X1 U9292 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7531) );
  XOR2_X1 U9293 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10431) );
  NAND2_X1 U9294 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7529) );
  AOI21_X1 U9295 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10386) );
  NAND2_X1 U9296 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n7526) );
  NOR2_X1 U9297 ( .A1(n6551), .A2(n7526), .ZN(n10385) );
  NOR2_X1 U9298 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10385), .ZN(n7527) );
  NOR2_X1 U9299 ( .A1(n10386), .A2(n7527), .ZN(n10429) );
  INV_X1 U9300 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n10242) );
  INV_X1 U9301 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n8964) );
  AOI22_X1 U9302 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .B1(n10242), .B2(n8964), .ZN(n10428) );
  NAND2_X1 U9303 ( .A1(n10429), .A2(n10428), .ZN(n7528) );
  NAND2_X1 U9304 ( .A1(n7529), .A2(n7528), .ZN(n10430) );
  NAND2_X1 U9305 ( .A1(n10431), .A2(n10430), .ZN(n7530) );
  NAND2_X1 U9306 ( .A1(n7531), .A2(n7530), .ZN(n10432) );
  NOR2_X1 U9307 ( .A1(n10433), .A2(n10432), .ZN(n7532) );
  NOR2_X1 U9308 ( .A1(n7533), .A2(n7532), .ZN(n7534) );
  NOR2_X1 U9309 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7534), .ZN(n10421) );
  AND2_X1 U9310 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7534), .ZN(n10422) );
  NOR2_X1 U9311 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10422), .ZN(n7535) );
  NOR2_X1 U9312 ( .A1(n10421), .A2(n7535), .ZN(n7536) );
  NAND2_X1 U9313 ( .A1(n7536), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n7538) );
  INV_X1 U9314 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10261) );
  XNOR2_X1 U9315 ( .A(n7536), .B(n10261), .ZN(n10420) );
  NAND2_X1 U9316 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10420), .ZN(n7537) );
  NAND2_X1 U9317 ( .A1(n7538), .A2(n7537), .ZN(n10425) );
  NAND2_X1 U9318 ( .A1(n10426), .A2(n10425), .ZN(n7539) );
  NAND2_X1 U9319 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7540), .ZN(n7542) );
  XOR2_X1 U9320 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7540), .Z(n10427) );
  NAND2_X1 U9321 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10427), .ZN(n7541) );
  NAND2_X1 U9322 ( .A1(n7542), .A2(n7541), .ZN(n7543) );
  NAND2_X1 U9323 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n7543), .ZN(n7545) );
  XOR2_X1 U9324 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7543), .Z(n10424) );
  NAND2_X1 U9325 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10424), .ZN(n7544) );
  NAND2_X1 U9326 ( .A1(n7545), .A2(n7544), .ZN(n10418) );
  AOI22_X1 U9327 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .B1(n10415), .B2(n10418), .ZN(n10414) );
  NAND2_X1 U9328 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7546) );
  OAI21_X1 U9329 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n7546), .ZN(n10413) );
  NOR2_X1 U9330 ( .A1(n10414), .A2(n10413), .ZN(n10412) );
  AOI21_X1 U9331 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n10412), .ZN(n10410) );
  NAND2_X1 U9332 ( .A1(n10411), .A2(n10410), .ZN(n10409) );
  OAI21_X1 U9333 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10409), .ZN(n10407) );
  NAND2_X1 U9334 ( .A1(n10408), .A2(n10407), .ZN(n10406) );
  OAI21_X1 U9335 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n10406), .ZN(n10404) );
  NAND2_X1 U9336 ( .A1(n10405), .A2(n10404), .ZN(n10403) );
  INV_X1 U9337 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n8934) );
  INV_X1 U9338 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8459) );
  OAI22_X1 U9339 ( .A1(n10400), .A2(n10401), .B1(n8934), .B2(n8459), .ZN(
        n10398) );
  AOI22_X1 U9340 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10395), .B2(n10398), .ZN(n10393) );
  NAND2_X1 U9341 ( .A1(n10394), .A2(n10393), .ZN(n10392) );
  OAI21_X1 U9342 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10392), .ZN(n10389) );
  NOR2_X1 U9343 ( .A1(n10390), .A2(n10389), .ZN(n7547) );
  NAND2_X1 U9344 ( .A1(n10390), .A2(n10389), .ZN(n10388) );
  OAI21_X1 U9345 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n7547), .A(n10388), .ZN(
        n7550) );
  XNOR2_X1 U9346 ( .A(n7548), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n7549) );
  XNOR2_X1 U9347 ( .A(n7550), .B(n7549), .ZN(ADD_1068_U4) );
  NAND2_X1 U9348 ( .A1(n7553), .A2(n7830), .ZN(n7819) );
  OAI21_X1 U9349 ( .B1(n7553), .B2(n7830), .A(n7819), .ZN(n7554) );
  INV_X1 U9350 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7809) );
  NOR2_X1 U9351 ( .A1(n7809), .A2(n7554), .ZN(n7820) );
  AOI21_X1 U9352 ( .B1(n7554), .B2(n7809), .A(n7820), .ZN(n7572) );
  MUX2_X1 U9353 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8376), .Z(n7824) );
  XNOR2_X1 U9354 ( .A(n7824), .B(n7562), .ZN(n7560) );
  OR2_X1 U9355 ( .A1(n7556), .A2(n7555), .ZN(n7558) );
  NAND2_X1 U9356 ( .A1(n7558), .A2(n7557), .ZN(n7559) );
  NAND2_X1 U9357 ( .A1(n7560), .A2(n7559), .ZN(n7825) );
  OAI21_X1 U9358 ( .B1(n7560), .B2(n7559), .A(n7825), .ZN(n7570) );
  NOR2_X1 U9359 ( .A1(n10284), .A2(n7830), .ZN(n7569) );
  INV_X1 U9360 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7567) );
  NOR2_X1 U9361 ( .A1(n7563), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7564) );
  OAI21_X1 U9362 ( .B1(n7833), .B2(n7564), .A(n10233), .ZN(n7566) );
  AND2_X1 U9363 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8101) );
  INV_X1 U9364 ( .A(n8101), .ZN(n7565) );
  OAI211_X1 U9365 ( .C1(n10283), .C2(n7567), .A(n7566), .B(n7565), .ZN(n7568)
         );
  AOI211_X1 U9366 ( .C1(n10298), .C2(n7570), .A(n7569), .B(n7568), .ZN(n7571)
         );
  OAI21_X1 U9367 ( .B1(n7572), .B2(n10293), .A(n7571), .ZN(P2_U3193) );
  AOI21_X1 U9368 ( .B1(n7575), .B2(n7574), .A(n7573), .ZN(n9687) );
  INV_X1 U9369 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9688) );
  XNOR2_X1 U9370 ( .A(n9689), .B(n9688), .ZN(n9686) );
  XNOR2_X1 U9371 ( .A(n9687), .B(n9686), .ZN(n7589) );
  NAND2_X1 U9372 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n7576), .ZN(n7578) );
  NAND2_X1 U9373 ( .A1(n7578), .A2(n7577), .ZN(n7581) );
  INV_X1 U9374 ( .A(n9689), .ZN(n7584) );
  NOR2_X1 U9375 ( .A1(n7584), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9696) );
  INV_X1 U9376 ( .A(n9696), .ZN(n7579) );
  OAI21_X1 U9377 ( .B1(n5547), .B2(n9689), .A(n7579), .ZN(n7580) );
  NOR2_X1 U9378 ( .A1(n7580), .A2(n7581), .ZN(n9695) );
  AOI21_X1 U9379 ( .B1(n7581), .B2(n7580), .A(n9695), .ZN(n7587) );
  NOR2_X1 U9380 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7582), .ZN(n7583) );
  AOI21_X1 U9381 ( .B1(n10155), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n7583), .ZN(
        n7586) );
  NAND2_X1 U9382 ( .A1(n10173), .A2(n7584), .ZN(n7585) );
  OAI211_X1 U9383 ( .C1(n7587), .C2(n10182), .A(n7586), .B(n7585), .ZN(n7588)
         );
  AOI21_X1 U9384 ( .B1(n7589), .B2(n10175), .A(n7588), .ZN(n7590) );
  INV_X1 U9385 ( .A(n7590), .ZN(P1_U3260) );
  OR2_X1 U9386 ( .A1(n7592), .A2(n8206), .ZN(n7689) );
  INV_X1 U9387 ( .A(n7689), .ZN(n7591) );
  AOI21_X1 U9388 ( .B1(n8206), .B2(n7592), .A(n7591), .ZN(n7597) );
  NAND2_X1 U9389 ( .A1(n7593), .A2(n8347), .ZN(n7594) );
  OAI22_X1 U9390 ( .A1(n7614), .A2(n8676), .B1(n7750), .B2(n8678), .ZN(n7595)
         );
  AOI21_X1 U9391 ( .B1(n10347), .B2(n7775), .A(n7595), .ZN(n7596) );
  OAI21_X1 U9392 ( .B1(n7597), .B2(n8673), .A(n7596), .ZN(n10351) );
  INV_X1 U9393 ( .A(n10351), .ZN(n7601) );
  AOI22_X1 U9394 ( .A1(n8741), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n10314), .B2(
        n7612), .ZN(n7598) );
  OAI21_X1 U9395 ( .B1(n10348), .B2(n8699), .A(n7598), .ZN(n7599) );
  AOI21_X1 U9396 ( .B1(n10347), .B2(n8548), .A(n7599), .ZN(n7600) );
  OAI21_X1 U9397 ( .B1(n7601), .B2(n8741), .A(n7600), .ZN(P2_U3226) );
  INV_X1 U9398 ( .A(n7602), .ZN(n7605) );
  OAI222_X1 U9399 ( .A1(n9171), .A2(n7604), .B1(P2_U3151), .B2(n7603), .C1(
        n9169), .C2(n7605), .ZN(P2_U3274) );
  OAI222_X1 U9400 ( .A1(n9535), .A2(P1_U3086), .B1(n7682), .B2(n8952), .C1(
        n7911), .C2(n7605), .ZN(P1_U3334) );
  INV_X1 U9401 ( .A(n7606), .ZN(n7607) );
  XNOR2_X1 U9402 ( .A(n8011), .B(n10348), .ZN(n7608) );
  OR2_X1 U9403 ( .A1(n7608), .A2(n8394), .ZN(n7737) );
  NAND2_X1 U9404 ( .A1(n7608), .A2(n8394), .ZN(n7609) );
  AND2_X1 U9405 ( .A1(n7737), .A2(n7609), .ZN(n7610) );
  OAI21_X1 U9406 ( .B1(n7611), .B2(n7610), .A(n7739), .ZN(n7620) );
  NAND2_X1 U9407 ( .A1(n8141), .A2(n7612), .ZN(n7618) );
  AND2_X1 U9408 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n10268) );
  AOI21_X1 U9409 ( .B1(n8137), .B2(n8393), .A(n10268), .ZN(n7617) );
  NAND2_X1 U9410 ( .A1(n8119), .A2(n7613), .ZN(n7616) );
  OR2_X1 U9411 ( .A1(n8139), .A2(n7614), .ZN(n7615) );
  NAND4_X1 U9412 ( .A1(n7618), .A2(n7617), .A3(n7616), .A4(n7615), .ZN(n7619)
         );
  AOI21_X1 U9413 ( .B1(n7620), .B2(n8133), .A(n7619), .ZN(n7621) );
  INV_X1 U9414 ( .A(n7621), .ZN(P2_U3153) );
  AOI211_X1 U9415 ( .C1(n7624), .C2(n10217), .A(n7623), .B(n7622), .ZN(n7629)
         );
  INV_X1 U9416 ( .A(n10067), .ZN(n7675) );
  INV_X1 U9417 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7625) );
  NOR2_X1 U9418 ( .A1(n10220), .A2(n7625), .ZN(n7626) );
  AOI21_X1 U9419 ( .B1(n9229), .B2(n7675), .A(n7626), .ZN(n7627) );
  OAI21_X1 U9420 ( .B1(n7629), .B2(n10218), .A(n7627), .ZN(P1_U3489) );
  AOI22_X1 U9421 ( .A1(n9229), .A2(n6494), .B1(n6496), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7628) );
  OAI21_X1 U9422 ( .B1(n7629), .B2(n6496), .A(n7628), .ZN(P1_U3534) );
  XNOR2_X1 U9423 ( .A(n7630), .B(n7636), .ZN(n7634) );
  OR2_X1 U9424 ( .A1(n7795), .A2(n9301), .ZN(n7632) );
  OR2_X1 U9425 ( .A1(n7666), .A2(n9300), .ZN(n7631) );
  NAND2_X1 U9426 ( .A1(n7632), .A2(n7631), .ZN(n9290) );
  INV_X1 U9427 ( .A(n9290), .ZN(n7633) );
  OAI21_X1 U9428 ( .B1(n7634), .B2(n9906), .A(n7633), .ZN(n7648) );
  INV_X1 U9429 ( .A(n7648), .ZN(n7645) );
  OAI21_X1 U9430 ( .B1(n7637), .B2(n7636), .A(n7635), .ZN(n7650) );
  NAND2_X1 U9431 ( .A1(n7650), .A2(n9876), .ZN(n7644) );
  AOI211_X1 U9432 ( .C1(n9294), .C2(n7638), .A(n9922), .B(n7697), .ZN(n7649)
         );
  NOR2_X1 U9433 ( .A1(n7639), .A2(n9927), .ZN(n7642) );
  OAI22_X1 U9434 ( .A1(n9916), .A2(n7640), .B1(n9292), .B2(n9774), .ZN(n7641)
         );
  AOI211_X1 U9435 ( .C1(n7649), .C2(n10189), .A(n7642), .B(n7641), .ZN(n7643)
         );
  OAI211_X1 U9436 ( .C1(n4415), .C2(n7645), .A(n7644), .B(n7643), .ZN(P1_U3280) );
  INV_X1 U9437 ( .A(n7646), .ZN(n7683) );
  OAI222_X1 U9438 ( .A1(n9169), .A2(n7683), .B1(P2_U3151), .B2(n8163), .C1(
        n7647), .C2(n9171), .ZN(P2_U3273) );
  AOI211_X1 U9439 ( .C1(n7650), .C2(n10217), .A(n7649), .B(n7648), .ZN(n7653)
         );
  AOI22_X1 U9440 ( .A1(n9294), .A2(n7675), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10218), .ZN(n7651) );
  OAI21_X1 U9441 ( .B1(n7653), .B2(n10218), .A(n7651), .ZN(P1_U3492) );
  AOI22_X1 U9442 ( .A1(n9294), .A2(n6494), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n6496), .ZN(n7652) );
  OAI21_X1 U9443 ( .B1(n7653), .B2(n6496), .A(n7652), .ZN(P1_U3535) );
  INV_X1 U9444 ( .A(n7657), .ZN(n7655) );
  NAND2_X1 U9445 ( .A1(n9166), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7654) );
  OAI211_X1 U9446 ( .C1(n7655), .C2(n9169), .A(n8381), .B(n7654), .ZN(P2_U3272) );
  NAND2_X1 U9447 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  OAI211_X1 U9448 ( .C1(n8783), .C2(n7682), .A(n7658), .B(n9617), .ZN(P1_U3332) );
  OAI21_X1 U9449 ( .B1(n7660), .B2(n9555), .A(n7659), .ZN(n10191) );
  INV_X1 U9450 ( .A(n7661), .ZN(n7664) );
  INV_X1 U9451 ( .A(n7662), .ZN(n7663) );
  AOI211_X1 U9452 ( .C1(n10187), .C2(n7664), .A(n9922), .B(n7663), .ZN(n10188)
         );
  OR2_X1 U9453 ( .A1(n7665), .A2(n9300), .ZN(n7668) );
  OR2_X1 U9454 ( .A1(n7666), .A2(n9301), .ZN(n7667) );
  NAND2_X1 U9455 ( .A1(n7668), .A2(n7667), .ZN(n9310) );
  INV_X1 U9456 ( .A(n7669), .ZN(n7670) );
  AOI211_X1 U9457 ( .C1(n9555), .C2(n4506), .A(n9906), .B(n7670), .ZN(n7671)
         );
  AOI211_X1 U9458 ( .C1(n7672), .C2(n10191), .A(n9310), .B(n7671), .ZN(n10194)
         );
  INV_X1 U9459 ( .A(n10194), .ZN(n7673) );
  AOI211_X1 U9460 ( .C1(n7674), .C2(n10191), .A(n10188), .B(n7673), .ZN(n7678)
         );
  AOI22_X1 U9461 ( .A1(n10187), .A2(n7675), .B1(n10218), .B2(
        P1_REG0_REG_11__SCAN_IN), .ZN(n7676) );
  OAI21_X1 U9462 ( .B1(n7678), .B2(n10218), .A(n7676), .ZN(P1_U3486) );
  AOI22_X1 U9463 ( .A1(n10187), .A2(n6494), .B1(n6496), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n7677) );
  OAI21_X1 U9464 ( .B1(n7678), .B2(n6496), .A(n7677), .ZN(P1_U3533) );
  INV_X1 U9465 ( .A(n7679), .ZN(n7712) );
  AOI22_X1 U9466 ( .A1(n7680), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10082), .ZN(n7681) );
  OAI21_X1 U9467 ( .B1(n7712), .B2(n10085), .A(n7681), .ZN(P1_U3331) );
  OAI222_X1 U9468 ( .A1(P1_U3086), .A2(n5850), .B1(n10085), .B2(n7683), .C1(
        n8977), .C2(n7682), .ZN(P1_U3333) );
  NAND2_X1 U9469 ( .A1(n7684), .A2(n8213), .ZN(n8348) );
  NAND2_X1 U9470 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  XOR2_X1 U9471 ( .A(n8348), .B(n7687), .Z(n10354) );
  NAND2_X1 U9472 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  XOR2_X1 U9473 ( .A(n8348), .B(n7690), .Z(n7691) );
  OAI222_X1 U9474 ( .A1(n8678), .A2(n7773), .B1(n8676), .B2(n7734), .C1(n8673), 
        .C2(n7691), .ZN(n10356) );
  NAND2_X1 U9475 ( .A1(n10356), .A2(n10317), .ZN(n7695) );
  INV_X1 U9476 ( .A(n7729), .ZN(n7692) );
  OAI22_X1 U9477 ( .A1(n10317), .A2(n7055), .B1(n7692), .B2(n8606), .ZN(n7693)
         );
  AOI21_X1 U9478 ( .B1(n10312), .B2(n7743), .A(n7693), .ZN(n7694) );
  OAI211_X1 U9479 ( .C1(n10354), .C2(n8728), .A(n7695), .B(n7694), .ZN(
        P2_U3225) );
  XNOR2_X1 U9480 ( .A(n7696), .B(n9559), .ZN(n10019) );
  AOI211_X1 U9481 ( .C1(n10015), .C2(n4723), .A(n9922), .B(n7800), .ZN(n10014)
         );
  INV_X1 U9482 ( .A(n9182), .ZN(n7698) );
  AOI22_X1 U9483 ( .A1(n4415), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7698), .B2(
        n10184), .ZN(n7699) );
  OAI21_X1 U9484 ( .B1(n7700), .B2(n9927), .A(n7699), .ZN(n7708) );
  NAND3_X1 U9485 ( .A1(n7701), .A2(n9487), .A3(n9469), .ZN(n7702) );
  AOI21_X1 U9486 ( .B1(n7793), .B2(n7702), .A(n9906), .ZN(n7706) );
  OR2_X1 U9487 ( .A1(n7703), .A2(n9300), .ZN(n7705) );
  OR2_X1 U9488 ( .A1(n7853), .A2(n9301), .ZN(n7704) );
  NAND2_X1 U9489 ( .A1(n7705), .A2(n7704), .ZN(n9180) );
  NOR2_X1 U9490 ( .A1(n7706), .A2(n9180), .ZN(n10017) );
  NOR2_X1 U9491 ( .A1(n10017), .A2(n4415), .ZN(n7707) );
  AOI211_X1 U9492 ( .C1(n10014), .C2(n10189), .A(n7708), .B(n7707), .ZN(n7709)
         );
  OAI21_X1 U9493 ( .B1(n9936), .B2(n10019), .A(n7709), .ZN(P1_U3279) );
  OAI222_X1 U9494 ( .A1(n9169), .A2(n7712), .B1(P2_U3151), .B2(n7711), .C1(
        n7710), .C2(n9171), .ZN(P2_U3271) );
  AOI21_X1 U9495 ( .B1(n7715), .B2(n7714), .A(n7713), .ZN(n7723) );
  AND2_X1 U9496 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9676) );
  AOI21_X1 U9497 ( .B1(n9346), .B2(n7716), .A(n9676), .ZN(n7719) );
  NAND2_X1 U9498 ( .A1(n9337), .A2(n7717), .ZN(n7718) );
  OAI211_X1 U9499 ( .C1(n9283), .C2(n7720), .A(n7719), .B(n7718), .ZN(n7721)
         );
  INV_X1 U9500 ( .A(n7721), .ZN(n7722) );
  OAI21_X1 U9501 ( .B1(n7723), .B2(n9354), .A(n7722), .ZN(P1_U3221) );
  INV_X1 U9502 ( .A(n7724), .ZN(n7728) );
  AOI22_X1 U9503 ( .A1(n7725), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10082), .ZN(n7726) );
  OAI21_X1 U9504 ( .B1(n7728), .B2(n10085), .A(n7726), .ZN(P1_U3330) );
  AOI22_X1 U9505 ( .A1(n6352), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9166), .ZN(n7727) );
  OAI21_X1 U9506 ( .B1(n7728), .B2(n9169), .A(n7727), .ZN(P2_U3270) );
  NAND2_X1 U9507 ( .A1(n8141), .A2(n7729), .ZN(n7733) );
  INV_X1 U9508 ( .A(n7730), .ZN(n7731) );
  AOI21_X1 U9509 ( .B1(n8137), .B2(n8392), .A(n7731), .ZN(n7732) );
  OAI211_X1 U9510 ( .C1(n7734), .C2(n8139), .A(n7733), .B(n7732), .ZN(n7742)
         );
  NAND2_X1 U9511 ( .A1(n7739), .A2(n7737), .ZN(n7735) );
  XNOR2_X1 U9512 ( .A(n8011), .B(n7743), .ZN(n7745) );
  XNOR2_X1 U9513 ( .A(n7745), .B(n8393), .ZN(n7736) );
  NAND2_X1 U9514 ( .A1(n7735), .A2(n7736), .ZN(n7747) );
  INV_X1 U9515 ( .A(n7736), .ZN(n7738) );
  NAND3_X1 U9516 ( .A1(n7739), .A2(n7738), .A3(n7737), .ZN(n7740) );
  AOI21_X1 U9517 ( .B1(n7747), .B2(n7740), .A(n8131), .ZN(n7741) );
  AOI211_X1 U9518 ( .C1(n8119), .C2(n7743), .A(n7742), .B(n7741), .ZN(n7744)
         );
  INV_X1 U9519 ( .A(n7744), .ZN(P2_U3161) );
  NAND2_X1 U9520 ( .A1(n7745), .A2(n7750), .ZN(n7746) );
  AND2_X2 U9521 ( .A1(n7747), .A2(n7746), .ZN(n7749) );
  XNOR2_X1 U9522 ( .A(n10313), .B(n8011), .ZN(n7890) );
  XNOR2_X1 U9523 ( .A(n7890), .B(n8392), .ZN(n7748) );
  OAI211_X1 U9524 ( .C1(n7749), .C2(n7748), .A(n7893), .B(n8133), .ZN(n7757)
         );
  OR2_X1 U9525 ( .A1(n8139), .A2(n7750), .ZN(n7753) );
  INV_X1 U9526 ( .A(n7751), .ZN(n7752) );
  OAI211_X1 U9527 ( .C1(n8127), .C2(n7754), .A(n7753), .B(n7752), .ZN(n7755)
         );
  AOI21_X1 U9528 ( .B1(n10315), .B2(n8141), .A(n7755), .ZN(n7756) );
  OAI211_X1 U9529 ( .C1(n7766), .C2(n8145), .A(n7757), .B(n7756), .ZN(P2_U3171) );
  OAI21_X1 U9530 ( .B1(n7759), .B2(n8353), .A(n7758), .ZN(n10310) );
  XOR2_X1 U9531 ( .A(n7760), .B(n8353), .Z(n7761) );
  AOI222_X1 U9532 ( .A1(n8722), .A2(n7761), .B1(n8391), .B2(n8717), .C1(n8393), 
        .C2(n8719), .ZN(n10309) );
  OAI21_X1 U9533 ( .B1(n10353), .B2(n10310), .A(n10309), .ZN(n7768) );
  OAI22_X1 U9534 ( .A1(n9075), .A2(n7766), .B1(n10384), .B2(n7762), .ZN(n7763)
         );
  AOI21_X1 U9535 ( .B1(n7768), .B2(n10384), .A(n7763), .ZN(n7764) );
  INV_X1 U9536 ( .A(n7764), .ZN(P2_U3468) );
  INV_X1 U9537 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7765) );
  OAI22_X1 U9538 ( .A1(n7766), .A2(n9147), .B1(n10367), .B2(n7765), .ZN(n7767)
         );
  AOI21_X1 U9539 ( .B1(n7768), .B2(n10367), .A(n7767), .ZN(n7769) );
  INV_X1 U9540 ( .A(n7769), .ZN(P2_U3417) );
  AND2_X1 U9541 ( .A1(n8222), .A2(n8215), .ZN(n8351) );
  XNOR2_X1 U9542 ( .A(n7770), .B(n8351), .ZN(n7777) );
  INV_X1 U9543 ( .A(n8351), .ZN(n7771) );
  XNOR2_X1 U9544 ( .A(n7772), .B(n7771), .ZN(n10358) );
  OAI22_X1 U9545 ( .A1(n7773), .A2(n8676), .B1(n7922), .B2(n8678), .ZN(n7774)
         );
  AOI21_X1 U9546 ( .B1(n10358), .B2(n7775), .A(n7774), .ZN(n7776) );
  OAI21_X1 U9547 ( .B1(n7777), .B2(n8673), .A(n7776), .ZN(n10364) );
  INV_X1 U9548 ( .A(n10364), .ZN(n7781) );
  INV_X1 U9549 ( .A(n7924), .ZN(n10360) );
  AOI22_X1 U9550 ( .A1(n8741), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10314), .B2(
        n7918), .ZN(n7778) );
  OAI21_X1 U9551 ( .B1(n10360), .B2(n8699), .A(n7778), .ZN(n7779) );
  AOI21_X1 U9552 ( .B1(n10358), .B2(n8548), .A(n7779), .ZN(n7780) );
  OAI21_X1 U9553 ( .B1(n7781), .B2(n8741), .A(n7780), .ZN(P2_U3223) );
  OAI21_X1 U9554 ( .B1(n7783), .B2(n7713), .A(n7782), .ZN(n7784) );
  NAND3_X1 U9555 ( .A1(n4513), .A2(n9329), .A3(n7784), .ZN(n7792) );
  INV_X1 U9556 ( .A(n7785), .ZN(n7790) );
  NOR2_X1 U9557 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7786), .ZN(n10110) );
  AOI21_X1 U9558 ( .B1(n7788), .B2(n7787), .A(n9323), .ZN(n7789) );
  AOI211_X1 U9559 ( .C1(n7790), .C2(n9337), .A(n10110), .B(n7789), .ZN(n7791)
         );
  OAI211_X1 U9560 ( .C1(n10213), .C2(n9283), .A(n7792), .B(n7791), .ZN(
        P1_U3231) );
  NAND2_X1 U9561 ( .A1(n7793), .A2(n9486), .ZN(n7794) );
  XOR2_X1 U9562 ( .A(n9561), .B(n7794), .Z(n7798) );
  OR2_X1 U9563 ( .A1(n7795), .A2(n9300), .ZN(n7797) );
  NAND2_X1 U9564 ( .A1(n9632), .A2(n9321), .ZN(n7796) );
  NAND2_X1 U9565 ( .A1(n7797), .A2(n7796), .ZN(n9345) );
  AOI21_X1 U9566 ( .B1(n7798), .B2(n9931), .A(n9345), .ZN(n7844) );
  XOR2_X1 U9567 ( .A(n7799), .B(n9561), .Z(n7847) );
  NAND2_X1 U9568 ( .A1(n7847), .A2(n9876), .ZN(n7804) );
  OAI22_X1 U9569 ( .A1(n9916), .A2(n8994), .B1(n9348), .B2(n9774), .ZN(n7802)
         );
  OAI211_X1 U9570 ( .C1(n7845), .C2(n7800), .A(n9777), .B(n7859), .ZN(n7843)
         );
  NOR2_X1 U9571 ( .A1(n7843), .A2(n9778), .ZN(n7801) );
  AOI211_X1 U9572 ( .C1(n10186), .C2(n9352), .A(n7802), .B(n7801), .ZN(n7803)
         );
  OAI211_X1 U9573 ( .C1(n4415), .C2(n7844), .A(n7804), .B(n7803), .ZN(P1_U3278) );
  NAND2_X1 U9574 ( .A1(n7805), .A2(n8215), .ZN(n7806) );
  XNOR2_X1 U9575 ( .A(n7806), .B(n7894), .ZN(n7818) );
  XNOR2_X1 U9576 ( .A(n7807), .B(n7894), .ZN(n7808) );
  AOI222_X1 U9577 ( .A1(n8722), .A2(n7808), .B1(n8389), .B2(n8717), .C1(n8391), 
        .C2(n8719), .ZN(n7815) );
  MUX2_X1 U9578 ( .A(n7809), .B(n7815), .S(n10384), .Z(n7811) );
  NAND2_X1 U9579 ( .A1(n8112), .A2(n9084), .ZN(n7810) );
  OAI211_X1 U9580 ( .C1(n9087), .C2(n7818), .A(n7811), .B(n7810), .ZN(P2_U3470) );
  INV_X1 U9581 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7812) );
  MUX2_X1 U9582 ( .A(n7812), .B(n7815), .S(n10367), .Z(n7814) );
  NAND2_X1 U9583 ( .A1(n9158), .A2(n8112), .ZN(n7813) );
  OAI211_X1 U9584 ( .C1(n7818), .C2(n9162), .A(n7814), .B(n7813), .ZN(P2_U3423) );
  INV_X1 U9585 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8955) );
  MUX2_X1 U9586 ( .A(n8955), .B(n7815), .S(n10317), .Z(n7817) );
  AOI22_X1 U9587 ( .A1(n8112), .A2(n10312), .B1(n10314), .B2(n8100), .ZN(n7816) );
  OAI211_X1 U9588 ( .C1(n7818), .C2(n8728), .A(n7817), .B(n7816), .ZN(P2_U3222) );
  INV_X1 U9589 ( .A(n7819), .ZN(n7821) );
  NOR2_X1 U9590 ( .A1(n7821), .A2(n7820), .ZN(n7823) );
  INV_X1 U9591 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7876) );
  AOI22_X1 U9592 ( .A1(n7834), .A2(P2_REG1_REG_12__SCAN_IN), .B1(n7876), .B2(
        n8414), .ZN(n7822) );
  NOR2_X1 U9593 ( .A1(n7823), .A2(n7822), .ZN(n8401) );
  AOI21_X1 U9594 ( .B1(n7823), .B2(n7822), .A(n8401), .ZN(n7842) );
  MUX2_X1 U9595 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8376), .Z(n8415) );
  XNOR2_X1 U9596 ( .A(n8415), .B(n7834), .ZN(n7828) );
  OR2_X1 U9597 ( .A1(n7824), .A2(n7830), .ZN(n7826) );
  NAND2_X1 U9598 ( .A1(n7826), .A2(n7825), .ZN(n7827) );
  NAND2_X1 U9599 ( .A1(n7828), .A2(n7827), .ZN(n8416) );
  OAI21_X1 U9600 ( .B1(n7828), .B2(n7827), .A(n8416), .ZN(n7840) );
  INV_X1 U9601 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n7829) );
  NOR2_X1 U9602 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7829), .ZN(n7965) );
  AND2_X1 U9603 ( .A1(n7831), .A2(n7830), .ZN(n7832) );
  INV_X1 U9604 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9037) );
  XNOR2_X1 U9605 ( .A(n7834), .B(n9037), .ZN(n7835) );
  AOI21_X1 U9606 ( .B1(n4504), .B2(n7835), .A(n8405), .ZN(n7836) );
  NOR2_X1 U9607 ( .A1(n10302), .A2(n7836), .ZN(n7837) );
  AOI211_X1 U9608 ( .C1(n10096), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7965), .B(
        n7837), .ZN(n7838) );
  OAI21_X1 U9609 ( .B1(n8414), .B2(n10284), .A(n7838), .ZN(n7839) );
  AOI21_X1 U9610 ( .B1(n10298), .B2(n7840), .A(n7839), .ZN(n7841) );
  OAI21_X1 U9611 ( .B1(n7842), .B2(n10293), .A(n7841), .ZN(P2_U3194) );
  INV_X1 U9612 ( .A(n10205), .ZN(n10212) );
  OAI211_X1 U9613 ( .C1(n7845), .C2(n10212), .A(n7844), .B(n7843), .ZN(n7846)
         );
  AOI21_X1 U9614 ( .B1(n7847), .B2(n10217), .A(n7846), .ZN(n7850) );
  NAND2_X1 U9615 ( .A1(n10218), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7848) );
  OAI21_X1 U9616 ( .B1(n7850), .B2(n10218), .A(n7848), .ZN(P1_U3498) );
  NAND2_X1 U9617 ( .A1(n6496), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n7849) );
  OAI21_X1 U9618 ( .B1(n7850), .B2(n6496), .A(n7849), .ZN(P1_U3537) );
  OAI211_X1 U9619 ( .C1(n7852), .C2(n9563), .A(n7851), .B(n9931), .ZN(n7856)
         );
  OAI22_X1 U9620 ( .A1(n7854), .A2(n9301), .B1(n7853), .B2(n9300), .ZN(n9248)
         );
  INV_X1 U9621 ( .A(n9248), .ZN(n7855) );
  NAND2_X1 U9622 ( .A1(n7856), .A2(n7855), .ZN(n10010) );
  INV_X1 U9623 ( .A(n10010), .ZN(n7866) );
  NAND2_X1 U9624 ( .A1(n7857), .A2(n9563), .ZN(n10007) );
  NAND3_X1 U9625 ( .A1(n10008), .A2(n10007), .A3(n9876), .ZN(n7865) );
  AOI211_X1 U9626 ( .C1(n10011), .C2(n7859), .A(n9922), .B(n7858), .ZN(n10009)
         );
  INV_X1 U9627 ( .A(n10011), .ZN(n7860) );
  NOR2_X1 U9628 ( .A1(n7860), .A2(n9927), .ZN(n7863) );
  OAI22_X1 U9629 ( .A1(n9916), .A2(n7861), .B1(n9251), .B2(n9774), .ZN(n7862)
         );
  AOI211_X1 U9630 ( .C1(n10009), .C2(n10189), .A(n7863), .B(n7862), .ZN(n7864)
         );
  OAI211_X1 U9631 ( .C1(n4415), .C2(n7866), .A(n7865), .B(n7864), .ZN(P1_U3277) );
  INV_X1 U9632 ( .A(n7867), .ZN(n7872) );
  AOI22_X1 U9633 ( .A1(n7868), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10082), .ZN(n7869) );
  OAI21_X1 U9634 ( .B1(n7872), .B2(n10085), .A(n7869), .ZN(P1_U3329) );
  OAI222_X1 U9635 ( .A1(n9169), .A2(n7872), .B1(P2_U3151), .B2(n7871), .C1(
        n7870), .C2(n9171), .ZN(P2_U3269) );
  XNOR2_X1 U9636 ( .A(n7873), .B(n8231), .ZN(n7884) );
  INV_X1 U9637 ( .A(n8231), .ZN(n8356) );
  XNOR2_X1 U9638 ( .A(n7874), .B(n8356), .ZN(n7875) );
  AOI222_X1 U9639 ( .A1(n8722), .A2(n7875), .B1(n8720), .B2(n8717), .C1(n8390), 
        .C2(n8719), .ZN(n7881) );
  MUX2_X1 U9640 ( .A(n7876), .B(n7881), .S(n10384), .Z(n7878) );
  NAND2_X1 U9641 ( .A1(n7969), .A2(n9084), .ZN(n7877) );
  OAI211_X1 U9642 ( .C1(n7884), .C2(n9087), .A(n7878), .B(n7877), .ZN(P2_U3471) );
  INV_X1 U9643 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n8785) );
  MUX2_X1 U9644 ( .A(n8785), .B(n7881), .S(n10367), .Z(n7880) );
  NAND2_X1 U9645 ( .A1(n9158), .A2(n7969), .ZN(n7879) );
  OAI211_X1 U9646 ( .C1(n7884), .C2(n9162), .A(n7880), .B(n7879), .ZN(P2_U3426) );
  MUX2_X1 U9647 ( .A(n9037), .B(n7881), .S(n10317), .Z(n7883) );
  AOI22_X1 U9648 ( .A1(n7969), .A2(n10312), .B1(n10314), .B2(n7964), .ZN(n7882) );
  OAI211_X1 U9649 ( .C1(n7884), .C2(n8728), .A(n7883), .B(n7882), .ZN(P2_U3221) );
  INV_X1 U9650 ( .A(n7885), .ZN(n7889) );
  AOI22_X1 U9651 ( .A1(n9610), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10082), .ZN(n7886) );
  OAI21_X1 U9652 ( .B1(n7889), .B2(n7911), .A(n7886), .ZN(P1_U3328) );
  AOI21_X1 U9653 ( .B1(n9166), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n7887), .ZN(
        n7888) );
  OAI21_X1 U9654 ( .B1(n7889), .B2(n9169), .A(n7888), .ZN(P2_U3268) );
  XOR2_X1 U9655 ( .A(n8011), .B(n7924), .Z(n7917) );
  INV_X1 U9656 ( .A(n8011), .ZN(n8008) );
  XNOR2_X1 U9657 ( .A(n8352), .B(n8008), .ZN(n8109) );
  INV_X1 U9658 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U9659 ( .A1(n7891), .A2(n8392), .ZN(n7892) );
  NOR3_X1 U9660 ( .A1(n10360), .A2(n8008), .A3(n8391), .ZN(n7895) );
  AOI211_X1 U9661 ( .C1(n7922), .C2(n8008), .A(n7895), .B(n7894), .ZN(n7898)
         );
  NOR3_X1 U9662 ( .A1(n7924), .A2(n8391), .A3(n8011), .ZN(n7896) );
  AOI211_X1 U9663 ( .C1(n7922), .C2(n8011), .A(n7896), .B(n8352), .ZN(n7897)
         );
  XNOR2_X1 U9664 ( .A(n7969), .B(n8011), .ZN(n7899) );
  NAND2_X1 U9665 ( .A1(n7899), .A2(n8104), .ZN(n7960) );
  OAI21_X1 U9666 ( .B1(n7898), .B2(n7897), .A(n7960), .ZN(n7901) );
  INV_X1 U9667 ( .A(n7899), .ZN(n7900) );
  NAND2_X1 U9668 ( .A1(n7900), .A2(n8389), .ZN(n7961) );
  XNOR2_X1 U9669 ( .A(n8732), .B(n8011), .ZN(n7949) );
  XNOR2_X1 U9670 ( .A(n7949), .B(n8235), .ZN(n7902) );
  XNOR2_X1 U9671 ( .A(n7948), .B(n7902), .ZN(n7907) );
  NAND2_X1 U9672 ( .A1(n8141), .A2(n8736), .ZN(n7904) );
  AND2_X1 U9673 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8408) );
  AOI21_X1 U9674 ( .B1(n8137), .B2(n8388), .A(n8408), .ZN(n7903) );
  OAI211_X1 U9675 ( .C1(n8104), .C2(n8139), .A(n7904), .B(n7903), .ZN(n7905)
         );
  AOI21_X1 U9676 ( .B1(n7936), .B2(n8119), .A(n7905), .ZN(n7906) );
  OAI21_X1 U9677 ( .B1(n7907), .B2(n8131), .A(n7906), .ZN(P2_U3174) );
  INV_X1 U9678 ( .A(n7908), .ZN(n7914) );
  AOI22_X1 U9679 ( .A1(n7909), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10082), .ZN(n7910) );
  OAI21_X1 U9680 ( .B1(n7914), .B2(n7911), .A(n7910), .ZN(P1_U3327) );
  AOI21_X1 U9681 ( .B1(n9166), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n7912), .ZN(
        n7913) );
  OAI21_X1 U9682 ( .B1(n7914), .B2(n9169), .A(n7913), .ZN(P2_U3267) );
  XNOR2_X1 U9683 ( .A(n7915), .B(n8391), .ZN(n7916) );
  NOR2_X1 U9684 ( .A1(n7916), .A2(n7917), .ZN(n8106) );
  AOI21_X1 U9685 ( .B1(n7917), .B2(n7916), .A(n8106), .ZN(n7926) );
  NAND2_X1 U9686 ( .A1(n8141), .A2(n7918), .ZN(n7921) );
  INV_X1 U9687 ( .A(n8139), .ZN(n8124) );
  AOI21_X1 U9688 ( .B1(n8124), .B2(n8392), .A(n7919), .ZN(n7920) );
  OAI211_X1 U9689 ( .C1(n7922), .C2(n8127), .A(n7921), .B(n7920), .ZN(n7923)
         );
  AOI21_X1 U9690 ( .B1(n8119), .B2(n7924), .A(n7923), .ZN(n7925) );
  OAI21_X1 U9691 ( .B1(n7926), .B2(n8131), .A(n7925), .ZN(P2_U3157) );
  XNOR2_X1 U9692 ( .A(n7927), .B(n7928), .ZN(n8737) );
  INV_X1 U9693 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8403) );
  INV_X1 U9694 ( .A(n7928), .ZN(n8357) );
  NAND2_X1 U9695 ( .A1(n7931), .A2(n8357), .ZN(n8714) );
  OAI21_X1 U9696 ( .B1(n8357), .B2(n7931), .A(n8714), .ZN(n7932) );
  AOI222_X1 U9697 ( .A1(n8722), .A2(n7932), .B1(n8388), .B2(n8717), .C1(n8389), 
        .C2(n8719), .ZN(n8733) );
  MUX2_X1 U9698 ( .A(n8403), .B(n8733), .S(n10384), .Z(n7934) );
  NAND2_X1 U9699 ( .A1(n7936), .A2(n9084), .ZN(n7933) );
  OAI211_X1 U9700 ( .C1(n9087), .C2(n8737), .A(n7934), .B(n7933), .ZN(P2_U3472) );
  INV_X1 U9701 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7935) );
  MUX2_X1 U9702 ( .A(n7935), .B(n8733), .S(n10367), .Z(n7938) );
  NAND2_X1 U9703 ( .A1(n7936), .A2(n9158), .ZN(n7937) );
  OAI211_X1 U9704 ( .C1(n8737), .C2(n9162), .A(n7938), .B(n7937), .ZN(P2_U3429) );
  XNOR2_X1 U9705 ( .A(n7939), .B(n8339), .ZN(n7975) );
  NAND2_X1 U9706 ( .A1(n7940), .A2(n8339), .ZN(n7941) );
  NAND3_X1 U9707 ( .A1(n7942), .A2(n8722), .A3(n7941), .ZN(n7944) );
  AOI22_X1 U9708 ( .A1(n8691), .A2(n8717), .B1(n8719), .B2(n8388), .ZN(n7943)
         );
  NAND2_X1 U9709 ( .A1(n7944), .A2(n7943), .ZN(n7974) );
  MUX2_X1 U9710 ( .A(n7974), .B(P2_REG2_REG_15__SCAN_IN), .S(n8741), .Z(n7945)
         );
  INV_X1 U9711 ( .A(n7945), .ZN(n7947) );
  AOI22_X1 U9712 ( .A1(n7980), .A2(n10312), .B1(n10314), .B2(n8142), .ZN(n7946) );
  OAI211_X1 U9713 ( .C1(n7975), .C2(n8728), .A(n7947), .B(n7946), .ZN(P2_U3218) );
  XNOR2_X1 U9714 ( .A(n9159), .B(n8011), .ZN(n7978) );
  XNOR2_X1 U9715 ( .A(n7978), .B(n8242), .ZN(n7953) );
  INV_X1 U9716 ( .A(n7949), .ZN(n7951) );
  OAI21_X1 U9717 ( .B1(n7949), .B2(n8720), .A(n7948), .ZN(n7950) );
  OAI21_X1 U9718 ( .B1(n8235), .B2(n7951), .A(n7950), .ZN(n7952) );
  AOI21_X1 U9719 ( .B1(n7953), .B2(n7952), .A(n7979), .ZN(n7959) );
  NAND2_X1 U9720 ( .A1(n8141), .A2(n8723), .ZN(n7956) );
  INV_X1 U9721 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7954) );
  NOR2_X1 U9722 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7954), .ZN(n8434) );
  AOI21_X1 U9723 ( .B1(n8137), .B2(n8718), .A(n8434), .ZN(n7955) );
  OAI211_X1 U9724 ( .C1(n8235), .C2(n8139), .A(n7956), .B(n7955), .ZN(n7957)
         );
  AOI21_X1 U9725 ( .B1(n9159), .B2(n8119), .A(n7957), .ZN(n7958) );
  OAI21_X1 U9726 ( .B1(n7959), .B2(n8131), .A(n7958), .ZN(P2_U3155) );
  NOR2_X1 U9727 ( .A1(n7915), .A2(n8391), .ZN(n8105) );
  NOR3_X1 U9728 ( .A1(n8106), .A2(n8105), .A3(n8109), .ZN(n8107) );
  AOI21_X1 U9729 ( .B1(n8390), .B2(n8109), .A(n8107), .ZN(n7963) );
  NAND2_X1 U9730 ( .A1(n7961), .A2(n7960), .ZN(n7962) );
  XNOR2_X1 U9731 ( .A(n7963), .B(n7962), .ZN(n7971) );
  NAND2_X1 U9732 ( .A1(n8141), .A2(n7964), .ZN(n7967) );
  AOI21_X1 U9733 ( .B1(n8124), .B2(n8390), .A(n7965), .ZN(n7966) );
  OAI211_X1 U9734 ( .C1(n8235), .C2(n8127), .A(n7967), .B(n7966), .ZN(n7968)
         );
  AOI21_X1 U9735 ( .B1(n8119), .B2(n7969), .A(n7968), .ZN(n7970) );
  OAI21_X1 U9736 ( .B1(n7971), .B2(n8131), .A(n7970), .ZN(P2_U3164) );
  MUX2_X1 U9737 ( .A(n7974), .B(P2_REG0_REG_15__SCAN_IN), .S(n10365), .Z(n7973) );
  INV_X1 U9738 ( .A(n7980), .ZN(n8146) );
  OAI22_X1 U9739 ( .A1(n7975), .A2(n9162), .B1(n8146), .B2(n9147), .ZN(n7972)
         );
  OR2_X1 U9740 ( .A1(n7973), .A2(n7972), .ZN(P2_U3435) );
  MUX2_X1 U9741 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n7974), .S(n10384), .Z(n7977) );
  OAI22_X1 U9742 ( .A1(n7975), .A2(n9087), .B1(n8146), .B2(n9075), .ZN(n7976)
         );
  OR2_X1 U9743 ( .A1(n7977), .A2(n7976), .ZN(P2_U3474) );
  XNOR2_X1 U9744 ( .A(n7980), .B(n8011), .ZN(n7982) );
  XNOR2_X1 U9745 ( .A(n7982), .B(n8718), .ZN(n8135) );
  NAND2_X1 U9746 ( .A1(n8136), .A2(n8135), .ZN(n8134) );
  OR2_X1 U9747 ( .A1(n7982), .A2(n7981), .ZN(n7983) );
  XOR2_X1 U9748 ( .A(n8011), .B(n9152), .Z(n8062) );
  INV_X1 U9749 ( .A(n8062), .ZN(n7984) );
  NOR2_X1 U9750 ( .A1(n7984), .A2(n8074), .ZN(n7986) );
  XNOR2_X1 U9751 ( .A(n9076), .B(n8011), .ZN(n7987) );
  XNOR2_X1 U9752 ( .A(n7987), .B(n8707), .ZN(n8070) );
  XNOR2_X1 U9753 ( .A(n8683), .B(n8011), .ZN(n7988) );
  XNOR2_X1 U9754 ( .A(n7988), .B(n8663), .ZN(n8114) );
  INV_X1 U9755 ( .A(n7988), .ZN(n7989) );
  XNOR2_X1 U9756 ( .A(n9139), .B(n8011), .ZN(n7990) );
  XNOR2_X1 U9757 ( .A(n7990), .B(n8677), .ZN(n8040) );
  INV_X1 U9758 ( .A(n7990), .ZN(n7991) );
  XNOR2_X1 U9759 ( .A(n9133), .B(n8011), .ZN(n7992) );
  XNOR2_X1 U9760 ( .A(n7992), .B(n8662), .ZN(n8086) );
  XNOR2_X1 U9761 ( .A(n8052), .B(n8011), .ZN(n7993) );
  XOR2_X1 U9762 ( .A(n8624), .B(n7993), .Z(n8048) );
  XNOR2_X1 U9763 ( .A(n8627), .B(n8011), .ZN(n7995) );
  XNOR2_X1 U9764 ( .A(n7995), .B(n8635), .ZN(n8094) );
  INV_X1 U9765 ( .A(n7995), .ZN(n7996) );
  XNOR2_X1 U9766 ( .A(n9119), .B(n8011), .ZN(n7997) );
  XNOR2_X1 U9767 ( .A(n8083), .B(n8011), .ZN(n8000) );
  XNOR2_X1 U9768 ( .A(n8000), .B(n8615), .ZN(n8079) );
  NAND2_X1 U9769 ( .A1(n8078), .A2(n8079), .ZN(n8002) );
  NAND2_X1 U9770 ( .A1(n8002), .A2(n8001), .ZN(n8055) );
  XNOR2_X1 U9771 ( .A(n8761), .B(n8011), .ZN(n8003) );
  XNOR2_X1 U9772 ( .A(n8003), .B(n8385), .ZN(n8056) );
  NAND2_X1 U9773 ( .A1(n8055), .A2(n8056), .ZN(n8005) );
  NAND2_X1 U9774 ( .A1(n8003), .A2(n8604), .ZN(n8004) );
  NAND2_X1 U9775 ( .A1(n8005), .A2(n8004), .ZN(n8122) );
  XNOR2_X1 U9776 ( .A(n8129), .B(n8011), .ZN(n8006) );
  XNOR2_X1 U9777 ( .A(n8006), .B(n8568), .ZN(n8123) );
  NAND2_X1 U9778 ( .A1(n8006), .A2(n8590), .ZN(n8007) );
  XNOR2_X1 U9779 ( .A(n9103), .B(n8008), .ZN(n8009) );
  NAND2_X1 U9780 ( .A1(n8009), .A2(n8557), .ZN(n8010) );
  OAI21_X1 U9781 ( .B1(n8009), .B2(n8557), .A(n8010), .ZN(n8024) );
  NAND2_X1 U9782 ( .A1(n8025), .A2(n8010), .ZN(n8013) );
  XNOR2_X1 U9783 ( .A(n8553), .B(n8011), .ZN(n8012) );
  XNOR2_X1 U9784 ( .A(n8013), .B(n8012), .ZN(n8020) );
  OAI22_X1 U9785 ( .A1(n8577), .A2(n8139), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8014), .ZN(n8015) );
  INV_X1 U9786 ( .A(n8015), .ZN(n8017) );
  NAND2_X1 U9787 ( .A1(n8562), .A2(n8141), .ZN(n8016) );
  OAI211_X1 U9788 ( .C1(n8384), .C2(n8127), .A(n8017), .B(n8016), .ZN(n8018)
         );
  AOI21_X1 U9789 ( .B1(n9097), .B2(n8119), .A(n8018), .ZN(n8019) );
  OAI21_X1 U9790 ( .B1(n8020), .B2(n8131), .A(n8019), .ZN(P2_U3160) );
  INV_X1 U9791 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n8021) );
  OAI222_X1 U9792 ( .A1(n9169), .A2(n6415), .B1(P2_U3151), .B2(n8022), .C1(
        n8021), .C2(n9171), .ZN(P2_U3266) );
  INV_X1 U9793 ( .A(n9103), .ZN(n8032) );
  AOI21_X1 U9794 ( .B1(n8023), .B2(n8024), .A(n8131), .ZN(n8026) );
  NAND2_X1 U9795 ( .A1(n8026), .A2(n8025), .ZN(n8031) );
  AOI22_X1 U9796 ( .A1(n8568), .A2(n8124), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8027) );
  OAI21_X1 U9797 ( .B1(n8028), .B2(n8127), .A(n8027), .ZN(n8029) );
  AOI21_X1 U9798 ( .B1(n8572), .B2(n8141), .A(n8029), .ZN(n8030) );
  OAI211_X1 U9799 ( .C1(n8032), .C2(n8145), .A(n8031), .B(n8030), .ZN(P2_U3154) );
  XNOR2_X1 U9800 ( .A(n8033), .B(n8623), .ZN(n8039) );
  INV_X1 U9801 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8034) );
  OAI22_X1 U9802 ( .A1(n8139), .A2(n8635), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8034), .ZN(n8036) );
  NOR2_X1 U9803 ( .A1(n8591), .A2(n8127), .ZN(n8035) );
  AOI211_X1 U9804 ( .C1(n8618), .C2(n8141), .A(n8036), .B(n8035), .ZN(n8038)
         );
  NAND2_X1 U9805 ( .A1(n9119), .A2(n8119), .ZN(n8037) );
  OAI211_X1 U9806 ( .C1(n8039), .C2(n8131), .A(n8038), .B(n8037), .ZN(P2_U3156) );
  XOR2_X1 U9807 ( .A(n8041), .B(n8040), .Z(n8046) );
  NAND2_X1 U9808 ( .A1(n8141), .A2(n8668), .ZN(n8043) );
  AOI22_X1 U9809 ( .A1(n8137), .A2(n8387), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8042) );
  OAI211_X1 U9810 ( .C1(n8663), .C2(n8139), .A(n8043), .B(n8042), .ZN(n8044)
         );
  AOI21_X1 U9811 ( .B1(n8669), .B2(n8119), .A(n8044), .ZN(n8045) );
  OAI21_X1 U9812 ( .B1(n8046), .B2(n8131), .A(n8045), .ZN(P2_U3159) );
  XOR2_X1 U9813 ( .A(n8048), .B(n8047), .Z(n8054) );
  NAND2_X1 U9814 ( .A1(n8141), .A2(n8640), .ZN(n8050) );
  AOI22_X1 U9815 ( .A1(n8137), .A2(n8614), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8049) );
  OAI211_X1 U9816 ( .C1(n8662), .C2(n8139), .A(n8050), .B(n8049), .ZN(n8051)
         );
  AOI21_X1 U9817 ( .B1(n8052), .B2(n8119), .A(n8051), .ZN(n8053) );
  OAI21_X1 U9818 ( .B1(n8054), .B2(n8131), .A(n8053), .ZN(P2_U3163) );
  XOR2_X1 U9819 ( .A(n8056), .B(n8055), .Z(n8061) );
  AOI22_X1 U9820 ( .A1(n8568), .A2(n8137), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8058) );
  NAND2_X1 U9821 ( .A1(n8141), .A2(n8592), .ZN(n8057) );
  OAI211_X1 U9822 ( .C1(n8591), .C2(n8139), .A(n8058), .B(n8057), .ZN(n8059)
         );
  AOI21_X1 U9823 ( .B1(n8761), .B2(n8119), .A(n8059), .ZN(n8060) );
  OAI21_X1 U9824 ( .B1(n8061), .B2(n8131), .A(n8060), .ZN(P2_U3165) );
  XNOR2_X1 U9825 ( .A(n8062), .B(n8074), .ZN(n8063) );
  XNOR2_X1 U9826 ( .A(n8064), .B(n8063), .ZN(n8069) );
  NAND2_X1 U9827 ( .A1(n8124), .A2(n8718), .ZN(n8065) );
  NAND2_X1 U9828 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8487) );
  OAI211_X1 U9829 ( .C1(n8675), .C2(n8127), .A(n8065), .B(n8487), .ZN(n8066)
         );
  AOI21_X1 U9830 ( .B1(n8710), .B2(n8141), .A(n8066), .ZN(n8068) );
  NAND2_X1 U9831 ( .A1(n9152), .A2(n8119), .ZN(n8067) );
  OAI211_X1 U9832 ( .C1(n8069), .C2(n8131), .A(n8068), .B(n8067), .ZN(P2_U3166) );
  XOR2_X1 U9833 ( .A(n8071), .B(n8070), .Z(n8077) );
  NAND2_X1 U9834 ( .A1(n8141), .A2(n8697), .ZN(n8073) );
  AOI22_X1 U9835 ( .A1(n8137), .A2(n8692), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8072) );
  OAI211_X1 U9836 ( .C1(n8074), .C2(n8139), .A(n8073), .B(n8072), .ZN(n8075)
         );
  AOI21_X1 U9837 ( .B1(n9076), .B2(n8119), .A(n8075), .ZN(n8076) );
  OAI21_X1 U9838 ( .B1(n8077), .B2(n8131), .A(n8076), .ZN(P2_U3168) );
  XOR2_X1 U9839 ( .A(n8079), .B(n8078), .Z(n8085) );
  AOI22_X1 U9840 ( .A1(n8385), .A2(n8137), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8081) );
  NAND2_X1 U9841 ( .A1(n8141), .A2(n8605), .ZN(n8080) );
  OAI211_X1 U9842 ( .C1(n8623), .C2(n8139), .A(n8081), .B(n8080), .ZN(n8082)
         );
  AOI21_X1 U9843 ( .B1(n8083), .B2(n8119), .A(n8082), .ZN(n8084) );
  OAI21_X1 U9844 ( .B1(n8085), .B2(n8131), .A(n8084), .ZN(P2_U3169) );
  XOR2_X1 U9845 ( .A(n8087), .B(n8086), .Z(n8092) );
  NAND2_X1 U9846 ( .A1(n8141), .A2(n8653), .ZN(n8089) );
  INV_X1 U9847 ( .A(n8624), .ZN(n8650) );
  AOI22_X1 U9848 ( .A1(n8137), .A2(n8650), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8088) );
  OAI211_X1 U9849 ( .C1(n8677), .C2(n8139), .A(n8089), .B(n8088), .ZN(n8090)
         );
  AOI21_X1 U9850 ( .B1(n9133), .B2(n8119), .A(n8090), .ZN(n8091) );
  OAI21_X1 U9851 ( .B1(n8092), .B2(n8131), .A(n8091), .ZN(P2_U3173) );
  XOR2_X1 U9852 ( .A(n8094), .B(n8093), .Z(n8099) );
  NOR2_X1 U9853 ( .A1(n8127), .A2(n8623), .ZN(n8096) );
  OAI22_X1 U9854 ( .A1(n8139), .A2(n8624), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8799), .ZN(n8095) );
  AOI211_X1 U9855 ( .C1(n8628), .C2(n8141), .A(n8096), .B(n8095), .ZN(n8098)
         );
  NAND2_X1 U9856 ( .A1(n8627), .A2(n8119), .ZN(n8097) );
  OAI211_X1 U9857 ( .C1(n8099), .C2(n8131), .A(n8098), .B(n8097), .ZN(P2_U3175) );
  NAND2_X1 U9858 ( .A1(n8141), .A2(n8100), .ZN(n8103) );
  AOI21_X1 U9859 ( .B1(n8124), .B2(n8391), .A(n8101), .ZN(n8102) );
  OAI211_X1 U9860 ( .C1(n8104), .C2(n8127), .A(n8103), .B(n8102), .ZN(n8111)
         );
  OR2_X1 U9861 ( .A1(n8106), .A2(n8105), .ZN(n8108) );
  AOI211_X1 U9862 ( .C1(n8109), .C2(n8108), .A(n8131), .B(n8107), .ZN(n8110)
         );
  AOI211_X1 U9863 ( .C1(n8119), .C2(n8112), .A(n8111), .B(n8110), .ZN(n8113)
         );
  INV_X1 U9864 ( .A(n8113), .ZN(P2_U3176) );
  XOR2_X1 U9865 ( .A(n8115), .B(n8114), .Z(n8121) );
  NAND2_X1 U9866 ( .A1(n8141), .A2(n8684), .ZN(n8117) );
  AOI22_X1 U9867 ( .A1(n8137), .A2(n8649), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3151), .ZN(n8116) );
  OAI211_X1 U9868 ( .C1(n8675), .C2(n8139), .A(n8117), .B(n8116), .ZN(n8118)
         );
  AOI21_X1 U9869 ( .B1(n8683), .B2(n8119), .A(n8118), .ZN(n8120) );
  OAI21_X1 U9870 ( .B1(n8121), .B2(n8131), .A(n8120), .ZN(P2_U3178) );
  XOR2_X1 U9871 ( .A(n8123), .B(n8122), .Z(n8132) );
  AOI22_X1 U9872 ( .A1(n8385), .A2(n8124), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8126) );
  NAND2_X1 U9873 ( .A1(n8141), .A2(n8581), .ZN(n8125) );
  OAI211_X1 U9874 ( .C1(n8577), .C2(n8127), .A(n8126), .B(n8125), .ZN(n8128)
         );
  AOI21_X1 U9875 ( .B1(n8129), .B2(n8119), .A(n8128), .ZN(n8130) );
  OAI21_X1 U9876 ( .B1(n8132), .B2(n8131), .A(n8130), .ZN(P2_U3180) );
  OAI211_X1 U9877 ( .C1(n8136), .C2(n8135), .A(n8134), .B(n8133), .ZN(n8144)
         );
  NAND2_X1 U9878 ( .A1(n8137), .A2(n8691), .ZN(n8138) );
  NAND2_X1 U9879 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8457) );
  OAI211_X1 U9880 ( .C1(n8242), .C2(n8139), .A(n8138), .B(n8457), .ZN(n8140)
         );
  AOI21_X1 U9881 ( .B1(n8142), .B2(n8141), .A(n8140), .ZN(n8143) );
  OAI211_X1 U9882 ( .C1(n8146), .C2(n8145), .A(n8144), .B(n8143), .ZN(P2_U3181) );
  AND2_X1 U9883 ( .A1(n8306), .A2(n8147), .ZN(n8148) );
  MUX2_X1 U9884 ( .A(n8152), .B(n8155), .S(n6332), .Z(n8153) );
  NAND2_X1 U9885 ( .A1(n8626), .A2(n8153), .ZN(n8278) );
  AND2_X1 U9886 ( .A1(n8155), .A2(n8154), .ZN(n8157) );
  OAI211_X1 U9887 ( .C1(n8278), .C2(n8157), .A(n8156), .B(n8279), .ZN(n8158)
         );
  AND2_X1 U9888 ( .A1(n8637), .A2(n8267), .ZN(n8161) );
  NOR2_X1 U9889 ( .A1(n8647), .A2(n8159), .ZN(n8160) );
  MUX2_X1 U9890 ( .A(n8161), .B(n8160), .S(n8312), .Z(n8274) );
  NAND2_X1 U9891 ( .A1(n8170), .A2(n6332), .ZN(n8175) );
  INV_X1 U9892 ( .A(n8164), .ZN(n8162) );
  OAI21_X1 U9893 ( .B1(n8342), .B2(n8162), .A(n8175), .ZN(n8169) );
  NAND2_X1 U9894 ( .A1(n8164), .A2(n8163), .ZN(n8166) );
  MUX2_X1 U9895 ( .A(n8167), .B(n8166), .S(n8165), .Z(n8168) );
  NAND2_X1 U9896 ( .A1(n8169), .A2(n8168), .ZN(n8174) );
  NOR2_X1 U9897 ( .A1(n8170), .A2(n6332), .ZN(n8172) );
  NOR2_X1 U9898 ( .A1(n8172), .A2(n8171), .ZN(n8173) );
  OAI211_X1 U9899 ( .C1(n8176), .C2(n8175), .A(n8174), .B(n8173), .ZN(n8183)
         );
  NAND2_X1 U9900 ( .A1(n8186), .A2(n8177), .ZN(n8180) );
  NAND2_X1 U9901 ( .A1(n8197), .A2(n8178), .ZN(n8179) );
  MUX2_X1 U9902 ( .A(n8180), .B(n8179), .S(n8285), .Z(n8181) );
  INV_X1 U9903 ( .A(n8181), .ZN(n8182) );
  NAND2_X1 U9904 ( .A1(n8183), .A2(n8182), .ZN(n8185) );
  NAND2_X1 U9905 ( .A1(n8185), .A2(n8184), .ZN(n8201) );
  INV_X1 U9906 ( .A(n8186), .ZN(n8188) );
  OAI21_X1 U9907 ( .B1(n8201), .B2(n8188), .A(n8187), .ZN(n8191) );
  AND2_X1 U9908 ( .A1(n8193), .A2(n8198), .ZN(n8190) );
  AOI21_X1 U9909 ( .B1(n8191), .B2(n8190), .A(n8189), .ZN(n8192) );
  MUX2_X1 U9910 ( .A(n8193), .B(n8192), .S(n8285), .Z(n8207) );
  NAND2_X1 U9911 ( .A1(n8214), .A2(n8213), .ZN(n8210) );
  MUX2_X1 U9912 ( .A(n8194), .B(n8210), .S(n8312), .Z(n8196) );
  NOR2_X1 U9913 ( .A1(n8196), .A2(n8195), .ZN(n8218) );
  INV_X1 U9914 ( .A(n8197), .ZN(n8200) );
  OAI211_X1 U9915 ( .C1(n8201), .C2(n8200), .A(n8199), .B(n8198), .ZN(n8204)
         );
  NAND4_X1 U9916 ( .A1(n8204), .A2(n8312), .A3(n8203), .A4(n8202), .ZN(n8205)
         );
  NAND4_X1 U9917 ( .A1(n8207), .A2(n8218), .A3(n8206), .A4(n8205), .ZN(n8221)
         );
  OAI211_X1 U9918 ( .C1(n8210), .C2(n8209), .A(n8222), .B(n8208), .ZN(n8211)
         );
  INV_X1 U9919 ( .A(n8211), .ZN(n8220) );
  NAND2_X1 U9920 ( .A1(n8213), .A2(n8212), .ZN(n8217) );
  NAND2_X1 U9921 ( .A1(n8215), .A2(n8214), .ZN(n8216) );
  AOI21_X1 U9922 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8219) );
  NAND2_X1 U9923 ( .A1(n8224), .A2(n8225), .ZN(n8230) );
  INV_X1 U9924 ( .A(n8225), .ZN(n8226) );
  AOI21_X1 U9925 ( .B1(n8228), .B2(n8227), .A(n8226), .ZN(n8229) );
  MUX2_X1 U9926 ( .A(n8233), .B(n8232), .S(n8285), .Z(n8234) );
  INV_X1 U9927 ( .A(n8237), .ZN(n8240) );
  MUX2_X1 U9928 ( .A(n8235), .B(n8732), .S(n8285), .Z(n8236) );
  OAI21_X1 U9929 ( .B1(n8240), .B2(n8239), .A(n8238), .ZN(n8241) );
  NAND2_X1 U9930 ( .A1(n8241), .A2(n8727), .ZN(n8246) );
  NAND2_X1 U9931 ( .A1(n9159), .A2(n8242), .ZN(n8243) );
  MUX2_X1 U9932 ( .A(n8244), .B(n8243), .S(n8312), .Z(n8245) );
  NAND3_X1 U9933 ( .A1(n8246), .A2(n8339), .A3(n8245), .ZN(n8258) );
  INV_X1 U9934 ( .A(n8247), .ZN(n8250) );
  INV_X1 U9935 ( .A(n8248), .ZN(n8249) );
  MUX2_X1 U9936 ( .A(n8250), .B(n8249), .S(n8312), .Z(n8251) );
  NOR2_X1 U9937 ( .A1(n8252), .A2(n8251), .ZN(n8257) );
  MUX2_X1 U9938 ( .A(n8254), .B(n8253), .S(n8312), .Z(n8255) );
  NAND2_X1 U9939 ( .A1(n8690), .A2(n8255), .ZN(n8256) );
  AOI21_X1 U9940 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8272) );
  NAND2_X1 U9941 ( .A1(n8259), .A2(n8680), .ZN(n8262) );
  NAND2_X1 U9942 ( .A1(n8263), .A2(n8260), .ZN(n8261) );
  MUX2_X1 U9943 ( .A(n8262), .B(n8261), .S(n8312), .Z(n8271) );
  NAND2_X1 U9944 ( .A1(n8264), .A2(n8263), .ZN(n8266) );
  MUX2_X1 U9945 ( .A(n8266), .B(n8265), .S(n6332), .Z(n8269) );
  INV_X1 U9946 ( .A(n8267), .ZN(n8268) );
  NOR2_X1 U9947 ( .A1(n8269), .A2(n8268), .ZN(n8270) );
  OAI21_X1 U9948 ( .B1(n8272), .B2(n8271), .A(n8270), .ZN(n8273) );
  NAND2_X1 U9949 ( .A1(n8598), .A2(n8276), .ZN(n8277) );
  AND2_X1 U9950 ( .A1(n8364), .A2(n8279), .ZN(n8281) );
  AOI21_X1 U9951 ( .B1(n8284), .B2(n8281), .A(n8280), .ZN(n8287) );
  INV_X1 U9952 ( .A(n8364), .ZN(n8282) );
  AOI21_X1 U9953 ( .B1(n8284), .B2(n8283), .A(n8282), .ZN(n8286) );
  MUX2_X1 U9954 ( .A(n8287), .B(n8286), .S(n8285), .Z(n8288) );
  NAND2_X1 U9955 ( .A1(n8288), .A2(n8587), .ZN(n8292) );
  MUX2_X1 U9956 ( .A(n8290), .B(n8289), .S(n8312), .Z(n8291) );
  MUX2_X1 U9957 ( .A(n8294), .B(n8293), .S(n8285), .Z(n8295) );
  INV_X1 U9958 ( .A(n8296), .ZN(n8298) );
  NAND2_X1 U9959 ( .A1(n8298), .A2(n8297), .ZN(n8299) );
  MUX2_X1 U9960 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n4525), .Z(n8321) );
  XNOR2_X1 U9961 ( .A(n8321), .B(SI_30_), .ZN(n8322) );
  NAND2_X1 U9962 ( .A1(n9408), .A2(n4418), .ZN(n8302) );
  NAND2_X1 U9963 ( .A1(n5963), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U9964 ( .A1(n8302), .A2(n8301), .ZN(n8744) );
  OR2_X1 U9965 ( .A1(n8744), .A2(n8303), .ZN(n8319) );
  OAI211_X1 U9966 ( .C1(n8304), .C2(n9097), .A(n8319), .B(n8334), .ZN(n8305)
         );
  NAND2_X1 U9967 ( .A1(n8305), .A2(n8285), .ZN(n8311) );
  NOR2_X1 U9968 ( .A1(n9094), .A2(n8383), .ZN(n8371) );
  INV_X1 U9969 ( .A(n8306), .ZN(n8307) );
  NOR2_X1 U9970 ( .A1(n8371), .A2(n8307), .ZN(n8330) );
  OAI21_X1 U9971 ( .B1(n8308), .B2(n8569), .A(n8330), .ZN(n8309) );
  NAND2_X1 U9972 ( .A1(n8309), .A2(n8312), .ZN(n8310) );
  NAND2_X1 U9973 ( .A1(n8311), .A2(n8310), .ZN(n8316) );
  MUX2_X1 U9974 ( .A(n8569), .B(n9097), .S(n8312), .Z(n8313) );
  AND2_X1 U9975 ( .A1(n8314), .A2(n8313), .ZN(n8315) );
  INV_X1 U9976 ( .A(n8320), .ZN(n8318) );
  INV_X1 U9977 ( .A(n8371), .ZN(n8317) );
  INV_X1 U9978 ( .A(n8319), .ZN(n8370) );
  OAI22_X1 U9979 ( .A1(n8323), .A2(n8322), .B1(SI_30_), .B2(n8321), .ZN(n8326)
         );
  MUX2_X1 U9980 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n4525), .Z(n8324) );
  INV_X1 U9981 ( .A(SI_31_), .ZN(n8954) );
  XNOR2_X1 U9982 ( .A(n8324), .B(n8954), .ZN(n8325) );
  XNOR2_X1 U9983 ( .A(n8326), .B(n8325), .ZN(n9357) );
  NAND2_X1 U9984 ( .A1(n9357), .A2(n4418), .ZN(n8328) );
  NAND2_X1 U9985 ( .A1(n5963), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8327) );
  NOR2_X1 U9986 ( .A1(n9088), .A2(n8539), .ZN(n8372) );
  INV_X1 U9987 ( .A(n8330), .ZN(n8333) );
  INV_X1 U9988 ( .A(n8372), .ZN(n8331) );
  OAI21_X1 U9989 ( .B1(n9094), .B2(n9088), .A(n8331), .ZN(n8332) );
  INV_X1 U9990 ( .A(n8578), .ZN(n8366) );
  INV_X1 U9991 ( .A(n8587), .ZN(n8588) );
  INV_X1 U9992 ( .A(n8598), .ZN(n8337) );
  NOR2_X1 U9993 ( .A1(n8338), .A2(n8337), .ZN(n8613) );
  INV_X1 U9994 ( .A(n8339), .ZN(n8358) );
  NOR4_X1 U9995 ( .A1(n8342), .A2(n8171), .A3(n8341), .A4(n8340), .ZN(n8346)
         );
  NAND4_X1 U9996 ( .A1(n8346), .A2(n8345), .A3(n8344), .A4(n8343), .ZN(n8350)
         );
  NOR4_X1 U9997 ( .A1(n8350), .A2(n8349), .A3(n8348), .A4(n8347), .ZN(n8354)
         );
  NAND4_X1 U9998 ( .A1(n8354), .A2(n8353), .A3(n8352), .A4(n8351), .ZN(n8355)
         );
  NOR4_X1 U9999 ( .A1(n8358), .A2(n8357), .A3(n8356), .A4(n8355), .ZN(n8359)
         );
  NAND4_X1 U10000 ( .A1(n8690), .A2(n8706), .A3(n8359), .A4(n8727), .ZN(n8360)
         );
  NOR4_X1 U10001 ( .A1(n8647), .A2(n8682), .A3(n8361), .A4(n8360), .ZN(n8362)
         );
  NAND4_X1 U10002 ( .A1(n8613), .A2(n8626), .A3(n8638), .A4(n8362), .ZN(n8365)
         );
  NAND2_X1 U10003 ( .A1(n8364), .A2(n8363), .ZN(n8601) );
  NOR4_X1 U10004 ( .A1(n8366), .A2(n8588), .A3(n8365), .A4(n8601), .ZN(n8367)
         );
  NAND4_X1 U10005 ( .A1(n8368), .A2(n8566), .A3(n8367), .A4(n8553), .ZN(n8369)
         );
  NOR4_X1 U10006 ( .A1(n8372), .A2(n8371), .A3(n8370), .A4(n8369), .ZN(n8373)
         );
  XNOR2_X1 U10007 ( .A(n8374), .B(n8509), .ZN(n8382) );
  NAND3_X1 U10008 ( .A1(n8377), .A2(n8376), .A3(n8375), .ZN(n8378) );
  OAI211_X1 U10009 ( .C1(n8379), .C2(n8381), .A(n8378), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8380) );
  OAI21_X1 U10010 ( .B1(n8382), .B2(n8381), .A(n8380), .ZN(P2_U3296) );
  MUX2_X1 U10011 ( .A(n8383), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8399), .Z(
        P2_U3521) );
  INV_X1 U10012 ( .A(n8384), .ZN(n8556) );
  MUX2_X1 U10013 ( .A(n8556), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8399), .Z(
        P2_U3520) );
  MUX2_X1 U10014 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8569), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8557), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8568), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8385), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10018 ( .A(n8615), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8399), .Z(
        P2_U3515) );
  MUX2_X1 U10019 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8386), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8614), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8650), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8387), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10023 ( .A(n8649), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8399), .Z(
        P2_U3510) );
  MUX2_X1 U10024 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8692), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10025 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8707), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10026 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8691), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U10027 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8718), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10028 ( .A(n8388), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8399), .Z(
        P2_U3505) );
  MUX2_X1 U10029 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8720), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10030 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8389), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U10031 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8390), .S(P2_U3893), .Z(
        P2_U3502) );
  MUX2_X1 U10032 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8391), .S(P2_U3893), .Z(
        P2_U3501) );
  MUX2_X1 U10033 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8392), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10034 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8393), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10035 ( .A(n8394), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8399), .Z(
        P2_U3498) );
  MUX2_X1 U10036 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8395), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10037 ( .A(n8396), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8399), .Z(
        P2_U3496) );
  MUX2_X1 U10038 ( .A(n8397), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8399), .Z(
        P2_U3495) );
  MUX2_X1 U10039 ( .A(n8398), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8399), .Z(
        P2_U3494) );
  MUX2_X1 U10040 ( .A(n8400), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8399), .Z(
        P2_U3493) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n5940), .S(P2_U3893), .Z(
        P2_U3492) );
  AOI21_X1 U10042 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8414), .A(n8401), .ZN(
        n8424) );
  AOI21_X1 U10043 ( .B1(n8403), .B2(n8402), .A(n8425), .ZN(n8423) );
  XNOR2_X1 U10044 ( .A(n8437), .B(n8438), .ZN(n8407) );
  INV_X1 U10045 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8406) );
  NOR2_X1 U10046 ( .A1(n8406), .A2(n8407), .ZN(n8439) );
  AOI21_X1 U10047 ( .B1(n8407), .B2(n8406), .A(n8439), .ZN(n8410) );
  INV_X1 U10048 ( .A(n8408), .ZN(n8409) );
  OAI21_X1 U10049 ( .B1(n10302), .B2(n8410), .A(n8409), .ZN(n8413) );
  NOR2_X1 U10050 ( .A1(n10283), .A2(n8411), .ZN(n8412) );
  AOI211_X1 U10051 ( .C1(n10270), .C2(n8438), .A(n8413), .B(n8412), .ZN(n8422)
         );
  MUX2_X1 U10052 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8376), .Z(n8428) );
  XNOR2_X1 U10053 ( .A(n8428), .B(n8438), .ZN(n8419) );
  OR2_X1 U10054 ( .A1(n8415), .A2(n8414), .ZN(n8417) );
  NAND2_X1 U10055 ( .A1(n8417), .A2(n8416), .ZN(n8418) );
  NAND2_X1 U10056 ( .A1(n8419), .A2(n8418), .ZN(n8430) );
  OAI21_X1 U10057 ( .B1(n8419), .B2(n8418), .A(n8430), .ZN(n8420) );
  NAND2_X1 U10058 ( .A1(n8420), .A2(n10298), .ZN(n8421) );
  OAI211_X1 U10059 ( .C1(n8423), .C2(n10293), .A(n8422), .B(n8421), .ZN(
        P2_U3195) );
  NOR2_X1 U10060 ( .A1(n8438), .A2(n8424), .ZN(n8426) );
  INV_X1 U10061 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9083) );
  AOI22_X1 U10062 ( .A1(n8463), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9083), .B2(
        n8451), .ZN(n8427) );
  AOI21_X1 U10063 ( .B1(n4509), .B2(n8427), .A(n8449), .ZN(n8448) );
  INV_X1 U10064 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n9010) );
  MUX2_X1 U10065 ( .A(n9010), .B(n9083), .S(n8376), .Z(n8462) );
  XNOR2_X1 U10066 ( .A(n8462), .B(n8451), .ZN(n8433) );
  INV_X1 U10067 ( .A(n8428), .ZN(n8429) );
  NAND2_X1 U10068 ( .A1(n8438), .A2(n8429), .ZN(n8431) );
  NAND2_X1 U10069 ( .A1(n8431), .A2(n8430), .ZN(n8432) );
  NAND2_X1 U10070 ( .A1(n8433), .A2(n8432), .ZN(n8464) );
  OAI21_X1 U10071 ( .B1(n8433), .B2(n8432), .A(n8464), .ZN(n8446) );
  NAND2_X1 U10072 ( .A1(n10096), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n8436) );
  INV_X1 U10073 ( .A(n8434), .ZN(n8435) );
  OAI211_X1 U10074 ( .C1(n10284), .C2(n8451), .A(n8436), .B(n8435), .ZN(n8445)
         );
  NOR2_X1 U10075 ( .A1(n8438), .A2(n8437), .ZN(n8440) );
  NOR2_X1 U10076 ( .A1(n8440), .A2(n8439), .ZN(n8442) );
  MUX2_X1 U10077 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n9010), .S(n8463), .Z(n8441) );
  AOI21_X1 U10078 ( .B1(n8442), .B2(n8441), .A(n8453), .ZN(n8443) );
  NOR2_X1 U10079 ( .A1(n8443), .A2(n10302), .ZN(n8444) );
  AOI211_X1 U10080 ( .C1(n10298), .C2(n8446), .A(n8445), .B(n8444), .ZN(n8447)
         );
  OAI21_X1 U10081 ( .B1(n8448), .B2(n10293), .A(n8447), .ZN(P2_U3196) );
  INV_X1 U10082 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8808) );
  AOI21_X1 U10083 ( .B1(n8808), .B2(n8450), .A(n8474), .ZN(n8471) );
  XNOR2_X1 U10084 ( .A(n8490), .B(n8489), .ZN(n8456) );
  INV_X1 U10085 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8455) );
  AOI21_X1 U10086 ( .B1(n8456), .B2(n8455), .A(n8454), .ZN(n8458) );
  OAI21_X1 U10087 ( .B1(n10302), .B2(n8458), .A(n8457), .ZN(n8461) );
  NOR2_X1 U10088 ( .A1(n10283), .A2(n8459), .ZN(n8460) );
  AOI211_X1 U10089 ( .C1(n10270), .C2(n8490), .A(n8461), .B(n8460), .ZN(n8470)
         );
  MUX2_X1 U10090 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8376), .Z(n8482) );
  XNOR2_X1 U10091 ( .A(n8482), .B(n8490), .ZN(n8467) );
  NAND2_X1 U10092 ( .A1(n8463), .A2(n8462), .ZN(n8465) );
  NAND2_X1 U10093 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  NAND2_X1 U10094 ( .A1(n8467), .A2(n8466), .ZN(n8483) );
  OAI21_X1 U10095 ( .B1(n8467), .B2(n8466), .A(n8483), .ZN(n8468) );
  NAND2_X1 U10096 ( .A1(n8468), .A2(n10298), .ZN(n8469) );
  OAI211_X1 U10097 ( .C1(n8471), .C2(n10293), .A(n8470), .B(n8469), .ZN(
        P2_U3197) );
  NOR2_X1 U10098 ( .A1(n8490), .A2(n8472), .ZN(n8473) );
  INV_X1 U10099 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9080) );
  OR2_X1 U10100 ( .A1(n8523), .A2(n9080), .ZN(n8504) );
  NAND2_X1 U10101 ( .A1(n8523), .A2(n9080), .ZN(n8475) );
  NAND2_X1 U10102 ( .A1(n8504), .A2(n8475), .ZN(n8479) );
  INV_X1 U10103 ( .A(n8479), .ZN(n8476) );
  INV_X1 U10104 ( .A(n8505), .ZN(n8478) );
  AOI21_X1 U10105 ( .B1(n8480), .B2(n8479), .A(n8478), .ZN(n8503) );
  MUX2_X1 U10106 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8376), .Z(n8521) );
  XNOR2_X1 U10107 ( .A(n8521), .B(n8523), .ZN(n8486) );
  OR2_X1 U10108 ( .A1(n8482), .A2(n8481), .ZN(n8484) );
  NAND2_X1 U10109 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U10110 ( .A1(n8486), .A2(n8485), .ZN(n8524) );
  OAI21_X1 U10111 ( .B1(n8486), .B2(n8485), .A(n8524), .ZN(n8501) );
  NAND2_X1 U10112 ( .A1(n10270), .A2(n8523), .ZN(n8488) );
  OAI211_X1 U10113 ( .C1(n10396), .C2(n10283), .A(n8488), .B(n8487), .ZN(n8500) );
  OR2_X1 U10114 ( .A1(n8523), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8493) );
  NAND2_X1 U10115 ( .A1(n8523), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8492) );
  AND2_X1 U10116 ( .A1(n8493), .A2(n8492), .ZN(n8496) );
  INV_X1 U10117 ( .A(n8496), .ZN(n8494) );
  INV_X1 U10118 ( .A(n8495), .ZN(n8497) );
  NAND2_X1 U10119 ( .A1(n8497), .A2(n8496), .ZN(n8498) );
  AOI21_X1 U10120 ( .B1(n8512), .B2(n8498), .A(n10302), .ZN(n8499) );
  AOI211_X1 U10121 ( .C1(n10298), .C2(n8501), .A(n8500), .B(n8499), .ZN(n8502)
         );
  OAI21_X1 U10122 ( .B1(n8503), .B2(n10293), .A(n8502), .ZN(P2_U3198) );
  INV_X1 U10123 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n10292) );
  NOR2_X1 U10124 ( .A1(n8527), .A2(n8506), .ZN(n8507) );
  INV_X1 U10125 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9073) );
  AOI22_X1 U10126 ( .A1(n10092), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n9073), 
        .B2(n10101), .ZN(n10095) );
  AOI21_X1 U10127 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n10101), .A(n10094), 
        .ZN(n8508) );
  XNOR2_X1 U10128 ( .A(n8509), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8519) );
  INV_X1 U10129 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8510) );
  MUX2_X1 U10130 ( .A(n8510), .B(P2_REG2_REG_19__SCAN_IN), .S(n8509), .Z(n8520) );
  INV_X1 U10131 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n10289) );
  INV_X1 U10132 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8709) );
  OR2_X1 U10133 ( .A1(n8523), .A2(n8709), .ZN(n8511) );
  XNOR2_X1 U10134 ( .A(n8527), .B(n8513), .ZN(n10288) );
  NOR2_X1 U10135 ( .A1(n8527), .A2(n8513), .ZN(n8514) );
  NAND2_X1 U10136 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n10101), .ZN(n8515) );
  OAI21_X1 U10137 ( .B1(n10101), .B2(P2_REG2_REG_18__SCAN_IN), .A(n8515), .ZN(
        n10098) );
  INV_X1 U10138 ( .A(n8515), .ZN(n8516) );
  XNOR2_X1 U10139 ( .A(n8520), .B(n8517), .ZN(n8518) );
  MUX2_X1 U10140 ( .A(n8520), .B(n8519), .S(n8376), .Z(n8532) );
  MUX2_X1 U10141 ( .A(n10289), .B(n10292), .S(n8376), .Z(n8528) );
  XNOR2_X1 U10142 ( .A(n8528), .B(n10285), .ZN(n10297) );
  INV_X1 U10143 ( .A(n8521), .ZN(n8522) );
  NAND2_X1 U10144 ( .A1(n8523), .A2(n8522), .ZN(n8525) );
  NAND2_X1 U10145 ( .A1(n8525), .A2(n8524), .ZN(n10296) );
  NAND2_X1 U10146 ( .A1(n10297), .A2(n10296), .ZN(n10295) );
  INV_X1 U10147 ( .A(n10295), .ZN(n8526) );
  AOI21_X1 U10148 ( .B1(n8528), .B2(n8527), .A(n8526), .ZN(n8530) );
  MUX2_X1 U10149 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8376), .Z(n8529) );
  NAND2_X1 U10150 ( .A1(n8530), .A2(n8529), .ZN(n10088) );
  NOR2_X1 U10151 ( .A1(n8530), .A2(n8529), .ZN(n10090) );
  AOI21_X1 U10152 ( .B1(n10092), .B2(n10088), .A(n10090), .ZN(n8531) );
  XOR2_X1 U10153 ( .A(n8532), .B(n8531), .Z(n8535) );
  NOR2_X1 U10154 ( .A1(n10284), .A2(n8533), .ZN(n8534) );
  INV_X1 U10155 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U10156 ( .A1(n9088), .A2(n10312), .ZN(n8541) );
  INV_X1 U10157 ( .A(n8537), .ZN(n8538) );
  NOR2_X1 U10158 ( .A1(n8539), .A2(n8538), .ZN(n9089) );
  NOR2_X1 U10159 ( .A1(n8540), .A2(n8606), .ZN(n8544) );
  AOI21_X1 U10160 ( .B1(n9089), .B2(n10317), .A(n8544), .ZN(n8543) );
  OAI211_X1 U10161 ( .C1(n10317), .C2(n8993), .A(n8541), .B(n8543), .ZN(
        P2_U3202) );
  NAND2_X1 U10162 ( .A1(n8741), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8542) );
  OAI211_X1 U10163 ( .C1(n9094), .C2(n8699), .A(n8543), .B(n8542), .ZN(
        P2_U3203) );
  INV_X1 U10164 ( .A(n6376), .ZN(n8546) );
  AOI21_X1 U10165 ( .B1(n8741), .B2(P2_REG2_REG_29__SCAN_IN), .A(n8544), .ZN(
        n8545) );
  OAI21_X1 U10166 ( .B1(n8546), .B2(n8699), .A(n8545), .ZN(n8547) );
  AOI21_X1 U10167 ( .B1(n8549), .B2(n8548), .A(n8547), .ZN(n8550) );
  OAI21_X1 U10168 ( .B1(n8551), .B2(n8741), .A(n8550), .ZN(P2_U3204) );
  XNOR2_X1 U10169 ( .A(n8552), .B(n8553), .ZN(n9100) );
  NAND2_X1 U10170 ( .A1(n8556), .A2(n8717), .ZN(n8559) );
  MUX2_X1 U10171 ( .A(n8830), .B(n9095), .S(n10317), .Z(n8564) );
  AOI22_X1 U10172 ( .A1(n9097), .A2(n10312), .B1(n10314), .B2(n8562), .ZN(
        n8563) );
  OAI211_X1 U10173 ( .C1(n9100), .C2(n8728), .A(n8564), .B(n8563), .ZN(
        P2_U3205) );
  XNOR2_X1 U10174 ( .A(n8565), .B(n8566), .ZN(n9106) );
  XNOR2_X1 U10175 ( .A(n8567), .B(n8566), .ZN(n8570) );
  AOI222_X1 U10176 ( .A1(n8722), .A2(n8570), .B1(n8569), .B2(n8717), .C1(n8568), .C2(n8719), .ZN(n9101) );
  MUX2_X1 U10177 ( .A(n8571), .B(n9101), .S(n10317), .Z(n8574) );
  AOI22_X1 U10178 ( .A1(n9103), .A2(n10312), .B1(n10314), .B2(n8572), .ZN(
        n8573) );
  OAI211_X1 U10179 ( .C1(n9106), .C2(n8728), .A(n8574), .B(n8573), .ZN(
        P2_U3206) );
  XNOR2_X1 U10180 ( .A(n8575), .B(n8578), .ZN(n8576) );
  OAI222_X1 U10181 ( .A1(n8678), .A2(n8577), .B1(n8676), .B2(n8604), .C1(n8673), .C2(n8576), .ZN(n8755) );
  NOR2_X1 U10182 ( .A1(n8579), .A2(n8578), .ZN(n8754) );
  INV_X1 U10183 ( .A(n8756), .ZN(n8580) );
  NOR3_X1 U10184 ( .A1(n8754), .A2(n8580), .A3(n8728), .ZN(n8584) );
  AOI22_X1 U10185 ( .A1(n8741), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8581), .B2(
        n10314), .ZN(n8582) );
  OAI21_X1 U10186 ( .B1(n9110), .B2(n8699), .A(n8582), .ZN(n8583) );
  AOI211_X1 U10187 ( .C1(n8755), .C2(n10317), .A(n8584), .B(n8583), .ZN(n8585)
         );
  INV_X1 U10188 ( .A(n8585), .ZN(P2_U3207) );
  XNOR2_X1 U10189 ( .A(n8586), .B(n8587), .ZN(n9114) );
  XNOR2_X1 U10190 ( .A(n4485), .B(n8588), .ZN(n8589) );
  OAI222_X1 U10191 ( .A1(n8676), .A2(n8591), .B1(n8678), .B2(n8590), .C1(n8673), .C2(n8589), .ZN(n8760) );
  INV_X1 U10192 ( .A(n8761), .ZN(n8594) );
  INV_X1 U10193 ( .A(n8592), .ZN(n8593) );
  OAI22_X1 U10194 ( .A1(n8594), .A2(n8731), .B1(n8593), .B2(n8606), .ZN(n8595)
         );
  OAI21_X1 U10195 ( .B1(n8760), .B2(n8595), .A(n10317), .ZN(n8597) );
  NAND2_X1 U10196 ( .A1(n8741), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8596) );
  OAI211_X1 U10197 ( .C1(n9114), .C2(n8728), .A(n8597), .B(n8596), .ZN(
        P2_U3208) );
  NAND2_X1 U10198 ( .A1(n8599), .A2(n8598), .ZN(n8600) );
  XNOR2_X1 U10199 ( .A(n8600), .B(n8601), .ZN(n8765) );
  XNOR2_X1 U10200 ( .A(n8602), .B(n8601), .ZN(n8603) );
  OAI222_X1 U10201 ( .A1(n8678), .A2(n8604), .B1(n8676), .B2(n8623), .C1(n8603), .C2(n8673), .ZN(n8767) );
  INV_X1 U10202 ( .A(n8605), .ZN(n8607) );
  OAI22_X1 U10203 ( .A1(n8764), .A2(n8731), .B1(n8607), .B2(n8606), .ZN(n8608)
         );
  OAI21_X1 U10204 ( .B1(n8767), .B2(n8608), .A(n10317), .ZN(n8610) );
  NAND2_X1 U10205 ( .A1(n8741), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8609) );
  OAI211_X1 U10206 ( .C1(n8765), .C2(n8728), .A(n8610), .B(n8609), .ZN(
        P2_U3209) );
  XNOR2_X1 U10207 ( .A(n8611), .B(n8613), .ZN(n9122) );
  INV_X1 U10208 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8617) );
  XOR2_X1 U10209 ( .A(n8613), .B(n8612), .Z(n8616) );
  AOI222_X1 U10210 ( .A1(n8722), .A2(n8616), .B1(n8615), .B2(n8717), .C1(n8614), .C2(n8719), .ZN(n9117) );
  MUX2_X1 U10211 ( .A(n8617), .B(n9117), .S(n10317), .Z(n8620) );
  AOI22_X1 U10212 ( .A1(n9119), .A2(n10312), .B1(n10314), .B2(n8618), .ZN(
        n8619) );
  OAI211_X1 U10213 ( .C1(n9122), .C2(n8728), .A(n8620), .B(n8619), .ZN(
        P2_U3210) );
  XOR2_X1 U10214 ( .A(n8621), .B(n8626), .Z(n8622) );
  OAI222_X1 U10215 ( .A1(n8676), .A2(n8624), .B1(n8678), .B2(n8623), .C1(n8673), .C2(n8622), .ZN(n9055) );
  INV_X1 U10216 ( .A(n9055), .ZN(n8632) );
  XOR2_X1 U10217 ( .A(n8625), .B(n8626), .Z(n9056) );
  INV_X1 U10218 ( .A(n8627), .ZN(n9126) );
  AOI22_X1 U10219 ( .A1(n8741), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n10314), 
        .B2(n8628), .ZN(n8629) );
  OAI21_X1 U10220 ( .B1(n9126), .B2(n8699), .A(n8629), .ZN(n8630) );
  AOI21_X1 U10221 ( .B1(n9056), .B2(n8738), .A(n8630), .ZN(n8631) );
  OAI21_X1 U10222 ( .B1(n8632), .B2(n8741), .A(n8631), .ZN(P2_U3211) );
  XNOR2_X1 U10223 ( .A(n8633), .B(n8638), .ZN(n8634) );
  OAI222_X1 U10224 ( .A1(n8678), .A2(n8635), .B1(n8676), .B2(n8662), .C1(n8673), .C2(n8634), .ZN(n9059) );
  INV_X1 U10225 ( .A(n9059), .ZN(n8644) );
  NAND2_X1 U10226 ( .A1(n8636), .A2(n8637), .ZN(n8639) );
  XNOR2_X1 U10227 ( .A(n8639), .B(n8638), .ZN(n9060) );
  AOI22_X1 U10228 ( .A1(n8741), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n10314), 
        .B2(n8640), .ZN(n8641) );
  OAI21_X1 U10229 ( .B1(n9130), .B2(n8699), .A(n8641), .ZN(n8642) );
  AOI21_X1 U10230 ( .B1(n9060), .B2(n8738), .A(n8642), .ZN(n8643) );
  OAI21_X1 U10231 ( .B1(n8644), .B2(n8741), .A(n8643), .ZN(P2_U3212) );
  XNOR2_X1 U10232 ( .A(n8645), .B(n8647), .ZN(n9136) );
  INV_X1 U10233 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8652) );
  OAI21_X1 U10234 ( .B1(n8648), .B2(n8647), .A(n8646), .ZN(n8651) );
  AOI222_X1 U10235 ( .A1(n8722), .A2(n8651), .B1(n8650), .B2(n8717), .C1(n8649), .C2(n8719), .ZN(n9131) );
  MUX2_X1 U10236 ( .A(n8652), .B(n9131), .S(n10317), .Z(n8655) );
  AOI22_X1 U10237 ( .A1(n9133), .A2(n10312), .B1(n10314), .B2(n8653), .ZN(
        n8654) );
  OAI211_X1 U10238 ( .C1(n9136), .C2(n8728), .A(n8655), .B(n8654), .ZN(
        P2_U3213) );
  XNOR2_X1 U10239 ( .A(n8656), .B(n8657), .ZN(n9140) );
  NAND2_X1 U10240 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  NAND2_X1 U10241 ( .A1(n8659), .A2(n8722), .ZN(n8660) );
  OR2_X1 U10242 ( .A1(n8661), .A2(n8660), .ZN(n8666) );
  OAI22_X1 U10243 ( .A1(n8663), .A2(n8676), .B1(n8662), .B2(n8678), .ZN(n8664)
         );
  INV_X1 U10244 ( .A(n8664), .ZN(n8665) );
  NAND2_X1 U10245 ( .A1(n8666), .A2(n8665), .ZN(n9137) );
  MUX2_X1 U10246 ( .A(n9137), .B(P2_REG2_REG_19__SCAN_IN), .S(n8741), .Z(n8667) );
  INV_X1 U10247 ( .A(n8667), .ZN(n8671) );
  AOI22_X1 U10248 ( .A1(n8669), .A2(n10312), .B1(n10314), .B2(n8668), .ZN(
        n8670) );
  OAI211_X1 U10249 ( .C1(n9140), .C2(n8728), .A(n8671), .B(n8670), .ZN(
        P2_U3214) );
  XNOR2_X1 U10250 ( .A(n8672), .B(n8682), .ZN(n8674) );
  OAI222_X1 U10251 ( .A1(n8678), .A2(n8677), .B1(n8676), .B2(n8675), .C1(n8674), .C2(n8673), .ZN(n9070) );
  INV_X1 U10252 ( .A(n9070), .ZN(n8688) );
  NAND2_X1 U10253 ( .A1(n8679), .A2(n8680), .ZN(n8681) );
  AOI21_X1 U10254 ( .B1(n8682), .B2(n8681), .A(n4505), .ZN(n9072) );
  INV_X1 U10255 ( .A(n8683), .ZN(n9148) );
  AOI22_X1 U10256 ( .A1(n8741), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n10314), 
        .B2(n8684), .ZN(n8685) );
  OAI21_X1 U10257 ( .B1(n9148), .B2(n8699), .A(n8685), .ZN(n8686) );
  AOI21_X1 U10258 ( .B1(n9072), .B2(n8738), .A(n8686), .ZN(n8687) );
  OAI21_X1 U10259 ( .B1(n8688), .B2(n8741), .A(n8687), .ZN(P2_U3215) );
  XNOR2_X1 U10260 ( .A(n8689), .B(n8690), .ZN(n8693) );
  AOI222_X1 U10261 ( .A1(n8722), .A2(n8693), .B1(n8692), .B2(n8717), .C1(n8691), .C2(n8719), .ZN(n9078) );
  INV_X1 U10262 ( .A(n8679), .ZN(n8694) );
  AOI21_X1 U10263 ( .B1(n8696), .B2(n8695), .A(n8694), .ZN(n9079) );
  INV_X1 U10264 ( .A(n9079), .ZN(n8702) );
  INV_X1 U10265 ( .A(n9076), .ZN(n8700) );
  AOI22_X1 U10266 ( .A1(n8741), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n10314), 
        .B2(n8697), .ZN(n8698) );
  OAI21_X1 U10267 ( .B1(n8700), .B2(n8699), .A(n8698), .ZN(n8701) );
  AOI21_X1 U10268 ( .B1(n8702), .B2(n8738), .A(n8701), .ZN(n8703) );
  OAI21_X1 U10269 ( .B1(n9078), .B2(n8741), .A(n8703), .ZN(P2_U3216) );
  XNOR2_X1 U10270 ( .A(n8704), .B(n8706), .ZN(n9155) );
  XNOR2_X1 U10271 ( .A(n8705), .B(n8706), .ZN(n8708) );
  AOI222_X1 U10272 ( .A1(n8722), .A2(n8708), .B1(n8707), .B2(n8717), .C1(n8718), .C2(n8719), .ZN(n9150) );
  MUX2_X1 U10273 ( .A(n8709), .B(n9150), .S(n10317), .Z(n8712) );
  AOI22_X1 U10274 ( .A1(n9152), .A2(n10312), .B1(n8710), .B2(n10314), .ZN(
        n8711) );
  OAI211_X1 U10275 ( .C1(n9155), .C2(n8728), .A(n8712), .B(n8711), .ZN(
        P2_U3217) );
  NAND2_X1 U10276 ( .A1(n8714), .A2(n8713), .ZN(n8716) );
  XNOR2_X1 U10277 ( .A(n8716), .B(n8715), .ZN(n8721) );
  AOI222_X1 U10278 ( .A1(n8722), .A2(n8721), .B1(n8720), .B2(n8719), .C1(n8718), .C2(n8717), .ZN(n9156) );
  INV_X1 U10279 ( .A(n8731), .ZN(n8724) );
  AOI22_X1 U10280 ( .A1(n9159), .A2(n8724), .B1(n10314), .B2(n8723), .ZN(n8725) );
  AOI21_X1 U10281 ( .B1(n9156), .B2(n8725), .A(n8741), .ZN(n8730) );
  XNOR2_X1 U10282 ( .A(n8726), .B(n8727), .ZN(n9163) );
  OAI22_X1 U10283 ( .A1(n9163), .A2(n8728), .B1(n9010), .B2(n10317), .ZN(n8729) );
  OR2_X1 U10284 ( .A1(n8730), .A2(n8729), .ZN(P2_U3219) );
  NOR2_X1 U10285 ( .A1(n8732), .A2(n8731), .ZN(n8735) );
  INV_X1 U10286 ( .A(n8733), .ZN(n8734) );
  AOI211_X1 U10287 ( .C1(n10314), .C2(n8736), .A(n8735), .B(n8734), .ZN(n8742)
         );
  INV_X1 U10288 ( .A(n8737), .ZN(n8739) );
  AOI22_X1 U10289 ( .A1(n8739), .A2(n8738), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n8741), .ZN(n8740) );
  OAI21_X1 U10290 ( .B1(n8742), .B2(n8741), .A(n8740), .ZN(P2_U3220) );
  NAND2_X1 U10291 ( .A1(n9088), .A2(n9084), .ZN(n8743) );
  NAND2_X1 U10292 ( .A1(n9089), .A2(n10384), .ZN(n8745) );
  OAI211_X1 U10293 ( .C1(n10384), .C2(n9038), .A(n8743), .B(n8745), .ZN(
        P2_U3490) );
  NAND2_X1 U10294 ( .A1(n8744), .A2(n9084), .ZN(n8746) );
  OAI211_X1 U10295 ( .C1(n10384), .C2(n8747), .A(n8746), .B(n8745), .ZN(
        P2_U3489) );
  INV_X1 U10296 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8748) );
  MUX2_X1 U10297 ( .A(n8748), .B(n9095), .S(n10384), .Z(n8750) );
  NAND2_X1 U10298 ( .A1(n9097), .A2(n9084), .ZN(n8749) );
  OAI211_X1 U10299 ( .C1(n9100), .C2(n9087), .A(n8750), .B(n8749), .ZN(
        P2_U3487) );
  INV_X1 U10300 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8751) );
  MUX2_X1 U10301 ( .A(n8751), .B(n9101), .S(n10384), .Z(n8753) );
  NAND2_X1 U10302 ( .A1(n9103), .A2(n9084), .ZN(n8752) );
  OAI211_X1 U10303 ( .C1(n9106), .C2(n9087), .A(n8753), .B(n8752), .ZN(
        P2_U3486) );
  NOR2_X1 U10304 ( .A1(n8754), .A2(n10353), .ZN(n8757) );
  AOI21_X1 U10305 ( .B1(n8757), .B2(n8756), .A(n8755), .ZN(n9107) );
  MUX2_X1 U10306 ( .A(n8758), .B(n9107), .S(n10384), .Z(n8759) );
  OAI21_X1 U10307 ( .B1(n9110), .B2(n9075), .A(n8759), .ZN(P2_U3485) );
  AOI21_X1 U10308 ( .B1(n10325), .B2(n8761), .A(n8760), .ZN(n9111) );
  MUX2_X1 U10309 ( .A(n8762), .B(n9111), .S(n10384), .Z(n8763) );
  OAI21_X1 U10310 ( .B1(n9114), .B2(n9087), .A(n8763), .ZN(P2_U3484) );
  OAI22_X1 U10311 ( .A1(n8765), .A2(n10353), .B1(n8764), .B2(n10359), .ZN(
        n8766) );
  NOR2_X1 U10312 ( .A1(n8767), .A2(n8766), .ZN(n9116) );
  MUX2_X1 U10313 ( .A(n8768), .B(n9116), .S(n10384), .Z(n9051) );
  AOI22_X1 U10314 ( .A1(n8770), .A2(keyinput84), .B1(n9015), .B2(keyinput67), 
        .ZN(n8769) );
  OAI221_X1 U10315 ( .B1(n8770), .B2(keyinput84), .C1(n9015), .C2(keyinput67), 
        .A(n8769), .ZN(n8780) );
  INV_X1 U10316 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9063) );
  AOI22_X1 U10317 ( .A1(n10376), .A2(keyinput29), .B1(n9063), .B2(keyinput0), 
        .ZN(n8771) );
  OAI221_X1 U10318 ( .B1(n10376), .B2(keyinput29), .C1(n9063), .C2(keyinput0), 
        .A(n8771), .ZN(n8779) );
  AOI22_X1 U10319 ( .A1(n8774), .A2(keyinput22), .B1(keyinput107), .B2(n8773), 
        .ZN(n8772) );
  OAI221_X1 U10320 ( .B1(n8774), .B2(keyinput22), .C1(n8773), .C2(keyinput107), 
        .A(n8772), .ZN(n8778) );
  INV_X1 U10321 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U10322 ( .A1(n8776), .A2(keyinput69), .B1(keyinput96), .B2(n10200), 
        .ZN(n8775) );
  OAI221_X1 U10323 ( .B1(n8776), .B2(keyinput69), .C1(n10200), .C2(keyinput96), 
        .A(n8775), .ZN(n8777) );
  NOR4_X1 U10324 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .ZN(n8793)
         );
  AOI22_X1 U10325 ( .A1(n8783), .A2(keyinput110), .B1(n8782), .B2(keyinput30), 
        .ZN(n8781) );
  OAI221_X1 U10326 ( .B1(n8783), .B2(keyinput110), .C1(n8782), .C2(keyinput30), 
        .A(n8781), .ZN(n8791) );
  AOI22_X1 U10327 ( .A1(n8785), .A2(keyinput125), .B1(n8976), .B2(keyinput41), 
        .ZN(n8784) );
  OAI221_X1 U10328 ( .B1(n8785), .B2(keyinput125), .C1(n8976), .C2(keyinput41), 
        .A(n8784), .ZN(n8790) );
  INV_X1 U10329 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U10330 ( .A1(n10198), .A2(keyinput82), .B1(n10289), .B2(keyinput19), 
        .ZN(n8786) );
  OAI221_X1 U10331 ( .B1(n10198), .B2(keyinput82), .C1(n10289), .C2(keyinput19), .A(n8786), .ZN(n8789) );
  INV_X1 U10332 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10195) );
  AOI22_X1 U10333 ( .A1(n9027), .A2(keyinput3), .B1(keyinput79), .B2(n10195), 
        .ZN(n8787) );
  OAI221_X1 U10334 ( .B1(n9027), .B2(keyinput3), .C1(n10195), .C2(keyinput79), 
        .A(n8787), .ZN(n8788) );
  NOR4_X1 U10335 ( .A1(n8791), .A2(n8790), .A3(n8789), .A4(n8788), .ZN(n8792)
         );
  AND2_X1 U10336 ( .A1(n8793), .A2(n8792), .ZN(n8949) );
  AOI22_X1 U10337 ( .A1(n7256), .A2(keyinput50), .B1(keyinput88), .B2(n10281), 
        .ZN(n8794) );
  OAI221_X1 U10338 ( .B1(n7256), .B2(keyinput50), .C1(n10281), .C2(keyinput88), 
        .A(n8794), .ZN(n8803) );
  INV_X1 U10339 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8796) );
  AOI22_X1 U10340 ( .A1(n8796), .A2(keyinput63), .B1(n9025), .B2(keyinput66), 
        .ZN(n8795) );
  OAI221_X1 U10341 ( .B1(n8796), .B2(keyinput63), .C1(n9025), .C2(keyinput66), 
        .A(n8795), .ZN(n8802) );
  AOI22_X1 U10342 ( .A1(n9948), .A2(keyinput77), .B1(keyinput78), .B2(n10416), 
        .ZN(n8797) );
  OAI221_X1 U10343 ( .B1(n9948), .B2(keyinput77), .C1(n10416), .C2(keyinput78), 
        .A(n8797), .ZN(n8801) );
  AOI22_X1 U10344 ( .A1(n8571), .A2(keyinput23), .B1(n8799), .B2(keyinput53), 
        .ZN(n8798) );
  OAI221_X1 U10345 ( .B1(n8571), .B2(keyinput23), .C1(n8799), .C2(keyinput53), 
        .A(n8798), .ZN(n8800) );
  NOR4_X1 U10346 ( .A1(n8803), .A2(n8802), .A3(n8801), .A4(n8800), .ZN(n8948)
         );
  AOI22_X1 U10347 ( .A1(n9191), .A2(keyinput109), .B1(n8805), .B2(keyinput65), 
        .ZN(n8804) );
  OAI221_X1 U10348 ( .B1(n9191), .B2(keyinput109), .C1(n8805), .C2(keyinput65), 
        .A(n8804), .ZN(n8806) );
  INV_X1 U10349 ( .A(n8806), .ZN(n8817) );
  AOI22_X1 U10350 ( .A1(n10041), .A2(keyinput5), .B1(n8808), .B2(keyinput124), 
        .ZN(n8807) );
  OAI221_X1 U10351 ( .B1(n10041), .B2(keyinput5), .C1(n8808), .C2(keyinput124), 
        .A(n8807), .ZN(n8809) );
  INV_X1 U10352 ( .A(n8809), .ZN(n8816) );
  AOI22_X1 U10353 ( .A1(n9018), .A2(keyinput48), .B1(n8974), .B2(keyinput16), 
        .ZN(n8810) );
  OAI221_X1 U10354 ( .B1(n9018), .B2(keyinput48), .C1(n8974), .C2(keyinput16), 
        .A(n8810), .ZN(n8811) );
  INV_X1 U10355 ( .A(n8811), .ZN(n8815) );
  XNOR2_X1 U10356 ( .A(keyinput104), .B(n10264), .ZN(n8813) );
  XNOR2_X1 U10357 ( .A(keyinput122), .B(n8991), .ZN(n8812) );
  NOR2_X1 U10358 ( .A1(n8813), .A2(n8812), .ZN(n8814) );
  AND4_X1 U10359 ( .A1(n8817), .A2(n8816), .A3(n8815), .A4(n8814), .ZN(n8840)
         );
  AOI22_X1 U10360 ( .A1(n4704), .A2(keyinput34), .B1(n8819), .B2(keyinput127), 
        .ZN(n8818) );
  OAI221_X1 U10361 ( .B1(n4704), .B2(keyinput34), .C1(n8819), .C2(keyinput127), 
        .A(n8818), .ZN(n8823) );
  AOI22_X1 U10362 ( .A1(n8975), .A2(keyinput92), .B1(n8821), .B2(keyinput37), 
        .ZN(n8820) );
  OAI221_X1 U10363 ( .B1(n8975), .B2(keyinput92), .C1(n8821), .C2(keyinput37), 
        .A(n8820), .ZN(n8822) );
  NOR2_X1 U10364 ( .A1(n8823), .A2(n8822), .ZN(n8839) );
  INV_X1 U10365 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U10366 ( .A1(n8993), .A2(keyinput114), .B1(n10199), .B2(keyinput64), 
        .ZN(n8824) );
  OAI221_X1 U10367 ( .B1(n8993), .B2(keyinput114), .C1(n10199), .C2(keyinput64), .A(n8824), .ZN(n8828) );
  INV_X1 U10368 ( .A(SI_4_), .ZN(n8826) );
  AOI22_X1 U10369 ( .A1(n10030), .A2(keyinput119), .B1(n8826), .B2(keyinput115), .ZN(n8825) );
  OAI221_X1 U10370 ( .B1(n10030), .B2(keyinput119), .C1(n8826), .C2(
        keyinput115), .A(n8825), .ZN(n8827) );
  NOR2_X1 U10371 ( .A1(n8828), .A2(n8827), .ZN(n8838) );
  AOI22_X1 U10372 ( .A1(n10380), .A2(keyinput60), .B1(n8830), .B2(keyinput80), 
        .ZN(n8829) );
  OAI221_X1 U10373 ( .B1(n10380), .B2(keyinput60), .C1(n8830), .C2(keyinput80), 
        .A(n8829), .ZN(n8836) );
  XNOR2_X1 U10374 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput12), .ZN(n8834) );
  XNOR2_X1 U10375 ( .A(P2_REG2_REG_15__SCAN_IN), .B(keyinput35), .ZN(n8833) );
  XNOR2_X1 U10376 ( .A(P1_REG1_REG_0__SCAN_IN), .B(keyinput74), .ZN(n8832) );
  XNOR2_X1 U10377 ( .A(keyinput112), .B(P1_ADDR_REG_6__SCAN_IN), .ZN(n8831) );
  NAND4_X1 U10378 ( .A1(n8834), .A2(n8833), .A3(n8832), .A4(n8831), .ZN(n8835)
         );
  NOR2_X1 U10379 ( .A1(n8836), .A2(n8835), .ZN(n8837) );
  NAND4_X1 U10380 ( .A1(n8840), .A2(n8839), .A3(n8838), .A4(n8837), .ZN(n8877)
         );
  XNOR2_X1 U10381 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput100), .ZN(n8844)
         );
  XNOR2_X1 U10382 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput61), .ZN(n8843) );
  XNOR2_X1 U10383 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput86), .ZN(n8842) );
  XNOR2_X1 U10384 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput38), .ZN(n8841) );
  NAND4_X1 U10385 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(n8850)
         );
  XNOR2_X1 U10386 ( .A(SI_21_), .B(keyinput17), .ZN(n8848) );
  XNOR2_X1 U10387 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput2), .ZN(n8847) );
  XNOR2_X1 U10388 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput89), .ZN(n8846) );
  XNOR2_X1 U10389 ( .A(P2_REG1_REG_31__SCAN_IN), .B(keyinput24), .ZN(n8845) );
  NAND4_X1 U10390 ( .A1(n8848), .A2(n8847), .A3(n8846), .A4(n8845), .ZN(n8849)
         );
  NOR2_X1 U10391 ( .A1(n8850), .A2(n8849), .ZN(n8875) );
  XNOR2_X1 U10392 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput9), .ZN(n8854) );
  XNOR2_X1 U10393 ( .A(P2_REG2_REG_12__SCAN_IN), .B(keyinput33), .ZN(n8853) );
  XNOR2_X1 U10394 ( .A(P2_IR_REG_16__SCAN_IN), .B(keyinput126), .ZN(n8852) );
  XNOR2_X1 U10395 ( .A(P2_IR_REG_19__SCAN_IN), .B(keyinput42), .ZN(n8851) );
  NAND4_X1 U10396 ( .A1(n8854), .A2(n8853), .A3(n8852), .A4(n8851), .ZN(n8860)
         );
  XNOR2_X1 U10397 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(keyinput59), .ZN(n8858) );
  XNOR2_X1 U10398 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput46), .ZN(n8857) );
  XNOR2_X1 U10399 ( .A(P1_REG1_REG_1__SCAN_IN), .B(keyinput18), .ZN(n8856) );
  XNOR2_X1 U10400 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput55), .ZN(n8855) );
  NAND4_X1 U10401 ( .A1(n8858), .A2(n8857), .A3(n8856), .A4(n8855), .ZN(n8859)
         );
  NOR2_X1 U10402 ( .A1(n8860), .A2(n8859), .ZN(n8874) );
  XNOR2_X1 U10403 ( .A(P2_IR_REG_4__SCAN_IN), .B(keyinput57), .ZN(n8864) );
  XNOR2_X1 U10404 ( .A(P1_REG2_REG_15__SCAN_IN), .B(keyinput56), .ZN(n8863) );
  XNOR2_X1 U10405 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(keyinput10), .ZN(n8862)
         );
  XNOR2_X1 U10406 ( .A(P2_IR_REG_29__SCAN_IN), .B(keyinput27), .ZN(n8861) );
  NAND4_X1 U10407 ( .A1(n8864), .A2(n8863), .A3(n8862), .A4(n8861), .ZN(n8870)
         );
  XNOR2_X1 U10408 ( .A(SI_3_), .B(keyinput11), .ZN(n8868) );
  XNOR2_X1 U10409 ( .A(SI_1_), .B(keyinput90), .ZN(n8867) );
  XNOR2_X1 U10410 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(keyinput13), .ZN(n8866) );
  XNOR2_X1 U10411 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput7), .ZN(n8865) );
  NAND4_X1 U10412 ( .A1(n8868), .A2(n8867), .A3(n8866), .A4(n8865), .ZN(n8869)
         );
  NOR2_X1 U10413 ( .A1(n8870), .A2(n8869), .ZN(n8873) );
  INV_X1 U10414 ( .A(keyinput58), .ZN(n8871) );
  XNOR2_X1 U10415 ( .A(n10396), .B(n8871), .ZN(n8872) );
  NAND4_X1 U10416 ( .A1(n8875), .A2(n8874), .A3(n8873), .A4(n8872), .ZN(n8876)
         );
  NOR2_X1 U10417 ( .A1(n8877), .A2(n8876), .ZN(n8947) );
  AOI22_X1 U10418 ( .A1(n9036), .A2(keyinput120), .B1(keyinput75), .B2(n10390), 
        .ZN(n8878) );
  OAI221_X1 U10419 ( .B1(n9036), .B2(keyinput120), .C1(n10390), .C2(keyinput75), .A(n8878), .ZN(n8884) );
  AOI22_X1 U10420 ( .A1(n8880), .A2(keyinput40), .B1(keyinput121), .B2(n9019), 
        .ZN(n8879) );
  OAI221_X1 U10421 ( .B1(n8880), .B2(keyinput40), .C1(n9019), .C2(keyinput121), 
        .A(n8879), .ZN(n8883) );
  INV_X1 U10422 ( .A(keyinput116), .ZN(n8881) );
  XNOR2_X1 U10423 ( .A(n8881), .B(P1_ADDR_REG_14__SCAN_IN), .ZN(n8882) );
  NOR3_X1 U10424 ( .A1(n8884), .A2(n8883), .A3(n8882), .ZN(n8914) );
  INV_X1 U10425 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9363) );
  AOI22_X1 U10426 ( .A1(n5613), .A2(keyinput52), .B1(keyinput4), .B2(n9363), 
        .ZN(n8885) );
  OAI221_X1 U10427 ( .B1(n5613), .B2(keyinput52), .C1(n9363), .C2(keyinput4), 
        .A(n8885), .ZN(n8891) );
  INV_X1 U10428 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n8887) );
  INV_X1 U10429 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9151) );
  AOI22_X1 U10430 ( .A1(n8887), .A2(keyinput39), .B1(n9151), .B2(keyinput85), 
        .ZN(n8886) );
  OAI221_X1 U10431 ( .B1(n8887), .B2(keyinput39), .C1(n9151), .C2(keyinput85), 
        .A(n8886), .ZN(n8890) );
  XNOR2_X1 U10432 ( .A(n8888), .B(keyinput25), .ZN(n8889) );
  NOR3_X1 U10433 ( .A1(n8891), .A2(n8890), .A3(n8889), .ZN(n8913) );
  AOI22_X1 U10434 ( .A1(n5119), .A2(keyinput72), .B1(n8893), .B2(keyinput8), 
        .ZN(n8892) );
  OAI221_X1 U10435 ( .B1(n5119), .B2(keyinput72), .C1(n8893), .C2(keyinput8), 
        .A(n8892), .ZN(n8899) );
  XNOR2_X1 U10436 ( .A(P1_REG3_REG_21__SCAN_IN), .B(keyinput93), .ZN(n8897) );
  XNOR2_X1 U10437 ( .A(P1_IR_REG_21__SCAN_IN), .B(keyinput105), .ZN(n8896) );
  XNOR2_X1 U10438 ( .A(P2_D_REG_0__SCAN_IN), .B(keyinput49), .ZN(n8895) );
  XNOR2_X1 U10439 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput95), .ZN(n8894) );
  NAND4_X1 U10440 ( .A1(n8897), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(n8898)
         );
  NOR2_X1 U10441 ( .A1(n8899), .A2(n8898), .ZN(n8905) );
  INV_X1 U10442 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U10443 ( .A1(n10196), .A2(keyinput117), .B1(n8992), .B2(keyinput47), 
        .ZN(n8900) );
  OAI221_X1 U10444 ( .B1(n10196), .B2(keyinput117), .C1(n8992), .C2(keyinput47), .A(n8900), .ZN(n8903) );
  INV_X1 U10445 ( .A(keyinput26), .ZN(n8901) );
  XNOR2_X1 U10446 ( .A(n8901), .B(P1_ADDR_REG_13__SCAN_IN), .ZN(n8902) );
  NOR2_X1 U10447 ( .A1(n8903), .A2(n8902), .ZN(n8904) );
  AND2_X1 U10448 ( .A1(n8905), .A2(n8904), .ZN(n8912) );
  AOI22_X1 U10449 ( .A1(n8652), .A2(keyinput99), .B1(keyinput103), .B2(n9010), 
        .ZN(n8906) );
  OAI221_X1 U10450 ( .B1(n8652), .B2(keyinput99), .C1(n9010), .C2(keyinput103), 
        .A(n8906), .ZN(n8910) );
  INV_X1 U10451 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8908) );
  AOI22_X1 U10452 ( .A1(n8908), .A2(keyinput54), .B1(keyinput97), .B2(n8990), 
        .ZN(n8907) );
  OAI221_X1 U10453 ( .B1(n8908), .B2(keyinput54), .C1(n8990), .C2(keyinput97), 
        .A(n8907), .ZN(n8909) );
  NOR2_X1 U10454 ( .A1(n8910), .A2(n8909), .ZN(n8911) );
  NAND4_X1 U10455 ( .A1(n8914), .A2(n8913), .A3(n8912), .A4(n8911), .ZN(n8945)
         );
  AOI22_X1 U10456 ( .A1(n8916), .A2(keyinput20), .B1(keyinput91), .B2(n10374), 
        .ZN(n8915) );
  OAI221_X1 U10457 ( .B1(n8916), .B2(keyinput20), .C1(n10374), .C2(keyinput91), 
        .A(n8915), .ZN(n8921) );
  INV_X1 U10458 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9057) );
  AOI22_X1 U10459 ( .A1(n9057), .A2(keyinput118), .B1(keyinput102), .B2(n9083), 
        .ZN(n8917) );
  OAI221_X1 U10460 ( .B1(n9057), .B2(keyinput118), .C1(n9083), .C2(keyinput102), .A(n8917), .ZN(n8920) );
  AOI22_X1 U10461 ( .A1(n9039), .A2(keyinput68), .B1(keyinput44), .B2(n9953), 
        .ZN(n8918) );
  OAI221_X1 U10462 ( .B1(n9039), .B2(keyinput68), .C1(n9953), .C2(keyinput44), 
        .A(n8918), .ZN(n8919) );
  NOR3_X1 U10463 ( .A1(n8921), .A2(n8920), .A3(n8919), .ZN(n8943) );
  AOI22_X1 U10464 ( .A1(n8923), .A2(keyinput70), .B1(n8709), .B2(keyinput94), 
        .ZN(n8922) );
  OAI221_X1 U10465 ( .B1(n8923), .B2(keyinput70), .C1(n8709), .C2(keyinput94), 
        .A(n8922), .ZN(n8926) );
  AOI22_X1 U10466 ( .A1(n6845), .A2(keyinput51), .B1(n7352), .B2(keyinput81), 
        .ZN(n8924) );
  OAI221_X1 U10467 ( .B1(n6845), .B2(keyinput51), .C1(n7352), .C2(keyinput81), 
        .A(n8924), .ZN(n8925) );
  NOR2_X1 U10468 ( .A1(n8926), .A2(n8925), .ZN(n8942) );
  INV_X1 U10469 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n8928) );
  AOI22_X1 U10470 ( .A1(n9021), .A2(keyinput98), .B1(keyinput32), .B2(n8928), 
        .ZN(n8927) );
  OAI221_X1 U10471 ( .B1(n9021), .B2(keyinput98), .C1(n8928), .C2(keyinput32), 
        .A(n8927), .ZN(n8932) );
  INV_X1 U10472 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U10473 ( .A1(n8930), .A2(keyinput113), .B1(keyinput62), .B2(n10197), 
        .ZN(n8929) );
  OAI221_X1 U10474 ( .B1(n8930), .B2(keyinput113), .C1(n10197), .C2(keyinput62), .A(n8929), .ZN(n8931) );
  NOR2_X1 U10475 ( .A1(n8932), .A2(n8931), .ZN(n8941) );
  AOI22_X1 U10476 ( .A1(n8999), .A2(keyinput123), .B1(keyinput45), .B2(n8934), 
        .ZN(n8933) );
  OAI221_X1 U10477 ( .B1(n8999), .B2(keyinput123), .C1(n8934), .C2(keyinput45), 
        .A(n8933), .ZN(n8939) );
  AOI22_X1 U10478 ( .A1(n8937), .A2(keyinput87), .B1(keyinput14), .B2(n8936), 
        .ZN(n8935) );
  OAI221_X1 U10479 ( .B1(n8937), .B2(keyinput87), .C1(n8936), .C2(keyinput14), 
        .A(n8935), .ZN(n8938) );
  NOR2_X1 U10480 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  NAND4_X1 U10481 ( .A1(n8943), .A2(n8942), .A3(n8941), .A4(n8940), .ZN(n8944)
         );
  NOR2_X1 U10482 ( .A1(n8945), .A2(n8944), .ZN(n8946) );
  AND4_X1 U10483 ( .A1(n8949), .A2(n8948), .A3(n8947), .A4(n8946), .ZN(n8973)
         );
  AOI22_X1 U10484 ( .A1(n8952), .A2(keyinput76), .B1(keyinput71), .B2(n8951), 
        .ZN(n8950) );
  OAI221_X1 U10485 ( .B1(n8952), .B2(keyinput76), .C1(n8951), .C2(keyinput71), 
        .A(n8950), .ZN(n8961) );
  AOI22_X1 U10486 ( .A1(n8955), .A2(keyinput83), .B1(keyinput15), .B2(n8954), 
        .ZN(n8953) );
  OAI221_X1 U10487 ( .B1(n8955), .B2(keyinput83), .C1(n8954), .C2(keyinput15), 
        .A(n8953), .ZN(n8960) );
  INV_X1 U10488 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9124) );
  AOI22_X1 U10489 ( .A1(n9984), .A2(keyinput106), .B1(n9124), .B2(keyinput36), 
        .ZN(n8956) );
  OAI221_X1 U10490 ( .B1(n9984), .B2(keyinput106), .C1(n9124), .C2(keyinput36), 
        .A(n8956), .ZN(n8959) );
  AOI22_X1 U10491 ( .A1(n8977), .A2(keyinput108), .B1(keyinput73), .B2(n10382), 
        .ZN(n8957) );
  OAI221_X1 U10492 ( .B1(n8977), .B2(keyinput108), .C1(n10382), .C2(keyinput73), .A(n8957), .ZN(n8958) );
  NOR4_X1 U10493 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n8972)
         );
  AOI22_X1 U10494 ( .A1(n7083), .A2(keyinput21), .B1(n6803), .B2(keyinput101), 
        .ZN(n8962) );
  OAI221_X1 U10495 ( .B1(n7083), .B2(keyinput21), .C1(n6803), .C2(keyinput101), 
        .A(n8962), .ZN(n8970) );
  AOI22_X1 U10496 ( .A1(n8964), .A2(keyinput1), .B1(n9020), .B2(keyinput6), 
        .ZN(n8963) );
  OAI221_X1 U10497 ( .B1(n8964), .B2(keyinput1), .C1(n9020), .C2(keyinput6), 
        .A(n8963), .ZN(n8969) );
  INV_X1 U10498 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9170) );
  AOI22_X1 U10499 ( .A1(n9170), .A2(keyinput111), .B1(n9974), .B2(keyinput31), 
        .ZN(n8965) );
  OAI221_X1 U10500 ( .B1(n9170), .B2(keyinput111), .C1(n9974), .C2(keyinput31), 
        .A(n8965), .ZN(n8968) );
  AOI22_X1 U10501 ( .A1(n9016), .A2(keyinput28), .B1(keyinput43), .B2(n10166), 
        .ZN(n8966) );
  OAI221_X1 U10502 ( .B1(n9016), .B2(keyinput28), .C1(n10166), .C2(keyinput43), 
        .A(n8966), .ZN(n8967) );
  NOR4_X1 U10503 ( .A1(n8970), .A2(n8969), .A3(n8968), .A4(n8967), .ZN(n8971)
         );
  NAND3_X1 U10504 ( .A1(n8973), .A2(n8972), .A3(n8971), .ZN(n9049) );
  NOR4_X1 U10505 ( .A1(n8977), .A2(n8976), .A3(n8975), .A4(n8974), .ZN(n9009)
         );
  NOR4_X1 U10506 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P1_ADDR_REG_19__SCAN_IN), .A4(P2_DATAO_REG_23__SCAN_IN), .ZN(n9008) );
  NOR4_X1 U10507 ( .A1(P2_D_REG_1__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .A3(
        P2_REG3_REG_22__SCAN_IN), .A4(n8978), .ZN(n8979) );
  NAND3_X1 U10508 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        n8979), .ZN(n8987) );
  NOR4_X1 U10509 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .A3(P1_ADDR_REG_2__SCAN_IN), .A4(P2_ADDR_REG_7__SCAN_IN), .ZN(n8983)
         );
  NAND2_X1 U10510 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8981) );
  NAND4_X1 U10511 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), 
        .A3(P2_IR_REG_10__SCAN_IN), .A4(P2_IR_REG_9__SCAN_IN), .ZN(n8980) );
  NOR4_X1 U10512 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .A3(
        n8981), .A4(n8980), .ZN(n8982) );
  NAND4_X1 U10513 ( .A1(n8985), .A2(n8984), .A3(n8983), .A4(n8982), .ZN(n8986)
         );
  NOR4_X1 U10514 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .A3(
        n8987), .A4(n8986), .ZN(n9007) );
  NOR4_X1 U10515 ( .A1(P1_REG1_REG_23__SCAN_IN), .A2(P1_REG2_REG_5__SCAN_IN), 
        .A3(n6803), .A4(n9170), .ZN(n8988) );
  NAND3_X1 U10516 ( .A1(P1_REG1_REG_28__SCAN_IN), .A2(n8988), .A3(n10416), 
        .ZN(n9005) );
  NAND4_X1 U10517 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_REG0_REG_25__SCAN_IN), 
        .A3(P1_REG2_REG_10__SCAN_IN), .A4(P1_REG2_REG_31__SCAN_IN), .ZN(n8989)
         );
  NOR3_X1 U10518 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_REG3_REG_20__SCAN_IN), 
        .A3(n8989), .ZN(n9003) );
  NOR4_X1 U10519 ( .A1(n8992), .A2(n8991), .A3(n8990), .A4(
        P1_REG1_REG_1__SCAN_IN), .ZN(n8998) );
  NAND4_X1 U10520 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .A3(n8994), .A4(n8993), .ZN(n8995) );
  NOR3_X1 U10521 ( .A1(n7523), .A2(P1_IR_REG_15__SCAN_IN), .A3(n8995), .ZN(
        n8997) );
  NAND4_X1 U10522 ( .A1(n8998), .A2(P1_REG0_REG_11__SCAN_IN), .A3(n8997), .A4(
        n8996), .ZN(n9001) );
  NAND4_X1 U10523 ( .A1(SI_26_), .A2(P1_ADDR_REG_15__SCAN_IN), .A3(n8999), 
        .A4(n8571), .ZN(n9000) );
  NOR2_X1 U10524 ( .A1(n9001), .A2(n9000), .ZN(n9002) );
  NAND4_X1 U10525 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), 
        .A3(n9003), .A4(n9002), .ZN(n9004) );
  NOR4_X1 U10526 ( .A1(P1_D_REG_1__SCAN_IN), .A2(P1_REG2_REG_18__SCAN_IN), 
        .A3(n9005), .A4(n9004), .ZN(n9006) );
  NAND4_X1 U10527 ( .A1(n9009), .A2(n9008), .A3(n9007), .A4(n9006), .ZN(n9033)
         );
  NOR4_X1 U10528 ( .A1(P2_REG0_REG_22__SCAN_IN), .A2(P2_REG2_REG_20__SCAN_IN), 
        .A3(P2_REG1_REG_20__SCAN_IN), .A4(n10289), .ZN(n9014) );
  NOR4_X1 U10529 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), 
        .A3(SI_21_), .A4(P2_REG1_REG_22__SCAN_IN), .ZN(n9013) );
  NOR4_X1 U10530 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(P2_REG2_REG_9__SCAN_IN), .A4(n9010), .ZN(n9012) );
  NOR4_X1 U10531 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(P2_REG2_REG_16__SCAN_IN), 
        .A3(P2_REG1_REG_15__SCAN_IN), .A4(n9151), .ZN(n9011) );
  NAND4_X1 U10532 ( .A1(n9014), .A2(n9013), .A3(n9012), .A4(n9011), .ZN(n9032)
         );
  INV_X1 U10533 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9015) );
  NAND4_X1 U10534 ( .A1(n10380), .A2(n9015), .A3(P2_REG2_REG_7__SCAN_IN), .A4(
        P2_REG0_REG_0__SCAN_IN), .ZN(n9031) );
  NOR4_X1 U10535 ( .A1(SI_9_), .A2(n9018), .A3(n9017), .A4(n9016), .ZN(n9024)
         );
  NOR4_X1 U10536 ( .A1(n9021), .A2(n9020), .A3(n9019), .A4(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n9023) );
  NOR4_X1 U10537 ( .A1(SI_4_), .A2(SI_3_), .A3(P1_DATAO_REG_2__SCAN_IN), .A4(
        SI_1_), .ZN(n9022) );
  NAND4_X1 U10538 ( .A1(n9025), .A2(n9024), .A3(n9023), .A4(n9022), .ZN(n9026)
         );
  NOR4_X1 U10539 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P2_DATAO_REG_7__SCAN_IN), 
        .A3(P1_DATAO_REG_5__SCAN_IN), .A4(n9026), .ZN(n9029) );
  NOR2_X1 U10540 ( .A1(n9027), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9028) );
  NAND4_X1 U10541 ( .A1(n9029), .A2(P2_REG1_REG_4__SCAN_IN), .A3(
        P2_DATAO_REG_5__SCAN_IN), .A4(n9028), .ZN(n9030) );
  NOR4_X1 U10542 ( .A1(n9033), .A2(n9032), .A3(n9031), .A4(n9030), .ZN(n9047)
         );
  NOR4_X1 U10543 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(P1_REG2_REG_20__SCAN_IN), 
        .A3(SI_31_), .A4(P2_ADDR_REG_16__SCAN_IN), .ZN(n9034) );
  NAND3_X1 U10544 ( .A1(P2_REG2_REG_28__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), 
        .A3(n9034), .ZN(n9045) );
  NOR4_X1 U10545 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .A3(n9036), .A4(n9035), .ZN(n9043) );
  NOR4_X1 U10546 ( .A1(P2_REG0_REG_12__SCAN_IN), .A2(P2_REG1_REG_10__SCAN_IN), 
        .A3(P2_REG1_REG_6__SCAN_IN), .A4(n9037), .ZN(n9042) );
  NOR4_X1 U10547 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_REG1_REG_27__SCAN_IN), 
        .A3(P1_REG0_REG_28__SCAN_IN), .A4(n10131), .ZN(n9041) );
  NOR4_X1 U10548 ( .A1(P1_REG2_REG_30__SCAN_IN), .A2(n10200), .A3(n9039), .A4(
        n9038), .ZN(n9040) );
  NAND4_X1 U10549 ( .A1(n9043), .A2(n9042), .A3(n9041), .A4(n9040), .ZN(n9044)
         );
  NOR4_X1 U10550 ( .A1(P1_B_REG_SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), .A3(
        n9045), .A4(n9044), .ZN(n9046) );
  NAND2_X1 U10551 ( .A1(n9047), .A2(n9046), .ZN(n9048) );
  XOR2_X1 U10552 ( .A(n9049), .B(n9048), .Z(n9050) );
  XNOR2_X1 U10553 ( .A(n9051), .B(n9050), .ZN(P2_U3483) );
  INV_X1 U10554 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9052) );
  MUX2_X1 U10555 ( .A(n9052), .B(n9117), .S(n10384), .Z(n9054) );
  NAND2_X1 U10556 ( .A1(n9119), .A2(n9084), .ZN(n9053) );
  OAI211_X1 U10557 ( .C1(n9122), .C2(n9087), .A(n9054), .B(n9053), .ZN(
        P2_U3482) );
  AOI21_X1 U10558 ( .B1(n9071), .B2(n9056), .A(n9055), .ZN(n9123) );
  MUX2_X1 U10559 ( .A(n9057), .B(n9123), .S(n10384), .Z(n9058) );
  OAI21_X1 U10560 ( .B1(n9126), .B2(n9075), .A(n9058), .ZN(P2_U3481) );
  INV_X1 U10561 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9061) );
  AOI21_X1 U10562 ( .B1(n9060), .B2(n9071), .A(n9059), .ZN(n9127) );
  MUX2_X1 U10563 ( .A(n9061), .B(n9127), .S(n10384), .Z(n9062) );
  OAI21_X1 U10564 ( .B1(n9130), .B2(n9075), .A(n9062), .ZN(P2_U3480) );
  MUX2_X1 U10565 ( .A(n9063), .B(n9131), .S(n10384), .Z(n9065) );
  NAND2_X1 U10566 ( .A1(n9133), .A2(n9084), .ZN(n9064) );
  OAI211_X1 U10567 ( .C1(n9087), .C2(n9136), .A(n9065), .B(n9064), .ZN(
        P2_U3479) );
  MUX2_X1 U10568 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9137), .S(n10384), .Z(
        n9066) );
  INV_X1 U10569 ( .A(n9066), .ZN(n9069) );
  OAI22_X1 U10570 ( .A1(n9140), .A2(n9087), .B1(n9139), .B2(n9075), .ZN(n9067)
         );
  INV_X1 U10571 ( .A(n9067), .ZN(n9068) );
  NAND2_X1 U10572 ( .A1(n9069), .A2(n9068), .ZN(P2_U3478) );
  AOI21_X1 U10573 ( .B1(n9072), .B2(n9071), .A(n9070), .ZN(n9144) );
  MUX2_X1 U10574 ( .A(n9073), .B(n9144), .S(n10384), .Z(n9074) );
  OAI21_X1 U10575 ( .B1(n9148), .B2(n9075), .A(n9074), .ZN(P2_U3477) );
  NAND2_X1 U10576 ( .A1(n9076), .A2(n10325), .ZN(n9077) );
  OAI211_X1 U10577 ( .C1(n10353), .C2(n9079), .A(n9078), .B(n9077), .ZN(n9149)
         );
  MUX2_X1 U10578 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9149), .S(n10384), .Z(
        P2_U3476) );
  MUX2_X1 U10579 ( .A(n9080), .B(n9150), .S(n10384), .Z(n9082) );
  NAND2_X1 U10580 ( .A1(n9152), .A2(n9084), .ZN(n9081) );
  OAI211_X1 U10581 ( .C1(n9155), .C2(n9087), .A(n9082), .B(n9081), .ZN(
        P2_U3475) );
  MUX2_X1 U10582 ( .A(n9083), .B(n9156), .S(n10384), .Z(n9086) );
  NAND2_X1 U10583 ( .A1(n9159), .A2(n9084), .ZN(n9085) );
  OAI211_X1 U10584 ( .C1(n9087), .C2(n9163), .A(n9086), .B(n9085), .ZN(
        P2_U3473) );
  INV_X1 U10585 ( .A(n9088), .ZN(n9091) );
  NAND2_X1 U10586 ( .A1(n9089), .A2(n10367), .ZN(n9092) );
  NAND2_X1 U10587 ( .A1(n10365), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9090) );
  OAI211_X1 U10588 ( .C1(n9091), .C2(n9147), .A(n9092), .B(n9090), .ZN(
        P2_U3458) );
  NAND2_X1 U10589 ( .A1(n10365), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9093) );
  OAI211_X1 U10590 ( .C1(n9094), .C2(n9147), .A(n9093), .B(n9092), .ZN(
        P2_U3457) );
  INV_X1 U10591 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9096) );
  MUX2_X1 U10592 ( .A(n9096), .B(n9095), .S(n10367), .Z(n9099) );
  NAND2_X1 U10593 ( .A1(n9097), .A2(n9158), .ZN(n9098) );
  OAI211_X1 U10594 ( .C1(n9100), .C2(n9162), .A(n9099), .B(n9098), .ZN(
        P2_U3455) );
  INV_X1 U10595 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9102) );
  MUX2_X1 U10596 ( .A(n9102), .B(n9101), .S(n10367), .Z(n9105) );
  NAND2_X1 U10597 ( .A1(n9103), .A2(n9158), .ZN(n9104) );
  OAI211_X1 U10598 ( .C1(n9106), .C2(n9162), .A(n9105), .B(n9104), .ZN(
        P2_U3454) );
  INV_X1 U10599 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9108) );
  MUX2_X1 U10600 ( .A(n9108), .B(n9107), .S(n10367), .Z(n9109) );
  OAI21_X1 U10601 ( .B1(n9110), .B2(n9147), .A(n9109), .ZN(P2_U3453) );
  INV_X1 U10602 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9112) );
  MUX2_X1 U10603 ( .A(n9112), .B(n9111), .S(n10367), .Z(n9113) );
  OAI21_X1 U10604 ( .B1(n9114), .B2(n9162), .A(n9113), .ZN(P2_U3452) );
  NAND2_X1 U10605 ( .A1(n10365), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9115) );
  OAI21_X1 U10606 ( .B1(n9116), .B2(n10365), .A(n9115), .ZN(P2_U3451) );
  INV_X1 U10607 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9118) );
  MUX2_X1 U10608 ( .A(n9118), .B(n9117), .S(n10367), .Z(n9121) );
  NAND2_X1 U10609 ( .A1(n9119), .A2(n9158), .ZN(n9120) );
  OAI211_X1 U10610 ( .C1(n9122), .C2(n9162), .A(n9121), .B(n9120), .ZN(
        P2_U3450) );
  MUX2_X1 U10611 ( .A(n9124), .B(n9123), .S(n10367), .Z(n9125) );
  OAI21_X1 U10612 ( .B1(n9126), .B2(n9147), .A(n9125), .ZN(P2_U3449) );
  INV_X1 U10613 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9128) );
  MUX2_X1 U10614 ( .A(n9128), .B(n9127), .S(n10367), .Z(n9129) );
  OAI21_X1 U10615 ( .B1(n9130), .B2(n9147), .A(n9129), .ZN(P2_U3448) );
  INV_X1 U10616 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9132) );
  MUX2_X1 U10617 ( .A(n9132), .B(n9131), .S(n10367), .Z(n9135) );
  NAND2_X1 U10618 ( .A1(n9133), .A2(n9158), .ZN(n9134) );
  OAI211_X1 U10619 ( .C1(n9136), .C2(n9162), .A(n9135), .B(n9134), .ZN(
        P2_U3447) );
  MUX2_X1 U10620 ( .A(n9137), .B(P2_REG0_REG_19__SCAN_IN), .S(n10365), .Z(
        n9138) );
  INV_X1 U10621 ( .A(n9138), .ZN(n9143) );
  OAI22_X1 U10622 ( .A1(n9140), .A2(n9162), .B1(n9139), .B2(n9147), .ZN(n9141)
         );
  INV_X1 U10623 ( .A(n9141), .ZN(n9142) );
  NAND2_X1 U10624 ( .A1(n9143), .A2(n9142), .ZN(P2_U3446) );
  INV_X1 U10625 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9145) );
  MUX2_X1 U10626 ( .A(n9145), .B(n9144), .S(n10367), .Z(n9146) );
  OAI21_X1 U10627 ( .B1(n9148), .B2(n9147), .A(n9146), .ZN(P2_U3444) );
  MUX2_X1 U10628 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9149), .S(n10367), .Z(
        P2_U3441) );
  MUX2_X1 U10629 ( .A(n9151), .B(n9150), .S(n10367), .Z(n9154) );
  NAND2_X1 U10630 ( .A1(n9152), .A2(n9158), .ZN(n9153) );
  OAI211_X1 U10631 ( .C1(n9155), .C2(n9162), .A(n9154), .B(n9153), .ZN(
        P2_U3438) );
  INV_X1 U10632 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9157) );
  MUX2_X1 U10633 ( .A(n9157), .B(n9156), .S(n10367), .Z(n9161) );
  NAND2_X1 U10634 ( .A1(n9159), .A2(n9158), .ZN(n9160) );
  OAI211_X1 U10635 ( .C1(n9163), .C2(n9162), .A(n9161), .B(n9160), .ZN(
        P2_U3432) );
  INV_X1 U10636 ( .A(n9357), .ZN(n10078) );
  NOR4_X1 U10637 ( .A1(n9164), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n6099), .ZN(n9165) );
  AOI21_X1 U10638 ( .B1(n9166), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9165), .ZN(
        n9167) );
  OAI21_X1 U10639 ( .B1(n10078), .B2(n9169), .A(n9167), .ZN(P2_U3264) );
  INV_X1 U10640 ( .A(n9408), .ZN(n10081) );
  OAI222_X1 U10641 ( .A1(n9171), .A2(n9170), .B1(n9169), .B2(n10081), .C1(
        P2_U3151), .C2(n9168), .ZN(P2_U3265) );
  MUX2_X1 U10642 ( .A(n9172), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10643 ( .A(n9173), .ZN(n9174) );
  NAND2_X1 U10644 ( .A1(n9175), .A2(n9174), .ZN(n9179) );
  XNOR2_X1 U10645 ( .A(n9177), .B(n9176), .ZN(n9178) );
  XNOR2_X1 U10646 ( .A(n9179), .B(n9178), .ZN(n9185) );
  NAND2_X1 U10647 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10143)
         );
  NAND2_X1 U10648 ( .A1(n9346), .A2(n9180), .ZN(n9181) );
  OAI211_X1 U10649 ( .C1(n9349), .C2(n9182), .A(n10143), .B(n9181), .ZN(n9183)
         );
  AOI21_X1 U10650 ( .B1(n10015), .B2(n9351), .A(n9183), .ZN(n9184) );
  OAI21_X1 U10651 ( .B1(n9185), .B2(n9354), .A(n9184), .ZN(P1_U3215) );
  AND3_X1 U10652 ( .A1(n9187), .A2(n9189), .A3(n9188), .ZN(n9190) );
  OAI21_X1 U10653 ( .B1(n9186), .B2(n9190), .A(n9329), .ZN(n9194) );
  OAI22_X1 U10654 ( .A1(n9235), .A2(n9301), .B1(n9217), .B2(n9300), .ZN(n9820)
         );
  OAI22_X1 U10655 ( .A1(n9828), .A2(n9349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9191), .ZN(n9192) );
  AOI21_X1 U10656 ( .B1(n9820), .B2(n9346), .A(n9192), .ZN(n9193) );
  OAI211_X1 U10657 ( .C1(n10050), .C2(n9283), .A(n9194), .B(n9193), .ZN(
        P1_U3216) );
  OAI21_X1 U10658 ( .B1(n9197), .B2(n9196), .A(n9195), .ZN(n9198) );
  NAND2_X1 U10659 ( .A1(n9198), .A2(n9329), .ZN(n9204) );
  NOR2_X1 U10660 ( .A1(n9349), .A2(n9199), .ZN(n9200) );
  AOI211_X1 U10661 ( .C1(n9346), .C2(n9202), .A(n9201), .B(n9200), .ZN(n9203)
         );
  OAI211_X1 U10662 ( .C1(n9205), .C2(n9283), .A(n9204), .B(n9203), .ZN(
        P1_U3217) );
  XNOR2_X1 U10663 ( .A(n9208), .B(n9207), .ZN(n9209) );
  XNOR2_X1 U10664 ( .A(n9206), .B(n9209), .ZN(n9213) );
  OAI22_X1 U10665 ( .A1(n9371), .A2(n9301), .B1(n9259), .B2(n9300), .ZN(n9898)
         );
  AOI22_X1 U10666 ( .A1(n9898), .A2(n9346), .B1(P1_REG3_REG_19__SCAN_IN), .B2(
        P1_U3086), .ZN(n9210) );
  OAI21_X1 U10667 ( .B1(n9349), .B2(n9889), .A(n9210), .ZN(n9211) );
  AOI21_X1 U10668 ( .B1(n9992), .B2(n9351), .A(n9211), .ZN(n9212) );
  OAI21_X1 U10669 ( .B1(n9213), .B2(n9354), .A(n9212), .ZN(P1_U3219) );
  OAI21_X1 U10670 ( .B1(n9216), .B2(n9215), .A(n9214), .ZN(n9221) );
  NAND2_X1 U10671 ( .A1(n9861), .A2(n9351), .ZN(n9219) );
  OAI22_X1 U10672 ( .A1(n9217), .A2(n9301), .B1(n9371), .B2(n9300), .ZN(n9853)
         );
  AOI22_X1 U10673 ( .A1(n9853), .A2(n9346), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9218) );
  OAI211_X1 U10674 ( .C1(n9349), .C2(n9862), .A(n9219), .B(n9218), .ZN(n9220)
         );
  AOI21_X1 U10675 ( .B1(n9221), .B2(n9329), .A(n9220), .ZN(n9222) );
  INV_X1 U10676 ( .A(n9222), .ZN(P1_U3223) );
  XOR2_X1 U10677 ( .A(n9223), .B(n9224), .Z(n9231) );
  AOI22_X1 U10678 ( .A1(n9346), .A2(n9225), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3086), .ZN(n9226) );
  OAI21_X1 U10679 ( .B1(n9349), .B2(n9227), .A(n9226), .ZN(n9228) );
  AOI21_X1 U10680 ( .B1(n9229), .B2(n9351), .A(n9228), .ZN(n9230) );
  OAI21_X1 U10681 ( .B1(n9231), .B2(n9354), .A(n9230), .ZN(P1_U3224) );
  OAI21_X1 U10682 ( .B1(n9233), .B2(n9232), .A(n5882), .ZN(n9234) );
  NAND2_X1 U10683 ( .A1(n9234), .A2(n9329), .ZN(n9241) );
  OAI22_X1 U10684 ( .A1(n9236), .A2(n9301), .B1(n9235), .B2(n9300), .ZN(n9786)
         );
  INV_X1 U10685 ( .A(n9793), .ZN(n9238) );
  OAI22_X1 U10686 ( .A1(n9238), .A2(n9349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9237), .ZN(n9239) );
  AOI21_X1 U10687 ( .B1(n9786), .B2(n9346), .A(n9239), .ZN(n9240) );
  OAI211_X1 U10688 ( .C1(n10043), .C2(n9283), .A(n9241), .B(n9240), .ZN(
        P1_U3225) );
  XNOR2_X1 U10689 ( .A(n9242), .B(n9243), .ZN(n9343) );
  NOR2_X1 U10690 ( .A1(n9343), .A2(n9344), .ZN(n9342) );
  AOI21_X1 U10691 ( .B1(n9243), .B2(n9242), .A(n9342), .ZN(n9247) );
  XNOR2_X1 U10692 ( .A(n9245), .B(n9244), .ZN(n9246) );
  XNOR2_X1 U10693 ( .A(n9247), .B(n9246), .ZN(n9254) );
  NAND2_X1 U10694 ( .A1(n9346), .A2(n9248), .ZN(n9249) );
  OAI211_X1 U10695 ( .C1(n9349), .C2(n9251), .A(n9250), .B(n9249), .ZN(n9252)
         );
  AOI21_X1 U10696 ( .B1(n10011), .B2(n9351), .A(n9252), .ZN(n9253) );
  OAI21_X1 U10697 ( .B1(n9254), .B2(n9354), .A(n9253), .ZN(P1_U3226) );
  NOR2_X1 U10698 ( .A1(n9256), .A2(n4517), .ZN(n9257) );
  XNOR2_X1 U10699 ( .A(n9255), .B(n9257), .ZN(n9263) );
  OAI22_X1 U10700 ( .A1(n9259), .A2(n9301), .B1(n9258), .B2(n9300), .ZN(n9930)
         );
  AOI22_X1 U10701 ( .A1(n9346), .A2(n9930), .B1(P1_REG3_REG_17__SCAN_IN), .B2(
        P1_U3086), .ZN(n9260) );
  OAI21_X1 U10702 ( .B1(n9349), .B2(n9924), .A(n9260), .ZN(n9261) );
  AOI21_X1 U10703 ( .B1(n10003), .B2(n9351), .A(n9261), .ZN(n9262) );
  OAI21_X1 U10704 ( .B1(n9263), .B2(n9354), .A(n9262), .ZN(P1_U3228) );
  INV_X1 U10705 ( .A(n9264), .ZN(n9268) );
  NOR3_X1 U10706 ( .A1(n9186), .A2(n9266), .A3(n9265), .ZN(n9267) );
  OAI21_X1 U10707 ( .B1(n9268), .B2(n9267), .A(n9329), .ZN(n9276) );
  OR2_X1 U10708 ( .A1(n9269), .A2(n9301), .ZN(n9271) );
  NAND2_X1 U10709 ( .A1(n9625), .A2(n9320), .ZN(n9270) );
  NAND2_X1 U10710 ( .A1(n9271), .A2(n9270), .ZN(n9802) );
  INV_X1 U10711 ( .A(n9811), .ZN(n9273) );
  OAI22_X1 U10712 ( .A1(n9273), .A2(n9349), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9272), .ZN(n9274) );
  AOI21_X1 U10713 ( .B1(n9802), .B2(n9346), .A(n9274), .ZN(n9275) );
  OAI211_X1 U10714 ( .C1(n4724), .C2(n9283), .A(n9276), .B(n9275), .ZN(
        P1_U3229) );
  OAI21_X1 U10715 ( .B1(n9279), .B2(n9278), .A(n9277), .ZN(n9285) );
  OAI22_X1 U10716 ( .A1(n9370), .A2(n9301), .B1(n9280), .B2(n9300), .ZN(n9871)
         );
  AOI22_X1 U10717 ( .A1(n9871), .A2(n9346), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9282) );
  NAND2_X1 U10718 ( .A1(n9337), .A2(n9879), .ZN(n9281) );
  OAI211_X1 U10719 ( .C1(n10062), .C2(n9283), .A(n9282), .B(n9281), .ZN(n9284)
         );
  AOI21_X1 U10720 ( .B1(n9285), .B2(n9329), .A(n9284), .ZN(n9286) );
  INV_X1 U10721 ( .A(n9286), .ZN(P1_U3233) );
  XOR2_X1 U10722 ( .A(n9287), .B(n9288), .Z(n9296) );
  NAND2_X1 U10723 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10130)
         );
  NAND2_X1 U10724 ( .A1(n9346), .A2(n9290), .ZN(n9291) );
  OAI211_X1 U10725 ( .C1(n9349), .C2(n9292), .A(n10130), .B(n9291), .ZN(n9293)
         );
  AOI21_X1 U10726 ( .B1(n9294), .B2(n9351), .A(n9293), .ZN(n9295) );
  OAI21_X1 U10727 ( .B1(n9296), .B2(n9354), .A(n9295), .ZN(P1_U3234) );
  INV_X1 U10728 ( .A(n9187), .ZN(n9298) );
  AOI21_X1 U10729 ( .B1(n4584), .B2(n9299), .A(n9298), .ZN(n9305) );
  OAI22_X1 U10730 ( .A1(n9512), .A2(n9301), .B1(n9370), .B2(n9300), .ZN(n9836)
         );
  AOI22_X1 U10731 ( .A1(n9836), .A2(n9346), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3086), .ZN(n9302) );
  OAI21_X1 U10732 ( .B1(n9349), .B2(n9843), .A(n9302), .ZN(n9303) );
  AOI21_X1 U10733 ( .B1(n9842), .B2(n9351), .A(n9303), .ZN(n9304) );
  OAI21_X1 U10734 ( .B1(n9305), .B2(n9354), .A(n9304), .ZN(P1_U3235) );
  AOI21_X1 U10735 ( .B1(n9307), .B2(n9309), .A(n9306), .ZN(n9308) );
  AOI21_X1 U10736 ( .B1(n4507), .B2(n9309), .A(n9308), .ZN(n9314) );
  AOI22_X1 U10737 ( .A1(n9346), .A2(n9310), .B1(P1_REG3_REG_11__SCAN_IN), .B2(
        P1_U3086), .ZN(n9311) );
  OAI21_X1 U10738 ( .B1(n9349), .B2(n10183), .A(n9311), .ZN(n9312) );
  AOI21_X1 U10739 ( .B1(n10187), .B2(n9351), .A(n9312), .ZN(n9313) );
  OAI21_X1 U10740 ( .B1(n9314), .B2(n9354), .A(n9313), .ZN(P1_U3236) );
  INV_X1 U10741 ( .A(n9316), .ZN(n9318) );
  NAND2_X1 U10742 ( .A1(n9318), .A2(n9317), .ZN(n9319) );
  XNOR2_X1 U10743 ( .A(n9315), .B(n9319), .ZN(n9327) );
  AOI22_X1 U10744 ( .A1(n9629), .A2(n9321), .B1(n9631), .B2(n9320), .ZN(n9908)
         );
  OAI22_X1 U10745 ( .A1(n9323), .A2(n9908), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9322), .ZN(n9324) );
  AOI21_X1 U10746 ( .B1(n9912), .B2(n9337), .A(n9324), .ZN(n9326) );
  NAND2_X1 U10747 ( .A1(n9911), .A2(n9351), .ZN(n9325) );
  OAI211_X1 U10748 ( .C1(n9327), .C2(n9354), .A(n9326), .B(n9325), .ZN(
        P1_U3238) );
  AND3_X1 U10749 ( .A1(n7177), .A2(n5237), .A3(n9328), .ZN(n9330) );
  OAI21_X1 U10750 ( .B1(n4520), .B2(n9330), .A(n9329), .ZN(n9341) );
  INV_X1 U10751 ( .A(n9331), .ZN(n9332) );
  AOI21_X1 U10752 ( .B1(n9346), .B2(n9333), .A(n9332), .ZN(n9340) );
  NAND2_X1 U10753 ( .A1(n9351), .A2(n9334), .ZN(n9339) );
  INV_X1 U10754 ( .A(n9335), .ZN(n9336) );
  NAND2_X1 U10755 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  NAND4_X1 U10756 ( .A1(n9341), .A2(n9340), .A3(n9339), .A4(n9338), .ZN(
        P1_U3239) );
  AOI21_X1 U10757 ( .B1(n9344), .B2(n9343), .A(n9342), .ZN(n9355) );
  AOI22_X1 U10758 ( .A1(n9346), .A2(n9345), .B1(P1_REG3_REG_15__SCAN_IN), .B2(
        P1_U3086), .ZN(n9347) );
  OAI21_X1 U10759 ( .B1(n9349), .B2(n9348), .A(n9347), .ZN(n9350) );
  AOI21_X1 U10760 ( .B1(n9352), .B2(n9351), .A(n9350), .ZN(n9353) );
  OAI21_X1 U10761 ( .B1(n9355), .B2(n9354), .A(n9353), .ZN(P1_U3241) );
  NAND2_X1 U10762 ( .A1(n9359), .A2(n9358), .ZN(n10024) );
  NAND2_X1 U10763 ( .A1(n9360), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n9362) );
  NAND2_X1 U10764 ( .A1(n4614), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n9361) );
  OAI211_X1 U10765 ( .C1(n9364), .C2(n9363), .A(n9362), .B(n9361), .ZN(n9713)
         );
  NAND2_X1 U10766 ( .A1(n10024), .A2(n9713), .ZN(n9593) );
  NAND2_X1 U10767 ( .A1(n9528), .A2(n9520), .ZN(n9381) );
  NAND2_X1 U10768 ( .A1(n4473), .A2(n9801), .ZN(n9367) );
  NAND2_X1 U10769 ( .A1(n9784), .A2(n9367), .ZN(n9368) );
  NAND2_X1 U10770 ( .A1(n9368), .A2(n9514), .ZN(n9369) );
  NAND2_X1 U10771 ( .A1(n9519), .A2(n9369), .ZN(n9380) );
  INV_X1 U10772 ( .A(n9380), .ZN(n9377) );
  OR2_X1 U10773 ( .A1(n9861), .A2(n9370), .ZN(n9507) );
  INV_X1 U10774 ( .A(n9507), .ZN(n9374) );
  NAND2_X1 U10775 ( .A1(n9878), .A2(n9371), .ZN(n9417) );
  NAND2_X1 U10776 ( .A1(n9503), .A2(n9417), .ZN(n9508) );
  INV_X1 U10777 ( .A(n9508), .ZN(n9373) );
  AND2_X1 U10778 ( .A1(n9801), .A2(n9372), .ZN(n9506) );
  OAI211_X1 U10779 ( .C1(n9374), .C2(n9373), .A(n9514), .B(n9506), .ZN(n9376)
         );
  INV_X1 U10780 ( .A(n9517), .ZN(n9375) );
  AOI21_X1 U10781 ( .B1(n9377), .B2(n9376), .A(n9375), .ZN(n9378) );
  NOR2_X1 U10782 ( .A1(n9381), .A2(n9378), .ZN(n9379) );
  OR2_X1 U10783 ( .A1(n4491), .A2(n9379), .ZN(n9582) );
  NAND2_X1 U10784 ( .A1(n9507), .A2(n9416), .ZN(n9504) );
  OR3_X1 U10785 ( .A1(n9381), .A2(n9380), .A3(n9504), .ZN(n9580) );
  NAND2_X1 U10786 ( .A1(n9497), .A2(n9495), .ZN(n9539) );
  AND2_X1 U10787 ( .A1(n9484), .A2(n9382), .ZN(n9490) );
  NAND2_X1 U10788 ( .A1(n9494), .A2(n9486), .ZN(n9470) );
  INV_X1 U10789 ( .A(n9470), .ZN(n9399) );
  AOI21_X1 U10790 ( .B1(n9645), .B2(n6383), .A(n9535), .ZN(n9386) );
  NAND2_X1 U10791 ( .A1(n6380), .A2(n9383), .ZN(n9384) );
  AND4_X1 U10792 ( .A1(n9386), .A2(n9385), .A3(n9384), .A4(n9428), .ZN(n9387)
         );
  AND3_X1 U10793 ( .A1(n9387), .A2(n9440), .A3(n9435), .ZN(n9389) );
  OAI211_X1 U10794 ( .C1(n9390), .C2(n9389), .A(n9388), .B(n9461), .ZN(n9392)
         );
  NAND2_X1 U10795 ( .A1(n9464), .A2(n9457), .ZN(n9451) );
  INV_X1 U10796 ( .A(n9451), .ZN(n9391) );
  NAND2_X1 U10797 ( .A1(n9392), .A2(n9391), .ZN(n9394) );
  NAND2_X1 U10798 ( .A1(n9466), .A2(n9460), .ZN(n9453) );
  INV_X1 U10799 ( .A(n9453), .ZN(n9393) );
  NAND2_X1 U10800 ( .A1(n9394), .A2(n9393), .ZN(n9395) );
  NAND3_X1 U10801 ( .A1(n9395), .A2(n9487), .A3(n9463), .ZN(n9397) );
  NAND3_X1 U10802 ( .A1(n9489), .A2(n9397), .A3(n9396), .ZN(n9398) );
  NAND2_X1 U10803 ( .A1(n9399), .A2(n9398), .ZN(n9401) );
  INV_X1 U10804 ( .A(n9492), .ZN(n9400) );
  AOI21_X1 U10805 ( .B1(n9490), .B2(n9401), .A(n9400), .ZN(n9402) );
  AND2_X1 U10806 ( .A1(n9481), .A2(n9478), .ZN(n9564) );
  OAI21_X1 U10807 ( .B1(n9539), .B2(n9402), .A(n9564), .ZN(n9403) );
  NAND3_X1 U10808 ( .A1(n9403), .A2(n9497), .A3(n9496), .ZN(n9404) );
  AND2_X1 U10809 ( .A1(n9404), .A2(n9475), .ZN(n9406) );
  INV_X1 U10810 ( .A(n9518), .ZN(n9405) );
  NAND2_X1 U10811 ( .A1(n9528), .A2(n9405), .ZN(n9579) );
  OAI21_X1 U10812 ( .B1(n9580), .B2(n9406), .A(n9579), .ZN(n9407) );
  NOR2_X1 U10813 ( .A1(n9582), .A2(n9407), .ZN(n9411) );
  NAND2_X1 U10814 ( .A1(n9529), .A2(n4494), .ZN(n9584) );
  NAND2_X1 U10815 ( .A1(n9408), .A2(n5214), .ZN(n9410) );
  NAND2_X1 U10816 ( .A1(n5610), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n9409) );
  AND2_X2 U10817 ( .A1(n9410), .A2(n9409), .ZN(n10028) );
  NAND2_X1 U10818 ( .A1(n9720), .A2(n9412), .ZN(n9589) );
  OAI211_X1 U10819 ( .C1(n9411), .C2(n9584), .A(n9589), .B(n9588), .ZN(n9413)
         );
  OR2_X1 U10820 ( .A1(n9720), .A2(n9412), .ZN(n9577) );
  NAND2_X1 U10821 ( .A1(n9413), .A2(n9577), .ZN(n9414) );
  NAND2_X1 U10822 ( .A1(n9593), .A2(n9414), .ZN(n9415) );
  OR2_X1 U10823 ( .A1(n10024), .A2(n9713), .ZN(n9594) );
  NAND2_X1 U10824 ( .A1(n9415), .A2(n9594), .ZN(n9609) );
  AOI21_X1 U10825 ( .B1(n9417), .B2(n9892), .A(n9533), .ZN(n9420) );
  NAND2_X1 U10826 ( .A1(n9416), .A2(n9496), .ZN(n9419) );
  INV_X1 U10827 ( .A(n9533), .ZN(n9534) );
  NAND3_X1 U10828 ( .A1(n9417), .A2(n9629), .A3(n9534), .ZN(n9418) );
  OAI21_X1 U10829 ( .B1(n9420), .B2(n9419), .A(n9418), .ZN(n9502) );
  NAND2_X1 U10830 ( .A1(n9423), .A2(n9533), .ZN(n9424) );
  NAND3_X1 U10831 ( .A1(n9425), .A2(n9533), .A3(n9428), .ZN(n9426) );
  NAND2_X1 U10832 ( .A1(n9427), .A2(n9426), .ZN(n9437) );
  OAI21_X1 U10833 ( .B1(n9437), .B2(n4618), .A(n9429), .ZN(n9431) );
  INV_X1 U10834 ( .A(n9442), .ZN(n9430) );
  AOI21_X1 U10835 ( .B1(n9431), .B2(n9440), .A(n9430), .ZN(n9434) );
  OAI21_X1 U10836 ( .B1(n9434), .B2(n9433), .A(n9432), .ZN(n9446) );
  OAI21_X1 U10837 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9439) );
  MUX2_X1 U10838 ( .A(n9446), .B(n9445), .S(n9533), .Z(n9450) );
  MUX2_X1 U10839 ( .A(n9448), .B(n9447), .S(n9534), .Z(n9449) );
  NAND2_X1 U10840 ( .A1(n9450), .A2(n9449), .ZN(n9456) );
  NAND2_X1 U10841 ( .A1(n9456), .A2(n9458), .ZN(n9452) );
  AOI21_X1 U10842 ( .B1(n9452), .B2(n9461), .A(n9451), .ZN(n9454) );
  OAI21_X1 U10843 ( .B1(n9454), .B2(n9453), .A(n9463), .ZN(n9468) );
  NAND2_X1 U10844 ( .A1(n9456), .A2(n9455), .ZN(n9459) );
  NAND3_X1 U10845 ( .A1(n9459), .A2(n9458), .A3(n9457), .ZN(n9462) );
  NAND3_X1 U10846 ( .A1(n9462), .A2(n9461), .A3(n9460), .ZN(n9465) );
  NAND3_X1 U10847 ( .A1(n9465), .A2(n9464), .A3(n9463), .ZN(n9467) );
  NAND2_X1 U10848 ( .A1(n9485), .A2(n9487), .ZN(n9472) );
  NOR2_X1 U10849 ( .A1(n9469), .A2(n9488), .ZN(n9471) );
  AOI21_X1 U10850 ( .B1(n9472), .B2(n9471), .A(n9470), .ZN(n9474) );
  OAI21_X1 U10851 ( .B1(n9474), .B2(n9473), .A(n9492), .ZN(n9477) );
  NAND4_X1 U10852 ( .A1(n9475), .A2(n9533), .A3(n9478), .A4(n9481), .ZN(n9476)
         );
  AOI21_X1 U10853 ( .B1(n9477), .B2(n9484), .A(n9476), .ZN(n9500) );
  OR2_X1 U10854 ( .A1(n9497), .A2(n9533), .ZN(n9483) );
  NAND2_X1 U10855 ( .A1(n9478), .A2(n9534), .ZN(n9479) );
  NAND2_X1 U10856 ( .A1(n9481), .A2(n9479), .ZN(n9480) );
  OAI21_X1 U10857 ( .B1(n9481), .B2(n9533), .A(n9480), .ZN(n9482) );
  OAI211_X1 U10858 ( .C1(n9539), .C2(n9534), .A(n9483), .B(n9482), .ZN(n9499)
         );
  NAND3_X1 U10859 ( .A1(n9491), .A2(n9490), .A3(n9489), .ZN(n9493) );
  AND2_X1 U10860 ( .A1(n9495), .A2(n9534), .ZN(n9498) );
  OAI21_X1 U10861 ( .B1(n9509), .B2(n9504), .A(n9503), .ZN(n9505) );
  OAI21_X1 U10862 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9510) );
  OR3_X1 U10863 ( .A1(n9827), .A2(n9512), .A3(n9533), .ZN(n9513) );
  MUX2_X1 U10864 ( .A(n9514), .B(n9784), .S(n9533), .Z(n9515) );
  NAND2_X1 U10865 ( .A1(n9518), .A2(n9517), .ZN(n9524) );
  OR2_X1 U10866 ( .A1(n9524), .A2(n9519), .ZN(n9521) );
  AND2_X1 U10867 ( .A1(n9521), .A2(n9520), .ZN(n9525) );
  INV_X1 U10868 ( .A(n9525), .ZN(n9527) );
  MUX2_X1 U10869 ( .A(n9588), .B(n9529), .S(n9534), .Z(n9530) );
  NAND2_X1 U10870 ( .A1(n9531), .A2(n9530), .ZN(n9532) );
  NAND2_X1 U10871 ( .A1(n9713), .A2(n9619), .ZN(n9591) );
  OAI22_X1 U10872 ( .A1(n9599), .A2(n5851), .B1(n9534), .B2(n9594), .ZN(n9538)
         );
  INV_X1 U10873 ( .A(n9593), .ZN(n9536) );
  AOI21_X1 U10874 ( .B1(n9536), .B2(n9705), .A(n9535), .ZN(n9537) );
  INV_X1 U10875 ( .A(n9539), .ZN(n9565) );
  NOR2_X1 U10876 ( .A1(n9540), .A2(n9601), .ZN(n9543) );
  NOR2_X1 U10877 ( .A1(n9545), .A2(n9544), .ZN(n9549) );
  NAND4_X1 U10878 ( .A1(n9549), .A2(n9548), .A3(n9547), .A4(n9546), .ZN(n9550)
         );
  OR4_X1 U10879 ( .A1(n9553), .A2(n9552), .A3(n9551), .A4(n9550), .ZN(n9554)
         );
  NOR2_X1 U10880 ( .A1(n9555), .A2(n9554), .ZN(n9556) );
  NAND4_X1 U10881 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(n9560)
         );
  NOR2_X1 U10882 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  NAND4_X1 U10883 ( .A1(n9565), .A2(n9564), .A3(n9563), .A4(n9562), .ZN(n9566)
         );
  NOR2_X1 U10884 ( .A1(n9894), .A2(n9566), .ZN(n9567) );
  NAND4_X1 U10885 ( .A1(n9840), .A2(n9567), .A3(n9875), .A4(n9856), .ZN(n9569)
         );
  INV_X1 U10886 ( .A(n9800), .ZN(n9806) );
  OR3_X1 U10887 ( .A1(n9569), .A2(n9806), .A3(n9568), .ZN(n9572) );
  OR4_X1 U10888 ( .A1(n9572), .A2(n9571), .A3(n9771), .A4(n9570), .ZN(n9573)
         );
  NOR2_X1 U10889 ( .A1(n9574), .A2(n9573), .ZN(n9575) );
  AND4_X1 U10890 ( .A1(n9577), .A2(n9589), .A3(n9576), .A4(n9575), .ZN(n9578)
         );
  AND3_X1 U10891 ( .A1(n9594), .A2(n9578), .A3(n9593), .ZN(n9600) );
  INV_X1 U10892 ( .A(n9600), .ZN(n9598) );
  OAI21_X1 U10893 ( .B1(n9580), .B2(n4445), .A(n9579), .ZN(n9581) );
  NOR2_X1 U10894 ( .A1(n9582), .A2(n9581), .ZN(n9583) );
  OR2_X1 U10895 ( .A1(n9584), .A2(n9583), .ZN(n9587) );
  INV_X1 U10896 ( .A(n9713), .ZN(n9585) );
  NAND2_X1 U10897 ( .A1(n9720), .A2(n9585), .ZN(n9586) );
  NAND4_X1 U10898 ( .A1(n9589), .A2(n9588), .A3(n9587), .A4(n9586), .ZN(n9590)
         );
  OAI21_X1 U10899 ( .B1(n9591), .B2(n9720), .A(n9590), .ZN(n9592) );
  NAND2_X1 U10900 ( .A1(n9593), .A2(n9592), .ZN(n9596) );
  NAND3_X1 U10901 ( .A1(n9596), .A2(n9595), .A3(n9594), .ZN(n9597) );
  NAND2_X1 U10902 ( .A1(n9598), .A2(n9597), .ZN(n9604) );
  NAND2_X1 U10903 ( .A1(n9599), .A2(n5851), .ZN(n9602) );
  AOI21_X1 U10904 ( .B1(n9602), .B2(n9601), .A(n9600), .ZN(n9603) );
  NAND2_X1 U10905 ( .A1(n9609), .A2(n9705), .ZN(n9606) );
  NAND2_X1 U10906 ( .A1(n9611), .A2(n9610), .ZN(n9612) );
  NOR4_X1 U10907 ( .A1(n9614), .A2(n9613), .A3(n5856), .A4(n9612), .ZN(n9616)
         );
  OAI21_X1 U10908 ( .B1(n9617), .B2(n5851), .A(P1_B_REG_SCAN_IN), .ZN(n9615)
         );
  OAI22_X1 U10909 ( .A1(n9618), .A2(n9617), .B1(n9616), .B2(n9615), .ZN(
        P1_U3242) );
  MUX2_X1 U10910 ( .A(n9713), .B(P1_DATAO_REG_31__SCAN_IN), .S(n9646), .Z(
        P1_U3585) );
  MUX2_X1 U10911 ( .A(n9619), .B(P1_DATAO_REG_30__SCAN_IN), .S(n9646), .Z(
        P1_U3584) );
  MUX2_X1 U10912 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9620), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10913 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9621), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10914 ( .A(n9622), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9646), .Z(
        P1_U3580) );
  MUX2_X1 U10915 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9623), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10916 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9624), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10917 ( .A(n9625), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9646), .Z(
        P1_U3577) );
  MUX2_X1 U10918 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9626), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10919 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9627), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10920 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9628), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10921 ( .A(n9629), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9646), .Z(
        P1_U3573) );
  MUX2_X1 U10922 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9630), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10923 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9631), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10924 ( .A(n9632), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9646), .Z(
        P1_U3570) );
  MUX2_X1 U10925 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9633), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10926 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9634), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10927 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9635), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10928 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9636), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10929 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9637), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10930 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9638), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10931 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9639), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10932 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9640), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10933 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9641), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10934 ( .A(n9642), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9646), .Z(
        P1_U3560) );
  MUX2_X1 U10935 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9643), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10936 ( .A(n9644), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9646), .Z(
        P1_U3558) );
  MUX2_X1 U10937 ( .A(n6385), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9646), .Z(
        P1_U3557) );
  MUX2_X1 U10938 ( .A(n9645), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9646), .Z(
        P1_U3556) );
  MUX2_X1 U10939 ( .A(n9647), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9646), .Z(
        P1_U3554) );
  NAND2_X1 U10940 ( .A1(n10173), .A2(n9648), .ZN(n9650) );
  OAI211_X1 U10941 ( .C1(n9651), .C2(n10171), .A(n9650), .B(n9649), .ZN(n9652)
         );
  INV_X1 U10942 ( .A(n9652), .ZN(n9667) );
  MUX2_X1 U10943 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6596), .S(n9659), .Z(n9655)
         );
  INV_X1 U10944 ( .A(n9653), .ZN(n9654) );
  NAND2_X1 U10945 ( .A1(n9655), .A2(n9654), .ZN(n9657) );
  OAI211_X1 U10946 ( .C1(n9658), .C2(n9657), .A(n10158), .B(n9656), .ZN(n9666)
         );
  MUX2_X1 U10947 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6605), .S(n9659), .Z(n9660)
         );
  NAND3_X1 U10948 ( .A1(n9662), .A2(n9661), .A3(n9660), .ZN(n9663) );
  NAND3_X1 U10949 ( .A1(n10175), .A2(n9664), .A3(n9663), .ZN(n9665) );
  NAND4_X1 U10950 ( .A1(n9668), .A2(n9667), .A3(n9666), .A4(n9665), .ZN(
        P1_U3247) );
  OR3_X1 U10951 ( .A1(n9671), .A2(n9670), .A3(n9669), .ZN(n9672) );
  NAND3_X1 U10952 ( .A1(n9673), .A2(n10158), .A3(n9672), .ZN(n9685) );
  NOR2_X1 U10953 ( .A1(n9674), .A2(n9677), .ZN(n9675) );
  AOI211_X1 U10954 ( .C1(n10155), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n9676), .B(
        n9675), .ZN(n9684) );
  MUX2_X1 U10955 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6680), .S(n9677), .Z(n9678)
         );
  NAND3_X1 U10956 ( .A1(n9680), .A2(n9679), .A3(n9678), .ZN(n9681) );
  NAND3_X1 U10957 ( .A1(n10175), .A2(n9682), .A3(n9681), .ZN(n9683) );
  NAND3_X1 U10958 ( .A1(n9685), .A2(n9684), .A3(n9683), .ZN(P1_U3251) );
  OR2_X1 U10959 ( .A1(n9687), .A2(n9686), .ZN(n9691) );
  NAND2_X1 U10960 ( .A1(n9689), .A2(n9688), .ZN(n9690) );
  AND2_X1 U10961 ( .A1(n9691), .A2(n9690), .ZN(n10178) );
  XNOR2_X1 U10962 ( .A(n10170), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10177) );
  NAND2_X1 U10963 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  INV_X1 U10964 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9999) );
  OR2_X1 U10965 ( .A1(n10170), .A2(n9999), .ZN(n9692) );
  NAND2_X1 U10966 ( .A1(n10176), .A2(n9692), .ZN(n9694) );
  XNOR2_X1 U10967 ( .A(n9694), .B(n9693), .ZN(n9702) );
  NOR2_X1 U10968 ( .A1(n9696), .A2(n9695), .ZN(n10169) );
  NOR2_X1 U10969 ( .A1(n10169), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9698) );
  INV_X1 U10970 ( .A(n10169), .ZN(n9697) );
  OAI22_X1 U10971 ( .A1(n10170), .A2(n9698), .B1(n10166), .B2(n9697), .ZN(
        n9699) );
  XNOR2_X1 U10972 ( .A(n9699), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9704) );
  INV_X1 U10973 ( .A(n9704), .ZN(n9700) );
  AOI22_X1 U10974 ( .A1(n9702), .A2(n10175), .B1(n10158), .B2(n9700), .ZN(
        n9707) );
  NOR2_X1 U10975 ( .A1(n9702), .A2(n9701), .ZN(n9703) );
  AOI211_X1 U10976 ( .C1(n9704), .C2(n10158), .A(n10173), .B(n9703), .ZN(n9706) );
  MUX2_X1 U10977 ( .A(n9707), .B(n9706), .S(n9705), .Z(n9709) );
  NAND2_X1 U10978 ( .A1(P1_REG3_REG_19__SCAN_IN), .A2(P1_U3086), .ZN(n9708) );
  OAI211_X1 U10979 ( .C1(n7548), .C2(n10171), .A(n9709), .B(n9708), .ZN(
        P1_U3262) );
  XNOR2_X1 U10980 ( .A(n9718), .B(n10024), .ZN(n9710) );
  NOR2_X1 U10981 ( .A1(n9710), .A2(n9922), .ZN(n9937) );
  INV_X1 U10982 ( .A(n9711), .ZN(n9712) );
  AND2_X1 U10983 ( .A1(n9713), .A2(n9712), .ZN(n9940) );
  INV_X1 U10984 ( .A(n9940), .ZN(n9714) );
  OR2_X1 U10985 ( .A1(n4415), .A2(n9714), .ZN(n9721) );
  NAND2_X1 U10986 ( .A1(n4415), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9715) );
  OAI211_X1 U10987 ( .C1(n10024), .C2(n9927), .A(n9721), .B(n9715), .ZN(n9716)
         );
  AOI21_X1 U10988 ( .B1(n9937), .B2(n10189), .A(n9716), .ZN(n9717) );
  INV_X1 U10989 ( .A(n9717), .ZN(P1_U3263) );
  AOI211_X1 U10990 ( .C1(n9720), .C2(n9719), .A(n9922), .B(n9718), .ZN(n9941)
         );
  NAND2_X1 U10991 ( .A1(n4415), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9722) );
  OAI211_X1 U10992 ( .C1(n10028), .C2(n9927), .A(n9722), .B(n9721), .ZN(n9723)
         );
  AOI21_X1 U10993 ( .B1(n9941), .B2(n10189), .A(n9723), .ZN(n9724) );
  INV_X1 U10994 ( .A(n9724), .ZN(P1_U3264) );
  NAND2_X1 U10995 ( .A1(n9725), .A2(n9876), .ZN(n9733) );
  NAND2_X1 U10996 ( .A1(n10184), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n9727) );
  INV_X1 U10997 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n9726) );
  OAI22_X1 U10998 ( .A1(n9728), .A2(n9727), .B1(n9726), .B2(n9916), .ZN(n9731)
         );
  NOR2_X1 U10999 ( .A1(n9729), .A2(n9778), .ZN(n9730) );
  AOI211_X1 U11000 ( .C1(n10186), .C2(n6452), .A(n9731), .B(n9730), .ZN(n9732)
         );
  OAI211_X1 U11001 ( .C1(n9734), .C2(n4415), .A(n9733), .B(n9732), .ZN(
        P1_U3356) );
  XNOR2_X1 U11002 ( .A(n9735), .B(n9738), .ZN(n9737) );
  AOI21_X1 U11003 ( .B1(n9737), .B2(n9931), .A(n9736), .ZN(n9945) );
  AND2_X1 U11004 ( .A1(n9739), .A2(n9738), .ZN(n9740) );
  NOR2_X1 U11005 ( .A1(n9741), .A2(n9740), .ZN(n9947) );
  NAND2_X1 U11006 ( .A1(n9947), .A2(n9876), .ZN(n9749) );
  AND2_X1 U11007 ( .A1(n9742), .A2(n9757), .ZN(n9743) );
  OR3_X1 U11008 ( .A1(n4439), .A2(n9743), .A3(n9922), .ZN(n9944) );
  INV_X1 U11009 ( .A(n9944), .ZN(n9747) );
  AOI22_X1 U11010 ( .A1(n9744), .A2(n10184), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n4415), .ZN(n9745) );
  OAI21_X1 U11011 ( .B1(n10032), .B2(n9927), .A(n9745), .ZN(n9746) );
  AOI21_X1 U11012 ( .B1(n9747), .B2(n10189), .A(n9746), .ZN(n9748) );
  OAI211_X1 U11013 ( .C1(n4415), .C2(n9945), .A(n9749), .B(n9748), .ZN(
        P1_U3265) );
  XNOR2_X1 U11014 ( .A(n9750), .B(n9755), .ZN(n9751) );
  NAND2_X1 U11015 ( .A1(n9751), .A2(n9931), .ZN(n9754) );
  INV_X1 U11016 ( .A(n9752), .ZN(n9753) );
  INV_X1 U11017 ( .A(n9950), .ZN(n9765) );
  XNOR2_X1 U11018 ( .A(n9756), .B(n9755), .ZN(n9952) );
  NAND2_X1 U11019 ( .A1(n9952), .A2(n9876), .ZN(n9764) );
  INV_X1 U11020 ( .A(n9757), .ZN(n9758) );
  AOI211_X1 U11021 ( .C1(n9759), .C2(n9776), .A(n9922), .B(n9758), .ZN(n9951)
         );
  AOI22_X1 U11022 ( .A1(n9760), .A2(n10184), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n4415), .ZN(n9761) );
  OAI21_X1 U11023 ( .B1(n10035), .B2(n9927), .A(n9761), .ZN(n9762) );
  AOI21_X1 U11024 ( .B1(n9951), .B2(n10189), .A(n9762), .ZN(n9763) );
  OAI211_X1 U11025 ( .C1(n4415), .C2(n9765), .A(n9764), .B(n9763), .ZN(
        P1_U3266) );
  OAI21_X1 U11026 ( .B1(n9768), .B2(n9767), .A(n9766), .ZN(n9770) );
  AOI21_X1 U11027 ( .B1(n9770), .B2(n9931), .A(n9769), .ZN(n9956) );
  XNOR2_X1 U11028 ( .A(n9772), .B(n9771), .ZN(n9958) );
  NAND2_X1 U11029 ( .A1(n9958), .A2(n9876), .ZN(n9783) );
  INV_X1 U11030 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n9773) );
  OAI22_X1 U11031 ( .A1(n9775), .A2(n9774), .B1(n9773), .B2(n9916), .ZN(n9780)
         );
  OAI211_X1 U11032 ( .C1(n10039), .C2(n9791), .A(n9777), .B(n9776), .ZN(n9955)
         );
  NOR2_X1 U11033 ( .A1(n9955), .A2(n9778), .ZN(n9779) );
  AOI211_X1 U11034 ( .C1(n10186), .C2(n9781), .A(n9780), .B(n9779), .ZN(n9782)
         );
  OAI211_X1 U11035 ( .C1(n4415), .C2(n9956), .A(n9783), .B(n9782), .ZN(
        P1_U3267) );
  NAND2_X1 U11036 ( .A1(n9799), .A2(n9784), .ZN(n9785) );
  XNOR2_X1 U11037 ( .A(n9785), .B(n9789), .ZN(n9788) );
  INV_X1 U11038 ( .A(n9786), .ZN(n9787) );
  OAI21_X1 U11039 ( .B1(n9788), .B2(n9906), .A(n9787), .ZN(n9961) );
  INV_X1 U11040 ( .A(n9961), .ZN(n9798) );
  XNOR2_X1 U11041 ( .A(n9790), .B(n9789), .ZN(n9963) );
  NAND2_X1 U11042 ( .A1(n9963), .A2(n9876), .ZN(n9797) );
  AOI211_X1 U11043 ( .C1(n9792), .C2(n9808), .A(n9922), .B(n9791), .ZN(n9962)
         );
  AOI22_X1 U11044 ( .A1(n9793), .A2(n10184), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n4415), .ZN(n9794) );
  OAI21_X1 U11045 ( .B1(n10043), .B2(n9927), .A(n9794), .ZN(n9795) );
  AOI21_X1 U11046 ( .B1(n9962), .B2(n10189), .A(n9795), .ZN(n9796) );
  OAI211_X1 U11047 ( .C1(n4415), .C2(n9798), .A(n9797), .B(n9796), .ZN(
        P1_U3268) );
  NAND2_X1 U11048 ( .A1(n9799), .A2(n9931), .ZN(n9805) );
  AOI21_X1 U11049 ( .B1(n9801), .B2(n9817), .A(n9800), .ZN(n9804) );
  INV_X1 U11050 ( .A(n9802), .ZN(n9803) );
  OAI21_X1 U11051 ( .B1(n9805), .B2(n9804), .A(n9803), .ZN(n9966) );
  INV_X1 U11052 ( .A(n9966), .ZN(n9816) );
  XNOR2_X1 U11053 ( .A(n9807), .B(n9806), .ZN(n9968) );
  NAND2_X1 U11054 ( .A1(n9968), .A2(n9876), .ZN(n9815) );
  INV_X1 U11055 ( .A(n9808), .ZN(n9809) );
  AOI211_X1 U11056 ( .C1(n9810), .C2(n9825), .A(n9922), .B(n9809), .ZN(n9967)
         );
  AOI22_X1 U11057 ( .A1(n9811), .A2(n10184), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n4415), .ZN(n9812) );
  OAI21_X1 U11058 ( .B1(n4724), .B2(n9927), .A(n9812), .ZN(n9813) );
  AOI21_X1 U11059 ( .B1(n9967), .B2(n10189), .A(n9813), .ZN(n9814) );
  OAI211_X1 U11060 ( .C1(n4415), .C2(n9816), .A(n9815), .B(n9814), .ZN(
        P1_U3269) );
  OAI21_X1 U11061 ( .B1(n9823), .B2(n9818), .A(n9817), .ZN(n9819) );
  NAND2_X1 U11062 ( .A1(n9819), .A2(n9931), .ZN(n9822) );
  INV_X1 U11063 ( .A(n9820), .ZN(n9821) );
  NAND2_X1 U11064 ( .A1(n9822), .A2(n9821), .ZN(n9971) );
  INV_X1 U11065 ( .A(n9971), .ZN(n9834) );
  XNOR2_X1 U11066 ( .A(n9824), .B(n9823), .ZN(n9973) );
  NAND2_X1 U11067 ( .A1(n9973), .A2(n9876), .ZN(n9833) );
  INV_X1 U11068 ( .A(n9825), .ZN(n9826) );
  INV_X1 U11069 ( .A(n9828), .ZN(n9829) );
  AOI22_X1 U11070 ( .A1(n9829), .A2(n10184), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n4415), .ZN(n9830) );
  OAI21_X1 U11071 ( .B1(n10050), .B2(n9927), .A(n9830), .ZN(n9831) );
  AOI21_X1 U11072 ( .B1(n9972), .B2(n10189), .A(n9831), .ZN(n9832) );
  OAI211_X1 U11073 ( .C1(n4415), .C2(n9834), .A(n9833), .B(n9832), .ZN(
        P1_U3270) );
  XOR2_X1 U11074 ( .A(n9840), .B(n9835), .Z(n9838) );
  INV_X1 U11075 ( .A(n9836), .ZN(n9837) );
  OAI21_X1 U11076 ( .B1(n9838), .B2(n9906), .A(n9837), .ZN(n9976) );
  INV_X1 U11077 ( .A(n9976), .ZN(n9849) );
  XOR2_X1 U11078 ( .A(n9840), .B(n9839), .Z(n9978) );
  NAND2_X1 U11079 ( .A1(n9978), .A2(n9876), .ZN(n9848) );
  AOI211_X1 U11080 ( .C1(n9842), .C2(n9859), .A(n9922), .B(n9841), .ZN(n9977)
         );
  INV_X1 U11081 ( .A(n9842), .ZN(n10054) );
  INV_X1 U11082 ( .A(n9843), .ZN(n9844) );
  AOI22_X1 U11083 ( .A1(n9844), .A2(n10184), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n4415), .ZN(n9845) );
  OAI21_X1 U11084 ( .B1(n10054), .B2(n9927), .A(n9845), .ZN(n9846) );
  AOI21_X1 U11085 ( .B1(n9977), .B2(n10189), .A(n9846), .ZN(n9847) );
  OAI211_X1 U11086 ( .C1(n4415), .C2(n9849), .A(n9848), .B(n9847), .ZN(
        P1_U3271) );
  OAI21_X1 U11087 ( .B1(n9851), .B2(n9856), .A(n9850), .ZN(n9852) );
  NAND2_X1 U11088 ( .A1(n9852), .A2(n9931), .ZN(n9855) );
  INV_X1 U11089 ( .A(n9853), .ZN(n9854) );
  NAND2_X1 U11090 ( .A1(n9855), .A2(n9854), .ZN(n9981) );
  INV_X1 U11091 ( .A(n9981), .ZN(n9868) );
  XNOR2_X1 U11092 ( .A(n9857), .B(n9856), .ZN(n9983) );
  NAND2_X1 U11093 ( .A1(n9983), .A2(n9876), .ZN(n9867) );
  INV_X1 U11094 ( .A(n9859), .ZN(n9860) );
  AOI211_X1 U11095 ( .C1(n9861), .C2(n9877), .A(n9922), .B(n9860), .ZN(n9982)
         );
  INV_X1 U11096 ( .A(n9861), .ZN(n10058) );
  INV_X1 U11097 ( .A(n9862), .ZN(n9863) );
  AOI22_X1 U11098 ( .A1(n9863), .A2(n10184), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n4415), .ZN(n9864) );
  OAI21_X1 U11099 ( .B1(n10058), .B2(n9927), .A(n9864), .ZN(n9865) );
  AOI21_X1 U11100 ( .B1(n9982), .B2(n10189), .A(n9865), .ZN(n9866) );
  OAI211_X1 U11101 ( .C1(n4415), .C2(n9868), .A(n9867), .B(n9866), .ZN(
        P1_U3272) );
  INV_X1 U11102 ( .A(n9875), .ZN(n9869) );
  XNOR2_X1 U11103 ( .A(n4445), .B(n9869), .ZN(n9870) );
  NAND2_X1 U11104 ( .A1(n9870), .A2(n9931), .ZN(n9873) );
  INV_X1 U11105 ( .A(n9871), .ZN(n9872) );
  NAND2_X1 U11106 ( .A1(n9873), .A2(n9872), .ZN(n9986) );
  INV_X1 U11107 ( .A(n9986), .ZN(n9884) );
  XOR2_X1 U11108 ( .A(n9875), .B(n9874), .Z(n9988) );
  NAND2_X1 U11109 ( .A1(n9988), .A2(n9876), .ZN(n9883) );
  AOI211_X1 U11110 ( .C1(n9878), .C2(n9886), .A(n9922), .B(n9858), .ZN(n9987)
         );
  AOI22_X1 U11111 ( .A1(n4415), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9879), .B2(
        n10184), .ZN(n9880) );
  OAI21_X1 U11112 ( .B1(n10062), .B2(n9927), .A(n9880), .ZN(n9881) );
  AOI21_X1 U11113 ( .B1(n9987), .B2(n10189), .A(n9881), .ZN(n9882) );
  OAI211_X1 U11114 ( .C1(n4415), .C2(n9884), .A(n9883), .B(n9882), .ZN(
        P1_U3273) );
  XOR2_X1 U11115 ( .A(n9894), .B(n9885), .Z(n9995) );
  INV_X1 U11116 ( .A(n9910), .ZN(n9888) );
  INV_X1 U11117 ( .A(n9886), .ZN(n9887) );
  AOI211_X1 U11118 ( .C1(n9992), .C2(n9888), .A(n9922), .B(n9887), .ZN(n9991)
         );
  INV_X1 U11119 ( .A(n9889), .ZN(n9890) );
  AOI22_X1 U11120 ( .A1(n4415), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9890), .B2(
        n10184), .ZN(n9891) );
  OAI21_X1 U11121 ( .B1(n9892), .B2(n9927), .A(n9891), .ZN(n9901) );
  INV_X1 U11122 ( .A(n9893), .ZN(n9897) );
  INV_X1 U11123 ( .A(n9894), .ZN(n9896) );
  OAI21_X1 U11124 ( .B1(n9897), .B2(n9896), .A(n9895), .ZN(n9899) );
  AOI21_X1 U11125 ( .B1(n9899), .B2(n9931), .A(n9898), .ZN(n9994) );
  NOR2_X1 U11126 ( .A1(n9994), .A2(n4415), .ZN(n9900) );
  AOI211_X1 U11127 ( .C1(n9991), .C2(n10189), .A(n9901), .B(n9900), .ZN(n9902)
         );
  OAI21_X1 U11128 ( .B1(n9995), .B2(n9936), .A(n9902), .ZN(P1_U3274) );
  XNOR2_X1 U11129 ( .A(n9903), .B(n9904), .ZN(n9998) );
  INV_X1 U11130 ( .A(n9998), .ZN(n9918) );
  XNOR2_X1 U11131 ( .A(n9905), .B(n9904), .ZN(n9907) );
  OR2_X1 U11132 ( .A1(n9907), .A2(n9906), .ZN(n9909) );
  NAND2_X1 U11133 ( .A1(n9909), .A2(n9908), .ZN(n9996) );
  INV_X1 U11134 ( .A(n9911), .ZN(n10068) );
  AOI211_X1 U11135 ( .C1(n9911), .C2(n9920), .A(n9922), .B(n9910), .ZN(n9997)
         );
  NAND2_X1 U11136 ( .A1(n9997), .A2(n10189), .ZN(n9914) );
  AOI22_X1 U11137 ( .A1(n4415), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9912), .B2(
        n10184), .ZN(n9913) );
  OAI211_X1 U11138 ( .C1(n10068), .C2(n9927), .A(n9914), .B(n9913), .ZN(n9915)
         );
  AOI21_X1 U11139 ( .B1(n9916), .B2(n9996), .A(n9915), .ZN(n9917) );
  OAI21_X1 U11140 ( .B1(n9918), .B2(n9936), .A(n9917), .ZN(P1_U3275) );
  XOR2_X1 U11141 ( .A(n9919), .B(n9929), .Z(n10006) );
  INV_X1 U11142 ( .A(n9920), .ZN(n9921) );
  AOI211_X1 U11143 ( .C1(n10003), .C2(n9923), .A(n9922), .B(n9921), .ZN(n10002) );
  INV_X1 U11144 ( .A(n9924), .ZN(n9925) );
  AOI22_X1 U11145 ( .A1(n4415), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9925), .B2(
        n10184), .ZN(n9926) );
  OAI21_X1 U11146 ( .B1(n6455), .B2(n9927), .A(n9926), .ZN(n9934) );
  XOR2_X1 U11147 ( .A(n9929), .B(n9928), .Z(n9932) );
  AOI21_X1 U11148 ( .B1(n9932), .B2(n9931), .A(n9930), .ZN(n10005) );
  NOR2_X1 U11149 ( .A1(n10005), .A2(n4415), .ZN(n9933) );
  AOI211_X1 U11150 ( .C1(n10002), .C2(n10189), .A(n9934), .B(n9933), .ZN(n9935) );
  OAI21_X1 U11151 ( .B1(n10006), .B2(n9936), .A(n9935), .ZN(P1_U3276) );
  INV_X1 U11152 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9938) );
  NOR2_X1 U11153 ( .A1(n9937), .A2(n9940), .ZN(n10021) );
  MUX2_X1 U11154 ( .A(n9938), .B(n10021), .S(n10223), .Z(n9939) );
  OAI21_X1 U11155 ( .B1(n10024), .B2(n10001), .A(n9939), .ZN(P1_U3553) );
  NOR2_X1 U11156 ( .A1(n9941), .A2(n9940), .ZN(n10025) );
  MUX2_X1 U11157 ( .A(n9942), .B(n10025), .S(n10223), .Z(n9943) );
  OAI21_X1 U11158 ( .B1(n10028), .B2(n10001), .A(n9943), .ZN(P1_U3552) );
  NAND2_X1 U11159 ( .A1(n9945), .A2(n9944), .ZN(n9946) );
  AOI21_X1 U11160 ( .B1(n9947), .B2(n10217), .A(n9946), .ZN(n10029) );
  MUX2_X1 U11161 ( .A(n9948), .B(n10029), .S(n10223), .Z(n9949) );
  OAI21_X1 U11162 ( .B1(n10032), .B2(n10001), .A(n9949), .ZN(P1_U3550) );
  MUX2_X1 U11163 ( .A(n9953), .B(n10033), .S(n10223), .Z(n9954) );
  OAI21_X1 U11164 ( .B1(n10035), .B2(n10001), .A(n9954), .ZN(P1_U3549) );
  NAND2_X1 U11165 ( .A1(n9956), .A2(n9955), .ZN(n9957) );
  AOI21_X1 U11166 ( .B1(n9958), .B2(n10217), .A(n9957), .ZN(n10036) );
  MUX2_X1 U11167 ( .A(n9959), .B(n10036), .S(n10223), .Z(n9960) );
  OAI21_X1 U11168 ( .B1(n10039), .B2(n10001), .A(n9960), .ZN(P1_U3548) );
  INV_X1 U11169 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9964) );
  AOI211_X1 U11170 ( .C1(n9963), .C2(n10217), .A(n9962), .B(n9961), .ZN(n10040) );
  MUX2_X1 U11171 ( .A(n9964), .B(n10040), .S(n10223), .Z(n9965) );
  OAI21_X1 U11172 ( .B1(n10043), .B2(n10001), .A(n9965), .ZN(P1_U3547) );
  AOI211_X1 U11173 ( .C1(n9968), .C2(n10217), .A(n9967), .B(n9966), .ZN(n10044) );
  MUX2_X1 U11174 ( .A(n9969), .B(n10044), .S(n10223), .Z(n9970) );
  OAI21_X1 U11175 ( .B1(n4724), .B2(n10001), .A(n9970), .ZN(P1_U3546) );
  AOI211_X1 U11176 ( .C1(n9973), .C2(n10217), .A(n9972), .B(n9971), .ZN(n10047) );
  MUX2_X1 U11177 ( .A(n9974), .B(n10047), .S(n10223), .Z(n9975) );
  OAI21_X1 U11178 ( .B1(n10050), .B2(n10001), .A(n9975), .ZN(P1_U3545) );
  AOI211_X1 U11179 ( .C1(n9978), .C2(n10217), .A(n9977), .B(n9976), .ZN(n10051) );
  MUX2_X1 U11180 ( .A(n9979), .B(n10051), .S(n10223), .Z(n9980) );
  OAI21_X1 U11181 ( .B1(n10054), .B2(n10001), .A(n9980), .ZN(P1_U3544) );
  AOI211_X1 U11182 ( .C1(n9983), .C2(n10217), .A(n9982), .B(n9981), .ZN(n10055) );
  MUX2_X1 U11183 ( .A(n9984), .B(n10055), .S(n10223), .Z(n9985) );
  OAI21_X1 U11184 ( .B1(n10058), .B2(n10001), .A(n9985), .ZN(P1_U3543) );
  INV_X1 U11185 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n9989) );
  AOI211_X1 U11186 ( .C1(n9988), .C2(n10217), .A(n9987), .B(n9986), .ZN(n10059) );
  MUX2_X1 U11187 ( .A(n9989), .B(n10059), .S(n10223), .Z(n9990) );
  OAI21_X1 U11188 ( .B1(n10062), .B2(n10001), .A(n9990), .ZN(P1_U3542) );
  AOI21_X1 U11189 ( .B1(n10205), .B2(n9992), .A(n9991), .ZN(n9993) );
  OAI211_X1 U11190 ( .C1(n9995), .C2(n10018), .A(n9994), .B(n9993), .ZN(n10063) );
  MUX2_X1 U11191 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10063), .S(n10223), .Z(
        P1_U3541) );
  AOI211_X1 U11192 ( .C1(n9998), .C2(n10217), .A(n9997), .B(n9996), .ZN(n10064) );
  MUX2_X1 U11193 ( .A(n9999), .B(n10064), .S(n10223), .Z(n10000) );
  OAI21_X1 U11194 ( .B1(n10068), .B2(n10001), .A(n10000), .ZN(P1_U3540) );
  AOI21_X1 U11195 ( .B1(n10205), .B2(n10003), .A(n10002), .ZN(n10004) );
  OAI211_X1 U11196 ( .C1(n10006), .C2(n10018), .A(n10005), .B(n10004), .ZN(
        n10069) );
  MUX2_X1 U11197 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10069), .S(n10223), .Z(
        P1_U3539) );
  NAND3_X1 U11198 ( .A1(n10008), .A2(n10007), .A3(n10217), .ZN(n10013) );
  AOI211_X1 U11199 ( .C1(n10205), .C2(n10011), .A(n10010), .B(n10009), .ZN(
        n10012) );
  NAND2_X1 U11200 ( .A1(n10013), .A2(n10012), .ZN(n10070) );
  MUX2_X1 U11201 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10070), .S(n10223), .Z(
        P1_U3538) );
  AOI21_X1 U11202 ( .B1(n10205), .B2(n10015), .A(n10014), .ZN(n10016) );
  OAI211_X1 U11203 ( .C1(n10019), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10071) );
  MUX2_X1 U11204 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10071), .S(n10223), .Z(
        P1_U3536) );
  MUX2_X1 U11205 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n10020), .S(n10223), .Z(
        P1_U3522) );
  INV_X1 U11206 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10022) );
  MUX2_X1 U11207 ( .A(n10022), .B(n10021), .S(n10220), .Z(n10023) );
  OAI21_X1 U11208 ( .B1(n10024), .B2(n10067), .A(n10023), .ZN(P1_U3521) );
  MUX2_X1 U11209 ( .A(n10026), .B(n10025), .S(n10220), .Z(n10027) );
  OAI21_X1 U11210 ( .B1(n10028), .B2(n10067), .A(n10027), .ZN(P1_U3520) );
  MUX2_X1 U11211 ( .A(n10030), .B(n10029), .S(n10220), .Z(n10031) );
  OAI21_X1 U11212 ( .B1(n10032), .B2(n10067), .A(n10031), .ZN(P1_U3518) );
  INV_X1 U11213 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n10034) );
  INV_X1 U11214 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10037) );
  MUX2_X1 U11215 ( .A(n10037), .B(n10036), .S(n10220), .Z(n10038) );
  OAI21_X1 U11216 ( .B1(n10039), .B2(n10067), .A(n10038), .ZN(P1_U3516) );
  MUX2_X1 U11217 ( .A(n10041), .B(n10040), .S(n10220), .Z(n10042) );
  OAI21_X1 U11218 ( .B1(n10043), .B2(n10067), .A(n10042), .ZN(P1_U3515) );
  INV_X1 U11219 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10045) );
  MUX2_X1 U11220 ( .A(n10045), .B(n10044), .S(n10220), .Z(n10046) );
  OAI21_X1 U11221 ( .B1(n4724), .B2(n10067), .A(n10046), .ZN(P1_U3514) );
  INV_X1 U11222 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10048) );
  MUX2_X1 U11223 ( .A(n10048), .B(n10047), .S(n10220), .Z(n10049) );
  OAI21_X1 U11224 ( .B1(n10050), .B2(n10067), .A(n10049), .ZN(P1_U3513) );
  INV_X1 U11225 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n10052) );
  MUX2_X1 U11226 ( .A(n10052), .B(n10051), .S(n10220), .Z(n10053) );
  OAI21_X1 U11227 ( .B1(n10054), .B2(n10067), .A(n10053), .ZN(P1_U3512) );
  INV_X1 U11228 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n10056) );
  MUX2_X1 U11229 ( .A(n10056), .B(n10055), .S(n10220), .Z(n10057) );
  OAI21_X1 U11230 ( .B1(n10058), .B2(n10067), .A(n10057), .ZN(P1_U3511) );
  INV_X1 U11231 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10060) );
  MUX2_X1 U11232 ( .A(n10060), .B(n10059), .S(n10220), .Z(n10061) );
  OAI21_X1 U11233 ( .B1(n10062), .B2(n10067), .A(n10061), .ZN(P1_U3510) );
  MUX2_X1 U11234 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10063), .S(n10220), .Z(
        P1_U3509) );
  INV_X1 U11235 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10065) );
  MUX2_X1 U11236 ( .A(n10065), .B(n10064), .S(n10220), .Z(n10066) );
  OAI21_X1 U11237 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(P1_U3507) );
  MUX2_X1 U11238 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10069), .S(n10220), .Z(
        P1_U3504) );
  MUX2_X1 U11239 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10070), .S(n10220), .Z(
        P1_U3501) );
  MUX2_X1 U11240 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10071), .S(n10220), .Z(
        P1_U3495) );
  MUX2_X1 U11241 ( .A(n10072), .B(P1_D_REG_1__SCAN_IN), .S(n10202), .Z(
        P1_U3440) );
  MUX2_X1 U11242 ( .A(n10073), .B(P1_D_REG_0__SCAN_IN), .S(n10202), .Z(
        P1_U3439) );
  NOR4_X1 U11243 ( .A1(n10075), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n10074), .ZN(n10076) );
  AOI21_X1 U11244 ( .B1(n10082), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n10076), 
        .ZN(n10077) );
  OAI21_X1 U11245 ( .B1(n10078), .B2(n10085), .A(n10077), .ZN(P1_U3324) );
  AOI22_X1 U11246 ( .A1(n10079), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10082), .ZN(n10080) );
  OAI21_X1 U11247 ( .B1(n10081), .B2(n10085), .A(n10080), .ZN(P1_U3325) );
  AOI22_X1 U11248 ( .A1(n10083), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10082), .ZN(n10084) );
  OAI21_X1 U11249 ( .B1(n6415), .B2(n10085), .A(n10084), .ZN(P1_U3326) );
  INV_X1 U11250 ( .A(n10086), .ZN(n10087) );
  MUX2_X1 U11251 ( .A(n10087), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U11252 ( .A(n10088), .ZN(n10089) );
  NOR2_X1 U11253 ( .A1(n10090), .A2(n10089), .ZN(n10093) );
  AOI21_X1 U11254 ( .B1(n10093), .B2(P2_U3893), .A(n10270), .ZN(n10102) );
  AOI21_X1 U11255 ( .B1(n4452), .B2(n10098), .A(n10097), .ZN(n10099) );
  OR2_X1 U11256 ( .A1(n10099), .A2(n10302), .ZN(n10100) );
  AOI21_X1 U11257 ( .B1(n10105), .B2(n10104), .A(n10103), .ZN(n10117) );
  AND2_X1 U11258 ( .A1(n10107), .A2(n10106), .ZN(n10108) );
  OAI21_X1 U11259 ( .B1(n10109), .B2(n10108), .A(n10175), .ZN(n10115) );
  AOI21_X1 U11260 ( .B1(n10155), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10110), .ZN(
        n10114) );
  INV_X1 U11261 ( .A(n10111), .ZN(n10112) );
  NAND2_X1 U11262 ( .A1(n10173), .A2(n10112), .ZN(n10113) );
  AND3_X1 U11263 ( .A1(n10115), .A2(n10114), .A3(n10113), .ZN(n10116) );
  OAI21_X1 U11264 ( .B1(n10117), .B2(n10182), .A(n10116), .ZN(P1_U3252) );
  XNOR2_X1 U11265 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11266 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U11267 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n10155), .B1(
        P1_REG3_REG_11__SCAN_IN), .B2(P1_U3086), .ZN(n10129) );
  INV_X1 U11268 ( .A(n10118), .ZN(n10119) );
  NAND2_X1 U11269 ( .A1(n10173), .A2(n10119), .ZN(n10128) );
  OAI211_X1 U11270 ( .C1(n10122), .C2(n10121), .A(n10120), .B(n10175), .ZN(
        n10127) );
  OAI211_X1 U11271 ( .C1(n10125), .C2(n10124), .A(n10123), .B(n10158), .ZN(
        n10126) );
  NAND4_X1 U11272 ( .A1(n10129), .A2(n10128), .A3(n10127), .A4(n10126), .ZN(
        P1_U3254) );
  OAI21_X1 U11273 ( .B1(n10171), .B2(n10131), .A(n10130), .ZN(n10132) );
  AOI21_X1 U11274 ( .B1(n10133), .B2(n10173), .A(n10132), .ZN(n10142) );
  OAI211_X1 U11275 ( .C1(n10136), .C2(n10135), .A(n10158), .B(n10134), .ZN(
        n10141) );
  OAI211_X1 U11276 ( .C1(n10139), .C2(n10138), .A(n10175), .B(n10137), .ZN(
        n10140) );
  NAND3_X1 U11277 ( .A1(n10142), .A2(n10141), .A3(n10140), .ZN(P1_U3256) );
  OAI21_X1 U11278 ( .B1(n10171), .B2(n7523), .A(n10143), .ZN(n10144) );
  AOI21_X1 U11279 ( .B1(n10145), .B2(n10173), .A(n10144), .ZN(n10154) );
  OAI211_X1 U11280 ( .C1(n10148), .C2(n10147), .A(n10158), .B(n10146), .ZN(
        n10153) );
  OAI211_X1 U11281 ( .C1(n10151), .C2(n10150), .A(n10175), .B(n10149), .ZN(
        n10152) );
  NAND3_X1 U11282 ( .A1(n10154), .A2(n10153), .A3(n10152), .ZN(P1_U3257) );
  AOI22_X1 U11283 ( .A1(n10155), .A2(P1_ADDR_REG_15__SCAN_IN), .B1(
        P1_REG3_REG_15__SCAN_IN), .B2(P1_U3086), .ZN(n10165) );
  NAND2_X1 U11284 ( .A1(n10173), .A2(n10156), .ZN(n10164) );
  OAI211_X1 U11285 ( .C1(P1_REG2_REG_15__SCAN_IN), .C2(n10159), .A(n10158), 
        .B(n10157), .ZN(n10163) );
  OAI211_X1 U11286 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n10161), .A(n10175), 
        .B(n10160), .ZN(n10162) );
  NAND4_X1 U11287 ( .A1(n10165), .A2(n10164), .A3(n10163), .A4(n10162), .ZN(
        P1_U3258) );
  MUX2_X1 U11288 ( .A(n10166), .B(P1_REG2_REG_18__SCAN_IN), .S(n10170), .Z(
        n10168) );
  NAND2_X1 U11289 ( .A1(n10168), .A2(n10169), .ZN(n10167) );
  OAI21_X1 U11290 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(n10181) );
  INV_X1 U11291 ( .A(n10170), .ZN(n10174) );
  OAI22_X1 U11292 ( .A1(n10171), .A2(n10390), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9322), .ZN(n10172) );
  AOI21_X1 U11293 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10180) );
  OAI211_X1 U11294 ( .C1(n10178), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10179) );
  OAI211_X1 U11295 ( .C1(n10182), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        P1_U3261) );
  INV_X1 U11296 ( .A(n10183), .ZN(n10185) );
  AOI222_X1 U11297 ( .A1(n10187), .A2(n10186), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n4415), .C1(n10185), .C2(n10184), .ZN(n10193) );
  AOI22_X1 U11298 ( .A1(n10191), .A2(n10190), .B1(n10189), .B2(n10188), .ZN(
        n10192) );
  OAI211_X1 U11299 ( .C1(n4415), .C2(n10194), .A(n10193), .B(n10192), .ZN(
        P1_U3282) );
  AND2_X1 U11300 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10202), .ZN(P1_U3294) );
  AND2_X1 U11301 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10202), .ZN(P1_U3295) );
  NOR2_X1 U11302 ( .A1(n10201), .A2(n10195), .ZN(P1_U3296) );
  AND2_X1 U11303 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10202), .ZN(P1_U3297) );
  NOR2_X1 U11304 ( .A1(n10201), .A2(n10196), .ZN(P1_U3298) );
  AND2_X1 U11305 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10202), .ZN(P1_U3299) );
  AND2_X1 U11306 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10202), .ZN(P1_U3300) );
  AND2_X1 U11307 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10202), .ZN(P1_U3301) );
  AND2_X1 U11308 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10202), .ZN(P1_U3302) );
  AND2_X1 U11309 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10202), .ZN(P1_U3303) );
  AND2_X1 U11310 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10202), .ZN(P1_U3304) );
  AND2_X1 U11311 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10202), .ZN(P1_U3305) );
  AND2_X1 U11312 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10202), .ZN(P1_U3306) );
  AND2_X1 U11313 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10202), .ZN(P1_U3307) );
  AND2_X1 U11314 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10202), .ZN(P1_U3308) );
  AND2_X1 U11315 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10202), .ZN(P1_U3309) );
  AND2_X1 U11316 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10202), .ZN(P1_U3310) );
  NOR2_X1 U11317 ( .A1(n10201), .A2(n10197), .ZN(P1_U3311) );
  AND2_X1 U11318 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10202), .ZN(P1_U3312) );
  AND2_X1 U11319 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10202), .ZN(P1_U3313) );
  AND2_X1 U11320 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10202), .ZN(P1_U3314) );
  NOR2_X1 U11321 ( .A1(n10201), .A2(n10198), .ZN(P1_U3315) );
  NOR2_X1 U11322 ( .A1(n10201), .A2(n10199), .ZN(P1_U3316) );
  AND2_X1 U11323 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10202), .ZN(P1_U3317) );
  AND2_X1 U11324 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10202), .ZN(P1_U3318) );
  NOR2_X1 U11325 ( .A1(n10201), .A2(n10200), .ZN(P1_U3319) );
  AND2_X1 U11326 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10202), .ZN(P1_U3320) );
  AND2_X1 U11327 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10202), .ZN(P1_U3321) );
  AND2_X1 U11328 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10202), .ZN(P1_U3322) );
  AND2_X1 U11329 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10202), .ZN(P1_U3323) );
  AOI21_X1 U11330 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(n10206) );
  OAI211_X1 U11331 ( .C1(n10209), .C2(n10208), .A(n10207), .B(n10206), .ZN(
        n10210) );
  INV_X1 U11332 ( .A(n10210), .ZN(n10221) );
  AOI22_X1 U11333 ( .A1(n10220), .A2(n10221), .B1(n5279), .B2(n10218), .ZN(
        P1_U3474) );
  OAI21_X1 U11334 ( .B1(n10213), .B2(n10212), .A(n10211), .ZN(n10215) );
  AOI211_X1 U11335 ( .C1(n10217), .C2(n10216), .A(n10215), .B(n10214), .ZN(
        n10222) );
  INV_X1 U11336 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U11337 ( .A1(n10220), .A2(n10222), .B1(n10219), .B2(n10218), .ZN(
        P1_U3480) );
  AOI22_X1 U11338 ( .A1(n10223), .A2(n10221), .B1(n6628), .B2(n6496), .ZN(
        P1_U3529) );
  AOI22_X1 U11339 ( .A1(n10223), .A2(n10222), .B1(n8990), .B2(n6496), .ZN(
        P1_U3531) );
  OAI21_X1 U11340 ( .B1(n10226), .B2(n10225), .A(n10224), .ZN(n10227) );
  AOI22_X1 U11341 ( .A1(n10228), .A2(n10227), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(P2_U3151), .ZN(n10235) );
  OAI21_X1 U11342 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(n10232) );
  NAND2_X1 U11343 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  OAI211_X1 U11344 ( .C1(n10284), .C2(n5959), .A(n10235), .B(n10234), .ZN(
        n10236) );
  INV_X1 U11345 ( .A(n10236), .ZN(n10241) );
  XOR2_X1 U11346 ( .A(n10238), .B(n10237), .Z(n10239) );
  NAND2_X1 U11347 ( .A1(n10239), .A2(n10298), .ZN(n10240) );
  OAI211_X1 U11348 ( .C1(n10242), .C2(n10283), .A(n10241), .B(n10240), .ZN(
        P2_U3184) );
  AOI21_X1 U11349 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(n10246) );
  NOR2_X1 U11350 ( .A1(n10246), .A2(n10293), .ZN(n10253) );
  AOI21_X1 U11351 ( .B1(n5042), .B2(n10248), .A(n10247), .ZN(n10251) );
  INV_X1 U11352 ( .A(n10249), .ZN(n10250) );
  OAI21_X1 U11353 ( .B1(n10251), .B2(n10302), .A(n10250), .ZN(n10252) );
  AOI211_X1 U11354 ( .C1(n10270), .C2(n10254), .A(n10253), .B(n10252), .ZN(
        n10260) );
  OAI21_X1 U11355 ( .B1(n10257), .B2(n10256), .A(n10255), .ZN(n10258) );
  NAND2_X1 U11356 ( .A1(n10258), .A2(n10298), .ZN(n10259) );
  OAI211_X1 U11357 ( .C1(n10261), .C2(n10283), .A(n10260), .B(n10259), .ZN(
        P2_U3188) );
  AOI21_X1 U11358 ( .B1(n10264), .B2(n10263), .A(n10262), .ZN(n10273) );
  AOI21_X1 U11359 ( .B1(n10378), .B2(n10266), .A(n10265), .ZN(n10267) );
  OR2_X1 U11360 ( .A1(n10267), .A2(n10293), .ZN(n10272) );
  AOI21_X1 U11361 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(n10271) );
  OAI211_X1 U11362 ( .C1(n10273), .C2(n10302), .A(n10272), .B(n10271), .ZN(
        n10274) );
  INV_X1 U11363 ( .A(n10274), .ZN(n10280) );
  OAI21_X1 U11364 ( .B1(n10277), .B2(n10276), .A(n10275), .ZN(n10278) );
  NAND2_X1 U11365 ( .A1(n10278), .A2(n10298), .ZN(n10279) );
  OAI211_X1 U11366 ( .C1(n10283), .C2(n10281), .A(n10280), .B(n10279), .ZN(
        P2_U3189) );
  INV_X1 U11367 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10307) );
  INV_X1 U11368 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10282) );
  OAI22_X1 U11369 ( .A1(n10285), .A2(n10284), .B1(n10283), .B2(n10282), .ZN(
        n10286) );
  INV_X1 U11370 ( .A(n10286), .ZN(n10306) );
  AOI21_X1 U11371 ( .B1(n10289), .B2(n10288), .A(n10287), .ZN(n10303) );
  AOI21_X1 U11372 ( .B1(n10292), .B2(n10291), .A(n10290), .ZN(n10294) );
  OR2_X1 U11373 ( .A1(n10294), .A2(n10293), .ZN(n10301) );
  OAI21_X1 U11374 ( .B1(n10297), .B2(n10296), .A(n10295), .ZN(n10299) );
  NAND2_X1 U11375 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  OAI211_X1 U11376 ( .C1(n10303), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10304) );
  INV_X1 U11377 ( .A(n10304), .ZN(n10305) );
  OAI211_X1 U11378 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10307), .A(n10306), .B(
        n10305), .ZN(P2_U3199) );
  INV_X1 U11379 ( .A(n10308), .ZN(n10311) );
  OAI21_X1 U11380 ( .B1(n10311), .B2(n10310), .A(n10309), .ZN(n10316) );
  AOI222_X1 U11381 ( .A1(n10317), .A2(n10316), .B1(n10315), .B2(n10314), .C1(
        n10313), .C2(n10312), .ZN(n10318) );
  OAI21_X1 U11382 ( .B1(n10317), .B2(n4704), .A(n10318), .ZN(P2_U3224) );
  OAI22_X1 U11383 ( .A1(n10320), .A2(n10361), .B1(n10319), .B2(n10359), .ZN(
        n10322) );
  NOR2_X1 U11384 ( .A1(n10322), .A2(n10321), .ZN(n10369) );
  INV_X1 U11385 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U11386 ( .A1(n10367), .A2(n10369), .B1(n10323), .B2(n10365), .ZN(
        P2_U3393) );
  AOI22_X1 U11387 ( .A1(n10326), .A2(n6278), .B1(n10325), .B2(n10324), .ZN(
        n10327) );
  NAND2_X1 U11388 ( .A1(n10328), .A2(n10327), .ZN(n10370) );
  OAI22_X1 U11389 ( .A1(n10365), .A2(n10370), .B1(P2_REG0_REG_2__SCAN_IN), 
        .B2(n10367), .ZN(n10329) );
  INV_X1 U11390 ( .A(n10329), .ZN(P2_U3396) );
  INV_X1 U11391 ( .A(n10330), .ZN(n10334) );
  OAI22_X1 U11392 ( .A1(n10332), .A2(n10353), .B1(n10331), .B2(n10359), .ZN(
        n10333) );
  NOR2_X1 U11393 ( .A1(n10334), .A2(n10333), .ZN(n10373) );
  INV_X1 U11394 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10335) );
  AOI22_X1 U11395 ( .A1(n10367), .A2(n10373), .B1(n10335), .B2(n10365), .ZN(
        P2_U3399) );
  OR2_X1 U11396 ( .A1(n10336), .A2(n10353), .ZN(n10339) );
  OR2_X1 U11397 ( .A1(n10337), .A2(n10359), .ZN(n10338) );
  INV_X1 U11398 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10341) );
  AOI22_X1 U11399 ( .A1(n10367), .A2(n10375), .B1(n10341), .B2(n10365), .ZN(
        P2_U3402) );
  OAI22_X1 U11400 ( .A1(n10343), .A2(n10353), .B1(n10342), .B2(n10359), .ZN(
        n10345) );
  NOR2_X1 U11401 ( .A1(n10345), .A2(n10344), .ZN(n10377) );
  INV_X1 U11402 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10346) );
  AOI22_X1 U11403 ( .A1(n10367), .A2(n10377), .B1(n10346), .B2(n10365), .ZN(
        P2_U3408) );
  INV_X1 U11404 ( .A(n10347), .ZN(n10349) );
  OAI22_X1 U11405 ( .A1(n10349), .A2(n10361), .B1(n10348), .B2(n10359), .ZN(
        n10350) );
  NOR2_X1 U11406 ( .A1(n10351), .A2(n10350), .ZN(n10379) );
  AOI22_X1 U11407 ( .A1(n10367), .A2(n10379), .B1(n9015), .B2(n10365), .ZN(
        P2_U3411) );
  OAI22_X1 U11408 ( .A1(n10354), .A2(n10353), .B1(n10352), .B2(n10359), .ZN(
        n10355) );
  NOR2_X1 U11409 ( .A1(n10356), .A2(n10355), .ZN(n10381) );
  INV_X1 U11410 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U11411 ( .A1(n10367), .A2(n10381), .B1(n10357), .B2(n10365), .ZN(
        P2_U3414) );
  INV_X1 U11412 ( .A(n10358), .ZN(n10362) );
  OAI22_X1 U11413 ( .A1(n10362), .A2(n10361), .B1(n10360), .B2(n10359), .ZN(
        n10363) );
  NOR2_X1 U11414 ( .A1(n10364), .A2(n10363), .ZN(n10383) );
  INV_X1 U11415 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U11416 ( .A1(n10367), .A2(n10383), .B1(n10366), .B2(n10365), .ZN(
        P2_U3420) );
  AOI22_X1 U11417 ( .A1(n10384), .A2(n10369), .B1(n10368), .B2(n6377), .ZN(
        P2_U3460) );
  OAI22_X1 U11418 ( .A1(n6377), .A2(n10370), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n10384), .ZN(n10371) );
  INV_X1 U11419 ( .A(n10371), .ZN(P2_U3461) );
  AOI22_X1 U11420 ( .A1(n10384), .A2(n10373), .B1(n10372), .B2(n6377), .ZN(
        P2_U3462) );
  AOI22_X1 U11421 ( .A1(n10384), .A2(n10375), .B1(n10374), .B2(n6377), .ZN(
        P2_U3463) );
  AOI22_X1 U11422 ( .A1(n10384), .A2(n10377), .B1(n10376), .B2(n6377), .ZN(
        P2_U3465) );
  AOI22_X1 U11423 ( .A1(n10384), .A2(n10379), .B1(n10378), .B2(n6377), .ZN(
        P2_U3466) );
  AOI22_X1 U11424 ( .A1(n10384), .A2(n10381), .B1(n10380), .B2(n6377), .ZN(
        P2_U3467) );
  AOI22_X1 U11425 ( .A1(n10384), .A2(n10383), .B1(n10382), .B2(n6377), .ZN(
        P2_U3469) );
  NOR2_X1 U11426 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  XOR2_X1 U11427 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10387), .Z(ADD_1068_U5) );
  XOR2_X1 U11428 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI21_X1 U11429 ( .B1(n10390), .B2(n10389), .A(n10388), .ZN(n10391) );
  XNOR2_X1 U11430 ( .A(n10391), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(ADD_1068_U55)
         );
  OAI21_X1 U11431 ( .B1(n10394), .B2(n10393), .A(n10392), .ZN(ADD_1068_U56) );
  OAI21_X1 U11432 ( .B1(n10397), .B2(n10396), .A(n10395), .ZN(n10399) );
  XNOR2_X1 U11433 ( .A(n10399), .B(n10398), .ZN(ADD_1068_U57) );
  AOI21_X1 U11434 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10400), .ZN(n10402) );
  XNOR2_X1 U11435 ( .A(n10402), .B(n10401), .ZN(ADD_1068_U58) );
  OAI21_X1 U11436 ( .B1(n10405), .B2(n10404), .A(n10403), .ZN(ADD_1068_U59) );
  OAI21_X1 U11437 ( .B1(n10408), .B2(n10407), .A(n10406), .ZN(ADD_1068_U60) );
  OAI21_X1 U11438 ( .B1(n10411), .B2(n10410), .A(n10409), .ZN(ADD_1068_U61) );
  AOI21_X1 U11439 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(ADD_1068_U62) );
  OAI21_X1 U11440 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10419) );
  XNOR2_X1 U11441 ( .A(n10419), .B(n10418), .ZN(ADD_1068_U63) );
  XOR2_X1 U11442 ( .A(n10420), .B(P1_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11443 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  XOR2_X1 U11444 ( .A(n10423), .B(P1_ADDR_REG_5__SCAN_IN), .Z(ADD_1068_U51) );
  XOR2_X1 U11445 ( .A(n10424), .B(P2_ADDR_REG_9__SCAN_IN), .Z(ADD_1068_U47) );
  XOR2_X1 U11446 ( .A(n10426), .B(n10425), .Z(ADD_1068_U49) );
  XOR2_X1 U11447 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10427), .Z(ADD_1068_U48) );
  XOR2_X1 U11448 ( .A(n10429), .B(n10428), .Z(ADD_1068_U54) );
  XOR2_X1 U11449 ( .A(n10431), .B(n10430), .Z(ADD_1068_U53) );
  XNOR2_X1 U11450 ( .A(n10433), .B(n10432), .ZN(ADD_1068_U52) );
  CLKBUF_X1 U4918 ( .A(n5994), .Z(n4414) );
  INV_X2 U4944 ( .A(n5387), .ZN(n9364) );
  CLKBUF_X1 U4922 ( .A(n5202), .Z(n5743) );
  CLKBUF_X1 U4924 ( .A(n5994), .Z(n4413) );
  CLKBUF_X1 U4929 ( .A(n5221), .Z(n9360) );
  NAND2_X2 U4940 ( .A1(n10079), .A2(n10083), .ZN(n5129) );
  NAND2_X1 U4947 ( .A1(n4930), .A2(n4928), .ZN(n8656) );
  CLKBUF_X1 U4949 ( .A(n9356), .Z(n4525) );
endmodule

