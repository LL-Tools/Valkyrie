

module b20_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4278, n4279, n4280, n4281, n4282, n4283, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10367;

  OR2_X1 U4784 ( .A1(n9739), .A2(n4390), .ZN(n5853) );
  INV_X1 U4785 ( .A(n10227), .ZN(n9973) );
  OR2_X1 U4786 ( .A1(n10202), .A2(n10201), .ZN(n10204) );
  NAND2_X1 U4787 ( .A1(n9811), .A2(n10083), .ZN(n9786) );
  INV_X1 U4788 ( .A(n9733), .ZN(n10075) );
  XNOR2_X1 U4789 ( .A(n5937), .B(n5936), .ZN(n10123) );
  NAND2_X1 U4790 ( .A1(n8295), .A2(n8296), .ZN(n8331) );
  NAND2_X1 U4791 ( .A1(n8939), .A2(n8938), .ZN(n8937) );
  NOR2_X1 U4792 ( .A1(n8342), .A2(n8343), .ZN(n8341) );
  OR2_X1 U4793 ( .A1(n7309), .A2(n7308), .ZN(n4888) );
  NAND2_X1 U4794 ( .A1(n7994), .A2(n9551), .ZN(n8250) );
  NAND2_X1 U4795 ( .A1(n5968), .A2(n6090), .ZN(n9904) );
  OR2_X1 U4796 ( .A1(n7282), .A2(n7283), .ZN(n4890) );
  NAND2_X1 U4797 ( .A1(n7891), .A2(n7896), .ZN(n7995) );
  NAND2_X1 U4798 ( .A1(n6916), .A2(n6785), .ZN(n6918) );
  NAND2_X1 U4799 ( .A1(n5502), .A2(n5501), .ZN(n10051) );
  CLKBUF_X2 U4800 ( .A(n6364), .Z(n4288) );
  AOI21_X1 U4801 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7676), .A(n7674), .ZN(
        n7664) );
  BUF_X1 U4803 ( .A(n6193), .Z(n6364) );
  CLKBUF_X1 U4804 ( .A(n5593), .Z(n4670) );
  INV_X2 U4805 ( .A(n6185), .ZN(n6419) );
  INV_X1 U4806 ( .A(n8515), .ZN(n4756) );
  NAND3_X1 U4807 ( .A1(n7143), .A2(n6166), .A3(n9968), .ZN(n6381) );
  AND4_X1 U4808 ( .A1(n5291), .A2(n5290), .A3(n5289), .A4(n5288), .ZN(n7736)
         );
  NAND2_X1 U4809 ( .A1(n7499), .A2(n4758), .ZN(n7059) );
  NOR2_X1 U4810 ( .A1(n5463), .A2(n8748), .ZN(n5483) );
  CLKBUF_X1 U4812 ( .A(n6760), .Z(n4300) );
  XNOR2_X1 U4813 ( .A(n5297), .B(n5294), .ZN(n7168) );
  NAND2_X1 U4814 ( .A1(n5277), .A2(n5318), .ZN(n5297) );
  NAND2_X1 U4815 ( .A1(n6622), .A2(n6623), .ZN(n7050) );
  BUF_X1 U4816 ( .A(n6760), .Z(n4301) );
  NAND2_X1 U4817 ( .A1(n5244), .A2(n7524), .ZN(n5247) );
  OR2_X1 U4818 ( .A1(n4292), .A2(n5234), .ZN(n5235) );
  BUF_X2 U4819 ( .A(n5751), .Z(n4290) );
  CLKBUF_X2 U4820 ( .A(n7156), .Z(n5035) );
  AND4_X1 U4821 ( .A1(n6542), .A2(n6538), .A3(n4429), .A4(n6533), .ZN(n4335)
         );
  XNOR2_X1 U4822 ( .A(n5207), .B(SI_2_), .ZN(n4514) );
  NAND4_X1 U4823 ( .A1(n5167), .A2(n5169), .A3(n5170), .A4(n5168), .ZN(n5478)
         );
  NAND4_X1 U4824 ( .A1(n4283), .A2(n5172), .A3(n5171), .A4(n5279), .ZN(n5173)
         );
  INV_X1 U4825 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5586) );
  OAI21_X2 U4826 ( .B1(n5640), .B2(n4704), .A(n5037), .ZN(n5683) );
  NOR2_X2 U4828 ( .A1(n5548), .A2(n5547), .ZN(n5565) );
  INV_X2 U4829 ( .A(n9778), .ZN(n4698) );
  NAND2_X2 U4830 ( .A1(n6918), .A2(n6917), .ZN(n9346) );
  OAI21_X1 U4831 ( .B1(n7586), .B2(n6796), .A(n6795), .ZN(n4279) );
  BUF_X1 U4833 ( .A(n9256), .Z(n4281) );
  OAI21_X1 U4834 ( .B1(n7586), .B2(n6796), .A(n6795), .ZN(n7923) );
  OAI21_X1 U4835 ( .B1(n9218), .B2(n6927), .A(n6926), .ZN(n9206) );
  OAI22_X1 U4836 ( .A1(n8351), .A2(n6886), .B1(n9257), .B2(n8357), .ZN(n9256)
         );
  OAI21_X1 U4837 ( .B1(n6652), .B2(n7175), .A(n8937), .ZN(n4282) );
  OAI21_X1 U4838 ( .B1(n6652), .B2(n7175), .A(n8937), .ZN(n7635) );
  XNOR2_X1 U4840 ( .A(n5241), .B(n4588), .ZN(n7153) );
  NOR2_X2 U4841 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n4283) );
  NAND2_X1 U4843 ( .A1(n5498), .A2(n10367), .ZN(n5863) );
  NAND2_X1 U4845 ( .A1(n5529), .A2(n5528), .ZN(n4286) );
  NOR2_X1 U4846 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5191) );
  INV_X1 U4847 ( .A(n6788), .ZN(n6760) );
  OR2_X1 U4848 ( .A1(n6800), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6810) );
  INV_X1 U4849 ( .A(n6381), .ZN(n6345) );
  OR2_X1 U4850 ( .A1(n10145), .A2(n4829), .ZN(n4828) );
  INV_X1 U4851 ( .A(n8934), .ZN(n7369) );
  NAND2_X1 U4852 ( .A1(n7078), .A2(n8099), .ZN(n7329) );
  AOI22_X1 U4853 ( .A1(n8999), .A2(n8998), .B1(n6663), .B2(n6866), .ZN(n9016)
         );
  OR2_X1 U4854 ( .A1(n8514), .A2(n8509), .ZN(n9120) );
  NAND2_X1 U4855 ( .A1(n8428), .A2(n8439), .ZN(n8426) );
  INV_X1 U4856 ( .A(n4667), .ZN(n5788) );
  AOI21_X1 U4857 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n7268), .A(n8341), .ZN(
        n10147) );
  NOR2_X1 U4858 ( .A1(n10178), .A2(n10177), .ZN(n10176) );
  NAND2_X1 U4859 ( .A1(n6167), .A2(n7856), .ZN(n9968) );
  INV_X1 U4860 ( .A(n7744), .ZN(n5969) );
  XNOR2_X1 U4861 ( .A(n8652), .B(n8650), .ZN(n8883) );
  NAND2_X1 U4862 ( .A1(n4434), .A2(n7557), .ZN(n7795) );
  AND2_X1 U4863 ( .A1(n4890), .A2(n4889), .ZN(n7309) );
  INV_X1 U4864 ( .A(n6623), .ZN(n7043) );
  OAI211_X1 U4865 ( .C1(n6145), .C2(n6144), .A(n6152), .B(n6143), .ZN(n6150)
         );
  AND2_X1 U4866 ( .A1(n4646), .A2(n4645), .ZN(n4321) );
  AOI21_X1 U4867 ( .B1(n6150), .B2(n6149), .A(n4803), .ZN(n4805) );
  AND2_X2 U4868 ( .A1(n5482), .A2(n5481), .ZN(n5832) );
  AND2_X2 U4869 ( .A1(n4420), .A2(n7833), .ZN(n4327) );
  AOI22_X2 U4870 ( .A1(n8967), .A2(n8966), .B1(n8965), .B2(n6660), .ZN(n8972)
         );
  NAND3_X2 U4871 ( .A1(n6485), .A2(n5194), .A3(n5195), .ZN(n5198) );
  NOR2_X2 U4872 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6553) );
  NAND2_X2 U4873 ( .A1(n8601), .A2(n8600), .ZN(n8857) );
  AND3_X4 U4874 ( .A1(n4436), .A2(n4335), .A3(n4435), .ZN(n6521) );
  INV_X4 U4875 ( .A(n7690), .ZN(n10239) );
  NOR2_X2 U4876 ( .A1(n7709), .A2(n7708), .ZN(n7711) );
  NAND2_X4 U4877 ( .A1(n5592), .A2(n5591), .ZN(n9871) );
  AND2_X2 U4878 ( .A1(n5588), .A2(n5587), .ZN(n5592) );
  NAND2_X2 U4879 ( .A1(n4458), .A2(n4457), .ZN(n7690) );
  NAND2_X4 U4880 ( .A1(n5305), .A2(n5304), .ZN(n10260) );
  INV_X2 U4881 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8679) );
  NAND2_X1 U4883 ( .A1(n8110), .A2(n9871), .ZN(n5884) );
  NAND2_X2 U4884 ( .A1(n8011), .A2(n6841), .ZN(n6845) );
  NAND2_X2 U4885 ( .A1(n7821), .A2(n6824), .ZN(n8011) );
  OAI222_X1 U4887 ( .A1(n5881), .A2(P1_U3086), .B1(n10134), .B2(n8590), .C1(
        n8589), .C2(n10128), .ZN(P1_U3331) );
  XNOR2_X2 U4888 ( .A(n5861), .B(n5860), .ZN(n5881) );
  NAND2_X2 U4889 ( .A1(n7884), .A2(n7888), .ZN(n5406) );
  NAND2_X2 U4890 ( .A1(n4455), .A2(n4978), .ZN(n7884) );
  NAND2_X2 U4891 ( .A1(n4587), .A2(n7757), .ZN(n6036) );
  OAI211_X4 U4892 ( .C1(n5248), .C2(n7524), .A(n5247), .B(n5246), .ZN(n7744)
         );
  AOI21_X1 U4893 ( .B1(n8840), .B2(n8841), .A(n4376), .ZN(n8900) );
  NAND2_X1 U4894 ( .A1(n4699), .A2(n4698), .ZN(n6121) );
  INV_X1 U4895 ( .A(n9173), .ZN(n8886) );
  OAI21_X1 U4896 ( .B1(n6045), .B2(n6044), .A(n6043), .ZN(n6046) );
  NAND2_X1 U4897 ( .A1(n5462), .A2(n5461), .ZN(n5470) );
  INV_X2 U4898 ( .A(n9971), .ZN(n4287) );
  BUF_X2 U4899 ( .A(n6177), .Z(n6379) );
  AND4_X1 U4902 ( .A1(n5363), .A2(n5362), .A3(n5361), .A4(n5360), .ZN(n8264)
         );
  AND4_X1 U4903 ( .A1(n6832), .A2(n6831), .A3(n6830), .A4(n6829), .ZN(n8103)
         );
  AND4_X1 U4904 ( .A1(n5314), .A2(n5313), .A3(n5312), .A4(n5311), .ZN(n7756)
         );
  INV_X2 U4905 ( .A(n9871), .ZN(n7856) );
  BUF_X4 U4906 ( .A(n5278), .Z(n5744) );
  BUF_X2 U4907 ( .A(n6785), .Z(n7010) );
  NAND2_X2 U4908 ( .A1(n4893), .A2(P1_U3086), .ZN(n10128) );
  XNOR2_X1 U4910 ( .A(n5212), .B(SI_3_), .ZN(n5211) );
  INV_X2 U4911 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6509) );
  AOI21_X1 U4912 ( .B1(n9645), .B2(n9646), .A(n9662), .ZN(n4686) );
  NOR2_X1 U4913 ( .A1(n6439), .A2(n6438), .ZN(n6440) );
  OAI21_X1 U4914 ( .B1(n9587), .B2(n4634), .A(n9589), .ZN(n4633) );
  OR2_X2 U4915 ( .A1(n7125), .A2(n7124), .ZN(n9739) );
  OR2_X1 U4916 ( .A1(n10080), .A2(n10289), .ZN(n4593) );
  NAND2_X1 U4917 ( .A1(n9620), .A2(n9618), .ZN(n9617) );
  XNOR2_X1 U4918 ( .A(n9759), .B(n9763), .ZN(n9989) );
  NAND2_X1 U4919 ( .A1(n9553), .A2(n9554), .ZN(n9552) );
  AOI21_X1 U4920 ( .B1(n9109), .B2(n9295), .A(n9108), .ZN(n9395) );
  OAI22_X1 U4921 ( .A1(n8900), .A2(n8901), .B1(n8620), .B2(n9133), .ZN(n8622)
         );
  OAI21_X1 U4922 ( .B1(n9785), .B2(n5716), .A(n4306), .ZN(n4616) );
  NAND2_X1 U4923 ( .A1(n4433), .A2(n8617), .ZN(n8840) );
  NAND2_X1 U4924 ( .A1(n6341), .A2(n6340), .ZN(n9511) );
  NAND2_X1 U4925 ( .A1(n4513), .A2(n9059), .ZN(n9033) );
  AND2_X1 U4926 ( .A1(n10075), .A2(n9664), .ZN(n6139) );
  OAI21_X1 U4927 ( .B1(n9519), .B2(n6325), .A(n6324), .ZN(n9598) );
  NAND2_X1 U4928 ( .A1(n6640), .A2(n9038), .ZN(n9059) );
  INV_X1 U4929 ( .A(n9499), .ZN(n9501) );
  NAND2_X1 U4930 ( .A1(n4843), .A2(n4842), .ZN(n4841) );
  AOI21_X1 U4931 ( .B1(n8632), .B2(n6785), .A(n4417), .ZN(n8801) );
  NAND2_X1 U4932 ( .A1(n9605), .A2(n9606), .ZN(n9604) );
  INV_X1 U4933 ( .A(n9120), .ZN(n9122) );
  XNOR2_X1 U4934 ( .A(n5933), .B(n5932), .ZN(n8632) );
  NAND2_X1 U4935 ( .A1(n4500), .A2(n4499), .ZN(n9023) );
  NAND2_X1 U4936 ( .A1(n7023), .A2(n7022), .ZN(n9391) );
  OAI21_X1 U4937 ( .B1(n5900), .B2(n5899), .A(n5898), .ZN(n5933) );
  AOI21_X1 U4938 ( .B1(n4986), .B2(n4984), .A(n4357), .ZN(n4983) );
  NAND2_X1 U4939 ( .A1(n5746), .A2(n5745), .ZN(n9987) );
  AND2_X1 U4940 ( .A1(n6971), .A2(n4840), .ZN(n4835) );
  NAND2_X1 U4941 ( .A1(n4502), .A2(n9002), .ZN(n9021) );
  NAND2_X1 U4942 ( .A1(n6254), .A2(n6257), .ZN(n5018) );
  AND2_X1 U4943 ( .A1(n4987), .A2(n5681), .ZN(n4986) );
  OR2_X1 U4944 ( .A1(n8659), .A2(n8886), .ZN(n5145) );
  NAND2_X1 U4945 ( .A1(n5023), .A2(n5724), .ZN(n9780) );
  XNOR2_X1 U4946 ( .A(n10009), .B(n9860), .ZN(n9846) );
  OR2_X1 U4947 ( .A1(n9421), .A2(n9173), .ZN(n4583) );
  AND2_X1 U4948 ( .A1(n8493), .A2(n8492), .ZN(n9197) );
  NAND2_X1 U4949 ( .A1(n6975), .A2(n6974), .ZN(n9415) );
  NAND3_X1 U4950 ( .A1(n5143), .A2(n5834), .A3(n6069), .ZN(n8373) );
  AND2_X1 U4951 ( .A1(n5697), .A2(n5696), .ZN(n9823) );
  AND2_X1 U4952 ( .A1(n6082), .A2(n6081), .ZN(n9946) );
  NAND2_X1 U4953 ( .A1(n6931), .A2(n6930), .ZN(n9443) );
  INV_X1 U4954 ( .A(n6074), .ZN(n6081) );
  NAND2_X1 U4955 ( .A1(n6939), .A2(n6938), .ZN(n9339) );
  NAND2_X1 U4956 ( .A1(n8245), .A2(n5831), .ZN(n9957) );
  NAND2_X1 U4957 ( .A1(n5546), .A2(n5545), .ZN(n10039) );
  INV_X1 U4958 ( .A(n6075), .ZN(n6082) );
  AND2_X1 U4959 ( .A1(n5707), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5725) );
  XNOR2_X1 U4960 ( .A(n4907), .B(n5574), .ZN(n6916) );
  OR2_X1 U4961 ( .A1(n10051), .A2(n9963), .ZN(n6073) );
  NAND2_X1 U4962 ( .A1(n4456), .A2(n5340), .ZN(n7932) );
  INV_X1 U4963 ( .A(n10108), .ZN(n9939) );
  INV_X1 U4964 ( .A(n6067), .ZN(n6069) );
  NAND2_X1 U4965 ( .A1(n6889), .A2(n6888), .ZN(n9464) );
  INV_X1 U4966 ( .A(n5830), .ZN(n8247) );
  INV_X1 U4967 ( .A(n5010), .ZN(n5009) );
  AND2_X2 U4968 ( .A1(n5518), .A2(n5517), .ZN(n10108) );
  NAND2_X1 U4969 ( .A1(n6897), .A2(n6896), .ZN(n9457) );
  AND2_X1 U4970 ( .A1(n5990), .A2(n9956), .ZN(n5830) );
  NOR2_X1 U4971 ( .A1(n8115), .A2(n6063), .ZN(n5828) );
  AOI21_X1 U4972 ( .B1(n4856), .B2(n4852), .A(n4368), .ZN(n4850) );
  NAND2_X1 U4973 ( .A1(n6878), .A2(n6877), .ZN(n8357) );
  NAND2_X1 U4974 ( .A1(n7343), .A2(n7342), .ZN(n8920) );
  AND2_X1 U4975 ( .A1(n8116), .A2(n5984), .ZN(n7989) );
  NAND2_X1 U4976 ( .A1(n5029), .A2(n5030), .ZN(n5532) );
  NAND2_X1 U4977 ( .A1(n4658), .A2(n7785), .ZN(n7784) );
  INV_X1 U4978 ( .A(n8370), .ZN(n10065) );
  AND2_X1 U4979 ( .A1(n5450), .A2(n9610), .ZN(n6063) );
  AND2_X1 U4980 ( .A1(n5423), .A2(n5422), .ZN(n8370) );
  NAND2_X1 U4981 ( .A1(n4534), .A2(n5477), .ZN(n5495) );
  NAND2_X1 U4982 ( .A1(n4955), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n4954) );
  NAND2_X1 U4983 ( .A1(n5475), .A2(n5474), .ZN(n4534) );
  AOI21_X1 U4984 ( .B1(n7312), .B2(n5152), .A(n8949), .ZN(n8951) );
  NAND2_X1 U4985 ( .A1(n5396), .A2(n5395), .ZN(n8325) );
  NAND2_X1 U4986 ( .A1(n6817), .A2(n6816), .ZN(n8004) );
  AOI22_X1 U4987 ( .A1(n7683), .A2(n7702), .B1(n7708), .B2(n9679), .ZN(n5275)
         );
  AND2_X1 U4988 ( .A1(n7828), .A2(n8449), .ZN(n9301) );
  NAND2_X1 U4989 ( .A1(n6039), .A2(n7934), .ZN(n7850) );
  NAND2_X1 U4990 ( .A1(n5229), .A2(n5228), .ZN(n7708) );
  AND2_X1 U4991 ( .A1(n6780), .A2(n6779), .ZN(n7574) );
  NOR2_X1 U4992 ( .A1(n6631), .A2(n7594), .ZN(n4945) );
  INV_X1 U4993 ( .A(n6632), .ZN(n8945) );
  OAI21_X1 U4994 ( .B1(n5297), .B2(n5296), .A(n5319), .ZN(n5299) );
  INV_X1 U4995 ( .A(n8936), .ZN(n4758) );
  NAND2_X1 U4996 ( .A1(n5098), .A2(n7447), .ZN(n8416) );
  AND2_X1 U4997 ( .A1(n5969), .A2(n7405), .ZN(n7403) );
  AND4_X1 U4998 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n8230)
         );
  AND2_X1 U4999 ( .A1(n6161), .A2(n6163), .ZN(n6162) );
  INV_X4 U5000 ( .A(n6151), .ZN(n4788) );
  NAND2_X1 U5001 ( .A1(n5441), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5463) );
  AND4_X1 U5002 ( .A1(n6815), .A2(n6814), .A3(n6813), .A4(n6812), .ZN(n7968)
         );
  AND4_X1 U5003 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n8071)
         );
  NAND2_X1 U5004 ( .A1(n4759), .A2(n4650), .ZN(n8936) );
  AND3_X2 U5005 ( .A1(n5272), .A2(n5271), .A3(n5157), .ZN(n10228) );
  AND2_X1 U5006 ( .A1(n6740), .A2(n6739), .ZN(n4650) );
  NAND4_X2 U5007 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n7911)
         );
  INV_X1 U5008 ( .A(n5609), .ZN(n5593) );
  OR3_X1 U5009 ( .A1(n5393), .A2(P1_IR_REG_9__SCAN_IN), .A3(
        P1_IR_REG_8__SCAN_IN), .ZN(n5418) );
  CLKBUF_X1 U5010 ( .A(n6160), .Z(n4294) );
  AND2_X1 U5011 ( .A1(n5270), .A2(n6735), .ZN(n5278) );
  NAND2_X1 U5012 ( .A1(n5805), .A2(n5806), .ZN(n8110) );
  NAND3_X1 U5013 ( .A1(n4629), .A2(n4628), .A3(n4832), .ZN(n7952) );
  OR2_X1 U5014 ( .A1(n8221), .A2(n7219), .ZN(n6740) );
  NOR2_X1 U5015 ( .A1(n7256), .A2(n4959), .ZN(n7255) );
  MUX2_X1 U5016 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5804), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5806) );
  OR2_X1 U5018 ( .A1(n10131), .A2(n10135), .ZN(n5880) );
  BUF_X1 U5019 ( .A(n6773), .Z(n4625) );
  INV_X2 U5020 ( .A(n8218), .ZN(n7044) );
  CLKBUF_X1 U5021 ( .A(n8531), .Z(n4657) );
  AND2_X1 U5022 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  NAND2_X1 U5023 ( .A1(n5322), .A2(SI_5_), .ZN(n5319) );
  INV_X1 U5024 ( .A(n6728), .ZN(n9479) );
  NAND2_X1 U5025 ( .A1(n4424), .A2(n4422), .ZN(n6512) );
  INV_X2 U5026 ( .A(n10122), .ZN(n10134) );
  AND2_X1 U5027 ( .A1(n4892), .A2(n4891), .ZN(n5322) );
  INV_X1 U5028 ( .A(n5473), .ZN(n5474) );
  OAI21_X1 U5029 ( .B1(n5298), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4608), .ZN(
        n5218) );
  XNOR2_X1 U5030 ( .A(n6727), .B(P2_IR_REG_29__SCAN_IN), .ZN(n6728) );
  XNOR2_X1 U5031 ( .A(n6530), .B(n6529), .ZN(n6623) );
  OR2_X1 U5032 ( .A1(n4425), .A2(n6726), .ZN(n4424) );
  NAND2_X1 U5033 ( .A1(n6527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6530) );
  XNOR2_X1 U5034 ( .A(n6570), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7286) );
  OR2_X1 U5035 ( .A1(n7040), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6524) );
  XNOR2_X1 U5036 ( .A(n5269), .B(n5268), .ZN(n7538) );
  AND2_X1 U5037 ( .A1(n5127), .A2(n6724), .ZN(n5126) );
  AND2_X1 U5038 ( .A1(n6529), .A2(n6528), .ZN(n5127) );
  NOR2_X1 U5039 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5167) );
  INV_X1 U5040 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5195) );
  INV_X1 U5041 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n6485) );
  INV_X4 U5042 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X4 U5043 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U5044 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6500) );
  INV_X1 U5045 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4429) );
  INV_X1 U5046 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6529) );
  NOR2_X1 U5047 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5096) );
  NOR2_X1 U5048 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5095) );
  INV_X1 U5049 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5279) );
  INV_X1 U5050 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6538) );
  INV_X1 U5051 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6497) );
  INV_X1 U5052 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6496) );
  INV_X1 U5053 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6495) );
  INV_X1 U5054 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6513) );
  OR2_X2 U5055 ( .A1(n5609), .A2(n7167), .ZN(n5157) );
  BUF_X2 U5056 ( .A(n5260), .Z(n4291) );
  NAND2_X1 U5057 ( .A1(n8633), .A2(n8388), .ZN(n5260) );
  NAND2_X1 U5058 ( .A1(n7397), .A2(n5258), .ZN(n7390) );
  NAND2_X1 U5059 ( .A1(n4596), .A2(n4595), .ZN(n7397) );
  NAND2_X2 U5060 ( .A1(n7581), .A2(n7582), .ZN(n7580) );
  XNOR2_X1 U5061 ( .A(n4616), .B(n4696), .ZN(n9992) );
  OR2_X2 U5062 ( .A1(n5251), .A2(n6465), .ZN(n5237) );
  NAND2_X1 U5063 ( .A1(n8144), .A2(n4401), .ZN(n6635) );
  NAND2_X4 U5064 ( .A1(n5270), .A2(n4893), .ZN(n5609) );
  AOI21_X2 U5066 ( .B1(n9151), .B2(n8501), .A(n7077), .ZN(n9139) );
  AOI21_X2 U5067 ( .B1(n9501), .B2(n9500), .A(n9561), .ZN(n9502) );
  NAND2_X1 U5068 ( .A1(n5181), .A2(n5182), .ZN(n5751) );
  INV_X2 U5069 ( .A(n10253), .ZN(n7757) );
  NAND2_X2 U5070 ( .A1(n5283), .A2(n5284), .ZN(n10253) );
  NAND2_X1 U5071 ( .A1(n8633), .A2(n5182), .ZN(n4292) );
  NAND2_X1 U5072 ( .A1(n5492), .A2(n5491), .ZN(n8371) );
  NAND2_X2 U5073 ( .A1(n7059), .A2(n8418), .ZN(n7491) );
  BUF_X4 U5074 ( .A(n6422), .Z(n4293) );
  NAND2_X1 U5075 ( .A1(n6162), .A2(n7143), .ZN(n6422) );
  OAI211_X2 U5076 ( .C1(n4475), .C2(n6218), .A(n4474), .B(n7732), .ZN(n7862)
         );
  NAND2_X1 U5077 ( .A1(n8633), .A2(n8388), .ZN(n4295) );
  NAND2_X1 U5078 ( .A1(n8633), .A2(n8388), .ZN(n4296) );
  INV_X4 U5079 ( .A(n4291), .ZN(n5306) );
  AOI21_X2 U5080 ( .B1(n8242), .B2(n5472), .A(n4387), .ZN(n9954) );
  OAI21_X2 U5081 ( .B1(n8371), .B2(n4316), .A(n5510), .ZN(n9945) );
  NAND3_X1 U5082 ( .A1(n4327), .A2(n4419), .A3(n7329), .ZN(n4297) );
  OAI21_X2 U5083 ( .B1(n9872), .B2(n5623), .A(n5622), .ZN(n9850) );
  BUF_X8 U5084 ( .A(n8221), .Z(n4298) );
  NAND2_X2 U5085 ( .A1(n6729), .A2(n9479), .ZN(n8221) );
  AOI21_X2 U5086 ( .B1(n7571), .B2(n6784), .A(n6783), .ZN(n7586) );
  MUX2_X1 U5087 ( .A(n9097), .B(n9389), .S(n9296), .Z(n9103) );
  OAI21_X2 U5088 ( .B1(n9801), .B2(n5699), .A(n5698), .ZN(n9785) );
  OAI21_X2 U5089 ( .B1(n9847), .B2(n4985), .A(n4983), .ZN(n9801) );
  OR2_X1 U5090 ( .A1(n9780), .A2(n9795), .ZN(n6115) );
  NAND2_X1 U5091 ( .A1(n4692), .A2(n4691), .ZN(n5434) );
  NOR2_X1 U5092 ( .A1(n5144), .A2(n5415), .ZN(n4691) );
  NOR2_X1 U5093 ( .A1(n4631), .A2(n8565), .ZN(n4630) );
  NAND2_X1 U5094 ( .A1(n5035), .A2(n7170), .ZN(n4891) );
  NAND2_X1 U5095 ( .A1(n4893), .A2(n7187), .ZN(n4892) );
  INV_X1 U5096 ( .A(n8820), .ZN(n6729) );
  NOR2_X1 U5097 ( .A1(n7000), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n4710) );
  NAND2_X1 U5098 ( .A1(n5099), .A2(n8418), .ZN(n4564) );
  NOR2_X1 U5099 ( .A1(n4365), .A2(n4860), .ZN(n4859) );
  INV_X1 U5100 ( .A(n5148), .ZN(n4860) );
  NOR2_X1 U5101 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5093) );
  NAND2_X1 U5102 ( .A1(n5725), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5749) );
  OR2_X1 U5103 ( .A1(n10031), .A2(n9917), .ZN(n5968) );
  NAND2_X1 U5104 ( .A1(n10031), .A2(n9917), .ZN(n6090) );
  AND2_X1 U5105 ( .A1(n5807), .A2(n4294), .ZN(n6444) );
  NAND2_X1 U5106 ( .A1(n5532), .A2(n5531), .ZN(n5535) );
  INV_X1 U5107 ( .A(n5530), .ZN(n5531) );
  AND2_X1 U5108 ( .A1(n5408), .A2(n5391), .ZN(n4693) );
  NAND2_X1 U5109 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5036) );
  INV_X1 U5110 ( .A(n4625), .ZN(n7033) );
  NAND2_X1 U5111 ( .A1(n8986), .A2(n6591), .ZN(n6596) );
  NAND2_X1 U5112 ( .A1(n4918), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4917) );
  NAND2_X1 U5113 ( .A1(n7050), .A2(n4893), .ZN(n6756) );
  XNOR2_X1 U5114 ( .A(n8641), .B(n9397), .ZN(n9113) );
  NAND2_X1 U5115 ( .A1(n5016), .A2(n5015), .ZN(n6418) );
  INV_X1 U5116 ( .A(n9554), .ZN(n4488) );
  AOI21_X1 U5117 ( .B1(n9753), .B2(n5793), .A(n5769), .ZN(n9766) );
  AND2_X1 U5118 ( .A1(n5924), .A2(n5908), .ZN(n6136) );
  NAND2_X1 U5119 ( .A1(n4462), .A2(n4972), .ZN(n7125) );
  AOI21_X1 U5120 ( .B1(n4973), .B2(n4976), .A(n4370), .ZN(n4972) );
  NAND2_X1 U5121 ( .A1(n9785), .A2(n4973), .ZN(n4462) );
  AND2_X1 U5122 ( .A1(n5554), .A2(n5553), .ZN(n9899) );
  AND2_X1 U5123 ( .A1(n7298), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6442) );
  NAND2_X1 U5124 ( .A1(n9780), .A2(n9659), .ZN(n4684) );
  AND2_X1 U5125 ( .A1(n6058), .A2(n6057), .ZN(n4786) );
  AND2_X1 U5126 ( .A1(n9196), .A2(n9195), .ZN(n4682) );
  INV_X1 U5127 ( .A(n8508), .ZN(n4519) );
  NOR2_X1 U5128 ( .A1(n4745), .A2(n4756), .ZN(n4744) );
  NOR2_X1 U5129 ( .A1(n4752), .A2(n7076), .ZN(n4745) );
  NAND2_X1 U5130 ( .A1(n8936), .A2(n7952), .ZN(n8418) );
  NAND2_X1 U5131 ( .A1(n7973), .A2(n6057), .ZN(n5824) );
  INV_X1 U5132 ( .A(n8082), .ZN(n5089) );
  NAND2_X1 U5133 ( .A1(n4561), .A2(n8537), .ZN(n8541) );
  NAND2_X1 U5134 ( .A1(n7780), .A2(n5155), .ZN(n6581) );
  INV_X1 U5135 ( .A(n7774), .ZN(n4883) );
  OAI21_X1 U5136 ( .B1(n4917), .B2(n4452), .A(n4450), .ZN(n6604) );
  INV_X1 U5137 ( .A(n4451), .ZN(n4450) );
  OAI21_X1 U5138 ( .B1(n9011), .B2(n4452), .A(n6599), .ZN(n4451) );
  NAND2_X1 U5139 ( .A1(n9062), .A2(n6641), .ZN(n6642) );
  OR2_X1 U5140 ( .A1(n7106), .A2(n8926), .ZN(n8537) );
  INV_X1 U5141 ( .A(n9207), .ZN(n4842) );
  NAND2_X1 U5142 ( .A1(n7568), .A2(n7061), .ZN(n4556) );
  AND2_X1 U5143 ( .A1(n8427), .A2(n8439), .ZN(n7061) );
  OR2_X1 U5144 ( .A1(n9403), .A2(n9133), .ZN(n7007) );
  OR2_X1 U5145 ( .A1(n9415), .A2(n9159), .ZN(n8505) );
  OR2_X1 U5146 ( .A1(n9421), .A2(n8886), .ZN(n8500) );
  OR2_X1 U5147 ( .A1(n7068), .A2(n8293), .ZN(n8460) );
  INV_X1 U5148 ( .A(n6517), .ZN(n4425) );
  NAND2_X1 U5149 ( .A1(n7864), .A2(n7863), .ZN(n5012) );
  AND2_X1 U5150 ( .A1(n6358), .A2(n9586), .ZN(n6359) );
  INV_X1 U5151 ( .A(n6139), .ZN(n6004) );
  OR2_X1 U5152 ( .A1(n10009), .A2(n10014), .ZN(n4942) );
  OR2_X1 U5153 ( .A1(n7708), .A2(n7577), .ZN(n6033) );
  NOR3_X1 U5154 ( .A1(n9786), .A2(n9780), .A3(n9987), .ZN(n7133) );
  NAND3_X1 U5155 ( .A1(n5784), .A2(n5783), .A3(n5782), .ZN(n5900) );
  NAND2_X1 U5156 ( .A1(n5771), .A2(n5146), .ZN(n5783) );
  OR2_X1 U5157 ( .A1(n5771), .A2(n5772), .ZN(n5784) );
  NAND2_X1 U5158 ( .A1(n5859), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5799) );
  NAND2_X1 U5159 ( .A1(n5538), .A2(n5537), .ZN(n5557) );
  INV_X1 U5160 ( .A(SI_17_), .ZN(n5537) );
  NAND2_X1 U5161 ( .A1(n5535), .A2(n4701), .ZN(n5558) );
  NAND2_X1 U5162 ( .A1(n5412), .A2(n5411), .ZN(n5433) );
  NAND3_X1 U5163 ( .A1(n4906), .A2(n4905), .A3(n5151), .ZN(n5392) );
  NAND2_X1 U5164 ( .A1(n5372), .A2(n4318), .ZN(n4905) );
  INV_X1 U5165 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5196) );
  INV_X1 U5166 ( .A(n9124), .ZN(n8641) );
  AND2_X1 U5167 ( .A1(n8610), .A2(n8609), .ZN(n8611) );
  OR2_X1 U5168 ( .A1(n8870), .A2(n9159), .ZN(n8609) );
  OR2_X1 U5169 ( .A1(n8599), .A2(n9220), .ZN(n8600) );
  XNOR2_X1 U5170 ( .A(n9421), .B(n7357), .ZN(n8868) );
  INV_X1 U5171 ( .A(n4301), .ZN(n6993) );
  NAND2_X1 U5172 ( .A1(n4652), .A2(n8965), .ZN(n4953) );
  INV_X1 U5173 ( .A(n6635), .ZN(n4652) );
  NAND2_X1 U5174 ( .A1(n6635), .A2(n7232), .ZN(n6636) );
  AND2_X1 U5175 ( .A1(n9021), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n4499) );
  NAND3_X1 U5176 ( .A1(n4921), .A2(P2_REG2_REG_17__SCAN_IN), .A3(n6696), .ZN(
        n9069) );
  NAND2_X1 U5177 ( .A1(n6642), .A2(n9080), .ZN(n6691) );
  NAND2_X1 U5178 ( .A1(n7015), .A2(n7024), .ZN(n9110) );
  INV_X1 U5179 ( .A(n9172), .ZN(n9194) );
  NAND2_X1 U5180 ( .A1(n4841), .A2(n4840), .ZN(n9167) );
  XNOR2_X1 U5181 ( .A(n8210), .B(n9276), .ZN(n8033) );
  OR2_X1 U5182 ( .A1(n8063), .A2(n8103), .ZN(n8434) );
  NAND2_X1 U5183 ( .A1(n8004), .A2(n8071), .ZN(n8450) );
  INV_X1 U5184 ( .A(n4627), .ZN(n5098) );
  AND2_X1 U5185 ( .A1(n5118), .A2(n8492), .ZN(n5117) );
  INV_X1 U5186 ( .A(n5123), .ZN(n5122) );
  OR2_X1 U5187 ( .A1(n9443), .A2(n9221), .ZN(n9196) );
  AND2_X1 U5188 ( .A1(n8515), .A2(n7347), .ZN(n9290) );
  NAND2_X1 U5189 ( .A1(n6723), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4626) );
  OR2_X1 U5190 ( .A1(n6572), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6549) );
  NAND2_X1 U5191 ( .A1(n6185), .A2(n7401), .ZN(n6174) );
  NOR2_X1 U5192 ( .A1(n5018), .A2(n4498), .ZN(n4495) );
  INV_X1 U5193 ( .A(n8361), .ZN(n4498) );
  NOR2_X1 U5194 ( .A1(n9532), .A2(n5020), .ZN(n5019) );
  INV_X1 U5195 ( .A(n6173), .ZN(n4601) );
  NAND2_X1 U5196 ( .A1(n6139), .A2(n6151), .ZN(n4783) );
  AND2_X1 U5197 ( .A1(n5963), .A2(n6153), .ZN(n6146) );
  NOR2_X1 U5198 ( .A1(n5962), .A2(n5961), .ZN(n5963) );
  NAND2_X1 U5199 ( .A1(n5960), .A2(n6136), .ZN(n5961) );
  AND2_X1 U5200 ( .A1(n5733), .A2(n5732), .ZN(n9795) );
  OR2_X1 U5201 ( .A1(n5839), .A2(n9667), .ZN(n5698) );
  AND2_X1 U5202 ( .A1(n5714), .A2(n5713), .ZN(n9810) );
  NAND2_X1 U5203 ( .A1(n4492), .A2(n4348), .ZN(n9894) );
  INV_X1 U5204 ( .A(n9904), .ZN(n5835) );
  INV_X1 U5205 ( .A(n7888), .ZN(n5827) );
  INV_X1 U5206 ( .A(n10015), .ZN(n9952) );
  INV_X1 U5207 ( .A(n5850), .ZN(n4584) );
  OR2_X1 U5208 ( .A1(n6151), .A2(n6393), .ZN(n10277) );
  NAND2_X1 U5209 ( .A1(n10117), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5176) );
  NAND2_X1 U5210 ( .A1(n5141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5178) );
  XNOR2_X1 U5211 ( .A(n5024), .B(n4405), .ZN(n9489) );
  NAND2_X1 U5212 ( .A1(n5025), .A2(n5718), .ZN(n5024) );
  NAND2_X1 U5213 ( .A1(n5720), .A2(n5719), .ZN(n5025) );
  AOI21_X1 U5214 ( .B1(n5040), .B2(n5043), .A(n5038), .ZN(n5037) );
  INV_X1 U5215 ( .A(n5040), .ZN(n4704) );
  INV_X1 U5216 ( .A(n5668), .ZN(n5038) );
  NAND2_X1 U5217 ( .A1(n5805), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5802) );
  OAI22_X1 U5218 ( .A1(n5078), .A2(n9173), .B1(n8886), .B2(n5074), .ZN(n5073)
         );
  INV_X1 U5219 ( .A(n5077), .ZN(n5074) );
  NAND2_X1 U5220 ( .A1(n7352), .A2(n9238), .ZN(n8908) );
  NOR2_X1 U5221 ( .A1(n4302), .A2(n8099), .ZN(n4661) );
  NAND2_X1 U5222 ( .A1(n8583), .A2(n4340), .ZN(n4603) );
  NAND2_X1 U5223 ( .A1(n7030), .A2(n7029), .ZN(n9105) );
  INV_X1 U5224 ( .A(n6596), .ZN(n4919) );
  NAND2_X1 U5225 ( .A1(n6596), .A2(n9002), .ZN(n9011) );
  NAND2_X1 U5226 ( .A1(n9395), .A2(n9383), .ZN(n9316) );
  NAND2_X1 U5227 ( .A1(n7012), .A2(n7011), .ZN(n9397) );
  OAI21_X1 U5228 ( .B1(n9644), .B2(n6387), .A(n6386), .ZN(n6392) );
  AND2_X1 U5229 ( .A1(n6408), .A2(n6407), .ZN(n9636) );
  NAND2_X1 U5230 ( .A1(n6399), .A2(n10221), .ZN(n9659) );
  NOR2_X1 U5231 ( .A1(n7809), .A2(n7810), .ZN(n7808) );
  NAND2_X1 U5232 ( .A1(n5939), .A2(n5938), .ZN(n9723) );
  NAND2_X1 U5233 ( .A1(n8425), .A2(n4756), .ZN(n4547) );
  NAND2_X1 U5234 ( .A1(n8424), .A2(n8515), .ZN(n4548) );
  NAND2_X1 U5235 ( .A1(n4678), .A2(n4677), .ZN(n8453) );
  NAND2_X1 U5236 ( .A1(n8447), .A2(n4756), .ZN(n4677) );
  NAND2_X1 U5237 ( .A1(n8435), .A2(n8515), .ZN(n4678) );
  INV_X1 U5238 ( .A(n8436), .ZN(n4544) );
  NOR2_X1 U5239 ( .A1(n8442), .A2(n8515), .ZN(n4543) );
  INV_X1 U5240 ( .A(n8437), .ZN(n4545) );
  NOR2_X1 U5241 ( .A1(n8443), .A2(n4756), .ZN(n4613) );
  INV_X1 U5242 ( .A(n8444), .ZN(n4614) );
  INV_X1 U5243 ( .A(n8442), .ZN(n4612) );
  OR2_X1 U5244 ( .A1(n6027), .A2(n6151), .ZN(n4819) );
  AND2_X1 U5245 ( .A1(n8468), .A2(n8469), .ZN(n4767) );
  INV_X1 U5246 ( .A(n8466), .ZN(n4768) );
  NAND2_X1 U5247 ( .A1(n4792), .A2(n5315), .ZN(n4791) );
  INV_X1 U5248 ( .A(n5824), .ZN(n6047) );
  NAND2_X1 U5249 ( .A1(n4817), .A2(n4816), .ZN(n4815) );
  NOR2_X1 U5250 ( .A1(n6063), .A2(n8115), .ZN(n4816) );
  NAND2_X1 U5251 ( .A1(n4332), .A2(n4813), .ZN(n4812) );
  NOR2_X1 U5252 ( .A1(n6074), .A2(n6075), .ZN(n4813) );
  NAND2_X1 U5253 ( .A1(n4536), .A2(n4756), .ZN(n4750) );
  NAND2_X1 U5254 ( .A1(n8493), .A2(n9196), .ZN(n4536) );
  NAND2_X1 U5255 ( .A1(n4681), .A2(n8515), .ZN(n4680) );
  INV_X1 U5256 ( .A(n8490), .ZN(n4748) );
  NOR2_X1 U5257 ( .A1(n4747), .A2(n8515), .ZN(n4746) );
  INV_X1 U5258 ( .A(n4754), .ZN(n4747) );
  AOI21_X1 U5259 ( .B1(n4750), .B2(n8489), .A(n4755), .ZN(n4754) );
  NAND2_X1 U5260 ( .A1(n8496), .A2(n8492), .ZN(n4755) );
  NOR2_X1 U5261 ( .A1(n8515), .A2(n4750), .ZN(n4749) );
  NOR2_X1 U5262 ( .A1(n9913), .A2(n4788), .ZN(n4777) );
  NOR2_X1 U5263 ( .A1(n4782), .A2(n9913), .ZN(n4776) );
  NOR2_X1 U5264 ( .A1(n4780), .A2(n5837), .ZN(n4779) );
  NAND2_X1 U5265 ( .A1(n4515), .A2(n4358), .ZN(n8513) );
  NOR2_X1 U5266 ( .A1(n5470), .A2(n9961), .ZN(n6066) );
  AND2_X1 U5267 ( .A1(n5106), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U5268 ( .A1(n5101), .A2(n8509), .ZN(n4558) );
  NAND2_X1 U5269 ( .A1(n5004), .A2(n6301), .ZN(n5003) );
  INV_X1 U5270 ( .A(n6293), .ZN(n5004) );
  NAND2_X1 U5271 ( .A1(n4799), .A2(n4788), .ZN(n4798) );
  NAND2_X1 U5272 ( .A1(n9802), .A2(n4328), .ZN(n4794) );
  NAND2_X1 U5273 ( .A1(n4971), .A2(n5556), .ZN(n4970) );
  INV_X1 U5274 ( .A(n5555), .ZN(n4971) );
  OR2_X1 U5275 ( .A1(n7140), .A2(n9766), .ZN(n6129) );
  INV_X1 U5276 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5560) );
  INV_X1 U5277 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5536) );
  INV_X1 U5278 ( .A(n5033), .ZN(n5032) );
  OAI21_X1 U5279 ( .B1(n5494), .B2(n5034), .A(n5512), .ZN(n5033) );
  INV_X1 U5280 ( .A(n5511), .ZN(n5512) );
  INV_X1 U5281 ( .A(n5497), .ZN(n5034) );
  NAND2_X1 U5282 ( .A1(n8294), .A2(n8928), .ZN(n5088) );
  XNOR2_X1 U5283 ( .A(n9350), .B(n7357), .ZN(n8599) );
  NAND2_X1 U5284 ( .A1(n8539), .A2(n8409), .ZN(n8573) );
  INV_X1 U5285 ( .A(n8573), .ZN(n4761) );
  NAND2_X1 U5286 ( .A1(n4551), .A2(n4354), .ZN(n4764) );
  INV_X1 U5287 ( .A(n8528), .ZN(n4617) );
  NOR2_X1 U5288 ( .A1(n7244), .A2(n6627), .ZN(n6628) );
  AND2_X1 U5289 ( .A1(n7253), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6627) );
  OR2_X1 U5290 ( .A1(n7240), .A2(n6565), .ZN(n4439) );
  NOR2_X1 U5291 ( .A1(n8951), .A2(n4346), .ZN(n6576) );
  NAND2_X1 U5292 ( .A1(n4924), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4443) );
  INV_X1 U5293 ( .A(n8137), .ZN(n4871) );
  AND2_X1 U5294 ( .A1(n6718), .A2(n4720), .ZN(n4719) );
  INV_X1 U5295 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n4720) );
  INV_X1 U5296 ( .A(n6907), .ZN(n6719) );
  AND2_X1 U5297 ( .A1(n6716), .A2(n4717), .ZN(n4716) );
  INV_X1 U5298 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n4717) );
  INV_X1 U5299 ( .A(n6869), .ZN(n6717) );
  NAND2_X1 U5300 ( .A1(n6714), .A2(n6713), .ZN(n6835) );
  INV_X1 U5301 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6713) );
  INV_X1 U5302 ( .A(n6827), .ZN(n6714) );
  NAND2_X1 U5303 ( .A1(n6708), .A2(n6707), .ZN(n6789) );
  INV_X1 U5304 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6708) );
  INV_X1 U5305 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6707) );
  INV_X1 U5306 ( .A(n7904), .ZN(n4623) );
  NAND2_X1 U5307 ( .A1(n4624), .A2(n9379), .ZN(n8421) );
  AND2_X1 U5308 ( .A1(n4302), .A2(n7079), .ZN(n7080) );
  AND2_X1 U5309 ( .A1(n8906), .A2(n9409), .ZN(n8504) );
  OR2_X1 U5310 ( .A1(n9409), .A2(n8906), .ZN(n8511) );
  OR2_X1 U5311 ( .A1(n9457), .A2(n9235), .ZN(n8478) );
  INV_X1 U5312 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6595) );
  NAND2_X1 U5313 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6557) );
  OAI21_X1 U5314 ( .B1(n5013), .B2(n5011), .A(n6236), .ZN(n5010) );
  NOR2_X1 U5315 ( .A1(n4483), .A2(n5002), .ZN(n4482) );
  NOR2_X1 U5316 ( .A1(n9606), .A2(n4484), .ZN(n4483) );
  INV_X1 U5317 ( .A(n6279), .ZN(n4484) );
  INV_X1 U5318 ( .A(n6301), .ZN(n5005) );
  OR2_X1 U5319 ( .A1(n5765), .A2(n6432), .ZN(n5787) );
  NAND2_X1 U5320 ( .A1(n5747), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5765) );
  INV_X1 U5321 ( .A(n5749), .ZN(n5747) );
  OAI21_X1 U5322 ( .B1(n6112), .B2(n5131), .A(n6115), .ZN(n4478) );
  OR2_X1 U5323 ( .A1(n9806), .A2(n6112), .ZN(n4479) );
  NOR2_X1 U5324 ( .A1(n9792), .A2(n6021), .ZN(n5131) );
  NAND2_X1 U5325 ( .A1(n9846), .A2(n5660), .ZN(n4987) );
  INV_X1 U5326 ( .A(n5660), .ZN(n4984) );
  NAND2_X1 U5327 ( .A1(n4490), .A2(n4642), .ZN(n9803) );
  AND2_X1 U5328 ( .A1(n5136), .A2(n9819), .ZN(n4642) );
  NAND2_X1 U5329 ( .A1(n9857), .A2(n5133), .ZN(n4490) );
  AND2_X1 U5330 ( .A1(n9904), .A2(n4970), .ZN(n4965) );
  NOR2_X1 U5331 ( .A1(n4968), .A2(n5556), .ZN(n4967) );
  INV_X1 U5332 ( .A(n4970), .ZN(n4968) );
  NOR2_X1 U5333 ( .A1(n10051), .A2(n10055), .ZN(n4929) );
  INV_X1 U5334 ( .A(n4981), .ZN(n4980) );
  OAI21_X1 U5335 ( .B1(n7933), .B2(n4982), .A(n7984), .ZN(n4981) );
  INV_X1 U5336 ( .A(n5364), .ZN(n4982) );
  AND2_X1 U5337 ( .A1(n7702), .A2(n7686), .ZN(n5273) );
  INV_X1 U5338 ( .A(n6388), .ZN(n7612) );
  INV_X1 U5339 ( .A(n5884), .ZN(n6164) );
  OR2_X1 U5340 ( .A1(n10114), .A2(n5879), .ZN(n6389) );
  NOR2_X1 U5341 ( .A1(n4942), .A2(n9825), .ZN(n4941) );
  AND2_X1 U5342 ( .A1(n6069), .A2(n6068), .ZN(n9958) );
  AND2_X1 U5343 ( .A1(n4590), .A2(n8238), .ZN(n6394) );
  NAND2_X1 U5344 ( .A1(n5720), .A2(n5717), .ZN(n5735) );
  AND2_X1 U5345 ( .A1(n5737), .A2(n5718), .ZN(n5734) );
  NOR2_X1 U5346 ( .A1(n5662), .A2(n5045), .ZN(n5044) );
  INV_X1 U5347 ( .A(n5645), .ZN(n5045) );
  OAI21_X1 U5348 ( .B1(n5535), .B2(n5049), .A(n4363), .ZN(n5627) );
  NAND2_X1 U5349 ( .A1(n5048), .A2(n4702), .ZN(n4700) );
  NAND2_X1 U5350 ( .A1(n5051), .A2(n5577), .ZN(n4527) );
  XNOR2_X1 U5351 ( .A(n5476), .B(SI_13_), .ZN(n5473) );
  NAND2_X1 U5352 ( .A1(n4531), .A2(n5454), .ZN(n5475) );
  NAND2_X1 U5353 ( .A1(n5434), .A2(n4532), .ZN(n4531) );
  XNOR2_X1 U5354 ( .A(n5452), .B(SI_12_), .ZN(n5451) );
  NAND2_X1 U5355 ( .A1(n5344), .A2(SI_8_), .ZN(n5368) );
  AND2_X1 U5356 ( .A1(n5326), .A2(n4378), .ZN(n5027) );
  NAND2_X1 U5357 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  INV_X1 U5358 ( .A(n5192), .ZN(n5226) );
  NAND2_X1 U5359 ( .A1(n5080), .A2(n8800), .ZN(n5078) );
  NAND2_X1 U5360 ( .A1(n4421), .A2(n4337), .ZN(n4419) );
  NAND2_X1 U5361 ( .A1(n5085), .A2(n5089), .ZN(n5084) );
  INV_X1 U5362 ( .A(n5086), .ZN(n5085) );
  INV_X1 U5363 ( .A(n8083), .ZN(n5087) );
  AND2_X1 U5364 ( .A1(n5060), .A2(n8823), .ZN(n5059) );
  XNOR2_X1 U5365 ( .A(n4297), .B(n7499), .ZN(n7360) );
  AND2_X1 U5366 ( .A1(n8890), .A2(n5066), .ZN(n5065) );
  OR2_X1 U5367 ( .A1(n8218), .A2(n6761), .ZN(n6762) );
  OAI22_X1 U5368 ( .A1(n8218), .A2(n6738), .B1(n6773), .B2(n7951), .ZN(n4757)
         );
  NAND2_X1 U5369 ( .A1(n4438), .A2(n6563), .ZN(n7218) );
  NAND2_X1 U5370 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(n4959), .ZN(n4958) );
  NOR2_X1 U5371 ( .A1(n7224), .A2(n7502), .ZN(n7223) );
  NOR2_X1 U5372 ( .A1(n7246), .A2(n7245), .ZN(n7244) );
  XNOR2_X1 U5373 ( .A(n7253), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n7242) );
  NOR2_X1 U5374 ( .A1(n7241), .A2(n7242), .ZN(n7240) );
  NAND2_X1 U5375 ( .A1(n6576), .A2(n7633), .ZN(n4924) );
  NAND2_X1 U5376 ( .A1(n4954), .A2(n4505), .ZN(n4658) );
  AOI21_X1 U5377 ( .B1(n4881), .B2(n4305), .A(n4379), .ZN(n4880) );
  NAND2_X1 U5378 ( .A1(n4914), .A2(n8164), .ZN(n4913) );
  NAND2_X1 U5379 ( .A1(n4874), .A2(n4886), .ZN(n4873) );
  INV_X1 U5380 ( .A(n4877), .ZN(n4874) );
  AOI21_X1 U5381 ( .B1(n4880), .B2(n4882), .A(n4878), .ZN(n4877) );
  INV_X1 U5382 ( .A(n8165), .ZN(n4878) );
  INV_X1 U5383 ( .A(n4880), .ZN(n4879) );
  INV_X1 U5384 ( .A(n4886), .ZN(n4875) );
  INV_X1 U5385 ( .A(n6582), .ZN(n8150) );
  INV_X1 U5386 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6584) );
  AND2_X1 U5387 ( .A1(n4317), .A2(n4953), .ZN(n8979) );
  NAND2_X1 U5388 ( .A1(n4442), .A2(n4440), .ZN(n8986) );
  AOI21_X1 U5389 ( .B1(n6587), .B2(n8957), .A(n4441), .ZN(n4440) );
  NAND2_X1 U5390 ( .A1(n8956), .A2(n6587), .ZN(n4442) );
  INV_X1 U5391 ( .A(n8987), .ZN(n4441) );
  INV_X1 U5392 ( .A(n6604), .ZN(n6605) );
  OAI21_X1 U5393 ( .B1(n9016), .B2(n9015), .A(n4410), .ZN(n9035) );
  NAND2_X1 U5394 ( .A1(n9051), .A2(n4664), .ZN(n6608) );
  NAND2_X1 U5395 ( .A1(n9058), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4664) );
  NAND2_X1 U5396 ( .A1(n4868), .A2(n6700), .ZN(n4867) );
  INV_X1 U5397 ( .A(n6701), .ZN(n4868) );
  NAND2_X1 U5398 ( .A1(n6988), .A2(n6987), .ZN(n7000) );
  INV_X1 U5399 ( .A(n6989), .ZN(n6988) );
  OR2_X1 U5400 ( .A1(n6959), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6961) );
  INV_X1 U5401 ( .A(n4280), .ZN(n4843) );
  OR2_X1 U5402 ( .A1(n6898), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6907) );
  INV_X1 U5403 ( .A(n4856), .ZN(n4855) );
  NOR2_X1 U5404 ( .A1(n8556), .A2(n5113), .ZN(n5112) );
  INV_X1 U5405 ( .A(n8450), .ZN(n5113) );
  AND4_X1 U5406 ( .A1(n6805), .A2(n6804), .A3(n6803), .A4(n6802), .ZN(n7588)
         );
  OAI211_X1 U5407 ( .C1(n6756), .C2(n7183), .A(n6755), .B(n6754), .ZN(n7409)
         );
  INV_X1 U5408 ( .A(n7230), .ZN(n6741) );
  NOR2_X1 U5409 ( .A1(n8803), .A2(n8802), .ZN(n8808) );
  NAND2_X1 U5410 ( .A1(n9092), .A2(n9290), .ZN(n9094) );
  AOI21_X1 U5411 ( .B1(n6971), .B2(n4838), .A(n6970), .ZN(n4836) );
  INV_X1 U5412 ( .A(n9290), .ZN(n9234) );
  NAND2_X1 U5413 ( .A1(n8498), .A2(n4579), .ZN(n4578) );
  INV_X1 U5414 ( .A(n8497), .ZN(n4579) );
  AND2_X1 U5415 ( .A1(n8498), .A2(n8494), .ZN(n4580) );
  OR2_X1 U5416 ( .A1(n8606), .A2(n9194), .ZN(n8494) );
  AND2_X1 U5417 ( .A1(n7075), .A2(n5121), .ZN(n5120) );
  AOI21_X1 U5418 ( .B1(n5115), .B2(n4571), .A(n8350), .ZN(n4570) );
  INV_X1 U5419 ( .A(n7069), .ZN(n4571) );
  AOI21_X1 U5420 ( .B1(n4377), .B2(n4850), .A(n4847), .ZN(n4846) );
  NOR2_X1 U5421 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5091) );
  NOR2_X1 U5422 ( .A1(P2_IR_REG_5__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5094) );
  NOR2_X1 U5423 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5092) );
  AND2_X1 U5424 ( .A1(n5095), .A2(n5096), .ZN(n4435) );
  INV_X1 U5425 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6503) );
  NAND2_X1 U5426 ( .A1(n4425), .A2(n6500), .ZN(n6508) );
  INV_X1 U5427 ( .A(n4423), .ZN(n4422) );
  OAI21_X1 U5428 ( .B1(n6500), .B2(n6726), .A(n6509), .ZN(n4423) );
  NAND2_X1 U5429 ( .A1(n6613), .A2(n6612), .ZN(n6619) );
  INV_X1 U5430 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U5431 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4503) );
  NAND2_X1 U5432 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4504) );
  INV_X1 U5433 ( .A(n4640), .ZN(n5691) );
  NAND2_X1 U5434 ( .A1(n4639), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5426) );
  INV_X1 U5435 ( .A(n5399), .ZN(n4639) );
  NAND2_X1 U5436 ( .A1(n8260), .A2(n4351), .ZN(n6254) );
  NAND2_X1 U5437 ( .A1(n4995), .A2(n4994), .ZN(n9553) );
  INV_X1 U5438 ( .A(n4641), .ZN(n5631) );
  NAND2_X1 U5439 ( .A1(n9542), .A2(n6271), .ZN(n9605) );
  OR2_X1 U5440 ( .A1(n5651), .A2(n9624), .ZN(n5674) );
  NAND2_X1 U5441 ( .A1(n4641), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5651) );
  NAND2_X1 U5442 ( .A1(n8260), .A2(n6247), .ZN(n6253) );
  XNOR2_X1 U5443 ( .A(n6184), .B(n6379), .ZN(n6189) );
  XNOR2_X1 U5444 ( .A(n7538), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n7541) );
  NAND2_X1 U5445 ( .A1(n7540), .A2(n7541), .ZN(n7539) );
  NAND2_X1 U5446 ( .A1(n4737), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U5447 ( .A1(n6470), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4736) );
  NAND2_X1 U5448 ( .A1(n4735), .A2(n4734), .ZN(n4733) );
  INV_X1 U5449 ( .A(n9708), .ZN(n4734) );
  NAND2_X1 U5450 ( .A1(n7644), .A2(n7643), .ZN(n4646) );
  AND2_X1 U5451 ( .A1(n7234), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4827) );
  NOR2_X1 U5452 ( .A1(n4831), .A2(n4722), .ZN(n4721) );
  INV_X1 U5453 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n4722) );
  INV_X1 U5454 ( .A(n4828), .ZN(n6474) );
  NAND2_X1 U5455 ( .A1(n10172), .A2(n6457), .ZN(n10190) );
  NAND2_X1 U5456 ( .A1(n5786), .A2(n5785), .ZN(n5817) );
  AND2_X1 U5457 ( .A1(n9806), .A2(n5131), .ZN(n9794) );
  INV_X1 U5458 ( .A(n9792), .ZN(n4594) );
  AOI21_X1 U5459 ( .B1(n9879), .B2(n4779), .A(n5836), .ZN(n9859) );
  INV_X1 U5460 ( .A(n6092), .ZN(n5836) );
  NAND2_X1 U5461 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  AND2_X1 U5462 ( .A1(n5601), .A2(n5600), .ZN(n9898) );
  NAND2_X1 U5463 ( .A1(n9930), .A2(n5128), .ZN(n4492) );
  NAND2_X1 U5464 ( .A1(n9938), .A2(n9926), .ZN(n9919) );
  AND2_X1 U5465 ( .A1(n5573), .A2(n5572), .ZN(n9917) );
  NAND2_X1 U5466 ( .A1(n5529), .A2(n5528), .ZN(n9912) );
  NAND2_X1 U5467 ( .A1(n8373), .A2(n6078), .ZN(n9931) );
  NAND2_X1 U5468 ( .A1(n9931), .A2(n9946), .ZN(n9930) );
  INV_X1 U5469 ( .A(n9669), .ZN(n9918) );
  NAND2_X1 U5470 ( .A1(n9957), .A2(n5833), .ZN(n5143) );
  AND2_X1 U5471 ( .A1(n9958), .A2(n9956), .ZN(n5833) );
  NAND2_X1 U5472 ( .A1(n4489), .A2(n5828), .ZN(n8245) );
  INV_X1 U5473 ( .A(n5443), .ZN(n5441) );
  INV_X1 U5474 ( .A(n9673), .ZN(n8320) );
  AND4_X1 U5475 ( .A1(n5389), .A2(n5388), .A3(n5387), .A4(n5386), .ZN(n7890)
         );
  NAND2_X1 U5476 ( .A1(n5982), .A2(n5825), .ZN(n5826) );
  NAND2_X1 U5477 ( .A1(n6058), .A2(n6061), .ZN(n7888) );
  NAND2_X1 U5478 ( .A1(n4510), .A2(n6033), .ZN(n4508) );
  AND2_X1 U5479 ( .A1(n7683), .A2(n6027), .ZN(n4507) );
  NAND2_X1 U5480 ( .A1(n5278), .A2(n7151), .ZN(n4457) );
  INV_X1 U5481 ( .A(n4459), .ZN(n4458) );
  INV_X1 U5482 ( .A(n5478), .ZN(n5175) );
  INV_X1 U5483 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U5484 ( .A(n5735), .B(n5734), .ZN(n9493) );
  INV_X1 U5485 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5857) );
  INV_X1 U5486 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5798) );
  INV_X1 U5487 ( .A(n5640), .ZN(n5642) );
  AND2_X1 U5488 ( .A1(n5682), .A2(n5667), .ZN(n5668) );
  AOI21_X1 U5489 ( .B1(n5044), .B2(n5042), .A(n5041), .ZN(n5040) );
  INV_X1 U5490 ( .A(n5661), .ZN(n5041) );
  INV_X1 U5491 ( .A(n5641), .ZN(n5042) );
  INV_X1 U5492 ( .A(n5044), .ZN(n5043) );
  OAI21_X1 U5493 ( .B1(n5558), .B2(n5050), .A(n5048), .ZN(n5625) );
  OAI211_X1 U5494 ( .C1(n5558), .C2(n4527), .A(n4523), .B(n4521), .ZN(n7875)
         );
  INV_X1 U5495 ( .A(n4524), .ZN(n4523) );
  NAND2_X1 U5496 ( .A1(n5558), .A2(n4522), .ZN(n4521) );
  OAI21_X1 U5497 ( .B1(n5052), .B2(n4527), .A(n4525), .ZN(n4524) );
  NAND2_X1 U5498 ( .A1(n5543), .A2(n5558), .ZN(n7566) );
  NAND2_X1 U5499 ( .A1(n4692), .A2(n4694), .ZN(n5416) );
  OR2_X1 U5500 ( .A1(n5479), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5349) );
  INV_X1 U5501 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U5502 ( .A1(n5298), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4589) );
  NAND2_X1 U5503 ( .A1(n7795), .A2(n7794), .ZN(n7798) );
  OAI21_X1 U5504 ( .B1(n5078), .B2(n8886), .A(n5071), .ZN(n5070) );
  NAND2_X1 U5505 ( .A1(n8886), .A2(n5077), .ZN(n5071) );
  NOR2_X1 U5506 ( .A1(n8912), .A2(n5079), .ZN(n5076) );
  INV_X1 U5507 ( .A(n9379), .ZN(n7484) );
  AND2_X1 U5508 ( .A1(n6947), .A2(n6946), .ZN(n8829) );
  AND2_X1 U5509 ( .A1(n6983), .A2(n6982), .ZN(n9159) );
  AOI21_X1 U5510 ( .B1(n9212), .B2(n7033), .A(n6936), .ZN(n9221) );
  INV_X1 U5511 ( .A(n9145), .ZN(n8906) );
  INV_X1 U5512 ( .A(n8908), .ZN(n8923) );
  INV_X1 U5513 ( .A(n4530), .ZN(n4529) );
  NAND2_X1 U5514 ( .A1(n7020), .A2(n7019), .ZN(n9124) );
  NAND2_X1 U5515 ( .A1(n6734), .A2(n6733), .ZN(n9173) );
  NAND2_X1 U5516 ( .A1(n6956), .A2(n6955), .ZN(n9172) );
  INV_X1 U5517 ( .A(n9220), .ZN(n9248) );
  OAI211_X1 U5518 ( .C1(n4298), .C2(n9260), .A(n6893), .B(n6892), .ZN(n9247)
         );
  OR2_X1 U5519 ( .A1(n4298), .A2(n6771), .ZN(n6777) );
  OR2_X1 U5520 ( .A1(n7334), .A2(n6519), .ZN(n8935) );
  NAND4_X2 U5521 ( .A1(n6743), .A2(n6745), .A3(n6746), .A4(n6744), .ZN(n4627)
         );
  OR2_X1 U5522 ( .A1(n8218), .A2(n6742), .ZN(n6743) );
  OR2_X1 U5523 ( .A1(n6773), .A2(n7257), .ZN(n6744) );
  INV_X1 U5524 ( .A(n8976), .ZN(n9077) );
  OR2_X1 U5525 ( .A1(P2_U3150), .A2(n6678), .ZN(n8976) );
  NAND2_X1 U5526 ( .A1(n6680), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9081) );
  NAND2_X1 U5527 ( .A1(n6650), .A2(n7178), .ZN(n4889) );
  NAND2_X1 U5528 ( .A1(n4500), .A2(n9021), .ZN(n9004) );
  INV_X1 U5529 ( .A(n4917), .ZN(n4916) );
  NAND2_X1 U5530 ( .A1(n4663), .A2(n6905), .ZN(n4921) );
  INV_X1 U5531 ( .A(n6608), .ZN(n4663) );
  AND2_X1 U5532 ( .A1(n4949), .A2(n6691), .ZN(n9072) );
  NAND2_X1 U5533 ( .A1(n4864), .A2(n4863), .ZN(n4862) );
  INV_X1 U5534 ( .A(n7654), .ZN(n4863) );
  NAND2_X1 U5535 ( .A1(n4867), .A2(n9066), .ZN(n4864) );
  OAI21_X1 U5536 ( .B1(n4867), .B2(n8935), .A(n4866), .ZN(n4865) );
  AND2_X1 U5537 ( .A1(n9081), .A2(n7654), .ZN(n4866) );
  OR2_X1 U5538 ( .A1(n6694), .A2(n6618), .ZN(n6621) );
  AND2_X1 U5539 ( .A1(n7254), .A2(n7043), .ZN(n9043) );
  NAND2_X1 U5540 ( .A1(n9112), .A2(n5101), .ZN(n5105) );
  INV_X1 U5541 ( .A(n9397), .ZN(n9116) );
  NOR2_X1 U5542 ( .A1(n9283), .A2(n5110), .ZN(n5109) );
  INV_X1 U5543 ( .A(n8462), .ZN(n5110) );
  OR2_X1 U5544 ( .A1(n8008), .A2(n7351), .ZN(n9238) );
  AND2_X1 U5545 ( .A1(n7446), .A2(n8273), .ZN(n9300) );
  INV_X1 U5546 ( .A(n9238), .ZN(n9299) );
  AND2_X1 U5547 ( .A1(n9383), .A2(n9376), .ZN(n9332) );
  NAND2_X1 U5548 ( .A1(n9383), .A2(n9378), .ZN(n9310) );
  NAND2_X1 U5549 ( .A1(n8533), .A2(n8532), .ZN(n9385) );
  NOR2_X1 U5550 ( .A1(n8813), .A2(n8805), .ZN(n7121) );
  NAND2_X1 U5551 ( .A1(n9107), .A2(n9106), .ZN(n9108) );
  NAND2_X1 U5552 ( .A1(n9133), .A2(n9292), .ZN(n9106) );
  NAND2_X1 U5553 ( .A1(n6737), .A2(n6736), .ZN(n9421) );
  OR2_X1 U5554 ( .A1(n10301), .A2(n9368), .ZN(n8805) );
  INV_X1 U5555 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U5556 ( .A1(n4635), .A2(n9586), .ZN(n4634) );
  INV_X1 U5557 ( .A(n9588), .ZN(n4635) );
  INV_X1 U5558 ( .A(n9659), .ZN(n9630) );
  INV_X1 U5559 ( .A(n4487), .ZN(n4486) );
  OAI21_X1 U5560 ( .B1(n4994), .B2(n4488), .A(n4324), .ZN(n4487) );
  NAND2_X1 U5561 ( .A1(n9552), .A2(n6370), .ZN(n9645) );
  INV_X1 U5562 ( .A(n9647), .ZN(n4685) );
  INV_X1 U5563 ( .A(n9636), .ZN(n9658) );
  NAND2_X1 U5564 ( .A1(n6159), .A2(n4804), .ZN(n4803) );
  NAND2_X1 U5565 ( .A1(n6149), .A2(n8238), .ZN(n4804) );
  NAND2_X1 U5566 ( .A1(n6153), .A2(n6138), .ZN(n6144) );
  OR2_X1 U5567 ( .A1(n5251), .A2(n5250), .ZN(n4471) );
  OAI21_X1 U5568 ( .B1(n7155), .B2(P1_REG1_REG_1__SCAN_IN), .A(n4467), .ZN(
        n9688) );
  NAND2_X1 U5569 ( .A1(n7155), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n4467) );
  OR2_X1 U5570 ( .A1(n7190), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4822) );
  NAND2_X1 U5571 ( .A1(n7504), .A2(n4466), .ZN(n7809) );
  XNOR2_X1 U5572 ( .A(n6455), .B(n7421), .ZN(n10161) );
  NOR2_X1 U5573 ( .A1(n10160), .A2(n10161), .ZN(n10159) );
  NOR2_X1 U5574 ( .A1(n9722), .A2(n9952), .ZN(n9977) );
  AOI211_X1 U5575 ( .C1(n9732), .C2(n9733), .A(n9952), .B(n9731), .ZN(n9981)
         );
  NAND2_X1 U5576 ( .A1(n9770), .A2(n9769), .ZN(n9985) );
  AND2_X1 U5577 ( .A1(n9768), .A2(n9767), .ZN(n9769) );
  OAI21_X1 U5578 ( .B1(n9785), .B2(n4976), .A(n4974), .ZN(n9759) );
  NAND2_X1 U5579 ( .A1(n4903), .A2(n4901), .ZN(n9990) );
  INV_X1 U5580 ( .A(n4902), .ZN(n4901) );
  NAND2_X1 U5581 ( .A1(n4311), .A2(n9966), .ZN(n4903) );
  OAI22_X1 U5582 ( .A1(n9778), .A2(n9962), .B1(n9960), .B2(n9810), .ZN(n4902)
         );
  NAND2_X1 U5583 ( .A1(n9489), .A2(n5744), .ZN(n5023) );
  OR2_X1 U5584 ( .A1(n4287), .A2(n7614), .ZN(n9929) );
  NAND2_X1 U5585 ( .A1(n6398), .A2(n10113), .ZN(n10221) );
  NOR2_X1 U5586 ( .A1(n9743), .A2(n4372), .ZN(n4463) );
  INV_X1 U5587 ( .A(n9752), .ZN(n4674) );
  AOI21_X1 U5588 ( .B1(n9994), .B2(n10250), .A(n4606), .ZN(n10080) );
  INV_X1 U5589 ( .A(n5839), .ZN(n10087) );
  NAND2_X1 U5590 ( .A1(n5099), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U5591 ( .A1(n4741), .A2(n4739), .ZN(n4738) );
  AND2_X1 U5592 ( .A1(n8414), .A2(n4743), .ZN(n4739) );
  NAND2_X1 U5593 ( .A1(n4546), .A2(n8550), .ZN(n8441) );
  OAI21_X1 U5594 ( .B1(n4550), .B2(n4549), .A(n4373), .ZN(n4546) );
  OAI21_X1 U5595 ( .B1(n4738), .B2(n7491), .A(n8548), .ZN(n4550) );
  NAND2_X1 U5596 ( .A1(n4740), .A2(n8419), .ZN(n4549) );
  NAND2_X1 U5597 ( .A1(n4676), .A2(n9301), .ZN(n8442) );
  INV_X1 U5598 ( .A(n8453), .ZN(n4676) );
  NAND2_X1 U5599 ( .A1(n4611), .A2(n4542), .ZN(n4541) );
  MUX2_X1 U5600 ( .A(n8465), .B(n8464), .S(n8515), .Z(n8466) );
  INV_X1 U5601 ( .A(n7850), .ZN(n4792) );
  NAND2_X1 U5602 ( .A1(n4648), .A2(n4647), .ZN(n6045) );
  NAND2_X1 U5603 ( .A1(n6035), .A2(n6151), .ZN(n4647) );
  NAND2_X1 U5604 ( .A1(n6034), .A2(n4788), .ZN(n4648) );
  INV_X1 U5605 ( .A(n8476), .ZN(n4631) );
  NAND2_X1 U5606 ( .A1(n4793), .A2(n4787), .ZN(n6059) );
  NAND2_X1 U5607 ( .A1(n4789), .A2(n4788), .ZN(n4787) );
  AOI21_X1 U5608 ( .B1(n4750), .B2(n4303), .A(n4313), .ZN(n4752) );
  INV_X1 U5609 ( .A(n8495), .ZN(n4753) );
  NOR2_X1 U5610 ( .A1(n4353), .A2(n6067), .ZN(n4814) );
  NAND2_X1 U5611 ( .A1(n4380), .A2(n4519), .ZN(n4516) );
  NAND2_X1 U5612 ( .A1(n8499), .A2(n9177), .ZN(n4518) );
  AOI22_X1 U5613 ( .A1(n4749), .A2(n4754), .B1(n4756), .B2(n4751), .ZN(n4662)
         );
  AND2_X1 U5614 ( .A1(n4519), .A2(n8499), .ZN(n4517) );
  NAND2_X1 U5615 ( .A1(n4775), .A2(n4342), .ZN(n4772) );
  INV_X1 U5616 ( .A(n4778), .ZN(n4773) );
  INV_X1 U5617 ( .A(n4779), .ZN(n4774) );
  NOR2_X1 U5618 ( .A1(n9283), .A2(n8412), .ZN(n8561) );
  AOI21_X1 U5619 ( .B1(n4708), .B2(n8519), .A(n4707), .ZN(n4706) );
  OR2_X1 U5620 ( .A1(n8523), .A2(n9391), .ZN(n4708) );
  INV_X1 U5621 ( .A(n8522), .ZN(n4707) );
  NAND2_X1 U5622 ( .A1(n8518), .A2(n4709), .ZN(n4632) );
  INV_X1 U5623 ( .A(n9113), .ZN(n4709) );
  INV_X1 U5624 ( .A(n6106), .ZN(n4799) );
  INV_X1 U5625 ( .A(n5101), .ZN(n4560) );
  NAND2_X1 U5626 ( .A1(n8538), .A2(n4756), .ZN(n4618) );
  INV_X1 U5627 ( .A(n9012), .ZN(n4452) );
  AOI22_X1 U5628 ( .A1(n9073), .A2(n9074), .B1(n6905), .B2(n6669), .ZN(n6671)
         );
  NOR2_X1 U5629 ( .A1(n6125), .A2(n5923), .ZN(n6003) );
  NAND2_X1 U5630 ( .A1(n6110), .A2(n6151), .ZN(n4795) );
  NOR4_X1 U5631 ( .A1(n9781), .A2(n4788), .A3(n9792), .A4(n6019), .ZN(n6023)
         );
  NAND2_X1 U5632 ( .A1(n5916), .A2(n5915), .ZN(n6125) );
  INV_X1 U5633 ( .A(n5917), .ZN(n5137) );
  NOR2_X1 U5634 ( .A1(n5137), .A2(n5134), .ZN(n5133) );
  INV_X1 U5635 ( .A(n5918), .ZN(n5134) );
  INV_X1 U5636 ( .A(SI_22_), .ZN(n8710) );
  AOI21_X1 U5637 ( .B1(n5048), .B2(n5050), .A(n5047), .ZN(n5046) );
  INV_X1 U5638 ( .A(n5624), .ZN(n5047) );
  INV_X1 U5639 ( .A(n5541), .ZN(n4703) );
  NOR2_X1 U5640 ( .A1(n5455), .A2(n4533), .ZN(n4532) );
  INV_X1 U5641 ( .A(n5433), .ZN(n4533) );
  NAND2_X1 U5642 ( .A1(n5298), .A2(n5217), .ZN(n4608) );
  NAND2_X1 U5643 ( .A1(n5218), .A2(n8677), .ZN(n5318) );
  INV_X1 U5644 ( .A(n7327), .ZN(n4421) );
  INV_X1 U5645 ( .A(n7357), .ZN(n8621) );
  OR2_X1 U5646 ( .A1(n7270), .A2(n6571), .ZN(n4447) );
  NOR2_X1 U5647 ( .A1(n7286), .A2(n6771), .ZN(n6571) );
  NOR2_X1 U5648 ( .A1(n4912), .A2(n8156), .ZN(n4910) );
  NAND2_X1 U5649 ( .A1(n4325), .A2(n6894), .ZN(n4834) );
  NOR2_X1 U5650 ( .A1(n6835), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n4713) );
  OR2_X1 U5651 ( .A1(n6818), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6827) );
  NAND2_X1 U5652 ( .A1(n6712), .A2(n6711), .ZN(n6818) );
  INV_X1 U5653 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6711) );
  INV_X1 U5654 ( .A(n6810), .ZN(n6712) );
  NAND2_X1 U5655 ( .A1(n6710), .A2(n6709), .ZN(n6800) );
  INV_X1 U5656 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U5657 ( .A1(n7574), .A2(n7911), .ZN(n8439) );
  OR2_X1 U5658 ( .A1(n7089), .A2(n7101), .ZN(n7115) );
  NOR3_X1 U5659 ( .A1(n8489), .A2(n7073), .A3(n5124), .ZN(n5123) );
  INV_X1 U5660 ( .A(n8546), .ZN(n5124) );
  NAND2_X1 U5661 ( .A1(n5123), .A2(n9230), .ZN(n5121) );
  OR2_X1 U5662 ( .A1(n9346), .A2(n9233), .ZN(n9195) );
  NOR2_X1 U5663 ( .A1(n6865), .A2(n4853), .ZN(n4852) );
  INV_X1 U5664 ( .A(n6854), .ZN(n4853) );
  NOR2_X1 U5665 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5097) );
  INV_X1 U5666 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6542) );
  NOR2_X1 U5667 ( .A1(n5674), .A2(n5673), .ZN(n4640) );
  INV_X1 U5668 ( .A(n6333), .ZN(n5020) );
  NOR2_X1 U5669 ( .A1(n5615), .A2(n5614), .ZN(n4641) );
  AND2_X1 U5670 ( .A1(n5817), .A2(n7729), .ZN(n6133) );
  NOR2_X1 U5671 ( .A1(n5959), .A2(n7127), .ZN(n5960) );
  INV_X1 U5672 ( .A(n5958), .ZN(n5959) );
  NOR2_X1 U5673 ( .A1(n5957), .A2(n9792), .ZN(n4695) );
  AND2_X1 U5674 ( .A1(n4974), .A2(n9763), .ZN(n4973) );
  OR2_X1 U5675 ( .A1(n9790), .A2(n9810), .ZN(n6116) );
  AND2_X1 U5676 ( .A1(n5503), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U5677 ( .A1(n10065), .A2(n8320), .ZN(n5984) );
  NOR2_X2 U5678 ( .A1(n5824), .A2(n5823), .ZN(n5980) );
  INV_X1 U5679 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5383) );
  AND3_X1 U5680 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5307) );
  AOI21_X1 U5681 ( .B1(n7128), .B2(n6129), .A(n5841), .ZN(n5842) );
  NOR2_X1 U5682 ( .A1(n4938), .A2(n9987), .ZN(n4937) );
  NAND2_X1 U5683 ( .A1(n5812), .A2(n10079), .ZN(n4938) );
  NAND2_X1 U5684 ( .A1(n7403), .A2(n10228), .ZN(n7691) );
  NAND2_X1 U5685 ( .A1(n5868), .A2(n10115), .ZN(n6388) );
  OR2_X1 U5686 ( .A1(n10114), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U5687 ( .A1(n5762), .A2(n5761), .ZN(n5771) );
  NAND2_X1 U5688 ( .A1(n4690), .A2(n5738), .ZN(n5762) );
  AND2_X1 U5689 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  NAND2_X1 U5690 ( .A1(n5735), .A2(n5734), .ZN(n4690) );
  NAND2_X1 U5691 ( .A1(n5683), .A2(n5682), .ZN(n5701) );
  AND2_X1 U5692 ( .A1(n5717), .A2(n5687), .ZN(n5700) );
  NAND2_X1 U5693 ( .A1(n5051), .A2(n5577), .ZN(n5050) );
  NOR2_X1 U5694 ( .A1(n5578), .A2(n5053), .ZN(n5052) );
  INV_X1 U5695 ( .A(n5557), .ZN(n5053) );
  NAND2_X1 U5696 ( .A1(n5604), .A2(n4526), .ZN(n4525) );
  INV_X1 U5697 ( .A(n5577), .ZN(n4526) );
  AND2_X1 U5698 ( .A1(n5052), .A2(n5604), .ZN(n4522) );
  NAND2_X1 U5699 ( .A1(n5544), .A2(n8679), .ZN(n5794) );
  AND2_X1 U5700 ( .A1(n5498), .A2(n8733), .ZN(n5544) );
  AOI21_X1 U5701 ( .B1(n5032), .B2(n5034), .A(n4366), .ZN(n5030) );
  XNOR2_X1 U5702 ( .A(n5514), .B(SI_15_), .ZN(n5511) );
  INV_X1 U5703 ( .A(n5493), .ZN(n5494) );
  XNOR2_X1 U5704 ( .A(n5496), .B(SI_14_), .ZN(n5493) );
  XNOR2_X1 U5705 ( .A(n5325), .B(SI_6_), .ZN(n5321) );
  INV_X1 U5706 ( .A(n5322), .ZN(n5295) );
  NOR2_X1 U5707 ( .A1(n8800), .A2(n8910), .ZN(n5077) );
  AOI21_X2 U5708 ( .B1(n5065), .B2(n5068), .A(n4307), .ZN(n5063) );
  INV_X1 U5709 ( .A(n5065), .ZN(n5064) );
  XNOR2_X1 U5710 ( .A(n8606), .B(n7357), .ZN(n8607) );
  NAND2_X1 U5711 ( .A1(n4430), .A2(n5081), .ZN(n8295) );
  NAND2_X1 U5712 ( .A1(n5082), .A2(n5088), .ZN(n5081) );
  NAND2_X1 U5713 ( .A1(n5084), .A2(n4359), .ZN(n5082) );
  OAI21_X1 U5714 ( .B1(n8078), .B2(n8077), .A(n8076), .ZN(n8199) );
  NAND2_X1 U5715 ( .A1(n6719), .A2(n6718), .ZN(n6919) );
  INV_X1 U5716 ( .A(n8905), .ZN(n8916) );
  NAND2_X1 U5717 ( .A1(n8576), .A2(n4742), .ZN(n8577) );
  NOR2_X1 U5718 ( .A1(n8571), .A2(n8515), .ZN(n4763) );
  AND2_X1 U5719 ( .A1(n8224), .A2(n7039), .ZN(n8926) );
  OR2_X1 U5720 ( .A1(n4298), .A2(n7453), .ZN(n6746) );
  XNOR2_X1 U5721 ( .A(n6647), .B(n7230), .ZN(n7222) );
  NOR2_X1 U5722 ( .A1(n7222), .A2(n7255), .ZN(n7221) );
  NOR2_X1 U5723 ( .A1(n7223), .A2(n6626), .ZN(n7245) );
  XNOR2_X1 U5724 ( .A(n4439), .B(n6767), .ZN(n7211) );
  NAND2_X1 U5725 ( .A1(n7209), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7275) );
  AOI21_X1 U5726 ( .B1(n7275), .B2(n4320), .A(n7274), .ZN(n7277) );
  NAND2_X1 U5727 ( .A1(n7211), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7272) );
  INV_X1 U5728 ( .A(n4439), .ZN(n6568) );
  OR2_X1 U5729 ( .A1(n4304), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6569) );
  NOR2_X1 U5730 ( .A1(n6630), .A2(n7316), .ZN(n6632) );
  AND2_X1 U5731 ( .A1(n6630), .A2(n7316), .ZN(n6631) );
  AND2_X1 U5732 ( .A1(n4445), .A2(n5152), .ZN(n7313) );
  NAND2_X1 U5733 ( .A1(n4446), .A2(n7316), .ZN(n4445) );
  INV_X1 U5734 ( .A(n4447), .ZN(n4446) );
  NAND2_X1 U5735 ( .A1(n4447), .A2(n4444), .ZN(n5152) );
  AND2_X1 U5736 ( .A1(n4888), .A2(n4887), .ZN(n8939) );
  NAND2_X1 U5737 ( .A1(n6651), .A2(n4444), .ZN(n4887) );
  INV_X1 U5738 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U5739 ( .A1(n4668), .A2(n6634), .ZN(n8159) );
  NAND2_X1 U5740 ( .A1(n6536), .A2(n6535), .ZN(n6583) );
  NAND2_X1 U5741 ( .A1(n4367), .A2(n4884), .ZN(n4869) );
  NAND2_X1 U5742 ( .A1(n4501), .A2(n6866), .ZN(n4500) );
  NAND2_X1 U5743 ( .A1(n9025), .A2(n6639), .ZN(n6640) );
  NAND2_X1 U5744 ( .A1(n4957), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9031) );
  AOI21_X1 U5745 ( .B1(n9035), .B2(n9034), .A(n4861), .ZN(n9055) );
  AND2_X1 U5746 ( .A1(n6887), .A2(n6666), .ZN(n4861) );
  NAND2_X1 U5747 ( .A1(n4448), .A2(n9049), .ZN(n9051) );
  NAND2_X1 U5748 ( .A1(n4926), .A2(n9048), .ZN(n4448) );
  NAND2_X1 U5749 ( .A1(n6606), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4926) );
  NAND2_X1 U5750 ( .A1(n6644), .A2(n6689), .ZN(n6693) );
  AOI21_X1 U5751 ( .B1(n9069), .B2(n6696), .A(n6695), .ZN(n6694) );
  AND2_X1 U5752 ( .A1(n8525), .A2(n4334), .ZN(n4857) );
  AND2_X1 U5753 ( .A1(n5108), .A2(n8520), .ZN(n5101) );
  NAND2_X1 U5754 ( .A1(n5108), .A2(n5100), .ZN(n5106) );
  NAND2_X1 U5755 ( .A1(n9100), .A2(n5107), .ZN(n5100) );
  INV_X1 U5756 ( .A(n5106), .ZN(n5104) );
  NAND2_X1 U5757 ( .A1(n4710), .A2(n7013), .ZN(n7024) );
  OR2_X1 U5758 ( .A1(n7024), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8807) );
  INV_X1 U5759 ( .A(n4710), .ZN(n7014) );
  NAND2_X1 U5760 ( .A1(n4714), .A2(n6976), .ZN(n6989) );
  INV_X1 U5761 ( .A(n4714), .ZN(n6977) );
  NAND2_X1 U5762 ( .A1(n6721), .A2(n6720), .ZN(n6959) );
  INV_X1 U5763 ( .A(n6950), .ZN(n6721) );
  INV_X1 U5764 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n4718) );
  NAND2_X1 U5765 ( .A1(n6719), .A2(n4719), .ZN(n6932) );
  AND3_X1 U5766 ( .A1(n6902), .A2(n6901), .A3(n6900), .ZN(n9235) );
  INV_X1 U5767 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n4715) );
  NAND2_X1 U5768 ( .A1(n6717), .A2(n4716), .ZN(n6890) );
  NAND2_X1 U5769 ( .A1(n6717), .A2(n6716), .ZN(n6882) );
  NAND2_X1 U5770 ( .A1(n4711), .A2(n6715), .ZN(n6869) );
  INV_X1 U5771 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6715) );
  INV_X1 U5772 ( .A(n6857), .ZN(n4711) );
  NAND2_X1 U5773 ( .A1(n4713), .A2(n4712), .ZN(n6857) );
  INV_X1 U5774 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4712) );
  INV_X1 U5775 ( .A(n4713), .ZN(n6848) );
  OR2_X1 U5776 ( .A1(n6842), .A2(n8044), .ZN(n6843) );
  INV_X1 U5777 ( .A(n8928), .ZN(n8293) );
  NAND2_X1 U5778 ( .A1(n7063), .A2(n8553), .ZN(n4554) );
  NAND2_X1 U5779 ( .A1(n4556), .A2(n7064), .ZN(n7591) );
  NAND2_X1 U5780 ( .A1(n7591), .A2(n8553), .ZN(n7920) );
  NAND2_X1 U5781 ( .A1(n4564), .A2(n7059), .ZN(n7408) );
  NAND2_X1 U5782 ( .A1(n4563), .A2(n7059), .ZN(n7498) );
  INV_X1 U5783 ( .A(n4564), .ZN(n4563) );
  OR2_X1 U5784 ( .A1(n7090), .A2(n9472), .ZN(n7444) );
  NAND2_X1 U5785 ( .A1(n9105), .A2(n9290), .ZN(n9107) );
  AND2_X1 U5786 ( .A1(n9415), .A2(n9134), .ZN(n6984) );
  AND2_X1 U5787 ( .A1(n8510), .A2(n8511), .ZN(n9140) );
  OAI21_X1 U5788 ( .B1(n4581), .B2(n4577), .A(n4575), .ZN(n9151) );
  INV_X1 U5789 ( .A(n4576), .ZN(n4575) );
  OAI21_X1 U5790 ( .B1(n4580), .B2(n4577), .A(n8500), .ZN(n4576) );
  INV_X1 U5791 ( .A(n4578), .ZN(n4577) );
  AND2_X1 U5792 ( .A1(n9195), .A2(n8546), .ZN(n9217) );
  NAND2_X1 U5793 ( .A1(n9228), .A2(n8481), .ZN(n5125) );
  NAND2_X1 U5794 ( .A1(n4565), .A2(n4566), .ZN(n9244) );
  AOI21_X1 U5795 ( .B1(n4308), .B2(n4572), .A(n4567), .ZN(n4566) );
  INV_X1 U5796 ( .A(n8475), .ZN(n4567) );
  INV_X1 U5797 ( .A(n4852), .ZN(n4851) );
  OR2_X1 U5798 ( .A1(n7329), .A2(n4756), .ZN(n7344) );
  OR2_X1 U5799 ( .A1(n7112), .A2(n7327), .ZN(n7338) );
  NOR2_X1 U5800 ( .A1(n7341), .A2(n9471), .ZN(n7345) );
  AND2_X1 U5801 ( .A1(n7334), .A2(n7149), .ZN(n7350) );
  INV_X1 U5802 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6610) );
  NOR2_X1 U5803 ( .A1(n6540), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n5090) );
  INV_X1 U5804 ( .A(n6553), .ZN(n6561) );
  NAND2_X1 U5805 ( .A1(n6560), .A2(n6559), .ZN(n6562) );
  INV_X1 U5806 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n6558) );
  NOR2_X1 U5807 ( .A1(n6376), .A2(n6375), .ZN(n6387) );
  OR2_X1 U5808 ( .A1(n5384), .A2(n5383), .ZN(n5399) );
  NAND2_X1 U5809 ( .A1(n5355), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5384) );
  INV_X1 U5810 ( .A(n5357), .ZN(n5355) );
  NAND2_X1 U5811 ( .A1(n7862), .A2(n5013), .ZN(n5008) );
  NAND2_X1 U5812 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  NAND2_X1 U5813 ( .A1(n6185), .A2(n5257), .ZN(n6168) );
  OR2_X1 U5814 ( .A1(n6260), .A2(n6259), .ZN(n9539) );
  NAND2_X1 U5815 ( .A1(n4640), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U5816 ( .A1(n9604), .A2(n6279), .ZN(n9499) );
  AND2_X1 U5817 ( .A1(n9588), .A2(n4997), .ZN(n4996) );
  NAND2_X1 U5818 ( .A1(n6359), .A2(n4349), .ZN(n4997) );
  INV_X1 U5819 ( .A(n6359), .ZN(n4998) );
  AOI21_X1 U5820 ( .B1(n5009), .B2(n5011), .A(n4375), .ZN(n5006) );
  NAND2_X1 U5821 ( .A1(n4654), .A2(n4653), .ZN(n9620) );
  INV_X1 U5822 ( .A(n9510), .ZN(n4653) );
  NAND2_X1 U5823 ( .A1(n5565), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5615) );
  NAND2_X1 U5824 ( .A1(n4485), .A2(n4999), .ZN(n9519) );
  AOI21_X1 U5825 ( .B1(n5001), .B2(n5005), .A(n4360), .ZN(n4999) );
  OAI21_X1 U5826 ( .B1(n9605), .B2(n4484), .A(n4482), .ZN(n4485) );
  INV_X1 U5827 ( .A(n6370), .ZN(n5014) );
  AOI21_X1 U5828 ( .B1(n4996), .B2(n4998), .A(n6363), .ZN(n4994) );
  NAND2_X1 U5829 ( .A1(n5483), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5505) );
  INV_X1 U5830 ( .A(n8110), .ZN(n6393) );
  AND2_X1 U5831 ( .A1(n5680), .A2(n5679), .ZN(n9625) );
  AND2_X1 U5832 ( .A1(n5621), .A2(n5620), .ZN(n9527) );
  NAND2_X1 U5833 ( .A1(n5653), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n4960) );
  OR2_X1 U5834 ( .A1(n5251), .A2(n5179), .ZN(n5185) );
  OR2_X1 U5835 ( .A1(n4296), .A2(n5249), .ZN(n4470) );
  OR2_X1 U5836 ( .A1(n5330), .A2(n6176), .ZN(n4469) );
  NOR2_X1 U5837 ( .A1(n7662), .A2(n4823), .ZN(n7509) );
  NOR2_X1 U5838 ( .A1(n4825), .A2(n4824), .ZN(n4823) );
  INV_X1 U5839 ( .A(n7665), .ZN(n4825) );
  AND2_X1 U5840 ( .A1(n7268), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n4723) );
  NOR2_X1 U5841 ( .A1(n4831), .A2(n4830), .ZN(n4829) );
  AND2_X1 U5842 ( .A1(n7518), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4821) );
  NAND2_X1 U5843 ( .A1(n10190), .A2(n10191), .ZN(n6460) );
  OR2_X1 U5844 ( .A1(n10208), .A2(n10207), .ZN(n10210) );
  XNOR2_X1 U5845 ( .A(n6480), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n6488) );
  AND2_X1 U5846 ( .A1(n5787), .A2(n5766), .ZN(n9753) );
  NAND2_X1 U5847 ( .A1(n4479), .A2(n4477), .ZN(n4481) );
  INV_X1 U5848 ( .A(n4478), .ZN(n4477) );
  INV_X1 U5849 ( .A(n4975), .ZN(n4974) );
  OAI22_X1 U5850 ( .A1(n4696), .A2(n4306), .B1(n9795), .B2(n10079), .ZN(n4975)
         );
  OR2_X1 U5851 ( .A1(n9761), .A2(n4290), .ZN(n5757) );
  NOR2_X1 U5852 ( .A1(n9794), .A2(n9776), .ZN(n9777) );
  AND2_X1 U5853 ( .A1(n5728), .A2(n5749), .ZN(n9774) );
  INV_X1 U5854 ( .A(n4986), .ZN(n4985) );
  NAND2_X1 U5855 ( .A1(n9834), .A2(n9846), .ZN(n5135) );
  AND2_X1 U5856 ( .A1(n5910), .A2(n6111), .ZN(n9819) );
  NAND2_X1 U5857 ( .A1(n4939), .A2(n4940), .ZN(n9838) );
  INV_X1 U5858 ( .A(n4942), .ZN(n4939) );
  AND2_X1 U5859 ( .A1(n9879), .A2(n6098), .ZN(n4904) );
  AND2_X1 U5860 ( .A1(n5637), .A2(n5636), .ZN(n9869) );
  INV_X1 U5861 ( .A(n4940), .ZN(n5159) );
  AND2_X1 U5862 ( .A1(n6093), .A2(n6098), .ZN(n9881) );
  NAND2_X1 U5863 ( .A1(n4461), .A2(n4966), .ZN(n9878) );
  AOI21_X1 U5864 ( .B1(n9904), .B2(n4967), .A(n4344), .ZN(n4966) );
  NAND2_X1 U5865 ( .A1(n9912), .A2(n4965), .ZN(n4461) );
  INV_X1 U5866 ( .A(n5565), .ZN(n5567) );
  NOR2_X1 U5867 ( .A1(n4928), .A2(n9939), .ZN(n4927) );
  INV_X1 U5868 ( .A(n4929), .ZN(n4928) );
  NAND2_X1 U5869 ( .A1(n9949), .A2(n5832), .ZN(n9950) );
  NAND2_X1 U5870 ( .A1(n4638), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5443) );
  INV_X1 U5871 ( .A(n5426), .ZN(n4638) );
  INV_X1 U5872 ( .A(n5984), .ZN(n8115) );
  INV_X1 U5873 ( .A(n6060), .ZN(n8116) );
  AOI21_X1 U5874 ( .B1(n7991), .B2(n4964), .A(n4364), .ZN(n4963) );
  INV_X1 U5875 ( .A(n5405), .ZN(n4964) );
  AOI21_X1 U5876 ( .B1(n4980), .B2(n4982), .A(n4362), .ZN(n4978) );
  AND4_X1 U5877 ( .A1(n5404), .A2(n5403), .A3(n5402), .A4(n5401), .ZN(n7993)
         );
  NOR2_X1 U5878 ( .A1(n10260), .A2(n4932), .ZN(n4931) );
  NAND2_X1 U5879 ( .A1(n10275), .A2(n4933), .ZN(n4932) );
  NOR2_X1 U5880 ( .A1(n7768), .A2(n4935), .ZN(n7941) );
  OR2_X1 U5881 ( .A1(n10260), .A2(n7868), .ZN(n4935) );
  NAND2_X1 U5882 ( .A1(n5307), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5333) );
  AND2_X2 U5883 ( .A1(n6036), .A2(n6037), .ZN(n7610) );
  NAND2_X1 U5884 ( .A1(n5810), .A2(n10239), .ZN(n7709) );
  INV_X1 U5885 ( .A(n7691), .ZN(n5810) );
  AOI22_X1 U5886 ( .A1(n5593), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n6443), .B2(
        n6470), .ZN(n5228) );
  NAND2_X1 U5887 ( .A1(n7683), .A2(n7684), .ZN(n7699) );
  OR2_X1 U5888 ( .A1(n5257), .A2(n5969), .ZN(n5819) );
  INV_X1 U5889 ( .A(n9962), .ZN(n9934) );
  INV_X1 U5890 ( .A(n10125), .ZN(n7524) );
  NAND2_X1 U5891 ( .A1(n6389), .A2(n5885), .ZN(n7136) );
  AND2_X1 U5892 ( .A1(n5817), .A2(n10261), .ZN(n4944) );
  AND3_X1 U5893 ( .A1(n6136), .A2(n10250), .A3(n5815), .ZN(n5816) );
  NAND2_X1 U5894 ( .A1(n5595), .A2(n5594), .ZN(n10027) );
  NAND2_X1 U5895 ( .A1(n4286), .A2(n5555), .ZN(n4969) );
  CLKBUF_X1 U5896 ( .A(n9954), .Z(n9955) );
  INV_X1 U5897 ( .A(n7136), .ZN(n7613) );
  NAND2_X1 U5898 ( .A1(n5886), .A2(n10116), .ZN(n7611) );
  OR2_X1 U5899 ( .A1(n10114), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5886) );
  AND2_X1 U5900 ( .A1(n6388), .A2(n6397), .ZN(n7137) );
  NAND2_X1 U5901 ( .A1(n5771), .A2(n5773), .ZN(n5894) );
  XNOR2_X1 U5902 ( .A(n5743), .B(n5758), .ZN(n8383) );
  NAND2_X1 U5903 ( .A1(n5762), .A2(n5760), .ZN(n5743) );
  OR2_X1 U5904 ( .A1(n5799), .A2(n5857), .ZN(n5800) );
  NAND2_X1 U5905 ( .A1(n5039), .A2(n5645), .ZN(n5663) );
  INV_X1 U5906 ( .A(n5794), .ZN(n5797) );
  NOR2_X1 U5907 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5796) );
  NAND2_X1 U5908 ( .A1(n5558), .A2(n5557), .ZN(n4907) );
  NAND2_X1 U5909 ( .A1(n5794), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5561) );
  NAND2_X1 U5910 ( .A1(n5434), .A2(n5433), .ZN(n5456) );
  NAND2_X1 U5911 ( .A1(n5392), .A2(n5391), .ZN(n5407) );
  XNOR2_X1 U5912 ( .A(n5348), .B(n5347), .ZN(n7163) );
  INV_X1 U5913 ( .A(n5227), .ZN(n5301) );
  INV_X1 U5914 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U5915 ( .A1(n5206), .A2(n5205), .ZN(n5265) );
  NAND2_X1 U5916 ( .A1(n7604), .A2(n7690), .ZN(n7698) );
  INV_X1 U5917 ( .A(n9133), .ZN(n8628) );
  OAI21_X1 U5918 ( .B1(n8859), .B2(n5064), .A(n5063), .ZN(n8825) );
  AND2_X1 U5919 ( .A1(n6967), .A2(n6966), .ZN(n9158) );
  NAND2_X1 U5920 ( .A1(n4426), .A2(n4355), .ZN(n8834) );
  NAND2_X1 U5921 ( .A1(n8078), .A2(n4309), .ZN(n5083) );
  NAND2_X1 U5922 ( .A1(n8612), .A2(n8611), .ZN(n4433) );
  OAI21_X1 U5923 ( .B1(n8615), .B2(n8614), .A(n8613), .ZN(n8616) );
  AOI21_X1 U5924 ( .B1(n8859), .B2(n8858), .A(n8857), .ZN(n8892) );
  NAND2_X1 U5925 ( .A1(n5061), .A2(n5059), .ZN(n4427) );
  NAND2_X1 U5926 ( .A1(n4432), .A2(n7361), .ZN(n7367) );
  NAND2_X1 U5927 ( .A1(n8859), .A2(n5067), .ZN(n5062) );
  INV_X1 U5928 ( .A(n7555), .ZN(n4434) );
  OR2_X1 U5929 ( .A1(n7348), .A2(n7347), .ZN(n8905) );
  AND2_X1 U5930 ( .A1(n8224), .A2(n8223), .ZN(n8803) );
  NAND2_X1 U5931 ( .A1(n6996), .A2(n6995), .ZN(n9145) );
  INV_X1 U5932 ( .A(n9159), .ZN(n9134) );
  INV_X1 U5933 ( .A(n9158), .ZN(n9185) );
  INV_X1 U5934 ( .A(n8829), .ZN(n9209) );
  INV_X1 U5935 ( .A(n9235), .ZN(n9258) );
  INV_X1 U5936 ( .A(n8071), .ZN(n9291) );
  OR2_X1 U5937 ( .A1(n4298), .A2(n7914), .ZN(n6766) );
  NOR2_X1 U5938 ( .A1(n7239), .A2(n7238), .ZN(n7237) );
  NAND2_X1 U5939 ( .A1(n7207), .A2(n7206), .ZN(n7205) );
  INV_X1 U5940 ( .A(n4890), .ZN(n7281) );
  NAND2_X1 U5941 ( .A1(n4923), .A2(n4924), .ZN(n7629) );
  NAND2_X1 U5942 ( .A1(n4955), .A2(n4505), .ZN(n7626) );
  AOI21_X1 U5943 ( .B1(n4282), .B2(n7634), .A(n4305), .ZN(n7773) );
  XNOR2_X1 U5944 ( .A(n6578), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7783) );
  NAND2_X1 U5945 ( .A1(n4876), .A2(n4880), .ZN(n8166) );
  NAND2_X1 U5946 ( .A1(n4282), .A2(n4881), .ZN(n4876) );
  NAND2_X1 U5947 ( .A1(n4913), .A2(n6582), .ZN(n8155) );
  NAND2_X1 U5948 ( .A1(n4872), .A2(n4873), .ZN(n8136) );
  NAND2_X1 U5949 ( .A1(n6582), .A2(n4915), .ZN(n4911) );
  NAND2_X1 U5950 ( .A1(n4453), .A2(n8965), .ZN(n6586) );
  INV_X1 U5951 ( .A(n4454), .ZN(n4453) );
  AND2_X1 U5952 ( .A1(n4951), .A2(n4950), .ZN(n8981) );
  NAND2_X1 U5953 ( .A1(n4917), .A2(n9011), .ZN(n4449) );
  AND2_X1 U5954 ( .A1(n6606), .A2(n9048), .ZN(n9042) );
  NAND2_X1 U5955 ( .A1(n4925), .A2(n9048), .ZN(n9041) );
  INV_X1 U5956 ( .A(n4926), .ZN(n4925) );
  NAND2_X1 U5957 ( .A1(n4841), .A2(n4844), .ZN(n9192) );
  NAND2_X1 U5958 ( .A1(n7566), .A2(n7010), .ZN(n4600) );
  NAND2_X1 U5959 ( .A1(n6845), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U5960 ( .A1(n6847), .A2(n6846), .ZN(n8210) );
  NAND2_X1 U5961 ( .A1(n5114), .A2(n8450), .ZN(n8009) );
  OR2_X1 U5962 ( .A1(n7050), .A2(n4920), .ZN(n6768) );
  OR2_X1 U5963 ( .A1(n7050), .A2(n6741), .ZN(n4832) );
  NOR2_X1 U5964 ( .A1(n8813), .A2(n9310), .ZN(n7107) );
  INV_X2 U5965 ( .A(n9307), .ZN(n9383) );
  NAND2_X1 U5966 ( .A1(n9094), .A2(n9093), .ZN(n9095) );
  NAND2_X1 U5967 ( .A1(n9124), .A2(n9292), .ZN(n9093) );
  NAND2_X1 U5968 ( .A1(n6999), .A2(n6998), .ZN(n9403) );
  NAND2_X1 U5969 ( .A1(n6986), .A2(n6985), .ZN(n9409) );
  NAND2_X1 U5970 ( .A1(n4574), .A2(n4578), .ZN(n9156) );
  NAND2_X1 U5971 ( .A1(n4573), .A2(n4580), .ZN(n4574) );
  NAND2_X1 U5972 ( .A1(n4573), .A2(n8494), .ZN(n9178) );
  NAND2_X1 U5973 ( .A1(n5119), .A2(n5117), .ZN(n9182) );
  NAND2_X1 U5974 ( .A1(n7875), .A2(n7010), .ZN(n6931) );
  OAI21_X1 U5975 ( .B1(n4281), .B2(n4325), .A(n6894), .ZN(n9246) );
  NAND2_X1 U5976 ( .A1(n4568), .A2(n4570), .ZN(n9254) );
  NAND2_X1 U5977 ( .A1(n4569), .A2(n5115), .ZN(n4568) );
  INV_X1 U5978 ( .A(n8275), .ZN(n4569) );
  NAND2_X1 U5979 ( .A1(n8275), .A2(n7069), .ZN(n5116) );
  NAND2_X1 U5980 ( .A1(n6868), .A2(n6867), .ZN(n8410) );
  INV_X1 U5981 ( .A(n9467), .ZN(n9428) );
  INV_X1 U5982 ( .A(n7447), .ZN(n7471) );
  NAND2_X1 U5983 ( .A1(n7089), .A2(n7350), .ZN(n7165) );
  NAND2_X1 U5984 ( .A1(n9473), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6725) );
  INV_X1 U5985 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9486) );
  NAND2_X1 U5986 ( .A1(n6512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6514) );
  INV_X1 U5987 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8382) );
  OR2_X1 U5988 ( .A1(n6510), .A2(n6509), .ZN(n6511) );
  NAND2_X1 U5989 ( .A1(n6508), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6510) );
  INV_X1 U5990 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n8722) );
  INV_X1 U5991 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8289) );
  INV_X1 U5992 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n8214) );
  INV_X1 U5993 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8098) );
  INV_X1 U5994 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n8785) );
  NAND2_X1 U5995 ( .A1(n6619), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5054) );
  INV_X1 U5996 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7597) );
  INV_X1 U5997 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7266) );
  INV_X1 U5998 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7233) );
  INV_X1 U5999 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7201) );
  INV_X1 U6000 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7194) );
  NAND2_X1 U6001 ( .A1(n6552), .A2(n6574), .ZN(n7175) );
  INV_X1 U6002 ( .A(n6767), .ZN(n4920) );
  NAND2_X2 U6003 ( .A1(n6556), .A2(n4304), .ZN(n7253) );
  INV_X1 U6004 ( .A(n7653), .ZN(n9494) );
  NAND2_X1 U6005 ( .A1(n6561), .A2(n6562), .ZN(n7230) );
  AND2_X1 U6006 ( .A1(n5659), .A2(n5658), .ZN(n9824) );
  INV_X1 U6007 ( .A(n5018), .ZN(n5017) );
  NAND2_X1 U6008 ( .A1(n6254), .A2(n8360), .ZN(n8317) );
  NOR2_X1 U6009 ( .A1(n6418), .A2(n4329), .ZN(n6439) );
  NAND2_X1 U6010 ( .A1(n4582), .A2(n6179), .ZN(n7474) );
  NAND2_X1 U6011 ( .A1(n5021), .A2(n6333), .ZN(n9533) );
  NAND2_X1 U6012 ( .A1(n5629), .A2(n5628), .ZN(n10014) );
  AND4_X1 U6013 ( .A1(n5468), .A2(n5467), .A3(n5466), .A4(n5465), .ZN(n9961)
         );
  NAND2_X1 U6014 ( .A1(n5000), .A2(n6301), .ZN(n9580) );
  NAND2_X1 U6015 ( .A1(n9499), .A2(n6293), .ZN(n5000) );
  INV_X1 U6016 ( .A(n9643), .ZN(n9652) );
  OR2_X1 U6017 ( .A1(n6412), .A2(n6411), .ZN(n9654) );
  AND4_X1 U6018 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n9610)
         );
  INV_X1 U6019 ( .A(n9654), .ZN(n9640) );
  NAND2_X1 U6020 ( .A1(n7580), .A2(n6213), .ZN(n4476) );
  AOI21_X1 U6021 ( .B1(n6146), .B2(n6147), .A(n4705), .ZN(n6149) );
  NAND2_X1 U6022 ( .A1(n6148), .A2(n6442), .ZN(n4705) );
  INV_X1 U6023 ( .A(n9823), .ZN(n9667) );
  INV_X1 U6024 ( .A(n9625), .ZN(n9835) );
  INV_X1 U6025 ( .A(n9824), .ZN(n9860) );
  INV_X1 U6026 ( .A(n9869), .ZN(n9836) );
  INV_X1 U6027 ( .A(n9527), .ZN(n9882) );
  INV_X1 U6028 ( .A(n9899), .ZN(n9935) );
  INV_X1 U6029 ( .A(n9963), .ZN(n9933) );
  INV_X1 U6030 ( .A(P1_U3973), .ZN(n9670) );
  INV_X1 U6031 ( .A(n9610), .ZN(n5449) );
  OR2_X1 U6032 ( .A1(n5251), .A2(n6467), .ZN(n5263) );
  BUF_X1 U6033 ( .A(n5257), .Z(n4643) );
  NAND2_X1 U6034 ( .A1(n9688), .A2(n9687), .ZN(n9686) );
  NAND2_X1 U6035 ( .A1(n7539), .A2(n6468), .ZN(n9699) );
  NAND2_X1 U6036 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  NAND2_X1 U6037 ( .A1(n9702), .A2(n9703), .ZN(n9701) );
  AND2_X1 U6038 ( .A1(n6484), .A2(n6483), .ZN(n10141) );
  INV_X1 U6039 ( .A(n4735), .ZN(n9709) );
  INV_X1 U6040 ( .A(n4733), .ZN(n9707) );
  XNOR2_X1 U6041 ( .A(n5282), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9714) );
  AND2_X1 U6042 ( .A1(n4733), .A2(n4732), .ZN(n7642) );
  NAND2_X1 U6043 ( .A1(n9714), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n4732) );
  INV_X1 U6044 ( .A(n4646), .ZN(n7646) );
  NAND2_X1 U6045 ( .A1(n7647), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4645) );
  AND2_X1 U6046 ( .A1(n7676), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n4727) );
  NOR2_X1 U6047 ( .A1(n7659), .A2(n4726), .ZN(n7506) );
  AND2_X1 U6048 ( .A1(n7665), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n4726) );
  NAND2_X1 U6049 ( .A1(n7506), .A2(n7505), .ZN(n7504) );
  AND2_X1 U6050 ( .A1(n7202), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4644) );
  AND2_X1 U6051 ( .A1(n7202), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4725) );
  NOR2_X1 U6052 ( .A1(n8020), .A2(n4724), .ZN(n8181) );
  AND2_X1 U6053 ( .A1(n7234), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4724) );
  NAND2_X1 U6054 ( .A1(n8181), .A2(n8182), .ZN(n8180) );
  NAND2_X1 U6055 ( .A1(n8184), .A2(n4826), .ZN(n8342) );
  OR2_X1 U6056 ( .A1(n7263), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4826) );
  NOR2_X1 U6057 ( .A1(n8339), .A2(n8340), .ZN(n8338) );
  NAND2_X1 U6058 ( .A1(n8180), .A2(n4465), .ZN(n8339) );
  OR2_X1 U6059 ( .A1(n7263), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n4465) );
  XNOR2_X1 U6060 ( .A(n4828), .B(n10167), .ZN(n10164) );
  NOR2_X1 U6061 ( .A1(n10164), .A2(n10163), .ZN(n10162) );
  INV_X1 U6062 ( .A(n10211), .ZN(n10158) );
  NOR2_X1 U6063 ( .A1(n10159), .A2(n6456), .ZN(n10174) );
  NAND2_X1 U6064 ( .A1(n10174), .A2(n10173), .ZN(n10172) );
  NOR2_X1 U6065 ( .A1(n10143), .A2(n5846), .ZN(n10211) );
  NAND2_X1 U6066 ( .A1(n6488), .A2(n9716), .ZN(n4602) );
  OAI21_X1 U6067 ( .B1(n10220), .B2(n6485), .A(n9525), .ZN(n6486) );
  NAND2_X2 U6068 ( .A1(n5906), .A2(n5905), .ZN(n9733) );
  AOI21_X1 U6069 ( .B1(n9806), .B2(n6020), .A(n4594), .ZN(n9793) );
  NAND2_X1 U6070 ( .A1(n5611), .A2(n5610), .ZN(n10020) );
  INV_X1 U6071 ( .A(n10027), .ZN(n9890) );
  NAND2_X1 U6072 ( .A1(n4492), .A2(n5967), .ZN(n9896) );
  NAND2_X1 U6073 ( .A1(n9930), .A2(n6081), .ZN(n9914) );
  NAND2_X1 U6074 ( .A1(n5138), .A2(n5826), .ZN(n7887) );
  NAND2_X1 U6075 ( .A1(n7932), .A2(n7933), .ZN(n4979) );
  INV_X1 U6076 ( .A(n10224), .ZN(n9944) );
  INV_X1 U6077 ( .A(n4596), .ZN(n7399) );
  INV_X1 U6078 ( .A(n7405), .ZN(n7725) );
  NOR2_X1 U6079 ( .A1(n10079), .A2(n10048), .ZN(n4896) );
  INV_X1 U6080 ( .A(n9723), .ZN(n10071) );
  NOR2_X1 U6081 ( .A1(n9985), .A2(n4659), .ZN(n9988) );
  OR2_X1 U6082 ( .A1(n9986), .A2(n4660), .ZN(n4659) );
  AND2_X1 U6083 ( .A1(n9987), .A2(n10261), .ZN(n4660) );
  INV_X1 U6084 ( .A(n9991), .ZN(n4899) );
  OAI21_X1 U6085 ( .B1(n5933), .B2(n5932), .A(n5931), .ZN(n5937) );
  AND2_X1 U6086 ( .A1(n5139), .A2(n5177), .ZN(n4656) );
  NAND2_X1 U6088 ( .A1(n5863), .A2(n5189), .ZN(n4464) );
  AOI21_X1 U6089 ( .B1(n5187), .B2(n5188), .A(n4809), .ZN(n4808) );
  INV_X1 U6090 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10132) );
  XNOR2_X1 U6091 ( .A(n5855), .B(n5854), .ZN(n10135) );
  INV_X1 U6092 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8589) );
  INV_X1 U6093 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5860) );
  INV_X1 U6094 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8306) );
  OAI21_X1 U6095 ( .B1(n5642), .B2(n5043), .A(n5040), .ZN(n5669) );
  INV_X1 U6096 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8287) );
  INV_X1 U6097 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8240) );
  INV_X1 U6098 ( .A(n4294), .ZN(n8238) );
  INV_X1 U6099 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8108) );
  INV_X1 U6100 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n8811) );
  INV_X1 U6101 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7204) );
  INV_X1 U6102 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U6103 ( .A1(n4731), .A2(n4730), .ZN(n4729) );
  INV_X1 U6104 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n4731) );
  NAND2_X1 U6105 ( .A1(n5975), .A2(n7698), .ZN(n4510) );
  OAI22_X1 U6106 ( .A1(n8660), .A2(n5076), .B1(n5079), .B2(n5080), .ZN(n5075)
         );
  INV_X1 U6107 ( .A(n5073), .ZN(n5072) );
  NAND2_X1 U6108 ( .A1(n7428), .A2(n7427), .ZN(n7551) );
  INV_X1 U6109 ( .A(n4888), .ZN(n7307) );
  NAND2_X1 U6110 ( .A1(n4918), .A2(n9011), .ZN(n8996) );
  NAND2_X1 U6111 ( .A1(n4921), .A2(n6696), .ZN(n9071) );
  NAND2_X1 U6112 ( .A1(n4865), .A2(n4862), .ZN(n6704) );
  INV_X1 U6113 ( .A(n6684), .ZN(n4651) );
  AND2_X1 U6114 ( .A1(n9395), .A2(n9111), .ZN(n9119) );
  NAND2_X1 U6115 ( .A1(n9316), .A2(n9315), .ZN(n9318) );
  NOR2_X1 U6116 ( .A1(n7121), .A2(n7120), .ZN(n7122) );
  NAND2_X1 U6117 ( .A1(n9987), .A2(n9659), .ZN(n6417) );
  NAND2_X1 U6118 ( .A1(n4633), .A2(n9621), .ZN(n9594) );
  AOI21_X1 U6119 ( .B1(n5016), .B2(n4686), .A(n4683), .ZN(n9648) );
  NAND2_X1 U6120 ( .A1(n4685), .A2(n4684), .ZN(n4683) );
  AND2_X1 U6121 ( .A1(n4494), .A2(n4493), .ZN(n9772) );
  AOI21_X1 U6122 ( .B1(n9973), .B2(n9987), .A(n9771), .ZN(n4493) );
  OAI21_X1 U6123 ( .B1(n9985), .B2(n4310), .A(n9971), .ZN(n4494) );
  NAND2_X1 U6124 ( .A1(n10289), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6125 ( .A1(n9984), .A2(n10291), .ZN(n4943) );
  OAI21_X1 U6126 ( .B1(n7141), .B2(n10289), .A(n4989), .ZN(P1_U3550) );
  NOR2_X1 U6127 ( .A1(n4990), .A2(n4408), .ZN(n4989) );
  NOR2_X1 U6128 ( .A1(n10291), .A2(n7139), .ZN(n4990) );
  NAND2_X1 U6129 ( .A1(n4897), .A2(n4894), .ZN(P1_U3548) );
  NOR2_X1 U6130 ( .A1(n4896), .A2(n4895), .ZN(n4894) );
  OR2_X1 U6131 ( .A1(n10077), .A2(n10289), .ZN(n4897) );
  NOR2_X1 U6132 ( .A1(n10291), .A2(n9993), .ZN(n4895) );
  NAND2_X1 U6133 ( .A1(n4593), .A2(n4591), .ZN(P1_U3547) );
  AOI21_X1 U6134 ( .B1(n9790), .B2(n8281), .A(n4592), .ZN(n4591) );
  NOR2_X1 U6135 ( .A1(n10291), .A2(n9997), .ZN(n4592) );
  OAI21_X1 U6136 ( .B1(n7141), .B2(n10282), .A(n4597), .ZN(P1_U3518) );
  NOR2_X1 U6137 ( .A1(n4407), .A2(n4598), .ZN(n4597) );
  NOR2_X1 U6138 ( .A1(n10283), .A2(n7142), .ZN(n4598) );
  OAI21_X1 U6139 ( .B1(n10077), .B2(n10282), .A(n4620), .ZN(P1_U3516) );
  NOR2_X1 U6140 ( .A1(n4622), .A2(n4621), .ZN(n4620) );
  NOR2_X1 U6141 ( .A1(n10283), .A2(n10078), .ZN(n4621) );
  NOR2_X1 U6142 ( .A1(n10079), .A2(n10107), .ZN(n4622) );
  NAND2_X1 U6143 ( .A1(n9790), .A2(n8283), .ZN(n4605) );
  INV_X1 U6144 ( .A(n4510), .ZN(n6030) );
  XNOR2_X1 U6145 ( .A(n5054), .B(n4429), .ZN(n7078) );
  NOR2_X1 U6146 ( .A1(n8495), .A2(n8491), .ZN(n4303) );
  NAND2_X1 U6147 ( .A1(n5093), .A2(n6494), .ZN(n4304) );
  XNOR2_X1 U6148 ( .A(n5802), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6160) );
  AND2_X1 U6149 ( .A1(n6654), .A2(n7633), .ZN(n4305) );
  XNOR2_X1 U6150 ( .A(n6525), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8542) );
  INV_X1 U6151 ( .A(n8542), .ZN(n4742) );
  NAND2_X1 U6152 ( .A1(n4916), .A2(n9011), .ZN(n8994) );
  NAND2_X1 U6153 ( .A1(n4431), .A2(n7371), .ZN(n7486) );
  NAND2_X1 U6154 ( .A1(n9790), .A2(n5715), .ZN(n4306) );
  AND2_X1 U6155 ( .A1(n9196), .A2(n8491), .ZN(n9207) );
  INV_X1 U6156 ( .A(n9781), .ZN(n4696) );
  AND2_X1 U6157 ( .A1(n8602), .A2(n9233), .ZN(n4307) );
  INV_X1 U6158 ( .A(n6098), .ZN(n4780) );
  AND2_X1 U6159 ( .A1(n4570), .A2(n4385), .ZN(n4308) );
  AND2_X1 U6160 ( .A1(n5089), .A2(n8076), .ZN(n4309) );
  AND2_X1 U6161 ( .A1(n9986), .A2(n9871), .ZN(n4310) );
  INV_X1 U6162 ( .A(n8469), .ZN(n4847) );
  INV_X1 U6163 ( .A(n8494), .ZN(n4751) );
  AND2_X1 U6164 ( .A1(n5757), .A2(n5756), .ZN(n9778) );
  OAI21_X1 U6165 ( .B1(n4842), .B2(n4839), .A(n4371), .ZN(n4838) );
  XOR2_X1 U6166 ( .A(n9777), .B(n4696), .Z(n4311) );
  NAND2_X1 U6167 ( .A1(n9781), .A2(n4977), .ZN(n4976) );
  INV_X1 U6168 ( .A(n5049), .ZN(n5048) );
  OAI21_X1 U6169 ( .B1(n5052), .B2(n5050), .A(n5603), .ZN(n5049) );
  OR2_X1 U6170 ( .A1(n8583), .A2(n7329), .ZN(n4312) );
  OR2_X1 U6171 ( .A1(n4751), .A2(n8488), .ZN(n4313) );
  AND2_X1 U6172 ( .A1(n5125), .A2(n8483), .ZN(n4314) );
  AND2_X1 U6173 ( .A1(n5063), .A2(n4404), .ZN(n4315) );
  NOR2_X1 U6174 ( .A1(n10051), .A2(n9933), .ZN(n4316) );
  NAND2_X1 U6175 ( .A1(n5882), .A2(n5800), .ZN(n6165) );
  INV_X1 U6176 ( .A(n7316), .ZN(n4444) );
  INV_X1 U6177 ( .A(n8910), .ZN(n8912) );
  AND2_X1 U6178 ( .A1(n7071), .A2(n7070), .ZN(n5115) );
  INV_X1 U6179 ( .A(n8149), .ZN(n4912) );
  AND2_X1 U6180 ( .A1(n6636), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4317) );
  NAND2_X1 U6181 ( .A1(n5329), .A2(n5328), .ZN(n7868) );
  INV_X1 U6182 ( .A(n7868), .ZN(n4933) );
  INV_X1 U6183 ( .A(n9075), .ZN(n9066) );
  INV_X1 U6184 ( .A(n4302), .ZN(n6620) );
  CLKBUF_X1 U6185 ( .A(n8936), .Z(n4637) );
  NAND2_X1 U6186 ( .A1(n6608), .A2(n9080), .ZN(n6696) );
  NAND2_X1 U6187 ( .A1(n5366), .A2(n5368), .ZN(n4318) );
  OR2_X1 U6188 ( .A1(n6568), .A2(n6767), .ZN(n4319) );
  OR2_X1 U6189 ( .A1(n6628), .A2(n6767), .ZN(n4320) );
  INV_X1 U6190 ( .A(n9913), .ZN(n4781) );
  INV_X1 U6191 ( .A(n8411), .ZN(n4849) );
  OR2_X1 U6192 ( .A1(n9847), .A2(n9846), .ZN(n9845) );
  OR2_X1 U6193 ( .A1(n7143), .A2(n6176), .ZN(n4322) );
  INV_X1 U6194 ( .A(n5068), .ZN(n5067) );
  NOR2_X1 U6195 ( .A1(n4290), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n4323) );
  NOR2_X1 U6196 ( .A1(n9646), .A2(n5014), .ZN(n4324) );
  NOR2_X1 U6197 ( .A1(n9464), .A2(n9247), .ZN(n4325) );
  NAND2_X1 U6198 ( .A1(n6856), .A2(n6855), .ZN(n7068) );
  OR2_X1 U6199 ( .A1(n9786), .A2(n9780), .ZN(n4326) );
  INV_X1 U6200 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6535) );
  OR3_X1 U6201 ( .A1(n9825), .A2(n4788), .A3(n9625), .ZN(n4328) );
  AND2_X2 U6202 ( .A1(n7143), .A2(n6167), .ZN(n6185) );
  NAND2_X1 U6203 ( .A1(n9857), .A2(n5918), .ZN(n9834) );
  NAND2_X1 U6204 ( .A1(n4969), .A2(n5556), .ZN(n9903) );
  NAND2_X1 U6205 ( .A1(n6729), .A2(n6728), .ZN(n6773) );
  OR2_X1 U6206 ( .A1(n9427), .A2(n9158), .ZN(n8498) );
  OR2_X1 U6207 ( .A1(n6428), .A2(n9662), .ZN(n4329) );
  XNOR2_X1 U6208 ( .A(n6575), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7633) );
  INV_X1 U6209 ( .A(n9987), .ZN(n4699) );
  INV_X1 U6210 ( .A(n5604), .ZN(n5051) );
  OR2_X1 U6211 ( .A1(n8210), .A2(n9276), .ZN(n4330) );
  AND2_X1 U6212 ( .A1(n4837), .A2(n4836), .ZN(n4331) );
  AND4_X1 U6213 ( .A1(n6073), .A2(n6072), .A3(n6071), .A4(n6070), .ZN(n4332)
         );
  NAND2_X1 U6214 ( .A1(n6925), .A2(n6924), .ZN(n9208) );
  NAND2_X1 U6215 ( .A1(n6536), .A2(n5090), .ZN(n4333) );
  NAND2_X1 U6216 ( .A1(n5650), .A2(n5649), .ZN(n10009) );
  INV_X1 U6217 ( .A(n9157), .ZN(n4520) );
  NAND2_X1 U6218 ( .A1(n9116), .A2(n8641), .ZN(n4334) );
  AND3_X1 U6219 ( .A1(n5230), .A2(n5231), .A3(n4960), .ZN(n4336) );
  AND2_X1 U6220 ( .A1(n7147), .A2(P2_D_REG_0__SCAN_IN), .ZN(n4337) );
  AND2_X1 U6221 ( .A1(n6090), .A2(n5993), .ZN(n4338) );
  NOR2_X1 U6222 ( .A1(n9301), .A2(n7824), .ZN(n4339) );
  AND2_X1 U6223 ( .A1(n8579), .A2(n8535), .ZN(n4340) );
  AND3_X1 U6224 ( .A1(n8513), .A2(n8512), .A3(n9122), .ZN(n4341) );
  INV_X1 U6225 ( .A(n4882), .ZN(n4881) );
  OAI21_X1 U6226 ( .B1(n4305), .B2(n7634), .A(n4883), .ZN(n4882) );
  AND2_X1 U6227 ( .A1(n4779), .A2(n4338), .ZN(n4342) );
  INV_X1 U6228 ( .A(n5832), .ZN(n10055) );
  AND2_X1 U6229 ( .A1(n5090), .A2(n6542), .ZN(n4343) );
  AND2_X1 U6230 ( .A1(n10031), .A2(n9883), .ZN(n4344) );
  INV_X1 U6231 ( .A(n9825), .ZN(n10091) );
  NAND2_X1 U6232 ( .A1(n5672), .A2(n5671), .ZN(n9825) );
  AND2_X1 U6233 ( .A1(n5062), .A2(n5065), .ZN(n4345) );
  AND2_X1 U6234 ( .A1(n7175), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4346) );
  AND2_X1 U6235 ( .A1(n9140), .A2(n8507), .ZN(n4347) );
  AND2_X1 U6236 ( .A1(n5835), .A2(n5967), .ZN(n4348) );
  OR2_X1 U6237 ( .A1(n6353), .A2(n6352), .ZN(n4349) );
  INV_X1 U6238 ( .A(n8565), .ZN(n9245) );
  AND2_X1 U6239 ( .A1(n7796), .A2(n7794), .ZN(n4350) );
  AND2_X1 U6240 ( .A1(n6251), .A2(n6247), .ZN(n4351) );
  AND2_X1 U6241 ( .A1(n6152), .A2(n6004), .ZN(n6147) );
  AND2_X1 U6242 ( .A1(n5135), .A2(n5917), .ZN(n4352) );
  OR2_X1 U6243 ( .A1(n6066), .A2(n6065), .ZN(n4353) );
  AND2_X1 U6244 ( .A1(n4618), .A2(n4617), .ZN(n4354) );
  INV_X1 U6245 ( .A(n5115), .ZN(n4572) );
  OR2_X1 U6246 ( .A1(n8605), .A2(n9209), .ZN(n4355) );
  INV_X1 U6247 ( .A(n7731), .ZN(n4475) );
  NAND2_X1 U6248 ( .A1(n9739), .A2(n7126), .ZN(n4356) );
  AND2_X1 U6249 ( .A1(n9825), .A2(n9835), .ZN(n4357) );
  AND2_X1 U6250 ( .A1(n4516), .A2(n4347), .ZN(n4358) );
  INV_X1 U6251 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n4730) );
  NAND2_X1 U6252 ( .A1(n8292), .A2(n8293), .ZN(n4359) );
  NAND4_X1 U6253 ( .A1(n6794), .A2(n6793), .A3(n6792), .A4(n6791), .ZN(n8932)
         );
  AND2_X1 U6254 ( .A1(n6308), .A2(n6307), .ZN(n4360) );
  OR2_X1 U6255 ( .A1(n5863), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4361) );
  NOR2_X1 U6256 ( .A1(n8128), .A2(n9675), .ZN(n4362) );
  INV_X1 U6257 ( .A(n4702), .ZN(n4701) );
  NAND2_X1 U6258 ( .A1(n4703), .A2(n5534), .ZN(n4702) );
  AND2_X1 U6259 ( .A1(n5046), .A2(n4700), .ZN(n4363) );
  AND2_X1 U6260 ( .A1(n8370), .A2(n8320), .ZN(n4364) );
  INV_X1 U6261 ( .A(n4845), .ZN(n4844) );
  NOR2_X1 U6262 ( .A1(n6937), .A2(n9221), .ZN(n4845) );
  INV_X1 U6263 ( .A(n5144), .ZN(n4694) );
  INV_X1 U6264 ( .A(n5016), .ZN(n9644) );
  OAI21_X1 U6265 ( .B1(n4995), .B2(n4488), .A(n4486), .ZN(n5016) );
  AND2_X1 U6266 ( .A1(n9397), .A2(n9124), .ZN(n4365) );
  AND2_X1 U6267 ( .A1(n5514), .A2(SI_15_), .ZN(n4366) );
  NAND2_X1 U6268 ( .A1(n4873), .A2(n4871), .ZN(n4367) );
  NOR2_X1 U6269 ( .A1(n7068), .A2(n8928), .ZN(n4368) );
  NAND2_X1 U6270 ( .A1(n5150), .A2(n5022), .ZN(n4369) );
  NOR2_X1 U6271 ( .A1(n9987), .A2(n4698), .ZN(n4370) );
  AND2_X1 U6272 ( .A1(n6968), .A2(n9168), .ZN(n4371) );
  INV_X1 U6273 ( .A(n5002), .ZN(n5001) );
  NAND2_X1 U6274 ( .A1(n5003), .A2(n9579), .ZN(n5002) );
  INV_X1 U6275 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n4806) );
  OR2_X1 U6276 ( .A1(n5816), .A2(n4944), .ZN(n4372) );
  OAI21_X1 U6277 ( .B1(n9511), .B2(n4998), .A(n4996), .ZN(n9589) );
  AND2_X1 U6278 ( .A1(n4548), .A2(n4547), .ZN(n4373) );
  NAND2_X1 U6279 ( .A1(n6115), .A2(n6117), .ZN(n9781) );
  OR2_X1 U6280 ( .A1(n6424), .A2(n7476), .ZN(n4374) );
  NAND2_X1 U6281 ( .A1(n8258), .A2(n6243), .ZN(n4375) );
  AND2_X1 U6282 ( .A1(n8619), .A2(n8906), .ZN(n4376) );
  AND2_X1 U6283 ( .A1(n4851), .A2(n4849), .ZN(n4377) );
  OR2_X1 U6284 ( .A1(n5214), .A2(n5213), .ZN(n4378) );
  NOR2_X1 U6285 ( .A1(n6655), .A2(n7184), .ZN(n4379) );
  OR2_X1 U6286 ( .A1(n9339), .A2(n8829), .ZN(n8493) );
  AND2_X1 U6287 ( .A1(n6567), .A2(n6569), .ZN(n6767) );
  NAND2_X1 U6288 ( .A1(n4520), .A2(n4518), .ZN(n4380) );
  INV_X1 U6289 ( .A(n9763), .ZN(n4697) );
  NAND2_X1 U6290 ( .A1(n9845), .A2(n5660), .ZN(n9818) );
  OR2_X1 U6291 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n7453), .ZN(n4381) );
  AND2_X1 U6292 ( .A1(n4850), .A2(n4849), .ZN(n4382) );
  AND2_X1 U6293 ( .A1(n7973), .A2(n6039), .ZN(n4383) );
  AND2_X1 U6294 ( .A1(n6093), .A2(n5968), .ZN(n4384) );
  NAND2_X1 U6295 ( .A1(n9464), .A2(n8334), .ZN(n4385) );
  NAND2_X1 U6296 ( .A1(n5440), .A2(n5439), .ZN(n5450) );
  INV_X1 U6297 ( .A(n5450), .ZN(n9551) );
  NAND2_X1 U6298 ( .A1(n8537), .A2(n8408), .ZN(n8570) );
  INV_X1 U6299 ( .A(n8570), .ZN(n4619) );
  AND2_X1 U6300 ( .A1(n8565), .A2(n4834), .ZN(n4386) );
  INV_X1 U6301 ( .A(n4840), .ZN(n4839) );
  NOR2_X1 U6302 ( .A1(n9197), .A2(n4845), .ZN(n4840) );
  NAND2_X1 U6303 ( .A1(n5915), .A2(n6121), .ZN(n9763) );
  NOR2_X1 U6304 ( .A1(n5471), .A2(n8247), .ZN(n4387) );
  AND2_X1 U6305 ( .A1(n4750), .A2(n4753), .ZN(n4388) );
  AND2_X1 U6306 ( .A1(n6213), .A2(n7731), .ZN(n4389) );
  AND2_X1 U6307 ( .A1(n9939), .A2(n9918), .ZN(n6074) );
  NAND2_X1 U6308 ( .A1(n6136), .A2(n10250), .ZN(n4390) );
  OR2_X1 U6309 ( .A1(n7527), .A2(n6471), .ZN(n4391) );
  OR2_X1 U6310 ( .A1(n7169), .A2(n7618), .ZN(n4392) );
  AND2_X1 U6311 ( .A1(n4309), .A2(n5088), .ZN(n4393) );
  AND2_X1 U6312 ( .A1(n5117), .A2(n8496), .ZN(n4394) );
  INV_X1 U6313 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5177) );
  AND2_X1 U6314 ( .A1(n5829), .A2(n6056), .ZN(n8118) );
  INV_X1 U6315 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6724) );
  INV_X1 U6316 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n6528) );
  INV_X1 U6317 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6726) );
  AND2_X1 U6318 ( .A1(n8470), .A2(n4849), .ZN(n4395) );
  INV_X1 U6319 ( .A(n7127), .ZN(n7124) );
  INV_X1 U6320 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6494) );
  INV_X1 U6321 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5022) );
  INV_X1 U6322 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6533) );
  AND2_X1 U6323 ( .A1(n8579), .A2(n4661), .ZN(n4396) );
  INV_X1 U6324 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4959) );
  XNOR2_X1 U6325 ( .A(n6514), .B(n6513), .ZN(n7085) );
  NOR2_X2 U6326 ( .A1(n8250), .A2(n5470), .ZN(n9949) );
  NAND2_X1 U6327 ( .A1(n5764), .A2(n5763), .ZN(n7140) );
  NOR2_X1 U6328 ( .A1(n8956), .A2(n8957), .ZN(n4397) );
  NAND2_X1 U6329 ( .A1(n6536), .A2(n4343), .ZN(n6609) );
  AND2_X1 U6330 ( .A1(n5017), .A2(n8360), .ZN(n4398) );
  AND2_X1 U6331 ( .A1(n4496), .A2(n8361), .ZN(n4399) );
  AND2_X1 U6332 ( .A1(n5008), .A2(n5012), .ZN(n4400) );
  NAND2_X2 U6333 ( .A1(n7619), .A2(n10221), .ZN(n9971) );
  OR2_X1 U6334 ( .A1(n8147), .A2(n8693), .ZN(n4401) );
  XOR2_X1 U6335 ( .A(n8604), .B(n8829), .Z(n4402) );
  NAND2_X1 U6336 ( .A1(n6517), .A2(n6523), .ZN(n8415) );
  INV_X1 U6337 ( .A(n8415), .ZN(n4743) );
  NAND2_X1 U6338 ( .A1(n4854), .A2(n6854), .ZN(n9275) );
  OAI21_X1 U6339 ( .B1(n5406), .B2(n7989), .A(n4963), .ZN(n8114) );
  NAND2_X1 U6340 ( .A1(n4476), .A2(n6218), .ZN(n7730) );
  NAND2_X1 U6341 ( .A1(n5406), .A2(n5405), .ZN(n7988) );
  NAND2_X1 U6342 ( .A1(n5116), .A2(n7070), .ZN(n8354) );
  NAND2_X1 U6343 ( .A1(n5083), .A2(n5084), .ZN(n8291) );
  NAND2_X1 U6344 ( .A1(n4979), .A2(n5364), .ZN(n7983) );
  OR2_X1 U6345 ( .A1(n8147), .A2(n8172), .ZN(n4403) );
  NAND2_X1 U6346 ( .A1(n4586), .A2(n7086), .ZN(n7089) );
  AND2_X1 U6347 ( .A1(n6588), .A2(n6585), .ZN(n8965) );
  OR2_X1 U6348 ( .A1(n8603), .A2(n8927), .ZN(n4404) );
  NAND2_X1 U6349 ( .A1(n5736), .A2(n5760), .ZN(n4405) );
  INV_X1 U6350 ( .A(n6866), .ZN(n9002) );
  NAND2_X1 U6351 ( .A1(n5143), .A2(n6069), .ZN(n8372) );
  AND2_X1 U6352 ( .A1(n4911), .A2(n8149), .ZN(n4406) );
  OAI21_X1 U6353 ( .B1(n7089), .B2(P2_D_REG_0__SCAN_IN), .A(n7147), .ZN(n7328)
         );
  NAND2_X1 U6354 ( .A1(n7795), .A2(n4350), .ZN(n7963) );
  NAND2_X1 U6355 ( .A1(n5111), .A2(n8462), .ZN(n9282) );
  NOR2_X1 U6357 ( .A1(n5812), .A2(n10107), .ZN(n4407) );
  NOR2_X1 U6358 ( .A1(n5812), .A2(n10048), .ZN(n4408) );
  NAND2_X1 U6359 ( .A1(n9949), .A2(n4929), .ZN(n4930) );
  AND2_X1 U6360 ( .A1(n4449), .A2(n9012), .ZN(n4409) );
  INV_X1 U6361 ( .A(n9790), .ZN(n10083) );
  NAND2_X1 U6362 ( .A1(n5706), .A2(n5705), .ZN(n9790) );
  OR2_X1 U6363 ( .A1(n9019), .A2(n6664), .ZN(n4410) );
  NAND2_X1 U6364 ( .A1(n5007), .A2(n5006), .ZN(n8260) );
  OR2_X1 U6365 ( .A1(n10087), .A2(n9630), .ZN(n4411) );
  OR2_X1 U6366 ( .A1(n6661), .A2(n6590), .ZN(n4412) );
  AND2_X1 U6367 ( .A1(n6417), .A2(n6416), .ZN(n4413) );
  AND2_X1 U6368 ( .A1(n4716), .A2(n4715), .ZN(n4414) );
  AND2_X1 U6369 ( .A1(n4719), .A2(n4718), .ZN(n4415) );
  INV_X1 U6370 ( .A(n4885), .ZN(n4884) );
  NOR2_X1 U6371 ( .A1(n6658), .A2(n7200), .ZN(n4885) );
  INV_X1 U6372 ( .A(n10153), .ZN(n4831) );
  NOR2_X1 U6373 ( .A1(n7786), .A2(n4954), .ZN(n7625) );
  INV_X1 U6374 ( .A(n8800), .ZN(n5079) );
  NAND2_X1 U6375 ( .A1(n6766), .A2(n6765), .ZN(n8933) );
  INV_X1 U6376 ( .A(n8933), .ZN(n4624) );
  NOR2_X1 U6377 ( .A1(n7768), .A2(n10260), .ZN(n4416) );
  NOR2_X1 U6378 ( .A1(n6576), .A2(n7633), .ZN(n7778) );
  NOR2_X1 U6379 ( .A1(n4657), .A2(n8822), .ZN(n4417) );
  NAND2_X1 U6380 ( .A1(n7313), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7312) );
  AND2_X1 U6381 ( .A1(n5844), .A2(n5843), .ZN(n9916) );
  INV_X1 U6382 ( .A(n9916), .ZN(n9966) );
  AND2_X1 U6383 ( .A1(n4509), .A2(n4508), .ZN(n7615) );
  AND2_X1 U6384 ( .A1(n7919), .A2(n8438), .ZN(n8553) );
  INV_X1 U6385 ( .A(n8553), .ZN(n4555) );
  XOR2_X1 U6386 ( .A(n9058), .B(n9353), .Z(n4418) );
  NAND2_X1 U6387 ( .A1(n10278), .A2(n10277), .ZN(n10250) );
  INV_X1 U6388 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6600) );
  XNOR2_X1 U6389 ( .A(n7041), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8581) );
  INV_X1 U6390 ( .A(n8581), .ZN(n8099) );
  AOI21_X1 U6391 ( .B1(n7272), .B2(n4319), .A(n7271), .ZN(n7270) );
  NAND2_X1 U6392 ( .A1(n7531), .A2(n7532), .ZN(n4737) );
  INV_X1 U6393 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n4956) );
  NAND4_X1 U6394 ( .A1(n4656), .A2(n5140), .A3(n5174), .A4(n5175), .ZN(n10117)
         );
  INV_X1 U6395 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n4824) );
  INV_X1 U6396 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n4830) );
  INV_X1 U6397 ( .A(n10291), .ZN(n10289) );
  NAND3_X4 U6398 ( .A1(n4327), .A2(n4419), .A3(n7329), .ZN(n7357) );
  NAND3_X1 U6399 ( .A1(n4421), .A2(n7147), .A3(n7089), .ZN(n4420) );
  NAND3_X1 U6400 ( .A1(n5061), .A2(n4402), .A3(n5059), .ZN(n4426) );
  XNOR2_X1 U6401 ( .A(n4427), .B(n4402), .ZN(n8882) );
  INV_X1 U6402 ( .A(n7485), .ZN(n4437) );
  NAND2_X1 U6403 ( .A1(n5055), .A2(n4428), .ZN(n5058) );
  NAND2_X1 U6404 ( .A1(n7485), .A2(n7427), .ZN(n4428) );
  NOR2_X2 U6405 ( .A1(n7486), .A2(n7487), .ZN(n7485) );
  AOI21_X2 U6406 ( .B1(n8331), .B2(n8329), .A(n8330), .ZN(n8591) );
  NAND2_X1 U6407 ( .A1(n8078), .A2(n4393), .ZN(n4430) );
  NAND2_X1 U6408 ( .A1(n7367), .A2(n7366), .ZN(n4431) );
  NAND2_X1 U6409 ( .A1(n7359), .A2(n7358), .ZN(n4432) );
  NAND2_X1 U6410 ( .A1(n5058), .A2(n7554), .ZN(n7555) );
  NAND3_X1 U6411 ( .A1(n6521), .A2(n6532), .A3(n6499), .ZN(n6517) );
  AND4_X2 U6412 ( .A1(n5091), .A2(n5093), .A3(n5094), .A4(n5092), .ZN(n6532)
         );
  AND2_X1 U6413 ( .A1(n6498), .A2(n5097), .ZN(n4436) );
  NAND2_X1 U6414 ( .A1(n4437), .A2(n7375), .ZN(n7428) );
  NAND2_X1 U6415 ( .A1(n4437), .A2(n7373), .ZN(n7377) );
  NAND3_X1 U6416 ( .A1(n6561), .A2(n6562), .A3(n4381), .ZN(n4438) );
  NOR2_X1 U6417 ( .A1(n7218), .A2(n7219), .ZN(n7217) );
  NOR2_X1 U6418 ( .A1(n4443), .A2(n7778), .ZN(n7777) );
  NAND2_X1 U6419 ( .A1(n4923), .A2(n4443), .ZN(n4922) );
  NAND2_X1 U6420 ( .A1(n4454), .A2(n7232), .ZN(n6587) );
  NAND3_X1 U6421 ( .A1(n4908), .A2(n4909), .A3(n4403), .ZN(n4454) );
  NAND2_X1 U6422 ( .A1(n7932), .A2(n4980), .ZN(n4455) );
  NAND2_X1 U6423 ( .A1(n7849), .A2(n7850), .ZN(n4456) );
  AND2_X2 U6424 ( .A1(n5974), .A2(n7698), .ZN(n7683) );
  OAI22_X1 U6425 ( .A1(n5609), .A2(n7152), .B1(n5270), .B2(n9693), .ZN(n4459)
         );
  NAND2_X1 U6426 ( .A1(n10239), .A2(n9680), .ZN(n5974) );
  INV_X1 U6427 ( .A(n7604), .ZN(n9680) );
  NOR2_X2 U6428 ( .A1(n4460), .A2(n4323), .ZN(n7604) );
  NAND3_X1 U6429 ( .A1(n5184), .A2(n5185), .A3(n5183), .ZN(n4460) );
  OAI22_X2 U6430 ( .A1(n9878), .A2(n5602), .B1(n10027), .B2(n9668), .ZN(n9872)
         );
  NAND4_X1 U6431 ( .A1(n5852), .A2(n9742), .A3(n5853), .A4(n4463), .ZN(n9984)
         );
  NAND2_X2 U6432 ( .A1(n4808), .A2(n4464), .ZN(n8384) );
  OR2_X1 U6433 ( .A1(n7190), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n4466) );
  NOR2_X1 U6434 ( .A1(n7661), .A2(n7660), .ZN(n7659) );
  NAND3_X1 U6435 ( .A1(n4728), .A2(n5267), .A3(n4729), .ZN(n7155) );
  NAND2_X1 U6436 ( .A1(n9686), .A2(n6445), .ZN(n7543) );
  NAND2_X2 U6437 ( .A1(n5252), .A2(n4468), .ZN(n7401) );
  AND3_X1 U6438 ( .A1(n4471), .A2(n4470), .A3(n4469), .ZN(n4468) );
  AND2_X1 U6439 ( .A1(n4473), .A2(n4472), .ZN(n6172) );
  NAND2_X1 U6440 ( .A1(n6185), .A2(n7744), .ZN(n4472) );
  NAND2_X1 U6441 ( .A1(n4643), .A2(n6345), .ZN(n4473) );
  NAND2_X1 U6442 ( .A1(n7580), .A2(n4389), .ZN(n4474) );
  NAND2_X1 U6443 ( .A1(n9764), .A2(n4480), .ZN(n9765) );
  NAND2_X1 U6444 ( .A1(n4481), .A2(n9763), .ZN(n4480) );
  INV_X1 U6445 ( .A(n7990), .ZN(n4489) );
  NAND2_X1 U6446 ( .A1(n7885), .A2(n6061), .ZN(n7990) );
  NAND2_X2 U6447 ( .A1(n4491), .A2(n5819), .ZN(n7392) );
  OAI21_X1 U6448 ( .B1(n5943), .B2(n7400), .A(n4491), .ZN(n7402) );
  NAND2_X1 U6449 ( .A1(n7400), .A2(n5943), .ZN(n4491) );
  OAI21_X1 U6450 ( .B1(n8360), .B2(n4498), .A(n9539), .ZN(n4497) );
  OAI21_X2 U6451 ( .B1(n4495), .B2(n4497), .A(n9540), .ZN(n9542) );
  NAND2_X1 U6452 ( .A1(n5018), .A2(n8360), .ZN(n4496) );
  INV_X1 U6453 ( .A(n4502), .ZN(n4501) );
  NAND3_X1 U6454 ( .A1(n4950), .A2(n4951), .A3(n6637), .ZN(n4502) );
  XNOR2_X1 U6455 ( .A(n6628), .B(n4920), .ZN(n7209) );
  NAND3_X1 U6456 ( .A1(n4504), .A2(n4503), .A3(P2_IR_REG_2__SCAN_IN), .ZN(
        n6555) );
  INV_X1 U6457 ( .A(n4505), .ZN(n7786) );
  OR2_X1 U6458 ( .A1(n4506), .A2(n7633), .ZN(n4505) );
  NAND2_X1 U6459 ( .A1(n4506), .A2(n7633), .ZN(n4955) );
  NOR2_X1 U6460 ( .A1(n8948), .A2(n5156), .ZN(n4506) );
  NAND3_X1 U6461 ( .A1(n6029), .A2(n6033), .A3(n4507), .ZN(n4509) );
  NAND2_X1 U6462 ( .A1(n7615), .A2(n7610), .ZN(n5820) );
  NAND2_X1 U6463 ( .A1(n6029), .A2(n6027), .ZN(n5973) );
  INV_X1 U6464 ( .A(n5973), .ZN(n7684) );
  NAND2_X1 U6465 ( .A1(n4512), .A2(n4511), .ZN(n9062) );
  AOI21_X1 U6466 ( .B1(n9059), .B2(n4956), .A(n4418), .ZN(n4511) );
  NAND2_X1 U6467 ( .A1(n9033), .A2(n9059), .ZN(n4512) );
  NAND2_X1 U6468 ( .A1(n4655), .A2(n6887), .ZN(n4513) );
  INV_X1 U6469 ( .A(n5801), .ZN(n5805) );
  NOR2_X2 U6470 ( .A1(n5794), .A2(n4369), .ZN(n5801) );
  NAND2_X1 U6471 ( .A1(n5265), .A2(n4514), .ZN(n5210) );
  XNOR2_X1 U6472 ( .A(n5265), .B(n4514), .ZN(n7183) );
  NAND4_X1 U6473 ( .A1(n4517), .A2(n4662), .A3(n4539), .A4(n4540), .ZN(n4515)
         );
  NAND2_X1 U6474 ( .A1(n4528), .A2(n8588), .ZN(P2_U3296) );
  NAND4_X1 U6475 ( .A1(n4312), .A2(n4552), .A3(n4529), .A4(n4603), .ZN(n4528)
         );
  OAI21_X1 U6476 ( .B1(n4553), .B2(n8582), .A(n8580), .ZN(n4530) );
  NAND4_X1 U6477 ( .A1(n5028), .A2(n4535), .A3(n5027), .A4(n5319), .ZN(n4688)
         );
  NAND2_X1 U6478 ( .A1(n5221), .A2(n5028), .ZN(n5277) );
  AND2_X1 U6479 ( .A1(n4535), .A2(n4378), .ZN(n5221) );
  NAND2_X1 U6480 ( .A1(n5216), .A2(n5215), .ZN(n4535) );
  NAND2_X1 U6481 ( .A1(n4537), .A2(n4619), .ZN(n4551) );
  NAND2_X1 U6482 ( .A1(n4538), .A2(n8527), .ZN(n4537) );
  OAI21_X1 U6483 ( .B1(n4341), .B2(n4632), .A(n4706), .ZN(n4538) );
  NAND2_X1 U6484 ( .A1(n4746), .A2(n4748), .ZN(n4539) );
  NAND2_X1 U6485 ( .A1(n4744), .A2(n4610), .ZN(n4540) );
  OAI21_X1 U6486 ( .B1(n4541), .B2(n8459), .A(n8458), .ZN(n8467) );
  OAI21_X1 U6487 ( .B1(n4545), .B2(n4544), .A(n4543), .ZN(n4542) );
  NAND4_X1 U6488 ( .A1(n6532), .A2(n6506), .A3(n6521), .A4(n5126), .ZN(n9473)
         );
  NAND3_X1 U6489 ( .A1(n6532), .A2(n6521), .A3(n6506), .ZN(n6527) );
  INV_X1 U6490 ( .A(n4764), .ZN(n8530) );
  NAND2_X1 U6491 ( .A1(n4553), .A2(n4396), .ZN(n4552) );
  NAND2_X1 U6492 ( .A1(n8578), .A2(n8577), .ZN(n4553) );
  OR2_X1 U6493 ( .A1(n8531), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4628) );
  NAND2_X2 U6494 ( .A1(n7050), .A2(n6735), .ZN(n8531) );
  OAI211_X1 U6495 ( .C1(n4556), .C2(n4555), .A(n8444), .B(n4554), .ZN(n7065)
         );
  NAND2_X1 U6496 ( .A1(n4559), .A2(n4557), .ZN(n4561) );
  OR2_X1 U6497 ( .A1(n4562), .A2(n4560), .ZN(n4559) );
  NAND2_X1 U6498 ( .A1(n4562), .A2(n8517), .ZN(n9112) );
  OR2_X1 U6499 ( .A1(n9121), .A2(n8514), .ZN(n4562) );
  NAND4_X1 U6500 ( .A1(n6521), .A2(n6532), .A3(n6506), .A4(n6529), .ZN(n6723)
         );
  NOR2_X2 U6501 ( .A1(n6504), .A2(n6505), .ZN(n6506) );
  NAND2_X1 U6502 ( .A1(n7408), .A2(n8548), .ZN(n7060) );
  NAND2_X1 U6503 ( .A1(n8275), .A2(n4308), .ZN(n4565) );
  NAND2_X1 U6505 ( .A1(n5119), .A2(n4394), .ZN(n4581) );
  XNOR2_X1 U6506 ( .A(n4626), .B(n6528), .ZN(n6622) );
  AOI21_X2 U6507 ( .B1(n9244), .B2(n8479), .A(n7072), .ZN(n9228) );
  NAND2_X1 U6508 ( .A1(n8032), .A2(n8033), .ZN(n5111) );
  NAND2_X1 U6509 ( .A1(n7827), .A2(n8448), .ZN(n5114) );
  INV_X2 U6510 ( .A(n7952), .ZN(n7499) );
  NAND2_X1 U6512 ( .A1(n7295), .A2(n7296), .ZN(n4582) );
  NAND2_X1 U6513 ( .A1(n6915), .A2(n6914), .ZN(n9218) );
  NAND2_X1 U6514 ( .A1(n4331), .A2(n4583), .ZN(n6972) );
  NAND2_X2 U6515 ( .A1(n5239), .A2(n5238), .ZN(n5257) );
  NAND2_X1 U6516 ( .A1(n7764), .A2(n5821), .ZN(n5138) );
  NAND2_X1 U6517 ( .A1(n4585), .A2(n5818), .ZN(n6029) );
  AOI21_X2 U6518 ( .B1(n5851), .B2(n9966), .A(n4584), .ZN(n9742) );
  INV_X1 U6519 ( .A(n7392), .ZN(n4585) );
  NAND2_X1 U6520 ( .A1(n9880), .A2(n9881), .ZN(n9879) );
  OAI21_X2 U6521 ( .B1(n9850), .B2(n5639), .A(n5638), .ZN(n9847) );
  NAND2_X1 U6522 ( .A1(n9764), .A2(n5915), .ZN(n7128) );
  NAND2_X1 U6523 ( .A1(n9894), .A2(n6090), .ZN(n9880) );
  NAND2_X1 U6524 ( .A1(n6512), .A2(n6511), .ZN(n7083) );
  NAND2_X1 U6525 ( .A1(n7084), .A2(n7085), .ZN(n4586) );
  NAND2_X1 U6526 ( .A1(n8625), .A2(n8624), .ZN(n8648) );
  INV_X1 U6527 ( .A(n7736), .ZN(n4587) );
  AND2_X1 U6528 ( .A1(n6175), .A2(n6174), .ZN(n6178) );
  INV_X1 U6529 ( .A(n7610), .ZN(n7616) );
  OAI21_X1 U6530 ( .B1(n5298), .B2(n7158), .A(n4589), .ZN(n4588) );
  NAND2_X1 U6531 ( .A1(n7725), .A2(n7401), .ZN(n4596) );
  OR2_X1 U6532 ( .A1(n5751), .A2(n7741), .ZN(n5238) );
  INV_X2 U6533 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8733) );
  INV_X1 U6534 ( .A(n5943), .ZN(n4595) );
  MUX2_X1 U6535 ( .A(n10139), .B(n10136), .S(n5270), .Z(n7405) );
  NAND2_X1 U6536 ( .A1(n9996), .A2(n9995), .ZN(n4606) );
  NAND2_X1 U6537 ( .A1(n9984), .A2(n10283), .ZN(n5888) );
  INV_X2 U6538 ( .A(n5182), .ZN(n8388) );
  XNOR2_X2 U6539 ( .A(n5178), .B(P1_IR_REG_29__SCAN_IN), .ZN(n5182) );
  NAND2_X1 U6540 ( .A1(n9681), .A2(n10228), .ZN(n6027) );
  OAI21_X1 U6541 ( .B1(n8972), .B2(n8973), .A(n4412), .ZN(n8999) );
  NAND2_X1 U6542 ( .A1(n4599), .A2(n4682), .ZN(n4681) );
  NAND3_X1 U6543 ( .A1(n8485), .A2(n8483), .A3(n8546), .ZN(n4599) );
  NOR2_X2 U6544 ( .A1(n9826), .A2(n5839), .ZN(n9811) );
  NAND2_X1 U6545 ( .A1(n4680), .A2(n4679), .ZN(n8490) );
  NAND2_X1 U6546 ( .A1(n4934), .A2(n4931), .ZN(n7977) );
  INV_X1 U6547 ( .A(n8445), .ZN(n4615) );
  NOR2_X2 U6548 ( .A1(n9886), .A2(n10020), .ZN(n4940) );
  OAI21_X1 U6549 ( .B1(n4766), .B2(n4395), .A(n8562), .ZN(n4765) );
  NAND2_X2 U6550 ( .A1(n4600), .A2(n6906), .ZN(n9350) );
  NAND2_X1 U6551 ( .A1(n4374), .A2(n4601), .ZN(n7296) );
  NAND2_X1 U6552 ( .A1(n8185), .A2(n8186), .ZN(n8184) );
  NAND2_X1 U6553 ( .A1(n9684), .A2(n9683), .ZN(n9682) );
  NAND3_X1 U6554 ( .A1(n6491), .A2(n10215), .A3(n4602), .ZN(n4636) );
  NAND2_X2 U6555 ( .A1(n6381), .A2(n6422), .ZN(n6193) );
  INV_X1 U6556 ( .A(n6163), .ZN(n6167) );
  NAND2_X1 U6557 ( .A1(n9715), .A2(n4392), .ZN(n7644) );
  NAND2_X1 U6558 ( .A1(n4820), .A2(n6477), .ZN(n10202) );
  INV_X1 U6559 ( .A(n6188), .ZN(n4671) );
  NOR2_X1 U6560 ( .A1(n7812), .A2(n7813), .ZN(n7811) );
  NAND2_X1 U6561 ( .A1(n5203), .A2(n5240), .ZN(n5206) );
  NOR2_X1 U6562 ( .A1(n8025), .A2(n8024), .ZN(n8023) );
  OAI21_X1 U6563 ( .B1(n9139), .B2(n8504), .A(n8511), .ZN(n9121) );
  NAND3_X1 U6564 ( .A1(n4604), .A2(n6687), .A3(n4651), .ZN(P2_U3201) );
  NAND2_X1 U6565 ( .A1(n6686), .A2(n6685), .ZN(n4604) );
  NAND2_X1 U6566 ( .A1(n5114), .A2(n5112), .ZN(n8039) );
  AOI21_X1 U6567 ( .B1(n7310), .B2(n8945), .A(n8946), .ZN(n8948) );
  NOR2_X2 U6568 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n5165) );
  NAND2_X1 U6569 ( .A1(n10082), .A2(n4605), .ZN(P1_U3515) );
  NAND2_X1 U6570 ( .A1(n4607), .A2(n5276), .ZN(n7609) );
  NAND2_X1 U6571 ( .A1(n5274), .A2(n5275), .ZN(n4607) );
  NAND2_X1 U6572 ( .A1(n7231), .A2(n5744), .ZN(n5423) );
  NAND2_X1 U6573 ( .A1(n5417), .A2(n5434), .ZN(n7231) );
  AOI21_X1 U6574 ( .B1(n4963), .B2(n7989), .A(n8118), .ZN(n4961) );
  AND2_X2 U6575 ( .A1(n4687), .A2(n4688), .ZN(n5365) );
  NAND2_X1 U6576 ( .A1(n4609), .A2(n6685), .ZN(n6706) );
  NAND2_X1 U6577 ( .A1(n6692), .A2(n6693), .ZN(n4609) );
  INV_X1 U6578 ( .A(n6640), .ZN(n4655) );
  NAND2_X1 U6579 ( .A1(n4949), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4948) );
  INV_X2 U6580 ( .A(n5181), .ZN(n8633) );
  NAND3_X1 U6581 ( .A1(n8490), .A2(n4388), .A3(n8496), .ZN(n4610) );
  OAI211_X1 U6582 ( .C1(n4615), .C2(n4614), .A(n4613), .B(n4612), .ZN(n4611)
         );
  NAND2_X1 U6583 ( .A1(n4900), .A2(n4899), .ZN(n4898) );
  NAND2_X1 U6584 ( .A1(n7963), .A2(n7962), .ZN(n8078) );
  NAND2_X1 U6585 ( .A1(n8932), .A2(n4623), .ZN(n8438) );
  AND2_X1 U6586 ( .A1(n6763), .A2(n6762), .ZN(n5158) );
  OR2_X1 U6587 ( .A1(n6756), .A2(n7153), .ZN(n4629) );
  NAND2_X1 U6588 ( .A1(n9302), .A2(n9301), .ZN(n7827) );
  NAND2_X1 U6589 ( .A1(n8467), .A2(n8561), .ZN(n4769) );
  NAND2_X1 U6590 ( .A1(n6460), .A2(n6459), .ZN(n10208) );
  NOR2_X1 U6591 ( .A1(n10148), .A2(n4721), .ZN(n6455) );
  AOI21_X1 U6592 ( .B1(P1_REG1_REG_6__SCAN_IN), .B2(n7647), .A(n7640), .ZN(
        n7673) );
  NAND2_X1 U6593 ( .A1(n7542), .A2(n6447), .ZN(n9702) );
  NAND2_X1 U6594 ( .A1(n8477), .A2(n4630), .ZN(n8482) );
  AOI21_X1 U6595 ( .B1(n6487), .B2(n9871), .A(n6486), .ZN(n6493) );
  OR2_X1 U6596 ( .A1(n5322), .A2(SI_5_), .ZN(n5323) );
  NAND2_X1 U6597 ( .A1(n8487), .A2(n4756), .ZN(n4679) );
  AOI21_X1 U6598 ( .B1(n8077), .B2(n8076), .A(n5087), .ZN(n5086) );
  NOR2_X1 U6599 ( .A1(n10150), .A2(n10149), .ZN(n10148) );
  NOR2_X1 U6600 ( .A1(n8021), .A2(n8022), .ZN(n8020) );
  AOI22_X2 U6601 ( .A1(n8834), .A2(n8833), .B1(n9194), .B2(n8607), .ZN(n8652)
         );
  NAND2_X1 U6602 ( .A1(n5799), .A2(n5857), .ZN(n5882) );
  NAND2_X1 U6603 ( .A1(n5149), .A2(n6428), .ZN(n6441) );
  NAND2_X1 U6604 ( .A1(n4636), .A2(n7856), .ZN(n6492) );
  NAND2_X1 U6605 ( .A1(n9717), .A2(n9718), .ZN(n9715) );
  NAND2_X1 U6606 ( .A1(n7508), .A2(n4822), .ZN(n7812) );
  XNOR2_X1 U6607 ( .A(n5193), .B(n5225), .ZN(n9693) );
  NOR2_X1 U6608 ( .A1(n7811), .A2(n4644), .ZN(n8025) );
  NOR2_X1 U6609 ( .A1(n8023), .A2(n4827), .ZN(n8185) );
  NAND2_X1 U6610 ( .A1(n10186), .A2(n10188), .ZN(n4820) );
  NAND2_X1 U6611 ( .A1(n4283), .A2(n5268), .ZN(n5192) );
  NAND2_X1 U6612 ( .A1(n5331), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5357) );
  NAND2_X1 U6613 ( .A1(n4988), .A2(n4674), .ZN(n4673) );
  INV_X2 U6614 ( .A(n5186), .ZN(n5140) );
  NAND2_X1 U6615 ( .A1(n6101), .A2(n6151), .ZN(n4801) );
  NAND2_X1 U6616 ( .A1(n4797), .A2(n6111), .ZN(n4796) );
  AOI21_X1 U6617 ( .B1(n4815), .B2(n4814), .A(n4812), .ZN(n4811) );
  NAND2_X1 U6618 ( .A1(n7528), .A2(n4391), .ZN(n9717) );
  NAND2_X1 U6619 ( .A1(n7509), .A2(n7510), .ZN(n7508) );
  NAND2_X1 U6620 ( .A1(n4784), .A2(n4783), .ZN(n6142) );
  NOR2_X1 U6621 ( .A1(n10176), .A2(n4821), .ZN(n10186) );
  NOR2_X1 U6622 ( .A1(n6475), .A2(n10162), .ZN(n10178) );
  NAND2_X1 U6623 ( .A1(n6059), .A2(n4786), .ZN(n6062) );
  INV_X1 U6624 ( .A(n6581), .ZN(n4914) );
  NOR2_X1 U6625 ( .A1(n10147), .A2(n10146), .ZN(n10145) );
  OAI211_X1 U6626 ( .C1(n6026), .C2(n4788), .A(n7683), .B(n4819), .ZN(n6032)
         );
  INV_X1 U6627 ( .A(n6064), .ZN(n4817) );
  OAI21_X1 U6628 ( .B1(n6038), .B2(n4791), .A(n4383), .ZN(n4790) );
  NAND2_X1 U6629 ( .A1(n5067), .A2(n8857), .ZN(n5066) );
  OAI21_X1 U6630 ( .B1(n8857), .B2(n8858), .A(n8601), .ZN(n5068) );
  NAND2_X1 U6631 ( .A1(n4649), .A2(n6625), .ZN(n7224) );
  NAND3_X1 U6632 ( .A1(n6561), .A2(n6562), .A3(n4958), .ZN(n4649) );
  AOI21_X1 U6633 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(n4766) );
  NAND2_X1 U6634 ( .A1(n8417), .A2(n4741), .ZN(n4740) );
  INV_X2 U6635 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5194) );
  NOR2_X1 U6636 ( .A1(n9757), .A2(n4673), .ZN(n7141) );
  INV_X1 U6637 ( .A(n9511), .ZN(n4654) );
  XNOR2_X1 U6638 ( .A(n6463), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U6639 ( .A1(n7543), .A2(n7544), .ZN(n7542) );
  NOR2_X1 U6640 ( .A1(n7808), .A2(n4725), .ZN(n8022) );
  NOR2_X1 U6641 ( .A1(n7671), .A2(n4727), .ZN(n7661) );
  NOR2_X1 U6642 ( .A1(n8338), .A2(n4723), .ZN(n10150) );
  INV_X1 U6643 ( .A(n6189), .ZN(n4672) );
  NAND2_X1 U6644 ( .A1(n4672), .A2(n4671), .ZN(n6190) );
  OAI21_X1 U6645 ( .B1(n8140), .B2(n8142), .A(n8141), .ZN(n8144) );
  XNOR2_X1 U6646 ( .A(n6170), .B(n6177), .ZN(n4993) );
  NAND2_X1 U6647 ( .A1(n9598), .A2(n6330), .ZN(n5021) );
  OR2_X1 U6648 ( .A1(n7911), .A2(n7836), .ZN(n6781) );
  NAND2_X1 U6649 ( .A1(n9289), .A2(n4339), .ZN(n7821) );
  AOI21_X1 U6650 ( .B1(n9132), .B2(n6997), .A(n5147), .ZN(n9123) );
  NAND2_X1 U6651 ( .A1(n6972), .A2(n5145), .ZN(n9144) );
  NAND2_X1 U6652 ( .A1(n4848), .A2(n4846), .ZN(n8351) );
  NAND2_X1 U6653 ( .A1(n4943), .A2(n5129), .ZN(P1_U3551) );
  NOR2_X1 U6654 ( .A1(n6782), .A2(n8426), .ZN(n6783) );
  NAND2_X1 U6655 ( .A1(n6181), .A2(n6180), .ZN(n7456) );
  NOR2_X2 U6656 ( .A1(n5478), .A2(n5173), .ZN(n5498) );
  AOI22_X2 U6657 ( .A1(n8869), .A2(n8886), .B1(n8867), .B2(n8868), .ZN(n8872)
         );
  XNOR2_X2 U6658 ( .A(n8866), .B(n8868), .ZN(n8869) );
  NAND2_X1 U6659 ( .A1(n6638), .A2(n9020), .ZN(n9025) );
  AOI21_X1 U6660 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(n8915) );
  INV_X1 U6661 ( .A(n5190), .ZN(n4809) );
  AOI21_X1 U6662 ( .B1(n8816), .B2(n9376), .A(n8812), .ZN(n7119) );
  NAND2_X1 U6663 ( .A1(n4919), .A2(n6866), .ZN(n4918) );
  NAND2_X1 U6664 ( .A1(n6605), .A2(n6887), .ZN(n6606) );
  NAND2_X1 U6665 ( .A1(n6557), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n6560) );
  NOR2_X1 U6666 ( .A1(n7217), .A2(n6564), .ZN(n7241) );
  NAND2_X1 U6667 ( .A1(n6586), .A2(n6587), .ZN(n8956) );
  NAND2_X2 U6668 ( .A1(n9803), .A2(n5840), .ZN(n9806) );
  NAND2_X1 U6669 ( .A1(n4665), .A2(n4413), .ZN(P1_U3214) );
  NAND2_X1 U6670 ( .A1(n4666), .A2(n9621), .ZN(n4665) );
  NAND2_X1 U6671 ( .A1(n6392), .A2(n6418), .ZN(n4666) );
  BUF_X2 U6672 ( .A(n5251), .Z(n4667) );
  NOR2_X1 U6673 ( .A1(n8159), .A2(n8160), .ZN(n8140) );
  NAND2_X1 U6674 ( .A1(n4669), .A2(n8164), .ZN(n4668) );
  INV_X1 U6675 ( .A(n6633), .ZN(n4669) );
  XNOR2_X2 U6676 ( .A(n4807), .B(n4806), .ZN(n10125) );
  NAND2_X1 U6677 ( .A1(n9992), .A2(n10250), .ZN(n4900) );
  XNOR2_X2 U6678 ( .A(n6725), .B(n9474), .ZN(n8820) );
  NAND3_X1 U6679 ( .A1(n9594), .A2(n9593), .A3(n4411), .ZN(P1_U3229) );
  XNOR2_X1 U6680 ( .A(n5865), .B(n5864), .ZN(n10131) );
  OAI21_X1 U6681 ( .B1(n6052), .B2(n6051), .A(n6058), .ZN(n6055) );
  NAND3_X1 U6682 ( .A1(n5138), .A2(n5826), .A3(n5827), .ZN(n7885) );
  NAND2_X1 U6683 ( .A1(n6141), .A2(n6140), .ZN(n4784) );
  AOI21_X1 U6684 ( .B1(n4796), .B2(n4795), .A(n4794), .ZN(n6127) );
  NAND2_X1 U6685 ( .A1(n4800), .A2(n4798), .ZN(n4797) );
  NAND2_X1 U6686 ( .A1(n6102), .A2(n4788), .ZN(n4802) );
  NAND2_X1 U6687 ( .A1(n6113), .A2(n5130), .ZN(n5132) );
  NAND2_X1 U6688 ( .A1(n4818), .A2(n6033), .ZN(n6034) );
  NAND2_X1 U6689 ( .A1(n4778), .A2(n4775), .ZN(n6096) );
  NAND2_X1 U6690 ( .A1(n6050), .A2(n6151), .ZN(n4793) );
  NAND2_X1 U6691 ( .A1(n6132), .A2(n6131), .ZN(n4785) );
  XNOR2_X2 U6692 ( .A(n8934), .B(n7409), .ZN(n8548) );
  NAND2_X1 U6693 ( .A1(n5495), .A2(n5494), .ZN(n5031) );
  NAND2_X1 U6694 ( .A1(n5031), .A2(n5497), .ZN(n5513) );
  NAND2_X1 U6695 ( .A1(n4962), .A2(n4961), .ZN(n8242) );
  NOR2_X1 U6696 ( .A1(n9990), .A2(n4898), .ZN(n10077) );
  NAND3_X1 U6697 ( .A1(n4762), .A2(n4760), .A3(n8574), .ZN(n8583) );
  NAND2_X1 U6698 ( .A1(n5132), .A2(n4697), .ZN(n9764) );
  NAND2_X2 U6699 ( .A1(n5353), .A2(n5352), .ZN(n8235) );
  NAND3_X1 U6700 ( .A1(n5026), .A2(n5323), .A3(n5324), .ZN(n4689) );
  NAND2_X1 U6701 ( .A1(n5365), .A2(n5372), .ZN(n4906) );
  NAND2_X1 U6702 ( .A1(n4689), .A2(n5326), .ZN(n4687) );
  INV_X1 U6703 ( .A(n5222), .ZN(n5028) );
  NAND2_X1 U6704 ( .A1(n5392), .A2(n4693), .ZN(n4692) );
  NAND3_X1 U6705 ( .A1(n4697), .A2(n4696), .A3(n4695), .ZN(n5962) );
  NAND2_X1 U6706 ( .A1(n5535), .A2(n5534), .ZN(n5542) );
  NOR2_X2 U6707 ( .A1(n6961), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n4714) );
  NAND2_X1 U6708 ( .A1(n6717), .A2(n4414), .ZN(n6898) );
  NAND2_X1 U6709 ( .A1(n6719), .A2(n4415), .ZN(n6940) );
  NAND3_X1 U6710 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n4728) );
  INV_X1 U6711 ( .A(n4757), .ZN(n4759) );
  OAI21_X1 U6712 ( .B1(n8530), .B2(n4761), .A(n8515), .ZN(n4760) );
  NAND2_X1 U6713 ( .A1(n4764), .A2(n4763), .ZN(n4762) );
  NAND3_X1 U6714 ( .A1(n4765), .A2(n8473), .A3(n8563), .ZN(n8477) );
  NAND2_X1 U6715 ( .A1(n4770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6727) );
  NAND4_X1 U6716 ( .A1(n6521), .A2(n6532), .A3(n6506), .A4(n5127), .ZN(n4770)
         );
  INV_X1 U6717 ( .A(n4771), .ZN(n6100) );
  OAI22_X1 U6718 ( .A1(n4773), .A2(n4772), .B1(n4384), .B2(n4774), .ZN(n4771)
         );
  NAND2_X1 U6719 ( .A1(n6087), .A2(n4781), .ZN(n4778) );
  AOI21_X1 U6720 ( .B1(n6089), .B2(n4777), .A(n4776), .ZN(n4775) );
  INV_X1 U6721 ( .A(n6088), .ZN(n4782) );
  AOI21_X2 U6722 ( .B1(n4785), .B2(n6136), .A(n6135), .ZN(n6141) );
  NAND3_X1 U6723 ( .A1(n4790), .A2(n6041), .A3(n6040), .ZN(n4789) );
  NAND3_X1 U6724 ( .A1(n4802), .A2(n4801), .A3(n9846), .ZN(n4800) );
  NAND2_X1 U6725 ( .A1(n6158), .A2(n4805), .ZN(P1_U3242) );
  NAND2_X1 U6726 ( .A1(n4811), .A2(n4810), .ZN(n6086) );
  OR2_X1 U6727 ( .A1(n6077), .A2(n6076), .ZN(n4810) );
  OAI21_X1 U6728 ( .B1(n6032), .B2(n6031), .A(n6030), .ZN(n4818) );
  NAND2_X1 U6729 ( .A1(n9256), .A2(n6894), .ZN(n4833) );
  NAND2_X1 U6730 ( .A1(n4833), .A2(n4386), .ZN(n6904) );
  NAND2_X1 U6731 ( .A1(n9206), .A2(n4835), .ZN(n4837) );
  NAND2_X1 U6732 ( .A1(n6845), .A2(n4382), .ZN(n4848) );
  OAI21_X1 U6733 ( .B1(n6845), .B2(n4851), .A(n4850), .ZN(n8271) );
  NAND2_X1 U6734 ( .A1(n6845), .A2(n6844), .ZN(n8034) );
  NAND2_X1 U6735 ( .A1(n6844), .A2(n4330), .ZN(n4856) );
  NAND2_X1 U6736 ( .A1(n7009), .A2(n4859), .ZN(n4858) );
  NAND2_X1 U6737 ( .A1(n4858), .A2(n4857), .ZN(n7058) );
  NAND2_X1 U6738 ( .A1(n7009), .A2(n5148), .ZN(n9104) );
  OR3_X1 U6739 ( .A1(n4282), .A2(n4879), .A3(n4875), .ZN(n4872) );
  AND2_X2 U6740 ( .A1(n4870), .A2(n4869), .ZN(n8967) );
  OR4_X2 U6741 ( .A1(n7635), .A2(n4879), .A3(n4875), .A4(n4885), .ZN(n4870) );
  NAND2_X1 U6742 ( .A1(n6657), .A2(n8164), .ZN(n4886) );
  MUX2_X1 U6743 ( .A(P2_REG1_REG_0__SCAN_IN), .B(P2_REG2_REG_0__SCAN_IN), .S(
        n7043), .Z(n7256) );
  MUX2_X1 U6744 ( .A(P2_REG1_REG_1__SCAN_IN), .B(P2_REG2_REG_1__SCAN_IN), .S(
        n7043), .Z(n6647) );
  NAND2_X2 U6745 ( .A1(n5564), .A2(n5563), .ZN(n10031) );
  INV_X2 U6746 ( .A(n5298), .ZN(n4893) );
  XNOR2_X1 U6747 ( .A(n4904), .B(n9873), .ZN(n9868) );
  OAI21_X1 U6748 ( .B1(n5997), .B2(n4904), .A(n6117), .ZN(n5913) );
  OAI21_X1 U6749 ( .B1(n5365), .B2(n4318), .A(n5372), .ZN(n5390) );
  NAND2_X1 U6750 ( .A1(n8150), .A2(n8149), .ZN(n4908) );
  NAND3_X1 U6751 ( .A1(n4913), .A2(n6582), .A3(P2_REG2_REG_9__SCAN_IN), .ZN(
        n4915) );
  NAND3_X1 U6752 ( .A1(n4913), .A2(n6582), .A3(n4910), .ZN(n4909) );
  INV_X1 U6753 ( .A(n4915), .ZN(n8148) );
  NAND2_X1 U6754 ( .A1(n4922), .A2(n7776), .ZN(n7780) );
  INV_X1 U6755 ( .A(n7778), .ZN(n4923) );
  NAND2_X1 U6756 ( .A1(n5142), .A2(n5498), .ZN(n5190) );
  NAND2_X1 U6757 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  AND2_X2 U6758 ( .A1(n4927), .A2(n9949), .ZN(n9938) );
  INV_X1 U6759 ( .A(n4930), .ZN(n9937) );
  INV_X1 U6760 ( .A(n7768), .ZN(n4934) );
  INV_X1 U6761 ( .A(n9786), .ZN(n4936) );
  NAND2_X1 U6762 ( .A1(n4936), .A2(n4937), .ZN(n7135) );
  INV_X1 U6763 ( .A(n7135), .ZN(n5813) );
  NAND2_X1 U6764 ( .A1(n4941), .A2(n4940), .ZN(n9826) );
  NOR2_X1 U6765 ( .A1(n5159), .A2(n10014), .ZN(n9852) );
  NOR2_X1 U6766 ( .A1(n6632), .A2(n6631), .ZN(n7311) );
  NAND2_X1 U6767 ( .A1(n8945), .A2(n4945), .ZN(n7310) );
  INV_X1 U6768 ( .A(n6642), .ZN(n4946) );
  INV_X1 U6769 ( .A(n6691), .ZN(n4947) );
  NAND2_X1 U6770 ( .A1(n4946), .A2(n6905), .ZN(n4949) );
  OR2_X1 U6771 ( .A1(n4948), .A2(n4947), .ZN(n6688) );
  NAND2_X1 U6772 ( .A1(n4948), .A2(n6691), .ZN(n6644) );
  NAND2_X1 U6773 ( .A1(n8978), .A2(n8977), .ZN(n4950) );
  NAND3_X1 U6774 ( .A1(n4953), .A2(n4952), .A3(n6636), .ZN(n4951) );
  AND2_X1 U6775 ( .A1(n8977), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4952) );
  NAND2_X1 U6776 ( .A1(n4953), .A2(n6636), .ZN(n8960) );
  INV_X1 U6777 ( .A(n9033), .ZN(n4957) );
  INV_X1 U6778 ( .A(n9679), .ZN(n7577) );
  NAND2_X2 U6779 ( .A1(n5232), .A2(n4336), .ZN(n9679) );
  NAND2_X1 U6780 ( .A1(n5406), .A2(n4963), .ZN(n4962) );
  INV_X1 U6781 ( .A(n5716), .ZN(n4977) );
  NAND4_X1 U6782 ( .A1(n5140), .A2(n5174), .A3(n5139), .A4(n5175), .ZN(n5141)
         );
  NAND3_X1 U6783 ( .A1(n9739), .A2(n7126), .A3(n10250), .ZN(n4988) );
  NAND2_X1 U6784 ( .A1(n4991), .A2(n7457), .ZN(n7472) );
  NAND2_X1 U6785 ( .A1(n4993), .A2(n6172), .ZN(n7457) );
  NAND2_X1 U6786 ( .A1(n4992), .A2(n6171), .ZN(n4991) );
  INV_X1 U6787 ( .A(n4993), .ZN(n4992) );
  NAND2_X1 U6788 ( .A1(n9511), .A2(n4996), .ZN(n4995) );
  NAND2_X1 U6789 ( .A1(n7862), .A2(n5009), .ZN(n5007) );
  INV_X1 U6790 ( .A(n5012), .ZN(n5011) );
  OR2_X1 U6791 ( .A1(n7864), .A2(n7863), .ZN(n5013) );
  NOR2_X1 U6792 ( .A1(n6386), .A2(n6387), .ZN(n5015) );
  NAND2_X1 U6793 ( .A1(n5021), .A2(n5019), .ZN(n6341) );
  NAND2_X1 U6794 ( .A1(n5797), .A2(n5150), .ZN(n5803) );
  INV_X1 U6795 ( .A(n5321), .ZN(n5026) );
  NAND2_X1 U6796 ( .A1(n5495), .A2(n5032), .ZN(n5029) );
  OAI21_X1 U6797 ( .B1(n7156), .B2(n5036), .A(n5255), .ZN(n5240) );
  NAND2_X1 U6798 ( .A1(n5642), .A2(n5641), .ZN(n5039) );
  INV_X1 U6799 ( .A(n5056), .ZN(n5055) );
  OAI21_X1 U6800 ( .B1(n7375), .B2(n5057), .A(n7550), .ZN(n5056) );
  INV_X1 U6801 ( .A(n7427), .ZN(n5057) );
  NAND2_X1 U6802 ( .A1(n4315), .A2(n8847), .ZN(n5061) );
  NAND3_X1 U6803 ( .A1(n5063), .A2(n5064), .A3(n4404), .ZN(n5060) );
  NAND2_X1 U6804 ( .A1(n8869), .A2(n5070), .ZN(n5069) );
  OAI211_X1 U6805 ( .C1(n8869), .C2(n5072), .A(n5075), .B(n5069), .ZN(P2_U3156) );
  INV_X1 U6806 ( .A(n8660), .ZN(n5080) );
  INV_X1 U6807 ( .A(n6609), .ZN(n6611) );
  INV_X1 U6808 ( .A(n8416), .ZN(n5099) );
  NAND3_X1 U6809 ( .A1(n8570), .A2(n5105), .A3(n5106), .ZN(n5102) );
  OAI211_X1 U6810 ( .C1(n5105), .C2(n8570), .A(n5103), .B(n5102), .ZN(n8816)
         );
  NAND2_X1 U6811 ( .A1(n5104), .A2(n4619), .ZN(n5103) );
  OAI21_X1 U6812 ( .B1(n9112), .B2(n9113), .A(n8520), .ZN(n9099) );
  NAND2_X1 U6813 ( .A1(n9113), .A2(n8520), .ZN(n5107) );
  NAND2_X1 U6814 ( .A1(n8526), .A2(n9105), .ZN(n5108) );
  NAND2_X1 U6815 ( .A1(n5111), .A2(n5109), .ZN(n9281) );
  NAND3_X1 U6816 ( .A1(n7075), .A2(n5121), .A3(n5122), .ZN(n5118) );
  NAND2_X1 U6817 ( .A1(n9228), .A2(n5120), .ZN(n5119) );
  NOR2_X1 U6818 ( .A1(n6074), .A2(n9913), .ZN(n5128) );
  NAND3_X1 U6819 ( .A1(n9806), .A2(n5131), .A3(n6115), .ZN(n5130) );
  OR2_X1 U6820 ( .A1(n9846), .A2(n5137), .ZN(n5136) );
  NOR2_X1 U6821 ( .A1(n5186), .A2(n5166), .ZN(n5142) );
  NOR2_X2 U6822 ( .A1(n5166), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n5139) );
  INV_X1 U6823 ( .A(n6125), .ZN(n6024) );
  NAND2_X1 U6824 ( .A1(n6558), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6559) );
  NAND2_X1 U6825 ( .A1(n6160), .A2(n8110), .ZN(n6163) );
  BUF_X4 U6826 ( .A(n7156), .Z(n5298) );
  NAND2_X1 U6827 ( .A1(n9765), .A2(n9966), .ZN(n9770) );
  XNOR2_X1 U6828 ( .A(n9391), .B(n9105), .ZN(n9100) );
  NAND2_X1 U6829 ( .A1(n8544), .A2(n8543), .ZN(n8578) );
  NAND2_X1 U6830 ( .A1(n8820), .A2(n6728), .ZN(n6788) );
  CLKBUF_X1 U6831 ( .A(n8847), .Z(n8859) );
  OAI21_X1 U6832 ( .B1(n6128), .B2(n6127), .A(n6126), .ZN(n6132) );
  NAND4_X2 U6833 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n5186)
         );
  NAND2_X1 U6834 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  AND2_X1 U6835 ( .A1(n5410), .A2(SI_10_), .ZN(n5144) );
  INV_X1 U6836 ( .A(n9662), .ZN(n9621) );
  OR2_X1 U6837 ( .A1(n6412), .A2(n6391), .ZN(n9662) );
  AND3_X1 U6838 ( .A1(n5895), .A2(n5773), .A3(n5896), .ZN(n5146) );
  INV_X1 U6839 ( .A(n7286), .ZN(n7178) );
  NAND2_X1 U6840 ( .A1(n9551), .A2(n5449), .ZN(n5829) );
  AND2_X1 U6841 ( .A1(n9131), .A2(n8906), .ZN(n5147) );
  OR2_X1 U6842 ( .A1(n7008), .A2(n8628), .ZN(n5148) );
  AND3_X1 U6843 ( .A1(n6418), .A2(n9621), .A3(n6429), .ZN(n5149) );
  AND2_X1 U6844 ( .A1(n5796), .A2(n5795), .ZN(n5150) );
  INV_X1 U6845 ( .A(n8984), .ZN(n6590) );
  AND2_X1 U6846 ( .A1(n5391), .A2(n5376), .ZN(n5151) );
  NOR2_X1 U6847 ( .A1(n9790), .A2(n5715), .ZN(n5716) );
  INV_X1 U6848 ( .A(n6136), .ZN(n9740) );
  AND3_X2 U6849 ( .A1(n7137), .A2(n7613), .A3(n7611), .ZN(n10283) );
  INV_X1 U6850 ( .A(n9932), .ZN(n9960) );
  AND3_X1 U6851 ( .A1(n8570), .A2(n8519), .A3(n9295), .ZN(n5153) );
  INV_X1 U6852 ( .A(n8556), .ZN(n7066) );
  OR2_X1 U6853 ( .A1(n7783), .A2(n7958), .ZN(n5154) );
  OR2_X1 U6854 ( .A1(n7783), .A2(n8709), .ZN(n5155) );
  AND2_X1 U6855 ( .A1(n7175), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5156) );
  INV_X1 U6856 ( .A(n7133), .ZN(n9762) );
  AND2_X1 U6857 ( .A1(n9307), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5160) );
  NAND2_X2 U6858 ( .A1(n7451), .A2(n9238), .ZN(n9296) );
  AND2_X1 U6859 ( .A1(n7118), .A2(n7117), .ZN(n10301) );
  INV_X1 U6860 ( .A(n10260), .ZN(n5811) );
  INV_X1 U6861 ( .A(n6029), .ZN(n6031) );
  NOR4_X1 U6862 ( .A1(n9781), .A2(n9792), .A3(n6021), .A4(n6151), .ZN(n6022)
         );
  INV_X1 U6863 ( .A(n9810), .ZN(n5715) );
  AND2_X1 U6864 ( .A1(n7253), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6565) );
  NOR2_X1 U6865 ( .A1(n9510), .A2(n9618), .ZN(n6352) );
  OR2_X1 U6866 ( .A1(n6876), .A2(n6879), .ZN(n6599) );
  INV_X1 U6867 ( .A(n4288), .ZN(n6371) );
  INV_X1 U6868 ( .A(n7140), .ZN(n5812) );
  AND2_X1 U6869 ( .A1(n5760), .A2(n5759), .ZN(n5761) );
  INV_X1 U6870 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5559) );
  INV_X1 U6871 ( .A(SI_9_), .ZN(n5373) );
  INV_X1 U6872 ( .A(n9289), .ZN(n7822) );
  INV_X1 U6873 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5398) );
  INV_X1 U6874 ( .A(n5505), .ZN(n5503) );
  NAND2_X1 U6875 ( .A1(n9733), .A2(n6151), .ZN(n6137) );
  AOI22_X1 U6876 ( .A1(n9665), .A2(n9932), .B1(n9725), .B2(n9664), .ZN(n5850)
         );
  INV_X1 U6877 ( .A(n8375), .ZN(n5834) );
  INV_X1 U6878 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5795) );
  INV_X1 U6879 ( .A(SI_11_), .ZN(n5411) );
  INV_X1 U6880 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6716) );
  NAND2_X1 U6881 ( .A1(n6590), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6591) );
  OR2_X1 U6882 ( .A1(n8004), .A2(n8071), .ZN(n8433) );
  OR2_X1 U6883 ( .A1(n6597), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n6598) );
  INV_X1 U6884 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5547) );
  OAI22_X1 U6885 ( .A1(n9778), .A2(n9960), .B1(n9962), .B2(n7729), .ZN(n7130)
         );
  NAND2_X1 U6886 ( .A1(n5519), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5548) );
  AND2_X1 U6887 ( .A1(n5808), .A2(n7717), .ZN(n5809) );
  AND2_X1 U6888 ( .A1(n10113), .A2(n6401), .ZN(n5885) );
  INV_X1 U6889 ( .A(n5544), .ZN(n5515) );
  INV_X1 U6890 ( .A(n5451), .ZN(n5455) );
  NAND2_X1 U6891 ( .A1(n7156), .A2(n7167), .ZN(n5199) );
  OR2_X1 U6892 ( .A1(n4297), .A2(n7447), .ZN(n7330) );
  INV_X1 U6893 ( .A(n8616), .ZN(n8617) );
  INV_X1 U6894 ( .A(n7556), .ZN(n7557) );
  INV_X1 U6895 ( .A(n9208), .ZN(n9233) );
  AND2_X1 U6896 ( .A1(n8041), .A2(n8040), .ZN(n8558) );
  NAND2_X1 U6897 ( .A1(n6620), .A2(n8099), .ZN(n8534) );
  AND2_X1 U6898 ( .A1(n7328), .A2(n7103), .ZN(n7116) );
  INV_X1 U6899 ( .A(n8545), .ZN(n9152) );
  OR2_X1 U6900 ( .A1(n8534), .A2(n4743), .ZN(n8008) );
  AND2_X1 U6901 ( .A1(n7331), .A2(n7350), .ZN(n7349) );
  OR2_X1 U6902 ( .A1(n6412), .A2(n6409), .ZN(n9643) );
  AND3_X1 U6903 ( .A1(n5892), .A2(n5891), .A3(n5890), .ZN(n5965) );
  OR2_X1 U6904 ( .A1(n4290), .A2(n7722), .ZN(n5252) );
  NAND2_X1 U6905 ( .A1(n6489), .A2(n10211), .ZN(n6491) );
  INV_X1 U6906 ( .A(n6063), .ZN(n6056) );
  INV_X1 U6907 ( .A(n7846), .ZN(n5315) );
  INV_X1 U6908 ( .A(n7389), .ZN(n7391) );
  AND2_X1 U6909 ( .A1(n9725), .A2(n9724), .ZN(n9980) );
  NAND2_X1 U6910 ( .A1(n5689), .A2(n5688), .ZN(n5839) );
  NAND2_X1 U6911 ( .A1(n6444), .A2(n4675), .ZN(n9962) );
  XNOR2_X1 U6912 ( .A(n5894), .B(n5893), .ZN(n7021) );
  AND2_X1 U6913 ( .A1(n5626), .A2(n5608), .ZN(n5624) );
  XNOR2_X1 U6914 ( .A(n5533), .B(SI_16_), .ZN(n5530) );
  INV_X1 U6915 ( .A(n8918), .ZN(n8902) );
  AND2_X1 U6916 ( .A1(n6913), .A2(n6912), .ZN(n9220) );
  INV_X1 U6917 ( .A(n9060), .ZN(n6685) );
  NAND2_X1 U6918 ( .A1(n9110), .A2(n9299), .ZN(n9111) );
  AND2_X1 U6919 ( .A1(n9296), .A2(n7835), .ZN(n9303) );
  INV_X1 U6920 ( .A(n9310), .ZN(n9356) );
  AND2_X1 U6921 ( .A1(n8415), .A2(n4742), .ZN(n9378) );
  INV_X1 U6922 ( .A(n8563), .ZN(n9255) );
  INV_X1 U6923 ( .A(n8805), .ZN(n9463) );
  NAND2_X1 U6924 ( .A1(n8050), .A2(n8008), .ZN(n9376) );
  OR2_X1 U6925 ( .A1(n7089), .A2(P2_D_REG_1__SCAN_IN), .ZN(n7088) );
  NAND2_X1 U6926 ( .A1(n6437), .A2(n6436), .ZN(n6438) );
  XNOR2_X1 U6927 ( .A(n5883), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7298) );
  INV_X1 U6928 ( .A(n4290), .ZN(n5793) );
  AND3_X1 U6929 ( .A1(n5509), .A2(n5508), .A3(n5507), .ZN(n9963) );
  NAND2_X1 U6930 ( .A1(n6490), .A2(n6481), .ZN(n10206) );
  INV_X1 U6931 ( .A(n10215), .ZN(n10168) );
  INV_X1 U6932 ( .A(n9929), .ZN(n10231) );
  AND2_X1 U6933 ( .A1(n6394), .A2(n5884), .ZN(n10261) );
  INV_X1 U6934 ( .A(n10250), .ZN(n10265) );
  NAND2_X1 U6935 ( .A1(n5867), .A2(n5866), .ZN(n10114) );
  NAND2_X1 U6936 ( .A1(n5590), .A2(n5796), .ZN(n5591) );
  AND2_X1 U6937 ( .A1(n5303), .A2(n5349), .ZN(n7647) );
  INV_X2 U6938 ( .A(n7050), .ZN(n6929) );
  OR2_X1 U6939 ( .A1(n7348), .A2(n7346), .ZN(n8918) );
  AND2_X1 U6940 ( .A1(n7326), .A2(n7325), .ZN(n8910) );
  INV_X1 U6941 ( .A(n9043), .ZN(n9086) );
  INV_X1 U6942 ( .A(n9296), .ZN(n9273) );
  INV_X1 U6943 ( .A(n9303), .ZN(n9264) );
  NOR2_X1 U6944 ( .A1(n7107), .A2(n5160), .ZN(n7108) );
  INV_X1 U6945 ( .A(n9332), .ZN(n9359) );
  NAND2_X1 U6946 ( .A1(n7105), .A2(n7104), .ZN(n9307) );
  OR2_X1 U6947 ( .A1(n10301), .A2(n7830), .ZN(n9467) );
  AND3_X1 U6948 ( .A1(n9374), .A2(n9373), .A3(n9372), .ZN(n10299) );
  INV_X2 U6949 ( .A(n10301), .ZN(n10298) );
  AND2_X1 U6950 ( .A1(n7088), .A2(n7087), .ZN(n9472) );
  AND2_X1 U6951 ( .A1(n8308), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7149) );
  INV_X1 U6952 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n9495) );
  INV_X1 U6953 ( .A(n8965), .ZN(n7232) );
  INV_X1 U6954 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7180) );
  INV_X1 U6955 ( .A(n7298), .ZN(n7144) );
  INV_X1 U6956 ( .A(n10009), .ZN(n9839) );
  INV_X1 U6957 ( .A(n9917), .ZN(n9883) );
  INV_X1 U6958 ( .A(n10141), .ZN(n10220) );
  OR2_X1 U6959 ( .A1(n7619), .A2(n7856), .ZN(n10224) );
  OR2_X1 U6960 ( .A1(n4287), .A2(n7621), .ZN(n10227) );
  NAND2_X1 U6961 ( .A1(n10291), .A2(n10261), .ZN(n10048) );
  AND2_X2 U6962 ( .A1(n7138), .A2(n7137), .ZN(n10291) );
  INV_X1 U6963 ( .A(n9780), .ZN(n10079) );
  NAND2_X1 U6964 ( .A1(n10283), .A2(n10261), .ZN(n10107) );
  INV_X1 U6965 ( .A(n10283), .ZN(n10282) );
  INV_X1 U6966 ( .A(n10235), .ZN(n10236) );
  AND2_X1 U6967 ( .A1(n10114), .A2(n10113), .ZN(n10235) );
  INV_X1 U6968 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7264) );
  INV_X1 U6969 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n7236) );
  INV_X1 U6970 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10306) );
  INV_X1 U6971 ( .A(n8935), .ZN(P2_U3893) );
  AND2_X2 U6972 ( .A1(n7145), .A2(n7144), .ZN(P1_U3973) );
  NAND2_X1 U6973 ( .A1(n6493), .A2(n6492), .ZN(P1_U3262) );
  NAND2_X1 U6974 ( .A1(n5888), .A2(n5887), .ZN(P1_U3519) );
  AND3_X2 U6975 ( .A1(n8679), .A2(n5022), .A3(n5586), .ZN(n5164) );
  NOR2_X1 U6976 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5163) );
  NOR2_X1 U6977 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5162) );
  NOR2_X1 U6978 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5161) );
  INV_X2 U6979 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5854) );
  NAND3_X1 U6980 ( .A1(n5165), .A2(n8733), .A3(n5854), .ZN(n5166) );
  NOR2_X2 U6981 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5170) );
  NOR2_X2 U6982 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5169) );
  NOR2_X2 U6983 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n5168) );
  INV_X1 U6986 ( .A(n5173), .ZN(n5174) );
  XNOR2_X2 U6987 ( .A(n5176), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5181) );
  NAND2_X2 U6988 ( .A1(n5181), .A2(n8388), .ZN(n5251) );
  INV_X1 U6989 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5179) );
  NAND2_X2 U6990 ( .A1(n8633), .A2(n5182), .ZN(n5330) );
  INV_X1 U6991 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6448) );
  OR2_X1 U6992 ( .A1(n5330), .A2(n6448), .ZN(n5184) );
  INV_X1 U6993 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5180) );
  OR2_X1 U6994 ( .A1(n4296), .A2(n5180), .ZN(n5183) );
  AND2_X1 U6995 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5189) );
  NAND3_X1 U6996 ( .A1(n5854), .A2(n5864), .A3(P1_IR_REG_27__SCAN_IN), .ZN(
        n5188) );
  XNOR2_X1 U6997 ( .A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_27__SCAN_IN), .ZN(
        n5187) );
  NAND2_X1 U6998 ( .A1(n5192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5193) );
  NAND3_X1 U6999 ( .A1(n5196), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n5197) );
  NAND2_X4 U7000 ( .A1(n5198), .A2(n5197), .ZN(n7156) );
  INV_X1 U7001 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8678) );
  INV_X1 U7002 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n7167) );
  INV_X1 U7004 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U7005 ( .A1(n7156), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5201) );
  INV_X1 U7006 ( .A(SI_1_), .ZN(n5200) );
  OAI211_X1 U7007 ( .C1(n7156), .C2(n7158), .A(n5201), .B(n5200), .ZN(n5203)
         );
  AND2_X1 U7008 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5202) );
  NAND2_X1 U7009 ( .A1(n7156), .A2(n5202), .ZN(n5255) );
  INV_X1 U7010 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7154) );
  NAND2_X1 U7011 ( .A1(n7156), .A2(n7154), .ZN(n5204) );
  OAI211_X1 U7012 ( .C1(n5298), .C2(P1_DATAO_REG_1__SCAN_IN), .A(n5204), .B(
        SI_1_), .ZN(n5205) );
  INV_X1 U7013 ( .A(n5207), .ZN(n5208) );
  NAND2_X1 U7014 ( .A1(n5208), .A2(SI_2_), .ZN(n5209) );
  NAND2_X1 U7015 ( .A1(n5210), .A2(n5209), .ZN(n5216) );
  MUX2_X1 U7016 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .S(n7156), .Z(n5212) );
  XNOR2_X1 U7017 ( .A(n5216), .B(n5211), .ZN(n7151) );
  INV_X1 U7018 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7152) );
  NAND2_X1 U7019 ( .A1(n7604), .A2(n10239), .ZN(n7702) );
  INV_X1 U7020 ( .A(n5211), .ZN(n5215) );
  INV_X1 U7021 ( .A(n5212), .ZN(n5214) );
  INV_X1 U7022 ( .A(SI_3_), .ZN(n5213) );
  INV_X1 U7023 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5217) );
  INV_X1 U7024 ( .A(SI_4_), .ZN(n8677) );
  INV_X1 U7025 ( .A(n5218), .ZN(n5219) );
  NAND2_X1 U7026 ( .A1(n5219), .A2(SI_4_), .ZN(n5220) );
  NAND2_X1 U7027 ( .A1(n5318), .A2(n5220), .ZN(n5222) );
  INV_X1 U7028 ( .A(n5221), .ZN(n5223) );
  NAND2_X1 U7029 ( .A1(n5223), .A2(n5222), .ZN(n5224) );
  NAND2_X1 U7030 ( .A1(n5277), .A2(n5224), .ZN(n7146) );
  NAND2_X1 U7031 ( .A1(n7146), .A2(n5744), .ZN(n5229) );
  INV_X2 U7032 ( .A(n5270), .ZN(n6443) );
  NAND2_X1 U7033 ( .A1(n5227), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5280) );
  XNOR2_X1 U7034 ( .A(n5280), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U7035 ( .A1(n5306), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5232) );
  INV_X1 U7036 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6471) );
  OR2_X1 U7037 ( .A1(n4667), .A2(n6471), .ZN(n5231) );
  XNOR2_X1 U7038 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n7706) );
  OR2_X1 U7039 ( .A1(n4290), .A2(n7706), .ZN(n5230) );
  INV_X1 U7041 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6450) );
  INV_X1 U7042 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5233) );
  OR2_X1 U7043 ( .A1(n4295), .A2(n5233), .ZN(n5236) );
  INV_X1 U7044 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5234) );
  AND3_X2 U7045 ( .A1(n5237), .A2(n5236), .A3(n5235), .ZN(n5239) );
  INV_X1 U7046 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7741) );
  INV_X1 U7047 ( .A(n5191), .ZN(n5267) );
  INV_X1 U7048 ( .A(n7155), .ZN(n9685) );
  NAND2_X1 U7049 ( .A1(n8384), .A2(n9685), .ZN(n5248) );
  XNOR2_X1 U7050 ( .A(n5240), .B(SI_1_), .ZN(n5241) );
  NAND2_X1 U7051 ( .A1(n7153), .A2(n5035), .ZN(n5243) );
  NAND2_X1 U7052 ( .A1(n4893), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5242) );
  NAND2_X1 U7053 ( .A1(n5243), .A2(n5242), .ZN(n5244) );
  INV_X2 U7054 ( .A(n8384), .ZN(n5846) );
  NAND2_X1 U7055 ( .A1(n4893), .A2(n7154), .ZN(n5245) );
  OAI211_X1 U7056 ( .C1(n7153), .C2(n4893), .A(n5846), .B(n5245), .ZN(n5246)
         );
  XNOR2_X2 U7057 ( .A(n5257), .B(n7744), .ZN(n5943) );
  INV_X1 U7058 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6176) );
  INV_X1 U7059 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5249) );
  INV_X1 U7060 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5250) );
  INV_X1 U7061 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7722) );
  INV_X1 U7062 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10139) );
  INV_X1 U7063 ( .A(SI_0_), .ZN(n5254) );
  INV_X1 U7064 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5253) );
  OAI21_X1 U7065 ( .B1(n4893), .B2(n5254), .A(n5253), .ZN(n5256) );
  NAND2_X1 U7066 ( .A1(n5256), .A2(n5255), .ZN(n10136) );
  OR2_X1 U7067 ( .A1(n5257), .A2(n7744), .ZN(n5258) );
  NAND2_X1 U7068 ( .A1(n5653), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5264) );
  INV_X1 U7069 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6467) );
  INV_X1 U7070 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10222) );
  OR2_X1 U7071 ( .A1(n4290), .A2(n10222), .ZN(n5262) );
  INV_X1 U7072 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5259) );
  OR2_X1 U7073 ( .A1(n5260), .A2(n5259), .ZN(n5261) );
  NAND4_X2 U7074 ( .A1(n5264), .A2(n5263), .A3(n5262), .A4(n5261), .ZN(n9681)
         );
  INV_X1 U7075 ( .A(n7183), .ZN(n5266) );
  NAND2_X1 U7076 ( .A1(n5278), .A2(n5266), .ZN(n5272) );
  NAND2_X1 U7077 ( .A1(n5267), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5269) );
  OR2_X1 U7078 ( .A1(n5270), .A2(n7538), .ZN(n5271) );
  OR2_X2 U7079 ( .A1(n9681), .A2(n10228), .ZN(n5818) );
  NAND2_X2 U7080 ( .A1(n5818), .A2(n6027), .ZN(n7389) );
  INV_X1 U7081 ( .A(n9681), .ZN(n7475) );
  NAND2_X1 U7082 ( .A1(n7475), .A2(n10228), .ZN(n7686) );
  NAND2_X1 U7083 ( .A1(n7687), .A2(n5273), .ZN(n5274) );
  INV_X1 U7084 ( .A(n7708), .ZN(n10245) );
  NAND2_X1 U7085 ( .A1(n10245), .A2(n7577), .ZN(n5276) );
  INV_X1 U7086 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7187) );
  INV_X1 U7087 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7170) );
  XNOR2_X1 U7088 ( .A(n5295), .B(SI_5_), .ZN(n5294) );
  NAND2_X1 U7089 ( .A1(n7168), .A2(n5744), .ZN(n5284) );
  NAND2_X1 U7090 ( .A1(n5280), .A2(n5279), .ZN(n5281) );
  NAND2_X1 U7091 ( .A1(n5281), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5282) );
  AOI22_X1 U7092 ( .A1(n5593), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6443), .B2(
        n9714), .ZN(n5283) );
  NAND2_X1 U7093 ( .A1(n5306), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5291) );
  INV_X1 U7094 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7618) );
  OR2_X1 U7095 ( .A1(n4667), .A2(n7618), .ZN(n5290) );
  INV_X1 U7096 ( .A(n5307), .ZN(n5309) );
  INV_X1 U7097 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5286) );
  NAND2_X1 U7098 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5285) );
  NAND2_X1 U7099 ( .A1(n5286), .A2(n5285), .ZN(n5287) );
  NAND2_X1 U7100 ( .A1(n5309), .A2(n5287), .ZN(n7762) );
  OR2_X1 U7101 ( .A1(n4290), .A2(n7762), .ZN(n5289) );
  INV_X1 U7102 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6451) );
  OR2_X1 U7103 ( .A1(n5330), .A2(n6451), .ZN(n5288) );
  NAND2_X1 U7104 ( .A1(n10253), .A2(n7736), .ZN(n6037) );
  NAND2_X1 U7105 ( .A1(n7609), .A2(n7616), .ZN(n5293) );
  OR2_X1 U7106 ( .A1(n10253), .A2(n4587), .ZN(n5292) );
  NAND2_X1 U7107 ( .A1(n5293), .A2(n5292), .ZN(n7763) );
  INV_X1 U7108 ( .A(n5294), .ZN(n5296) );
  MUX2_X1 U7109 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n7156), .Z(n5325) );
  XNOR2_X1 U7110 ( .A(n5299), .B(n5321), .ZN(n7159) );
  NAND2_X1 U7111 ( .A1(n7159), .A2(n5744), .ZN(n5305) );
  NOR2_X1 U7112 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5300) );
  NAND2_X1 U7113 ( .A1(n5301), .A2(n5300), .ZN(n5479) );
  NAND2_X1 U7114 ( .A1(n5479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5302) );
  MUX2_X1 U7115 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5302), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5303) );
  AOI22_X1 U7116 ( .A1(n5593), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6443), .B2(
        n7647), .ZN(n5304) );
  NAND2_X1 U7117 ( .A1(n5306), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5314) );
  INV_X1 U7118 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7767) );
  OR2_X1 U7119 ( .A1(n4667), .A2(n7767), .ZN(n5313) );
  INV_X1 U7120 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U7121 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U7122 ( .A1(n5333), .A2(n5310), .ZN(n7769) );
  OR2_X1 U7123 ( .A1(n4290), .A2(n7769), .ZN(n5312) );
  INV_X1 U7124 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6452) );
  OR2_X1 U7125 ( .A1(n5889), .A2(n6452), .ZN(n5311) );
  OR2_X1 U7126 ( .A1(n10260), .A2(n7756), .ZN(n7845) );
  AND2_X2 U7127 ( .A1(n10260), .A2(n7756), .ZN(n7846) );
  NAND2_X1 U7128 ( .A1(n7845), .A2(n5315), .ZN(n7765) );
  NAND2_X1 U7129 ( .A1(n7763), .A2(n7765), .ZN(n5317) );
  INV_X1 U7130 ( .A(n7756), .ZN(n9678) );
  OR2_X1 U7131 ( .A1(n10260), .A2(n9678), .ZN(n5316) );
  NAND2_X1 U7132 ( .A1(n5317), .A2(n5316), .ZN(n7849) );
  INV_X1 U7133 ( .A(n5318), .ZN(n5320) );
  NAND2_X1 U7134 ( .A1(n5320), .A2(n5319), .ZN(n5324) );
  NAND2_X1 U7135 ( .A1(n5325), .A2(SI_6_), .ZN(n5326) );
  MUX2_X1 U7136 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n5035), .Z(n5367) );
  XNOR2_X1 U7137 ( .A(n5367), .B(SI_7_), .ZN(n5341) );
  XNOR2_X1 U7138 ( .A(n5365), .B(n5341), .ZN(n7161) );
  NAND2_X1 U7139 ( .A1(n7161), .A2(n5744), .ZN(n5329) );
  NAND2_X1 U7140 ( .A1(n5349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5327) );
  XNOR2_X1 U7141 ( .A(n5327), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7676) );
  AOI22_X1 U7142 ( .A1(n5593), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6443), .B2(
        n7676), .ZN(n5328) );
  NAND2_X1 U7143 ( .A1(n5788), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5339) );
  INV_X1 U7144 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6453) );
  OR2_X1 U7145 ( .A1(n5889), .A2(n6453), .ZN(n5338) );
  INV_X1 U7146 ( .A(n5333), .ZN(n5331) );
  INV_X1 U7147 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5332) );
  NAND2_X1 U7148 ( .A1(n5333), .A2(n5332), .ZN(n5334) );
  NAND2_X1 U7149 ( .A1(n5357), .A2(n5334), .ZN(n7866) );
  OR2_X1 U7150 ( .A1(n4290), .A2(n7866), .ZN(n5337) );
  INV_X1 U7151 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5335) );
  OR2_X1 U7152 ( .A1(n4291), .A2(n5335), .ZN(n5336) );
  OR2_X1 U7153 ( .A1(n7868), .A2(n8230), .ZN(n6039) );
  NAND2_X1 U7154 ( .A1(n7868), .A2(n8230), .ZN(n7934) );
  INV_X1 U7155 ( .A(n8230), .ZN(n9677) );
  OR2_X1 U7156 ( .A1(n7868), .A2(n9677), .ZN(n5340) );
  INV_X1 U7157 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U7158 ( .A1(n5365), .A2(n5342), .ZN(n5343) );
  NAND2_X1 U7159 ( .A1(n5367), .A2(SI_7_), .ZN(n5366) );
  NAND2_X1 U7160 ( .A1(n5343), .A2(n5366), .ZN(n5348) );
  MUX2_X1 U7161 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n5035), .Z(n5344) );
  INV_X1 U7162 ( .A(n5344), .ZN(n5346) );
  INV_X1 U7163 ( .A(SI_8_), .ZN(n5345) );
  NAND2_X1 U7164 ( .A1(n5346), .A2(n5345), .ZN(n5370) );
  NAND2_X1 U7165 ( .A1(n5368), .A2(n5370), .ZN(n5347) );
  NAND2_X1 U7166 ( .A1(n7163), .A2(n5744), .ZN(n5353) );
  INV_X1 U7167 ( .A(n5349), .ZN(n5351) );
  INV_X1 U7168 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U7169 ( .A1(n5351), .A2(n5350), .ZN(n5393) );
  NAND2_X1 U7170 ( .A1(n5393), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U7171 ( .A(n5378), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7665) );
  AOI22_X1 U7172 ( .A1(n5593), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6443), .B2(
        n7665), .ZN(n5352) );
  NAND2_X1 U7173 ( .A1(n5788), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5363) );
  INV_X1 U7174 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5354) );
  OR2_X1 U7175 ( .A1(n5889), .A2(n5354), .ZN(n5362) );
  INV_X1 U7176 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U7177 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  NAND2_X1 U7178 ( .A1(n5384), .A2(n5358), .ZN(n8233) );
  OR2_X1 U7179 ( .A1(n4290), .A2(n8233), .ZN(n5361) );
  INV_X1 U7180 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5359) );
  OR2_X1 U7181 ( .A1(n4291), .A2(n5359), .ZN(n5360) );
  OR2_X1 U7182 ( .A1(n8235), .A2(n8264), .ZN(n7973) );
  NAND2_X1 U7183 ( .A1(n8235), .A2(n8264), .ZN(n6040) );
  NAND2_X1 U7184 ( .A1(n7973), .A2(n6040), .ZN(n7933) );
  INV_X1 U7185 ( .A(n8264), .ZN(n9676) );
  OR2_X1 U7186 ( .A1(n8235), .A2(n9676), .ZN(n5364) );
  NOR2_X1 U7187 ( .A1(n5367), .A2(SI_7_), .ZN(n5369) );
  NAND2_X1 U7188 ( .A1(n5369), .A2(n5368), .ZN(n5371) );
  MUX2_X1 U7189 ( .A(n7194), .B(n7191), .S(n5035), .Z(n5374) );
  NAND2_X1 U7190 ( .A1(n5374), .A2(n5373), .ZN(n5391) );
  INV_X1 U7191 ( .A(n5374), .ZN(n5375) );
  NAND2_X1 U7192 ( .A1(n5375), .A2(SI_9_), .ZN(n5376) );
  XNOR2_X1 U7193 ( .A(n5390), .B(n5151), .ZN(n7189) );
  NAND2_X1 U7194 ( .A1(n7189), .A2(n5744), .ZN(n5382) );
  INV_X1 U7195 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U7196 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  NAND2_X1 U7197 ( .A1(n5379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U7198 ( .A(n5380), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7190) );
  AOI22_X1 U7199 ( .A1(n6443), .A2(n7190), .B1(n5593), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n5381) );
  NAND2_X2 U7200 ( .A1(n5382), .A2(n5381), .ZN(n8128) );
  NAND2_X1 U7201 ( .A1(n5306), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5389) );
  INV_X1 U7202 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6472) );
  OR2_X1 U7203 ( .A1(n4667), .A2(n6472), .ZN(n5388) );
  NAND2_X1 U7204 ( .A1(n5384), .A2(n5383), .ZN(n5385) );
  NAND2_X1 U7205 ( .A1(n5399), .A2(n5385), .ZN(n8265) );
  OR2_X1 U7206 ( .A1(n4290), .A2(n8265), .ZN(n5387) );
  INV_X1 U7207 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6454) );
  OR2_X1 U7208 ( .A1(n5889), .A2(n6454), .ZN(n5386) );
  OR2_X1 U7209 ( .A1(n8128), .A2(n7890), .ZN(n6057) );
  NAND2_X1 U7210 ( .A1(n8128), .A2(n7890), .ZN(n6041) );
  NAND2_X1 U7211 ( .A1(n6057), .A2(n6041), .ZN(n7984) );
  INV_X1 U7212 ( .A(n7890), .ZN(n9675) );
  MUX2_X1 U7213 ( .A(n7201), .B(n7204), .S(n5035), .Z(n5409) );
  XNOR2_X1 U7214 ( .A(n5409), .B(SI_10_), .ZN(n5408) );
  XNOR2_X1 U7215 ( .A(n5407), .B(n5408), .ZN(n7199) );
  NAND2_X1 U7216 ( .A1(n7199), .A2(n5744), .ZN(n5396) );
  NAND2_X1 U7217 ( .A1(n5418), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U7218 ( .A(n5394), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7202) );
  AOI22_X1 U7219 ( .A1(n4670), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n7202), .B2(
        n6443), .ZN(n5395) );
  NAND2_X1 U7220 ( .A1(n5788), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5404) );
  INV_X1 U7221 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5397) );
  OR2_X1 U7222 ( .A1(n4291), .A2(n5397), .ZN(n5403) );
  NAND2_X1 U7223 ( .A1(n5399), .A2(n5398), .ZN(n5400) );
  NAND2_X1 U7224 ( .A1(n5426), .A2(n5400), .ZN(n8323) );
  OR2_X1 U7225 ( .A1(n4290), .A2(n8323), .ZN(n5402) );
  INV_X1 U7226 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n8778) );
  OR2_X1 U7227 ( .A1(n5889), .A2(n8778), .ZN(n5401) );
  OR2_X1 U7228 ( .A1(n8325), .A2(n7993), .ZN(n6058) );
  NAND2_X1 U7229 ( .A1(n8325), .A2(n7993), .ZN(n6061) );
  INV_X1 U7230 ( .A(n7993), .ZN(n9674) );
  OR2_X1 U7231 ( .A1(n8325), .A2(n9674), .ZN(n5405) );
  INV_X1 U7232 ( .A(n5409), .ZN(n5410) );
  MUX2_X1 U7233 ( .A(n7233), .B(n7236), .S(n5035), .Z(n5412) );
  INV_X1 U7234 ( .A(n5412), .ZN(n5413) );
  NAND2_X1 U7235 ( .A1(n5413), .A2(SI_11_), .ZN(n5414) );
  NAND2_X1 U7236 ( .A1(n5433), .A2(n5414), .ZN(n5415) );
  NAND2_X1 U7237 ( .A1(n5416), .A2(n5415), .ZN(n5417) );
  INV_X1 U7238 ( .A(n5418), .ZN(n5420) );
  INV_X1 U7239 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U7240 ( .A1(n5420), .A2(n5419), .ZN(n5435) );
  NAND2_X1 U7241 ( .A1(n5435), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5421) );
  XNOR2_X1 U7242 ( .A(n5421), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7234) );
  AOI22_X1 U7243 ( .A1(n7234), .A2(n6443), .B1(n4670), .B2(
        P2_DATAO_REG_11__SCAN_IN), .ZN(n5422) );
  NAND2_X1 U7244 ( .A1(n5788), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5432) );
  INV_X1 U7245 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5424) );
  OR2_X1 U7246 ( .A1(n5889), .A2(n5424), .ZN(n5431) );
  INV_X1 U7247 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5425) );
  NAND2_X1 U7248 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  NAND2_X1 U7249 ( .A1(n5443), .A2(n5427), .ZN(n8365) );
  OR2_X1 U7250 ( .A1(n4290), .A2(n8365), .ZN(n5430) );
  INV_X1 U7251 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5428) );
  OR2_X1 U7252 ( .A1(n4291), .A2(n5428), .ZN(n5429) );
  NAND4_X1 U7253 ( .A1(n5432), .A2(n5431), .A3(n5430), .A4(n5429), .ZN(n9673)
         );
  AND2_X1 U7254 ( .A1(n8370), .A2(n9673), .ZN(n6060) );
  INV_X1 U7255 ( .A(n7989), .ZN(n7991) );
  MUX2_X1 U7256 ( .A(n7266), .B(n7264), .S(n6735), .Z(n5452) );
  XNOR2_X1 U7257 ( .A(n5456), .B(n5451), .ZN(n7262) );
  NAND2_X1 U7258 ( .A1(n7262), .A2(n5744), .ZN(n5440) );
  INV_X1 U7259 ( .A(n5435), .ZN(n5437) );
  INV_X1 U7260 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5436) );
  NAND2_X1 U7261 ( .A1(n5437), .A2(n5436), .ZN(n5438) );
  NAND2_X1 U7262 ( .A1(n5438), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5458) );
  XNOR2_X1 U7263 ( .A(n5458), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7263) );
  AOI22_X1 U7264 ( .A1(n7263), .A2(n6443), .B1(n4670), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U7265 ( .A1(n5306), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5448) );
  INV_X1 U7266 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8122) );
  OR2_X1 U7267 ( .A1(n4667), .A2(n8122), .ZN(n5447) );
  INV_X1 U7268 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n8712) );
  OR2_X1 U7269 ( .A1(n5889), .A2(n8712), .ZN(n5446) );
  INV_X1 U7270 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7271 ( .A1(n5443), .A2(n5442), .ZN(n5444) );
  NAND2_X1 U7272 ( .A1(n5463), .A2(n5444), .ZN(n9546) );
  OR2_X1 U7273 ( .A1(n4290), .A2(n9546), .ZN(n5445) );
  OR2_X1 U7274 ( .A1(n5450), .A2(n5449), .ZN(n8241) );
  INV_X1 U7275 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U7276 ( .A1(n5453), .A2(SI_12_), .ZN(n5454) );
  MUX2_X1 U7277 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n5035), .Z(n5476) );
  XNOR2_X1 U7278 ( .A(n5475), .B(n5473), .ZN(n7267) );
  NAND2_X1 U7279 ( .A1(n7267), .A2(n5744), .ZN(n5462) );
  INV_X1 U7280 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5457) );
  NAND2_X1 U7281 ( .A1(n5458), .A2(n5457), .ZN(n5459) );
  NAND2_X1 U7282 ( .A1(n5459), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5460) );
  XNOR2_X1 U7283 ( .A(n5460), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7268) );
  AOI22_X1 U7284 ( .A1(n7268), .A2(n6443), .B1(n4670), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5461) );
  INV_X1 U7285 ( .A(n5483), .ZN(n5485) );
  INV_X1 U7286 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U7287 ( .A1(n5463), .A2(n8748), .ZN(n5464) );
  AND2_X1 U7288 ( .A1(n5485), .A2(n5464), .ZN(n9612) );
  NAND2_X1 U7289 ( .A1(n9612), .A2(n5793), .ZN(n5468) );
  NAND2_X1 U7290 ( .A1(n5788), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U7291 ( .A1(n5306), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U7292 ( .A1(n5653), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n5465) );
  INV_X1 U7293 ( .A(n9961), .ZN(n9672) );
  OR2_X1 U7294 ( .A1(n5470), .A2(n9672), .ZN(n5469) );
  AND2_X1 U7295 ( .A1(n8241), .A2(n5469), .ZN(n5472) );
  INV_X1 U7296 ( .A(n5469), .ZN(n5471) );
  INV_X1 U7297 ( .A(n6066), .ZN(n5990) );
  NAND2_X1 U7298 ( .A1(n5470), .A2(n9961), .ZN(n9956) );
  NAND2_X1 U7299 ( .A1(n5476), .A2(SI_13_), .ZN(n5477) );
  MUX2_X1 U7300 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6735), .Z(n5496) );
  XNOR2_X1 U7301 ( .A(n5495), .B(n5493), .ZN(n6875) );
  NAND2_X1 U7302 ( .A1(n6875), .A2(n5744), .ZN(n5482) );
  OAI21_X1 U7303 ( .B1(n5479), .B2(n5478), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5480) );
  XNOR2_X1 U7304 ( .A(n5480), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U7305 ( .A1(n4670), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6443), .B2(
        n10153), .ZN(n5481) );
  INV_X1 U7306 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5489) );
  AOI22_X1 U7307 ( .A1(n5653), .A2(P1_REG1_REG_14__SCAN_IN), .B1(n5788), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n5488) );
  INV_X1 U7308 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7309 ( .A1(n5485), .A2(n5484), .ZN(n5486) );
  NAND2_X1 U7310 ( .A1(n5505), .A2(n5486), .ZN(n9970) );
  OR2_X1 U7311 ( .A1(n9970), .A2(n4290), .ZN(n5487) );
  OAI211_X1 U7312 ( .C1(n4291), .C2(n5489), .A(n5488), .B(n5487), .ZN(n9671)
         );
  INV_X1 U7313 ( .A(n9671), .ZN(n9655) );
  OR2_X1 U7314 ( .A1(n5832), .A2(n9655), .ZN(n5490) );
  NAND2_X1 U7315 ( .A1(n9954), .A2(n5490), .ZN(n5492) );
  NAND2_X1 U7316 ( .A1(n5832), .A2(n9655), .ZN(n5491) );
  NAND2_X1 U7317 ( .A1(n5496), .A2(SI_14_), .ZN(n5497) );
  MUX2_X1 U7318 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6735), .Z(n5514) );
  XNOR2_X1 U7319 ( .A(n5513), .B(n5511), .ZN(n7420) );
  NAND2_X1 U7320 ( .A1(n7420), .A2(n5744), .ZN(n5502) );
  INV_X1 U7321 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7322 ( .A1(n5499), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5500) );
  XNOR2_X1 U7323 ( .A(n5500), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10167) );
  AOI22_X1 U7324 ( .A1(n4670), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6443), .B2(
        n10167), .ZN(n5501) );
  INV_X1 U7325 ( .A(n5519), .ZN(n5521) );
  INV_X1 U7326 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5504) );
  NAND2_X1 U7327 ( .A1(n5505), .A2(n5504), .ZN(n5506) );
  AND2_X1 U7328 ( .A1(n5521), .A2(n5506), .ZN(n9657) );
  NAND2_X1 U7329 ( .A1(n9657), .A2(n5793), .ZN(n5509) );
  AOI22_X1 U7330 ( .A1(n5653), .A2(P1_REG1_REG_15__SCAN_IN), .B1(n5788), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n5508) );
  INV_X1 U7331 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n8701) );
  OR2_X1 U7332 ( .A1(n4291), .A2(n8701), .ZN(n5507) );
  NAND2_X1 U7333 ( .A1(n10051), .A2(n9933), .ZN(n5510) );
  MUX2_X1 U7334 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n6735), .Z(n5533) );
  XNOR2_X1 U7335 ( .A(n5532), .B(n5530), .ZN(n7517) );
  NAND2_X1 U7336 ( .A1(n7517), .A2(n5744), .ZN(n5518) );
  NAND2_X1 U7337 ( .A1(n5515), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5516) );
  XNOR2_X1 U7338 ( .A(n5516), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7518) );
  AOI22_X1 U7339 ( .A1(n4670), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6443), .B2(
        n7518), .ZN(n5517) );
  INV_X1 U7340 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5520) );
  NAND2_X1 U7341 ( .A1(n5521), .A2(n5520), .ZN(n5522) );
  NAND2_X1 U7342 ( .A1(n5548), .A2(n5522), .ZN(n9940) );
  OR2_X1 U7343 ( .A1(n9940), .A2(n4290), .ZN(n5527) );
  INV_X1 U7344 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10046) );
  NAND2_X1 U7345 ( .A1(n5306), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5524) );
  INV_X1 U7346 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9941) );
  OR2_X1 U7347 ( .A1(n4667), .A2(n9941), .ZN(n5523) );
  OAI211_X1 U7348 ( .C1(n10046), .C2(n5889), .A(n5524), .B(n5523), .ZN(n5525)
         );
  INV_X1 U7349 ( .A(n5525), .ZN(n5526) );
  NAND2_X1 U7350 ( .A1(n5527), .A2(n5526), .ZN(n9669) );
  AND2_X1 U7351 ( .A1(n10108), .A2(n9669), .ZN(n6075) );
  INV_X1 U7352 ( .A(n9946), .ZN(n5953) );
  NAND2_X1 U7353 ( .A1(n9945), .A2(n5953), .ZN(n5529) );
  OR2_X1 U7354 ( .A1(n10108), .A2(n9918), .ZN(n5528) );
  NAND2_X1 U7355 ( .A1(n5533), .A2(SI_16_), .ZN(n5534) );
  MUX2_X1 U7356 ( .A(n7597), .B(n5536), .S(n6735), .Z(n5538) );
  INV_X1 U7357 ( .A(n5538), .ZN(n5539) );
  NAND2_X1 U7358 ( .A1(n5539), .A2(SI_17_), .ZN(n5540) );
  NAND2_X1 U7359 ( .A1(n5557), .A2(n5540), .ZN(n5541) );
  NAND2_X1 U7360 ( .A1(n5542), .A2(n5541), .ZN(n5543) );
  NAND2_X1 U7361 ( .A1(n7566), .A2(n5744), .ZN(n5546) );
  XNOR2_X1 U7362 ( .A(n5561), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U7363 ( .A1(n4670), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6443), .B2(
        n10185), .ZN(n5545) );
  NAND2_X1 U7364 ( .A1(n5548), .A2(n5547), .ZN(n5549) );
  AND2_X1 U7365 ( .A1(n5567), .A2(n5549), .ZN(n9923) );
  NAND2_X1 U7366 ( .A1(n9923), .A2(n5793), .ZN(n5554) );
  INV_X1 U7367 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U7368 ( .A1(n5306), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5551) );
  INV_X1 U7369 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6464) );
  OR2_X1 U7370 ( .A1(n4667), .A2(n6464), .ZN(n5550) );
  OAI211_X1 U7371 ( .C1(n5889), .C2(n6458), .A(n5551), .B(n5550), .ZN(n5552)
         );
  INV_X1 U7372 ( .A(n5552), .ZN(n5553) );
  OR2_X1 U7373 ( .A1(n10039), .A2(n9935), .ZN(n5555) );
  NAND2_X1 U7374 ( .A1(n10039), .A2(n9935), .ZN(n5556) );
  MUX2_X1 U7375 ( .A(n5560), .B(n5559), .S(n6735), .Z(n5575) );
  XNOR2_X1 U7376 ( .A(n5575), .B(SI_18_), .ZN(n5574) );
  NAND2_X1 U7377 ( .A1(n6916), .A2(n5744), .ZN(n5564) );
  NAND2_X1 U7378 ( .A1(n5561), .A2(n5795), .ZN(n5589) );
  NAND2_X1 U7379 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5562) );
  XNOR2_X1 U7380 ( .A(n5562), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U7381 ( .A1(n4670), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n6443), .B2(
        n10200), .ZN(n5563) );
  INV_X1 U7382 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7383 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  NAND2_X1 U7384 ( .A1(n5615), .A2(n5568), .ZN(n9901) );
  OR2_X1 U7385 ( .A1(n9901), .A2(n4290), .ZN(n5573) );
  INV_X1 U7386 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n10035) );
  NAND2_X1 U7387 ( .A1(n5788), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7388 ( .A1(n5306), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5569) );
  OAI211_X1 U7389 ( .C1(n10035), .C2(n5889), .A(n5570), .B(n5569), .ZN(n5571)
         );
  INV_X1 U7390 ( .A(n5571), .ZN(n5572) );
  INV_X1 U7391 ( .A(n5574), .ZN(n5578) );
  INV_X1 U7392 ( .A(n5575), .ZN(n5576) );
  NAND2_X1 U7393 ( .A1(n5576), .A2(SI_18_), .ZN(n5577) );
  MUX2_X1 U7394 ( .A(n8785), .B(n8811), .S(n6735), .Z(n5580) );
  INV_X1 U7395 ( .A(SI_19_), .ZN(n5579) );
  NAND2_X1 U7396 ( .A1(n5580), .A2(n5579), .ZN(n5603) );
  INV_X1 U7397 ( .A(n5580), .ZN(n5581) );
  NAND2_X1 U7398 ( .A1(n5581), .A2(SI_19_), .ZN(n5582) );
  NAND2_X1 U7399 ( .A1(n5603), .A2(n5582), .ZN(n5604) );
  NAND2_X1 U7400 ( .A1(n7875), .A2(n5744), .ZN(n5595) );
  AND2_X1 U7401 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5583) );
  NAND2_X1 U7402 ( .A1(n5589), .A2(n5583), .ZN(n5588) );
  NAND2_X1 U7403 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5584) );
  NAND2_X1 U7404 ( .A1(n5584), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5585) );
  OAI21_X1 U7405 ( .B1(n5586), .B2(P1_IR_REG_31__SCAN_IN), .A(n5585), .ZN(
        n5587) );
  INV_X1 U7406 ( .A(n5589), .ZN(n5590) );
  AOI22_X1 U7407 ( .A1(n4670), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7856), .B2(
        n6443), .ZN(n5594) );
  XNOR2_X1 U7408 ( .A(n5615), .B(P1_REG3_REG_19__SCAN_IN), .ZN(n9887) );
  NAND2_X1 U7409 ( .A1(n9887), .A2(n5793), .ZN(n5601) );
  INV_X1 U7410 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5598) );
  NAND2_X1 U7411 ( .A1(n5306), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U7412 ( .A1(n5788), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5596) );
  OAI211_X1 U7413 ( .C1(n5598), .C2(n5889), .A(n5597), .B(n5596), .ZN(n5599)
         );
  INV_X1 U7414 ( .A(n5599), .ZN(n5600) );
  INV_X1 U7415 ( .A(n9898), .ZN(n9668) );
  AND2_X1 U7416 ( .A1(n10027), .A2(n9668), .ZN(n5602) );
  MUX2_X1 U7417 ( .A(n8098), .B(n8108), .S(n6735), .Z(n5606) );
  INV_X1 U7418 ( .A(SI_20_), .ZN(n5605) );
  NAND2_X1 U7419 ( .A1(n5606), .A2(n5605), .ZN(n5626) );
  INV_X1 U7420 ( .A(n5606), .ZN(n5607) );
  NAND2_X1 U7421 ( .A1(n5607), .A2(SI_20_), .ZN(n5608) );
  XNOR2_X1 U7422 ( .A(n5625), .B(n5624), .ZN(n8097) );
  NAND2_X1 U7423 ( .A1(n8097), .A2(n5744), .ZN(n5611) );
  OR2_X1 U7424 ( .A1(n5609), .A2(n8108), .ZN(n5610) );
  INV_X1 U7425 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5613) );
  INV_X1 U7426 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n5612) );
  OAI21_X1 U7427 ( .B1(n5615), .B2(n5613), .A(n5612), .ZN(n5616) );
  NAND2_X1 U7428 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5614) );
  NAND2_X1 U7429 ( .A1(n5616), .A2(n5631), .ZN(n9867) );
  OR2_X1 U7430 ( .A1(n9867), .A2(n4290), .ZN(n5621) );
  INV_X1 U7431 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10024) );
  NAND2_X1 U7432 ( .A1(n5306), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5618) );
  NAND2_X1 U7433 ( .A1(n5788), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5617) );
  OAI211_X1 U7434 ( .C1(n10024), .C2(n5889), .A(n5618), .B(n5617), .ZN(n5619)
         );
  INV_X1 U7435 ( .A(n5619), .ZN(n5620) );
  NOR2_X1 U7436 ( .A1(n10020), .A2(n9882), .ZN(n5623) );
  NAND2_X1 U7437 ( .A1(n10020), .A2(n9882), .ZN(n5622) );
  NAND2_X1 U7438 ( .A1(n5627), .A2(n5626), .ZN(n5640) );
  MUX2_X1 U7439 ( .A(n8214), .B(n8240), .S(n6735), .Z(n5643) );
  XNOR2_X1 U7440 ( .A(n5643), .B(SI_21_), .ZN(n5641) );
  XNOR2_X1 U7441 ( .A(n5640), .B(n5641), .ZN(n8213) );
  NAND2_X1 U7442 ( .A1(n8213), .A2(n5744), .ZN(n5629) );
  OR2_X1 U7443 ( .A1(n5609), .A2(n8240), .ZN(n5628) );
  INV_X1 U7444 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7445 ( .A1(n5631), .A2(n5630), .ZN(n5632) );
  NAND2_X1 U7446 ( .A1(n5651), .A2(n5632), .ZN(n9853) );
  OR2_X1 U7447 ( .A1(n9853), .A2(n4290), .ZN(n5637) );
  INV_X1 U7448 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U7449 ( .A1(n5788), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U7450 ( .A1(n5306), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5633) );
  OAI211_X1 U7451 ( .C1(n8758), .C2(n5889), .A(n5634), .B(n5633), .ZN(n5635)
         );
  INV_X1 U7452 ( .A(n5635), .ZN(n5636) );
  AND2_X1 U7453 ( .A1(n10014), .A2(n9836), .ZN(n5639) );
  OR2_X1 U7454 ( .A1(n10014), .A2(n9836), .ZN(n5638) );
  INV_X1 U7455 ( .A(n5643), .ZN(n5644) );
  NAND2_X1 U7456 ( .A1(n5644), .A2(SI_21_), .ZN(n5645) );
  MUX2_X1 U7457 ( .A(n8289), .B(n8287), .S(n6735), .Z(n5646) );
  NAND2_X1 U7458 ( .A1(n5646), .A2(n8710), .ZN(n5661) );
  INV_X1 U7459 ( .A(n5646), .ZN(n5647) );
  NAND2_X1 U7460 ( .A1(n5647), .A2(SI_22_), .ZN(n5648) );
  NAND2_X1 U7461 ( .A1(n5661), .A2(n5648), .ZN(n5662) );
  XNOR2_X1 U7462 ( .A(n5663), .B(n5662), .ZN(n8286) );
  NAND2_X1 U7463 ( .A1(n8286), .A2(n5744), .ZN(n5650) );
  OR2_X1 U7464 ( .A1(n5609), .A2(n8287), .ZN(n5649) );
  INV_X1 U7465 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9624) );
  NAND2_X1 U7466 ( .A1(n5651), .A2(n9624), .ZN(n5652) );
  NAND2_X1 U7467 ( .A1(n5674), .A2(n5652), .ZN(n9840) );
  OR2_X1 U7468 ( .A1(n9840), .A2(n4290), .ZN(n5659) );
  INV_X1 U7469 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U7470 ( .A1(n5306), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U7471 ( .A1(n5653), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n5654) );
  OAI211_X1 U7472 ( .C1(n4667), .C2(n5656), .A(n5655), .B(n5654), .ZN(n5657)
         );
  INV_X1 U7473 ( .A(n5657), .ZN(n5658) );
  NAND2_X1 U7474 ( .A1(n10009), .A2(n9860), .ZN(n5660) );
  MUX2_X1 U7475 ( .A(n8722), .B(n8306), .S(n6735), .Z(n5665) );
  INV_X1 U7476 ( .A(SI_23_), .ZN(n5664) );
  NAND2_X1 U7477 ( .A1(n5665), .A2(n5664), .ZN(n5682) );
  INV_X1 U7478 ( .A(n5665), .ZN(n5666) );
  NAND2_X1 U7479 ( .A1(n5666), .A2(SI_23_), .ZN(n5667) );
  OR2_X1 U7480 ( .A1(n5669), .A2(n5668), .ZN(n5670) );
  NAND2_X1 U7481 ( .A1(n5683), .A2(n5670), .ZN(n8307) );
  NAND2_X1 U7482 ( .A1(n8307), .A2(n5744), .ZN(n5672) );
  OR2_X1 U7483 ( .A1(n5609), .A2(n8306), .ZN(n5671) );
  INV_X1 U7484 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5673) );
  NAND2_X1 U7485 ( .A1(n5674), .A2(n5673), .ZN(n5675) );
  AND2_X1 U7486 ( .A1(n5691), .A2(n5675), .ZN(n9828) );
  NAND2_X1 U7487 ( .A1(n9828), .A2(n5793), .ZN(n5680) );
  INV_X1 U7488 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U7489 ( .A1(n5788), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U7490 ( .A1(n5306), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5676) );
  OAI211_X1 U7491 ( .C1(n10006), .C2(n5889), .A(n5677), .B(n5676), .ZN(n5678)
         );
  INV_X1 U7492 ( .A(n5678), .ZN(n5679) );
  OR2_X1 U7493 ( .A1(n9825), .A2(n9835), .ZN(n5681) );
  MUX2_X1 U7494 ( .A(n8382), .B(n8589), .S(n6735), .Z(n5685) );
  INV_X1 U7495 ( .A(SI_24_), .ZN(n5684) );
  NAND2_X1 U7496 ( .A1(n5685), .A2(n5684), .ZN(n5717) );
  INV_X1 U7497 ( .A(n5685), .ZN(n5686) );
  NAND2_X1 U7498 ( .A1(n5686), .A2(SI_24_), .ZN(n5687) );
  XNOR2_X1 U7499 ( .A(n5701), .B(n5700), .ZN(n6973) );
  NAND2_X1 U7500 ( .A1(n6973), .A2(n5744), .ZN(n5689) );
  OR2_X1 U7501 ( .A1(n5609), .A2(n8589), .ZN(n5688) );
  INV_X1 U7502 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7503 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  NAND2_X1 U7504 ( .A1(n5708), .A2(n5692), .ZN(n9590) );
  OR2_X1 U7505 ( .A1(n9590), .A2(n4290), .ZN(n5697) );
  INV_X1 U7506 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n10001) );
  NAND2_X1 U7507 ( .A1(n5788), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5694) );
  NAND2_X1 U7508 ( .A1(n5306), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U7509 ( .C1(n5889), .C2(n10001), .A(n5694), .B(n5693), .ZN(n5695)
         );
  INV_X1 U7510 ( .A(n5695), .ZN(n5696) );
  AND2_X1 U7511 ( .A1(n5839), .A2(n9667), .ZN(n5699) );
  NAND2_X1 U7512 ( .A1(n5701), .A2(n5700), .ZN(n5720) );
  MUX2_X1 U7513 ( .A(n9495), .B(n10132), .S(n6735), .Z(n5703) );
  INV_X1 U7514 ( .A(SI_25_), .ZN(n5702) );
  NAND2_X1 U7515 ( .A1(n5703), .A2(n5702), .ZN(n5737) );
  INV_X1 U7516 ( .A(n5703), .ZN(n5704) );
  NAND2_X1 U7517 ( .A1(n5704), .A2(SI_25_), .ZN(n5718) );
  NAND2_X1 U7518 ( .A1(n9493), .A2(n5744), .ZN(n5706) );
  OR2_X1 U7519 ( .A1(n5609), .A2(n10132), .ZN(n5705) );
  INV_X1 U7520 ( .A(n5708), .ZN(n5707) );
  INV_X1 U7521 ( .A(n5725), .ZN(n5727) );
  INV_X1 U7522 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9556) );
  NAND2_X1 U7523 ( .A1(n5708), .A2(n9556), .ZN(n5709) );
  NAND2_X1 U7524 ( .A1(n5727), .A2(n5709), .ZN(n9788) );
  OR2_X1 U7525 ( .A1(n9788), .A2(n4290), .ZN(n5714) );
  INV_X1 U7526 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U7527 ( .A1(n5788), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5711) );
  NAND2_X1 U7528 ( .A1(n5306), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5710) );
  OAI211_X1 U7529 ( .C1(n5889), .C2(n9997), .A(n5711), .B(n5710), .ZN(n5712)
         );
  INV_X1 U7530 ( .A(n5712), .ZN(n5713) );
  AND2_X1 U7531 ( .A1(n5717), .A2(n5737), .ZN(n5719) );
  INV_X1 U7532 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9491) );
  INV_X1 U7533 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n10129) );
  MUX2_X1 U7534 ( .A(n9491), .B(n10129), .S(n6735), .Z(n5722) );
  INV_X1 U7535 ( .A(SI_26_), .ZN(n5721) );
  NAND2_X1 U7536 ( .A1(n5722), .A2(n5721), .ZN(n5736) );
  INV_X1 U7537 ( .A(n5722), .ZN(n5723) );
  NAND2_X1 U7538 ( .A1(n5723), .A2(SI_26_), .ZN(n5760) );
  OR2_X1 U7539 ( .A1(n5609), .A2(n10129), .ZN(n5724) );
  INV_X1 U7540 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5726) );
  NAND2_X1 U7541 ( .A1(n5727), .A2(n5726), .ZN(n5728) );
  NAND2_X1 U7542 ( .A1(n9774), .A2(n5793), .ZN(n5733) );
  INV_X1 U7543 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U7544 ( .A1(n5788), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5730) );
  NAND2_X1 U7545 ( .A1(n5306), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5729) );
  OAI211_X1 U7546 ( .C1(n9993), .C2(n5889), .A(n5730), .B(n5729), .ZN(n5731)
         );
  INV_X1 U7547 ( .A(n5731), .ZN(n5732) );
  NAND2_X1 U7548 ( .A1(n9780), .A2(n9795), .ZN(n6117) );
  INV_X1 U7549 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8385) );
  MUX2_X1 U7550 ( .A(n9486), .B(n8385), .S(n6735), .Z(n5740) );
  INV_X1 U7551 ( .A(SI_27_), .ZN(n5739) );
  NAND2_X1 U7552 ( .A1(n5740), .A2(n5739), .ZN(n5773) );
  INV_X1 U7553 ( .A(n5740), .ZN(n5741) );
  NAND2_X1 U7554 ( .A1(n5741), .A2(SI_27_), .ZN(n5742) );
  NAND2_X1 U7555 ( .A1(n5773), .A2(n5742), .ZN(n5758) );
  NAND2_X1 U7556 ( .A1(n8383), .A2(n5744), .ZN(n5746) );
  OR2_X1 U7557 ( .A1(n5609), .A2(n8385), .ZN(n5745) );
  INV_X1 U7558 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U7559 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7560 ( .A1(n5765), .A2(n5750), .ZN(n9761) );
  INV_X1 U7561 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5754) );
  NAND2_X1 U7562 ( .A1(n5788), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5753) );
  NAND2_X1 U7563 ( .A1(n5306), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5752) );
  OAI211_X1 U7564 ( .C1(n5754), .C2(n5889), .A(n5753), .B(n5752), .ZN(n5755)
         );
  INV_X1 U7565 ( .A(n5755), .ZN(n5756) );
  NAND2_X1 U7566 ( .A1(n9987), .A2(n9778), .ZN(n5915) );
  INV_X1 U7567 ( .A(n5758), .ZN(n5759) );
  INV_X1 U7568 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9485) );
  INV_X1 U7569 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10127) );
  MUX2_X1 U7570 ( .A(n9485), .B(n10127), .S(n6735), .Z(n5777) );
  XNOR2_X1 U7571 ( .A(n5777), .B(SI_28_), .ZN(n5893) );
  NAND2_X1 U7572 ( .A1(n7021), .A2(n5744), .ZN(n5764) );
  OR2_X1 U7573 ( .A1(n5609), .A2(n10127), .ZN(n5763) );
  INV_X1 U7574 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U7575 ( .A1(n5765), .A2(n6432), .ZN(n5766) );
  INV_X1 U7576 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n7139) );
  NAND2_X1 U7577 ( .A1(n5788), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7578 ( .A1(n5306), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5767) );
  OAI211_X1 U7579 ( .C1(n7139), .C2(n5889), .A(n5768), .B(n5767), .ZN(n5769)
         );
  NAND2_X1 U7580 ( .A1(n7140), .A2(n9766), .ZN(n5916) );
  NAND2_X1 U7581 ( .A1(n6129), .A2(n5916), .ZN(n7127) );
  INV_X1 U7582 ( .A(n5777), .ZN(n5774) );
  NAND2_X1 U7583 ( .A1(n5774), .A2(SI_28_), .ZN(n5770) );
  MUX2_X1 U7584 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n6735), .Z(n5896) );
  INV_X1 U7585 ( .A(n5896), .ZN(n5776) );
  NAND2_X1 U7586 ( .A1(n5770), .A2(n5776), .ZN(n5772) );
  INV_X1 U7587 ( .A(SI_28_), .ZN(n5775) );
  NAND2_X1 U7588 ( .A1(n5777), .A2(n5775), .ZN(n5895) );
  INV_X1 U7589 ( .A(n5772), .ZN(n5781) );
  INV_X1 U7590 ( .A(n5773), .ZN(n5780) );
  OAI21_X1 U7591 ( .B1(n5776), .B2(n5775), .A(n5774), .ZN(n5779) );
  OAI21_X1 U7592 ( .B1(n5896), .B2(SI_28_), .A(n5777), .ZN(n5778) );
  AOI22_X1 U7593 ( .A1(n5781), .A2(n5780), .B1(n5779), .B2(n5778), .ZN(n5782)
         );
  XNOR2_X1 U7594 ( .A(n5900), .B(SI_29_), .ZN(n8386) );
  NAND2_X1 U7595 ( .A1(n8386), .A2(n5744), .ZN(n5786) );
  INV_X1 U7596 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8387) );
  OR2_X1 U7597 ( .A1(n5609), .A2(n8387), .ZN(n5785) );
  INV_X1 U7598 ( .A(n5787), .ZN(n9744) );
  INV_X1 U7599 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7600 ( .A1(n5306), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7601 ( .A1(n5788), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5789) );
  OAI211_X1 U7602 ( .C1(n5791), .C2(n5889), .A(n5790), .B(n5789), .ZN(n5792)
         );
  AOI21_X1 U7603 ( .B1(n9744), .B2(n5793), .A(n5792), .ZN(n7729) );
  NOR2_X1 U7604 ( .A1(n5817), .A2(n7729), .ZN(n6134) );
  INV_X1 U7605 ( .A(n6134), .ZN(n5924) );
  INV_X1 U7606 ( .A(n6133), .ZN(n5908) );
  NAND2_X1 U7607 ( .A1(n5801), .A2(n5798), .ZN(n5859) );
  NAND2_X1 U7608 ( .A1(n5803), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5804) );
  NAND2_X1 U7609 ( .A1(n6444), .A2(n6164), .ZN(n7718) );
  INV_X1 U7610 ( .A(n6165), .ZN(n5807) );
  NAND2_X1 U7611 ( .A1(n5807), .A2(n9871), .ZN(n6161) );
  NAND2_X1 U7612 ( .A1(n6161), .A2(n5884), .ZN(n5808) );
  INV_X1 U7613 ( .A(n6394), .ZN(n7717) );
  NAND2_X1 U7614 ( .A1(n7718), .A2(n5809), .ZN(n10278) );
  NAND2_X4 U7615 ( .A1(n4590), .A2(n7856), .ZN(n6151) );
  INV_X1 U7616 ( .A(n9766), .ZN(n9665) );
  NAND2_X1 U7617 ( .A1(n7140), .A2(n9665), .ZN(n9738) );
  NAND4_X1 U7618 ( .A1(n9739), .A2(n9740), .A3(n10250), .A4(n9738), .ZN(n5852)
         );
  INV_X1 U7619 ( .A(n5817), .ZN(n9747) );
  NAND2_X1 U7620 ( .A1(n7711), .A2(n7757), .ZN(n7768) );
  INV_X1 U7621 ( .A(n8235), .ZN(n10275) );
  NOR2_X2 U7622 ( .A1(n7977), .A2(n8128), .ZN(n7891) );
  INV_X1 U7623 ( .A(n10039), .ZN(n9926) );
  NOR2_X2 U7624 ( .A1(n9919), .A2(n10031), .ZN(n9907) );
  NAND2_X1 U7625 ( .A1(n9890), .A2(n9907), .ZN(n9886) );
  NAND2_X1 U7626 ( .A1(n9747), .A2(n5813), .ZN(n9732) );
  AND2_X1 U7627 ( .A1(n6394), .A2(n8110), .ZN(n10015) );
  AOI21_X1 U7628 ( .B1(n5817), .B2(n7135), .A(n9952), .ZN(n5814) );
  AND2_X1 U7629 ( .A1(n9732), .A2(n5814), .ZN(n9743) );
  INV_X1 U7630 ( .A(n9738), .ZN(n5815) );
  INV_X1 U7631 ( .A(n5818), .ZN(n6025) );
  NOR2_X2 U7632 ( .A1(n7401), .A2(n7405), .ZN(n7400) );
  NAND2_X1 U7633 ( .A1(n7708), .A2(n7577), .ZN(n5975) );
  NAND2_X1 U7634 ( .A1(n5820), .A2(n6036), .ZN(n7764) );
  INV_X1 U7635 ( .A(n6041), .ZN(n6051) );
  NAND2_X1 U7636 ( .A1(n6040), .A2(n7934), .ZN(n6048) );
  OR2_X1 U7637 ( .A1(n6051), .A2(n6048), .ZN(n5941) );
  NOR2_X1 U7638 ( .A1(n5941), .A2(n7846), .ZN(n5821) );
  NAND2_X1 U7639 ( .A1(n5824), .A2(n6041), .ZN(n5822) );
  NAND2_X1 U7640 ( .A1(n5822), .A2(n5941), .ZN(n5982) );
  NAND2_X1 U7641 ( .A1(n7845), .A2(n6039), .ZN(n5823) );
  INV_X1 U7642 ( .A(n5980), .ZN(n5825) );
  NAND2_X1 U7643 ( .A1(n5829), .A2(n8116), .ZN(n6053) );
  INV_X1 U7644 ( .A(n6053), .ZN(n5985) );
  OR2_X1 U7645 ( .A1(n6063), .A2(n5985), .ZN(n8244) );
  AND2_X1 U7646 ( .A1(n5830), .A2(n8244), .ZN(n5831) );
  AND2_X1 U7647 ( .A1(n5832), .A2(n9671), .ZN(n6067) );
  NAND2_X1 U7648 ( .A1(n10055), .A2(n9655), .ZN(n6068) );
  NAND2_X1 U7649 ( .A1(n10051), .A2(n9963), .ZN(n6078) );
  NAND2_X1 U7650 ( .A1(n6073), .A2(n6078), .ZN(n8375) );
  XNOR2_X1 U7651 ( .A(n10039), .B(n9899), .ZN(n9913) );
  OR2_X1 U7652 ( .A1(n10039), .A2(n9899), .ZN(n5967) );
  OR2_X1 U7653 ( .A1(n10027), .A2(n9898), .ZN(n6093) );
  NAND2_X1 U7654 ( .A1(n10027), .A2(n9898), .ZN(n6098) );
  NAND2_X1 U7655 ( .A1(n10020), .A2(n9527), .ZN(n6097) );
  OR2_X1 U7656 ( .A1(n10020), .A2(n9527), .ZN(n6092) );
  XNOR2_X1 U7657 ( .A(n10014), .B(n9836), .ZN(n9858) );
  OR2_X1 U7658 ( .A1(n10014), .A2(n9869), .ZN(n6103) );
  INV_X1 U7659 ( .A(n6097), .ZN(n5837) );
  NAND2_X1 U7660 ( .A1(n6103), .A2(n5837), .ZN(n5838) );
  NAND2_X1 U7661 ( .A1(n10014), .A2(n9869), .ZN(n6108) );
  AND2_X1 U7662 ( .A1(n5838), .A2(n6108), .ZN(n5918) );
  NAND2_X1 U7663 ( .A1(n10009), .A2(n9824), .ZN(n5917) );
  OR2_X1 U7664 ( .A1(n9825), .A2(n9625), .ZN(n5910) );
  NAND2_X1 U7665 ( .A1(n9825), .A2(n9625), .ZN(n6111) );
  OR2_X1 U7666 ( .A1(n5839), .A2(n9823), .ZN(n6020) );
  NAND2_X1 U7667 ( .A1(n5839), .A2(n9823), .ZN(n6018) );
  NAND2_X1 U7668 ( .A1(n6020), .A2(n6018), .ZN(n9804) );
  INV_X1 U7669 ( .A(n6111), .ZN(n9805) );
  NOR2_X1 U7670 ( .A1(n9804), .A2(n9805), .ZN(n5840) );
  NAND2_X1 U7671 ( .A1(n9790), .A2(n9810), .ZN(n9775) );
  NAND2_X1 U7672 ( .A1(n6116), .A2(n9775), .ZN(n9792) );
  NAND2_X1 U7673 ( .A1(n6117), .A2(n9775), .ZN(n6112) );
  INV_X1 U7674 ( .A(n5916), .ZN(n5841) );
  XNOR2_X1 U7675 ( .A(n5842), .B(n9740), .ZN(n5851) );
  OR2_X1 U7676 ( .A1(n4590), .A2(n9871), .ZN(n5844) );
  NAND2_X1 U7677 ( .A1(n4294), .A2(n6393), .ZN(n5843) );
  INV_X1 U7678 ( .A(n6444), .ZN(n5845) );
  NOR2_X2 U7679 ( .A1(n5845), .A2(n4675), .ZN(n9932) );
  AND2_X1 U7680 ( .A1(n5846), .A2(P1_B_REG_SCAN_IN), .ZN(n5847) );
  NOR2_X1 U7681 ( .A1(n9962), .A2(n5847), .ZN(n9725) );
  INV_X1 U7682 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9982) );
  NAND2_X1 U7683 ( .A1(n5788), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5849) );
  NAND2_X1 U7684 ( .A1(n5306), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5848) );
  OAI211_X1 U7685 ( .C1(n5889), .C2(n9982), .A(n5849), .B(n5848), .ZN(n9664)
         );
  NAND2_X1 U7686 ( .A1(n5863), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5855) );
  NAND2_X1 U7687 ( .A1(n10135), .A2(P1_B_REG_SCAN_IN), .ZN(n5862) );
  INV_X1 U7688 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7689 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  OAI21_X2 U7690 ( .B1(n5859), .B2(n5858), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5861) );
  MUX2_X1 U7691 ( .A(P1_B_REG_SCAN_IN), .B(n5862), .S(n5881), .Z(n5867) );
  NAND2_X1 U7692 ( .A1(n4361), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5865) );
  INV_X1 U7693 ( .A(n10131), .ZN(n5866) );
  NAND2_X1 U7694 ( .A1(n10131), .A2(n10135), .ZN(n10115) );
  NAND2_X1 U7695 ( .A1(n10015), .A2(n7856), .ZN(n6397) );
  NOR2_X1 U7696 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n5872) );
  NOR4_X1 U7697 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5871) );
  NOR4_X1 U7698 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5870) );
  NOR4_X1 U7699 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5869) );
  NAND4_X1 U7700 ( .A1(n5872), .A2(n5871), .A3(n5870), .A4(n5869), .ZN(n5878)
         );
  NOR4_X1 U7701 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5876) );
  NOR4_X1 U7702 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5875) );
  NOR4_X1 U7703 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5874) );
  NOR4_X1 U7704 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5873) );
  NAND4_X1 U7705 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n5877)
         );
  NOR2_X1 U7706 ( .A1(n5878), .A2(n5877), .ZN(n5879) );
  OR2_X4 U7707 ( .A1(n5881), .A2(n5880), .ZN(n7143) );
  NAND2_X1 U7708 ( .A1(n5882), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5883) );
  AND3_X1 U7709 ( .A1(n7143), .A2(P1_STATE_REG_SCAN_IN), .A3(n7144), .ZN(
        n10113) );
  NAND2_X1 U7710 ( .A1(n6444), .A2(n5884), .ZN(n6401) );
  NAND2_X1 U7711 ( .A1(n5881), .A2(n10131), .ZN(n10116) );
  NAND2_X1 U7712 ( .A1(n10282), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5887) );
  INV_X1 U7713 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9978) );
  OR2_X1 U7714 ( .A1(n5889), .A2(n9978), .ZN(n5892) );
  INV_X1 U7715 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9728) );
  OR2_X1 U7716 ( .A1(n4667), .A2(n9728), .ZN(n5891) );
  INV_X1 U7717 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10069) );
  OR2_X1 U7718 ( .A1(n4291), .A2(n10069), .ZN(n5890) );
  INV_X1 U7719 ( .A(n5965), .ZN(n9724) );
  NAND2_X1 U7720 ( .A1(n9664), .A2(n9724), .ZN(n6138) );
  INV_X1 U7721 ( .A(SI_29_), .ZN(n5899) );
  NAND2_X1 U7722 ( .A1(n5894), .A2(n5893), .ZN(n5897) );
  NAND3_X1 U7723 ( .A1(n5897), .A2(n5896), .A3(n5895), .ZN(n5898) );
  INV_X1 U7724 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8634) );
  INV_X1 U7725 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8822) );
  MUX2_X1 U7726 ( .A(n8634), .B(n8822), .S(n4893), .Z(n5902) );
  INV_X1 U7727 ( .A(SI_30_), .ZN(n5901) );
  NAND2_X1 U7728 ( .A1(n5902), .A2(n5901), .ZN(n5931) );
  INV_X1 U7729 ( .A(n5902), .ZN(n5903) );
  NAND2_X1 U7730 ( .A1(n5903), .A2(SI_30_), .ZN(n5904) );
  NAND2_X1 U7731 ( .A1(n5931), .A2(n5904), .ZN(n5932) );
  NAND2_X1 U7732 ( .A1(n8632), .A2(n5744), .ZN(n5906) );
  OR2_X1 U7733 ( .A1(n5609), .A2(n8634), .ZN(n5905) );
  INV_X1 U7734 ( .A(n9664), .ZN(n5907) );
  NAND2_X1 U7735 ( .A1(n9733), .A2(n5907), .ZN(n5958) );
  NAND2_X1 U7736 ( .A1(n5958), .A2(n5908), .ZN(n6005) );
  INV_X1 U7737 ( .A(n6005), .ZN(n5929) );
  NAND2_X1 U7738 ( .A1(n6121), .A2(n6115), .ZN(n5966) );
  OR2_X1 U7739 ( .A1(n10009), .A2(n9824), .ZN(n5909) );
  NAND2_X1 U7740 ( .A1(n5910), .A2(n5909), .ZN(n6104) );
  NAND2_X1 U7741 ( .A1(n6104), .A2(n6111), .ZN(n5911) );
  NAND2_X1 U7742 ( .A1(n6020), .A2(n5911), .ZN(n5912) );
  NAND2_X1 U7743 ( .A1(n5912), .A2(n6018), .ZN(n5920) );
  AND2_X1 U7744 ( .A1(n6103), .A2(n6092), .ZN(n6099) );
  NAND3_X1 U7745 ( .A1(n6116), .A2(n5920), .A3(n6099), .ZN(n5997) );
  INV_X1 U7746 ( .A(n5913), .ZN(n5914) );
  NOR2_X1 U7747 ( .A1(n5966), .A2(n5914), .ZN(n5927) );
  AND2_X1 U7748 ( .A1(n6111), .A2(n5917), .ZN(n6107) );
  NAND3_X1 U7749 ( .A1(n6018), .A2(n6107), .A3(n5918), .ZN(n5919) );
  NAND3_X1 U7750 ( .A1(n6116), .A2(n5920), .A3(n5919), .ZN(n5921) );
  AND2_X1 U7751 ( .A1(n5921), .A2(n9775), .ZN(n5922) );
  NOR2_X1 U7752 ( .A1(n5966), .A2(n5922), .ZN(n5923) );
  INV_X1 U7753 ( .A(n6003), .ZN(n5926) );
  NAND2_X1 U7754 ( .A1(n5924), .A2(n6129), .ZN(n6001) );
  INV_X1 U7755 ( .A(n6001), .ZN(n5925) );
  OAI21_X1 U7756 ( .B1(n5927), .B2(n5926), .A(n5925), .ZN(n5928) );
  OAI211_X1 U7757 ( .C1(n10075), .C2(n9724), .A(n5929), .B(n5928), .ZN(n5930)
         );
  OAI21_X1 U7758 ( .B1(n6138), .B2(n9733), .A(n5930), .ZN(n5940) );
  MUX2_X1 U7759 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4893), .Z(n5935) );
  INV_X1 U7760 ( .A(SI_31_), .ZN(n5934) );
  XNOR2_X1 U7761 ( .A(n5935), .B(n5934), .ZN(n5936) );
  NAND2_X1 U7762 ( .A1(n10123), .A2(n5744), .ZN(n5939) );
  INV_X1 U7763 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10119) );
  OR2_X1 U7764 ( .A1(n5609), .A2(n10119), .ZN(n5938) );
  OR2_X1 U7765 ( .A1(n9723), .A2(n5965), .ZN(n6153) );
  NAND2_X1 U7766 ( .A1(n5940), .A2(n6153), .ZN(n5964) );
  INV_X1 U7767 ( .A(n9804), .ZN(n9802) );
  INV_X1 U7768 ( .A(n9881), .ZN(n9877) );
  INV_X1 U7769 ( .A(n5941), .ZN(n5947) );
  INV_X1 U7770 ( .A(n7400), .ZN(n5942) );
  NAND2_X1 U7771 ( .A1(n7401), .A2(n7405), .ZN(n5971) );
  NAND2_X1 U7772 ( .A1(n5942), .A2(n5971), .ZN(n7719) );
  INV_X1 U7773 ( .A(n7719), .ZN(n5944) );
  NAND4_X1 U7774 ( .A1(n7391), .A2(n5944), .A3(n8238), .A4(n5943), .ZN(n5945)
         );
  NAND2_X1 U7775 ( .A1(n6033), .A2(n5975), .ZN(n7704) );
  INV_X1 U7776 ( .A(n7683), .ZN(n7688) );
  NOR3_X1 U7777 ( .A1(n5945), .A2(n7704), .A3(n7688), .ZN(n5946) );
  NAND4_X1 U7778 ( .A1(n5947), .A2(n7610), .A3(n5946), .A4(n5315), .ZN(n5948)
         );
  NOR2_X1 U7779 ( .A1(n5948), .A2(n7888), .ZN(n5949) );
  NAND4_X1 U7780 ( .A1(n5980), .A2(n8118), .A3(n7989), .A4(n5949), .ZN(n5950)
         );
  NOR2_X1 U7781 ( .A1(n8247), .A2(n5950), .ZN(n5951) );
  NAND3_X1 U7782 ( .A1(n5834), .A2(n9958), .A3(n5951), .ZN(n5952) );
  OR4_X1 U7783 ( .A1(n9904), .A2(n9913), .A3(n5953), .A4(n5952), .ZN(n5954) );
  NOR2_X1 U7784 ( .A1(n9877), .A2(n5954), .ZN(n5955) );
  XNOR2_X1 U7785 ( .A(n10020), .B(n9882), .ZN(n9873) );
  AND4_X1 U7786 ( .A1(n9819), .A2(n5955), .A3(n9858), .A4(n9873), .ZN(n5956)
         );
  NAND3_X1 U7787 ( .A1(n9802), .A2(n5956), .A3(n9846), .ZN(n5957) );
  AOI22_X1 U7788 ( .A1(n5964), .A2(n6444), .B1(n6146), .B2(n6004), .ZN(n6016)
         );
  NAND2_X1 U7789 ( .A1(n9723), .A2(n5965), .ZN(n6152) );
  NAND4_X1 U7790 ( .A1(n6152), .A2(n6442), .A3(n6393), .A4(n9871), .ZN(n6015)
         );
  INV_X1 U7791 ( .A(n5966), .ZN(n6000) );
  NAND2_X1 U7792 ( .A1(n5968), .A2(n5967), .ZN(n6091) );
  NAND2_X1 U7793 ( .A1(n6078), .A2(n6068), .ZN(n6085) );
  NAND2_X1 U7794 ( .A1(n4643), .A2(n5969), .ZN(n5970) );
  NAND4_X1 U7795 ( .A1(n6027), .A2(n5971), .A3(n4294), .A4(n5970), .ZN(n5972)
         );
  NAND3_X1 U7796 ( .A1(n5973), .A2(n7698), .A3(n5972), .ZN(n5976) );
  AND2_X1 U7797 ( .A1(n5974), .A2(n6033), .ZN(n6028) );
  NAND2_X1 U7798 ( .A1(n6037), .A2(n5975), .ZN(n6044) );
  AOI21_X1 U7799 ( .B1(n5976), .B2(n6028), .A(n6044), .ZN(n5978) );
  INV_X1 U7800 ( .A(n6036), .ZN(n5977) );
  OAI21_X1 U7801 ( .B1(n5978), .B2(n5977), .A(n5315), .ZN(n5979) );
  NAND2_X1 U7802 ( .A1(n5980), .A2(n5979), .ZN(n5983) );
  INV_X1 U7803 ( .A(n6058), .ZN(n5981) );
  AOI21_X1 U7804 ( .B1(n5983), .B2(n5982), .A(n5981), .ZN(n5987) );
  AND2_X1 U7805 ( .A1(n5984), .A2(n6061), .ZN(n6054) );
  INV_X1 U7806 ( .A(n6054), .ZN(n5986) );
  OAI21_X1 U7807 ( .B1(n5987), .B2(n5986), .A(n5985), .ZN(n5988) );
  NAND3_X1 U7808 ( .A1(n5988), .A2(n9956), .A3(n6056), .ZN(n5989) );
  AND3_X1 U7809 ( .A1(n5990), .A2(n6069), .A3(n5989), .ZN(n5991) );
  OAI211_X1 U7810 ( .C1(n6085), .C2(n5991), .A(n6082), .B(n6073), .ZN(n5992)
         );
  AND2_X1 U7811 ( .A1(n5992), .A2(n6081), .ZN(n5994) );
  NAND2_X1 U7812 ( .A1(n10039), .A2(n9899), .ZN(n5993) );
  OAI21_X1 U7813 ( .B1(n6091), .B2(n5994), .A(n4338), .ZN(n5995) );
  AOI21_X1 U7814 ( .B1(n4384), .B2(n5995), .A(n4780), .ZN(n5996) );
  NOR2_X1 U7815 ( .A1(n5997), .A2(n5996), .ZN(n5999) );
  INV_X1 U7816 ( .A(n6117), .ZN(n5998) );
  AOI22_X1 U7817 ( .A1(n6000), .A2(n5999), .B1(n5998), .B2(n6121), .ZN(n6002)
         );
  AOI21_X1 U7818 ( .B1(n6003), .B2(n6002), .A(n6001), .ZN(n6006) );
  OAI21_X1 U7819 ( .B1(n6006), .B2(n6005), .A(n6147), .ZN(n6007) );
  NAND2_X1 U7820 ( .A1(n6007), .A2(n6153), .ZN(n6008) );
  XNOR2_X1 U7821 ( .A(n6008), .B(n9871), .ZN(n6009) );
  NAND3_X1 U7822 ( .A1(n6009), .A2(n6442), .A3(n8110), .ZN(n6014) );
  NAND2_X1 U7823 ( .A1(n10113), .A2(n6164), .ZN(n6410) );
  NAND2_X1 U7824 ( .A1(n9932), .A2(n5846), .ZN(n6012) );
  INV_X1 U7825 ( .A(P1_B_REG_SCAN_IN), .ZN(n6010) );
  AOI21_X1 U7826 ( .B1(n6442), .B2(n4590), .A(n6010), .ZN(n6011) );
  OAI21_X1 U7827 ( .B1(n6410), .B2(n6012), .A(n6011), .ZN(n6013) );
  OAI211_X1 U7828 ( .C1(n6016), .C2(n6015), .A(n6014), .B(n6013), .ZN(n6017)
         );
  INV_X1 U7829 ( .A(n6017), .ZN(n6159) );
  INV_X1 U7830 ( .A(n6018), .ZN(n6019) );
  INV_X1 U7831 ( .A(n6020), .ZN(n6021) );
  AOI22_X1 U7832 ( .A1(n6024), .A2(n6023), .B1(n6022), .B2(n6121), .ZN(n6128)
         );
  AOI21_X1 U7833 ( .B1(n7392), .B2(n6027), .A(n6025), .ZN(n6026) );
  AND2_X1 U7834 ( .A1(n6032), .A2(n6028), .ZN(n6035) );
  NAND2_X1 U7835 ( .A1(n7845), .A2(n6036), .ZN(n6042) );
  AOI21_X1 U7836 ( .B1(n6045), .B2(n6037), .A(n6042), .ZN(n6038) );
  INV_X1 U7837 ( .A(n6042), .ZN(n6043) );
  AOI21_X1 U7838 ( .B1(n6046), .B2(n5315), .A(n7850), .ZN(n6049) );
  OAI21_X1 U7839 ( .B1(n6049), .B2(n6048), .A(n6047), .ZN(n6050) );
  INV_X1 U7840 ( .A(n6059), .ZN(n6052) );
  AOI21_X1 U7841 ( .B1(n6055), .B2(n6054), .A(n6053), .ZN(n6077) );
  NAND4_X1 U7842 ( .A1(n6068), .A2(n6151), .A3(n9956), .A4(n6056), .ZN(n6076)
         );
  AOI21_X1 U7843 ( .B1(n6062), .B2(n6061), .A(n6060), .ZN(n6064) );
  NAND2_X1 U7844 ( .A1(n5829), .A2(n4788), .ZN(n6065) );
  NAND4_X1 U7845 ( .A1(n6069), .A2(n4788), .A3(n9961), .A4(n5470), .ZN(n6072)
         );
  INV_X1 U7846 ( .A(n5470), .ZN(n9615) );
  NAND4_X1 U7847 ( .A1(n6068), .A2(n9615), .A3(n6151), .A4(n9672), .ZN(n6071)
         );
  OR2_X1 U7848 ( .A1(n6069), .A2(n4788), .ZN(n6070) );
  INV_X1 U7849 ( .A(n6086), .ZN(n6089) );
  INV_X1 U7850 ( .A(n6078), .ZN(n6080) );
  OAI21_X1 U7851 ( .B1(n6151), .B2(n10051), .A(n6081), .ZN(n6079) );
  AOI21_X1 U7852 ( .B1(n6080), .B2(n6082), .A(n6079), .ZN(n6084) );
  AOI21_X1 U7853 ( .B1(n6081), .B2(n9933), .A(n6151), .ZN(n6083) );
  OAI22_X1 U7854 ( .A1(n6084), .A2(n6083), .B1(n6151), .B2(n6082), .ZN(n6088)
         );
  NOR2_X1 U7855 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  OAI211_X1 U7856 ( .C1(n6096), .C2(n6091), .A(n6098), .B(n6090), .ZN(n6094)
         );
  NAND3_X1 U7857 ( .A1(n6094), .A2(n6093), .A3(n6092), .ZN(n6095) );
  NAND3_X1 U7858 ( .A1(n6095), .A2(n6108), .A3(n6097), .ZN(n6102) );
  NAND2_X1 U7859 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  INV_X1 U7860 ( .A(n9846), .ZN(n6109) );
  INV_X1 U7861 ( .A(n6103), .ZN(n6105) );
  AOI21_X1 U7862 ( .B1(n6105), .B2(n9846), .A(n6104), .ZN(n6106) );
  OAI21_X1 U7863 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(n6110) );
  INV_X1 U7864 ( .A(n6121), .ZN(n6114) );
  NAND2_X1 U7865 ( .A1(n6112), .A2(n6115), .ZN(n6113) );
  OAI21_X1 U7866 ( .B1(n6114), .B2(n6113), .A(n4788), .ZN(n6124) );
  NAND3_X1 U7867 ( .A1(n6125), .A2(n6129), .A3(n6151), .ZN(n6123) );
  INV_X1 U7868 ( .A(n6115), .ZN(n6119) );
  INV_X1 U7869 ( .A(n6116), .ZN(n6118) );
  OAI21_X1 U7870 ( .B1(n6119), .B2(n6118), .A(n6117), .ZN(n6120) );
  NAND4_X1 U7871 ( .A1(n6129), .A2(n6151), .A3(n6121), .A4(n6120), .ZN(n6122)
         );
  OAI211_X1 U7872 ( .C1(n6125), .C2(n6124), .A(n6123), .B(n6122), .ZN(n6126)
         );
  INV_X1 U7873 ( .A(n6129), .ZN(n6130) );
  NAND2_X1 U7874 ( .A1(n6130), .A2(n4788), .ZN(n6131) );
  MUX2_X1 U7875 ( .A(n6134), .B(n6133), .S(n6151), .Z(n6135) );
  OAI21_X1 U7876 ( .B1(n6141), .B2(n9733), .A(n6137), .ZN(n6145) );
  AND2_X1 U7877 ( .A1(n9733), .A2(n9664), .ZN(n6140) );
  NAND2_X1 U7878 ( .A1(n6142), .A2(n9723), .ZN(n6143) );
  AOI211_X1 U7879 ( .C1(n4788), .C2(n4294), .A(n9871), .B(n8110), .ZN(n6148)
         );
  OAI21_X1 U7880 ( .B1(n6152), .B2(n6151), .A(n6150), .ZN(n6157) );
  INV_X1 U7881 ( .A(n6153), .ZN(n6155) );
  INV_X1 U7882 ( .A(n6442), .ZN(n8304) );
  NAND3_X1 U7883 ( .A1(n4590), .A2(n4294), .A3(n6393), .ZN(n6154) );
  AOI211_X1 U7884 ( .C1(n6155), .C2(n7856), .A(n8304), .B(n6154), .ZN(n6156)
         );
  NAND2_X1 U7885 ( .A1(n6157), .A2(n6156), .ZN(n6158) );
  NAND2_X1 U7886 ( .A1(n6165), .A2(n6164), .ZN(n6166) );
  NAND2_X1 U7887 ( .A1(n6193), .A2(n7744), .ZN(n6169) );
  INV_X1 U7888 ( .A(n4293), .ZN(n6177) );
  INV_X1 U7889 ( .A(n6172), .ZN(n6171) );
  INV_X1 U7890 ( .A(n7472), .ZN(n6181) );
  INV_X1 U7891 ( .A(n7401), .ZN(n7476) );
  OAI22_X1 U7892 ( .A1(n6419), .A2(n7405), .B1(n10139), .B2(n7143), .ZN(n6173)
         );
  NAND2_X1 U7893 ( .A1(n6364), .A2(n7725), .ZN(n6175) );
  NAND2_X1 U7894 ( .A1(n6178), .A2(n4322), .ZN(n7295) );
  NAND2_X1 U7895 ( .A1(n6178), .A2(n6379), .ZN(n6179) );
  INV_X1 U7896 ( .A(n7474), .ZN(n6180) );
  NAND2_X1 U7897 ( .A1(n7456), .A2(n7457), .ZN(n6191) );
  INV_X1 U7898 ( .A(n10228), .ZN(n7465) );
  NAND2_X1 U7899 ( .A1(n6364), .A2(n7465), .ZN(n6183) );
  OR2_X1 U7900 ( .A1(n6419), .A2(n7475), .ZN(n6182) );
  NAND2_X1 U7901 ( .A1(n6183), .A2(n6182), .ZN(n6184) );
  NAND2_X1 U7902 ( .A1(n6345), .A2(n9681), .ZN(n6187) );
  OR2_X1 U7903 ( .A1(n6419), .A2(n10228), .ZN(n6186) );
  AND2_X1 U7904 ( .A1(n6187), .A2(n6186), .ZN(n6188) );
  NAND2_X1 U7905 ( .A1(n6189), .A2(n6188), .ZN(n6192) );
  AND2_X1 U7906 ( .A1(n6190), .A2(n6192), .ZN(n7458) );
  NAND2_X1 U7907 ( .A1(n6191), .A2(n7458), .ZN(n7460) );
  NAND2_X1 U7908 ( .A1(n7460), .A2(n6192), .ZN(n7581) );
  NAND2_X1 U7909 ( .A1(n6193), .A2(n7690), .ZN(n6195) );
  OR2_X1 U7910 ( .A1(n6419), .A2(n7604), .ZN(n6194) );
  NAND2_X1 U7911 ( .A1(n6195), .A2(n6194), .ZN(n6196) );
  XNOR2_X1 U7912 ( .A(n6196), .B(n6379), .ZN(n6210) );
  OR2_X1 U7913 ( .A1(n6419), .A2(n10239), .ZN(n6197) );
  OAI21_X1 U7914 ( .B1(n6424), .B2(n7604), .A(n6197), .ZN(n6208) );
  XNOR2_X1 U7915 ( .A(n6210), .B(n6208), .ZN(n7582) );
  NAND2_X1 U7916 ( .A1(n6193), .A2(n7708), .ZN(n6199) );
  OR2_X1 U7917 ( .A1(n6419), .A2(n7577), .ZN(n6198) );
  NAND2_X1 U7918 ( .A1(n6199), .A2(n6198), .ZN(n6200) );
  XNOR2_X1 U7919 ( .A(n4293), .B(n6200), .ZN(n7600) );
  NAND2_X1 U7920 ( .A1(n6345), .A2(n9679), .ZN(n6202) );
  NAND2_X1 U7921 ( .A1(n4289), .A2(n7708), .ZN(n6201) );
  NAND2_X1 U7922 ( .A1(n6202), .A2(n6201), .ZN(n7598) );
  NAND2_X1 U7923 ( .A1(n10253), .A2(n6193), .ZN(n6204) );
  OR2_X1 U7924 ( .A1(n6419), .A2(n7736), .ZN(n6203) );
  NAND2_X1 U7925 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  XNOR2_X1 U7926 ( .A(n6205), .B(n6379), .ZN(n7752) );
  NAND2_X1 U7927 ( .A1(n10253), .A2(n4289), .ZN(n6207) );
  NAND2_X1 U7928 ( .A1(n6345), .A2(n4587), .ZN(n6206) );
  AND2_X1 U7929 ( .A1(n6207), .A2(n6206), .ZN(n7751) );
  NAND2_X1 U7930 ( .A1(n7752), .A2(n7751), .ZN(n6211) );
  INV_X1 U7931 ( .A(n6208), .ZN(n6209) );
  NAND2_X1 U7932 ( .A1(n6210), .A2(n6209), .ZN(n7601) );
  OAI211_X1 U7933 ( .C1(n7600), .C2(n7598), .A(n6211), .B(n7601), .ZN(n6212)
         );
  INV_X1 U7934 ( .A(n6212), .ZN(n6213) );
  INV_X1 U7935 ( .A(n7752), .ZN(n6217) );
  NAND2_X1 U7936 ( .A1(n7600), .A2(n7598), .ZN(n7749) );
  NAND2_X1 U7937 ( .A1(n7749), .A2(n7751), .ZN(n6216) );
  INV_X1 U7938 ( .A(n7749), .ZN(n6215) );
  INV_X1 U7939 ( .A(n7751), .ZN(n6214) );
  AOI22_X1 U7940 ( .A1(n6217), .A2(n6216), .B1(n6215), .B2(n6214), .ZN(n6218)
         );
  NAND2_X1 U7941 ( .A1(n10260), .A2(n4288), .ZN(n6220) );
  OR2_X1 U7942 ( .A1(n6419), .A2(n7756), .ZN(n6219) );
  NAND2_X1 U7943 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  XNOR2_X1 U7944 ( .A(n6221), .B(n6379), .ZN(n6223) );
  NOR2_X1 U7945 ( .A1(n6424), .A2(n7756), .ZN(n6222) );
  AOI21_X1 U7946 ( .B1(n10260), .B2(n4289), .A(n6222), .ZN(n6224) );
  NAND2_X1 U7947 ( .A1(n6223), .A2(n6224), .ZN(n7731) );
  INV_X1 U7948 ( .A(n6223), .ZN(n6226) );
  INV_X1 U7949 ( .A(n6224), .ZN(n6225) );
  NAND2_X1 U7950 ( .A1(n6226), .A2(n6225), .ZN(n7732) );
  NAND2_X1 U7951 ( .A1(n7868), .A2(n4289), .ZN(n6228) );
  NAND2_X1 U7952 ( .A1(n6345), .A2(n9677), .ZN(n6227) );
  NAND2_X1 U7953 ( .A1(n6228), .A2(n6227), .ZN(n7863) );
  NAND2_X1 U7954 ( .A1(n7868), .A2(n4288), .ZN(n6230) );
  OR2_X1 U7955 ( .A1(n6419), .A2(n8230), .ZN(n6229) );
  NAND2_X1 U7956 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  XNOR2_X1 U7957 ( .A(n4293), .B(n6231), .ZN(n7864) );
  NAND2_X1 U7958 ( .A1(n8235), .A2(n4288), .ZN(n6233) );
  OR2_X1 U7959 ( .A1(n6419), .A2(n8264), .ZN(n6232) );
  NAND2_X1 U7960 ( .A1(n6233), .A2(n6232), .ZN(n6234) );
  XNOR2_X1 U7961 ( .A(n6234), .B(n6379), .ZN(n8226) );
  NOR2_X1 U7962 ( .A1(n6424), .A2(n8264), .ZN(n6235) );
  AOI21_X1 U7963 ( .B1(n8235), .B2(n4289), .A(n6235), .ZN(n6241) );
  NAND2_X1 U7964 ( .A1(n8226), .A2(n6241), .ZN(n6236) );
  NAND2_X1 U7965 ( .A1(n8128), .A2(n4288), .ZN(n6238) );
  OR2_X1 U7966 ( .A1(n6419), .A2(n7890), .ZN(n6237) );
  NAND2_X1 U7967 ( .A1(n6238), .A2(n6237), .ZN(n6239) );
  XNOR2_X1 U7968 ( .A(n4293), .B(n6239), .ZN(n6244) );
  NOR2_X1 U7969 ( .A1(n6424), .A2(n7890), .ZN(n6240) );
  AOI21_X1 U7970 ( .B1(n8128), .B2(n4289), .A(n6240), .ZN(n6245) );
  XNOR2_X1 U7971 ( .A(n6244), .B(n6245), .ZN(n8258) );
  INV_X1 U7972 ( .A(n8226), .ZN(n6242) );
  INV_X1 U7973 ( .A(n6241), .ZN(n8228) );
  NAND2_X1 U7974 ( .A1(n6242), .A2(n8228), .ZN(n6243) );
  INV_X1 U7975 ( .A(n6244), .ZN(n6246) );
  NAND2_X1 U7976 ( .A1(n6246), .A2(n6245), .ZN(n6247) );
  NAND2_X1 U7977 ( .A1(n8325), .A2(n4288), .ZN(n6249) );
  OR2_X1 U7978 ( .A1(n6419), .A2(n7993), .ZN(n6248) );
  NAND2_X1 U7979 ( .A1(n6249), .A2(n6248), .ZN(n6250) );
  XNOR2_X1 U7980 ( .A(n6250), .B(n6379), .ZN(n6252) );
  INV_X1 U7981 ( .A(n6252), .ZN(n6251) );
  NAND2_X1 U7982 ( .A1(n6253), .A2(n6252), .ZN(n8360) );
  NAND2_X1 U7983 ( .A1(n8325), .A2(n4289), .ZN(n6256) );
  NAND2_X1 U7984 ( .A1(n6345), .A2(n9674), .ZN(n6255) );
  NAND2_X1 U7985 ( .A1(n6256), .A2(n6255), .ZN(n8318) );
  INV_X1 U7986 ( .A(n8318), .ZN(n6257) );
  OAI22_X1 U7987 ( .A1(n8370), .A2(n6371), .B1(n8320), .B2(n6419), .ZN(n6258)
         );
  XNOR2_X1 U7988 ( .A(n4293), .B(n6258), .ZN(n6260) );
  OAI22_X1 U7989 ( .A1(n8370), .A2(n6419), .B1(n8320), .B2(n6424), .ZN(n6259)
         );
  NAND2_X1 U7990 ( .A1(n6260), .A2(n6259), .ZN(n6261) );
  AND2_X1 U7991 ( .A1(n9539), .A2(n6261), .ZN(n8361) );
  NAND2_X1 U7992 ( .A1(n5450), .A2(n4288), .ZN(n6263) );
  OR2_X1 U7993 ( .A1(n6419), .A2(n9610), .ZN(n6262) );
  NAND2_X1 U7994 ( .A1(n6263), .A2(n6262), .ZN(n6264) );
  XNOR2_X1 U7995 ( .A(n6264), .B(n6379), .ZN(n6266) );
  NOR2_X1 U7996 ( .A1(n6424), .A2(n9610), .ZN(n6265) );
  AOI21_X1 U7997 ( .B1(n5450), .B2(n4289), .A(n6265), .ZN(n6267) );
  NAND2_X1 U7998 ( .A1(n6266), .A2(n6267), .ZN(n6271) );
  INV_X1 U7999 ( .A(n6266), .ZN(n6269) );
  INV_X1 U8000 ( .A(n6267), .ZN(n6268) );
  NAND2_X1 U8001 ( .A1(n6269), .A2(n6268), .ZN(n6270) );
  AND2_X1 U8002 ( .A1(n6271), .A2(n6270), .ZN(n9540) );
  NAND2_X1 U8003 ( .A1(n5470), .A2(n4288), .ZN(n6273) );
  OR2_X1 U8004 ( .A1(n6419), .A2(n9961), .ZN(n6272) );
  NAND2_X1 U8005 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  XNOR2_X1 U8006 ( .A(n4293), .B(n6274), .ZN(n6276) );
  NOR2_X1 U8007 ( .A1(n6424), .A2(n9961), .ZN(n6275) );
  AOI21_X1 U8008 ( .B1(n5470), .B2(n4289), .A(n6275), .ZN(n6277) );
  XNOR2_X1 U8009 ( .A(n6276), .B(n6277), .ZN(n9606) );
  INV_X1 U8010 ( .A(n6276), .ZN(n6278) );
  NAND2_X1 U8011 ( .A1(n6278), .A2(n6277), .ZN(n6279) );
  OAI22_X1 U8012 ( .A1(n10108), .A2(n6371), .B1(n9918), .B2(n6419), .ZN(n6280)
         );
  XNOR2_X1 U8013 ( .A(n4293), .B(n6280), .ZN(n6295) );
  OR2_X1 U8014 ( .A1(n10108), .A2(n6419), .ZN(n6282) );
  NAND2_X1 U8015 ( .A1(n9669), .A2(n6345), .ZN(n6281) );
  NAND2_X1 U8016 ( .A1(n6282), .A2(n6281), .ZN(n6296) );
  NAND2_X1 U8017 ( .A1(n6295), .A2(n6296), .ZN(n9569) );
  NAND2_X1 U8018 ( .A1(n10051), .A2(n4288), .ZN(n6284) );
  NAND2_X1 U8019 ( .A1(n9933), .A2(n4289), .ZN(n6283) );
  NAND2_X1 U8020 ( .A1(n6284), .A2(n6283), .ZN(n6285) );
  XNOR2_X1 U8021 ( .A(n4293), .B(n6285), .ZN(n9564) );
  NAND2_X1 U8022 ( .A1(n10051), .A2(n4289), .ZN(n6287) );
  NAND2_X1 U8023 ( .A1(n9933), .A2(n6345), .ZN(n6286) );
  NAND2_X1 U8024 ( .A1(n6287), .A2(n6286), .ZN(n9651) );
  NAND2_X1 U8025 ( .A1(n9564), .A2(n9651), .ZN(n6288) );
  NAND2_X1 U8026 ( .A1(n9569), .A2(n6288), .ZN(n6294) );
  OAI22_X1 U8027 ( .A1(n5832), .A2(n6371), .B1(n9655), .B2(n6419), .ZN(n6289)
         );
  XNOR2_X1 U8028 ( .A(n4293), .B(n6289), .ZN(n9500) );
  OR2_X1 U8029 ( .A1(n5832), .A2(n6419), .ZN(n6291) );
  NAND2_X1 U8030 ( .A1(n6345), .A2(n9671), .ZN(n6290) );
  NAND2_X1 U8031 ( .A1(n6291), .A2(n6290), .ZN(n9498) );
  AND2_X1 U8032 ( .A1(n9500), .A2(n9498), .ZN(n6292) );
  NOR2_X1 U8033 ( .A1(n6294), .A2(n6292), .ZN(n6293) );
  INV_X1 U8034 ( .A(n6294), .ZN(n6300) );
  OAI22_X1 U8035 ( .A1(n9564), .A2(n9651), .B1(n9500), .B2(n9498), .ZN(n6299)
         );
  INV_X1 U8036 ( .A(n6295), .ZN(n6298) );
  INV_X1 U8037 ( .A(n6296), .ZN(n6297) );
  AND2_X1 U8038 ( .A1(n6298), .A2(n6297), .ZN(n9570) );
  AOI21_X1 U8039 ( .B1(n6300), .B2(n6299), .A(n9570), .ZN(n6301) );
  NAND2_X1 U8040 ( .A1(n10039), .A2(n4288), .ZN(n6303) );
  NAND2_X1 U8041 ( .A1(n9935), .A2(n4289), .ZN(n6302) );
  NAND2_X1 U8042 ( .A1(n6303), .A2(n6302), .ZN(n6304) );
  XNOR2_X1 U8043 ( .A(n4293), .B(n6304), .ZN(n6306) );
  NOR2_X1 U8044 ( .A1(n9899), .A2(n6424), .ZN(n6305) );
  AOI21_X1 U8045 ( .B1(n10039), .B2(n4289), .A(n6305), .ZN(n6307) );
  XNOR2_X1 U8046 ( .A(n6306), .B(n6307), .ZN(n9579) );
  INV_X1 U8047 ( .A(n6306), .ZN(n6308) );
  NAND2_X1 U8048 ( .A1(n10027), .A2(n4288), .ZN(n6310) );
  OR2_X1 U8049 ( .A1(n9898), .A2(n6419), .ZN(n6309) );
  NAND2_X1 U8050 ( .A1(n6310), .A2(n6309), .ZN(n6311) );
  XNOR2_X1 U8051 ( .A(n4293), .B(n6311), .ZN(n9522) );
  NAND2_X1 U8052 ( .A1(n10027), .A2(n4289), .ZN(n6313) );
  OR2_X1 U8053 ( .A1(n9898), .A2(n6424), .ZN(n6312) );
  NAND2_X1 U8054 ( .A1(n6313), .A2(n6312), .ZN(n6320) );
  NAND2_X1 U8055 ( .A1(n10031), .A2(n4288), .ZN(n6315) );
  NAND2_X1 U8056 ( .A1(n9883), .A2(n4289), .ZN(n6314) );
  NAND2_X1 U8057 ( .A1(n6315), .A2(n6314), .ZN(n6316) );
  XNOR2_X1 U8058 ( .A(n4293), .B(n6316), .ZN(n6321) );
  NAND2_X1 U8059 ( .A1(n10031), .A2(n4289), .ZN(n6318) );
  NAND2_X1 U8060 ( .A1(n9883), .A2(n6345), .ZN(n6317) );
  NAND2_X1 U8061 ( .A1(n6318), .A2(n6317), .ZN(n9632) );
  OAI22_X1 U8062 ( .A1(n9522), .A2(n6320), .B1(n6321), .B2(n9632), .ZN(n6325)
         );
  INV_X1 U8063 ( .A(n6321), .ZN(n9520) );
  INV_X1 U8064 ( .A(n9632), .ZN(n6319) );
  INV_X1 U8065 ( .A(n6320), .ZN(n9521) );
  OAI21_X1 U8066 ( .B1(n9520), .B2(n6319), .A(n9521), .ZN(n6323) );
  AND2_X1 U8067 ( .A1(n6320), .A2(n9632), .ZN(n6322) );
  AOI22_X1 U8068 ( .A1(n9522), .A2(n6323), .B1(n6322), .B2(n6321), .ZN(n6324)
         );
  NAND2_X1 U8069 ( .A1(n10020), .A2(n4288), .ZN(n6327) );
  NAND2_X1 U8070 ( .A1(n9882), .A2(n4289), .ZN(n6326) );
  NAND2_X1 U8071 ( .A1(n6327), .A2(n6326), .ZN(n6328) );
  XNOR2_X1 U8072 ( .A(n6328), .B(n6379), .ZN(n9596) );
  NOR2_X1 U8073 ( .A1(n9527), .A2(n6424), .ZN(n6329) );
  AOI21_X1 U8074 ( .B1(n10020), .B2(n4289), .A(n6329), .ZN(n6331) );
  NAND2_X1 U8075 ( .A1(n9596), .A2(n6331), .ZN(n6330) );
  INV_X1 U8076 ( .A(n9596), .ZN(n6332) );
  INV_X1 U8077 ( .A(n6331), .ZN(n9595) );
  NAND2_X1 U8078 ( .A1(n6332), .A2(n9595), .ZN(n6333) );
  NAND2_X1 U8079 ( .A1(n10014), .A2(n4288), .ZN(n6335) );
  NAND2_X1 U8080 ( .A1(n9836), .A2(n4289), .ZN(n6334) );
  NAND2_X1 U8081 ( .A1(n6335), .A2(n6334), .ZN(n6336) );
  XNOR2_X1 U8082 ( .A(n6336), .B(n6379), .ZN(n6339) );
  NOR2_X1 U8083 ( .A1(n9869), .A2(n6424), .ZN(n6337) );
  AOI21_X1 U8084 ( .B1(n10014), .B2(n4289), .A(n6337), .ZN(n6338) );
  XNOR2_X1 U8085 ( .A(n6339), .B(n6338), .ZN(n9532) );
  NAND2_X1 U8086 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  NAND2_X1 U8087 ( .A1(n9825), .A2(n4288), .ZN(n6343) );
  NAND2_X1 U8088 ( .A1(n9835), .A2(n4289), .ZN(n6342) );
  NAND2_X1 U8089 ( .A1(n6343), .A2(n6342), .ZN(n6344) );
  XNOR2_X1 U8090 ( .A(n4293), .B(n6344), .ZN(n6354) );
  NAND2_X1 U8091 ( .A1(n9825), .A2(n4289), .ZN(n6347) );
  NAND2_X1 U8092 ( .A1(n9835), .A2(n6345), .ZN(n6346) );
  NAND2_X1 U8093 ( .A1(n6347), .A2(n6346), .ZN(n6355) );
  NAND2_X1 U8094 ( .A1(n6354), .A2(n6355), .ZN(n9512) );
  INV_X1 U8095 ( .A(n9512), .ZN(n6353) );
  NAND2_X1 U8096 ( .A1(n10009), .A2(n4288), .ZN(n6349) );
  NAND2_X1 U8097 ( .A1(n9860), .A2(n4289), .ZN(n6348) );
  NAND2_X1 U8098 ( .A1(n6349), .A2(n6348), .ZN(n6350) );
  XNOR2_X1 U8099 ( .A(n6350), .B(n6379), .ZN(n9510) );
  NOR2_X1 U8100 ( .A1(n9824), .A2(n6424), .ZN(n6351) );
  AOI21_X1 U8101 ( .B1(n10009), .B2(n4289), .A(n6351), .ZN(n9618) );
  NAND3_X1 U8102 ( .A1(n9512), .A2(n9618), .A3(n9510), .ZN(n6358) );
  INV_X1 U8103 ( .A(n6354), .ZN(n6357) );
  INV_X1 U8104 ( .A(n6355), .ZN(n6356) );
  NAND2_X1 U8105 ( .A1(n6357), .A2(n6356), .ZN(n9586) );
  AOI22_X1 U8106 ( .A1(n5839), .A2(n4288), .B1(n4289), .B2(n9667), .ZN(n6360)
         );
  XOR2_X1 U8107 ( .A(n4293), .B(n6360), .Z(n6362) );
  OAI22_X1 U8108 ( .A1(n10087), .A2(n6419), .B1(n9823), .B2(n6424), .ZN(n6361)
         );
  NOR2_X1 U8109 ( .A1(n6362), .A2(n6361), .ZN(n6363) );
  AOI21_X1 U8110 ( .B1(n6362), .B2(n6361), .A(n6363), .ZN(n9588) );
  OAI22_X1 U8111 ( .A1(n10083), .A2(n6419), .B1(n9810), .B2(n6424), .ZN(n6368)
         );
  NAND2_X1 U8112 ( .A1(n9790), .A2(n4288), .ZN(n6366) );
  NAND2_X1 U8113 ( .A1(n5715), .A2(n4289), .ZN(n6365) );
  NAND2_X1 U8114 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  XNOR2_X1 U8115 ( .A(n4293), .B(n6367), .ZN(n6369) );
  XOR2_X1 U8116 ( .A(n6368), .B(n6369), .Z(n9554) );
  OR2_X1 U8117 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  OAI22_X1 U8118 ( .A1(n10079), .A2(n6371), .B1(n9795), .B2(n6419), .ZN(n6372)
         );
  XNOR2_X1 U8119 ( .A(n4293), .B(n6372), .ZN(n6373) );
  OAI22_X1 U8120 ( .A1(n10079), .A2(n6419), .B1(n9795), .B2(n6424), .ZN(n6374)
         );
  XNOR2_X1 U8121 ( .A(n6373), .B(n6374), .ZN(n9646) );
  INV_X1 U8122 ( .A(n6373), .ZN(n6376) );
  INV_X1 U8123 ( .A(n6374), .ZN(n6375) );
  NAND2_X1 U8124 ( .A1(n9987), .A2(n4288), .ZN(n6378) );
  NAND2_X1 U8125 ( .A1(n4698), .A2(n4289), .ZN(n6377) );
  NAND2_X1 U8126 ( .A1(n6378), .A2(n6377), .ZN(n6380) );
  XNOR2_X1 U8127 ( .A(n6380), .B(n6379), .ZN(n6384) );
  NOR2_X1 U8128 ( .A1(n9778), .A2(n6424), .ZN(n6382) );
  AOI21_X1 U8129 ( .B1(n9987), .B2(n4289), .A(n6382), .ZN(n6383) );
  NAND2_X1 U8130 ( .A1(n6384), .A2(n6383), .ZN(n6429) );
  OR2_X1 U8131 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  NAND2_X1 U8132 ( .A1(n6429), .A2(n6385), .ZN(n6386) );
  INV_X1 U8133 ( .A(n7611), .ZN(n6390) );
  NAND3_X1 U8134 ( .A1(n6390), .A2(n7612), .A3(n6389), .ZN(n6412) );
  NOR2_X1 U8135 ( .A1(n10261), .A2(n6444), .ZN(n6400) );
  NAND2_X1 U8136 ( .A1(n6400), .A2(n10113), .ZN(n6391) );
  NAND2_X1 U8137 ( .A1(n6394), .A2(n6393), .ZN(n7621) );
  INV_X1 U8138 ( .A(n7621), .ZN(n6395) );
  NAND2_X1 U8139 ( .A1(n10113), .A2(n6395), .ZN(n6396) );
  OR2_X1 U8140 ( .A1(n6412), .A2(n6396), .ZN(n6399) );
  INV_X1 U8141 ( .A(n6397), .ZN(n6398) );
  NAND2_X1 U8142 ( .A1(n6412), .A2(n6400), .ZN(n6403) );
  AND2_X1 U8143 ( .A1(n6401), .A2(n7143), .ZN(n6402) );
  NAND2_X1 U8144 ( .A1(n6403), .A2(n6402), .ZN(n7299) );
  NAND2_X1 U8145 ( .A1(n7299), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6408) );
  INV_X1 U8146 ( .A(n7718), .ZN(n6404) );
  NAND2_X1 U8147 ( .A1(n10113), .A2(n6404), .ZN(n6405) );
  OAI21_X1 U8148 ( .B1(n7621), .B2(P1_U3086), .A(n6405), .ZN(n6406) );
  NAND2_X1 U8149 ( .A1(n6412), .A2(n6406), .ZN(n7297) );
  AND2_X1 U8150 ( .A1(n7297), .A2(n8304), .ZN(n6407) );
  OR2_X1 U8151 ( .A1(n6410), .A2(n9962), .ZN(n6409) );
  NAND2_X1 U8152 ( .A1(n9665), .A2(n9652), .ZN(n6414) );
  INV_X1 U8153 ( .A(n9795), .ZN(n9666) );
  OR2_X1 U8154 ( .A1(n6410), .A2(n9960), .ZN(n6411) );
  AOI22_X1 U8155 ( .A1(n9666), .A2(n9640), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3086), .ZN(n6413) );
  OAI211_X1 U8156 ( .C1(n9636), .C2(n9761), .A(n6414), .B(n6413), .ZN(n6415)
         );
  INV_X1 U8157 ( .A(n6415), .ZN(n6416) );
  NAND2_X1 U8158 ( .A1(n7140), .A2(n4288), .ZN(n6421) );
  OR2_X1 U8159 ( .A1(n9766), .A2(n6419), .ZN(n6420) );
  NAND2_X1 U8160 ( .A1(n6421), .A2(n6420), .ZN(n6423) );
  XNOR2_X1 U8161 ( .A(n4293), .B(n6423), .ZN(n6427) );
  NOR2_X1 U8162 ( .A1(n9766), .A2(n6424), .ZN(n6425) );
  AOI21_X1 U8163 ( .B1(n7140), .B2(n4289), .A(n6425), .ZN(n6426) );
  XNOR2_X1 U8164 ( .A(n6427), .B(n6426), .ZN(n6431) );
  INV_X1 U8165 ( .A(n6431), .ZN(n6428) );
  INV_X1 U8166 ( .A(n6429), .ZN(n6430) );
  NAND3_X1 U8167 ( .A1(n6431), .A2(n9621), .A3(n6430), .ZN(n6437) );
  INV_X1 U8168 ( .A(n9753), .ZN(n6433) );
  OAI22_X1 U8169 ( .A1(n6433), .A2(n9636), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6432), .ZN(n6435) );
  OAI22_X1 U8170 ( .A1(n7729), .A2(n9643), .B1(n9778), .B2(n9654), .ZN(n6434)
         );
  AOI211_X1 U8171 ( .C1(n7140), .C2(n9659), .A(n6435), .B(n6434), .ZN(n6436)
         );
  NAND2_X1 U8172 ( .A1(n6441), .A2(n6440), .ZN(P1_U3220) );
  OR2_X1 U8173 ( .A1(n10113), .A2(n6442), .ZN(n6483) );
  AOI21_X1 U8174 ( .B1(n7144), .B2(n6444), .A(n6443), .ZN(n6482) );
  NAND2_X1 U8175 ( .A1(n6483), .A2(n6482), .ZN(n10143) );
  OR2_X1 U8176 ( .A1(n7518), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U8177 ( .A(n7518), .B(n10046), .ZN(n10173) );
  AND2_X1 U8178 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9687) );
  NAND2_X1 U8179 ( .A1(n9685), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6445) );
  XNOR2_X1 U8180 ( .A(n7538), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n7544) );
  INV_X1 U8181 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6446) );
  OR2_X1 U8182 ( .A1(n7538), .A2(n6446), .ZN(n6447) );
  XNOR2_X1 U8183 ( .A(n9693), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n9703) );
  OR2_X1 U8184 ( .A1(n9693), .A2(n6448), .ZN(n6449) );
  NAND2_X1 U8185 ( .A1(n9701), .A2(n6449), .ZN(n7531) );
  XNOR2_X1 U8186 ( .A(n6470), .B(n6450), .ZN(n7532) );
  MUX2_X1 U8187 ( .A(n6451), .B(P1_REG1_REG_5__SCAN_IN), .S(n9714), .Z(n9708)
         );
  MUX2_X1 U8188 ( .A(n6452), .B(P1_REG1_REG_6__SCAN_IN), .S(n7647), .Z(n7641)
         );
  NOR2_X1 U8189 ( .A1(n7642), .A2(n7641), .ZN(n7640) );
  MUX2_X1 U8190 ( .A(n6453), .B(P1_REG1_REG_7__SCAN_IN), .S(n7676), .Z(n7672)
         );
  NOR2_X1 U8191 ( .A1(n7673), .A2(n7672), .ZN(n7671) );
  XNOR2_X1 U8192 ( .A(n7665), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n7660) );
  MUX2_X1 U8193 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n6454), .S(n7190), .Z(n7505)
         );
  XNOR2_X1 U8194 ( .A(n7202), .B(P1_REG1_REG_10__SCAN_IN), .ZN(n7810) );
  XNOR2_X1 U8195 ( .A(n7234), .B(P1_REG1_REG_11__SCAN_IN), .ZN(n8021) );
  XOR2_X1 U8196 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7263), .Z(n8182) );
  XNOR2_X1 U8197 ( .A(n7268), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n8340) );
  XNOR2_X1 U8198 ( .A(n10153), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n10149) );
  INV_X1 U8199 ( .A(n10167), .ZN(n7421) );
  NOR2_X1 U8200 ( .A1(n6455), .A2(n7421), .ZN(n6456) );
  INV_X1 U8201 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10160) );
  XNOR2_X1 U8202 ( .A(n10185), .B(n6458), .ZN(n10191) );
  OR2_X1 U8203 ( .A1(n10185), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n6459) );
  NAND2_X1 U8204 ( .A1(n10200), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6462) );
  OR2_X1 U8205 ( .A1(n10200), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n6461) );
  NAND2_X1 U8206 ( .A1(n6462), .A2(n6461), .ZN(n10207) );
  NAND2_X1 U8207 ( .A1(n10210), .A2(n6462), .ZN(n6463) );
  XNOR2_X1 U8208 ( .A(n10185), .B(n6464), .ZN(n10188) );
  INV_X1 U8209 ( .A(n9714), .ZN(n7169) );
  INV_X1 U8210 ( .A(n6470), .ZN(n7527) );
  INV_X1 U8211 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6465) );
  MUX2_X1 U8212 ( .A(n6465), .B(P1_REG2_REG_1__SCAN_IN), .S(n7155), .Z(n9684)
         );
  AND2_X1 U8213 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9683) );
  NAND2_X1 U8214 ( .A1(n9685), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6466) );
  NAND2_X1 U8215 ( .A1(n9682), .A2(n6466), .ZN(n7540) );
  OR2_X1 U8216 ( .A1(n7538), .A2(n6467), .ZN(n6468) );
  XNOR2_X1 U8217 ( .A(n9693), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n9700) );
  OR2_X1 U8218 ( .A1(n9693), .A2(n5179), .ZN(n6469) );
  NAND2_X1 U8219 ( .A1(n9698), .A2(n6469), .ZN(n7529) );
  XNOR2_X1 U8220 ( .A(n6470), .B(n6471), .ZN(n7530) );
  NAND2_X1 U8221 ( .A1(n7529), .A2(n7530), .ZN(n7528) );
  MUX2_X1 U8222 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7618), .S(n9714), .Z(n9718)
         );
  MUX2_X1 U8223 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7767), .S(n7647), .Z(n7643)
         );
  XNOR2_X1 U8224 ( .A(n7676), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n7675) );
  NOR2_X1 U8225 ( .A1(n4321), .A2(n7675), .ZN(n7674) );
  XNOR2_X1 U8226 ( .A(n7665), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n7663) );
  NOR2_X1 U8227 ( .A1(n7664), .A2(n7663), .ZN(n7662) );
  XNOR2_X1 U8228 ( .A(n7190), .B(n6472), .ZN(n7510) );
  XNOR2_X1 U8229 ( .A(n7202), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n7813) );
  XNOR2_X1 U8230 ( .A(n7234), .B(P1_REG2_REG_11__SCAN_IN), .ZN(n8024) );
  XNOR2_X1 U8231 ( .A(n7263), .B(n8122), .ZN(n8186) );
  XNOR2_X1 U8232 ( .A(n7268), .B(P1_REG2_REG_13__SCAN_IN), .ZN(n8343) );
  NAND2_X1 U8233 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n10153), .ZN(n6473) );
  OAI21_X1 U8234 ( .B1(n10153), .B2(P1_REG2_REG_14__SCAN_IN), .A(n6473), .ZN(
        n10146) );
  NOR2_X1 U8235 ( .A1(n6474), .A2(n7421), .ZN(n6475) );
  INV_X1 U8236 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n10163) );
  NAND2_X1 U8237 ( .A1(n7518), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n6476) );
  OAI21_X1 U8238 ( .B1(n7518), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6476), .ZN(
        n10177) );
  OR2_X1 U8239 ( .A1(n10185), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6477) );
  NAND2_X1 U8240 ( .A1(n10200), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6479) );
  OR2_X1 U8241 ( .A1(n10200), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8242 ( .A1(n6479), .A2(n6478), .ZN(n10201) );
  NAND2_X1 U8243 ( .A1(n10204), .A2(n6479), .ZN(n6480) );
  INV_X1 U8244 ( .A(n10143), .ZN(n6490) );
  AND2_X1 U8245 ( .A1(n5846), .A2(n7524), .ZN(n6481) );
  OAI22_X1 U8246 ( .A1(n10158), .A2(n6489), .B1(n6488), .B2(n10206), .ZN(n6487) );
  INV_X1 U8247 ( .A(n6482), .ZN(n6484) );
  NAND2_X1 U8248 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9525) );
  NAND2_X1 U8249 ( .A1(n6490), .A2(n4675), .ZN(n10215) );
  NAND3_X1 U8250 ( .A1(n6497), .A2(n6496), .A3(n6495), .ZN(n6505) );
  INV_X1 U8251 ( .A(n6505), .ZN(n6499) );
  NOR2_X1 U8252 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n6498) );
  NAND2_X1 U8253 ( .A1(n6509), .A2(n6513), .ZN(n6501) );
  OAI21_X1 U8254 ( .B1(n6508), .B2(n6501), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6502) );
  MUX2_X1 U8255 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6502), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6507) );
  NAND4_X1 U8256 ( .A1(n6509), .A2(n6513), .A3(n6500), .A4(n6503), .ZN(n6504)
         );
  NAND2_X1 U8257 ( .A1(n6507), .A2(n6527), .ZN(n9492) );
  NOR2_X1 U8258 ( .A1(n9492), .A2(n7083), .ZN(n6516) );
  INV_X1 U8259 ( .A(n7085), .ZN(n6515) );
  NAND2_X1 U8260 ( .A1(n6516), .A2(n6515), .ZN(n7334) );
  NAND2_X1 U8261 ( .A1(n6517), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6518) );
  XNOR2_X1 U8262 ( .A(n6518), .B(n6500), .ZN(n8308) );
  INV_X1 U8263 ( .A(n7149), .ZN(n6519) );
  INV_X1 U8264 ( .A(n8308), .ZN(n6520) );
  OR2_X1 U8265 ( .A1(n7334), .A2(n6520), .ZN(n6676) );
  NAND2_X1 U8266 ( .A1(n6532), .A2(n6521), .ZN(n7040) );
  OAI21_X1 U8267 ( .B1(n6524), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6522) );
  MUX2_X1 U8268 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6522), .S(
        P2_IR_REG_22__SCAN_IN), .Z(n6523) );
  NAND2_X1 U8269 ( .A1(n6524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6525) );
  NOR2_X4 U8270 ( .A1(n8415), .A2(n4742), .ZN(n8515) );
  NAND2_X1 U8271 ( .A1(n8515), .A2(n8308), .ZN(n6526) );
  NAND2_X1 U8272 ( .A1(n6676), .A2(n6526), .ZN(n6677) );
  OAI21_X1 U8273 ( .B1(n6677), .B2(n6929), .A(P2_STATE_REG_SCAN_IN), .ZN(
        P2_U3150) );
  NAND2_X1 U8274 ( .A1(n6532), .A2(n6531), .ZN(n6579) );
  INV_X1 U8275 ( .A(n6579), .ZN(n6534) );
  NAND2_X1 U8276 ( .A1(n6534), .A2(n6533), .ZN(n6544) );
  INV_X1 U8277 ( .A(n6544), .ZN(n6536) );
  INV_X1 U8278 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6537) );
  NAND2_X1 U8279 ( .A1(n6584), .A2(n6537), .ZN(n6592) );
  INV_X1 U8280 ( .A(n6592), .ZN(n6539) );
  NAND4_X1 U8281 ( .A1(n6539), .A2(n6538), .A3(n6595), .A4(n6600), .ZN(n6540)
         );
  NAND2_X1 U8282 ( .A1(n4333), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6541) );
  MUX2_X1 U8283 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6541), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6543) );
  NAND2_X1 U8284 ( .A1(n6543), .A2(n6609), .ZN(n9058) );
  INV_X1 U8285 ( .A(n9058), .ZN(n6895) );
  INV_X1 U8286 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9250) );
  NAND2_X1 U8287 ( .A1(n6544), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6545) );
  XNOR2_X1 U8288 ( .A(n6545), .B(P2_IR_REG_10__SCAN_IN), .ZN(n8147) );
  INV_X1 U8289 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8172) );
  INV_X1 U8290 ( .A(n6569), .ZN(n6547) );
  INV_X1 U8291 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U8292 ( .A1(n6547), .A2(n6546), .ZN(n6572) );
  NAND2_X1 U8293 ( .A1(n6549), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6548) );
  MUX2_X1 U8294 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6548), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n6552) );
  INV_X1 U8295 ( .A(n6549), .ZN(n6551) );
  NAND2_X1 U8296 ( .A1(n6551), .A2(n6550), .ZN(n6574) );
  NAND2_X1 U8297 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6494), .ZN(n6554) );
  INV_X1 U8298 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7453) );
  NAND2_X1 U8299 ( .A1(n6553), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6563) );
  INV_X1 U8300 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7219) );
  INV_X1 U8301 ( .A(n6563), .ZN(n6564) );
  NAND2_X1 U8302 ( .A1(n4304), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6566) );
  MUX2_X1 U8303 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6566), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6567) );
  NAND2_X1 U8304 ( .A1(n6569), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6570) );
  INV_X1 U8305 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6771) );
  XNOR2_X1 U8306 ( .A(n7286), .B(n6771), .ZN(n7271) );
  NAND2_X1 U8307 ( .A1(n6572), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6573) );
  XNOR2_X1 U8308 ( .A(n6573), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7316) );
  XNOR2_X1 U8309 ( .A(n7175), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n8949) );
  NAND2_X1 U8310 ( .A1(n6574), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6575) );
  INV_X1 U8311 ( .A(n7633), .ZN(n7172) );
  INV_X1 U8312 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9297) );
  INV_X1 U8313 ( .A(n6532), .ZN(n6577) );
  NAND2_X1 U8314 ( .A1(n6577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6578) );
  XNOR2_X1 U8315 ( .A(n7783), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n7776) );
  INV_X1 U8316 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U8317 ( .A1(n6579), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6580) );
  XNOR2_X1 U8318 ( .A(n6580), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8164) );
  INV_X1 U8319 ( .A(n8164), .ZN(n7193) );
  NAND2_X1 U8320 ( .A1(n6581), .A2(n7193), .ZN(n6582) );
  INV_X1 U8321 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8156) );
  XNOR2_X1 U8322 ( .A(n8147), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n8149) );
  NAND2_X1 U8323 ( .A1(n6583), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8324 ( .A1(n6594), .A2(n6584), .ZN(n6588) );
  OR2_X1 U8325 ( .A1(n6594), .A2(n6584), .ZN(n6585) );
  INV_X1 U8326 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8957) );
  INV_X1 U8327 ( .A(n6587), .ZN(n8988) );
  NAND2_X1 U8328 ( .A1(n6588), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6589) );
  XNOR2_X1 U8329 ( .A(n6589), .B(P2_IR_REG_12__SCAN_IN), .ZN(n8984) );
  XNOR2_X1 U8330 ( .A(n8984), .B(P2_REG2_REG_12__SCAN_IN), .ZN(n8987) );
  INV_X1 U8331 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U8332 ( .A1(n6592), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6593) );
  NAND2_X1 U8333 ( .A1(n6594), .A2(n6593), .ZN(n6597) );
  XNOR2_X1 U8334 ( .A(n6597), .B(n6595), .ZN(n6866) );
  INV_X1 U8335 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U8336 ( .A1(n6598), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6601) );
  XNOR2_X1 U8337 ( .A(n6601), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6876) );
  XNOR2_X1 U8338 ( .A(n6876), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9012) );
  INV_X1 U8339 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U8340 ( .A1(n6601), .A2(n6600), .ZN(n6602) );
  NAND2_X1 U8341 ( .A1(n6602), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6603) );
  XNOR2_X1 U8342 ( .A(n6603), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6887) );
  INV_X1 U8343 ( .A(n6887), .ZN(n9038) );
  NAND2_X1 U8344 ( .A1(n6604), .A2(n9038), .ZN(n9048) );
  XNOR2_X1 U8345 ( .A(n9058), .B(n9250), .ZN(n9049) );
  NAND2_X1 U8346 ( .A1(n6609), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6607) );
  XNOR2_X1 U8347 ( .A(n6607), .B(P2_IR_REG_17__SCAN_IN), .ZN(n6905) );
  INV_X1 U8348 ( .A(n6905), .ZN(n9080) );
  INV_X1 U8349 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9240) );
  AOI21_X1 U8350 ( .B1(n6611), .B2(n6610), .A(n6726), .ZN(n6614) );
  INV_X1 U8351 ( .A(n6614), .ZN(n6613) );
  INV_X1 U8352 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6612) );
  NAND2_X1 U8353 ( .A1(n6614), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n6615) );
  AND2_X1 U8354 ( .A1(n6619), .A2(n6615), .ZN(n7654) );
  INV_X1 U8355 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9224) );
  OR2_X1 U8356 ( .A1(n7654), .A2(n9224), .ZN(n6617) );
  NAND2_X1 U8357 ( .A1(n7654), .A2(n9224), .ZN(n6616) );
  NAND2_X1 U8358 ( .A1(n6617), .A2(n6616), .ZN(n6695) );
  INV_X1 U8359 ( .A(n6617), .ZN(n6618) );
  XNOR2_X1 U8360 ( .A(n6620), .B(P2_REG2_REG_19__SCAN_IN), .ZN(n6672) );
  XNOR2_X1 U8361 ( .A(n6621), .B(n6672), .ZN(n6624) );
  OR2_X1 U8362 ( .A1(n6622), .A2(P2_U3151), .ZN(n9483) );
  NOR2_X1 U8363 ( .A1(n6677), .A2(n9483), .ZN(n7254) );
  NAND2_X1 U8364 ( .A1(n6624), .A2(n9043), .ZN(n6687) );
  INV_X1 U8365 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8693) );
  INV_X1 U8366 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8780) );
  NAND2_X1 U8367 ( .A1(n6553), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6625) );
  INV_X1 U8368 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7502) );
  INV_X1 U8369 ( .A(n6625), .ZN(n6626) );
  XNOR2_X1 U8370 ( .A(n7253), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n7246) );
  INV_X1 U8371 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6629) );
  XNOR2_X1 U8372 ( .A(n7286), .B(n6629), .ZN(n7274) );
  AOI21_X1 U8373 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n7178), .A(n7277), .ZN(
        n6630) );
  XNOR2_X1 U8374 ( .A(n7175), .B(P2_REG1_REG_6__SCAN_IN), .ZN(n8946) );
  INV_X1 U8375 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7627) );
  XNOR2_X1 U8376 ( .A(n7783), .B(P2_REG1_REG_8__SCAN_IN), .ZN(n7785) );
  INV_X1 U8377 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n7958) );
  NAND2_X1 U8378 ( .A1(n7784), .A2(n5154), .ZN(n6633) );
  NAND2_X1 U8379 ( .A1(n6633), .A2(n7193), .ZN(n6634) );
  INV_X1 U8380 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8160) );
  INV_X1 U8381 ( .A(n6634), .ZN(n8142) );
  XNOR2_X1 U8382 ( .A(n8147), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n8141) );
  INV_X1 U8383 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8961) );
  INV_X1 U8384 ( .A(n6636), .ZN(n8978) );
  XNOR2_X1 U8385 ( .A(n8984), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n8977) );
  INV_X1 U8386 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6859) );
  NAND2_X1 U8387 ( .A1(n6590), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6637) );
  INV_X1 U8388 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n9003) );
  NAND2_X1 U8389 ( .A1(n9023), .A2(n9021), .ZN(n6638) );
  XNOR2_X1 U8390 ( .A(n6876), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n9020) );
  INV_X1 U8391 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8698) );
  OR2_X1 U8392 ( .A1(n6876), .A2(n8698), .ZN(n6639) );
  INV_X1 U8393 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9353) );
  NAND2_X1 U8394 ( .A1(n9058), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6641) );
  INV_X1 U8395 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9347) );
  OR2_X1 U8396 ( .A1(n7654), .A2(n9347), .ZN(n6645) );
  NAND2_X1 U8397 ( .A1(n7654), .A2(n9347), .ZN(n6643) );
  AND2_X1 U8398 ( .A1(n6645), .A2(n6643), .ZN(n6689) );
  NAND2_X1 U8399 ( .A1(n6693), .A2(n6645), .ZN(n6646) );
  XNOR2_X1 U8400 ( .A(n6620), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6673) );
  XNOR2_X1 U8401 ( .A(n6646), .B(n6673), .ZN(n6686) );
  INV_X4 U8402 ( .A(n7043), .ZN(n9487) );
  NAND2_X1 U8403 ( .A1(n7254), .A2(n9487), .ZN(n9060) );
  MUX2_X1 U8404 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n9487), .Z(n6652) );
  MUX2_X1 U8405 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n9487), .Z(n6651) );
  MUX2_X1 U8406 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n9487), .Z(n6650) );
  MUX2_X1 U8407 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n9487), .Z(n6649) );
  MUX2_X1 U8408 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n9487), .Z(n6648) );
  AOI21_X1 U8409 ( .B1(n6647), .B2(n7230), .A(n7221), .ZN(n7239) );
  XNOR2_X1 U8410 ( .A(n6648), .B(n7253), .ZN(n7238) );
  AOI21_X1 U8411 ( .B1(n6648), .B2(n7253), .A(n7237), .ZN(n7207) );
  XNOR2_X1 U8412 ( .A(n6649), .B(n6767), .ZN(n7206) );
  OAI21_X1 U8413 ( .B1(n6649), .B2(n4920), .A(n7205), .ZN(n7282) );
  XOR2_X1 U8414 ( .A(n7286), .B(n6650), .Z(n7283) );
  XOR2_X1 U8415 ( .A(n7316), .B(n6651), .Z(n7308) );
  INV_X1 U8416 ( .A(n7175), .ZN(n8944) );
  XNOR2_X1 U8417 ( .A(n6652), .B(n8944), .ZN(n8938) );
  MUX2_X1 U8418 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n9487), .Z(n6653) );
  XNOR2_X1 U8419 ( .A(n6653), .B(n7633), .ZN(n7634) );
  INV_X1 U8420 ( .A(n6653), .ZN(n6654) );
  MUX2_X1 U8421 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n9487), .Z(n6655) );
  XOR2_X1 U8422 ( .A(n7783), .B(n6655), .Z(n7774) );
  INV_X1 U8423 ( .A(n7783), .ZN(n7184) );
  MUX2_X1 U8424 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n9487), .Z(n6656) );
  XNOR2_X1 U8425 ( .A(n6656), .B(n8164), .ZN(n8165) );
  INV_X1 U8426 ( .A(n6656), .ZN(n6657) );
  MUX2_X1 U8427 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n9487), .Z(n6658) );
  XOR2_X1 U8428 ( .A(n8147), .B(n6658), .Z(n8137) );
  INV_X1 U8429 ( .A(n8147), .ZN(n7200) );
  MUX2_X1 U8430 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n9487), .Z(n6659) );
  XNOR2_X1 U8431 ( .A(n6659), .B(n8965), .ZN(n8966) );
  INV_X1 U8432 ( .A(n6659), .ZN(n6660) );
  MUX2_X1 U8433 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n9487), .Z(n6661) );
  XOR2_X1 U8434 ( .A(n6661), .B(n8984), .Z(n8973) );
  MUX2_X1 U8435 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n9487), .Z(n6662) );
  XNOR2_X1 U8436 ( .A(n6866), .B(n6662), .ZN(n8998) );
  INV_X1 U8437 ( .A(n6662), .ZN(n6663) );
  MUX2_X1 U8438 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n9487), .Z(n6664) );
  XOR2_X1 U8439 ( .A(n6664), .B(n6876), .Z(n9015) );
  INV_X1 U8440 ( .A(n6876), .ZN(n9019) );
  MUX2_X1 U8441 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n9487), .Z(n6665) );
  XNOR2_X1 U8442 ( .A(n6887), .B(n6665), .ZN(n9034) );
  INV_X1 U8443 ( .A(n6665), .ZN(n6666) );
  MUX2_X1 U8444 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n9487), .Z(n6667) );
  XNOR2_X1 U8445 ( .A(n9058), .B(n6667), .ZN(n9054) );
  OAI22_X1 U8446 ( .A1(n9055), .A2(n9054), .B1(n6667), .B2(n9058), .ZN(n9073)
         );
  MUX2_X1 U8447 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n9487), .Z(n6668) );
  XNOR2_X1 U8448 ( .A(n6905), .B(n6668), .ZN(n9074) );
  INV_X1 U8449 ( .A(n6668), .ZN(n6669) );
  MUX2_X1 U8450 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n9487), .Z(n6670) );
  NOR2_X1 U8451 ( .A1(n6671), .A2(n6670), .ZN(n6701) );
  NAND2_X1 U8452 ( .A1(n6671), .A2(n6670), .ZN(n6700) );
  OAI21_X1 U8453 ( .B1(n6701), .B2(n7654), .A(n6700), .ZN(n6675) );
  MUX2_X1 U8454 ( .A(n6673), .B(n6672), .S(n7043), .Z(n6674) );
  XNOR2_X1 U8455 ( .A(n6675), .B(n6674), .ZN(n6683) );
  NAND2_X1 U8456 ( .A1(P2_U3893), .A2(n6622), .ZN(n9075) );
  INV_X1 U8457 ( .A(n6676), .ZN(n6678) );
  AND2_X1 U8458 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8826) );
  NOR2_X1 U8459 ( .A1(n6677), .A2(n9487), .ZN(n6679) );
  INV_X1 U8460 ( .A(n6622), .ZN(n8584) );
  MUX2_X1 U8461 ( .A(n6679), .B(n6678), .S(n8584), .Z(n6680) );
  NOR2_X1 U8462 ( .A1(n9081), .A2(n4302), .ZN(n6681) );
  AOI211_X1 U8463 ( .C1(P2_ADDR_REG_19__SCAN_IN), .C2(n9077), .A(n8826), .B(
        n6681), .ZN(n6682) );
  OAI21_X1 U8464 ( .B1(n6683), .B2(n9075), .A(n6682), .ZN(n6684) );
  INV_X1 U8465 ( .A(n6689), .ZN(n6690) );
  NAND3_X1 U8466 ( .A1(n6688), .A2(n6691), .A3(n6690), .ZN(n6692) );
  INV_X1 U8467 ( .A(n6694), .ZN(n6698) );
  NAND3_X1 U8468 ( .A1(n9069), .A2(n6696), .A3(n6695), .ZN(n6697) );
  AOI21_X1 U8469 ( .B1(n6698), .B2(n6697), .A(n9086), .ZN(n6699) );
  INV_X1 U8470 ( .A(n6699), .ZN(n6705) );
  INV_X1 U8471 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10314) );
  NAND2_X1 U8472 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8894) );
  OAI21_X1 U8473 ( .B1(n8976), .B2(n10314), .A(n8894), .ZN(n6702) );
  INV_X1 U8474 ( .A(n6702), .ZN(n6703) );
  NAND4_X1 U8475 ( .A1(n6706), .A2(n6705), .A3(n6704), .A4(n6703), .ZN(
        P2_U3200) );
  INV_X1 U8476 ( .A(n6789), .ZN(n6710) );
  INV_X1 U8477 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6718) );
  OR2_X2 U8478 ( .A1(n6940), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6950) );
  INV_X1 U8479 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6720) );
  NAND2_X1 U8480 ( .A1(n6961), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U8481 ( .A1(n6977), .A2(n6722), .ZN(n9163) );
  NAND2_X1 U8482 ( .A1(n9163), .A2(n7033), .ZN(n6734) );
  INV_X1 U8483 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9328) );
  INV_X1 U8484 ( .A(n4298), .ZN(n7035) );
  NAND2_X1 U8485 ( .A1(n7035), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6731) );
  NAND2_X2 U8486 ( .A1(n8820), .A2(n9479), .ZN(n8218) );
  NAND2_X1 U8487 ( .A1(n7044), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6730) );
  OAI211_X1 U8488 ( .C1(n6993), .C2(n9328), .A(n6731), .B(n6730), .ZN(n6732)
         );
  INV_X1 U8489 ( .A(n6732), .ZN(n6733) );
  INV_X2 U8490 ( .A(n6756), .ZN(n6785) );
  NAND2_X1 U8491 ( .A1(n8307), .A2(n7010), .ZN(n6737) );
  OR2_X1 U8492 ( .A1(n4657), .A2(n8722), .ZN(n6736) );
  INV_X1 U8493 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U8494 ( .A1(n6760), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6739) );
  INV_X1 U8495 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7951) );
  OR2_X1 U8496 ( .A1(n6788), .A2(n8780), .ZN(n6745) );
  INV_X1 U8497 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7257) );
  INV_X1 U8498 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8499 ( .A1(n4893), .A2(SI_0_), .ZN(n6747) );
  XNOR2_X1 U8500 ( .A(n6747), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9497) );
  MUX2_X1 U8501 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9497), .S(n7050), .Z(n7447) );
  NAND2_X1 U8502 ( .A1(n4627), .A2(n7447), .ZN(n7492) );
  AND2_X2 U8503 ( .A1(n7491), .A2(n7492), .ZN(n7494) );
  NAND2_X1 U8504 ( .A1(n4300), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6753) );
  INV_X1 U8505 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6748) );
  OR2_X1 U8506 ( .A1(n6773), .A2(n6748), .ZN(n6752) );
  INV_X1 U8507 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7881) );
  OR2_X1 U8508 ( .A1(n4298), .A2(n7881), .ZN(n6751) );
  INV_X1 U8509 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6749) );
  OR2_X1 U8510 ( .A1(n8218), .A2(n6749), .ZN(n6750) );
  NAND4_X2 U8511 ( .A1(n6753), .A2(n6752), .A3(n6751), .A4(n6750), .ZN(n8934)
         );
  OR2_X1 U8512 ( .A1(n8531), .A2(n8678), .ZN(n6755) );
  OR2_X1 U8513 ( .A1(n7050), .A2(n7253), .ZN(n6754) );
  NAND2_X1 U8514 ( .A1(n8934), .A2(n7409), .ZN(n6757) );
  NAND2_X1 U8515 ( .A1(n7494), .A2(n6757), .ZN(n6759) );
  NOR2_X1 U8516 ( .A1(n4637), .A2(n7499), .ZN(n7410) );
  INV_X1 U8517 ( .A(n7409), .ZN(n8422) );
  AOI22_X1 U8518 ( .A1(n7410), .A2(n6757), .B1(n7369), .B2(n8422), .ZN(n6758)
         );
  NAND2_X1 U8519 ( .A1(n6759), .A2(n6758), .ZN(n7909) );
  INV_X1 U8520 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7914) );
  OR2_X1 U8521 ( .A1(n6773), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6764) );
  NAND2_X1 U8522 ( .A1(n4301), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6763) );
  INV_X1 U8523 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6761) );
  AND2_X1 U8524 ( .A1(n6764), .A2(n5158), .ZN(n6765) );
  INV_X1 U8525 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n7182) );
  NAND2_X1 U8526 ( .A1(n7151), .A2(n6785), .ZN(n6769) );
  OAI211_X1 U8527 ( .C1(n8531), .C2(n7182), .A(n6769), .B(n6768), .ZN(n9379)
         );
  NAND2_X1 U8528 ( .A1(n8933), .A2(n9379), .ZN(n6770) );
  NAND2_X1 U8529 ( .A1(n7909), .A2(n6770), .ZN(n7571) );
  OR2_X1 U8530 ( .A1(n8933), .A2(n9379), .ZN(n7570) );
  NAND2_X1 U8531 ( .A1(n4300), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8532 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n6772) );
  AND2_X1 U8533 ( .A1(n6789), .A2(n6772), .ZN(n7382) );
  OR2_X1 U8534 ( .A1(n6773), .A2(n7382), .ZN(n6776) );
  INV_X1 U8535 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6774) );
  OR2_X1 U8536 ( .A1(n8218), .A2(n6774), .ZN(n6775) );
  NAND2_X1 U8537 ( .A1(n7146), .A2(n6785), .ZN(n6780) );
  AOI22_X1 U8538 ( .A1(n6928), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6929), .B2(
        n7286), .ZN(n6779) );
  INV_X1 U8539 ( .A(n7574), .ZN(n7836) );
  AND2_X1 U8540 ( .A1(n7570), .A2(n6781), .ZN(n6784) );
  INV_X1 U8541 ( .A(n6781), .ZN(n6782) );
  OR2_X1 U8542 ( .A1(n7911), .A2(n7574), .ZN(n8428) );
  NAND2_X1 U8543 ( .A1(n7168), .A2(n6785), .ZN(n6787) );
  INV_X2 U8544 ( .A(n8531), .ZN(n6928) );
  AOI22_X1 U8545 ( .A1(n6928), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6929), .B2(
        n7316), .ZN(n6786) );
  NAND2_X1 U8546 ( .A1(n6787), .A2(n6786), .ZN(n7904) );
  NAND2_X1 U8547 ( .A1(n7044), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6794) );
  INV_X1 U8548 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7594) );
  OR2_X1 U8549 ( .A1(n6788), .A2(n7594), .ZN(n6793) );
  NAND2_X1 U8550 ( .A1(n6789), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6790) );
  AND2_X1 U8551 ( .A1(n6800), .A2(n6790), .ZN(n7429) );
  OR2_X1 U8552 ( .A1(n6773), .A2(n7429), .ZN(n6792) );
  INV_X1 U8553 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7902) );
  OR2_X1 U8554 ( .A1(n4298), .A2(n7902), .ZN(n6791) );
  NOR2_X1 U8555 ( .A1(n7904), .A2(n8932), .ZN(n6796) );
  NAND2_X1 U8556 ( .A1(n7904), .A2(n8932), .ZN(n6795) );
  NAND2_X1 U8557 ( .A1(n7159), .A2(n6785), .ZN(n6798) );
  AOI22_X1 U8558 ( .A1(n6928), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6929), .B2(
        n8944), .ZN(n6797) );
  NAND2_X1 U8559 ( .A1(n6798), .A2(n6797), .ZN(n9371) );
  NAND2_X1 U8560 ( .A1(n7044), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6805) );
  INV_X1 U8561 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6799) );
  OR2_X1 U8562 ( .A1(n6993), .A2(n6799), .ZN(n6804) );
  NAND2_X1 U8563 ( .A1(n6800), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6801) );
  AND2_X1 U8564 ( .A1(n6810), .A2(n6801), .ZN(n7559) );
  OR2_X1 U8565 ( .A1(n4625), .A2(n7559), .ZN(n6803) );
  INV_X1 U8566 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7927) );
  OR2_X1 U8567 ( .A1(n4298), .A2(n7927), .ZN(n6802) );
  OR2_X1 U8568 ( .A1(n9371), .A2(n7588), .ZN(n8430) );
  NAND2_X1 U8569 ( .A1(n9371), .A2(n7588), .ZN(n8431) );
  NAND2_X1 U8570 ( .A1(n8430), .A2(n8431), .ZN(n7921) );
  NAND2_X1 U8571 ( .A1(n7923), .A2(n7921), .ZN(n6807) );
  INV_X1 U8572 ( .A(n7588), .ZN(n9293) );
  NAND2_X1 U8573 ( .A1(n9371), .A2(n9293), .ZN(n6806) );
  AND2_X2 U8574 ( .A1(n6807), .A2(n6806), .ZN(n9289) );
  NAND2_X1 U8575 ( .A1(n7161), .A2(n6785), .ZN(n6809) );
  AOI22_X1 U8576 ( .A1(n6928), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6929), .B2(
        n7633), .ZN(n6808) );
  NAND2_X1 U8577 ( .A1(n6809), .A2(n6808), .ZN(n9364) );
  NAND2_X1 U8578 ( .A1(n7044), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n6815) );
  OR2_X1 U8579 ( .A1(n6993), .A2(n7627), .ZN(n6814) );
  NAND2_X1 U8580 ( .A1(n6810), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6811) );
  AND2_X1 U8581 ( .A1(n6818), .A2(n6811), .ZN(n7800) );
  OR2_X1 U8582 ( .A1(n4625), .A2(n7800), .ZN(n6813) );
  OR2_X1 U8583 ( .A1(n4298), .A2(n9297), .ZN(n6812) );
  OR2_X1 U8584 ( .A1(n9364), .A2(n7968), .ZN(n7828) );
  NAND2_X1 U8585 ( .A1(n9364), .A2(n7968), .ZN(n8449) );
  NAND2_X1 U8586 ( .A1(n7163), .A2(n7010), .ZN(n6817) );
  AOI22_X1 U8587 ( .A1(n6928), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6929), .B2(
        n7783), .ZN(n6816) );
  NAND2_X1 U8588 ( .A1(n7044), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6823) );
  OR2_X1 U8589 ( .A1(n6993), .A2(n7958), .ZN(n6822) );
  NAND2_X1 U8590 ( .A1(n6818), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6819) );
  AND2_X1 U8591 ( .A1(n6827), .A2(n6819), .ZN(n7964) );
  OR2_X1 U8592 ( .A1(n4625), .A2(n7964), .ZN(n6821) );
  OR2_X1 U8593 ( .A1(n4298), .A2(n8709), .ZN(n6820) );
  NAND2_X1 U8594 ( .A1(n8433), .A2(n8450), .ZN(n8555) );
  INV_X1 U8595 ( .A(n8555), .ZN(n7824) );
  OR2_X1 U8596 ( .A1(n8004), .A2(n9291), .ZN(n8012) );
  INV_X1 U8597 ( .A(n7968), .ZN(n8931) );
  OR2_X1 U8598 ( .A1(n9364), .A2(n8931), .ZN(n7823) );
  OR2_X1 U8599 ( .A1(n7824), .A2(n7823), .ZN(n7820) );
  AND2_X1 U8600 ( .A1(n8012), .A2(n7820), .ZN(n6824) );
  NAND2_X1 U8601 ( .A1(n7189), .A2(n7010), .ZN(n6826) );
  AOI22_X1 U8602 ( .A1(n6928), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6929), .B2(
        n8164), .ZN(n6825) );
  NAND2_X1 U8603 ( .A1(n6826), .A2(n6825), .ZN(n8063) );
  NAND2_X1 U8604 ( .A1(n7044), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6832) );
  OR2_X1 U8605 ( .A1(n6993), .A2(n8160), .ZN(n6831) );
  NAND2_X1 U8606 ( .A1(n6827), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6828) );
  AND2_X1 U8607 ( .A1(n6835), .A2(n6828), .ZN(n8056) );
  OR2_X1 U8608 ( .A1(n6773), .A2(n8056), .ZN(n6830) );
  OR2_X1 U8609 ( .A1(n4298), .A2(n8156), .ZN(n6829) );
  NAND2_X1 U8610 ( .A1(n8063), .A2(n8103), .ZN(n8451) );
  NAND2_X1 U8611 ( .A1(n8434), .A2(n8451), .ZN(n8556) );
  NAND2_X1 U8612 ( .A1(n7199), .A2(n7010), .ZN(n6834) );
  AOI22_X1 U8613 ( .A1(n6928), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6929), .B2(
        n8147), .ZN(n6833) );
  NAND2_X1 U8614 ( .A1(n6834), .A2(n6833), .ZN(n8175) );
  NAND2_X1 U8615 ( .A1(n7044), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6840) );
  OR2_X1 U8616 ( .A1(n6993), .A2(n8693), .ZN(n6839) );
  NAND2_X1 U8617 ( .A1(n6835), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6836) );
  AND2_X1 U8618 ( .A1(n6848), .A2(n6836), .ZN(n8101) );
  OR2_X1 U8619 ( .A1(n6773), .A2(n8101), .ZN(n6838) );
  OR2_X1 U8620 ( .A1(n4298), .A2(n8172), .ZN(n6837) );
  NAND4_X1 U8621 ( .A1(n6840), .A2(n6839), .A3(n6838), .A4(n6837), .ZN(n8929)
         );
  NAND2_X1 U8622 ( .A1(n8175), .A2(n8929), .ZN(n8040) );
  AND2_X1 U8623 ( .A1(n8556), .A2(n8040), .ZN(n6841) );
  OR2_X1 U8624 ( .A1(n8175), .A2(n8929), .ZN(n8041) );
  INV_X1 U8625 ( .A(n8040), .ZN(n6842) );
  INV_X1 U8626 ( .A(n8103), .ZN(n8930) );
  OR2_X1 U8627 ( .A1(n8063), .A2(n8930), .ZN(n8044) );
  AND2_X1 U8628 ( .A1(n8041), .A2(n6843), .ZN(n6844) );
  NAND2_X1 U8629 ( .A1(n7231), .A2(n7010), .ZN(n6847) );
  AOI22_X1 U8630 ( .A1(n6928), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6929), .B2(
        n8965), .ZN(n6846) );
  NAND2_X1 U8631 ( .A1(n6848), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6849) );
  AND2_X1 U8632 ( .A1(n6857), .A2(n6849), .ZN(n8208) );
  OR2_X1 U8633 ( .A1(n4625), .A2(n8208), .ZN(n6853) );
  NAND2_X1 U8634 ( .A1(n7044), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6852) );
  OR2_X1 U8635 ( .A1(n6993), .A2(n8961), .ZN(n6851) );
  OR2_X1 U8636 ( .A1(n4298), .A2(n8957), .ZN(n6850) );
  NAND4_X1 U8637 ( .A1(n6853), .A2(n6852), .A3(n6851), .A4(n6850), .ZN(n9276)
         );
  NAND2_X1 U8638 ( .A1(n8210), .A2(n9276), .ZN(n6854) );
  NAND2_X1 U8639 ( .A1(n7262), .A2(n6785), .ZN(n6856) );
  AOI22_X1 U8640 ( .A1(n8984), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8641 ( .A1(n6857), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6858) );
  NAND2_X1 U8642 ( .A1(n6869), .A2(n6858), .ZN(n9280) );
  NAND2_X1 U8643 ( .A1(n7033), .A2(n9280), .ZN(n6864) );
  OR2_X1 U8644 ( .A1(n6993), .A2(n6859), .ZN(n6863) );
  OR2_X1 U8645 ( .A1(n4298), .A2(n9279), .ZN(n6862) );
  INV_X1 U8646 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6860) );
  OR2_X1 U8647 ( .A1(n8218), .A2(n6860), .ZN(n6861) );
  NAND4_X1 U8648 ( .A1(n6864), .A2(n6863), .A3(n6862), .A4(n6861), .ZN(n8928)
         );
  AND2_X1 U8649 ( .A1(n7068), .A2(n8928), .ZN(n6865) );
  NAND2_X1 U8650 ( .A1(n7267), .A2(n7010), .ZN(n6868) );
  AOI22_X1 U8651 ( .A1(n6928), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6866), .B2(
        n6929), .ZN(n6867) );
  NAND2_X1 U8652 ( .A1(n6869), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6870) );
  NAND2_X1 U8653 ( .A1(n6882), .A2(n6870), .ZN(n8300) );
  NAND2_X1 U8654 ( .A1(n7033), .A2(n8300), .ZN(n6874) );
  INV_X1 U8655 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n8310) );
  OR2_X1 U8656 ( .A1(n8218), .A2(n8310), .ZN(n6873) );
  OR2_X1 U8657 ( .A1(n6993), .A2(n9003), .ZN(n6872) );
  OR2_X1 U8658 ( .A1(n4298), .A2(n8997), .ZN(n6871) );
  NAND4_X1 U8659 ( .A1(n6874), .A2(n6873), .A3(n6872), .A4(n6871), .ZN(n9277)
         );
  NOR2_X1 U8660 ( .A1(n8410), .A2(n9277), .ZN(n8411) );
  NAND2_X1 U8661 ( .A1(n8410), .A2(n9277), .ZN(n8469) );
  NAND2_X1 U8662 ( .A1(n6875), .A2(n7010), .ZN(n6878) );
  AOI22_X1 U8663 ( .A1(n6876), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6877) );
  INV_X1 U8664 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8353) );
  OR2_X1 U8665 ( .A1(n6993), .A2(n8698), .ZN(n6881) );
  OR2_X1 U8666 ( .A1(n4298), .A2(n6879), .ZN(n6880) );
  AND2_X1 U8667 ( .A1(n6881), .A2(n6880), .ZN(n6885) );
  NAND2_X1 U8668 ( .A1(n6882), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6883) );
  NAND2_X1 U8669 ( .A1(n6890), .A2(n6883), .ZN(n9270) );
  NAND2_X1 U8670 ( .A1(n9270), .A2(n7033), .ZN(n6884) );
  OAI211_X1 U8671 ( .C1(n8218), .C2(n8353), .A(n6885), .B(n6884), .ZN(n9257)
         );
  AND2_X1 U8672 ( .A1(n8357), .A2(n9257), .ZN(n6886) );
  NAND2_X1 U8673 ( .A1(n7420), .A2(n7010), .ZN(n6889) );
  AOI22_X1 U8674 ( .A1(n6887), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6888) );
  INV_X1 U8675 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U8676 ( .A1(n6890), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U8677 ( .A1(n6898), .A2(n6891), .ZN(n9261) );
  NAND2_X1 U8678 ( .A1(n9261), .A2(n7033), .ZN(n6893) );
  AOI22_X1 U8679 ( .A1(n7044), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n4301), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n6892) );
  NAND2_X1 U8680 ( .A1(n9464), .A2(n9247), .ZN(n6894) );
  NAND2_X1 U8681 ( .A1(n7517), .A2(n7010), .ZN(n6897) );
  AOI22_X1 U8682 ( .A1(n6895), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U8683 ( .A1(n6898), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8684 ( .A1(n6907), .A2(n6899), .ZN(n9251) );
  NAND2_X1 U8685 ( .A1(n9251), .A2(n7033), .ZN(n6902) );
  AOI22_X1 U8686 ( .A1(n7044), .A2(P2_REG0_REG_16__SCAN_IN), .B1(n4301), .B2(
        P2_REG1_REG_16__SCAN_IN), .ZN(n6901) );
  NAND2_X1 U8687 ( .A1(n7035), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6900) );
  NAND2_X1 U8688 ( .A1(n9457), .A2(n9235), .ZN(n8479) );
  NAND2_X1 U8689 ( .A1(n8478), .A2(n8479), .ZN(n8565) );
  NAND2_X1 U8690 ( .A1(n9457), .A2(n9258), .ZN(n6903) );
  NAND2_X1 U8691 ( .A1(n6904), .A2(n6903), .ZN(n9229) );
  AOI22_X1 U8692 ( .A1(n6905), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U8693 ( .A1(n6907), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6908) );
  NAND2_X1 U8694 ( .A1(n6919), .A2(n6908), .ZN(n9237) );
  NAND2_X1 U8695 ( .A1(n9237), .A2(n7033), .ZN(n6913) );
  NAND2_X1 U8696 ( .A1(n7044), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6910) );
  NAND2_X1 U8697 ( .A1(n4300), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6909) );
  OAI211_X1 U8698 ( .C1(n9240), .C2(n4298), .A(n6910), .B(n6909), .ZN(n6911)
         );
  INV_X1 U8699 ( .A(n6911), .ZN(n6912) );
  OR2_X1 U8700 ( .A1(n9350), .A2(n9220), .ZN(n8484) );
  NAND2_X1 U8701 ( .A1(n9350), .A2(n9220), .ZN(n8483) );
  NAND2_X1 U8702 ( .A1(n8484), .A2(n8483), .ZN(n9230) );
  NAND2_X1 U8703 ( .A1(n9229), .A2(n9230), .ZN(n6915) );
  NAND2_X1 U8704 ( .A1(n9350), .A2(n9248), .ZN(n6914) );
  AOI22_X1 U8705 ( .A1(n7654), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6917) );
  NAND2_X1 U8706 ( .A1(n6919), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6920) );
  NAND2_X1 U8707 ( .A1(n6932), .A2(n6920), .ZN(n9222) );
  NAND2_X1 U8708 ( .A1(n9222), .A2(n7033), .ZN(n6925) );
  NAND2_X1 U8709 ( .A1(n4300), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6922) );
  NAND2_X1 U8710 ( .A1(n7044), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6921) );
  OAI211_X1 U8711 ( .C1(n9224), .C2(n4298), .A(n6922), .B(n6921), .ZN(n6923)
         );
  INV_X1 U8712 ( .A(n6923), .ZN(n6924) );
  AND2_X1 U8713 ( .A1(n9346), .A2(n9208), .ZN(n6927) );
  OR2_X1 U8714 ( .A1(n9346), .A2(n9208), .ZN(n6926) );
  AOI22_X1 U8715 ( .A1(n6620), .A2(n6929), .B1(n6928), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6930) );
  NAND2_X1 U8716 ( .A1(n6932), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U8717 ( .A1(n6940), .A2(n6933), .ZN(n9212) );
  INV_X1 U8718 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U8719 ( .A1(n4301), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6935) );
  NAND2_X1 U8720 ( .A1(n7044), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6934) );
  OAI211_X1 U8721 ( .C1(n4298), .C2(n9211), .A(n6935), .B(n6934), .ZN(n6936)
         );
  NAND2_X1 U8722 ( .A1(n9443), .A2(n9221), .ZN(n8491) );
  INV_X1 U8723 ( .A(n9443), .ZN(n6937) );
  NAND2_X1 U8724 ( .A1(n8097), .A2(n7010), .ZN(n6939) );
  OR2_X1 U8725 ( .A1(n4657), .A2(n8098), .ZN(n6938) );
  NAND2_X1 U8726 ( .A1(n6940), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6941) );
  NAND2_X1 U8727 ( .A1(n6950), .A2(n6941), .ZN(n9199) );
  NAND2_X1 U8728 ( .A1(n9199), .A2(n7033), .ZN(n6947) );
  INV_X1 U8729 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n6944) );
  NAND2_X1 U8730 ( .A1(n7044), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8731 ( .A1(n4301), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6942) );
  OAI211_X1 U8732 ( .C1(n6944), .C2(n4298), .A(n6943), .B(n6942), .ZN(n6945)
         );
  INV_X1 U8733 ( .A(n6945), .ZN(n6946) );
  NAND2_X1 U8734 ( .A1(n9339), .A2(n8829), .ZN(n8492) );
  OR2_X1 U8735 ( .A1(n9339), .A2(n9209), .ZN(n9168) );
  NAND2_X1 U8736 ( .A1(n8213), .A2(n7010), .ZN(n6949) );
  OR2_X1 U8737 ( .A1(n4657), .A2(n8214), .ZN(n6948) );
  NAND2_X2 U8738 ( .A1(n6949), .A2(n6948), .ZN(n8606) );
  NAND2_X1 U8739 ( .A1(n6950), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6951) );
  NAND2_X1 U8740 ( .A1(n6959), .A2(n6951), .ZN(n9188) );
  NAND2_X1 U8741 ( .A1(n9188), .A2(n7033), .ZN(n6956) );
  INV_X1 U8742 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U8743 ( .A1(n7044), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6953) );
  NAND2_X1 U8744 ( .A1(n4301), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n6952) );
  OAI211_X1 U8745 ( .C1(n9187), .C2(n4298), .A(n6953), .B(n6952), .ZN(n6954)
         );
  INV_X1 U8746 ( .A(n6954), .ZN(n6955) );
  OR2_X1 U8747 ( .A1(n8606), .A2(n9172), .ZN(n6968) );
  NAND2_X1 U8748 ( .A1(n8286), .A2(n6785), .ZN(n6958) );
  OR2_X1 U8749 ( .A1(n4657), .A2(n8289), .ZN(n6957) );
  NAND2_X2 U8750 ( .A1(n6958), .A2(n6957), .ZN(n9427) );
  NAND2_X1 U8751 ( .A1(n6959), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6960) );
  NAND2_X1 U8752 ( .A1(n6961), .A2(n6960), .ZN(n9176) );
  NAND2_X1 U8753 ( .A1(n9176), .A2(n7033), .ZN(n6967) );
  INV_X1 U8754 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6964) );
  NAND2_X1 U8755 ( .A1(n7044), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6963) );
  NAND2_X1 U8756 ( .A1(n4300), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6962) );
  OAI211_X1 U8757 ( .C1(n6964), .C2(n4298), .A(n6963), .B(n6962), .ZN(n6965)
         );
  INV_X1 U8758 ( .A(n6965), .ZN(n6966) );
  NAND2_X1 U8759 ( .A1(n9427), .A2(n9158), .ZN(n8497) );
  NAND2_X1 U8760 ( .A1(n8498), .A2(n8497), .ZN(n9177) );
  NAND2_X1 U8761 ( .A1(n8606), .A2(n9194), .ZN(n8496) );
  NAND2_X1 U8762 ( .A1(n8494), .A2(n8496), .ZN(n9183) );
  INV_X1 U8763 ( .A(n6968), .ZN(n9169) );
  OR2_X1 U8764 ( .A1(n9183), .A2(n9169), .ZN(n6969) );
  AND2_X1 U8765 ( .A1(n9177), .A2(n6969), .ZN(n6971) );
  NOR2_X1 U8766 ( .A1(n9427), .A2(n9185), .ZN(n6970) );
  INV_X1 U8767 ( .A(n9421), .ZN(n8659) );
  NAND2_X1 U8768 ( .A1(n6973), .A2(n6785), .ZN(n6975) );
  OR2_X1 U8769 ( .A1(n4657), .A2(n8382), .ZN(n6974) );
  INV_X1 U8770 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6976) );
  NAND2_X1 U8771 ( .A1(n6977), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6978) );
  NAND2_X1 U8772 ( .A1(n6989), .A2(n6978), .ZN(n9149) );
  NAND2_X1 U8773 ( .A1(n9149), .A2(n7033), .ZN(n6983) );
  INV_X1 U8774 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9325) );
  NAND2_X1 U8775 ( .A1(n7035), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8776 ( .A1(n7044), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6979) );
  OAI211_X1 U8777 ( .C1(n6993), .C2(n9325), .A(n6980), .B(n6979), .ZN(n6981)
         );
  INV_X1 U8778 ( .A(n6981), .ZN(n6982) );
  NAND2_X1 U8779 ( .A1(n9415), .A2(n9159), .ZN(n8506) );
  NAND2_X1 U8780 ( .A1(n8505), .A2(n8506), .ZN(n8545) );
  AOI21_X2 U8781 ( .B1(n9144), .B2(n8545), .A(n6984), .ZN(n9132) );
  NAND2_X1 U8782 ( .A1(n9493), .A2(n7010), .ZN(n6986) );
  OR2_X1 U8783 ( .A1(n4657), .A2(n9495), .ZN(n6985) );
  INV_X1 U8784 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6987) );
  NAND2_X1 U8785 ( .A1(n6989), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6990) );
  NAND2_X1 U8786 ( .A1(n7000), .A2(n6990), .ZN(n9138) );
  NAND2_X1 U8787 ( .A1(n9138), .A2(n7033), .ZN(n6996) );
  INV_X1 U8788 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U8789 ( .A1(n7044), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U8790 ( .A1(n7035), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6991) );
  OAI211_X1 U8791 ( .C1(n6993), .C2(n9322), .A(n6992), .B(n6991), .ZN(n6994)
         );
  INV_X1 U8792 ( .A(n6994), .ZN(n6995) );
  NAND2_X1 U8793 ( .A1(n9409), .A2(n9145), .ZN(n6997) );
  INV_X1 U8794 ( .A(n9409), .ZN(n9131) );
  NAND2_X1 U8795 ( .A1(n9489), .A2(n6785), .ZN(n6999) );
  OR2_X1 U8796 ( .A1(n4657), .A2(n9491), .ZN(n6998) );
  NAND2_X1 U8797 ( .A1(n7000), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n7001) );
  NAND2_X1 U8798 ( .A1(n7014), .A2(n7001), .ZN(n9127) );
  NAND2_X1 U8799 ( .A1(n9127), .A2(n7033), .ZN(n7006) );
  INV_X1 U8800 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n9126) );
  NAND2_X1 U8801 ( .A1(n7044), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n7003) );
  NAND2_X1 U8802 ( .A1(n4301), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n7002) );
  OAI211_X1 U8803 ( .C1(n9126), .C2(n4298), .A(n7003), .B(n7002), .ZN(n7004)
         );
  INV_X1 U8804 ( .A(n7004), .ZN(n7005) );
  NAND2_X2 U8805 ( .A1(n7006), .A2(n7005), .ZN(n9133) );
  NAND2_X1 U8806 ( .A1(n9123), .A2(n7007), .ZN(n7009) );
  INV_X1 U8807 ( .A(n9403), .ZN(n7008) );
  NAND2_X1 U8808 ( .A1(n8383), .A2(n7010), .ZN(n7012) );
  OR2_X1 U8809 ( .A1(n4657), .A2(n9486), .ZN(n7011) );
  INV_X1 U8810 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7013) );
  NAND2_X1 U8811 ( .A1(n7014), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U8812 ( .A1(n9110), .A2(n7033), .ZN(n7020) );
  INV_X1 U8813 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9114) );
  NAND2_X1 U8814 ( .A1(n4300), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n7017) );
  NAND2_X1 U8815 ( .A1(n7044), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n7016) );
  OAI211_X1 U8816 ( .C1(n4298), .C2(n9114), .A(n7017), .B(n7016), .ZN(n7018)
         );
  INV_X1 U8817 ( .A(n7018), .ZN(n7019) );
  NAND2_X1 U8818 ( .A1(n7021), .A2(n6785), .ZN(n7023) );
  OR2_X1 U8819 ( .A1(n4657), .A2(n9485), .ZN(n7022) );
  NAND2_X1 U8820 ( .A1(n7024), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U8821 ( .A1(n8807), .A2(n7025), .ZN(n9098) );
  NAND2_X1 U8822 ( .A1(n9098), .A2(n7033), .ZN(n7030) );
  INV_X1 U8823 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n9097) );
  NAND2_X1 U8824 ( .A1(n7044), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n7027) );
  NAND2_X1 U8825 ( .A1(n4301), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n7026) );
  OAI211_X1 U8826 ( .C1(n9097), .C2(n4298), .A(n7027), .B(n7026), .ZN(n7028)
         );
  INV_X1 U8827 ( .A(n7028), .ZN(n7029) );
  OR2_X1 U8828 ( .A1(n9391), .A2(n9105), .ZN(n8525) );
  NAND2_X1 U8829 ( .A1(n8386), .A2(n6785), .ZN(n7032) );
  INV_X1 U8830 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9478) );
  OR2_X1 U8831 ( .A1(n4657), .A2(n9478), .ZN(n7031) );
  NAND2_X1 U8832 ( .A1(n7032), .A2(n7031), .ZN(n7106) );
  INV_X1 U8833 ( .A(n8807), .ZN(n7034) );
  NAND2_X1 U8834 ( .A1(n7034), .A2(n7033), .ZN(n8224) );
  INV_X1 U8835 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U8836 ( .A1(n4300), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n7037) );
  NAND2_X1 U8837 ( .A1(n7035), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n7036) );
  OAI211_X1 U8838 ( .C1(n8777), .C2(n8218), .A(n7037), .B(n7036), .ZN(n7038)
         );
  INV_X1 U8839 ( .A(n7038), .ZN(n7039) );
  NAND2_X1 U8840 ( .A1(n7106), .A2(n8926), .ZN(n8408) );
  NAND2_X1 U8841 ( .A1(n6620), .A2(n4743), .ZN(n7112) );
  NAND2_X1 U8842 ( .A1(n7040), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7041) );
  NAND2_X1 U8843 ( .A1(n8542), .A2(n8581), .ZN(n7042) );
  NAND2_X2 U8844 ( .A1(n7112), .A2(n7042), .ZN(n9295) );
  NAND2_X1 U8845 ( .A1(n4619), .A2(n9295), .ZN(n7057) );
  XNOR2_X1 U8846 ( .A(n8584), .B(n7043), .ZN(n7347) );
  INV_X1 U8847 ( .A(n7347), .ZN(n7346) );
  AND2_X2 U8848 ( .A1(n8515), .A2(n7346), .ZN(n9292) );
  INV_X1 U8849 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8850 ( .A1(n7044), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7046) );
  NAND2_X1 U8851 ( .A1(n4301), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7045) );
  OAI211_X1 U8852 ( .C1(n7047), .C2(n4298), .A(n7046), .B(n7045), .ZN(n7048)
         );
  INV_X1 U8853 ( .A(n7048), .ZN(n7049) );
  AND2_X1 U8854 ( .A1(n8224), .A2(n7049), .ZN(n8409) );
  NAND2_X1 U8855 ( .A1(n7050), .A2(P2_B_REG_SCAN_IN), .ZN(n7051) );
  NAND2_X1 U8856 ( .A1(n9290), .A2(n7051), .ZN(n8802) );
  NOR2_X1 U8857 ( .A1(n8409), .A2(n8802), .ZN(n7054) );
  INV_X1 U8858 ( .A(n9391), .ZN(n8526) );
  INV_X1 U8859 ( .A(n9105), .ZN(n7052) );
  INV_X1 U8860 ( .A(n9295), .ZN(n9231) );
  NOR4_X1 U8861 ( .A1(n8570), .A2(n8526), .A3(n7052), .A4(n9231), .ZN(n7053)
         );
  AOI211_X1 U8862 ( .C1(n9292), .C2(n9105), .A(n7054), .B(n7053), .ZN(n7056)
         );
  NAND2_X1 U8863 ( .A1(n9391), .A2(n9105), .ZN(n8519) );
  NAND2_X1 U8864 ( .A1(n7058), .A2(n5153), .ZN(n7055) );
  OAI211_X1 U8865 ( .C1(n7058), .C2(n7057), .A(n7056), .B(n7055), .ZN(n8812)
         );
  OR2_X1 U8866 ( .A1(n8934), .A2(n8422), .ZN(n8420) );
  NAND2_X1 U8867 ( .A1(n7060), .A2(n8420), .ZN(n7568) );
  NAND2_X1 U8868 ( .A1(n8933), .A2(n7484), .ZN(n8427) );
  INV_X1 U8869 ( .A(n8439), .ZN(n7062) );
  OAI21_X1 U8870 ( .B1(n7062), .B2(n8421), .A(n8428), .ZN(n7063) );
  INV_X1 U8871 ( .A(n7063), .ZN(n7064) );
  INV_X1 U8872 ( .A(n8932), .ZN(n7552) );
  NAND2_X1 U8873 ( .A1(n7904), .A2(n7552), .ZN(n7919) );
  AND2_X1 U8874 ( .A1(n8431), .A2(n7919), .ZN(n8444) );
  NAND2_X1 U8875 ( .A1(n7065), .A2(n8430), .ZN(n9302) );
  AND2_X1 U8876 ( .A1(n8433), .A2(n7828), .ZN(n8448) );
  INV_X1 U8877 ( .A(n8929), .ZN(n8079) );
  OR2_X1 U8878 ( .A1(n8175), .A2(n8079), .ZN(n8456) );
  AND2_X1 U8879 ( .A1(n8434), .A2(n8456), .ZN(n8446) );
  NAND2_X1 U8880 ( .A1(n8039), .A2(n8446), .ZN(n7067) );
  NAND2_X1 U8881 ( .A1(n8175), .A2(n8079), .ZN(n8457) );
  NAND2_X1 U8882 ( .A1(n7067), .A2(n8457), .ZN(n8032) );
  INV_X1 U8883 ( .A(n9276), .ZN(n8202) );
  NAND2_X1 U8884 ( .A1(n8210), .A2(n8202), .ZN(n8462) );
  NAND2_X1 U8885 ( .A1(n7068), .A2(n8293), .ZN(n8463) );
  NAND2_X1 U8886 ( .A1(n8460), .A2(n8463), .ZN(n9283) );
  NAND2_X1 U8887 ( .A1(n9281), .A2(n8460), .ZN(n8275) );
  INV_X1 U8888 ( .A(n9277), .ZN(n8086) );
  NAND2_X1 U8889 ( .A1(n8410), .A2(n8086), .ZN(n7069) );
  OR2_X1 U8890 ( .A1(n8410), .A2(n8086), .ZN(n7070) );
  INV_X1 U8891 ( .A(n9257), .ZN(n8593) );
  NOR2_X1 U8892 ( .A1(n8357), .A2(n8593), .ZN(n8471) );
  INV_X1 U8893 ( .A(n8471), .ZN(n7071) );
  NAND2_X1 U8894 ( .A1(n8357), .A2(n8593), .ZN(n8472) );
  INV_X1 U8895 ( .A(n9247), .ZN(n8334) );
  OR2_X1 U8896 ( .A1(n9464), .A2(n8334), .ZN(n8475) );
  INV_X1 U8897 ( .A(n8478), .ZN(n7072) );
  INV_X1 U8898 ( .A(n9230), .ZN(n8481) );
  INV_X1 U8899 ( .A(n8483), .ZN(n7073) );
  NAND2_X1 U8900 ( .A1(n9346), .A2(n9233), .ZN(n8546) );
  INV_X1 U8901 ( .A(n8491), .ZN(n8489) );
  OAI211_X1 U8902 ( .C1(n8489), .C2(n9195), .A(n8493), .B(n9196), .ZN(n7074)
         );
  INV_X1 U8903 ( .A(n7074), .ZN(n7075) );
  INV_X1 U8904 ( .A(n8496), .ZN(n7076) );
  NAND2_X1 U8905 ( .A1(n9421), .A2(n8886), .ZN(n9150) );
  AND2_X1 U8906 ( .A1(n8506), .A2(n9150), .ZN(n8501) );
  INV_X1 U8907 ( .A(n8505), .ZN(n7077) );
  NOR2_X1 U8908 ( .A1(n9403), .A2(n8628), .ZN(n8514) );
  NAND2_X1 U8909 ( .A1(n9403), .A2(n8628), .ZN(n8517) );
  NAND2_X1 U8910 ( .A1(n9116), .A2(n9124), .ZN(n8520) );
  NAND2_X1 U8911 ( .A1(n8542), .A2(n8099), .ZN(n7833) );
  NAND2_X1 U8912 ( .A1(n7833), .A2(n8415), .ZN(n7079) );
  NAND2_X1 U8913 ( .A1(n7344), .A2(n7080), .ZN(n8050) );
  INV_X1 U8914 ( .A(n7080), .ZN(n7081) );
  OR2_X1 U8915 ( .A1(n7081), .A2(n8099), .ZN(n7082) );
  NAND2_X1 U8916 ( .A1(n7082), .A2(n4756), .ZN(n7090) );
  XNOR2_X1 U8917 ( .A(n7083), .B(P2_B_REG_SCAN_IN), .ZN(n7084) );
  INV_X1 U8918 ( .A(n9492), .ZN(n7086) );
  NAND2_X1 U8919 ( .A1(n7085), .A2(n9492), .ZN(n7087) );
  NOR2_X1 U8920 ( .A1(n8008), .A2(n8542), .ZN(n7091) );
  NAND2_X1 U8921 ( .A1(n9492), .A2(n7083), .ZN(n7147) );
  NAND2_X1 U8922 ( .A1(n7090), .A2(n7328), .ZN(n7443) );
  OAI21_X1 U8923 ( .B1(n7444), .B2(n7091), .A(n7443), .ZN(n7105) );
  NAND2_X1 U8924 ( .A1(n7329), .A2(n8515), .ZN(n7335) );
  NOR2_X1 U8925 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .ZN(
        n8687) );
  NOR4_X1 U8926 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n7094) );
  NOR4_X1 U8927 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_27__SCAN_IN), .ZN(n7093) );
  NOR4_X1 U8928 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n7092) );
  NAND4_X1 U8929 ( .A1(n8687), .A2(n7094), .A3(n7093), .A4(n7092), .ZN(n7100)
         );
  NOR4_X1 U8930 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n7098) );
  NOR4_X1 U8931 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n7097) );
  NOR4_X1 U8932 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n7096) );
  NOR4_X1 U8933 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_20__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_10__SCAN_IN), .ZN(n7095) );
  NAND4_X1 U8934 ( .A1(n7098), .A2(n7097), .A3(n7096), .A4(n7095), .ZN(n7099)
         );
  NOR2_X1 U8935 ( .A1(n7100), .A2(n7099), .ZN(n7101) );
  AND2_X1 U8936 ( .A1(n7350), .A2(n7115), .ZN(n7102) );
  NAND2_X1 U8937 ( .A1(n7335), .A2(n7102), .ZN(n7442) );
  INV_X1 U8938 ( .A(n9472), .ZN(n7103) );
  NOR2_X1 U8939 ( .A1(n7442), .A2(n7116), .ZN(n7104) );
  OR2_X1 U8940 ( .A1(n7119), .A2(n9307), .ZN(n7109) );
  INV_X1 U8941 ( .A(n7106), .ZN(n8813) );
  NAND2_X1 U8942 ( .A1(n7109), .A2(n7108), .ZN(P2_U3488) );
  INV_X1 U8943 ( .A(n7328), .ZN(n7110) );
  NAND2_X1 U8944 ( .A1(n7110), .A2(n9472), .ZN(n7440) );
  INV_X1 U8945 ( .A(n7115), .ZN(n7111) );
  NOR2_X1 U8946 ( .A1(n7440), .A2(n7111), .ZN(n7331) );
  OR2_X1 U8947 ( .A1(n8542), .A2(n8099), .ZN(n7327) );
  NAND2_X1 U8948 ( .A1(n7344), .A2(n7338), .ZN(n7113) );
  NAND2_X1 U8949 ( .A1(n7349), .A2(n7113), .ZN(n7118) );
  NOR2_X1 U8950 ( .A1(n8515), .A2(n9378), .ZN(n7114) );
  NAND2_X1 U8951 ( .A1(n7338), .A2(n7114), .ZN(n7322) );
  NAND2_X1 U8952 ( .A1(n8534), .A2(n9378), .ZN(n9265) );
  NAND2_X1 U8953 ( .A1(n7322), .A2(n9265), .ZN(n7333) );
  NAND2_X1 U8954 ( .A1(n7116), .A2(n7115), .ZN(n7341) );
  INV_X1 U8955 ( .A(n7350), .ZN(n9471) );
  NAND2_X1 U8956 ( .A1(n7333), .A2(n7345), .ZN(n7117) );
  OR2_X1 U8957 ( .A1(n7119), .A2(n10301), .ZN(n7123) );
  INV_X1 U8958 ( .A(n9378), .ZN(n9368) );
  NOR2_X1 U8959 ( .A1(n10298), .A2(n8777), .ZN(n7120) );
  NAND2_X1 U8960 ( .A1(n7123), .A2(n7122), .ZN(P2_U3456) );
  XNOR2_X1 U8961 ( .A(n7128), .B(n7124), .ZN(n7129) );
  NAND2_X1 U8962 ( .A1(n7129), .A2(n9966), .ZN(n7132) );
  INV_X1 U8963 ( .A(n7130), .ZN(n7131) );
  NAND2_X1 U8964 ( .A1(n7132), .A2(n7131), .ZN(n9757) );
  AOI21_X1 U8965 ( .B1(n7140), .B2(n9762), .A(n9952), .ZN(n7134) );
  AND2_X1 U8966 ( .A1(n7135), .A2(n7134), .ZN(n9752) );
  NOR2_X1 U8967 ( .A1(n7136), .A2(n7611), .ZN(n7138) );
  INV_X1 U8968 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7142) );
  NOR2_X1 U8969 ( .A1(n7143), .A2(P1_U3086), .ZN(n7145) );
  NOR2_X1 U8970 ( .A1(n4893), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10122) );
  INV_X1 U8971 ( .A(n7146), .ZN(n7179) );
  OAI222_X1 U8972 ( .A1(P1_U3086), .A2(n7527), .B1(n10134), .B2(n7179), .C1(
        n10128), .C2(n5217), .ZN(P1_U3351) );
  INV_X1 U8973 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n7150) );
  INV_X1 U8974 ( .A(n7147), .ZN(n7148) );
  AOI22_X1 U8975 ( .A1(n7165), .A2(n7150), .B1(n7149), .B2(n7148), .ZN(
        P2_U3376) );
  INV_X1 U8976 ( .A(n7151), .ZN(n7181) );
  OAI222_X1 U8977 ( .A1(n10128), .A2(n7152), .B1(n10134), .B2(n7181), .C1(
        P1_U3086), .C2(n9693), .ZN(P1_U3352) );
  INV_X1 U8978 ( .A(n7153), .ZN(n7157) );
  OAI222_X1 U8979 ( .A1(n7155), .A2(P1_U3086), .B1(n10134), .B2(n7157), .C1(
        n7154), .C2(n10128), .ZN(P1_U3354) );
  AND2_X1 U8980 ( .A1(n7165), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8981 ( .A1(n7165), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8982 ( .A1(n7165), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8983 ( .A1(n7165), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8984 ( .A1(n7165), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8985 ( .A1(n7165), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8986 ( .A1(n7165), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8987 ( .A1(n7165), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8988 ( .A1(n7165), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8989 ( .A1(n7165), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8990 ( .A1(n7165), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8991 ( .A1(n7165), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8992 ( .A1(n7165), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8993 ( .A1(n7165), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8994 ( .A1(n7165), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8995 ( .A1(n7165), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8996 ( .A1(n7165), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8997 ( .A1(n7165), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8998 ( .A1(n7165), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8999 ( .A1(n7165), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U9000 ( .A1(n7165), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U9001 ( .A1(n7165), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U9002 ( .A1(n7165), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U9003 ( .A1(n7165), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U9004 ( .A1(n7165), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  NAND2_X1 U9005 ( .A1(n6735), .A2(P2_U3151), .ZN(n9490) );
  NAND2_X1 U9006 ( .A1(n4893), .A2(P2_U3151), .ZN(n9496) );
  INV_X1 U9007 ( .A(n9496), .ZN(n9482) );
  INV_X1 U9008 ( .A(n9482), .ZN(n9481) );
  OAI222_X1 U9009 ( .A1(n9490), .A2(n7158), .B1(n9481), .B2(n7157), .C1(
        P2_U3151), .C2(n7230), .ZN(P2_U3294) );
  INV_X1 U9010 ( .A(n7159), .ZN(n7176) );
  INV_X1 U9011 ( .A(n10128), .ZN(n7656) );
  AOI22_X1 U9012 ( .A1(n7647), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n7656), .ZN(n7160) );
  OAI21_X1 U9013 ( .B1(n7176), .B2(n10134), .A(n7160), .ZN(P1_U3349) );
  INV_X1 U9014 ( .A(n7161), .ZN(n7173) );
  AOI22_X1 U9015 ( .A1(n7676), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n7656), .ZN(n7162) );
  OAI21_X1 U9016 ( .B1(n7173), .B2(n10134), .A(n7162), .ZN(P1_U3348) );
  INV_X1 U9017 ( .A(n7163), .ZN(n7185) );
  AOI22_X1 U9018 ( .A1(n7665), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7656), .ZN(n7164) );
  OAI21_X1 U9019 ( .B1(n7185), .B2(n10134), .A(n7164), .ZN(P1_U3347) );
  INV_X1 U9020 ( .A(n7165), .ZN(n7166) );
  INV_X1 U9021 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n8749) );
  NOR2_X1 U9022 ( .A1(n7166), .A2(n8749), .ZN(P2_U3251) );
  INV_X1 U9023 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n8745) );
  NOR2_X1 U9024 ( .A1(n7166), .A2(n8745), .ZN(P2_U3244) );
  INV_X1 U9025 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n8702) );
  NOR2_X1 U9026 ( .A1(n7166), .A2(n8702), .ZN(P2_U3252) );
  INV_X1 U9027 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n8787) );
  NOR2_X1 U9028 ( .A1(n7166), .A2(n8787), .ZN(P2_U3258) );
  INV_X1 U9029 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n8723) );
  NOR2_X1 U9030 ( .A1(n7166), .A2(n8723), .ZN(P2_U3253) );
  OAI222_X1 U9031 ( .A1(n10128), .A2(n7167), .B1(n10134), .B2(n7183), .C1(
        P1_U3086), .C2(n7538), .ZN(P1_U3353) );
  INV_X1 U9032 ( .A(n7168), .ZN(n7188) );
  OAI222_X1 U9033 ( .A1(n10128), .A2(n7170), .B1(n10134), .B2(n7188), .C1(
        n7169), .C2(P1_U3086), .ZN(P1_U3350) );
  NAND2_X1 U9034 ( .A1(n7911), .A2(P2_U3893), .ZN(n7171) );
  OAI21_X1 U9035 ( .B1(P2_U3893), .B2(n5217), .A(n7171), .ZN(P2_U3495) );
  INV_X1 U9036 ( .A(n9490), .ZN(n7653) );
  INV_X1 U9037 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7174) );
  OAI222_X1 U9038 ( .A1(n9494), .A2(n7174), .B1(n9496), .B2(n7173), .C1(
        P2_U3151), .C2(n7172), .ZN(P2_U3288) );
  INV_X1 U9039 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7177) );
  OAI222_X1 U9040 ( .A1(n9494), .A2(n7177), .B1(n9496), .B2(n7176), .C1(
        P2_U3151), .C2(n7175), .ZN(P2_U3289) );
  OAI222_X1 U9041 ( .A1(n9494), .A2(n7180), .B1(n9496), .B2(n7179), .C1(
        P2_U3151), .C2(n7178), .ZN(P2_U3291) );
  OAI222_X1 U9042 ( .A1(n9494), .A2(n7182), .B1(n9496), .B2(n7181), .C1(
        P2_U3151), .C2(n4920), .ZN(P2_U3292) );
  OAI222_X1 U9043 ( .A1(n9494), .A2(n8678), .B1(n9496), .B2(n7183), .C1(
        P2_U3151), .C2(n7253), .ZN(P2_U3293) );
  INV_X1 U9044 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n7186) );
  OAI222_X1 U9045 ( .A1(n9494), .A2(n7186), .B1(n9496), .B2(n7185), .C1(
        P2_U3151), .C2(n7184), .ZN(P2_U3287) );
  OAI222_X1 U9046 ( .A1(n9481), .A2(n7188), .B1(n4444), .B2(P2_U3151), .C1(
        n7187), .C2(n9494), .ZN(P2_U3290) );
  INV_X1 U9047 ( .A(n7189), .ZN(n7192) );
  INV_X1 U9048 ( .A(n7190), .ZN(n7512) );
  OAI222_X1 U9049 ( .A1(n10128), .A2(n7191), .B1(n10134), .B2(n7192), .C1(
        n7512), .C2(P1_U3086), .ZN(P1_U3346) );
  OAI222_X1 U9050 ( .A1(n9494), .A2(n7194), .B1(n7193), .B2(P2_U3151), .C1(
        n9481), .C2(n7192), .ZN(P2_U3286) );
  INV_X1 U9051 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n7196) );
  NAND2_X1 U9052 ( .A1(P1_U3973), .A2(n9724), .ZN(n7195) );
  OAI21_X1 U9053 ( .B1(P1_U3973), .B2(n7196), .A(n7195), .ZN(P1_U3585) );
  INV_X1 U9054 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7198) );
  NAND2_X1 U9055 ( .A1(P1_U3973), .A2(n7401), .ZN(n7197) );
  OAI21_X1 U9056 ( .B1(P1_U3973), .B2(n7198), .A(n7197), .ZN(P1_U3554) );
  NOR2_X1 U9057 ( .A1(n10141), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U9058 ( .A(n7199), .ZN(n7203) );
  OAI222_X1 U9059 ( .A1(n9494), .A2(n7201), .B1(n7200), .B2(P2_U3151), .C1(
        n9481), .C2(n7203), .ZN(P2_U3285) );
  INV_X1 U9060 ( .A(n7202), .ZN(n7816) );
  OAI222_X1 U9061 ( .A1(P1_U3086), .A2(n7816), .B1(n10128), .B2(n7204), .C1(
        n10134), .C2(n7203), .ZN(P1_U3345) );
  OAI21_X1 U9062 ( .B1(n7207), .B2(n7206), .A(n7205), .ZN(n7208) );
  NAND2_X1 U9063 ( .A1(n7208), .A2(n9066), .ZN(n7216) );
  OAI21_X1 U9064 ( .B1(P2_REG1_REG_3__SCAN_IN), .B2(n7209), .A(n7275), .ZN(
        n7210) );
  AOI22_X1 U9065 ( .A1(n7210), .A2(n6685), .B1(n9077), .B2(
        P2_ADDR_REG_3__SCAN_IN), .ZN(n7214) );
  NAND2_X1 U9066 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n7482) );
  OAI21_X1 U9067 ( .B1(P2_REG2_REG_3__SCAN_IN), .B2(n7211), .A(n7272), .ZN(
        n7212) );
  NAND2_X1 U9068 ( .A1(n7212), .A2(n9043), .ZN(n7213) );
  AND3_X1 U9069 ( .A1(n7214), .A2(n7482), .A3(n7213), .ZN(n7215) );
  OAI211_X1 U9070 ( .C1(n9081), .C2(n4920), .A(n7216), .B(n7215), .ZN(P2_U3185) );
  AOI21_X1 U9071 ( .B1(n7219), .B2(n7218), .A(n7217), .ZN(n7220) );
  OAI22_X1 U9072 ( .A1(n9086), .A2(n7220), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7951), .ZN(n7228) );
  AOI211_X1 U9073 ( .C1(n7222), .C2(n7255), .A(n9075), .B(n7221), .ZN(n7227)
         );
  AOI21_X1 U9074 ( .B1(n7502), .B2(n7224), .A(n7223), .ZN(n7225) );
  OAI22_X1 U9075 ( .A1(n8976), .A2(n10306), .B1(n9060), .B2(n7225), .ZN(n7226)
         );
  NOR3_X1 U9076 ( .A1(n7228), .A2(n7227), .A3(n7226), .ZN(n7229) );
  OAI21_X1 U9077 ( .B1(n7230), .B2(n9081), .A(n7229), .ZN(P2_U3183) );
  INV_X1 U9078 ( .A(n7231), .ZN(n7235) );
  OAI222_X1 U9079 ( .A1(n9494), .A2(n7233), .B1(n9496), .B2(n7235), .C1(
        P2_U3151), .C2(n7232), .ZN(P2_U3284) );
  INV_X1 U9080 ( .A(n7234), .ZN(n8028) );
  OAI222_X1 U9081 ( .A1(n10128), .A2(n7236), .B1(n10134), .B2(n7235), .C1(
        P1_U3086), .C2(n8028), .ZN(P1_U3344) );
  AOI211_X1 U9082 ( .C1(n7239), .C2(n7238), .A(n9075), .B(n7237), .ZN(n7251)
         );
  AOI21_X1 U9083 ( .B1(n7242), .B2(n7241), .A(n7240), .ZN(n7243) );
  OAI22_X1 U9084 ( .A1(n9086), .A2(n7243), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6748), .ZN(n7250) );
  INV_X1 U9085 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7248) );
  AOI21_X1 U9086 ( .B1(n7246), .B2(n7245), .A(n7244), .ZN(n7247) );
  OAI22_X1 U9087 ( .A1(n8976), .A2(n7248), .B1(n9060), .B2(n7247), .ZN(n7249)
         );
  NOR3_X1 U9088 ( .A1(n7251), .A2(n7250), .A3(n7249), .ZN(n7252) );
  OAI21_X1 U9089 ( .B1(n7253), .B2(n9081), .A(n7252), .ZN(P2_U3184) );
  NOR2_X1 U9090 ( .A1(n7254), .A2(n9066), .ZN(n7259) );
  AOI21_X1 U9091 ( .B1(n7256), .B2(n4959), .A(n7255), .ZN(n7258) );
  OAI22_X1 U9092 ( .A1(n7259), .A2(n7258), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7257), .ZN(n7260) );
  AOI21_X1 U9093 ( .B1(n9077), .B2(P2_ADDR_REG_0__SCAN_IN), .A(n7260), .ZN(
        n7261) );
  OAI21_X1 U9094 ( .B1(n4959), .B2(n9081), .A(n7261), .ZN(P2_U3182) );
  INV_X1 U9095 ( .A(n7262), .ZN(n7265) );
  INV_X1 U9096 ( .A(n7263), .ZN(n8188) );
  OAI222_X1 U9097 ( .A1(n10128), .A2(n7264), .B1(n10134), .B2(n7265), .C1(
        n8188), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U9098 ( .A1(n9494), .A2(n7266), .B1(n6590), .B2(P2_U3151), .C1(
        n9481), .C2(n7265), .ZN(P2_U3283) );
  INV_X1 U9099 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7269) );
  INV_X1 U9100 ( .A(n7267), .ZN(n7288) );
  INV_X1 U9101 ( .A(n7268), .ZN(n8346) );
  OAI222_X1 U9102 ( .A1(n10128), .A2(n7269), .B1(n10134), .B2(n7288), .C1(
        P1_U3086), .C2(n8346), .ZN(P1_U3342) );
  INV_X1 U9103 ( .A(n9081), .ZN(n8985) );
  AND3_X1 U9104 ( .A1(n7272), .A2(n7271), .A3(n4319), .ZN(n7273) );
  OAI21_X1 U9105 ( .B1(n7270), .B2(n7273), .A(n9043), .ZN(n7280) );
  AND3_X1 U9106 ( .A1(n7275), .A2(n7274), .A3(n4320), .ZN(n7276) );
  OAI21_X1 U9107 ( .B1(n7277), .B2(n7276), .A(n6685), .ZN(n7279) );
  NAND2_X1 U9108 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7379) );
  NAND2_X1 U9109 ( .A1(n9077), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7278) );
  NAND4_X1 U9110 ( .A1(n7280), .A2(n7279), .A3(n7379), .A4(n7278), .ZN(n7285)
         );
  AOI211_X1 U9111 ( .C1(n7283), .C2(n7282), .A(n9075), .B(n7281), .ZN(n7284)
         );
  AOI211_X1 U9112 ( .C1(n8985), .C2(n7286), .A(n7285), .B(n7284), .ZN(n7287)
         );
  INV_X1 U9113 ( .A(n7287), .ZN(P2_U3186) );
  INV_X1 U9114 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7289) );
  OAI222_X1 U9115 ( .A1(n9490), .A2(n7289), .B1(P2_U3151), .B2(n9002), .C1(
        n9481), .C2(n7288), .ZN(P2_U3282) );
  INV_X1 U9116 ( .A(n6875), .ZN(n7303) );
  AOI22_X1 U9117 ( .A1(n10153), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7656), .ZN(n7290) );
  OAI21_X1 U9118 ( .B1(n7303), .B2(n10134), .A(n7290), .ZN(P1_U3341) );
  OAI21_X1 U9119 ( .B1(n10250), .B2(n9966), .A(n7719), .ZN(n7293) );
  INV_X1 U9120 ( .A(n4643), .ZN(n7463) );
  OR2_X1 U9121 ( .A1(n9962), .A2(n7463), .ZN(n7720) );
  OAI21_X1 U9122 ( .B1(n7717), .B2(n7405), .A(n7720), .ZN(n7291) );
  INV_X1 U9123 ( .A(n7291), .ZN(n7292) );
  AND2_X1 U9124 ( .A1(n7293), .A2(n7292), .ZN(n10237) );
  NAND2_X1 U9125 ( .A1(n10289), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7294) );
  OAI21_X1 U9126 ( .B1(n10289), .B2(n10237), .A(n7294), .ZN(P1_U3522) );
  XNOR2_X1 U9127 ( .A(n7295), .B(n7296), .ZN(n7522) );
  INV_X1 U9128 ( .A(n7297), .ZN(n7300) );
  NOR4_X1 U9129 ( .A1(n7300), .A2(n7299), .A3(n7298), .A4(P1_U3086), .ZN(n7468) );
  INV_X1 U9130 ( .A(n7468), .ZN(n7479) );
  NAND2_X1 U9131 ( .A1(n7479), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7302) );
  AOI22_X1 U9132 ( .A1(n9652), .A2(n4643), .B1(n9659), .B2(n7725), .ZN(n7301)
         );
  OAI211_X1 U9133 ( .C1(n7522), .C2(n9662), .A(n7302), .B(n7301), .ZN(P1_U3232) );
  INV_X1 U9134 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7304) );
  OAI222_X1 U9135 ( .A1(n9490), .A2(n7304), .B1(n9481), .B2(n7303), .C1(
        P2_U3151), .C2(n9019), .ZN(P2_U3281) );
  INV_X1 U9136 ( .A(n9376), .ZN(n7830) );
  NAND2_X1 U9137 ( .A1(n7830), .A2(n9231), .ZN(n7305) );
  NAND2_X1 U9138 ( .A1(n4627), .A2(n7471), .ZN(n8414) );
  NAND2_X1 U9139 ( .A1(n8416), .A2(n8414), .ZN(n8547) );
  NOR2_X1 U9140 ( .A1(n4758), .A2(n9234), .ZN(n7449) );
  AOI21_X1 U9141 ( .B1(n7305), .B2(n8547), .A(n7449), .ZN(n7469) );
  MUX2_X1 U9142 ( .A(n7469), .B(n6742), .S(n10301), .Z(n7306) );
  OAI21_X1 U9143 ( .B1(n7471), .B2(n8805), .A(n7306), .ZN(P2_U3390) );
  AOI211_X1 U9144 ( .C1(n7309), .C2(n7308), .A(n9075), .B(n7307), .ZN(n7321)
         );
  OAI21_X1 U9145 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(n7311), .A(n7310), .ZN(
        n7315) );
  OAI21_X1 U9146 ( .B1(P2_REG2_REG_5__SCAN_IN), .B2(n7313), .A(n7312), .ZN(
        n7314) );
  AOI22_X1 U9147 ( .A1(n6685), .A2(n7315), .B1(n7314), .B2(n9043), .ZN(n7319)
         );
  NAND2_X1 U9148 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7430) );
  NAND2_X1 U9149 ( .A1(n8985), .A2(n7316), .ZN(n7318) );
  NAND2_X1 U9150 ( .A1(n9077), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7317) );
  NAND4_X1 U9151 ( .A1(n7319), .A2(n7430), .A3(n7318), .A4(n7317), .ZN(n7320)
         );
  OR2_X1 U9152 ( .A1(n7321), .A2(n7320), .ZN(P2_U3187) );
  INV_X1 U9153 ( .A(n7322), .ZN(n7323) );
  NAND2_X1 U9154 ( .A1(n7349), .A2(n7323), .ZN(n7326) );
  INV_X1 U9155 ( .A(n7338), .ZN(n7324) );
  NAND2_X1 U9156 ( .A1(n7345), .A2(n7324), .ZN(n7325) );
  XNOR2_X1 U9157 ( .A(n7360), .B(n4637), .ZN(n7359) );
  NAND2_X1 U9158 ( .A1(n7330), .A2(n8416), .ZN(n7358) );
  XOR2_X1 U9159 ( .A(n7359), .B(n7358), .Z(n7356) );
  INV_X1 U9160 ( .A(n7341), .ZN(n7339) );
  INV_X1 U9161 ( .A(n7331), .ZN(n7332) );
  NAND2_X1 U9162 ( .A1(n7333), .A2(n7332), .ZN(n7337) );
  AND3_X1 U9163 ( .A1(n7335), .A2(n7334), .A3(n8308), .ZN(n7336) );
  OAI211_X1 U9164 ( .C1(n7339), .C2(n7338), .A(n7337), .B(n7336), .ZN(n7340)
         );
  NAND2_X1 U9165 ( .A1(n7340), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7343) );
  NOR2_X1 U9166 ( .A1(n7344), .A2(n9471), .ZN(n8585) );
  NAND2_X1 U9167 ( .A1(n8585), .A2(n7341), .ZN(n7342) );
  INV_X1 U9168 ( .A(n8920), .ZN(n8655) );
  NAND2_X1 U9169 ( .A1(n8655), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7386) );
  INV_X1 U9170 ( .A(n7344), .ZN(n7448) );
  NAND2_X1 U9171 ( .A1(n7345), .A2(n7448), .ZN(n7348) );
  INV_X1 U9172 ( .A(n9265), .ZN(n8273) );
  NAND2_X1 U9173 ( .A1(n7349), .A2(n8273), .ZN(n7352) );
  NAND2_X1 U9174 ( .A1(n7350), .A2(n4742), .ZN(n7351) );
  AOI22_X1 U9175 ( .A1(n8916), .A2(n4627), .B1(n8908), .B2(n7499), .ZN(n7353)
         );
  OAI21_X1 U9176 ( .B1(n7369), .B2(n8918), .A(n7353), .ZN(n7354) );
  AOI21_X1 U9177 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n7386), .A(n7354), .ZN(
        n7355) );
  OAI21_X1 U9178 ( .B1(n8910), .B2(n7356), .A(n7355), .ZN(P2_U3162) );
  XNOR2_X1 U9179 ( .A(n8422), .B(n4297), .ZN(n7368) );
  XNOR2_X1 U9180 ( .A(n7368), .B(n7369), .ZN(n7366) );
  NAND2_X1 U9181 ( .A1(n7360), .A2(n4758), .ZN(n7361) );
  XOR2_X1 U9182 ( .A(n7367), .B(n7366), .Z(n7365) );
  AOI22_X1 U9183 ( .A1(n8916), .A2(n4637), .B1(n8908), .B2(n7409), .ZN(n7362)
         );
  OAI21_X1 U9184 ( .B1(n4624), .B2(n8918), .A(n7362), .ZN(n7363) );
  AOI21_X1 U9185 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7386), .A(n7363), .ZN(
        n7364) );
  OAI21_X1 U9186 ( .B1(n7365), .B2(n8910), .A(n7364), .ZN(P2_U3177) );
  XNOR2_X1 U9187 ( .A(n7357), .B(n7574), .ZN(n7424) );
  XNOR2_X1 U9188 ( .A(n7424), .B(n7911), .ZN(n7378) );
  INV_X1 U9189 ( .A(n7368), .ZN(n7370) );
  NAND2_X1 U9190 ( .A1(n7370), .A2(n7369), .ZN(n7371) );
  XNOR2_X1 U9191 ( .A(n7484), .B(n7357), .ZN(n7372) );
  XNOR2_X1 U9192 ( .A(n7372), .B(n8933), .ZN(n7487) );
  NAND2_X1 U9193 ( .A1(n7372), .A2(n8933), .ZN(n7373) );
  INV_X1 U9194 ( .A(n7373), .ZN(n7374) );
  NOR2_X1 U9195 ( .A1(n7378), .A2(n7374), .ZN(n7375) );
  INV_X1 U9196 ( .A(n7428), .ZN(n7376) );
  AOI21_X1 U9197 ( .B1(n7378), .B2(n7377), .A(n7376), .ZN(n7385) );
  INV_X1 U9198 ( .A(n7379), .ZN(n7381) );
  OAI22_X1 U9199 ( .A1(n7552), .A2(n8918), .B1(n8905), .B2(n4624), .ZN(n7380)
         );
  AOI211_X1 U9200 ( .C1(n7836), .C2(n8908), .A(n7381), .B(n7380), .ZN(n7384)
         );
  INV_X1 U9201 ( .A(n7382), .ZN(n7837) );
  NAND2_X1 U9202 ( .A1(n8920), .A2(n7837), .ZN(n7383) );
  OAI211_X1 U9203 ( .C1(n7385), .C2(n8910), .A(n7384), .B(n7383), .ZN(P2_U3170) );
  NAND2_X1 U9204 ( .A1(n7386), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7388) );
  AOI22_X1 U9205 ( .A1(n8912), .A2(n8547), .B1(n7447), .B2(n8908), .ZN(n7387)
         );
  OAI211_X1 U9206 ( .C1(n4758), .C2(n8918), .A(n7388), .B(n7387), .ZN(P2_U3172) );
  OAI21_X1 U9207 ( .B1(n7390), .B2(n7389), .A(n7687), .ZN(n10230) );
  INV_X1 U9208 ( .A(n10230), .ZN(n7394) );
  XNOR2_X1 U9209 ( .A(n7392), .B(n7391), .ZN(n7393) );
  AOI222_X1 U9210 ( .A1(n9966), .A2(n7393), .B1(n9680), .B2(n9934), .C1(n4643), 
        .C2(n9932), .ZN(n10233) );
  OAI211_X1 U9211 ( .C1(n7403), .C2(n10228), .A(n10015), .B(n7691), .ZN(n10223) );
  OAI211_X1 U9212 ( .C1(n10265), .C2(n7394), .A(n10233), .B(n10223), .ZN(n7418) );
  INV_X1 U9213 ( .A(n7418), .ZN(n7396) );
  INV_X1 U9214 ( .A(n10107), .ZN(n8283) );
  AOI22_X1 U9215 ( .A1(n8283), .A2(n7465), .B1(n10282), .B2(
        P1_REG0_REG_2__SCAN_IN), .ZN(n7395) );
  OAI21_X1 U9216 ( .B1(n7396), .B2(n10282), .A(n7395), .ZN(P1_U3459) );
  INV_X1 U9217 ( .A(n7397), .ZN(n7398) );
  AOI21_X1 U9218 ( .B1(n7399), .B2(n5943), .A(n7398), .ZN(n7748) );
  AOI222_X1 U9219 ( .A1(n9966), .A2(n7402), .B1(n9681), .B2(n9934), .C1(n7401), 
        .C2(n9932), .ZN(n7745) );
  INV_X1 U9220 ( .A(n7403), .ZN(n7404) );
  OAI211_X1 U9221 ( .C1(n5969), .C2(n7405), .A(n7404), .B(n10015), .ZN(n7742)
         );
  OAI211_X1 U9222 ( .C1(n10265), .C2(n7748), .A(n7745), .B(n7742), .ZN(n7438)
         );
  OAI22_X1 U9223 ( .A1(n10107), .A2(n5969), .B1(n10283), .B2(n5233), .ZN(n7406) );
  AOI21_X1 U9224 ( .B1(n10283), .B2(n7438), .A(n7406), .ZN(n7407) );
  INV_X1 U9225 ( .A(n7407), .ZN(P1_U3456) );
  INV_X1 U9226 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n7416) );
  XNOR2_X1 U9227 ( .A(n7408), .B(n8548), .ZN(n7876) );
  AND2_X1 U9228 ( .A1(n7409), .A2(n9378), .ZN(n7879) );
  NOR2_X1 U9229 ( .A1(n7494), .A2(n7410), .ZN(n7411) );
  XNOR2_X1 U9230 ( .A(n7411), .B(n8548), .ZN(n7412) );
  NAND2_X1 U9231 ( .A1(n7412), .A2(n9295), .ZN(n7414) );
  AOI22_X1 U9232 ( .A1(n9292), .A2(n4637), .B1(n8933), .B2(n9290), .ZN(n7413)
         );
  NAND2_X1 U9233 ( .A1(n7414), .A2(n7413), .ZN(n7877) );
  AOI211_X1 U9234 ( .C1(n9376), .C2(n7876), .A(n7879), .B(n7877), .ZN(n10293)
         );
  OR2_X1 U9235 ( .A1(n10293), .A2(n9307), .ZN(n7415) );
  OAI21_X1 U9236 ( .B1(n9383), .B2(n7416), .A(n7415), .ZN(P2_U3461) );
  OAI22_X1 U9237 ( .A1(n10048), .A2(n10228), .B1(n10291), .B2(n6446), .ZN(
        n7417) );
  AOI21_X1 U9238 ( .B1(n7418), .B2(n10291), .A(n7417), .ZN(n7419) );
  INV_X1 U9239 ( .A(n7419), .ZN(P1_U3524) );
  INV_X1 U9240 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n8669) );
  INV_X1 U9241 ( .A(n7420), .ZN(n7422) );
  OAI222_X1 U9242 ( .A1(n9490), .A2(n8669), .B1(n9481), .B2(n7422), .C1(
        P2_U3151), .C2(n9038), .ZN(P2_U3280) );
  INV_X1 U9243 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7423) );
  OAI222_X1 U9244 ( .A1(n10128), .A2(n7423), .B1(n10134), .B2(n7422), .C1(
        P1_U3086), .C2(n7421), .ZN(P1_U3340) );
  INV_X1 U9245 ( .A(n7424), .ZN(n7426) );
  INV_X1 U9246 ( .A(n7911), .ZN(n7425) );
  NAND2_X1 U9247 ( .A1(n7426), .A2(n7425), .ZN(n7427) );
  XNOR2_X1 U9248 ( .A(n7357), .B(n7904), .ZN(n7553) );
  XNOR2_X1 U9249 ( .A(n7553), .B(n8932), .ZN(n7550) );
  XOR2_X1 U9250 ( .A(n7551), .B(n7550), .Z(n7436) );
  INV_X1 U9251 ( .A(n7429), .ZN(n7903) );
  NAND2_X1 U9252 ( .A1(n8920), .A2(n7903), .ZN(n7433) );
  INV_X1 U9253 ( .A(n7430), .ZN(n7431) );
  AOI21_X1 U9254 ( .B1(n8916), .B2(n7911), .A(n7431), .ZN(n7432) );
  OAI211_X1 U9255 ( .C1(n7588), .C2(n8918), .A(n7433), .B(n7432), .ZN(n7434)
         );
  AOI21_X1 U9256 ( .B1(n7904), .B2(n8908), .A(n7434), .ZN(n7435) );
  OAI21_X1 U9257 ( .B1(n7436), .B2(n8910), .A(n7435), .ZN(P2_U3167) );
  OAI22_X1 U9258 ( .A1(n10048), .A2(n5969), .B1(n10291), .B2(n5234), .ZN(n7437) );
  AOI21_X1 U9259 ( .B1(n10291), .B2(n7438), .A(n7437), .ZN(n7439) );
  INV_X1 U9260 ( .A(n7439), .ZN(P1_U3523) );
  INV_X1 U9261 ( .A(n7440), .ZN(n7441) );
  NOR2_X1 U9262 ( .A1(n7442), .A2(n7441), .ZN(n7445) );
  NAND3_X1 U9263 ( .A1(n7445), .A2(n7444), .A3(n7443), .ZN(n7451) );
  INV_X1 U9264 ( .A(n7451), .ZN(n7446) );
  AOI22_X1 U9265 ( .A1(n9300), .A2(n7447), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n9299), .ZN(n7455) );
  NOR2_X1 U9266 ( .A1(n7448), .A2(n9378), .ZN(n7450) );
  AOI21_X1 U9267 ( .B1(n7450), .B2(n8547), .A(n7449), .ZN(n7452) );
  MUX2_X1 U9268 ( .A(n7453), .B(n7452), .S(n9296), .Z(n7454) );
  NAND2_X1 U9269 ( .A1(n7455), .A2(n7454), .ZN(P2_U3233) );
  INV_X1 U9270 ( .A(n7456), .ZN(n7473) );
  INV_X1 U9271 ( .A(n7457), .ZN(n7459) );
  NOR3_X1 U9272 ( .A1(n7473), .A2(n7459), .A3(n7458), .ZN(n7462) );
  INV_X1 U9273 ( .A(n7460), .ZN(n7461) );
  OAI21_X1 U9274 ( .B1(n7462), .B2(n7461), .A(n9621), .ZN(n7467) );
  OAI22_X1 U9275 ( .A1(n7463), .A2(n9654), .B1(n9643), .B2(n7604), .ZN(n7464)
         );
  AOI21_X1 U9276 ( .B1(n7465), .B2(n9659), .A(n7464), .ZN(n7466) );
  OAI211_X1 U9277 ( .C1(n7468), .C2(n10222), .A(n7467), .B(n7466), .ZN(
        P1_U3237) );
  MUX2_X1 U9278 ( .A(n8780), .B(n7469), .S(n9383), .Z(n7470) );
  OAI21_X1 U9279 ( .B1(n9310), .B2(n7471), .A(n7470), .ZN(P2_U3459) );
  AOI21_X1 U9280 ( .B1(n7474), .B2(n7472), .A(n7473), .ZN(n7481) );
  NOR2_X1 U9281 ( .A1(n9630), .A2(n5969), .ZN(n7478) );
  OAI22_X1 U9282 ( .A1(n7476), .A2(n9654), .B1(n9643), .B2(n7475), .ZN(n7477)
         );
  AOI211_X1 U9283 ( .C1(n7479), .C2(P1_REG3_REG_1__SCAN_IN), .A(n7478), .B(
        n7477), .ZN(n7480) );
  OAI21_X1 U9284 ( .B1(n7481), .B2(n9662), .A(n7480), .ZN(P1_U3222) );
  INV_X1 U9285 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7915) );
  AOI22_X1 U9286 ( .A1(n8916), .A2(n8934), .B1(n8902), .B2(n7911), .ZN(n7483)
         );
  OAI211_X1 U9287 ( .C1(n7484), .C2(n8923), .A(n7483), .B(n7482), .ZN(n7489)
         );
  AOI211_X1 U9288 ( .C1(n7487), .C2(n7486), .A(n8910), .B(n7485), .ZN(n7488)
         );
  AOI211_X1 U9289 ( .C1(n7915), .C2(n8920), .A(n7489), .B(n7488), .ZN(n7490)
         );
  INV_X1 U9290 ( .A(n7490), .ZN(P2_U3158) );
  NOR2_X1 U9291 ( .A1(n7491), .A2(n7492), .ZN(n7493) );
  OAI21_X1 U9292 ( .B1(n7494), .B2(n7493), .A(n9295), .ZN(n7496) );
  AOI22_X1 U9293 ( .A1(n9290), .A2(n8934), .B1(n4627), .B2(n9292), .ZN(n7495)
         );
  AND2_X1 U9294 ( .A1(n7496), .A2(n7495), .ZN(n7948) );
  NAND2_X1 U9295 ( .A1(n7491), .A2(n8416), .ZN(n7497) );
  AND2_X1 U9296 ( .A1(n7498), .A2(n7497), .ZN(n7949) );
  INV_X1 U9297 ( .A(n7949), .ZN(n7955) );
  NAND2_X1 U9298 ( .A1(n7955), .A2(n9376), .ZN(n7501) );
  NAND2_X1 U9299 ( .A1(n7499), .A2(n9378), .ZN(n7500) );
  AND3_X1 U9300 ( .A1(n7948), .A2(n7501), .A3(n7500), .ZN(n10292) );
  MUX2_X1 U9301 ( .A(n10292), .B(n7502), .S(n9307), .Z(n7503) );
  INV_X1 U9302 ( .A(n7503), .ZN(P2_U3460) );
  OAI21_X1 U9303 ( .B1(n7506), .B2(n7505), .A(n7504), .ZN(n7507) );
  NAND2_X1 U9304 ( .A1(n7507), .A2(n10211), .ZN(n7516) );
  OAI21_X1 U9305 ( .B1(n7510), .B2(n7509), .A(n7508), .ZN(n7514) );
  INV_X1 U9306 ( .A(n10206), .ZN(n9716) );
  NAND2_X1 U9307 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U9308 ( .A1(n10141), .A2(P1_ADDR_REG_9__SCAN_IN), .ZN(n7511) );
  OAI211_X1 U9309 ( .C1(n10215), .C2(n7512), .A(n8263), .B(n7511), .ZN(n7513)
         );
  AOI21_X1 U9310 ( .B1(n7514), .B2(n9716), .A(n7513), .ZN(n7515) );
  NAND2_X1 U9311 ( .A1(n7516), .A2(n7515), .ZN(P1_U3252) );
  INV_X1 U9312 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7519) );
  INV_X1 U9313 ( .A(n7517), .ZN(n7520) );
  INV_X1 U9314 ( .A(n7518), .ZN(n10175) );
  OAI222_X1 U9315 ( .A1(n10128), .A2(n7519), .B1(n10134), .B2(n7520), .C1(
        P1_U3086), .C2(n10175), .ZN(P1_U3339) );
  INV_X1 U9316 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7521) );
  OAI222_X1 U9317 ( .A1(n9490), .A2(n7521), .B1(n9481), .B2(n7520), .C1(
        P2_U3151), .C2(n9058), .ZN(P2_U3279) );
  MUX2_X1 U9318 ( .A(n7522), .B(n9683), .S(n5846), .Z(n7525) );
  AOI21_X1 U9319 ( .B1(n5846), .B2(n5250), .A(n4675), .ZN(n10138) );
  OAI21_X1 U9320 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10138), .A(P1_U3973), .ZN(
        n7523) );
  AOI21_X1 U9321 ( .B1(n7525), .B2(n7524), .A(n7523), .ZN(n7549) );
  AND2_X1 U9322 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n7606) );
  AOI21_X1 U9323 ( .B1(n10141), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n7606), .ZN(
        n7526) );
  OAI21_X1 U9324 ( .B1(n10215), .B2(n7527), .A(n7526), .ZN(n7536) );
  OAI21_X1 U9325 ( .B1(n7530), .B2(n7529), .A(n7528), .ZN(n7534) );
  OAI211_X1 U9326 ( .C1(n7532), .C2(n7531), .A(n10211), .B(n4737), .ZN(n7533)
         );
  OAI21_X1 U9327 ( .B1(n10206), .B2(n7534), .A(n7533), .ZN(n7535) );
  OR3_X1 U9328 ( .A1(n7549), .A2(n7536), .A3(n7535), .ZN(P1_U3247) );
  AOI22_X1 U9329 ( .A1(n10141), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n7537) );
  OAI21_X1 U9330 ( .B1(n7538), .B2(n10215), .A(n7537), .ZN(n7548) );
  OAI21_X1 U9331 ( .B1(n7541), .B2(n7540), .A(n7539), .ZN(n7546) );
  OAI211_X1 U9332 ( .C1(n7544), .C2(n7543), .A(n10211), .B(n7542), .ZN(n7545)
         );
  OAI21_X1 U9333 ( .B1(n7546), .B2(n10206), .A(n7545), .ZN(n7547) );
  OR3_X1 U9334 ( .A1(n7549), .A2(n7548), .A3(n7547), .ZN(P1_U3245) );
  NAND2_X1 U9335 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  XNOR2_X1 U9336 ( .A(n9371), .B(n7357), .ZN(n7792) );
  XNOR2_X1 U9337 ( .A(n7792), .B(n7588), .ZN(n7556) );
  AOI21_X1 U9338 ( .B1(n7555), .B2(n7556), .A(n8910), .ZN(n7558) );
  NAND2_X1 U9339 ( .A1(n7558), .A2(n7795), .ZN(n7565) );
  INV_X1 U9340 ( .A(n7559), .ZN(n7928) );
  INV_X1 U9341 ( .A(n9371), .ZN(n7560) );
  NOR2_X1 U9342 ( .A1(n8923), .A2(n7560), .ZN(n7563) );
  NAND2_X1 U9343 ( .A1(n8916), .A2(n8932), .ZN(n7561) );
  NAND2_X1 U9344 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8941) );
  OAI211_X1 U9345 ( .C1(n7968), .C2(n8918), .A(n7561), .B(n8941), .ZN(n7562)
         );
  AOI211_X1 U9346 ( .C1(n7928), .C2(n8920), .A(n7563), .B(n7562), .ZN(n7564)
         );
  NAND2_X1 U9347 ( .A1(n7565), .A2(n7564), .ZN(P2_U3179) );
  INV_X1 U9348 ( .A(n7566), .ZN(n7596) );
  AOI22_X1 U9349 ( .A1(n10185), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n7656), .ZN(n7567) );
  OAI21_X1 U9350 ( .B1(n7596), .B2(n10134), .A(n7567), .ZN(P1_U3338) );
  XNOR2_X1 U9351 ( .A(n8933), .B(n9379), .ZN(n8549) );
  INV_X1 U9352 ( .A(n8421), .ZN(n8440) );
  AOI21_X1 U9353 ( .B1(n7568), .B2(n8549), .A(n8440), .ZN(n7569) );
  XNOR2_X1 U9354 ( .A(n7569), .B(n8426), .ZN(n7843) );
  NAND2_X1 U9355 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  XNOR2_X1 U9356 ( .A(n7572), .B(n8426), .ZN(n7573) );
  AOI222_X1 U9357 ( .A1(n9295), .A2(n7573), .B1(n8933), .B2(n9292), .C1(n8932), 
        .C2(n9290), .ZN(n7840) );
  OAI21_X1 U9358 ( .B1(n7574), .B2(n9368), .A(n7840), .ZN(n7575) );
  AOI21_X1 U9359 ( .B1(n7843), .B2(n9376), .A(n7575), .ZN(n10295) );
  OR2_X1 U9360 ( .A1(n9383), .A2(n6629), .ZN(n7576) );
  OAI21_X1 U9361 ( .B1(n10295), .B2(n9307), .A(n7576), .ZN(P2_U3463) );
  NAND2_X1 U9362 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9694) );
  INV_X1 U9363 ( .A(n9694), .ZN(n7579) );
  OAI22_X1 U9364 ( .A1(n9630), .A2(n10239), .B1(n7577), .B2(n9643), .ZN(n7578)
         );
  AOI211_X1 U9365 ( .C1(n9640), .C2(n9681), .A(n7579), .B(n7578), .ZN(n7585)
         );
  OAI21_X1 U9366 ( .B1(n7582), .B2(n7581), .A(n7580), .ZN(n7583) );
  NAND2_X1 U9367 ( .A1(n7583), .A2(n9621), .ZN(n7584) );
  OAI211_X1 U9368 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9636), .A(n7585), .B(
        n7584), .ZN(P1_U3218) );
  XNOR2_X1 U9369 ( .A(n7586), .B(n4555), .ZN(n7590) );
  NAND2_X1 U9370 ( .A1(n7911), .A2(n9292), .ZN(n7587) );
  OAI21_X1 U9371 ( .B1(n7588), .B2(n9234), .A(n7587), .ZN(n7589) );
  AOI21_X1 U9372 ( .B1(n7590), .B2(n9295), .A(n7589), .ZN(n7901) );
  OR2_X1 U9373 ( .A1(n7591), .A2(n8553), .ZN(n7592) );
  NAND2_X1 U9374 ( .A1(n7920), .A2(n7592), .ZN(n7900) );
  AOI22_X1 U9375 ( .A1(n7900), .A2(n9376), .B1(n9378), .B2(n7904), .ZN(n7593)
         );
  AND2_X1 U9376 ( .A1(n7901), .A2(n7593), .ZN(n10296) );
  MUX2_X1 U9377 ( .A(n7594), .B(n10296), .S(n9383), .Z(n7595) );
  INV_X1 U9378 ( .A(n7595), .ZN(P2_U3464) );
  OAI222_X1 U9379 ( .A1(n9490), .A2(n7597), .B1(n9481), .B2(n7596), .C1(
        P2_U3151), .C2(n9080), .ZN(P2_U3278) );
  AND2_X1 U9380 ( .A1(n7580), .A2(n7601), .ZN(n7603) );
  INV_X1 U9381 ( .A(n7598), .ZN(n7599) );
  XNOR2_X1 U9382 ( .A(n7600), .B(n7599), .ZN(n7602) );
  NAND3_X1 U9383 ( .A1(n7580), .A2(n7602), .A3(n7601), .ZN(n7750) );
  OAI211_X1 U9384 ( .C1(n7603), .C2(n7602), .A(n9621), .B(n7750), .ZN(n7608)
         );
  OAI22_X1 U9385 ( .A1(n9630), .A2(n10245), .B1(n7604), .B2(n9654), .ZN(n7605)
         );
  AOI211_X1 U9386 ( .C1(n9652), .C2(n4587), .A(n7606), .B(n7605), .ZN(n7607)
         );
  OAI211_X1 U9387 ( .C1(n9636), .C2(n7706), .A(n7608), .B(n7607), .ZN(P1_U3230) );
  XNOR2_X1 U9388 ( .A(n7610), .B(n7609), .ZN(n10256) );
  NAND3_X1 U9389 ( .A1(n7613), .A2(n7612), .A3(n7611), .ZN(n7619) );
  AND2_X1 U9390 ( .A1(n10278), .A2(n9968), .ZN(n7614) );
  XNOR2_X1 U9391 ( .A(n7616), .B(n7615), .ZN(n7617) );
  AOI222_X1 U9392 ( .A1(n9966), .A2(n7617), .B1(n9678), .B2(n9934), .C1(n9679), 
        .C2(n9932), .ZN(n10255) );
  MUX2_X1 U9393 ( .A(n7618), .B(n10255), .S(n9971), .Z(n7624) );
  INV_X1 U9394 ( .A(n7711), .ZN(n7620) );
  AOI211_X1 U9395 ( .C1(n10253), .C2(n7620), .A(n9952), .B(n4934), .ZN(n10252)
         );
  OAI22_X1 U9396 ( .A1(n10227), .A2(n7757), .B1(n10221), .B2(n7762), .ZN(n7622) );
  AOI21_X1 U9397 ( .B1(n9944), .B2(n10252), .A(n7622), .ZN(n7623) );
  OAI211_X1 U9398 ( .C1(n10256), .C2(n9929), .A(n7624), .B(n7623), .ZN(
        P1_U3288) );
  AOI21_X1 U9399 ( .B1(n7627), .B2(n7626), .A(n7625), .ZN(n7639) );
  INV_X1 U9400 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7628) );
  NAND2_X1 U9401 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7801) );
  OAI21_X1 U9402 ( .B1(n8976), .B2(n7628), .A(n7801), .ZN(n7632) );
  AOI21_X1 U9403 ( .B1(n9297), .B2(n7629), .A(n7777), .ZN(n7630) );
  NOR2_X1 U9404 ( .A1(n7630), .A2(n9086), .ZN(n7631) );
  AOI211_X1 U9405 ( .C1(n8985), .C2(n7633), .A(n7632), .B(n7631), .ZN(n7638)
         );
  XNOR2_X1 U9406 ( .A(n4282), .B(n7634), .ZN(n7636) );
  NAND2_X1 U9407 ( .A1(n7636), .A2(n9066), .ZN(n7637) );
  OAI211_X1 U9408 ( .C1(n7639), .C2(n9060), .A(n7638), .B(n7637), .ZN(P2_U3189) );
  AOI211_X1 U9409 ( .C1(n7642), .C2(n7641), .A(n7640), .B(n10158), .ZN(n7652)
         );
  NOR2_X1 U9410 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  NOR3_X1 U9411 ( .A1(n10206), .A2(n7646), .A3(n7645), .ZN(n7651) );
  INV_X1 U9412 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n7649) );
  NAND2_X1 U9413 ( .A1(n10168), .A2(n7647), .ZN(n7648) );
  NAND2_X1 U9414 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7735) );
  OAI211_X1 U9415 ( .C1(n7649), .C2(n10220), .A(n7648), .B(n7735), .ZN(n7650)
         );
  OR3_X1 U9416 ( .A1(n7652), .A2(n7651), .A3(n7650), .ZN(P1_U3249) );
  INV_X1 U9417 ( .A(n6916), .ZN(n7658) );
  AOI22_X1 U9418 ( .A1(n7654), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7653), .ZN(n7655) );
  OAI21_X1 U9419 ( .B1(n7658), .B2(n9496), .A(n7655), .ZN(P2_U3277) );
  AOI22_X1 U9420 ( .A1(n10200), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7656), .ZN(n7657) );
  OAI21_X1 U9421 ( .B1(n7658), .B2(n10134), .A(n7657), .ZN(P1_U3337) );
  AOI211_X1 U9422 ( .C1(n7661), .C2(n7660), .A(n10158), .B(n7659), .ZN(n7670)
         );
  AOI211_X1 U9423 ( .C1(n7664), .C2(n7663), .A(n10206), .B(n7662), .ZN(n7669)
         );
  INV_X1 U9424 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n7667) );
  NAND2_X1 U9425 ( .A1(n10168), .A2(n7665), .ZN(n7666) );
  NAND2_X1 U9426 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n8229) );
  OAI211_X1 U9427 ( .C1(n7667), .C2(n10220), .A(n7666), .B(n8229), .ZN(n7668)
         );
  OR3_X1 U9428 ( .A1(n7670), .A2(n7669), .A3(n7668), .ZN(P1_U3251) );
  AOI211_X1 U9429 ( .C1(n7673), .C2(n7672), .A(n10158), .B(n7671), .ZN(n7682)
         );
  AOI211_X1 U9430 ( .C1(n4321), .C2(n7675), .A(n10206), .B(n7674), .ZN(n7681)
         );
  INV_X1 U9431 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7679) );
  NAND2_X1 U9432 ( .A1(n10168), .A2(n7676), .ZN(n7678) );
  NOR2_X1 U9433 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5332), .ZN(n7867) );
  INV_X1 U9434 ( .A(n7867), .ZN(n7677) );
  OAI211_X1 U9435 ( .C1(n7679), .C2(n10220), .A(n7678), .B(n7677), .ZN(n7680)
         );
  OR3_X1 U9436 ( .A1(n7682), .A2(n7681), .A3(n7680), .ZN(P1_U3250) );
  OAI21_X1 U9437 ( .B1(n7684), .B2(n7683), .A(n7699), .ZN(n7685) );
  AOI222_X1 U9438 ( .A1(n9966), .A2(n7685), .B1(n9679), .B2(n9934), .C1(n9681), 
        .C2(n9932), .ZN(n10240) );
  NAND2_X1 U9439 ( .A1(n7687), .A2(n7686), .ZN(n7689) );
  NAND2_X1 U9440 ( .A1(n7689), .A2(n7688), .ZN(n7703) );
  OAI21_X1 U9441 ( .B1(n7689), .B2(n7688), .A(n7703), .ZN(n10243) );
  NAND2_X1 U9442 ( .A1(n7691), .A2(n7690), .ZN(n7692) );
  NAND3_X1 U9443 ( .A1(n7709), .A2(n10015), .A3(n7692), .ZN(n10238) );
  OAI22_X1 U9444 ( .A1(n10224), .A2(n10238), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10221), .ZN(n7693) );
  INV_X1 U9445 ( .A(n7693), .ZN(n7695) );
  NAND2_X1 U9446 ( .A1(n4287), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n7694) );
  OAI211_X1 U9447 ( .C1(n10227), .C2(n10239), .A(n7695), .B(n7694), .ZN(n7696)
         );
  AOI21_X1 U9448 ( .B1(n10231), .B2(n10243), .A(n7696), .ZN(n7697) );
  OAI21_X1 U9449 ( .B1(n10240), .B2(n4287), .A(n7697), .ZN(P1_U3290) );
  NAND2_X1 U9450 ( .A1(n7699), .A2(n7698), .ZN(n7700) );
  XOR2_X1 U9451 ( .A(n7704), .B(n7700), .Z(n7701) );
  AOI222_X1 U9452 ( .A1(n9966), .A2(n7701), .B1(n4587), .B2(n9934), .C1(n9680), 
        .C2(n9932), .ZN(n10246) );
  NAND2_X1 U9453 ( .A1(n7703), .A2(n7702), .ZN(n7705) );
  XNOR2_X1 U9454 ( .A(n7705), .B(n7704), .ZN(n10249) );
  NOR2_X1 U9455 ( .A1(n10221), .A2(n7706), .ZN(n7707) );
  AOI21_X1 U9456 ( .B1(n4287), .B2(P1_REG2_REG_4__SCAN_IN), .A(n7707), .ZN(
        n7714) );
  NAND2_X1 U9457 ( .A1(n7709), .A2(n7708), .ZN(n7710) );
  NAND2_X1 U9458 ( .A1(n7710), .A2(n10015), .ZN(n7712) );
  OR2_X1 U9459 ( .A1(n7712), .A2(n7711), .ZN(n10244) );
  OR2_X1 U9460 ( .A1(n10224), .A2(n10244), .ZN(n7713) );
  OAI211_X1 U9461 ( .C1(n10227), .C2(n10245), .A(n7714), .B(n7713), .ZN(n7715)
         );
  AOI21_X1 U9462 ( .B1(n10231), .B2(n10249), .A(n7715), .ZN(n7716) );
  OAI21_X1 U9463 ( .B1(n10246), .B2(n4287), .A(n7716), .ZN(P1_U3289) );
  NAND3_X1 U9464 ( .A1(n7719), .A2(n7718), .A3(n7717), .ZN(n7721) );
  AND2_X1 U9465 ( .A1(n7721), .A2(n7720), .ZN(n7723) );
  OAI22_X1 U9466 ( .A1(n4287), .A2(n7723), .B1(n7722), .B2(n10221), .ZN(n7724)
         );
  AOI21_X1 U9467 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n4287), .A(n7724), .ZN(
        n7727) );
  NOR2_X1 U9468 ( .A1(n10224), .A2(n9952), .ZN(n9864) );
  OAI21_X1 U9469 ( .B1(n9973), .B2(n9864), .A(n7725), .ZN(n7726) );
  NAND2_X1 U9470 ( .A1(n7727), .A2(n7726), .ZN(P1_U3293) );
  NAND2_X1 U9471 ( .A1(n9670), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7728) );
  OAI21_X1 U9472 ( .B1(n7729), .B2(n9670), .A(n7728), .ZN(P1_U3583) );
  NAND2_X1 U9473 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  XNOR2_X1 U9474 ( .A(n7730), .B(n7733), .ZN(n7734) );
  NAND2_X1 U9475 ( .A1(n7734), .A2(n9621), .ZN(n7740) );
  NOR2_X1 U9476 ( .A1(n9643), .A2(n8230), .ZN(n7738) );
  OAI21_X1 U9477 ( .B1(n9654), .B2(n7736), .A(n7735), .ZN(n7737) );
  AOI211_X1 U9478 ( .C1(n10260), .C2(n9659), .A(n7738), .B(n7737), .ZN(n7739)
         );
  OAI211_X1 U9479 ( .C1(n9636), .C2(n7769), .A(n7740), .B(n7739), .ZN(P1_U3239) );
  OAI22_X1 U9480 ( .A1(n10224), .A2(n7742), .B1(n7741), .B2(n10221), .ZN(n7743) );
  AOI21_X1 U9481 ( .B1(n9973), .B2(n7744), .A(n7743), .ZN(n7747) );
  MUX2_X1 U9482 ( .A(n7745), .B(n6465), .S(n4287), .Z(n7746) );
  OAI211_X1 U9483 ( .C1(n7748), .C2(n9929), .A(n7747), .B(n7746), .ZN(P1_U3292) );
  NAND2_X1 U9484 ( .A1(n7750), .A2(n7749), .ZN(n7754) );
  XNOR2_X1 U9485 ( .A(n7752), .B(n7751), .ZN(n7753) );
  XNOR2_X1 U9486 ( .A(n7754), .B(n7753), .ZN(n7755) );
  NAND2_X1 U9487 ( .A1(n7755), .A2(n9621), .ZN(n7761) );
  NAND2_X1 U9488 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9711) );
  INV_X1 U9489 ( .A(n9711), .ZN(n7759) );
  OAI22_X1 U9490 ( .A1(n9630), .A2(n7757), .B1(n7756), .B2(n9643), .ZN(n7758)
         );
  AOI211_X1 U9491 ( .C1(n9640), .C2(n9679), .A(n7759), .B(n7758), .ZN(n7760)
         );
  OAI211_X1 U9492 ( .C1(n9636), .C2(n7762), .A(n7761), .B(n7760), .ZN(P1_U3227) );
  XOR2_X1 U9493 ( .A(n7763), .B(n7765), .Z(n10264) );
  XNOR2_X1 U9494 ( .A(n7764), .B(n7765), .ZN(n7766) );
  AOI222_X1 U9495 ( .A1(n9966), .A2(n7766), .B1(n9677), .B2(n9934), .C1(n4587), 
        .C2(n9932), .ZN(n10263) );
  MUX2_X1 U9496 ( .A(n7767), .B(n10263), .S(n9971), .Z(n7772) );
  AOI211_X1 U9497 ( .C1(n10260), .C2(n7768), .A(n9952), .B(n4416), .ZN(n10259)
         );
  OAI22_X1 U9498 ( .A1(n10227), .A2(n5811), .B1(n10221), .B2(n7769), .ZN(n7770) );
  AOI21_X1 U9499 ( .B1(n10259), .B2(n9944), .A(n7770), .ZN(n7771) );
  OAI211_X1 U9500 ( .C1(n10264), .C2(n9929), .A(n7772), .B(n7771), .ZN(
        P1_U3287) );
  XOR2_X1 U9501 ( .A(n7774), .B(n7773), .Z(n7791) );
  INV_X1 U9502 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n7775) );
  NAND2_X1 U9503 ( .A1(P2_U3151), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n7966) );
  OAI21_X1 U9504 ( .B1(n8976), .B2(n7775), .A(n7966), .ZN(n7782) );
  OR3_X1 U9505 ( .A1(n7778), .A2(n7777), .A3(n7776), .ZN(n7779) );
  AOI21_X1 U9506 ( .B1(n7780), .B2(n7779), .A(n9086), .ZN(n7781) );
  AOI211_X1 U9507 ( .C1(n8985), .C2(n7783), .A(n7782), .B(n7781), .ZN(n7790)
         );
  INV_X1 U9508 ( .A(n7784), .ZN(n7788) );
  NOR3_X1 U9509 ( .A1(n7786), .A2(n7625), .A3(n7785), .ZN(n7787) );
  OAI21_X1 U9510 ( .B1(n7788), .B2(n7787), .A(n6685), .ZN(n7789) );
  OAI211_X1 U9511 ( .C1(n7791), .C2(n9075), .A(n7790), .B(n7789), .ZN(P2_U3190) );
  XNOR2_X1 U9512 ( .A(n9364), .B(n7357), .ZN(n7961) );
  XNOR2_X1 U9513 ( .A(n7961), .B(n7968), .ZN(n7799) );
  INV_X1 U9514 ( .A(n7792), .ZN(n7793) );
  NAND2_X1 U9515 ( .A1(n7793), .A2(n9293), .ZN(n7794) );
  INV_X1 U9516 ( .A(n7799), .ZN(n7796) );
  INV_X1 U9517 ( .A(n7963), .ZN(n7797) );
  AOI21_X1 U9518 ( .B1(n7799), .B2(n7798), .A(n7797), .ZN(n7807) );
  INV_X1 U9519 ( .A(n7800), .ZN(n9298) );
  NAND2_X1 U9520 ( .A1(n8920), .A2(n9298), .ZN(n7804) );
  INV_X1 U9521 ( .A(n7801), .ZN(n7802) );
  AOI21_X1 U9522 ( .B1(n8916), .B2(n9293), .A(n7802), .ZN(n7803) );
  OAI211_X1 U9523 ( .C1(n8071), .C2(n8918), .A(n7804), .B(n7803), .ZN(n7805)
         );
  AOI21_X1 U9524 ( .B1(n9364), .B2(n8908), .A(n7805), .ZN(n7806) );
  OAI21_X1 U9525 ( .B1(n7807), .B2(n8910), .A(n7806), .ZN(P2_U3153) );
  AOI211_X1 U9526 ( .C1(n7810), .C2(n7809), .A(n10158), .B(n7808), .ZN(n7819)
         );
  AOI211_X1 U9527 ( .C1(n7813), .C2(n7812), .A(n10206), .B(n7811), .ZN(n7818)
         );
  NAND2_X1 U9528 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8319) );
  INV_X1 U9529 ( .A(n8319), .ZN(n7814) );
  AOI21_X1 U9530 ( .B1(n10141), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n7814), .ZN(
        n7815) );
  OAI21_X1 U9531 ( .B1(n10215), .B2(n7816), .A(n7815), .ZN(n7817) );
  OR3_X1 U9532 ( .A1(n7819), .A2(n7818), .A3(n7817), .ZN(P1_U3253) );
  AND2_X1 U9533 ( .A1(n7821), .A2(n7820), .ZN(n8013) );
  OR2_X1 U9534 ( .A1(n7822), .A2(n9301), .ZN(n9287) );
  NAND3_X1 U9535 ( .A1(n9287), .A2(n7824), .A3(n7823), .ZN(n7825) );
  NAND2_X1 U9536 ( .A1(n8013), .A2(n7825), .ZN(n7826) );
  AOI222_X1 U9537 ( .A1(n9295), .A2(n7826), .B1(n8931), .B2(n9292), .C1(n8930), 
        .C2(n9290), .ZN(n8002) );
  AOI22_X1 U9538 ( .A1(n9463), .A2(n8004), .B1(P2_REG0_REG_8__SCAN_IN), .B2(
        n10301), .ZN(n7832) );
  NAND2_X1 U9539 ( .A1(n7827), .A2(n7828), .ZN(n7829) );
  XNOR2_X1 U9540 ( .A(n7829), .B(n8555), .ZN(n8001) );
  NAND2_X1 U9541 ( .A1(n8001), .A2(n9428), .ZN(n7831) );
  OAI211_X1 U9542 ( .C1(n8002), .C2(n10301), .A(n7832), .B(n7831), .ZN(
        P2_U3414) );
  INV_X1 U9543 ( .A(n7833), .ZN(n7834) );
  NAND2_X1 U9544 ( .A1(n6620), .A2(n7834), .ZN(n7946) );
  NAND2_X1 U9545 ( .A1(n8050), .A2(n7946), .ZN(n7835) );
  NAND2_X1 U9546 ( .A1(n9300), .A2(n7836), .ZN(n7839) );
  NAND2_X1 U9547 ( .A1(n9299), .A2(n7837), .ZN(n7838) );
  OAI211_X1 U9548 ( .C1(n6771), .C2(n9296), .A(n7839), .B(n7838), .ZN(n7842)
         );
  NOR2_X1 U9549 ( .A1(n7840), .A2(n9273), .ZN(n7841) );
  AOI211_X1 U9550 ( .C1(n7843), .C2(n9303), .A(n7842), .B(n7841), .ZN(n7844)
         );
  INV_X1 U9551 ( .A(n7844), .ZN(P2_U3229) );
  INV_X1 U9552 ( .A(n7764), .ZN(n7847) );
  OAI21_X1 U9553 ( .B1(n7847), .B2(n7846), .A(n7845), .ZN(n7848) );
  NOR2_X1 U9554 ( .A1(n7848), .A2(n7850), .ZN(n7936) );
  AOI21_X1 U9555 ( .B1(n7850), .B2(n7848), .A(n7936), .ZN(n7854) );
  AOI22_X1 U9556 ( .A1(n9934), .A2(n9676), .B1(n9678), .B2(n9932), .ZN(n7853)
         );
  XNOR2_X1 U9557 ( .A(n7849), .B(n7850), .ZN(n10271) );
  INV_X1 U9558 ( .A(n10278), .ZN(n7851) );
  NAND2_X1 U9559 ( .A1(n10271), .A2(n7851), .ZN(n7852) );
  OAI211_X1 U9560 ( .C1(n7854), .C2(n9916), .A(n7853), .B(n7852), .ZN(n10269)
         );
  INV_X1 U9561 ( .A(n10271), .ZN(n7857) );
  INV_X1 U9562 ( .A(n7941), .ZN(n7855) );
  OAI211_X1 U9563 ( .C1(n4933), .C2(n4416), .A(n7855), .B(n10015), .ZN(n10268)
         );
  OAI22_X1 U9564 ( .A1(n7857), .A2(n9968), .B1(n7856), .B2(n10268), .ZN(n7858)
         );
  OAI21_X1 U9565 ( .B1(n10269), .B2(n7858), .A(n9971), .ZN(n7861) );
  INV_X1 U9566 ( .A(n7866), .ZN(n7859) );
  INV_X1 U9567 ( .A(n10221), .ZN(n9922) );
  AOI22_X1 U9568 ( .A1(n4287), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7859), .B2(
        n9922), .ZN(n7860) );
  OAI211_X1 U9569 ( .C1(n4933), .C2(n10227), .A(n7861), .B(n7860), .ZN(
        P1_U3286) );
  XNOR2_X1 U9570 ( .A(n7864), .B(n7863), .ZN(n7865) );
  XNOR2_X1 U9571 ( .A(n7862), .B(n7865), .ZN(n7873) );
  NOR2_X1 U9572 ( .A1(n9636), .A2(n7866), .ZN(n7872) );
  AOI21_X1 U9573 ( .B1(n9640), .B2(n9678), .A(n7867), .ZN(n7870) );
  NAND2_X1 U9574 ( .A1(n9659), .A2(n7868), .ZN(n7869) );
  OAI211_X1 U9575 ( .C1(n8264), .C2(n9643), .A(n7870), .B(n7869), .ZN(n7871)
         );
  AOI211_X1 U9576 ( .C1(n7873), .C2(n9621), .A(n7872), .B(n7871), .ZN(n7874)
         );
  INV_X1 U9577 ( .A(n7874), .ZN(P1_U3213) );
  INV_X1 U9578 ( .A(n7875), .ZN(n8810) );
  OAI222_X1 U9579 ( .A1(n9490), .A2(n8785), .B1(n9481), .B2(n8810), .C1(
        P2_U3151), .C2(n4302), .ZN(P2_U3276) );
  INV_X1 U9580 ( .A(n7876), .ZN(n7883) );
  NOR2_X1 U9581 ( .A1(n9238), .A2(n6748), .ZN(n7878) );
  AOI211_X1 U9582 ( .C1(n7879), .C2(n8534), .A(n7878), .B(n7877), .ZN(n7880)
         );
  MUX2_X1 U9583 ( .A(n7881), .B(n7880), .S(n9296), .Z(n7882) );
  OAI21_X1 U9584 ( .B1(n7883), .B2(n9264), .A(n7882), .ZN(P2_U3231) );
  XNOR2_X1 U9585 ( .A(n7884), .B(n7888), .ZN(n8093) );
  INV_X1 U9586 ( .A(n8093), .ZN(n7899) );
  INV_X1 U9587 ( .A(n7885), .ZN(n7886) );
  AOI21_X1 U9588 ( .B1(n7888), .B2(n7887), .A(n7886), .ZN(n7889) );
  OAI222_X1 U9589 ( .A1(n9962), .A2(n8320), .B1(n9960), .B2(n7890), .C1(n9916), 
        .C2(n7889), .ZN(n8091) );
  INV_X1 U9590 ( .A(n8325), .ZN(n7896) );
  INV_X1 U9591 ( .A(n7891), .ZN(n7978) );
  INV_X1 U9592 ( .A(n7995), .ZN(n7892) );
  AOI211_X1 U9593 ( .C1(n8325), .C2(n7978), .A(n9952), .B(n7892), .ZN(n8092)
         );
  NAND2_X1 U9594 ( .A1(n8092), .A2(n9944), .ZN(n7895) );
  INV_X1 U9595 ( .A(n8323), .ZN(n7893) );
  AOI22_X1 U9596 ( .A1(n4287), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7893), .B2(
        n9922), .ZN(n7894) );
  OAI211_X1 U9597 ( .C1(n7896), .C2(n10227), .A(n7895), .B(n7894), .ZN(n7897)
         );
  AOI21_X1 U9598 ( .B1(n8091), .B2(n9971), .A(n7897), .ZN(n7898) );
  OAI21_X1 U9599 ( .B1(n7899), .B2(n9929), .A(n7898), .ZN(P1_U3283) );
  INV_X1 U9600 ( .A(n7900), .ZN(n7907) );
  MUX2_X1 U9601 ( .A(n7902), .B(n7901), .S(n9296), .Z(n7906) );
  AOI22_X1 U9602 ( .A1(n9300), .A2(n7904), .B1(n9299), .B2(n7903), .ZN(n7905)
         );
  OAI211_X1 U9603 ( .C1(n7907), .C2(n9264), .A(n7906), .B(n7905), .ZN(P2_U3228) );
  XNOR2_X1 U9604 ( .A(n7568), .B(n8549), .ZN(n9377) );
  INV_X1 U9605 ( .A(n9377), .ZN(n7918) );
  INV_X1 U9606 ( .A(n8549), .ZN(n7908) );
  XNOR2_X1 U9607 ( .A(n7909), .B(n7908), .ZN(n7910) );
  NAND2_X1 U9608 ( .A1(n7910), .A2(n9295), .ZN(n7913) );
  AOI22_X1 U9609 ( .A1(n9292), .A2(n8934), .B1(n7911), .B2(n9290), .ZN(n7912)
         );
  AND2_X1 U9610 ( .A1(n7913), .A2(n7912), .ZN(n9382) );
  MUX2_X1 U9611 ( .A(n9382), .B(n7914), .S(n9273), .Z(n7917) );
  AOI22_X1 U9612 ( .A1(n9300), .A2(n9379), .B1(n7915), .B2(n9299), .ZN(n7916)
         );
  OAI211_X1 U9613 ( .C1(n7918), .C2(n9264), .A(n7917), .B(n7916), .ZN(P2_U3230) );
  NAND2_X1 U9614 ( .A1(n7920), .A2(n7919), .ZN(n7922) );
  INV_X1 U9615 ( .A(n7921), .ZN(n8554) );
  XNOR2_X1 U9616 ( .A(n7922), .B(n8554), .ZN(n9370) );
  INV_X1 U9617 ( .A(n9370), .ZN(n7931) );
  XNOR2_X1 U9618 ( .A(n4279), .B(n8554), .ZN(n7926) );
  NAND2_X1 U9619 ( .A1(n8932), .A2(n9292), .ZN(n7924) );
  OAI21_X1 U9620 ( .B1(n7968), .B2(n9234), .A(n7924), .ZN(n7925) );
  AOI21_X1 U9621 ( .B1(n7926), .B2(n9295), .A(n7925), .ZN(n9374) );
  MUX2_X1 U9622 ( .A(n9374), .B(n7927), .S(n9273), .Z(n7930) );
  AOI22_X1 U9623 ( .A1(n9300), .A2(n9371), .B1(n9299), .B2(n7928), .ZN(n7929)
         );
  OAI211_X1 U9624 ( .C1(n7931), .C2(n9264), .A(n7930), .B(n7929), .ZN(P2_U3227) );
  INV_X1 U9625 ( .A(n7933), .ZN(n7937) );
  XNOR2_X1 U9626 ( .A(n7932), .B(n7937), .ZN(n10276) );
  INV_X1 U9627 ( .A(n7934), .ZN(n7935) );
  NOR2_X1 U9628 ( .A1(n7936), .A2(n7935), .ZN(n7938) );
  NAND2_X1 U9629 ( .A1(n7938), .A2(n7937), .ZN(n7974) );
  OAI211_X1 U9630 ( .C1(n7938), .C2(n7937), .A(n7974), .B(n9966), .ZN(n7940)
         );
  AOI22_X1 U9631 ( .A1(n9934), .A2(n9675), .B1(n9677), .B2(n9932), .ZN(n7939)
         );
  NAND2_X1 U9632 ( .A1(n7940), .A2(n7939), .ZN(n10281) );
  NAND2_X1 U9633 ( .A1(n10281), .A2(n9971), .ZN(n7945) );
  OAI22_X1 U9634 ( .A1(n9971), .A2(n4824), .B1(n8233), .B2(n10221), .ZN(n7943)
         );
  OAI211_X1 U9635 ( .C1(n7941), .C2(n10275), .A(n7977), .B(n10015), .ZN(n10273) );
  NOR2_X1 U9636 ( .A1(n10273), .A2(n10224), .ZN(n7942) );
  AOI211_X1 U9637 ( .C1(n9973), .C2(n8235), .A(n7943), .B(n7942), .ZN(n7944)
         );
  OAI211_X1 U9638 ( .C1(n10276), .C2(n9929), .A(n7945), .B(n7944), .ZN(
        P1_U3285) );
  INV_X1 U9639 ( .A(n7946), .ZN(n7947) );
  NAND2_X1 U9640 ( .A1(n9296), .A2(n7947), .ZN(n8178) );
  INV_X1 U9641 ( .A(n8178), .ZN(n7956) );
  OAI21_X1 U9642 ( .B1(n7949), .B2(n8050), .A(n7948), .ZN(n7950) );
  MUX2_X1 U9643 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7950), .S(n9296), .Z(n7954)
         );
  INV_X1 U9644 ( .A(n9300), .ZN(n9115) );
  OAI22_X1 U9645 ( .A1(n9115), .A2(n7952), .B1(n7951), .B2(n9238), .ZN(n7953)
         );
  AOI211_X1 U9646 ( .C1(n7956), .C2(n7955), .A(n7954), .B(n7953), .ZN(n7957)
         );
  INV_X1 U9647 ( .A(n7957), .ZN(P2_U3232) );
  MUX2_X1 U9648 ( .A(n7958), .B(n8002), .S(n9383), .Z(n7960) );
  AOI22_X1 U9649 ( .A1(n8001), .A2(n9332), .B1(n9356), .B2(n8004), .ZN(n7959)
         );
  NAND2_X1 U9650 ( .A1(n7960), .A2(n7959), .ZN(P2_U3467) );
  NAND2_X1 U9651 ( .A1(n7961), .A2(n7968), .ZN(n7962) );
  XNOR2_X1 U9652 ( .A(n8004), .B(n7357), .ZN(n8072) );
  INV_X1 U9653 ( .A(n8072), .ZN(n8070) );
  XNOR2_X1 U9654 ( .A(n8078), .B(n8070), .ZN(n8060) );
  XNOR2_X1 U9655 ( .A(n8060), .B(n9291), .ZN(n7972) );
  INV_X1 U9656 ( .A(n7964), .ZN(n8003) );
  INV_X1 U9657 ( .A(n8004), .ZN(n7965) );
  NOR2_X1 U9658 ( .A1(n8923), .A2(n7965), .ZN(n7970) );
  NAND2_X1 U9659 ( .A1(n8902), .A2(n8930), .ZN(n7967) );
  OAI211_X1 U9660 ( .C1(n7968), .C2(n8905), .A(n7967), .B(n7966), .ZN(n7969)
         );
  AOI211_X1 U9661 ( .C1(n8003), .C2(n8920), .A(n7970), .B(n7969), .ZN(n7971)
         );
  OAI21_X1 U9662 ( .B1(n7972), .B2(n8910), .A(n7971), .ZN(P2_U3161) );
  NAND2_X1 U9663 ( .A1(n7974), .A2(n7973), .ZN(n7975) );
  XNOR2_X1 U9664 ( .A(n7975), .B(n7984), .ZN(n7976) );
  AOI22_X1 U9665 ( .A1(n7976), .A2(n9966), .B1(n9932), .B2(n9676), .ZN(n8130)
         );
  INV_X1 U9666 ( .A(n7977), .ZN(n7979) );
  INV_X1 U9667 ( .A(n8128), .ZN(n8270) );
  OAI211_X1 U9668 ( .C1(n7979), .C2(n8270), .A(n10015), .B(n7978), .ZN(n7980)
         );
  OAI21_X1 U9669 ( .B1(n7993), .B2(n9962), .A(n7980), .ZN(n8127) );
  NOR2_X1 U9670 ( .A1(n10221), .A2(n8265), .ZN(n7981) );
  AOI21_X1 U9671 ( .B1(n4287), .B2(P1_REG2_REG_9__SCAN_IN), .A(n7981), .ZN(
        n7982) );
  OAI21_X1 U9672 ( .B1(n10227), .B2(n8270), .A(n7982), .ZN(n7986) );
  XOR2_X1 U9673 ( .A(n7983), .B(n7984), .Z(n8131) );
  NOR2_X1 U9674 ( .A1(n8131), .A2(n9929), .ZN(n7985) );
  AOI211_X1 U9675 ( .C1(n9944), .C2(n8127), .A(n7986), .B(n7985), .ZN(n7987)
         );
  OAI21_X1 U9676 ( .B1(n8130), .B2(n4287), .A(n7987), .ZN(P1_U3284) );
  XNOR2_X1 U9677 ( .A(n7988), .B(n7989), .ZN(n10067) );
  XNOR2_X1 U9678 ( .A(n7990), .B(n7991), .ZN(n7992) );
  OAI222_X1 U9679 ( .A1(n9962), .A2(n9610), .B1(n9960), .B2(n7993), .C1(n7992), 
        .C2(n9916), .ZN(n10063) );
  AOI211_X1 U9680 ( .C1(n10065), .C2(n7995), .A(n9952), .B(n7994), .ZN(n10064)
         );
  NAND2_X1 U9681 ( .A1(n10064), .A2(n9944), .ZN(n7998) );
  INV_X1 U9682 ( .A(n8365), .ZN(n7996) );
  AOI22_X1 U9683 ( .A1(n4287), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7996), .B2(
        n9922), .ZN(n7997) );
  OAI211_X1 U9684 ( .C1(n8370), .C2(n10227), .A(n7998), .B(n7997), .ZN(n7999)
         );
  AOI21_X1 U9685 ( .B1(n9971), .B2(n10063), .A(n7999), .ZN(n8000) );
  OAI21_X1 U9686 ( .B1(n10067), .B2(n9929), .A(n8000), .ZN(P1_U3282) );
  INV_X1 U9687 ( .A(n8001), .ZN(n8007) );
  MUX2_X1 U9688 ( .A(n8709), .B(n8002), .S(n9296), .Z(n8006) );
  AOI22_X1 U9689 ( .A1(n9300), .A2(n8004), .B1(n9299), .B2(n8003), .ZN(n8005)
         );
  OAI211_X1 U9690 ( .C1(n8007), .C2(n9264), .A(n8006), .B(n8005), .ZN(P2_U3225) );
  INV_X1 U9691 ( .A(n8008), .ZN(n8052) );
  NAND2_X1 U9692 ( .A1(n8009), .A2(n8556), .ZN(n8010) );
  NAND2_X1 U9693 ( .A1(n8039), .A2(n8010), .ZN(n8059) );
  INV_X1 U9694 ( .A(n8059), .ZN(n8018) );
  NAND2_X1 U9695 ( .A1(n8011), .A2(n8556), .ZN(n8045) );
  INV_X1 U9696 ( .A(n8045), .ZN(n8015) );
  AND3_X1 U9697 ( .A1(n8013), .A2(n7066), .A3(n8012), .ZN(n8014) );
  OAI21_X1 U9698 ( .B1(n8015), .B2(n8014), .A(n9295), .ZN(n8017) );
  AOI22_X1 U9699 ( .A1(n9291), .A2(n9292), .B1(n9290), .B2(n8929), .ZN(n8016)
         );
  OAI211_X1 U9700 ( .C1(n8059), .C2(n8050), .A(n8017), .B(n8016), .ZN(n8054)
         );
  AOI21_X1 U9701 ( .B1(n8052), .B2(n8018), .A(n8054), .ZN(n8111) );
  AOI22_X1 U9702 ( .A1(n9463), .A2(n8063), .B1(P2_REG0_REG_9__SCAN_IN), .B2(
        n10301), .ZN(n8019) );
  OAI21_X1 U9703 ( .B1(n8111), .B2(n10301), .A(n8019), .ZN(P2_U3417) );
  AOI211_X1 U9704 ( .C1(n8022), .C2(n8021), .A(n10158), .B(n8020), .ZN(n8031)
         );
  AOI211_X1 U9705 ( .C1(n8025), .C2(n8024), .A(n10206), .B(n8023), .ZN(n8030)
         );
  NAND2_X1 U9706 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n8364) );
  INV_X1 U9707 ( .A(n8364), .ZN(n8026) );
  AOI21_X1 U9708 ( .B1(n10141), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n8026), .ZN(
        n8027) );
  OAI21_X1 U9709 ( .B1(n10215), .B2(n8028), .A(n8027), .ZN(n8029) );
  OR3_X1 U9710 ( .A1(n8031), .A2(n8030), .A3(n8029), .ZN(P1_U3254) );
  INV_X1 U9711 ( .A(n8033), .ZN(n8412) );
  XNOR2_X1 U9712 ( .A(n8032), .B(n8412), .ZN(n8198) );
  INV_X1 U9713 ( .A(n9292), .ZN(n9236) );
  XNOR2_X1 U9714 ( .A(n8034), .B(n8033), .ZN(n8035) );
  OAI222_X1 U9715 ( .A1(n9236), .A2(n8079), .B1(n9234), .B2(n8293), .C1(n8035), 
        .C2(n9231), .ZN(n8193) );
  NAND2_X1 U9716 ( .A1(n8193), .A2(n9296), .ZN(n8038) );
  OAI22_X1 U9717 ( .A1(n9296), .A2(n8957), .B1(n8208), .B2(n9238), .ZN(n8036)
         );
  AOI21_X1 U9718 ( .B1(n8210), .B2(n9300), .A(n8036), .ZN(n8037) );
  OAI211_X1 U9719 ( .C1(n8198), .C2(n9264), .A(n8038), .B(n8037), .ZN(P2_U3222) );
  NAND2_X1 U9720 ( .A1(n8039), .A2(n8434), .ZN(n8043) );
  INV_X1 U9721 ( .A(n8558), .ZN(n8042) );
  XNOR2_X1 U9722 ( .A(n8043), .B(n8042), .ZN(n8179) );
  INV_X1 U9723 ( .A(n8179), .ZN(n8051) );
  NAND2_X1 U9724 ( .A1(n8045), .A2(n8044), .ZN(n8046) );
  XNOR2_X1 U9725 ( .A(n8046), .B(n8558), .ZN(n8047) );
  NAND2_X1 U9726 ( .A1(n8047), .A2(n9295), .ZN(n8049) );
  AOI22_X1 U9727 ( .A1(n8930), .A2(n9292), .B1(n9290), .B2(n9276), .ZN(n8048)
         );
  OAI211_X1 U9728 ( .C1(n8179), .C2(n8050), .A(n8049), .B(n8048), .ZN(n8171)
         );
  AOI21_X1 U9729 ( .B1(n8052), .B2(n8051), .A(n8171), .ZN(n8215) );
  AOI22_X1 U9730 ( .A1(n9463), .A2(n8175), .B1(P2_REG0_REG_10__SCAN_IN), .B2(
        n10301), .ZN(n8053) );
  OAI21_X1 U9731 ( .B1(n8215), .B2(n10301), .A(n8053), .ZN(P2_U3420) );
  INV_X1 U9732 ( .A(n8054), .ZN(n8055) );
  MUX2_X1 U9733 ( .A(n8055), .B(n8156), .S(n9273), .Z(n8058) );
  INV_X1 U9734 ( .A(n8056), .ZN(n8067) );
  AOI22_X1 U9735 ( .A1(n9300), .A2(n8063), .B1(n9299), .B2(n8067), .ZN(n8057)
         );
  OAI211_X1 U9736 ( .C1(n8059), .C2(n8178), .A(n8058), .B(n8057), .ZN(P2_U3224) );
  AOI22_X1 U9737 ( .A1(n8060), .A2(n8071), .B1(n8078), .B2(n8072), .ZN(n8062)
         );
  XOR2_X1 U9738 ( .A(n7357), .B(n8063), .Z(n8075) );
  XNOR2_X1 U9739 ( .A(n8075), .B(n8103), .ZN(n8061) );
  XNOR2_X1 U9740 ( .A(n8062), .B(n8061), .ZN(n8069) );
  INV_X1 U9741 ( .A(n8063), .ZN(n8113) );
  NOR2_X1 U9742 ( .A1(n8923), .A2(n8113), .ZN(n8066) );
  NAND2_X1 U9743 ( .A1(n8902), .A2(n8929), .ZN(n8064) );
  NAND2_X1 U9744 ( .A1(P2_U3151), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8157) );
  OAI211_X1 U9745 ( .C1(n8071), .C2(n8905), .A(n8064), .B(n8157), .ZN(n8065)
         );
  AOI211_X1 U9746 ( .C1(n8067), .C2(n8920), .A(n8066), .B(n8065), .ZN(n8068)
         );
  OAI21_X1 U9747 ( .B1(n8069), .B2(n8910), .A(n8068), .ZN(P2_U3171) );
  OAI22_X1 U9748 ( .A1(n8075), .A2(n8930), .B1(n8070), .B2(n9291), .ZN(n8077)
         );
  OAI21_X1 U9749 ( .B1(n8072), .B2(n8071), .A(n8103), .ZN(n8074) );
  NOR3_X1 U9750 ( .A1(n8072), .A2(n8071), .A3(n8103), .ZN(n8073) );
  AOI21_X1 U9751 ( .B1(n8075), .B2(n8074), .A(n8073), .ZN(n8076) );
  XNOR2_X1 U9752 ( .A(n8210), .B(n7357), .ZN(n8203) );
  XNOR2_X1 U9753 ( .A(n8175), .B(n7357), .ZN(n8100) );
  AOI22_X1 U9754 ( .A1(n8203), .A2(n8202), .B1(n8079), .B2(n8100), .ZN(n8083)
         );
  INV_X1 U9755 ( .A(n8100), .ZN(n8200) );
  AOI21_X1 U9756 ( .B1(n8200), .B2(n8929), .A(n9276), .ZN(n8081) );
  NAND2_X1 U9757 ( .A1(n9276), .A2(n8929), .ZN(n8080) );
  OAI22_X1 U9758 ( .A1(n8203), .A2(n8081), .B1(n8100), .B2(n8080), .ZN(n8082)
         );
  XNOR2_X1 U9759 ( .A(n7068), .B(n7357), .ZN(n8292) );
  XNOR2_X1 U9760 ( .A(n8292), .B(n8293), .ZN(n8084) );
  XNOR2_X1 U9761 ( .A(n8291), .B(n8084), .ZN(n8090) );
  NAND2_X1 U9762 ( .A1(n8916), .A2(n9276), .ZN(n8085) );
  NAND2_X1 U9763 ( .A1(P2_U3151), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8974) );
  OAI211_X1 U9764 ( .C1(n8086), .C2(n8918), .A(n8085), .B(n8974), .ZN(n8088)
         );
  INV_X1 U9765 ( .A(n7068), .ZN(n9363) );
  NOR2_X1 U9766 ( .A1(n9363), .A2(n8923), .ZN(n8087) );
  AOI211_X1 U9767 ( .C1(n9280), .C2(n8920), .A(n8088), .B(n8087), .ZN(n8089)
         );
  OAI21_X1 U9768 ( .B1(n8090), .B2(n8910), .A(n8089), .ZN(P2_U3164) );
  AOI211_X1 U9769 ( .C1(n10250), .C2(n8093), .A(n8092), .B(n8091), .ZN(n8096)
         );
  AOI22_X1 U9770 ( .A1(n8283), .A2(n8325), .B1(P1_REG0_REG_10__SCAN_IN), .B2(
        n10282), .ZN(n8094) );
  OAI21_X1 U9771 ( .B1(n8096), .B2(n10282), .A(n8094), .ZN(P1_U3483) );
  INV_X1 U9772 ( .A(n10048), .ZN(n8281) );
  AOI22_X1 U9773 ( .A1(n8281), .A2(n8325), .B1(P1_REG1_REG_10__SCAN_IN), .B2(
        n10289), .ZN(n8095) );
  OAI21_X1 U9774 ( .B1(n8096), .B2(n10289), .A(n8095), .ZN(P1_U3532) );
  INV_X1 U9775 ( .A(n8097), .ZN(n8109) );
  OAI222_X1 U9776 ( .A1(n9481), .A2(n8109), .B1(n8099), .B2(P2_U3151), .C1(
        n8098), .C2(n9494), .ZN(P2_U3275) );
  XNOR2_X1 U9777 ( .A(n8199), .B(n8929), .ZN(n8201) );
  XNOR2_X1 U9778 ( .A(n8201), .B(n8100), .ZN(n8107) );
  INV_X1 U9779 ( .A(n8101), .ZN(n8174) );
  NAND2_X1 U9780 ( .A1(n8902), .A2(n9276), .ZN(n8102) );
  NAND2_X1 U9781 ( .A1(P2_U3151), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n8138) );
  OAI211_X1 U9782 ( .C1(n8103), .C2(n8905), .A(n8102), .B(n8138), .ZN(n8105)
         );
  INV_X1 U9783 ( .A(n8175), .ZN(n8217) );
  NOR2_X1 U9784 ( .A1(n8217), .A2(n8923), .ZN(n8104) );
  AOI211_X1 U9785 ( .C1(n8174), .C2(n8920), .A(n8105), .B(n8104), .ZN(n8106)
         );
  OAI21_X1 U9786 ( .B1(n8107), .B2(n8910), .A(n8106), .ZN(P2_U3157) );
  OAI222_X1 U9787 ( .A1(n8110), .A2(P1_U3086), .B1(n10134), .B2(n8109), .C1(
        n8108), .C2(n10128), .ZN(P1_U3335) );
  MUX2_X1 U9788 ( .A(n8160), .B(n8111), .S(n9383), .Z(n8112) );
  OAI21_X1 U9789 ( .B1(n8113), .B2(n9310), .A(n8112), .ZN(P2_U3468) );
  XNOR2_X1 U9790 ( .A(n8114), .B(n8118), .ZN(n10062) );
  OR2_X1 U9791 ( .A1(n7990), .A2(n8115), .ZN(n8117) );
  NAND2_X1 U9792 ( .A1(n8117), .A2(n8116), .ZN(n8119) );
  XNOR2_X1 U9793 ( .A(n8119), .B(n8118), .ZN(n8120) );
  OAI222_X1 U9794 ( .A1(n9960), .A2(n8320), .B1(n9962), .B2(n9961), .C1(n9916), 
        .C2(n8120), .ZN(n10059) );
  NAND2_X1 U9795 ( .A1(n10059), .A2(n9971), .ZN(n8126) );
  XNOR2_X1 U9796 ( .A(n7994), .B(n9551), .ZN(n8121) );
  NOR2_X1 U9797 ( .A1(n8121), .A2(n9952), .ZN(n10060) );
  NOR2_X1 U9798 ( .A1(n9551), .A2(n10227), .ZN(n8124) );
  OAI22_X1 U9799 ( .A1(n9971), .A2(n8122), .B1(n9546), .B2(n10221), .ZN(n8123)
         );
  AOI211_X1 U9800 ( .C1(n10060), .C2(n9944), .A(n8124), .B(n8123), .ZN(n8125)
         );
  OAI211_X1 U9801 ( .C1(n10062), .C2(n9929), .A(n8126), .B(n8125), .ZN(
        P1_U3281) );
  INV_X1 U9802 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n8133) );
  AOI21_X1 U9803 ( .B1(n10261), .B2(n8128), .A(n8127), .ZN(n8129) );
  OAI211_X1 U9804 ( .C1(n10265), .C2(n8131), .A(n8130), .B(n8129), .ZN(n8134)
         );
  NAND2_X1 U9805 ( .A1(n8134), .A2(n10283), .ZN(n8132) );
  OAI21_X1 U9806 ( .B1(n10283), .B2(n8133), .A(n8132), .ZN(P1_U3480) );
  NAND2_X1 U9807 ( .A1(n8134), .A2(n10291), .ZN(n8135) );
  OAI21_X1 U9808 ( .B1(n10291), .B2(n6454), .A(n8135), .ZN(P1_U3531) );
  XOR2_X1 U9809 ( .A(n8137), .B(n8136), .Z(n8154) );
  INV_X1 U9810 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n8139) );
  OAI21_X1 U9811 ( .B1(n8976), .B2(n8139), .A(n8138), .ZN(n8146) );
  OR3_X1 U9812 ( .A1(n8140), .A2(n8142), .A3(n8141), .ZN(n8143) );
  AOI21_X1 U9813 ( .B1(n8144), .B2(n8143), .A(n9060), .ZN(n8145) );
  AOI211_X1 U9814 ( .C1(n8985), .C2(n8147), .A(n8146), .B(n8145), .ZN(n8153)
         );
  NOR3_X1 U9815 ( .A1(n8148), .A2(n8150), .A3(n8149), .ZN(n8151) );
  OAI21_X1 U9816 ( .B1(n4406), .B2(n8151), .A(n9043), .ZN(n8152) );
  OAI211_X1 U9817 ( .C1(n8154), .C2(n9075), .A(n8153), .B(n8152), .ZN(P2_U3192) );
  AOI21_X1 U9818 ( .B1(n8156), .B2(n8155), .A(n8148), .ZN(n8170) );
  INV_X1 U9819 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n8158) );
  OAI21_X1 U9820 ( .B1(n8976), .B2(n8158), .A(n8157), .ZN(n8163) );
  AOI21_X1 U9821 ( .B1(n8160), .B2(n8159), .A(n8140), .ZN(n8161) );
  NOR2_X1 U9822 ( .A1(n8161), .A2(n9060), .ZN(n8162) );
  AOI211_X1 U9823 ( .C1(n8985), .C2(n8164), .A(n8163), .B(n8162), .ZN(n8169)
         );
  XNOR2_X1 U9824 ( .A(n8166), .B(n8165), .ZN(n8167) );
  NAND2_X1 U9825 ( .A1(n8167), .A2(n9066), .ZN(n8168) );
  OAI211_X1 U9826 ( .C1(n8170), .C2(n9086), .A(n8169), .B(n8168), .ZN(P2_U3191) );
  INV_X1 U9827 ( .A(n8171), .ZN(n8173) );
  MUX2_X1 U9828 ( .A(n8173), .B(n8172), .S(n9273), .Z(n8177) );
  AOI22_X1 U9829 ( .A1(n9300), .A2(n8175), .B1(n9299), .B2(n8174), .ZN(n8176)
         );
  OAI211_X1 U9830 ( .C1(n8179), .C2(n8178), .A(n8177), .B(n8176), .ZN(P2_U3223) );
  OAI21_X1 U9831 ( .B1(n8182), .B2(n8181), .A(n8180), .ZN(n8183) );
  NAND2_X1 U9832 ( .A1(n8183), .A2(n10211), .ZN(n8192) );
  OAI21_X1 U9833 ( .B1(n8186), .B2(n8185), .A(n8184), .ZN(n8190) );
  NAND2_X1 U9834 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U9835 ( .A1(n10141), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n8187) );
  OAI211_X1 U9836 ( .C1(n10215), .C2(n8188), .A(n9545), .B(n8187), .ZN(n8189)
         );
  AOI21_X1 U9837 ( .B1(n8190), .B2(n9716), .A(n8189), .ZN(n8191) );
  NAND2_X1 U9838 ( .A1(n8192), .A2(n8191), .ZN(P1_U3255) );
  AOI21_X1 U9839 ( .B1(n9378), .B2(n8210), .A(n8193), .ZN(n8195) );
  MUX2_X1 U9840 ( .A(n8961), .B(n8195), .S(n9383), .Z(n8194) );
  OAI21_X1 U9841 ( .B1(n8198), .B2(n9359), .A(n8194), .ZN(P2_U3470) );
  INV_X1 U9842 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n8196) );
  MUX2_X1 U9843 ( .A(n8196), .B(n8195), .S(n10298), .Z(n8197) );
  OAI21_X1 U9844 ( .B1(n8198), .B2(n9467), .A(n8197), .ZN(P2_U3423) );
  OAI22_X1 U9845 ( .A1(n8201), .A2(n8200), .B1(n8199), .B2(n8929), .ZN(n8205)
         );
  XNOR2_X1 U9846 ( .A(n8203), .B(n8202), .ZN(n8204) );
  XNOR2_X1 U9847 ( .A(n8205), .B(n8204), .ZN(n8212) );
  NAND2_X1 U9848 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8958) );
  OAI21_X1 U9849 ( .B1(n8918), .B2(n8293), .A(n8958), .ZN(n8206) );
  AOI21_X1 U9850 ( .B1(n8916), .B2(n8929), .A(n8206), .ZN(n8207) );
  OAI21_X1 U9851 ( .B1(n8208), .B2(n8655), .A(n8207), .ZN(n8209) );
  AOI21_X1 U9852 ( .B1(n8210), .B2(n8908), .A(n8209), .ZN(n8211) );
  OAI21_X1 U9853 ( .B1(n8212), .B2(n8910), .A(n8211), .ZN(P2_U3176) );
  INV_X1 U9854 ( .A(n8213), .ZN(n8239) );
  OAI222_X1 U9855 ( .A1(n9481), .A2(n8239), .B1(n4742), .B2(P2_U3151), .C1(
        n8214), .C2(n9494), .ZN(P2_U3274) );
  MUX2_X1 U9856 ( .A(n8693), .B(n8215), .S(n9383), .Z(n8216) );
  OAI21_X1 U9857 ( .B1(n8217), .B2(n9310), .A(n8216), .ZN(P2_U3469) );
  INV_X1 U9858 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9090) );
  NAND2_X1 U9859 ( .A1(n4300), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n8220) );
  INV_X1 U9860 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9388) );
  OR2_X1 U9861 ( .A1(n8218), .A2(n9388), .ZN(n8219) );
  OAI211_X1 U9862 ( .C1(n9090), .C2(n4298), .A(n8220), .B(n8219), .ZN(n8222)
         );
  INV_X1 U9863 ( .A(n8222), .ZN(n8223) );
  NAND2_X1 U9864 ( .A1(n8935), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n8225) );
  OAI21_X1 U9865 ( .B1(n8803), .B2(n8935), .A(n8225), .ZN(P2_U3522) );
  NAND2_X1 U9866 ( .A1(n4400), .A2(n8226), .ZN(n8256) );
  OAI21_X1 U9867 ( .B1(n4400), .B2(n8226), .A(n8256), .ZN(n8227) );
  NOR2_X1 U9868 ( .A1(n8227), .A2(n8228), .ZN(n8259) );
  AOI21_X1 U9869 ( .B1(n8228), .B2(n8227), .A(n8259), .ZN(n8237) );
  OAI21_X1 U9870 ( .B1(n9654), .B2(n8230), .A(n8229), .ZN(n8231) );
  AOI21_X1 U9871 ( .B1(n9652), .B2(n9675), .A(n8231), .ZN(n8232) );
  OAI21_X1 U9872 ( .B1(n9636), .B2(n8233), .A(n8232), .ZN(n8234) );
  AOI21_X1 U9873 ( .B1(n8235), .B2(n9659), .A(n8234), .ZN(n8236) );
  OAI21_X1 U9874 ( .B1(n8237), .B2(n9662), .A(n8236), .ZN(P1_U3221) );
  OAI222_X1 U9875 ( .A1(n10128), .A2(n8240), .B1(n10134), .B2(n8239), .C1(
        n8238), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U9876 ( .A1(n8242), .A2(n8241), .ZN(n8243) );
  XNOR2_X1 U9877 ( .A(n8243), .B(n8247), .ZN(n8280) );
  INV_X1 U9878 ( .A(n8280), .ZN(n8255) );
  NAND2_X1 U9879 ( .A1(n8245), .A2(n8244), .ZN(n8248) );
  INV_X1 U9880 ( .A(n9957), .ZN(n8246) );
  AOI21_X1 U9881 ( .B1(n8248), .B2(n8247), .A(n8246), .ZN(n8249) );
  OAI222_X1 U9882 ( .A1(n9960), .A2(n9610), .B1(n9962), .B2(n9655), .C1(n9916), 
        .C2(n8249), .ZN(n8278) );
  AOI211_X1 U9883 ( .C1(n5470), .C2(n8250), .A(n9952), .B(n9949), .ZN(n8279)
         );
  NAND2_X1 U9884 ( .A1(n8279), .A2(n9944), .ZN(n8252) );
  AOI22_X1 U9885 ( .A1(n4287), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n9612), .B2(
        n9922), .ZN(n8251) );
  OAI211_X1 U9886 ( .C1(n9615), .C2(n10227), .A(n8252), .B(n8251), .ZN(n8253)
         );
  AOI21_X1 U9887 ( .B1(n8278), .B2(n9971), .A(n8253), .ZN(n8254) );
  OAI21_X1 U9888 ( .B1(n8255), .B2(n9929), .A(n8254), .ZN(P1_U3280) );
  INV_X1 U9889 ( .A(n8256), .ZN(n8257) );
  NOR3_X1 U9890 ( .A1(n8259), .A2(n8258), .A3(n8257), .ZN(n8262) );
  INV_X1 U9891 ( .A(n8260), .ZN(n8261) );
  OAI21_X1 U9892 ( .B1(n8262), .B2(n8261), .A(n9621), .ZN(n8269) );
  OAI21_X1 U9893 ( .B1(n9654), .B2(n8264), .A(n8263), .ZN(n8267) );
  NOR2_X1 U9894 ( .A1(n9636), .A2(n8265), .ZN(n8266) );
  AOI211_X1 U9895 ( .C1(n9652), .C2(n9674), .A(n8267), .B(n8266), .ZN(n8268)
         );
  OAI211_X1 U9896 ( .C1(n8270), .C2(n9630), .A(n8269), .B(n8268), .ZN(P1_U3231) );
  OR2_X1 U9897 ( .A1(n8411), .A2(n4847), .ZN(n8559) );
  XOR2_X1 U9898 ( .A(n8271), .B(n8559), .Z(n8272) );
  AOI222_X1 U9899 ( .A1(n9295), .A2(n8272), .B1(n9257), .B2(n9290), .C1(n8928), 
        .C2(n9292), .ZN(n8313) );
  AOI22_X1 U9900 ( .A1(n8410), .A2(n8273), .B1(n9299), .B2(n8300), .ZN(n8274)
         );
  AOI21_X1 U9901 ( .B1(n8313), .B2(n8274), .A(n9273), .ZN(n8277) );
  XNOR2_X1 U9902 ( .A(n8275), .B(n8559), .ZN(n8316) );
  OAI22_X1 U9903 ( .A1(n8316), .A2(n9264), .B1(n8997), .B2(n9296), .ZN(n8276)
         );
  OR2_X1 U9904 ( .A1(n8277), .A2(n8276), .ZN(P2_U3220) );
  AOI211_X1 U9905 ( .C1(n10250), .C2(n8280), .A(n8279), .B(n8278), .ZN(n8285)
         );
  AOI22_X1 U9906 ( .A1(n5470), .A2(n8281), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n10289), .ZN(n8282) );
  OAI21_X1 U9907 ( .B1(n8285), .B2(n10289), .A(n8282), .ZN(P1_U3535) );
  AOI22_X1 U9908 ( .A1(n5470), .A2(n8283), .B1(P1_REG0_REG_13__SCAN_IN), .B2(
        n10282), .ZN(n8284) );
  OAI21_X1 U9909 ( .B1(n8285), .B2(n10282), .A(n8284), .ZN(P1_U3492) );
  INV_X1 U9910 ( .A(n8286), .ZN(n8288) );
  OAI222_X1 U9911 ( .A1(n10128), .A2(n8287), .B1(n10134), .B2(n8288), .C1(
        P1_U3086), .C2(n4590), .ZN(P1_U3333) );
  OAI222_X1 U9912 ( .A1(n9494), .A2(n8289), .B1(n9481), .B2(n8288), .C1(
        P2_U3151), .C2(n8415), .ZN(P2_U3273) );
  INV_X1 U9913 ( .A(n8410), .ZN(n8303) );
  XNOR2_X1 U9914 ( .A(n8410), .B(n8621), .ZN(n8290) );
  NOR2_X1 U9915 ( .A1(n8290), .A2(n9277), .ZN(n8328) );
  AOI21_X1 U9916 ( .B1(n8290), .B2(n9277), .A(n8328), .ZN(n8296) );
  INV_X1 U9917 ( .A(n8292), .ZN(n8294) );
  OAI21_X1 U9918 ( .B1(n8296), .B2(n8295), .A(n8331), .ZN(n8297) );
  NAND2_X1 U9919 ( .A1(n8297), .A2(n8912), .ZN(n8302) );
  NAND2_X1 U9920 ( .A1(n8916), .A2(n8928), .ZN(n8298) );
  NAND2_X1 U9921 ( .A1(P2_U3151), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n9000) );
  OAI211_X1 U9922 ( .C1(n8593), .C2(n8918), .A(n8298), .B(n9000), .ZN(n8299)
         );
  AOI21_X1 U9923 ( .B1(n8300), .B2(n8920), .A(n8299), .ZN(n8301) );
  OAI211_X1 U9924 ( .C1(n8303), .C2(n8923), .A(n8302), .B(n8301), .ZN(P2_U3174) );
  NAND2_X1 U9925 ( .A1(n8307), .A2(n10122), .ZN(n8305) );
  OAI211_X1 U9926 ( .C1(n8306), .C2(n10128), .A(n8305), .B(n8304), .ZN(
        P1_U3332) );
  NAND2_X1 U9927 ( .A1(n8307), .A2(n9482), .ZN(n8309) );
  OR2_X1 U9928 ( .A1(n8308), .A2(P2_U3151), .ZN(n8587) );
  OAI211_X1 U9929 ( .C1(n8722), .C2(n9494), .A(n8309), .B(n8587), .ZN(P2_U3272) );
  MUX2_X1 U9930 ( .A(n8310), .B(n8313), .S(n10298), .Z(n8312) );
  NAND2_X1 U9931 ( .A1(n8410), .A2(n9463), .ZN(n8311) );
  OAI211_X1 U9932 ( .C1(n8316), .C2(n9467), .A(n8312), .B(n8311), .ZN(P2_U3429) );
  MUX2_X1 U9933 ( .A(n9003), .B(n8313), .S(n9383), .Z(n8315) );
  NAND2_X1 U9934 ( .A1(n8410), .A2(n9356), .ZN(n8314) );
  OAI211_X1 U9935 ( .C1(n9359), .C2(n8316), .A(n8315), .B(n8314), .ZN(P2_U3472) );
  AOI21_X1 U9936 ( .B1(n8318), .B2(n8317), .A(n4398), .ZN(n8327) );
  OAI21_X1 U9937 ( .B1(n9643), .B2(n8320), .A(n8319), .ZN(n8321) );
  AOI21_X1 U9938 ( .B1(n9640), .B2(n9675), .A(n8321), .ZN(n8322) );
  OAI21_X1 U9939 ( .B1(n9636), .B2(n8323), .A(n8322), .ZN(n8324) );
  AOI21_X1 U9940 ( .B1(n8325), .B2(n9659), .A(n8324), .ZN(n8326) );
  OAI21_X1 U9941 ( .B1(n8327), .B2(n9662), .A(n8326), .ZN(P1_U3217) );
  INV_X1 U9942 ( .A(n8357), .ZN(n9266) );
  INV_X1 U9943 ( .A(n8328), .ZN(n8329) );
  XNOR2_X1 U9944 ( .A(n8357), .B(n7357), .ZN(n8592) );
  XNOR2_X1 U9945 ( .A(n8592), .B(n8593), .ZN(n8330) );
  AND3_X1 U9946 ( .A1(n8331), .A2(n8330), .A3(n8329), .ZN(n8332) );
  OAI21_X1 U9947 ( .B1(n8591), .B2(n8332), .A(n8912), .ZN(n8337) );
  NAND2_X1 U9948 ( .A1(n8916), .A2(n9277), .ZN(n8333) );
  NAND2_X1 U9949 ( .A1(P2_U3151), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n9017) );
  OAI211_X1 U9950 ( .C1(n8334), .C2(n8918), .A(n8333), .B(n9017), .ZN(n8335)
         );
  AOI21_X1 U9951 ( .B1(n9270), .B2(n8920), .A(n8335), .ZN(n8336) );
  OAI211_X1 U9952 ( .C1(n9266), .C2(n8923), .A(n8337), .B(n8336), .ZN(P2_U3155) );
  AOI211_X1 U9953 ( .C1(n8340), .C2(n8339), .A(n10158), .B(n8338), .ZN(n8349)
         );
  AOI211_X1 U9954 ( .C1(n8343), .C2(n8342), .A(n10206), .B(n8341), .ZN(n8348)
         );
  NAND2_X1 U9955 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9608) );
  INV_X1 U9956 ( .A(n9608), .ZN(n8344) );
  AOI21_X1 U9957 ( .B1(n10141), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n8344), .ZN(
        n8345) );
  OAI21_X1 U9958 ( .B1(n10215), .B2(n8346), .A(n8345), .ZN(n8347) );
  OR3_X1 U9959 ( .A1(n8349), .A2(n8348), .A3(n8347), .ZN(P1_U3256) );
  INV_X1 U9960 ( .A(n8472), .ZN(n8350) );
  OR2_X1 U9961 ( .A1(n8471), .A2(n8350), .ZN(n8474) );
  INV_X1 U9962 ( .A(n8474), .ZN(n8562) );
  XNOR2_X1 U9963 ( .A(n8351), .B(n8562), .ZN(n8352) );
  AOI222_X1 U9964 ( .A1(n9295), .A2(n8352), .B1(n9247), .B2(n9290), .C1(n9277), 
        .C2(n9292), .ZN(n9267) );
  MUX2_X1 U9965 ( .A(n8353), .B(n9267), .S(n10298), .Z(n8356) );
  XNOR2_X1 U9966 ( .A(n8354), .B(n8474), .ZN(n9271) );
  AOI22_X1 U9967 ( .A1(n9271), .A2(n9428), .B1(n9463), .B2(n8357), .ZN(n8355)
         );
  NAND2_X1 U9968 ( .A1(n8356), .A2(n8355), .ZN(P2_U3432) );
  MUX2_X1 U9969 ( .A(n8698), .B(n9267), .S(n9383), .Z(n8359) );
  AOI22_X1 U9970 ( .A1(n9271), .A2(n9332), .B1(n9356), .B2(n8357), .ZN(n8358)
         );
  NAND2_X1 U9971 ( .A1(n8359), .A2(n8358), .ZN(P2_U3473) );
  INV_X1 U9972 ( .A(n8360), .ZN(n8362) );
  NOR3_X1 U9973 ( .A1(n4398), .A2(n8362), .A3(n8361), .ZN(n8363) );
  OAI21_X1 U9974 ( .B1(n8363), .B2(n4399), .A(n9621), .ZN(n8369) );
  OAI21_X1 U9975 ( .B1(n9643), .B2(n9610), .A(n8364), .ZN(n8367) );
  NOR2_X1 U9976 ( .A1(n9636), .A2(n8365), .ZN(n8366) );
  AOI211_X1 U9977 ( .C1(n9640), .C2(n9674), .A(n8367), .B(n8366), .ZN(n8368)
         );
  OAI211_X1 U9978 ( .C1(n8370), .C2(n9630), .A(n8369), .B(n8368), .ZN(P1_U3236) );
  XNOR2_X1 U9979 ( .A(n8371), .B(n5834), .ZN(n10053) );
  INV_X1 U9980 ( .A(n8373), .ZN(n8374) );
  AOI21_X1 U9981 ( .B1(n8375), .B2(n8372), .A(n8374), .ZN(n8376) );
  OAI222_X1 U9982 ( .A1(n9960), .A2(n9655), .B1(n9962), .B2(n9918), .C1(n9916), 
        .C2(n8376), .ZN(n10049) );
  INV_X1 U9983 ( .A(n10051), .ZN(n8379) );
  AOI211_X1 U9984 ( .C1(n10051), .C2(n9950), .A(n9952), .B(n9937), .ZN(n10050)
         );
  NAND2_X1 U9985 ( .A1(n10050), .A2(n9944), .ZN(n8378) );
  AOI22_X1 U9986 ( .A1(n4287), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9657), .B2(
        n9922), .ZN(n8377) );
  OAI211_X1 U9987 ( .C1(n8379), .C2(n10227), .A(n8378), .B(n8377), .ZN(n8380)
         );
  AOI21_X1 U9988 ( .B1(n10049), .B2(n9971), .A(n8380), .ZN(n8381) );
  OAI21_X1 U9989 ( .B1(n10053), .B2(n9929), .A(n8381), .ZN(P1_U3278) );
  INV_X1 U9990 ( .A(n6973), .ZN(n8590) );
  OAI222_X1 U9991 ( .A1(n9496), .A2(n8590), .B1(P2_U3151), .B2(n7083), .C1(
        n8382), .C2(n9494), .ZN(P2_U3271) );
  INV_X1 U9992 ( .A(n8383), .ZN(n9488) );
  OAI222_X1 U9993 ( .A1(n10128), .A2(n8385), .B1(n10134), .B2(n9488), .C1(
        n8384), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U9994 ( .A(n8386), .ZN(n9480) );
  OAI222_X1 U9995 ( .A1(P1_U3086), .A2(n8388), .B1(n10134), .B2(n9480), .C1(
        n8387), .C2(n10128), .ZN(P1_U3326) );
  INV_X1 U9996 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10219) );
  INV_X1 U9997 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10199) );
  INV_X1 U9998 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8389) );
  AOI22_X1 U9999 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .B1(n10199), .B2(n8389), .ZN(n10317) );
  INV_X1 U10000 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10184) );
  INV_X1 U10001 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n8390) );
  AOI22_X1 U10002 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .B1(n10184), .B2(n8390), .ZN(n10320) );
  INV_X1 U10003 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n8391) );
  INV_X1 U10004 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U10005 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .B1(n8391), .B2(n10171), .ZN(n10323) );
  NOR2_X1 U10006 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n8392) );
  AOI21_X1 U10007 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n8392), .ZN(n10326) );
  NOR2_X1 U10008 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8393) );
  AOI21_X1 U10009 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n8393), .ZN(n10329) );
  NOR2_X1 U10010 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n8394) );
  AOI21_X1 U10011 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n8394), .ZN(n10332) );
  NOR2_X1 U10012 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n8395) );
  AOI21_X1 U10013 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n8395), .ZN(n10335) );
  NOR2_X1 U10014 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n8396) );
  AOI21_X1 U10015 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n8396), .ZN(n10338) );
  NOR2_X1 U10016 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n8397) );
  AOI21_X1 U10017 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n8397), .ZN(n10347) );
  NOR2_X1 U10018 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8398) );
  AOI21_X1 U10019 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n8398), .ZN(n10353) );
  NOR2_X1 U10020 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n8399) );
  AOI21_X1 U10021 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n8399), .ZN(n10350) );
  NOR2_X1 U10022 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n8400) );
  AOI21_X1 U10023 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n8400), .ZN(n10341) );
  NOR2_X1 U10024 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n8401) );
  AOI21_X1 U10025 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n8401), .ZN(n10344) );
  INV_X1 U10026 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10309) );
  INV_X1 U10027 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10308) );
  NOR2_X1 U10028 ( .A1(n10309), .A2(n10308), .ZN(n10307) );
  NOR2_X1 U10029 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10307), .ZN(n10303) );
  INV_X1 U10030 ( .A(n10303), .ZN(n10304) );
  NAND3_X1 U10031 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U10032 ( .A1(n10306), .A2(n10305), .ZN(n10302) );
  NAND2_X1 U10033 ( .A1(n10304), .A2(n10302), .ZN(n10356) );
  NAND2_X1 U10034 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n8402) );
  OAI21_X1 U10035 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n8402), .ZN(n10355) );
  NOR2_X1 U10036 ( .A1(n10356), .A2(n10355), .ZN(n10354) );
  AOI21_X1 U10037 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10354), .ZN(n10359) );
  NAND2_X1 U10038 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n8403) );
  OAI21_X1 U10039 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n8403), .ZN(n10358) );
  NOR2_X1 U10040 ( .A1(n10359), .A2(n10358), .ZN(n10357) );
  AOI21_X1 U10041 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10357), .ZN(n10362) );
  NOR2_X1 U10042 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n8404) );
  AOI21_X1 U10043 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n8404), .ZN(n10361) );
  NAND2_X1 U10044 ( .A1(n10362), .A2(n10361), .ZN(n10360) );
  OAI21_X1 U10045 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10360), .ZN(n10343) );
  NAND2_X1 U10046 ( .A1(n10344), .A2(n10343), .ZN(n10342) );
  OAI21_X1 U10047 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10342), .ZN(n10340) );
  NAND2_X1 U10048 ( .A1(n10341), .A2(n10340), .ZN(n10339) );
  OAI21_X1 U10049 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10339), .ZN(n10349) );
  NAND2_X1 U10050 ( .A1(n10350), .A2(n10349), .ZN(n10348) );
  OAI21_X1 U10051 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10348), .ZN(n10352) );
  NAND2_X1 U10052 ( .A1(n10353), .A2(n10352), .ZN(n10351) );
  OAI21_X1 U10053 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10351), .ZN(n10346) );
  NAND2_X1 U10054 ( .A1(n10347), .A2(n10346), .ZN(n10345) );
  OAI21_X1 U10055 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10345), .ZN(n10337) );
  NAND2_X1 U10056 ( .A1(n10338), .A2(n10337), .ZN(n10336) );
  OAI21_X1 U10057 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10336), .ZN(n10334) );
  NAND2_X1 U10058 ( .A1(n10335), .A2(n10334), .ZN(n10333) );
  OAI21_X1 U10059 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10333), .ZN(n10331) );
  NAND2_X1 U10060 ( .A1(n10332), .A2(n10331), .ZN(n10330) );
  OAI21_X1 U10061 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10330), .ZN(n10328) );
  NAND2_X1 U10062 ( .A1(n10329), .A2(n10328), .ZN(n10327) );
  OAI21_X1 U10063 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10327), .ZN(n10325) );
  NAND2_X1 U10064 ( .A1(n10326), .A2(n10325), .ZN(n10324) );
  OAI21_X1 U10065 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10324), .ZN(n10322) );
  NAND2_X1 U10066 ( .A1(n10323), .A2(n10322), .ZN(n10321) );
  OAI21_X1 U10067 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10321), .ZN(n10319) );
  NAND2_X1 U10068 ( .A1(n10320), .A2(n10319), .ZN(n10318) );
  OAI21_X1 U10069 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10318), .ZN(n10316) );
  NAND2_X1 U10070 ( .A1(n10317), .A2(n10316), .ZN(n10315) );
  OAI21_X1 U10071 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10315), .ZN(n8405) );
  OR2_X1 U10072 ( .A1(n10219), .A2(n8405), .ZN(n10313) );
  NAND2_X1 U10073 ( .A1(n10314), .A2(n10313), .ZN(n10310) );
  NAND2_X1 U10074 ( .A1(n10219), .A2(n8405), .ZN(n10312) );
  NAND2_X1 U10075 ( .A1(n10310), .A2(n10312), .ZN(n8407) );
  XNOR2_X1 U10076 ( .A(n5194), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n8406) );
  XNOR2_X1 U10077 ( .A(n8407), .B(n8406), .ZN(ADD_1068_U4) );
  INV_X1 U10078 ( .A(n8801), .ZN(n8539) );
  NAND2_X1 U10079 ( .A1(n8573), .A2(n8408), .ZN(n8538) );
  INV_X1 U10080 ( .A(n8409), .ZN(n8925) );
  NAND2_X1 U10081 ( .A1(n8801), .A2(n8925), .ZN(n8529) );
  AOI21_X1 U10082 ( .B1(n8529), .B2(n8537), .A(n4756), .ZN(n8528) );
  MUX2_X1 U10083 ( .A(n9277), .B(n8410), .S(n8515), .Z(n8468) );
  INV_X1 U10084 ( .A(n8468), .ZN(n8470) );
  INV_X1 U10085 ( .A(n7059), .ZN(n8413) );
  AOI211_X1 U10086 ( .C1(n8542), .C2(n8414), .A(n8515), .B(n8413), .ZN(n8417)
         );
  MUX2_X1 U10087 ( .A(n8418), .B(n7059), .S(n8515), .Z(n8419) );
  NAND2_X1 U10088 ( .A1(n8421), .A2(n8420), .ZN(n8425) );
  NAND2_X1 U10089 ( .A1(n8934), .A2(n8422), .ZN(n8423) );
  NAND2_X1 U10090 ( .A1(n8427), .A2(n8423), .ZN(n8424) );
  INV_X1 U10091 ( .A(n8426), .ZN(n8550) );
  INV_X1 U10092 ( .A(n8427), .ZN(n8429) );
  OAI211_X1 U10093 ( .C1(n8441), .C2(n8429), .A(n8444), .B(n8428), .ZN(n8437)
         );
  INV_X1 U10094 ( .A(n8430), .ZN(n8443) );
  INV_X1 U10095 ( .A(n8438), .ZN(n8432) );
  OAI21_X1 U10096 ( .B1(n8443), .B2(n8432), .A(n8431), .ZN(n8436) );
  NAND2_X1 U10097 ( .A1(n8434), .A2(n8433), .ZN(n8435) );
  NAND2_X1 U10098 ( .A1(n8451), .A2(n8450), .ZN(n8447) );
  OAI211_X1 U10099 ( .C1(n8441), .C2(n8440), .A(n8439), .B(n8438), .ZN(n8445)
         );
  OAI21_X1 U10100 ( .B1(n8448), .B2(n8447), .A(n8446), .ZN(n8455) );
  AND2_X1 U10101 ( .A1(n8450), .A2(n8449), .ZN(n8452) );
  OAI211_X1 U10102 ( .C1(n8453), .C2(n8452), .A(n8451), .B(n8457), .ZN(n8454)
         );
  MUX2_X1 U10103 ( .A(n8455), .B(n8454), .S(n8515), .Z(n8459) );
  MUX2_X1 U10104 ( .A(n8457), .B(n8456), .S(n8515), .Z(n8458) );
  INV_X1 U10105 ( .A(n8460), .ZN(n8461) );
  AOI21_X1 U10106 ( .B1(n8463), .B2(n8462), .A(n8461), .ZN(n8465) );
  NOR2_X1 U10107 ( .A1(n8465), .A2(n8561), .ZN(n8464) );
  MUX2_X1 U10108 ( .A(n8472), .B(n7071), .S(n8515), .Z(n8473) );
  XNOR2_X1 U10109 ( .A(n9464), .B(n9247), .ZN(n8563) );
  MUX2_X1 U10110 ( .A(n8475), .B(n4385), .S(n8515), .Z(n8476) );
  MUX2_X1 U10111 ( .A(n8479), .B(n8478), .S(n8515), .Z(n8480) );
  NAND3_X1 U10112 ( .A1(n8482), .A2(n8481), .A3(n8480), .ZN(n8485) );
  NAND3_X1 U10113 ( .A1(n8485), .A2(n8484), .A3(n9195), .ZN(n8486) );
  NAND2_X1 U10114 ( .A1(n8486), .A2(n8546), .ZN(n8487) );
  INV_X1 U10115 ( .A(n8493), .ZN(n8488) );
  NAND2_X1 U10116 ( .A1(n8492), .A2(n8491), .ZN(n8495) );
  INV_X1 U10117 ( .A(n9177), .ZN(n9170) );
  MUX2_X1 U10118 ( .A(n8498), .B(n8497), .S(n8515), .Z(n8499) );
  NAND2_X1 U10119 ( .A1(n8500), .A2(n9150), .ZN(n9157) );
  NAND2_X1 U10120 ( .A1(n8505), .A2(n8500), .ZN(n8503) );
  INV_X1 U10121 ( .A(n8501), .ZN(n8502) );
  MUX2_X1 U10122 ( .A(n8503), .B(n8502), .S(n8515), .Z(n8508) );
  INV_X1 U10123 ( .A(n8504), .ZN(n8510) );
  MUX2_X1 U10124 ( .A(n8506), .B(n8505), .S(n8515), .Z(n8507) );
  INV_X1 U10125 ( .A(n8517), .ZN(n8509) );
  MUX2_X1 U10126 ( .A(n8511), .B(n8510), .S(n8515), .Z(n8512) );
  INV_X1 U10127 ( .A(n8514), .ZN(n8516) );
  MUX2_X1 U10128 ( .A(n8517), .B(n8516), .S(n8515), .Z(n8518) );
  AND2_X1 U10129 ( .A1(n9105), .A2(n4756), .ZN(n8523) );
  NAND2_X1 U10130 ( .A1(n9397), .A2(n8641), .ZN(n8521) );
  MUX2_X1 U10131 ( .A(n8521), .B(n8520), .S(n4756), .Z(n8522) );
  INV_X1 U10132 ( .A(n8523), .ZN(n8524) );
  OAI211_X1 U10133 ( .C1(n8526), .C2(n4756), .A(n8525), .B(n8524), .ZN(n8527)
         );
  INV_X1 U10134 ( .A(n8529), .ZN(n8571) );
  NAND2_X1 U10135 ( .A1(n10123), .A2(n6785), .ZN(n8533) );
  OR2_X1 U10136 ( .A1(n4657), .A2(n7196), .ZN(n8532) );
  NOR2_X1 U10137 ( .A1(n9385), .A2(n8803), .ZN(n8572) );
  NAND2_X1 U10138 ( .A1(n9385), .A2(n8803), .ZN(n8579) );
  INV_X1 U10139 ( .A(n8534), .ZN(n8535) );
  INV_X1 U10140 ( .A(n8579), .ZN(n8536) );
  AOI21_X1 U10141 ( .B1(n8536), .B2(n4302), .A(n8587), .ZN(n8580) );
  INV_X1 U10142 ( .A(n9385), .ZN(n9311) );
  AOI211_X1 U10143 ( .C1(n9311), .C2(n8539), .A(n8538), .B(n8572), .ZN(n8540)
         );
  NAND2_X1 U10144 ( .A1(n8541), .A2(n8540), .ZN(n8544) );
  AOI21_X1 U10145 ( .B1(n8571), .B2(n9385), .A(n4742), .ZN(n8543) );
  NOR2_X1 U10146 ( .A1(n8547), .A2(n7491), .ZN(n8551) );
  AND4_X1 U10147 ( .A1(n8551), .A2(n8550), .A3(n8549), .A4(n8548), .ZN(n8552)
         );
  NAND4_X1 U10148 ( .A1(n8554), .A2(n9301), .A3(n8553), .A4(n8552), .ZN(n8557)
         );
  NOR4_X1 U10149 ( .A1(n8558), .A2(n8557), .A3(n8556), .A4(n8555), .ZN(n8560)
         );
  NAND4_X1 U10150 ( .A1(n8562), .A2(n8561), .A3(n8560), .A4(n8559), .ZN(n8564)
         );
  NOR4_X1 U10151 ( .A1(n9230), .A2(n8565), .A3(n8564), .A4(n9255), .ZN(n8566)
         );
  NAND4_X1 U10152 ( .A1(n9197), .A2(n9207), .A3(n9217), .A4(n8566), .ZN(n8567)
         );
  NOR4_X1 U10153 ( .A1(n9157), .A2(n9177), .A3(n9183), .A4(n8567), .ZN(n8568)
         );
  NAND4_X1 U10154 ( .A1(n9122), .A2(n9140), .A3(n9152), .A4(n8568), .ZN(n8569)
         );
  NOR4_X1 U10155 ( .A1(n8571), .A2(n8570), .A3(n9113), .A4(n8569), .ZN(n8575)
         );
  INV_X1 U10156 ( .A(n8572), .ZN(n8574) );
  AND4_X1 U10157 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n9100), .ZN(n8576)
         );
  NAND2_X1 U10158 ( .A1(n4302), .A2(n8581), .ZN(n8582) );
  NAND3_X1 U10159 ( .A1(n8585), .A2(n8584), .A3(n9487), .ZN(n8586) );
  OAI211_X1 U10160 ( .C1(n4743), .C2(n8587), .A(n8586), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8588) );
  XNOR2_X1 U10161 ( .A(n9427), .B(n7357), .ZN(n8650) );
  INV_X1 U10162 ( .A(n8650), .ZN(n8651) );
  XNOR2_X1 U10163 ( .A(n9346), .B(n7357), .ZN(n8602) );
  XNOR2_X1 U10164 ( .A(n9464), .B(n7357), .ZN(n8595) );
  XNOR2_X1 U10165 ( .A(n8595), .B(n9247), .ZN(n8914) );
  NAND2_X1 U10166 ( .A1(n8915), .A2(n8914), .ZN(n8913) );
  XNOR2_X1 U10167 ( .A(n9457), .B(n8621), .ZN(n8594) );
  NOR2_X1 U10168 ( .A1(n8594), .A2(n9258), .ZN(n8598) );
  AOI21_X1 U10169 ( .B1(n8594), .B2(n9258), .A(n8598), .ZN(n8848) );
  INV_X1 U10170 ( .A(n8595), .ZN(n8596) );
  NAND2_X1 U10171 ( .A1(n8596), .A2(n9247), .ZN(n8849) );
  AND2_X1 U10172 ( .A1(n8848), .A2(n8849), .ZN(n8597) );
  NAND2_X1 U10173 ( .A1(n8913), .A2(n8597), .ZN(n8847) );
  INV_X1 U10174 ( .A(n8598), .ZN(n8858) );
  NAND2_X1 U10175 ( .A1(n8599), .A2(n9220), .ZN(n8601) );
  INV_X1 U10176 ( .A(n8601), .ZN(n8891) );
  XNOR2_X1 U10177 ( .A(n8602), .B(n9208), .ZN(n8890) );
  XNOR2_X1 U10178 ( .A(n9443), .B(n8621), .ZN(n8603) );
  INV_X1 U10179 ( .A(n9221), .ZN(n8927) );
  NAND2_X1 U10180 ( .A1(n8603), .A2(n8927), .ZN(n8823) );
  XNOR2_X1 U10181 ( .A(n9339), .B(n7357), .ZN(n8604) );
  INV_X1 U10182 ( .A(n8604), .ZN(n8605) );
  XNOR2_X1 U10183 ( .A(n8607), .B(n9172), .ZN(n8833) );
  OAI21_X1 U10184 ( .B1(n8651), .B2(n9185), .A(n8652), .ZN(n8612) );
  INV_X1 U10185 ( .A(n8868), .ZN(n8608) );
  AOI22_X1 U10186 ( .A1(n8608), .A2(n9173), .B1(n8651), .B2(n9185), .ZN(n8610)
         );
  XNOR2_X1 U10187 ( .A(n9415), .B(n7357), .ZN(n8870) );
  INV_X1 U10188 ( .A(n8870), .ZN(n8615) );
  AOI21_X1 U10189 ( .B1(n8868), .B2(n8886), .A(n9159), .ZN(n8614) );
  NAND3_X1 U10190 ( .A1(n8868), .A2(n8886), .A3(n9159), .ZN(n8613) );
  XNOR2_X1 U10191 ( .A(n9409), .B(n8621), .ZN(n8618) );
  XNOR2_X1 U10192 ( .A(n8618), .B(n8906), .ZN(n8841) );
  INV_X1 U10193 ( .A(n8618), .ZN(n8619) );
  XNOR2_X1 U10194 ( .A(n9403), .B(n8621), .ZN(n8620) );
  XNOR2_X1 U10195 ( .A(n8620), .B(n9133), .ZN(n8901) );
  XNOR2_X1 U10196 ( .A(n9397), .B(n8621), .ZN(n8640) );
  NAND2_X1 U10197 ( .A1(n8640), .A2(n9124), .ZN(n8637) );
  OAI21_X1 U10198 ( .B1(n8640), .B2(n9124), .A(n8637), .ZN(n8623) );
  AOI21_X1 U10199 ( .B1(n8622), .B2(n8623), .A(n8910), .ZN(n8626) );
  INV_X1 U10200 ( .A(n8622), .ZN(n8625) );
  INV_X1 U10201 ( .A(n8623), .ZN(n8624) );
  NAND2_X1 U10202 ( .A1(n8626), .A2(n8648), .ZN(n8631) );
  AOI22_X1 U10203 ( .A1(n9110), .A2(n8920), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8627) );
  OAI21_X1 U10204 ( .B1(n8628), .B2(n8905), .A(n8627), .ZN(n8629) );
  AOI21_X1 U10205 ( .B1(n8902), .B2(n9105), .A(n8629), .ZN(n8630) );
  OAI211_X1 U10206 ( .C1(n8923), .C2(n9116), .A(n8631), .B(n8630), .ZN(
        P2_U3154) );
  INV_X1 U10207 ( .A(n8632), .ZN(n8821) );
  OAI222_X1 U10208 ( .A1(n10128), .A2(n8634), .B1(n10134), .B2(n8821), .C1(
        P1_U3086), .C2(n8633), .ZN(P1_U3325) );
  XNOR2_X1 U10209 ( .A(n9105), .B(n7357), .ZN(n8635) );
  XNOR2_X1 U10210 ( .A(n9391), .B(n8635), .ZN(n8643) );
  INV_X1 U10211 ( .A(n8643), .ZN(n8636) );
  NAND2_X1 U10212 ( .A1(n8636), .A2(n8912), .ZN(n8649) );
  NAND4_X1 U10213 ( .A1(n8648), .A2(n8912), .A3(n8637), .A4(n8643), .ZN(n8647)
         );
  AOI22_X1 U10214 ( .A1(n9098), .A2(n8920), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8639) );
  NAND2_X1 U10215 ( .A1(n9124), .A2(n8916), .ZN(n8638) );
  OAI211_X1 U10216 ( .C1(n8926), .C2(n8918), .A(n8639), .B(n8638), .ZN(n8645)
         );
  INV_X1 U10217 ( .A(n8640), .ZN(n8642) );
  NOR4_X1 U10218 ( .A1(n8643), .A2(n8642), .A3(n8910), .A4(n8641), .ZN(n8644)
         );
  AOI211_X1 U10219 ( .C1(n8908), .C2(n9391), .A(n8645), .B(n8644), .ZN(n8646)
         );
  OAI211_X1 U10220 ( .C1(n8649), .C2(n8648), .A(n8647), .B(n8646), .ZN(
        P2_U3160) );
  NOR2_X1 U10221 ( .A1(n8652), .A2(n8651), .ZN(n8653) );
  AOI21_X2 U10222 ( .B1(n8883), .B2(n9158), .A(n8653), .ZN(n8866) );
  INV_X1 U10223 ( .A(n9163), .ZN(n8656) );
  AOI22_X1 U10224 ( .A1(n9185), .A2(n8916), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8654) );
  OAI21_X1 U10225 ( .B1(n8656), .B2(n8655), .A(n8654), .ZN(n8657) );
  AOI21_X1 U10226 ( .B1(n8902), .B2(n9134), .A(n8657), .ZN(n8658) );
  OAI21_X1 U10227 ( .B1(n8659), .B2(n8923), .A(n8658), .ZN(n8660) );
  NAND3_X1 U10228 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), 
        .A3(P2_D_REG_14__SCAN_IN), .ZN(n8662) );
  NAND3_X1 U10229 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(P2_REG0_REG_15__SCAN_IN), 
        .A3(P2_REG1_REG_14__SCAN_IN), .ZN(n8661) );
  NOR4_X1 U10230 ( .A1(SI_1_), .A2(P2_REG1_REG_13__SCAN_IN), .A3(n8662), .A4(
        n8661), .ZN(n8799) );
  OR4_X1 U10231 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), 
        .A3(P2_REG1_REG_24__SCAN_IN), .A4(n9187), .ZN(n8691) );
  NOR3_X1 U10232 ( .A1(SI_31_), .A2(P2_WR_REG_SCAN_IN), .A3(n8748), .ZN(n8664)
         );
  NOR3_X1 U10233 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_REG1_REG_10__SCAN_IN), 
        .A3(n8777), .ZN(n8663) );
  NAND4_X1 U10234 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_REG2_REG_22__SCAN_IN), 
        .A3(n8664), .A4(n8663), .ZN(n8690) );
  INV_X1 U10235 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8699) );
  AND4_X1 U10236 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P2_REG1_REG_25__SCAN_IN), 
        .A3(n8699), .A4(n10171), .ZN(n8686) );
  INV_X1 U10237 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n8959) );
  AND2_X1 U10238 ( .A1(n8959), .A2(n10309), .ZN(n8685) );
  NAND4_X1 U10239 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(P2_REG1_REG_23__SCAN_IN), 
        .A3(P2_REG1_REG_10__SCAN_IN), .A4(P2_REG2_REG_8__SCAN_IN), .ZN(n8666)
         );
  NAND4_X1 U10240 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(P2_REG2_REG_11__SCAN_IN), 
        .A3(P2_REG0_REG_2__SCAN_IN), .A4(P2_REG1_REG_0__SCAN_IN), .ZN(n8665)
         );
  NOR2_X1 U10241 ( .A1(n8666), .A2(n8665), .ZN(n8674) );
  NAND4_X1 U10242 ( .A1(P1_REG1_REG_21__SCAN_IN), .A2(P1_REG1_REG_12__SCAN_IN), 
        .A3(n9486), .A4(n9478), .ZN(n8668) );
  NAND4_X1 U10243 ( .A1(P1_REG0_REG_15__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), 
        .A3(P1_REG0_REG_2__SCAN_IN), .A4(n6453), .ZN(n8667) );
  NOR2_X1 U10244 ( .A1(n8668), .A2(n8667), .ZN(n8673) );
  NAND4_X1 U10245 ( .A1(SI_22_), .A2(P1_DATAO_REG_19__SCAN_IN), .A3(n8811), 
        .A4(n8669), .ZN(n8671) );
  NAND3_X1 U10246 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_1__SCAN_IN), 
        .A3(n8722), .ZN(n8670) );
  NOR2_X1 U10247 ( .A1(n8671), .A2(n8670), .ZN(n8672) );
  INV_X1 U10248 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n8718) );
  NAND4_X1 U10249 ( .A1(n8674), .A2(n8673), .A3(n8672), .A4(n8718), .ZN(n8675)
         );
  NOR2_X1 U10250 ( .A1(P2_DATAO_REG_13__SCAN_IN), .A2(n8675), .ZN(n8676) );
  AND4_X1 U10251 ( .A1(n8676), .A2(P1_REG0_REG_8__SCAN_IN), .A3(n8745), .A4(
        P1_D_REG_1__SCAN_IN), .ZN(n8684) );
  INV_X1 U10252 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8731) );
  NAND4_X1 U10253 ( .A1(n8678), .A2(n6509), .A3(n8677), .A4(n8731), .ZN(n8682)
         );
  INV_X1 U10254 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8680) );
  NAND4_X1 U10255 ( .A1(n8680), .A2(n8679), .A3(P2_B_REG_SCAN_IN), .A4(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n8681) );
  NOR2_X1 U10256 ( .A1(n8682), .A2(n8681), .ZN(n8683) );
  NAND4_X1 U10257 ( .A1(n8686), .A2(n8685), .A3(n8684), .A4(n8683), .ZN(n8689)
         );
  INV_X1 U10258 ( .A(n8687), .ZN(n8688) );
  NOR4_X1 U10259 ( .A1(n8691), .A2(n8690), .A3(n8689), .A4(n8688), .ZN(n8798)
         );
  INV_X1 U10260 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n10234) );
  AOI22_X1 U10261 ( .A1(n10234), .A2(keyinput13), .B1(keyinput23), .B2(n8693), 
        .ZN(n8692) );
  OAI221_X1 U10262 ( .B1(n10234), .B2(keyinput13), .C1(n8693), .C2(keyinput23), 
        .A(n8692), .ZN(n8696) );
  INV_X1 U10263 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9462) );
  AOI22_X1 U10264 ( .A1(n9187), .A2(keyinput44), .B1(keyinput62), .B2(n9462), 
        .ZN(n8694) );
  OAI221_X1 U10265 ( .B1(n9187), .B2(keyinput44), .C1(n9462), .C2(keyinput62), 
        .A(n8694), .ZN(n8695) );
  NOR2_X1 U10266 ( .A1(n8696), .A2(n8695), .ZN(n8706) );
  AOI22_X1 U10267 ( .A1(n8699), .A2(keyinput15), .B1(keyinput51), .B2(n8698), 
        .ZN(n8697) );
  OAI221_X1 U10268 ( .B1(n8699), .B2(keyinput15), .C1(n8698), .C2(keyinput51), 
        .A(n8697), .ZN(n8704) );
  AOI22_X1 U10269 ( .A1(n8702), .A2(keyinput47), .B1(n8701), .B2(keyinput26), 
        .ZN(n8700) );
  OAI221_X1 U10270 ( .B1(n8702), .B2(keyinput47), .C1(n8701), .C2(keyinput26), 
        .A(n8700), .ZN(n8703) );
  NOR2_X1 U10271 ( .A1(n8704), .A2(n8703), .ZN(n8705) );
  AND2_X1 U10272 ( .A1(n8706), .A2(n8705), .ZN(n8729) );
  AOI22_X1 U10273 ( .A1(n10160), .A2(keyinput14), .B1(keyinput40), .B2(n8959), 
        .ZN(n8707) );
  OAI221_X1 U10274 ( .B1(n10160), .B2(keyinput14), .C1(n8959), .C2(keyinput40), 
        .A(n8707), .ZN(n8715) );
  AOI22_X1 U10275 ( .A1(n8710), .A2(keyinput36), .B1(keyinput45), .B2(n8709), 
        .ZN(n8708) );
  OAI221_X1 U10276 ( .B1(n8710), .B2(keyinput36), .C1(n8709), .C2(keyinput45), 
        .A(n8708), .ZN(n8714) );
  AOI22_X1 U10277 ( .A1(n9486), .A2(keyinput34), .B1(keyinput59), .B2(n8712), 
        .ZN(n8711) );
  OAI221_X1 U10278 ( .B1(n9486), .B2(keyinput34), .C1(n8712), .C2(keyinput59), 
        .A(n8711), .ZN(n8713) );
  NOR3_X1 U10279 ( .A1(n8715), .A2(n8714), .A3(n8713), .ZN(n8728) );
  AOI22_X1 U10280 ( .A1(n5259), .A2(keyinput63), .B1(n6453), .B2(keyinput24), 
        .ZN(n8716) );
  OAI221_X1 U10281 ( .B1(n5259), .B2(keyinput63), .C1(n6453), .C2(keyinput24), 
        .A(n8716), .ZN(n8720) );
  AOI22_X1 U10282 ( .A1(n9279), .A2(keyinput2), .B1(keyinput58), .B2(n8718), 
        .ZN(n8717) );
  OAI221_X1 U10283 ( .B1(n9279), .B2(keyinput2), .C1(n8718), .C2(keyinput58), 
        .A(n8717), .ZN(n8719) );
  NOR2_X1 U10284 ( .A1(n8720), .A2(n8719), .ZN(n8727) );
  AOI22_X1 U10285 ( .A1(n8722), .A2(keyinput38), .B1(keyinput1), .B2(n10306), 
        .ZN(n8721) );
  OAI221_X1 U10286 ( .B1(n8722), .B2(keyinput38), .C1(n10306), .C2(keyinput1), 
        .A(n8721), .ZN(n8725) );
  XNOR2_X1 U10287 ( .A(n8723), .B(keyinput20), .ZN(n8724) );
  NOR2_X1 U10288 ( .A1(n8725), .A2(n8724), .ZN(n8726) );
  NAND4_X1 U10289 ( .A1(n8729), .A2(n8728), .A3(n8727), .A4(n8726), .ZN(n8797)
         );
  AOI22_X1 U10290 ( .A1(n8731), .A2(keyinput19), .B1(keyinput30), .B2(n6724), 
        .ZN(n8730) );
  OAI221_X1 U10291 ( .B1(n8731), .B2(keyinput19), .C1(n6724), .C2(keyinput30), 
        .A(n8730), .ZN(n8737) );
  AOI22_X1 U10292 ( .A1(n8957), .A2(keyinput55), .B1(n9478), .B2(keyinput37), 
        .ZN(n8732) );
  OAI221_X1 U10293 ( .B1(n8957), .B2(keyinput55), .C1(n9478), .C2(keyinput37), 
        .A(n8732), .ZN(n8736) );
  XNOR2_X1 U10294 ( .A(keyinput43), .B(n8733), .ZN(n8735) );
  XNOR2_X1 U10295 ( .A(keyinput0), .B(n5934), .ZN(n8734) );
  OR4_X1 U10296 ( .A1(n8737), .A2(n8736), .A3(n8735), .A4(n8734), .ZN(n8743)
         );
  INV_X1 U10297 ( .A(P2_WR_REG_SCAN_IN), .ZN(n8739) );
  AOI22_X1 U10298 ( .A1(n5656), .A2(keyinput60), .B1(keyinput25), .B2(n8739), 
        .ZN(n8738) );
  OAI221_X1 U10299 ( .B1(n5656), .B2(keyinput60), .C1(n8739), .C2(keyinput25), 
        .A(n8738), .ZN(n8742) );
  AOI22_X1 U10300 ( .A1(n10171), .A2(keyinput21), .B1(n6600), .B2(keyinput18), 
        .ZN(n8740) );
  OAI221_X1 U10301 ( .B1(n10171), .B2(keyinput21), .C1(n6600), .C2(keyinput18), 
        .A(n8740), .ZN(n8741) );
  NOR3_X1 U10302 ( .A1(n8743), .A2(n8742), .A3(n8741), .ZN(n8795) );
  AOI22_X1 U10303 ( .A1(n8745), .A2(keyinput49), .B1(keyinput56), .B2(n9003), 
        .ZN(n8744) );
  OAI221_X1 U10304 ( .B1(n8745), .B2(keyinput49), .C1(n9003), .C2(keyinput56), 
        .A(n8744), .ZN(n8756) );
  AOI22_X1 U10305 ( .A1(n5332), .A2(keyinput12), .B1(keyinput48), .B2(n9328), 
        .ZN(n8746) );
  OAI221_X1 U10306 ( .B1(n5332), .B2(keyinput12), .C1(n9328), .C2(keyinput48), 
        .A(n8746), .ZN(n8755) );
  AOI22_X1 U10307 ( .A1(n8749), .A2(keyinput53), .B1(n8748), .B2(keyinput35), 
        .ZN(n8747) );
  OAI221_X1 U10308 ( .B1(n8749), .B2(keyinput53), .C1(n8748), .C2(keyinput35), 
        .A(n8747), .ZN(n8754) );
  XOR2_X1 U10309 ( .A(n5359), .B(keyinput29), .Z(n8752) );
  XNOR2_X1 U10310 ( .A(SI_1_), .B(keyinput6), .ZN(n8751) );
  XNOR2_X1 U10311 ( .A(P2_B_REG_SCAN_IN), .B(keyinput5), .ZN(n8750) );
  NAND3_X1 U10312 ( .A1(n8752), .A2(n8751), .A3(n8750), .ZN(n8753) );
  NOR4_X1 U10313 ( .A1(n8756), .A2(n8755), .A3(n8754), .A4(n8753), .ZN(n8794)
         );
  AOI22_X1 U10314 ( .A1(n10309), .A2(keyinput3), .B1(n8758), .B2(keyinput61), 
        .ZN(n8757) );
  OAI221_X1 U10315 ( .B1(n10309), .B2(keyinput3), .C1(n8758), .C2(keyinput61), 
        .A(n8757), .ZN(n8774) );
  XNOR2_X1 U10316 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(keyinput10), .ZN(n8762)
         );
  XNOR2_X1 U10317 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput7), .ZN(n8761) );
  XNOR2_X1 U10318 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput11), .ZN(n8760) );
  XNOR2_X1 U10319 ( .A(SI_4_), .B(keyinput42), .ZN(n8759) );
  NAND4_X1 U10320 ( .A1(n8762), .A2(n8761), .A3(n8760), .A4(n8759), .ZN(n8773)
         );
  XNOR2_X1 U10321 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput41), .ZN(n8766) );
  XNOR2_X1 U10322 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput4), .ZN(n8765) );
  XNOR2_X1 U10323 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput17), .ZN(n8764)
         );
  XNOR2_X1 U10324 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(keyinput33), .ZN(n8763) );
  NAND4_X1 U10325 ( .A1(n8766), .A2(n8765), .A3(n8764), .A4(n8763), .ZN(n8772)
         );
  XNOR2_X1 U10326 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput57), .ZN(n8770)
         );
  XNOR2_X1 U10327 ( .A(P2_REG1_REG_24__SCAN_IN), .B(keyinput32), .ZN(n8769) );
  XNOR2_X1 U10328 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput52), .ZN(n8768) );
  XNOR2_X1 U10329 ( .A(P2_REG2_REG_15__SCAN_IN), .B(keyinput22), .ZN(n8767) );
  NAND4_X1 U10330 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n8771)
         );
  NOR4_X1 U10331 ( .A1(n8774), .A2(n8773), .A3(n8772), .A4(n8771), .ZN(n8793)
         );
  AOI22_X1 U10332 ( .A1(n9322), .A2(keyinput46), .B1(keyinput50), .B2(n6749), 
        .ZN(n8775) );
  OAI221_X1 U10333 ( .B1(n9322), .B2(keyinput46), .C1(n6749), .C2(keyinput50), 
        .A(n8775), .ZN(n8783) );
  AOI22_X1 U10334 ( .A1(n8778), .A2(keyinput31), .B1(keyinput8), .B2(n8777), 
        .ZN(n8776) );
  OAI221_X1 U10335 ( .B1(n8778), .B2(keyinput31), .C1(n8777), .C2(keyinput8), 
        .A(n8776), .ZN(n8782) );
  AOI22_X1 U10336 ( .A1(n8780), .A2(keyinput28), .B1(n8811), .B2(keyinput16), 
        .ZN(n8779) );
  OAI221_X1 U10337 ( .B1(n8780), .B2(keyinput28), .C1(n8811), .C2(keyinput16), 
        .A(n8779), .ZN(n8781) );
  OR3_X1 U10338 ( .A1(n8783), .A2(n8782), .A3(n8781), .ZN(n8791) );
  AOI22_X1 U10339 ( .A1(n8785), .A2(keyinput27), .B1(keyinput9), .B2(n6509), 
        .ZN(n8784) );
  OAI221_X1 U10340 ( .B1(n8785), .B2(keyinput27), .C1(n6509), .C2(keyinput9), 
        .A(n8784), .ZN(n8790) );
  INV_X1 U10341 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8788) );
  AOI22_X1 U10342 ( .A1(n8788), .A2(keyinput39), .B1(keyinput54), .B2(n8787), 
        .ZN(n8786) );
  OAI221_X1 U10343 ( .B1(n8788), .B2(keyinput39), .C1(n8787), .C2(keyinput54), 
        .A(n8786), .ZN(n8789) );
  NOR3_X1 U10344 ( .A1(n8791), .A2(n8790), .A3(n8789), .ZN(n8792) );
  NAND4_X1 U10345 ( .A1(n8795), .A2(n8794), .A3(n8793), .A4(n8792), .ZN(n8796)
         );
  AOI211_X1 U10346 ( .C1(n8799), .C2(n8798), .A(n8797), .B(n8796), .ZN(n8800)
         );
  NAND2_X1 U10347 ( .A1(n10301), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n8804) );
  NAND2_X1 U10348 ( .A1(n8808), .A2(n10298), .ZN(n9386) );
  OAI211_X1 U10349 ( .C1(n8801), .C2(n8805), .A(n8804), .B(n9386), .ZN(
        P2_U3457) );
  NAND2_X1 U10350 ( .A1(n9307), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U10351 ( .A1(n8808), .A2(n9383), .ZN(n9309) );
  OAI211_X1 U10352 ( .C1(n8801), .C2(n9310), .A(n8806), .B(n9309), .ZN(
        P2_U3489) );
  NOR2_X1 U10353 ( .A1(n8807), .A2(n9238), .ZN(n8815) );
  AOI21_X1 U10354 ( .B1(n8808), .B2(n9296), .A(n8815), .ZN(n9088) );
  NAND2_X1 U10355 ( .A1(n9273), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8809) );
  OAI211_X1 U10356 ( .C1(n8801), .C2(n9115), .A(n9088), .B(n8809), .ZN(
        P2_U3203) );
  OAI222_X1 U10357 ( .A1(n10128), .A2(n8811), .B1(n10134), .B2(n8810), .C1(
        P1_U3086), .C2(n9871), .ZN(P1_U3336) );
  INV_X1 U10358 ( .A(n8812), .ZN(n8819) );
  NOR2_X1 U10359 ( .A1(n8813), .A2(n9115), .ZN(n8814) );
  AOI211_X1 U10360 ( .C1(n9273), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8815), .B(
        n8814), .ZN(n8818) );
  NAND2_X1 U10361 ( .A1(n8816), .A2(n9303), .ZN(n8817) );
  OAI211_X1 U10362 ( .C1(n8819), .C2(n9273), .A(n8818), .B(n8817), .ZN(
        P2_U3204) );
  OAI222_X1 U10363 ( .A1(n9494), .A2(n8822), .B1(n9496), .B2(n8821), .C1(
        P2_U3151), .C2(n8820), .ZN(P2_U3265) );
  NAND2_X1 U10364 ( .A1(n4404), .A2(n8823), .ZN(n8824) );
  XNOR2_X1 U10365 ( .A(n8825), .B(n8824), .ZN(n8832) );
  AOI21_X1 U10366 ( .B1(n8916), .B2(n9208), .A(n8826), .ZN(n8828) );
  NAND2_X1 U10367 ( .A1(n8920), .A2(n9212), .ZN(n8827) );
  OAI211_X1 U10368 ( .C1(n8829), .C2(n8918), .A(n8828), .B(n8827), .ZN(n8830)
         );
  AOI21_X1 U10369 ( .B1(n9443), .B2(n8908), .A(n8830), .ZN(n8831) );
  OAI21_X1 U10370 ( .B1(n8832), .B2(n8910), .A(n8831), .ZN(P2_U3159) );
  XOR2_X1 U10371 ( .A(n8834), .B(n8833), .Z(n8839) );
  AOI22_X1 U10372 ( .A1(n9209), .A2(n8916), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8836) );
  NAND2_X1 U10373 ( .A1(n9188), .A2(n8920), .ZN(n8835) );
  OAI211_X1 U10374 ( .C1(n9158), .C2(n8918), .A(n8836), .B(n8835), .ZN(n8837)
         );
  AOI21_X1 U10375 ( .B1(n8606), .B2(n8908), .A(n8837), .ZN(n8838) );
  OAI21_X1 U10376 ( .B1(n8839), .B2(n8910), .A(n8838), .ZN(P2_U3163) );
  XOR2_X1 U10377 ( .A(n8841), .B(n8840), .Z(n8846) );
  NAND2_X1 U10378 ( .A1(n9133), .A2(n8902), .ZN(n8843) );
  AOI22_X1 U10379 ( .A1(n9138), .A2(n8920), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8842) );
  OAI211_X1 U10380 ( .C1(n9159), .C2(n8905), .A(n8843), .B(n8842), .ZN(n8844)
         );
  AOI21_X1 U10381 ( .B1(n9409), .B2(n8908), .A(n8844), .ZN(n8845) );
  OAI21_X1 U10382 ( .B1(n8846), .B2(n8910), .A(n8845), .ZN(P2_U3165) );
  INV_X1 U10383 ( .A(n9457), .ZN(n8856) );
  INV_X1 U10384 ( .A(n8859), .ZN(n8851) );
  AOI21_X1 U10385 ( .B1(n8913), .B2(n8849), .A(n8848), .ZN(n8850) );
  OAI21_X1 U10386 ( .B1(n8851), .B2(n8850), .A(n8912), .ZN(n8855) );
  NAND2_X1 U10387 ( .A1(n8916), .A2(n9247), .ZN(n8852) );
  NAND2_X1 U10388 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n9056) );
  OAI211_X1 U10389 ( .C1(n9220), .C2(n8918), .A(n8852), .B(n9056), .ZN(n8853)
         );
  AOI21_X1 U10390 ( .B1(n9251), .B2(n8920), .A(n8853), .ZN(n8854) );
  OAI211_X1 U10391 ( .C1(n8856), .C2(n8923), .A(n8855), .B(n8854), .ZN(
        P2_U3166) );
  INV_X1 U10392 ( .A(n9350), .ZN(n8865) );
  AND3_X1 U10393 ( .A1(n8859), .A2(n8858), .A3(n8857), .ZN(n8860) );
  OAI21_X1 U10394 ( .B1(n8892), .B2(n8860), .A(n8912), .ZN(n8864) );
  NAND2_X1 U10395 ( .A1(n8902), .A2(n9208), .ZN(n8861) );
  NAND2_X1 U10396 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n9078) );
  OAI211_X1 U10397 ( .C1(n9235), .C2(n8905), .A(n8861), .B(n9078), .ZN(n8862)
         );
  AOI21_X1 U10398 ( .B1(n9237), .B2(n8920), .A(n8862), .ZN(n8863) );
  OAI211_X1 U10399 ( .C1(n8865), .C2(n8923), .A(n8864), .B(n8863), .ZN(
        P2_U3168) );
  INV_X1 U10400 ( .A(n8866), .ZN(n8867) );
  XNOR2_X1 U10401 ( .A(n8870), .B(n9134), .ZN(n8871) );
  XNOR2_X1 U10402 ( .A(n8872), .B(n8871), .ZN(n8877) );
  NOR2_X1 U10403 ( .A1(n8906), .A2(n8918), .ZN(n8875) );
  AOI22_X1 U10404 ( .A1(n9149), .A2(n8920), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8873) );
  OAI21_X1 U10405 ( .B1(n8886), .B2(n8905), .A(n8873), .ZN(n8874) );
  AOI211_X1 U10406 ( .C1(n9415), .C2(n8908), .A(n8875), .B(n8874), .ZN(n8876)
         );
  OAI21_X1 U10407 ( .B1(n8877), .B2(n8910), .A(n8876), .ZN(P2_U3169) );
  AOI22_X1 U10408 ( .A1(n9172), .A2(n8902), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8879) );
  NAND2_X1 U10409 ( .A1(n8920), .A2(n9199), .ZN(n8878) );
  OAI211_X1 U10410 ( .C1(n9221), .C2(n8905), .A(n8879), .B(n8878), .ZN(n8880)
         );
  AOI21_X1 U10411 ( .B1(n9339), .B2(n8908), .A(n8880), .ZN(n8881) );
  OAI21_X1 U10412 ( .B1(n8882), .B2(n8910), .A(n8881), .ZN(P2_U3173) );
  XNOR2_X1 U10413 ( .A(n8883), .B(n9185), .ZN(n8889) );
  AOI22_X1 U10414 ( .A1(n9172), .A2(n8916), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8885) );
  NAND2_X1 U10415 ( .A1(n9176), .A2(n8920), .ZN(n8884) );
  OAI211_X1 U10416 ( .C1(n8886), .C2(n8918), .A(n8885), .B(n8884), .ZN(n8887)
         );
  AOI21_X1 U10417 ( .B1(n9427), .B2(n8908), .A(n8887), .ZN(n8888) );
  OAI21_X1 U10418 ( .B1(n8889), .B2(n8910), .A(n8888), .ZN(P2_U3175) );
  INV_X1 U10419 ( .A(n9346), .ZN(n8899) );
  NOR3_X1 U10420 ( .A1(n8892), .A2(n8891), .A3(n8890), .ZN(n8893) );
  OAI21_X1 U10421 ( .B1(n4345), .B2(n8893), .A(n8912), .ZN(n8898) );
  NAND2_X1 U10422 ( .A1(n8916), .A2(n9248), .ZN(n8895) );
  OAI211_X1 U10423 ( .C1(n9221), .C2(n8918), .A(n8895), .B(n8894), .ZN(n8896)
         );
  AOI21_X1 U10424 ( .B1(n9222), .B2(n8920), .A(n8896), .ZN(n8897) );
  OAI211_X1 U10425 ( .C1(n8899), .C2(n8923), .A(n8898), .B(n8897), .ZN(
        P2_U3178) );
  XOR2_X1 U10426 ( .A(n8901), .B(n8900), .Z(n8911) );
  NAND2_X1 U10427 ( .A1(n9124), .A2(n8902), .ZN(n8904) );
  AOI22_X1 U10428 ( .A1(n9127), .A2(n8920), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8903) );
  OAI211_X1 U10429 ( .C1(n8906), .C2(n8905), .A(n8904), .B(n8903), .ZN(n8907)
         );
  AOI21_X1 U10430 ( .B1(n9403), .B2(n8908), .A(n8907), .ZN(n8909) );
  OAI21_X1 U10431 ( .B1(n8911), .B2(n8910), .A(n8909), .ZN(P2_U3180) );
  INV_X1 U10432 ( .A(n9464), .ZN(n8924) );
  OAI211_X1 U10433 ( .C1(n8915), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8922)
         );
  NAND2_X1 U10434 ( .A1(n8916), .A2(n9257), .ZN(n8917) );
  NAND2_X1 U10435 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9036) );
  OAI211_X1 U10436 ( .C1(n9235), .C2(n8918), .A(n8917), .B(n9036), .ZN(n8919)
         );
  AOI21_X1 U10437 ( .B1(n9261), .B2(n8920), .A(n8919), .ZN(n8921) );
  OAI211_X1 U10438 ( .C1(n8924), .C2(n8923), .A(n8922), .B(n8921), .ZN(
        P2_U3181) );
  MUX2_X1 U10439 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8925), .S(P2_U3893), .Z(
        P2_U3521) );
  INV_X1 U10440 ( .A(n8926), .ZN(n9092) );
  MUX2_X1 U10441 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9092), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10442 ( .A(n9105), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8935), .Z(
        P2_U3519) );
  MUX2_X1 U10443 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9124), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10444 ( .A(n9133), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8935), .Z(
        P2_U3517) );
  MUX2_X1 U10445 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n9145), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10446 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9134), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10447 ( .A(n9173), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8935), .Z(
        P2_U3514) );
  MUX2_X1 U10448 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9185), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10449 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9172), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U10450 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9209), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U10451 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8927), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10452 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n9208), .S(P2_U3893), .Z(
        P2_U3509) );
  MUX2_X1 U10453 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9248), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U10454 ( .A(n9258), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8935), .Z(
        P2_U3507) );
  MUX2_X1 U10455 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9247), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U10456 ( .A(n9257), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8935), .Z(
        P2_U3505) );
  MUX2_X1 U10457 ( .A(n9277), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8935), .Z(
        P2_U3504) );
  MUX2_X1 U10458 ( .A(n8928), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8935), .Z(
        P2_U3503) );
  MUX2_X1 U10459 ( .A(n9276), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8935), .Z(
        P2_U3502) );
  MUX2_X1 U10460 ( .A(n8929), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8935), .Z(
        P2_U3501) );
  MUX2_X1 U10461 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8930), .S(P2_U3893), .Z(
        P2_U3500) );
  MUX2_X1 U10462 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9291), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U10463 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8931), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U10464 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n9293), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U10465 ( .A(n8932), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8935), .Z(
        P2_U3496) );
  MUX2_X1 U10466 ( .A(n8933), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8935), .Z(
        P2_U3494) );
  MUX2_X1 U10467 ( .A(n8934), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8935), .Z(
        P2_U3493) );
  MUX2_X1 U10468 ( .A(n4637), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8935), .Z(
        P2_U3492) );
  MUX2_X1 U10469 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n4627), .S(P2_U3893), .Z(
        P2_U3491) );
  OAI21_X1 U10470 ( .B1(n8939), .B2(n8938), .A(n8937), .ZN(n8940) );
  NAND2_X1 U10471 ( .A1(n8940), .A2(n9066), .ZN(n8955) );
  INV_X1 U10472 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8942) );
  OAI21_X1 U10473 ( .B1(n8976), .B2(n8942), .A(n8941), .ZN(n8943) );
  AOI21_X1 U10474 ( .B1(n8944), .B2(n8985), .A(n8943), .ZN(n8954) );
  AND3_X1 U10475 ( .A1(n7310), .A2(n8946), .A3(n8945), .ZN(n8947) );
  OAI21_X1 U10476 ( .B1(n8948), .B2(n8947), .A(n6685), .ZN(n8953) );
  AND3_X1 U10477 ( .A1(n7312), .A2(n8949), .A3(n5152), .ZN(n8950) );
  OAI21_X1 U10478 ( .B1(n8951), .B2(n8950), .A(n9043), .ZN(n8952) );
  NAND4_X1 U10479 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(
        P2_U3188) );
  AOI21_X1 U10480 ( .B1(n8957), .B2(n8956), .A(n4397), .ZN(n8971) );
  OAI21_X1 U10481 ( .B1(n8976), .B2(n8959), .A(n8958), .ZN(n8964) );
  AOI21_X1 U10482 ( .B1(n8961), .B2(n8960), .A(n8979), .ZN(n8962) );
  NOR2_X1 U10483 ( .A1(n8962), .A2(n9060), .ZN(n8963) );
  AOI211_X1 U10484 ( .C1(n8985), .C2(n8965), .A(n8964), .B(n8963), .ZN(n8970)
         );
  XNOR2_X1 U10485 ( .A(n8967), .B(n8966), .ZN(n8968) );
  NAND2_X1 U10486 ( .A1(n8968), .A2(n9066), .ZN(n8969) );
  OAI211_X1 U10487 ( .C1(n8971), .C2(n9086), .A(n8970), .B(n8969), .ZN(
        P2_U3193) );
  XOR2_X1 U10488 ( .A(n8973), .B(n8972), .Z(n8993) );
  INV_X1 U10489 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n8975) );
  OAI21_X1 U10490 ( .B1(n8976), .B2(n8975), .A(n8974), .ZN(n8983) );
  OR3_X1 U10491 ( .A1(n8979), .A2(n8978), .A3(n8977), .ZN(n8980) );
  AOI21_X1 U10492 ( .B1(n8981), .B2(n8980), .A(n9060), .ZN(n8982) );
  AOI211_X1 U10493 ( .C1(n8985), .C2(n8984), .A(n8983), .B(n8982), .ZN(n8992)
         );
  INV_X1 U10494 ( .A(n8986), .ZN(n8990) );
  NOR3_X1 U10495 ( .A1(n4397), .A2(n8988), .A3(n8987), .ZN(n8989) );
  OAI21_X1 U10496 ( .B1(n8990), .B2(n8989), .A(n9043), .ZN(n8991) );
  OAI211_X1 U10497 ( .C1(n8993), .C2(n9075), .A(n8992), .B(n8991), .ZN(
        P2_U3194) );
  INV_X1 U10498 ( .A(n8994), .ZN(n8995) );
  AOI21_X1 U10499 ( .B1(n8997), .B2(n8996), .A(n8995), .ZN(n9010) );
  XNOR2_X1 U10500 ( .A(n8999), .B(n8998), .ZN(n9008) );
  NAND2_X1 U10501 ( .A1(n9077), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n9001) );
  OAI211_X1 U10502 ( .C1(n9081), .C2(n9002), .A(n9001), .B(n9000), .ZN(n9007)
         );
  NAND2_X1 U10503 ( .A1(n9004), .A2(n9003), .ZN(n9005) );
  AOI21_X1 U10504 ( .B1(n9023), .B2(n9005), .A(n9060), .ZN(n9006) );
  AOI211_X1 U10505 ( .C1(n9066), .C2(n9008), .A(n9007), .B(n9006), .ZN(n9009)
         );
  OAI21_X1 U10506 ( .B1(n9010), .B2(n9086), .A(n9009), .ZN(P2_U3195) );
  INV_X1 U10507 ( .A(n9011), .ZN(n9013) );
  NOR2_X1 U10508 ( .A1(n9013), .A2(n9012), .ZN(n9014) );
  AOI21_X1 U10509 ( .B1(n9014), .B2(n8994), .A(n4409), .ZN(n9030) );
  XNOR2_X1 U10510 ( .A(n9016), .B(n9015), .ZN(n9028) );
  NAND2_X1 U10511 ( .A1(n9077), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n9018) );
  OAI211_X1 U10512 ( .C1(n9081), .C2(n9019), .A(n9018), .B(n9017), .ZN(n9027)
         );
  INV_X1 U10513 ( .A(n9020), .ZN(n9022) );
  NAND3_X1 U10514 ( .A1(n9023), .A2(n9022), .A3(n9021), .ZN(n9024) );
  AOI21_X1 U10515 ( .B1(n9025), .B2(n9024), .A(n9060), .ZN(n9026) );
  AOI211_X1 U10516 ( .C1(n9066), .C2(n9028), .A(n9027), .B(n9026), .ZN(n9029)
         );
  OAI21_X1 U10517 ( .B1(n9030), .B2(n9086), .A(n9029), .ZN(P2_U3196) );
  INV_X1 U10518 ( .A(n9031), .ZN(n9032) );
  AOI21_X1 U10519 ( .B1(n4956), .B2(n9033), .A(n9032), .ZN(n9047) );
  XNOR2_X1 U10520 ( .A(n9035), .B(n9034), .ZN(n9040) );
  NAND2_X1 U10521 ( .A1(n9077), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n9037) );
  OAI211_X1 U10522 ( .C1(n9081), .C2(n9038), .A(n9037), .B(n9036), .ZN(n9039)
         );
  AOI21_X1 U10523 ( .B1(n9040), .B2(n9066), .A(n9039), .ZN(n9046) );
  OAI21_X1 U10524 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n9042), .A(n9041), .ZN(
        n9044) );
  NAND2_X1 U10525 ( .A1(n9044), .A2(n9043), .ZN(n9045) );
  OAI211_X1 U10526 ( .C1(n9047), .C2(n9060), .A(n9046), .B(n9045), .ZN(
        P2_U3197) );
  INV_X1 U10527 ( .A(n9048), .ZN(n9050) );
  NOR2_X1 U10528 ( .A1(n9050), .A2(n9049), .ZN(n9053) );
  INV_X1 U10529 ( .A(n9051), .ZN(n9052) );
  AOI21_X1 U10530 ( .B1(n9053), .B2(n9041), .A(n9052), .ZN(n9068) );
  XNOR2_X1 U10531 ( .A(n9055), .B(n9054), .ZN(n9065) );
  NAND2_X1 U10532 ( .A1(n9077), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n9057) );
  OAI211_X1 U10533 ( .C1(n9081), .C2(n9058), .A(n9057), .B(n9056), .ZN(n9064)
         );
  NAND3_X1 U10534 ( .A1(n9031), .A2(n4418), .A3(n9059), .ZN(n9061) );
  AOI21_X1 U10535 ( .B1(n9062), .B2(n9061), .A(n9060), .ZN(n9063) );
  AOI211_X1 U10536 ( .C1(n9066), .C2(n9065), .A(n9064), .B(n9063), .ZN(n9067)
         );
  OAI21_X1 U10537 ( .B1(n9068), .B2(n9086), .A(n9067), .ZN(P2_U3198) );
  INV_X1 U10538 ( .A(n9069), .ZN(n9070) );
  AOI21_X1 U10539 ( .B1(n9240), .B2(n9071), .A(n9070), .ZN(n9087) );
  OAI21_X1 U10540 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9072), .A(n6688), .ZN(
        n9084) );
  XOR2_X1 U10541 ( .A(n9074), .B(n9073), .Z(n9076) );
  NOR2_X1 U10542 ( .A1(n9076), .A2(n9075), .ZN(n9083) );
  NAND2_X1 U10543 ( .A1(n9077), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n9079) );
  OAI211_X1 U10544 ( .C1(n9081), .C2(n9080), .A(n9079), .B(n9078), .ZN(n9082)
         );
  AOI211_X1 U10545 ( .C1(n9084), .C2(n6685), .A(n9083), .B(n9082), .ZN(n9085)
         );
  OAI21_X1 U10546 ( .B1(n9087), .B2(n9086), .A(n9085), .ZN(P2_U3199) );
  NAND2_X1 U10547 ( .A1(n9385), .A2(n9300), .ZN(n9089) );
  OAI211_X1 U10548 ( .C1(n9296), .C2(n9090), .A(n9089), .B(n9088), .ZN(
        P2_U3202) );
  XNOR2_X1 U10549 ( .A(n9091), .B(n9100), .ZN(n9096) );
  AOI21_X1 U10550 ( .B1(n9096), .B2(n9295), .A(n9095), .ZN(n9389) );
  AOI22_X1 U10551 ( .A1(n9391), .A2(n9300), .B1(n9299), .B2(n9098), .ZN(n9102)
         );
  XOR2_X1 U10552 ( .A(n9100), .B(n9099), .Z(n9392) );
  NAND2_X1 U10553 ( .A1(n9392), .A2(n9303), .ZN(n9101) );
  NAND3_X1 U10554 ( .A1(n9103), .A2(n9102), .A3(n9101), .ZN(P2_U3205) );
  XOR2_X1 U10555 ( .A(n9104), .B(n9113), .Z(n9109) );
  XOR2_X1 U10556 ( .A(n9113), .B(n9112), .Z(n9398) );
  OAI22_X1 U10557 ( .A1(n9116), .A2(n9115), .B1(n9114), .B2(n9296), .ZN(n9117)
         );
  AOI21_X1 U10558 ( .B1(n9398), .B2(n9303), .A(n9117), .ZN(n9118) );
  OAI21_X1 U10559 ( .B1(n9119), .B2(n9273), .A(n9118), .ZN(P2_U3206) );
  XNOR2_X1 U10560 ( .A(n9121), .B(n9120), .ZN(n9404) );
  INV_X1 U10561 ( .A(n9404), .ZN(n9130) );
  XNOR2_X1 U10562 ( .A(n9123), .B(n9122), .ZN(n9125) );
  AOI222_X1 U10563 ( .A1(n9295), .A2(n9125), .B1(n9124), .B2(n9290), .C1(n9145), .C2(n9292), .ZN(n9401) );
  MUX2_X1 U10564 ( .A(n9126), .B(n9401), .S(n9296), .Z(n9129) );
  AOI22_X1 U10565 ( .A1(n9403), .A2(n9300), .B1(n9299), .B2(n9127), .ZN(n9128)
         );
  OAI211_X1 U10566 ( .C1(n9130), .C2(n9264), .A(n9129), .B(n9128), .ZN(
        P2_U3207) );
  NOR2_X1 U10567 ( .A1(n9131), .A2(n9265), .ZN(n9137) );
  XOR2_X1 U10568 ( .A(n9140), .B(n9132), .Z(n9135) );
  AOI222_X1 U10569 ( .A1(n9295), .A2(n9135), .B1(n9134), .B2(n9292), .C1(n9133), .C2(n9290), .ZN(n9407) );
  INV_X1 U10570 ( .A(n9407), .ZN(n9136) );
  AOI211_X1 U10571 ( .C1(n9299), .C2(n9138), .A(n9137), .B(n9136), .ZN(n9142)
         );
  XNOR2_X1 U10572 ( .A(n9139), .B(n9140), .ZN(n9410) );
  AOI22_X1 U10573 ( .A1(n9410), .A2(n9303), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9273), .ZN(n9141) );
  OAI21_X1 U10574 ( .B1(n9142), .B2(n9273), .A(n9141), .ZN(P2_U3208) );
  INV_X1 U10575 ( .A(n9415), .ZN(n9143) );
  NOR2_X1 U10576 ( .A1(n9143), .A2(n9265), .ZN(n9148) );
  XNOR2_X1 U10577 ( .A(n9144), .B(n9152), .ZN(n9146) );
  AOI222_X1 U10578 ( .A1(n9295), .A2(n9146), .B1(n9173), .B2(n9292), .C1(n9145), .C2(n9290), .ZN(n9413) );
  INV_X1 U10579 ( .A(n9413), .ZN(n9147) );
  AOI211_X1 U10580 ( .C1(n9299), .C2(n9149), .A(n9148), .B(n9147), .ZN(n9155)
         );
  NAND2_X1 U10581 ( .A1(n9151), .A2(n9150), .ZN(n9153) );
  XNOR2_X1 U10582 ( .A(n9153), .B(n9152), .ZN(n9416) );
  AOI22_X1 U10583 ( .A1(n9416), .A2(n9303), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9273), .ZN(n9154) );
  OAI21_X1 U10584 ( .B1(n9155), .B2(n9273), .A(n9154), .ZN(P2_U3209) );
  XOR2_X1 U10585 ( .A(n9156), .B(n9157), .Z(n9422) );
  INV_X1 U10586 ( .A(n9422), .ZN(n9166) );
  INV_X1 U10587 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n9162) );
  XNOR2_X1 U10588 ( .A(n4331), .B(n4520), .ZN(n9161) );
  OAI22_X1 U10589 ( .A1(n9159), .A2(n9234), .B1(n9158), .B2(n9236), .ZN(n9160)
         );
  AOI21_X1 U10590 ( .B1(n9161), .B2(n9295), .A(n9160), .ZN(n9419) );
  MUX2_X1 U10591 ( .A(n9162), .B(n9419), .S(n9296), .Z(n9165) );
  AOI22_X1 U10592 ( .A1(n9421), .A2(n9300), .B1(n9299), .B2(n9163), .ZN(n9164)
         );
  OAI211_X1 U10593 ( .C1(n9166), .C2(n9264), .A(n9165), .B(n9164), .ZN(
        P2_U3210) );
  NAND2_X1 U10594 ( .A1(n9167), .A2(n9168), .ZN(n9184) );
  AOI21_X1 U10595 ( .B1(n9184), .B2(n9183), .A(n9169), .ZN(n9171) );
  XNOR2_X1 U10596 ( .A(n9171), .B(n9170), .ZN(n9174) );
  AOI222_X1 U10597 ( .A1(n9295), .A2(n9174), .B1(n9173), .B2(n9290), .C1(n9172), .C2(n9292), .ZN(n9425) );
  INV_X1 U10598 ( .A(n9425), .ZN(n9175) );
  AOI21_X1 U10599 ( .B1(n9299), .B2(n9176), .A(n9175), .ZN(n9181) );
  AOI22_X1 U10600 ( .A1(n9427), .A2(n9300), .B1(P2_REG2_REG_22__SCAN_IN), .B2(
        n9273), .ZN(n9180) );
  XNOR2_X1 U10601 ( .A(n9178), .B(n9177), .ZN(n9429) );
  NAND2_X1 U10602 ( .A1(n9429), .A2(n9303), .ZN(n9179) );
  OAI211_X1 U10603 ( .C1(n9181), .C2(n9273), .A(n9180), .B(n9179), .ZN(
        P2_U3211) );
  XNOR2_X1 U10604 ( .A(n9182), .B(n9183), .ZN(n9436) );
  XNOR2_X1 U10605 ( .A(n9184), .B(n9183), .ZN(n9186) );
  AOI222_X1 U10606 ( .A1(n9295), .A2(n9186), .B1(n9185), .B2(n9290), .C1(n9209), .C2(n9292), .ZN(n9432) );
  MUX2_X1 U10607 ( .A(n9187), .B(n9432), .S(n9296), .Z(n9190) );
  AOI22_X1 U10608 ( .A1(n8606), .A2(n9300), .B1(n9299), .B2(n9188), .ZN(n9189)
         );
  OAI211_X1 U10609 ( .C1(n9436), .C2(n9264), .A(n9190), .B(n9189), .ZN(
        P2_U3212) );
  INV_X1 U10610 ( .A(n9167), .ZN(n9191) );
  AOI21_X1 U10611 ( .B1(n9197), .B2(n9192), .A(n9191), .ZN(n9193) );
  OAI222_X1 U10612 ( .A1(n9236), .A2(n9221), .B1(n9234), .B2(n9194), .C1(n9231), .C2(n9193), .ZN(n9338) );
  NAND2_X1 U10613 ( .A1(n4314), .A2(n9217), .ZN(n9216) );
  NAND2_X1 U10614 ( .A1(n9216), .A2(n9195), .ZN(n9205) );
  NAND2_X1 U10615 ( .A1(n9205), .A2(n9207), .ZN(n9204) );
  NAND2_X1 U10616 ( .A1(n9204), .A2(n9196), .ZN(n9198) );
  XNOR2_X1 U10617 ( .A(n9198), .B(n9197), .ZN(n9440) );
  AOI22_X1 U10618 ( .A1(n9273), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9199), .B2(
        n9299), .ZN(n9201) );
  NAND2_X1 U10619 ( .A1(n9339), .A2(n9300), .ZN(n9200) );
  OAI211_X1 U10620 ( .C1(n9440), .C2(n9264), .A(n9201), .B(n9200), .ZN(n9202)
         );
  AOI21_X1 U10621 ( .B1(n9338), .B2(n9296), .A(n9202), .ZN(n9203) );
  INV_X1 U10622 ( .A(n9203), .ZN(P2_U3213) );
  OAI21_X1 U10623 ( .B1(n9205), .B2(n9207), .A(n9204), .ZN(n9446) );
  XOR2_X1 U10624 ( .A(n4280), .B(n9207), .Z(n9210) );
  AOI222_X1 U10625 ( .A1(n9295), .A2(n9210), .B1(n9209), .B2(n9290), .C1(n9208), .C2(n9292), .ZN(n9441) );
  MUX2_X1 U10626 ( .A(n9211), .B(n9441), .S(n9296), .Z(n9214) );
  AOI22_X1 U10627 ( .A1(n9443), .A2(n9300), .B1(n9299), .B2(n9212), .ZN(n9213)
         );
  OAI211_X1 U10628 ( .C1(n9446), .C2(n9264), .A(n9214), .B(n9213), .ZN(
        P2_U3214) );
  OR2_X1 U10629 ( .A1(n4314), .A2(n9217), .ZN(n9215) );
  NAND2_X1 U10630 ( .A1(n9216), .A2(n9215), .ZN(n9450) );
  XOR2_X1 U10631 ( .A(n9218), .B(n9217), .Z(n9219) );
  OAI222_X1 U10632 ( .A1(n9234), .A2(n9221), .B1(n9236), .B2(n9220), .C1(n9219), .C2(n9231), .ZN(n9345) );
  NAND2_X1 U10633 ( .A1(n9345), .A2(n9296), .ZN(n9227) );
  INV_X1 U10634 ( .A(n9222), .ZN(n9223) );
  OAI22_X1 U10635 ( .A1(n9296), .A2(n9224), .B1(n9223), .B2(n9238), .ZN(n9225)
         );
  AOI21_X1 U10636 ( .B1(n9346), .B2(n9300), .A(n9225), .ZN(n9226) );
  OAI211_X1 U10637 ( .C1(n9450), .C2(n9264), .A(n9227), .B(n9226), .ZN(
        P2_U3215) );
  XNOR2_X1 U10638 ( .A(n9228), .B(n9230), .ZN(n9454) );
  XNOR2_X1 U10639 ( .A(n9229), .B(n9230), .ZN(n9232) );
  OAI222_X1 U10640 ( .A1(n9236), .A2(n9235), .B1(n9234), .B2(n9233), .C1(n9232), .C2(n9231), .ZN(n9349) );
  NAND2_X1 U10641 ( .A1(n9349), .A2(n9296), .ZN(n9243) );
  INV_X1 U10642 ( .A(n9237), .ZN(n9239) );
  OAI22_X1 U10643 ( .A1(n9296), .A2(n9240), .B1(n9239), .B2(n9238), .ZN(n9241)
         );
  AOI21_X1 U10644 ( .B1(n9350), .B2(n9300), .A(n9241), .ZN(n9242) );
  OAI211_X1 U10645 ( .C1(n9454), .C2(n9264), .A(n9243), .B(n9242), .ZN(
        P2_U3216) );
  XNOR2_X1 U10646 ( .A(n9244), .B(n9245), .ZN(n9460) );
  XNOR2_X1 U10647 ( .A(n9246), .B(n9245), .ZN(n9249) );
  AOI222_X1 U10648 ( .A1(n9295), .A2(n9249), .B1(n9248), .B2(n9290), .C1(n9247), .C2(n9292), .ZN(n9455) );
  MUX2_X1 U10649 ( .A(n9250), .B(n9455), .S(n9296), .Z(n9253) );
  AOI22_X1 U10650 ( .A1(n9457), .A2(n9300), .B1(n9299), .B2(n9251), .ZN(n9252)
         );
  OAI211_X1 U10651 ( .C1(n9460), .C2(n9264), .A(n9253), .B(n9252), .ZN(
        P2_U3217) );
  XNOR2_X1 U10652 ( .A(n9254), .B(n9255), .ZN(n9468) );
  XNOR2_X1 U10653 ( .A(n4281), .B(n9255), .ZN(n9259) );
  AOI222_X1 U10654 ( .A1(n9295), .A2(n9259), .B1(n9258), .B2(n9290), .C1(n9257), .C2(n9292), .ZN(n9461) );
  MUX2_X1 U10655 ( .A(n9260), .B(n9461), .S(n9296), .Z(n9263) );
  AOI22_X1 U10656 ( .A1(n9464), .A2(n9300), .B1(n9299), .B2(n9261), .ZN(n9262)
         );
  OAI211_X1 U10657 ( .C1(n9468), .C2(n9264), .A(n9263), .B(n9262), .ZN(
        P2_U3218) );
  NOR2_X1 U10658 ( .A1(n9266), .A2(n9265), .ZN(n9269) );
  INV_X1 U10659 ( .A(n9267), .ZN(n9268) );
  AOI211_X1 U10660 ( .C1(n9299), .C2(n9270), .A(n9269), .B(n9268), .ZN(n9274)
         );
  AOI22_X1 U10661 ( .A1(n9271), .A2(n9303), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9273), .ZN(n9272) );
  OAI21_X1 U10662 ( .B1(n9274), .B2(n9273), .A(n9272), .ZN(P2_U3219) );
  XOR2_X1 U10663 ( .A(n9275), .B(n9283), .Z(n9278) );
  AOI222_X1 U10664 ( .A1(n9295), .A2(n9278), .B1(n9277), .B2(n9290), .C1(n9276), .C2(n9292), .ZN(n9362) );
  MUX2_X1 U10665 ( .A(n9279), .B(n9362), .S(n9296), .Z(n9286) );
  AOI22_X1 U10666 ( .A1(n7068), .A2(n9300), .B1(n9299), .B2(n9280), .ZN(n9285)
         );
  NAND2_X1 U10667 ( .A1(n9282), .A2(n9283), .ZN(n9360) );
  NAND3_X1 U10668 ( .A1(n9281), .A2(n9360), .A3(n9303), .ZN(n9284) );
  NAND3_X1 U10669 ( .A1(n9286), .A2(n9285), .A3(n9284), .ZN(P2_U3221) );
  INV_X1 U10670 ( .A(n9301), .ZN(n9288) );
  OAI21_X1 U10671 ( .B1(n9289), .B2(n9288), .A(n9287), .ZN(n9294) );
  AOI222_X1 U10672 ( .A1(n9295), .A2(n9294), .B1(n9293), .B2(n9292), .C1(n9291), .C2(n9290), .ZN(n9367) );
  MUX2_X1 U10673 ( .A(n9297), .B(n9367), .S(n9296), .Z(n9306) );
  AOI22_X1 U10674 ( .A1(n9300), .A2(n9364), .B1(n9299), .B2(n9298), .ZN(n9305)
         );
  OR2_X1 U10675 ( .A1(n9302), .A2(n9301), .ZN(n9365) );
  NAND3_X1 U10676 ( .A1(n9365), .A2(n9303), .A3(n7827), .ZN(n9304) );
  NAND3_X1 U10677 ( .A1(n9306), .A2(n9305), .A3(n9304), .ZN(P2_U3226) );
  NAND2_X1 U10678 ( .A1(n9307), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9308) );
  OAI211_X1 U10679 ( .C1(n9311), .C2(n9310), .A(n9309), .B(n9308), .ZN(
        P2_U3490) );
  INV_X1 U10680 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9312) );
  MUX2_X1 U10681 ( .A(n9312), .B(n9389), .S(n9383), .Z(n9314) );
  AOI22_X1 U10682 ( .A1(n9392), .A2(n9332), .B1(n9356), .B2(n9391), .ZN(n9313)
         );
  NAND2_X1 U10683 ( .A1(n9314), .A2(n9313), .ZN(P2_U3487) );
  OR2_X1 U10684 ( .A1(n9383), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n9315) );
  AOI22_X1 U10685 ( .A1(n9398), .A2(n9332), .B1(n9356), .B2(n9397), .ZN(n9317)
         );
  NAND2_X1 U10686 ( .A1(n9318), .A2(n9317), .ZN(P2_U3486) );
  INV_X1 U10687 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9319) );
  MUX2_X1 U10688 ( .A(n9319), .B(n9401), .S(n9383), .Z(n9321) );
  AOI22_X1 U10689 ( .A1(n9404), .A2(n9332), .B1(n9356), .B2(n9403), .ZN(n9320)
         );
  NAND2_X1 U10690 ( .A1(n9321), .A2(n9320), .ZN(P2_U3485) );
  MUX2_X1 U10691 ( .A(n9322), .B(n9407), .S(n9383), .Z(n9324) );
  AOI22_X1 U10692 ( .A1(n9410), .A2(n9332), .B1(n9356), .B2(n9409), .ZN(n9323)
         );
  NAND2_X1 U10693 ( .A1(n9324), .A2(n9323), .ZN(P2_U3484) );
  MUX2_X1 U10694 ( .A(n9325), .B(n9413), .S(n9383), .Z(n9327) );
  AOI22_X1 U10695 ( .A1(n9416), .A2(n9332), .B1(n9356), .B2(n9415), .ZN(n9326)
         );
  NAND2_X1 U10696 ( .A1(n9327), .A2(n9326), .ZN(P2_U3483) );
  MUX2_X1 U10697 ( .A(n9328), .B(n9419), .S(n9383), .Z(n9330) );
  AOI22_X1 U10698 ( .A1(n9422), .A2(n9332), .B1(n9356), .B2(n9421), .ZN(n9329)
         );
  NAND2_X1 U10699 ( .A1(n9330), .A2(n9329), .ZN(P2_U3482) );
  INV_X1 U10700 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9331) );
  MUX2_X1 U10701 ( .A(n9331), .B(n9425), .S(n9383), .Z(n9334) );
  AOI22_X1 U10702 ( .A1(n9429), .A2(n9332), .B1(n9356), .B2(n9427), .ZN(n9333)
         );
  NAND2_X1 U10703 ( .A1(n9334), .A2(n9333), .ZN(P2_U3481) );
  INV_X1 U10704 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9335) );
  MUX2_X1 U10705 ( .A(n9335), .B(n9432), .S(n9383), .Z(n9337) );
  NAND2_X1 U10706 ( .A1(n8606), .A2(n9356), .ZN(n9336) );
  OAI211_X1 U10707 ( .C1(n9359), .C2(n9436), .A(n9337), .B(n9336), .ZN(
        P2_U3480) );
  INV_X1 U10708 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9340) );
  AOI21_X1 U10709 ( .B1(n9378), .B2(n9339), .A(n9338), .ZN(n9437) );
  MUX2_X1 U10710 ( .A(n9340), .B(n9437), .S(n9383), .Z(n9341) );
  OAI21_X1 U10711 ( .B1(n9440), .B2(n9359), .A(n9341), .ZN(P2_U3479) );
  INV_X1 U10712 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9342) );
  MUX2_X1 U10713 ( .A(n9342), .B(n9441), .S(n9383), .Z(n9344) );
  NAND2_X1 U10714 ( .A1(n9443), .A2(n9356), .ZN(n9343) );
  OAI211_X1 U10715 ( .C1(n9359), .C2(n9446), .A(n9344), .B(n9343), .ZN(
        P2_U3478) );
  AOI21_X1 U10716 ( .B1(n9378), .B2(n9346), .A(n9345), .ZN(n9447) );
  MUX2_X1 U10717 ( .A(n9347), .B(n9447), .S(n9383), .Z(n9348) );
  OAI21_X1 U10718 ( .B1(n9359), .B2(n9450), .A(n9348), .ZN(P2_U3477) );
  INV_X1 U10719 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9351) );
  AOI21_X1 U10720 ( .B1(n9378), .B2(n9350), .A(n9349), .ZN(n9451) );
  MUX2_X1 U10721 ( .A(n9351), .B(n9451), .S(n9383), .Z(n9352) );
  OAI21_X1 U10722 ( .B1(n9454), .B2(n9359), .A(n9352), .ZN(P2_U3476) );
  MUX2_X1 U10723 ( .A(n9353), .B(n9455), .S(n9383), .Z(n9355) );
  NAND2_X1 U10724 ( .A1(n9457), .A2(n9356), .ZN(n9354) );
  OAI211_X1 U10725 ( .C1(n9460), .C2(n9359), .A(n9355), .B(n9354), .ZN(
        P2_U3475) );
  MUX2_X1 U10726 ( .A(n4956), .B(n9461), .S(n9383), .Z(n9358) );
  NAND2_X1 U10727 ( .A1(n9464), .A2(n9356), .ZN(n9357) );
  OAI211_X1 U10728 ( .C1(n9468), .C2(n9359), .A(n9358), .B(n9357), .ZN(
        P2_U3474) );
  NAND3_X1 U10729 ( .A1(n9281), .A2(n9360), .A3(n9376), .ZN(n9361) );
  OAI211_X1 U10730 ( .C1(n9363), .C2(n9368), .A(n9362), .B(n9361), .ZN(n9469)
         );
  MUX2_X1 U10731 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9469), .S(n9383), .Z(
        P2_U3471) );
  INV_X1 U10732 ( .A(n9364), .ZN(n9369) );
  NAND3_X1 U10733 ( .A1(n9365), .A2(n7827), .A3(n9376), .ZN(n9366) );
  OAI211_X1 U10734 ( .C1(n9369), .C2(n9368), .A(n9367), .B(n9366), .ZN(n9470)
         );
  MUX2_X1 U10735 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n9470), .S(n9383), .Z(
        P2_U3466) );
  NAND2_X1 U10736 ( .A1(n9370), .A2(n9376), .ZN(n9373) );
  NAND2_X1 U10737 ( .A1(n9371), .A2(n9378), .ZN(n9372) );
  INV_X1 U10738 ( .A(n10299), .ZN(n9375) );
  MUX2_X1 U10739 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n9375), .S(n9383), .Z(
        P2_U3465) );
  NAND2_X1 U10740 ( .A1(n9377), .A2(n9376), .ZN(n9381) );
  NAND2_X1 U10741 ( .A1(n9379), .A2(n9378), .ZN(n9380) );
  AND3_X1 U10742 ( .A1(n9382), .A2(n9381), .A3(n9380), .ZN(n10294) );
  INV_X1 U10743 ( .A(n10294), .ZN(n9384) );
  MUX2_X1 U10744 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n9384), .S(n9383), .Z(
        P2_U3462) );
  NAND2_X1 U10745 ( .A1(n9385), .A2(n9463), .ZN(n9387) );
  OAI211_X1 U10746 ( .C1(n10298), .C2(n9388), .A(n9387), .B(n9386), .ZN(
        P2_U3458) );
  INV_X1 U10747 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9390) );
  MUX2_X1 U10748 ( .A(n9390), .B(n9389), .S(n10298), .Z(n9394) );
  AOI22_X1 U10749 ( .A1(n9392), .A2(n9428), .B1(n9463), .B2(n9391), .ZN(n9393)
         );
  NAND2_X1 U10750 ( .A1(n9394), .A2(n9393), .ZN(P2_U3455) );
  INV_X1 U10751 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9396) );
  MUX2_X1 U10752 ( .A(n9396), .B(n9395), .S(n10298), .Z(n9400) );
  AOI22_X1 U10753 ( .A1(n9398), .A2(n9428), .B1(n9463), .B2(n9397), .ZN(n9399)
         );
  NAND2_X1 U10754 ( .A1(n9400), .A2(n9399), .ZN(P2_U3454) );
  INV_X1 U10755 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9402) );
  MUX2_X1 U10756 ( .A(n9402), .B(n9401), .S(n10298), .Z(n9406) );
  AOI22_X1 U10757 ( .A1(n9404), .A2(n9428), .B1(n9463), .B2(n9403), .ZN(n9405)
         );
  NAND2_X1 U10758 ( .A1(n9406), .A2(n9405), .ZN(P2_U3453) );
  INV_X1 U10759 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9408) );
  MUX2_X1 U10760 ( .A(n9408), .B(n9407), .S(n10298), .Z(n9412) );
  AOI22_X1 U10761 ( .A1(n9410), .A2(n9428), .B1(n9463), .B2(n9409), .ZN(n9411)
         );
  NAND2_X1 U10762 ( .A1(n9412), .A2(n9411), .ZN(P2_U3452) );
  INV_X1 U10763 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9414) );
  MUX2_X1 U10764 ( .A(n9414), .B(n9413), .S(n10298), .Z(n9418) );
  AOI22_X1 U10765 ( .A1(n9416), .A2(n9428), .B1(n9463), .B2(n9415), .ZN(n9417)
         );
  NAND2_X1 U10766 ( .A1(n9418), .A2(n9417), .ZN(P2_U3451) );
  INV_X1 U10767 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9420) );
  MUX2_X1 U10768 ( .A(n9420), .B(n9419), .S(n10298), .Z(n9424) );
  AOI22_X1 U10769 ( .A1(n9422), .A2(n9428), .B1(n9463), .B2(n9421), .ZN(n9423)
         );
  NAND2_X1 U10770 ( .A1(n9424), .A2(n9423), .ZN(P2_U3450) );
  INV_X1 U10771 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n9426) );
  MUX2_X1 U10772 ( .A(n9426), .B(n9425), .S(n10298), .Z(n9431) );
  AOI22_X1 U10773 ( .A1(n9429), .A2(n9428), .B1(n9463), .B2(n9427), .ZN(n9430)
         );
  NAND2_X1 U10774 ( .A1(n9431), .A2(n9430), .ZN(P2_U3449) );
  INV_X1 U10775 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9433) );
  MUX2_X1 U10776 ( .A(n9433), .B(n9432), .S(n10298), .Z(n9435) );
  NAND2_X1 U10777 ( .A1(n8606), .A2(n9463), .ZN(n9434) );
  OAI211_X1 U10778 ( .C1(n9436), .C2(n9467), .A(n9435), .B(n9434), .ZN(
        P2_U3448) );
  INV_X1 U10779 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9438) );
  MUX2_X1 U10780 ( .A(n9438), .B(n9437), .S(n10298), .Z(n9439) );
  OAI21_X1 U10781 ( .B1(n9440), .B2(n9467), .A(n9439), .ZN(P2_U3447) );
  INV_X1 U10782 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9442) );
  MUX2_X1 U10783 ( .A(n9442), .B(n9441), .S(n10298), .Z(n9445) );
  NAND2_X1 U10784 ( .A1(n9443), .A2(n9463), .ZN(n9444) );
  OAI211_X1 U10785 ( .C1(n9446), .C2(n9467), .A(n9445), .B(n9444), .ZN(
        P2_U3446) );
  INV_X1 U10786 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9448) );
  MUX2_X1 U10787 ( .A(n9448), .B(n9447), .S(n10298), .Z(n9449) );
  OAI21_X1 U10788 ( .B1(n9450), .B2(n9467), .A(n9449), .ZN(P2_U3444) );
  INV_X1 U10789 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9452) );
  MUX2_X1 U10790 ( .A(n9452), .B(n9451), .S(n10298), .Z(n9453) );
  OAI21_X1 U10791 ( .B1(n9454), .B2(n9467), .A(n9453), .ZN(P2_U3441) );
  INV_X1 U10792 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9456) );
  MUX2_X1 U10793 ( .A(n9456), .B(n9455), .S(n10298), .Z(n9459) );
  NAND2_X1 U10794 ( .A1(n9457), .A2(n9463), .ZN(n9458) );
  OAI211_X1 U10795 ( .C1(n9460), .C2(n9467), .A(n9459), .B(n9458), .ZN(
        P2_U3438) );
  MUX2_X1 U10796 ( .A(n9462), .B(n9461), .S(n10298), .Z(n9466) );
  NAND2_X1 U10797 ( .A1(n9464), .A2(n9463), .ZN(n9465) );
  OAI211_X1 U10798 ( .C1(n9468), .C2(n9467), .A(n9466), .B(n9465), .ZN(
        P2_U3435) );
  MUX2_X1 U10799 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9469), .S(n10298), .Z(
        P2_U3426) );
  MUX2_X1 U10800 ( .A(P2_REG0_REG_7__SCAN_IN), .B(n9470), .S(n10298), .Z(
        P2_U3411) );
  MUX2_X1 U10801 ( .A(n9472), .B(P2_D_REG_1__SCAN_IN), .S(n9471), .Z(P2_U3377)
         );
  NAND3_X1 U10802 ( .A1(n9474), .A2(P2_STATE_REG_SCAN_IN), .A3(
        P2_IR_REG_31__SCAN_IN), .ZN(n9475) );
  OAI22_X1 U10803 ( .A1(n9473), .A2(n9475), .B1(n7196), .B2(n9494), .ZN(n9476)
         );
  AOI21_X1 U10804 ( .B1(n10123), .B2(n9482), .A(n9476), .ZN(n9477) );
  INV_X1 U10805 ( .A(n9477), .ZN(P2_U3264) );
  OAI222_X1 U10806 ( .A1(n9481), .A2(n9480), .B1(n9479), .B2(P2_U3151), .C1(
        n9478), .C2(n9494), .ZN(P2_U3266) );
  NAND2_X1 U10807 ( .A1(n7021), .A2(n9482), .ZN(n9484) );
  OAI211_X1 U10808 ( .C1(n9490), .C2(n9485), .A(n9484), .B(n9483), .ZN(
        P2_U3267) );
  OAI222_X1 U10809 ( .A1(n9496), .A2(n9488), .B1(n9487), .B2(P2_U3151), .C1(
        n9486), .C2(n9494), .ZN(P2_U3268) );
  INV_X1 U10810 ( .A(n9489), .ZN(n10130) );
  OAI222_X1 U10811 ( .A1(n9496), .A2(n10130), .B1(P2_U3151), .B2(n9492), .C1(
        n9491), .C2(n9490), .ZN(P2_U3269) );
  INV_X1 U10812 ( .A(n9493), .ZN(n10133) );
  OAI222_X1 U10813 ( .A1(n9496), .A2(n10133), .B1(P2_U3151), .B2(n7085), .C1(
        n9495), .C2(n9494), .ZN(P2_U3270) );
  MUX2_X1 U10814 ( .A(n9497), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  INV_X1 U10815 ( .A(n9498), .ZN(n9503) );
  NOR2_X1 U10816 ( .A1(n9501), .A2(n9500), .ZN(n9561) );
  NAND2_X1 U10817 ( .A1(n9502), .A2(n9503), .ZN(n9563) );
  OAI21_X1 U10818 ( .B1(n9503), .B2(n9502), .A(n9563), .ZN(n9504) );
  NAND2_X1 U10819 ( .A1(n9504), .A2(n9621), .ZN(n9509) );
  INV_X1 U10820 ( .A(n9970), .ZN(n9507) );
  AND2_X1 U10821 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n10154) );
  AOI21_X1 U10822 ( .B1(n9640), .B2(n9672), .A(n10154), .ZN(n9505) );
  OAI21_X1 U10823 ( .B1(n9963), .B2(n9643), .A(n9505), .ZN(n9506) );
  AOI21_X1 U10824 ( .B1(n9507), .B2(n9658), .A(n9506), .ZN(n9508) );
  OAI211_X1 U10825 ( .C1(n5832), .C2(n9630), .A(n9509), .B(n9508), .ZN(
        P1_U3215) );
  NAND2_X1 U10826 ( .A1(n9511), .A2(n9510), .ZN(n9619) );
  NAND2_X1 U10827 ( .A1(n9512), .A2(n9586), .ZN(n9513) );
  AOI21_X1 U10828 ( .B1(n9617), .B2(n9619), .A(n9513), .ZN(n9587) );
  AND3_X1 U10829 ( .A1(n9617), .A2(n9619), .A3(n9513), .ZN(n9514) );
  OAI21_X1 U10830 ( .B1(n9587), .B2(n9514), .A(n9621), .ZN(n9518) );
  AOI22_X1 U10831 ( .A1(n9667), .A2(n9652), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3086), .ZN(n9515) );
  OAI21_X1 U10832 ( .B1(n9824), .B2(n9654), .A(n9515), .ZN(n9516) );
  AOI21_X1 U10833 ( .B1(n9828), .B2(n9658), .A(n9516), .ZN(n9517) );
  OAI211_X1 U10834 ( .C1(n10091), .C2(n9630), .A(n9518), .B(n9517), .ZN(
        P1_U3216) );
  XNOR2_X1 U10835 ( .A(n9519), .B(n9520), .ZN(n9633) );
  NOR2_X1 U10836 ( .A1(n9633), .A2(n9632), .ZN(n9631) );
  AOI21_X1 U10837 ( .B1(n9520), .B2(n9519), .A(n9631), .ZN(n9524) );
  XNOR2_X1 U10838 ( .A(n9522), .B(n9521), .ZN(n9523) );
  XNOR2_X1 U10839 ( .A(n9524), .B(n9523), .ZN(n9531) );
  NAND2_X1 U10840 ( .A1(n9640), .A2(n9883), .ZN(n9526) );
  OAI211_X1 U10841 ( .C1(n9527), .C2(n9643), .A(n9526), .B(n9525), .ZN(n9529)
         );
  NOR2_X1 U10842 ( .A1(n9890), .A2(n9630), .ZN(n9528) );
  AOI211_X1 U10843 ( .C1(n9887), .C2(n9658), .A(n9529), .B(n9528), .ZN(n9530)
         );
  OAI21_X1 U10844 ( .B1(n9531), .B2(n9662), .A(n9530), .ZN(P1_U3219) );
  XOR2_X1 U10845 ( .A(n9533), .B(n9532), .Z(n9538) );
  AOI22_X1 U10846 ( .A1(n9860), .A2(n9652), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n9535) );
  NAND2_X1 U10847 ( .A1(n9882), .A2(n9640), .ZN(n9534) );
  OAI211_X1 U10848 ( .C1(n9636), .C2(n9853), .A(n9535), .B(n9534), .ZN(n9536)
         );
  AOI21_X1 U10849 ( .B1(n10014), .B2(n9659), .A(n9536), .ZN(n9537) );
  OAI21_X1 U10850 ( .B1(n9538), .B2(n9662), .A(n9537), .ZN(P1_U3223) );
  INV_X1 U10851 ( .A(n9539), .ZN(n9541) );
  NOR3_X1 U10852 ( .A1(n4399), .A2(n9541), .A3(n9540), .ZN(n9544) );
  INV_X1 U10853 ( .A(n9542), .ZN(n9543) );
  OAI21_X1 U10854 ( .B1(n9544), .B2(n9543), .A(n9621), .ZN(n9550) );
  OAI21_X1 U10855 ( .B1(n9643), .B2(n9961), .A(n9545), .ZN(n9548) );
  NOR2_X1 U10856 ( .A1(n9636), .A2(n9546), .ZN(n9547) );
  AOI211_X1 U10857 ( .C1(n9640), .C2(n9673), .A(n9548), .B(n9547), .ZN(n9549)
         );
  OAI211_X1 U10858 ( .C1(n9551), .C2(n9630), .A(n9550), .B(n9549), .ZN(
        P1_U3224) );
  OAI21_X1 U10859 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9555) );
  NAND2_X1 U10860 ( .A1(n9555), .A2(n9621), .ZN(n9560) );
  NOR2_X1 U10861 ( .A1(n9788), .A2(n9636), .ZN(n9558) );
  OAI22_X1 U10862 ( .A1(n9823), .A2(n9654), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9556), .ZN(n9557) );
  AOI211_X1 U10863 ( .C1(n9666), .C2(n9652), .A(n9558), .B(n9557), .ZN(n9559)
         );
  OAI211_X1 U10864 ( .C1(n10083), .C2(n9630), .A(n9560), .B(n9559), .ZN(
        P1_U3225) );
  INV_X1 U10865 ( .A(n9561), .ZN(n9562) );
  NAND2_X1 U10866 ( .A1(n9563), .A2(n9562), .ZN(n9566) );
  INV_X1 U10867 ( .A(n9564), .ZN(n9565) );
  NAND2_X1 U10868 ( .A1(n9566), .A2(n9565), .ZN(n9567) );
  OAI21_X1 U10869 ( .B1(n9566), .B2(n9565), .A(n9567), .ZN(n9650) );
  NOR2_X1 U10870 ( .A1(n9650), .A2(n9651), .ZN(n9649) );
  INV_X1 U10871 ( .A(n9567), .ZN(n9568) );
  NOR2_X1 U10872 ( .A1(n9649), .A2(n9568), .ZN(n9573) );
  INV_X1 U10873 ( .A(n9569), .ZN(n9571) );
  NOR2_X1 U10874 ( .A1(n9571), .A2(n9570), .ZN(n9572) );
  XNOR2_X1 U10875 ( .A(n9573), .B(n9572), .ZN(n9578) );
  NAND2_X1 U10876 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10182)
         );
  OAI21_X1 U10877 ( .B1(n9643), .B2(n9899), .A(n10182), .ZN(n9574) );
  AOI21_X1 U10878 ( .B1(n9640), .B2(n9933), .A(n9574), .ZN(n9575) );
  OAI21_X1 U10879 ( .B1(n9636), .B2(n9940), .A(n9575), .ZN(n9576) );
  AOI21_X1 U10880 ( .B1(n9939), .B2(n9659), .A(n9576), .ZN(n9577) );
  OAI21_X1 U10881 ( .B1(n9578), .B2(n9662), .A(n9577), .ZN(P1_U3226) );
  XOR2_X1 U10882 ( .A(n9580), .B(n9579), .Z(n9585) );
  NAND2_X1 U10883 ( .A1(n9652), .A2(n9883), .ZN(n9581) );
  NAND2_X1 U10884 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10197)
         );
  OAI211_X1 U10885 ( .C1(n9918), .C2(n9654), .A(n9581), .B(n10197), .ZN(n9583)
         );
  NOR2_X1 U10886 ( .A1(n9926), .A2(n9630), .ZN(n9582) );
  AOI211_X1 U10887 ( .C1(n9923), .C2(n9658), .A(n9583), .B(n9582), .ZN(n9584)
         );
  OAI21_X1 U10888 ( .B1(n9585), .B2(n9662), .A(n9584), .ZN(P1_U3228) );
  INV_X1 U10889 ( .A(n9590), .ZN(n9812) );
  AOI22_X1 U10890 ( .A1(n9835), .A2(n9640), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n9591) );
  OAI21_X1 U10891 ( .B1(n9810), .B2(n9643), .A(n9591), .ZN(n9592) );
  AOI21_X1 U10892 ( .B1(n9812), .B2(n9658), .A(n9592), .ZN(n9593) );
  XNOR2_X1 U10893 ( .A(n9596), .B(n9595), .ZN(n9597) );
  XNOR2_X1 U10894 ( .A(n9598), .B(n9597), .ZN(n9603) );
  AOI22_X1 U10895 ( .A1(n9836), .A2(n9652), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3086), .ZN(n9600) );
  NAND2_X1 U10896 ( .A1(n9668), .A2(n9640), .ZN(n9599) );
  OAI211_X1 U10897 ( .C1(n9636), .C2(n9867), .A(n9600), .B(n9599), .ZN(n9601)
         );
  AOI21_X1 U10898 ( .B1(n10020), .B2(n9659), .A(n9601), .ZN(n9602) );
  OAI21_X1 U10899 ( .B1(n9603), .B2(n9662), .A(n9602), .ZN(P1_U3233) );
  OAI21_X1 U10900 ( .B1(n9606), .B2(n9605), .A(n9604), .ZN(n9607) );
  NAND2_X1 U10901 ( .A1(n9607), .A2(n9621), .ZN(n9614) );
  NAND2_X1 U10902 ( .A1(n9652), .A2(n9671), .ZN(n9609) );
  OAI211_X1 U10903 ( .C1(n9610), .C2(n9654), .A(n9609), .B(n9608), .ZN(n9611)
         );
  AOI21_X1 U10904 ( .B1(n9658), .B2(n9612), .A(n9611), .ZN(n9613) );
  OAI211_X1 U10905 ( .C1(n9615), .C2(n9630), .A(n9614), .B(n9613), .ZN(
        P1_U3234) );
  INV_X1 U10906 ( .A(n9619), .ZN(n9616) );
  NOR2_X1 U10907 ( .A1(n9617), .A2(n9616), .ZN(n9623) );
  AOI21_X1 U10908 ( .B1(n9620), .B2(n9619), .A(n9618), .ZN(n9622) );
  OAI21_X1 U10909 ( .B1(n9623), .B2(n9622), .A(n9621), .ZN(n9629) );
  NOR2_X1 U10910 ( .A1(n9636), .A2(n9840), .ZN(n9627) );
  OAI22_X1 U10911 ( .A1(n9625), .A2(n9643), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9624), .ZN(n9626) );
  AOI211_X1 U10912 ( .C1(n9640), .C2(n9836), .A(n9627), .B(n9626), .ZN(n9628)
         );
  OAI211_X1 U10913 ( .C1(n9839), .C2(n9630), .A(n9629), .B(n9628), .ZN(
        P1_U3235) );
  AOI21_X1 U10914 ( .B1(n9633), .B2(n9632), .A(n9631), .ZN(n9639) );
  NAND2_X1 U10915 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10217)
         );
  OAI21_X1 U10916 ( .B1(n9898), .B2(n9643), .A(n10217), .ZN(n9634) );
  AOI21_X1 U10917 ( .B1(n9640), .B2(n9935), .A(n9634), .ZN(n9635) );
  OAI21_X1 U10918 ( .B1(n9636), .B2(n9901), .A(n9635), .ZN(n9637) );
  AOI21_X1 U10919 ( .B1(n10031), .B2(n9659), .A(n9637), .ZN(n9638) );
  OAI21_X1 U10920 ( .B1(n9639), .B2(n9662), .A(n9638), .ZN(P1_U3238) );
  AOI22_X1 U10921 ( .A1(n5715), .A2(n9640), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3086), .ZN(n9642) );
  NAND2_X1 U10922 ( .A1(n9774), .A2(n9658), .ZN(n9641) );
  OAI211_X1 U10923 ( .C1(n9778), .C2(n9643), .A(n9642), .B(n9641), .ZN(n9647)
         );
  INV_X1 U10924 ( .A(n9648), .ZN(P1_U3240) );
  AOI21_X1 U10925 ( .B1(n9651), .B2(n9650), .A(n9649), .ZN(n9663) );
  NAND2_X1 U10926 ( .A1(n9652), .A2(n9669), .ZN(n9653) );
  NAND2_X1 U10927 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10169)
         );
  OAI211_X1 U10928 ( .C1(n9655), .C2(n9654), .A(n9653), .B(n10169), .ZN(n9656)
         );
  AOI21_X1 U10929 ( .B1(n9658), .B2(n9657), .A(n9656), .ZN(n9661) );
  NAND2_X1 U10930 ( .A1(n10051), .A2(n9659), .ZN(n9660) );
  OAI211_X1 U10931 ( .C1(n9663), .C2(n9662), .A(n9661), .B(n9660), .ZN(
        P1_U3241) );
  MUX2_X1 U10932 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9664), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10933 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9665), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10934 ( .A(n4698), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9670), .Z(
        P1_U3581) );
  MUX2_X1 U10935 ( .A(n9666), .B(P1_DATAO_REG_26__SCAN_IN), .S(n9670), .Z(
        P1_U3580) );
  MUX2_X1 U10936 ( .A(n5715), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9670), .Z(
        P1_U3579) );
  MUX2_X1 U10937 ( .A(n9667), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9670), .Z(
        P1_U3578) );
  MUX2_X1 U10938 ( .A(n9835), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9670), .Z(
        P1_U3577) );
  MUX2_X1 U10939 ( .A(n9860), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9670), .Z(
        P1_U3576) );
  MUX2_X1 U10940 ( .A(n9836), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9670), .Z(
        P1_U3575) );
  MUX2_X1 U10941 ( .A(n9882), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9670), .Z(
        P1_U3574) );
  MUX2_X1 U10942 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9668), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10943 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9883), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10944 ( .A(n9935), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9670), .Z(
        P1_U3571) );
  MUX2_X1 U10945 ( .A(n9669), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9670), .Z(
        P1_U3570) );
  MUX2_X1 U10946 ( .A(n9933), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9670), .Z(
        P1_U3569) );
  MUX2_X1 U10947 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9671), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10948 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9672), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10949 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n5449), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10950 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9673), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10951 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9674), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10952 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9675), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10953 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9676), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10954 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9677), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10955 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9678), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10956 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n4587), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10957 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9679), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10958 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9680), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10959 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9681), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10960 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n4643), .S(P1_U3973), .Z(
        P1_U3555) );
  OAI211_X1 U10961 ( .C1(n9684), .C2(n9683), .A(n9716), .B(n9682), .ZN(n9692)
         );
  AOI22_X1 U10962 ( .A1(n10141), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n9691) );
  NAND2_X1 U10963 ( .A1(n10168), .A2(n9685), .ZN(n9690) );
  OAI211_X1 U10964 ( .C1(n9688), .C2(n9687), .A(n10211), .B(n9686), .ZN(n9689)
         );
  NAND4_X1 U10965 ( .A1(n9692), .A2(n9691), .A3(n9690), .A4(n9689), .ZN(
        P1_U3244) );
  INV_X1 U10966 ( .A(n9693), .ZN(n9697) );
  INV_X1 U10967 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9695) );
  OAI21_X1 U10968 ( .B1(n10220), .B2(n9695), .A(n9694), .ZN(n9696) );
  AOI21_X1 U10969 ( .B1(n9697), .B2(n10168), .A(n9696), .ZN(n9706) );
  OAI211_X1 U10970 ( .C1(n9700), .C2(n9699), .A(n9716), .B(n9698), .ZN(n9705)
         );
  OAI211_X1 U10971 ( .C1(n9703), .C2(n9702), .A(n10211), .B(n9701), .ZN(n9704)
         );
  NAND3_X1 U10972 ( .A1(n9706), .A2(n9705), .A3(n9704), .ZN(P1_U3246) );
  AOI211_X1 U10973 ( .C1(n9709), .C2(n9708), .A(n9707), .B(n10158), .ZN(n9710)
         );
  INV_X1 U10974 ( .A(n9710), .ZN(n9721) );
  INV_X1 U10975 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9712) );
  OAI21_X1 U10976 ( .B1(n10220), .B2(n9712), .A(n9711), .ZN(n9713) );
  AOI21_X1 U10977 ( .B1(n9714), .B2(n10168), .A(n9713), .ZN(n9720) );
  OAI211_X1 U10978 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9715), .ZN(n9719)
         );
  NAND3_X1 U10979 ( .A1(n9721), .A2(n9720), .A3(n9719), .ZN(P1_U3248) );
  NOR2_X2 U10980 ( .A1(n9732), .A2(n9733), .ZN(n9731) );
  XNOR2_X1 U10981 ( .A(n10071), .B(n9731), .ZN(n9722) );
  NAND2_X1 U10982 ( .A1(n9723), .A2(n9973), .ZN(n9727) );
  INV_X1 U10983 ( .A(n9980), .ZN(n9726) );
  OR2_X1 U10984 ( .A1(n4287), .A2(n9726), .ZN(n9736) );
  OAI211_X1 U10985 ( .C1(n9971), .C2(n9728), .A(n9727), .B(n9736), .ZN(n9729)
         );
  AOI21_X1 U10986 ( .B1(n9977), .B2(n9944), .A(n9729), .ZN(n9730) );
  INV_X1 U10987 ( .A(n9730), .ZN(P1_U3263) );
  NAND2_X1 U10988 ( .A1(n9981), .A2(n9944), .ZN(n9737) );
  NAND2_X1 U10989 ( .A1(n9733), .A2(n9973), .ZN(n9735) );
  NAND2_X1 U10990 ( .A1(n4287), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n9734) );
  NAND4_X1 U10991 ( .A1(n9737), .A2(n9736), .A3(n9735), .A4(n9734), .ZN(
        P1_U3264) );
  NAND2_X1 U10992 ( .A1(n9739), .A2(n9738), .ZN(n9741) );
  XNOR2_X1 U10993 ( .A(n9741), .B(n9740), .ZN(n9751) );
  INV_X1 U10994 ( .A(n9742), .ZN(n9749) );
  NAND2_X1 U10995 ( .A1(n9743), .A2(n9944), .ZN(n9746) );
  AOI22_X1 U10996 ( .A1(n9744), .A2(n9922), .B1(P1_REG2_REG_29__SCAN_IN), .B2(
        n4287), .ZN(n9745) );
  OAI211_X1 U10997 ( .C1(n9747), .C2(n10227), .A(n9746), .B(n9745), .ZN(n9748)
         );
  AOI21_X1 U10998 ( .B1(n9749), .B2(n9971), .A(n9748), .ZN(n9750) );
  OAI21_X1 U10999 ( .B1(n9751), .B2(n9929), .A(n9750), .ZN(P1_U3356) );
  NAND2_X1 U11000 ( .A1(n9752), .A2(n9944), .ZN(n9755) );
  AOI22_X1 U11001 ( .A1(n9753), .A2(n9922), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n4287), .ZN(n9754) );
  OAI211_X1 U11002 ( .C1(n5812), .C2(n10227), .A(n9755), .B(n9754), .ZN(n9756)
         );
  AOI21_X1 U11003 ( .B1(n9757), .B2(n9971), .A(n9756), .ZN(n9758) );
  OAI21_X1 U11004 ( .B1(n4356), .B2(n9929), .A(n9758), .ZN(P1_U3265) );
  INV_X1 U11005 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n9760) );
  OAI22_X1 U11006 ( .A1(n9761), .A2(n10221), .B1(n9760), .B2(n9971), .ZN(n9771) );
  AOI211_X1 U11007 ( .C1(n9987), .C2(n4326), .A(n9952), .B(n7133), .ZN(n9986)
         );
  OR2_X1 U11008 ( .A1(n9766), .A2(n9962), .ZN(n9768) );
  NAND2_X1 U11009 ( .A1(n9666), .A2(n9932), .ZN(n9767) );
  OAI21_X1 U11010 ( .B1(n9989), .B2(n9929), .A(n9772), .ZN(P1_U3266) );
  AOI21_X1 U11011 ( .B1(n9786), .B2(n9780), .A(n9952), .ZN(n9773) );
  AND2_X1 U11012 ( .A1(n9773), .A2(n4326), .ZN(n9991) );
  AND2_X1 U11013 ( .A1(n9774), .A2(n9922), .ZN(n9779) );
  INV_X1 U11014 ( .A(n9775), .ZN(n9776) );
  AOI211_X1 U11015 ( .C1(n9991), .C2(n9871), .A(n9779), .B(n9990), .ZN(n9784)
         );
  AOI22_X1 U11016 ( .A1(n9780), .A2(n9973), .B1(n4287), .B2(
        P1_REG2_REG_26__SCAN_IN), .ZN(n9783) );
  NAND2_X1 U11017 ( .A1(n9992), .A2(n10231), .ZN(n9782) );
  OAI211_X1 U11018 ( .C1(n9784), .C2(n4287), .A(n9783), .B(n9782), .ZN(
        P1_U3267) );
  XNOR2_X1 U11019 ( .A(n9785), .B(n9792), .ZN(n9994) );
  OAI211_X1 U11020 ( .C1(n10083), .C2(n9811), .A(n10015), .B(n9786), .ZN(n9995) );
  INV_X1 U11021 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9787) );
  OAI22_X1 U11022 ( .A1(n9788), .A2(n10221), .B1(n9787), .B2(n9971), .ZN(n9789) );
  AOI21_X1 U11023 ( .B1(n9790), .B2(n9973), .A(n9789), .ZN(n9791) );
  OAI21_X1 U11024 ( .B1(n9995), .B2(n10224), .A(n9791), .ZN(n9799) );
  OR2_X1 U11025 ( .A1(n9794), .A2(n9793), .ZN(n9797) );
  OAI22_X1 U11026 ( .A1(n9795), .A2(n9962), .B1(n9823), .B2(n9960), .ZN(n9796)
         );
  AOI21_X1 U11027 ( .B1(n9797), .B2(n9966), .A(n9796), .ZN(n9996) );
  NOR2_X1 U11028 ( .A1(n9996), .A2(n4287), .ZN(n9798) );
  AOI211_X1 U11029 ( .C1(n10231), .C2(n9994), .A(n9799), .B(n9798), .ZN(n9800)
         );
  INV_X1 U11030 ( .A(n9800), .ZN(P1_U3268) );
  XNOR2_X1 U11031 ( .A(n9801), .B(n9802), .ZN(n10000) );
  INV_X1 U11032 ( .A(n10000), .ZN(n9817) );
  INV_X1 U11033 ( .A(n4278), .ZN(n9820) );
  OAI21_X1 U11034 ( .B1(n9820), .B2(n9805), .A(n9804), .ZN(n9807) );
  NAND3_X1 U11035 ( .A1(n9807), .A2(n9966), .A3(n9806), .ZN(n9809) );
  NAND2_X1 U11036 ( .A1(n9835), .A2(n9932), .ZN(n9808) );
  OAI211_X1 U11037 ( .C1(n9810), .C2(n9962), .A(n9809), .B(n9808), .ZN(n9998)
         );
  AOI211_X1 U11038 ( .C1(n5839), .C2(n9826), .A(n9952), .B(n9811), .ZN(n9999)
         );
  NAND2_X1 U11039 ( .A1(n9999), .A2(n9944), .ZN(n9814) );
  AOI22_X1 U11040 ( .A1(n9812), .A2(n9922), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4287), .ZN(n9813) );
  OAI211_X1 U11041 ( .C1(n10087), .C2(n10227), .A(n9814), .B(n9813), .ZN(n9815) );
  AOI21_X1 U11042 ( .B1(n9971), .B2(n9998), .A(n9815), .ZN(n9816) );
  OAI21_X1 U11043 ( .B1(n9929), .B2(n9817), .A(n9816), .ZN(P1_U3269) );
  XNOR2_X1 U11044 ( .A(n9818), .B(n9819), .ZN(n10005) );
  INV_X1 U11045 ( .A(n10005), .ZN(n9833) );
  INV_X1 U11046 ( .A(n9819), .ZN(n9821) );
  AOI21_X1 U11047 ( .B1(n4352), .B2(n9821), .A(n9820), .ZN(n9822) );
  OAI222_X1 U11048 ( .A1(n9960), .A2(n9824), .B1(n9962), .B2(n9823), .C1(n9916), .C2(n9822), .ZN(n10003) );
  AOI21_X1 U11049 ( .B1(n9838), .B2(n9825), .A(n9952), .ZN(n9827) );
  AND2_X1 U11050 ( .A1(n9827), .A2(n9826), .ZN(n10004) );
  NAND2_X1 U11051 ( .A1(n10004), .A2(n9944), .ZN(n9830) );
  AOI22_X1 U11052 ( .A1(n9828), .A2(n9922), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4287), .ZN(n9829) );
  OAI211_X1 U11053 ( .C1(n10091), .C2(n10227), .A(n9830), .B(n9829), .ZN(n9831) );
  AOI21_X1 U11054 ( .B1(n10003), .B2(n9971), .A(n9831), .ZN(n9832) );
  OAI21_X1 U11055 ( .B1(n9929), .B2(n9833), .A(n9832), .ZN(P1_U3270) );
  XNOR2_X1 U11056 ( .A(n9834), .B(n9846), .ZN(n9837) );
  AOI222_X1 U11057 ( .A1(n9966), .A2(n9837), .B1(n9836), .B2(n9932), .C1(n9835), .C2(n9934), .ZN(n10013) );
  OAI211_X1 U11058 ( .C1(n9839), .C2(n9852), .A(n10015), .B(n9838), .ZN(n10012) );
  INV_X1 U11059 ( .A(n9840), .ZN(n9841) );
  AOI22_X1 U11060 ( .A1(n9841), .A2(n9922), .B1(n4287), .B2(
        P1_REG2_REG_22__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U11061 ( .A1(n10009), .A2(n9973), .ZN(n9842) );
  OAI211_X1 U11062 ( .C1(n10012), .C2(n10224), .A(n9843), .B(n9842), .ZN(n9844) );
  INV_X1 U11063 ( .A(n9844), .ZN(n9849) );
  NAND2_X1 U11064 ( .A1(n9847), .A2(n9846), .ZN(n10008) );
  NAND3_X1 U11065 ( .A1(n9845), .A2(n10008), .A3(n10231), .ZN(n9848) );
  OAI211_X1 U11066 ( .C1(n10013), .C2(n4287), .A(n9849), .B(n9848), .ZN(
        P1_U3271) );
  INV_X1 U11067 ( .A(n9858), .ZN(n9851) );
  XNOR2_X1 U11068 ( .A(n9850), .B(n9851), .ZN(n10019) );
  AOI21_X1 U11069 ( .B1(n10014), .B2(n5159), .A(n9852), .ZN(n10016) );
  INV_X1 U11070 ( .A(n10014), .ZN(n9856) );
  INV_X1 U11071 ( .A(n9853), .ZN(n9854) );
  AOI22_X1 U11072 ( .A1(n4287), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n9854), .B2(
        n9922), .ZN(n9855) );
  OAI21_X1 U11073 ( .B1(n9856), .B2(n10227), .A(n9855), .ZN(n9863) );
  OAI21_X1 U11074 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9861) );
  AOI222_X1 U11075 ( .A1(n9966), .A2(n9861), .B1(n9860), .B2(n9934), .C1(n9882), .C2(n9932), .ZN(n10018) );
  NOR2_X1 U11076 ( .A1(n10018), .A2(n4287), .ZN(n9862) );
  AOI211_X1 U11077 ( .C1(n10016), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9865)
         );
  OAI21_X1 U11078 ( .B1(n10019), .B2(n9929), .A(n9865), .ZN(P1_U3272) );
  AOI21_X1 U11079 ( .B1(n9886), .B2(n10020), .A(n9952), .ZN(n9866) );
  AND2_X1 U11080 ( .A1(n9866), .A2(n5159), .ZN(n10022) );
  NOR2_X1 U11081 ( .A1(n9867), .A2(n10221), .ZN(n9870) );
  OAI222_X1 U11082 ( .A1(n9962), .A2(n9869), .B1(n9960), .B2(n9898), .C1(n9916), .C2(n9868), .ZN(n10021) );
  AOI211_X1 U11083 ( .C1(n10022), .C2(n9871), .A(n9870), .B(n10021), .ZN(n9876) );
  AOI22_X1 U11084 ( .A1(n10020), .A2(n9973), .B1(n4287), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9875) );
  XOR2_X1 U11085 ( .A(n9872), .B(n9873), .Z(n10023) );
  NAND2_X1 U11086 ( .A1(n10023), .A2(n10231), .ZN(n9874) );
  OAI211_X1 U11087 ( .C1(n9876), .C2(n4287), .A(n9875), .B(n9874), .ZN(
        P1_U3273) );
  XNOR2_X1 U11088 ( .A(n9878), .B(n9877), .ZN(n10030) );
  OAI21_X1 U11089 ( .B1(n9881), .B2(n9880), .A(n9879), .ZN(n9884) );
  AOI222_X1 U11090 ( .A1(n9966), .A2(n9884), .B1(n9883), .B2(n9932), .C1(n9882), .C2(n9934), .ZN(n10029) );
  INV_X1 U11091 ( .A(n10029), .ZN(n9892) );
  OR2_X1 U11092 ( .A1(n9890), .A2(n9907), .ZN(n9885) );
  AND3_X1 U11093 ( .A1(n9886), .A2(n9885), .A3(n10015), .ZN(n10026) );
  NAND2_X1 U11094 ( .A1(n10026), .A2(n9944), .ZN(n9889) );
  AOI22_X1 U11095 ( .A1(n4287), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9887), .B2(
        n9922), .ZN(n9888) );
  OAI211_X1 U11096 ( .C1(n9890), .C2(n10227), .A(n9889), .B(n9888), .ZN(n9891)
         );
  AOI21_X1 U11097 ( .B1(n9892), .B2(n9971), .A(n9891), .ZN(n9893) );
  OAI21_X1 U11098 ( .B1(n9929), .B2(n10030), .A(n9893), .ZN(P1_U3274) );
  INV_X1 U11099 ( .A(n9894), .ZN(n9895) );
  AOI21_X1 U11100 ( .B1(n9904), .B2(n9896), .A(n9895), .ZN(n9897) );
  OAI222_X1 U11101 ( .A1(n9960), .A2(n9899), .B1(n9962), .B2(n9898), .C1(n9916), .C2(n9897), .ZN(n10032) );
  NAND2_X1 U11102 ( .A1(n10032), .A2(n9971), .ZN(n9911) );
  NAND2_X1 U11103 ( .A1(n4287), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9900) );
  OAI21_X1 U11104 ( .B1(n10221), .B2(n9901), .A(n9900), .ZN(n9902) );
  AOI21_X1 U11105 ( .B1(n10031), .B2(n9973), .A(n9902), .ZN(n9910) );
  XOR2_X1 U11106 ( .A(n9903), .B(n9904), .Z(n10034) );
  NAND2_X1 U11107 ( .A1(n10034), .A2(n10231), .ZN(n9909) );
  NAND2_X1 U11108 ( .A1(n10031), .A2(n9919), .ZN(n9905) );
  NAND2_X1 U11109 ( .A1(n9905), .A2(n10015), .ZN(n9906) );
  NOR2_X1 U11110 ( .A1(n9907), .A2(n9906), .ZN(n10033) );
  NAND2_X1 U11111 ( .A1(n10033), .A2(n9944), .ZN(n9908) );
  NAND4_X1 U11112 ( .A1(n9911), .A2(n9910), .A3(n9909), .A4(n9908), .ZN(
        P1_U3275) );
  XNOR2_X1 U11113 ( .A(n4286), .B(n9913), .ZN(n10041) );
  XNOR2_X1 U11114 ( .A(n9914), .B(n9913), .ZN(n9915) );
  OAI222_X1 U11115 ( .A1(n9960), .A2(n9918), .B1(n9962), .B2(n9917), .C1(n9916), .C2(n9915), .ZN(n10037) );
  INV_X1 U11116 ( .A(n9938), .ZN(n9921) );
  INV_X1 U11117 ( .A(n9919), .ZN(n9920) );
  AOI211_X1 U11118 ( .C1(n10039), .C2(n9921), .A(n9952), .B(n9920), .ZN(n10038) );
  NAND2_X1 U11119 ( .A1(n10038), .A2(n9944), .ZN(n9925) );
  AOI22_X1 U11120 ( .A1(n4287), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9923), .B2(
        n9922), .ZN(n9924) );
  OAI211_X1 U11121 ( .C1(n9926), .C2(n10227), .A(n9925), .B(n9924), .ZN(n9927)
         );
  AOI21_X1 U11122 ( .B1(n9971), .B2(n10037), .A(n9927), .ZN(n9928) );
  OAI21_X1 U11123 ( .B1(n10041), .B2(n9929), .A(n9928), .ZN(P1_U3276) );
  OAI21_X1 U11124 ( .B1(n9946), .B2(n9931), .A(n9930), .ZN(n9936) );
  AOI222_X1 U11125 ( .A1(n9966), .A2(n9936), .B1(n9935), .B2(n9934), .C1(n9933), .C2(n9932), .ZN(n10042) );
  AOI211_X1 U11126 ( .C1(n9939), .C2(n4930), .A(n9952), .B(n9938), .ZN(n10044)
         );
  NOR2_X1 U11127 ( .A1(n10108), .A2(n10227), .ZN(n9943) );
  OAI22_X1 U11128 ( .A1(n9971), .A2(n9941), .B1(n9940), .B2(n10221), .ZN(n9942) );
  AOI211_X1 U11129 ( .C1(n10044), .C2(n9944), .A(n9943), .B(n9942), .ZN(n9948)
         );
  XNOR2_X1 U11130 ( .A(n9945), .B(n9946), .ZN(n10045) );
  NAND2_X1 U11131 ( .A1(n10045), .A2(n10231), .ZN(n9947) );
  OAI211_X1 U11132 ( .C1(n10042), .C2(n4287), .A(n9948), .B(n9947), .ZN(
        P1_U3277) );
  INV_X1 U11133 ( .A(n9949), .ZN(n9953) );
  INV_X1 U11134 ( .A(n9950), .ZN(n9951) );
  AOI211_X1 U11135 ( .C1(n10055), .C2(n9953), .A(n9952), .B(n9951), .ZN(n10054) );
  INV_X1 U11136 ( .A(n10054), .ZN(n9976) );
  XNOR2_X1 U11137 ( .A(n9955), .B(n9958), .ZN(n10058) );
  NAND2_X1 U11138 ( .A1(n9957), .A2(n9956), .ZN(n9959) );
  XNOR2_X1 U11139 ( .A(n9959), .B(n9958), .ZN(n9967) );
  OAI22_X1 U11140 ( .A1(n9963), .A2(n9962), .B1(n9961), .B2(n9960), .ZN(n9965)
         );
  NOR2_X1 U11141 ( .A1(n10058), .A2(n10278), .ZN(n9964) );
  AOI211_X1 U11142 ( .C1(n9967), .C2(n9966), .A(n9965), .B(n9964), .ZN(n10057)
         );
  OAI21_X1 U11143 ( .B1(n10058), .B2(n9968), .A(n10057), .ZN(n9969) );
  NAND2_X1 U11144 ( .A1(n9969), .A2(n9971), .ZN(n9975) );
  OAI22_X1 U11145 ( .A1(n9971), .A2(n4830), .B1(n9970), .B2(n10221), .ZN(n9972) );
  AOI21_X1 U11146 ( .B1(n10055), .B2(n9973), .A(n9972), .ZN(n9974) );
  OAI211_X1 U11147 ( .C1(n9976), .C2(n10224), .A(n9975), .B(n9974), .ZN(
        P1_U3279) );
  NOR2_X1 U11148 ( .A1(n9977), .A2(n9980), .ZN(n10068) );
  MUX2_X1 U11149 ( .A(n9978), .B(n10068), .S(n10291), .Z(n9979) );
  OAI21_X1 U11150 ( .B1(n10071), .B2(n10048), .A(n9979), .ZN(P1_U3553) );
  NOR2_X1 U11151 ( .A1(n9981), .A2(n9980), .ZN(n10072) );
  MUX2_X1 U11152 ( .A(n9982), .B(n10072), .S(n10291), .Z(n9983) );
  OAI21_X1 U11153 ( .B1(n10075), .B2(n10048), .A(n9983), .ZN(P1_U3552) );
  OAI21_X1 U11154 ( .B1(n10265), .B2(n9989), .A(n9988), .ZN(n10076) );
  MUX2_X1 U11155 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10076), .S(n10291), .Z(
        P1_U3549) );
  AOI211_X1 U11156 ( .C1(n10000), .C2(n10250), .A(n9999), .B(n9998), .ZN(
        n10084) );
  MUX2_X1 U11157 ( .A(n10001), .B(n10084), .S(n10291), .Z(n10002) );
  OAI21_X1 U11158 ( .B1(n10087), .B2(n10048), .A(n10002), .ZN(P1_U3546) );
  AOI211_X1 U11159 ( .C1(n10005), .C2(n10250), .A(n10004), .B(n10003), .ZN(
        n10088) );
  MUX2_X1 U11160 ( .A(n10006), .B(n10088), .S(n10291), .Z(n10007) );
  OAI21_X1 U11161 ( .B1(n10091), .B2(n10048), .A(n10007), .ZN(P1_U3545) );
  NAND3_X1 U11162 ( .A1(n9845), .A2(n10008), .A3(n10250), .ZN(n10011) );
  NAND2_X1 U11163 ( .A1(n10009), .A2(n10261), .ZN(n10010) );
  NAND4_X1 U11164 ( .A1(n10013), .A2(n10012), .A3(n10011), .A4(n10010), .ZN(
        n10092) );
  MUX2_X1 U11165 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10092), .S(n10291), .Z(
        P1_U3544) );
  AOI22_X1 U11166 ( .A1(n10016), .A2(n10015), .B1(n10261), .B2(n10014), .ZN(
        n10017) );
  OAI211_X1 U11167 ( .C1(n10265), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        n10093) );
  MUX2_X1 U11168 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10093), .S(n10291), .Z(
        P1_U3543) );
  INV_X1 U11169 ( .A(n10020), .ZN(n10097) );
  AOI211_X1 U11170 ( .C1(n10023), .C2(n10250), .A(n10022), .B(n10021), .ZN(
        n10094) );
  MUX2_X1 U11171 ( .A(n10024), .B(n10094), .S(n10291), .Z(n10025) );
  OAI21_X1 U11172 ( .B1(n10097), .B2(n10048), .A(n10025), .ZN(P1_U3542) );
  AOI21_X1 U11173 ( .B1(n10261), .B2(n10027), .A(n10026), .ZN(n10028) );
  OAI211_X1 U11174 ( .C1(n10265), .C2(n10030), .A(n10029), .B(n10028), .ZN(
        n10098) );
  MUX2_X1 U11175 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10098), .S(n10291), .Z(
        P1_U3541) );
  INV_X1 U11176 ( .A(n10031), .ZN(n10102) );
  AOI211_X1 U11177 ( .C1(n10034), .C2(n10250), .A(n10033), .B(n10032), .ZN(
        n10099) );
  MUX2_X1 U11178 ( .A(n10035), .B(n10099), .S(n10291), .Z(n10036) );
  OAI21_X1 U11179 ( .B1(n10102), .B2(n10048), .A(n10036), .ZN(P1_U3540) );
  AOI211_X1 U11180 ( .C1(n10261), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10040) );
  OAI21_X1 U11181 ( .B1(n10265), .B2(n10041), .A(n10040), .ZN(n10103) );
  MUX2_X1 U11182 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10103), .S(n10291), .Z(
        P1_U3539) );
  INV_X1 U11183 ( .A(n10042), .ZN(n10043) );
  AOI211_X1 U11184 ( .C1(n10045), .C2(n10250), .A(n10044), .B(n10043), .ZN(
        n10104) );
  MUX2_X1 U11185 ( .A(n10046), .B(n10104), .S(n10291), .Z(n10047) );
  OAI21_X1 U11186 ( .B1(n10108), .B2(n10048), .A(n10047), .ZN(P1_U3538) );
  AOI211_X1 U11187 ( .C1(n10261), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        n10052) );
  OAI21_X1 U11188 ( .B1(n10265), .B2(n10053), .A(n10052), .ZN(n10109) );
  MUX2_X1 U11189 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n10109), .S(n10291), .Z(
        P1_U3537) );
  AOI21_X1 U11190 ( .B1(n10261), .B2(n10055), .A(n10054), .ZN(n10056) );
  OAI211_X1 U11191 ( .C1(n10058), .C2(n10277), .A(n10057), .B(n10056), .ZN(
        n10110) );
  MUX2_X1 U11192 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n10110), .S(n10291), .Z(
        P1_U3536) );
  AOI211_X1 U11193 ( .C1(n10261), .C2(n5450), .A(n10060), .B(n10059), .ZN(
        n10061) );
  OAI21_X1 U11194 ( .B1(n10265), .B2(n10062), .A(n10061), .ZN(n10111) );
  MUX2_X1 U11195 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10111), .S(n10291), .Z(
        P1_U3534) );
  AOI211_X1 U11196 ( .C1(n10261), .C2(n10065), .A(n10064), .B(n10063), .ZN(
        n10066) );
  OAI21_X1 U11197 ( .B1(n10265), .B2(n10067), .A(n10066), .ZN(n10112) );
  MUX2_X1 U11198 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10112), .S(n10291), .Z(
        P1_U3533) );
  MUX2_X1 U11199 ( .A(n10069), .B(n10068), .S(n10283), .Z(n10070) );
  OAI21_X1 U11200 ( .B1(n10071), .B2(n10107), .A(n10070), .ZN(P1_U3521) );
  INV_X1 U11201 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10073) );
  MUX2_X1 U11202 ( .A(n10073), .B(n10072), .S(n10283), .Z(n10074) );
  OAI21_X1 U11203 ( .B1(n10075), .B2(n10107), .A(n10074), .ZN(P1_U3520) );
  MUX2_X1 U11204 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10076), .S(n10283), .Z(
        P1_U3517) );
  INV_X1 U11205 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n10078) );
  INV_X1 U11206 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n10081) );
  MUX2_X1 U11207 ( .A(n10081), .B(n10080), .S(n10283), .Z(n10082) );
  INV_X1 U11208 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n10085) );
  MUX2_X1 U11209 ( .A(n10085), .B(n10084), .S(n10283), .Z(n10086) );
  OAI21_X1 U11210 ( .B1(n10087), .B2(n10107), .A(n10086), .ZN(P1_U3514) );
  INV_X1 U11211 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n10089) );
  MUX2_X1 U11212 ( .A(n10089), .B(n10088), .S(n10283), .Z(n10090) );
  OAI21_X1 U11213 ( .B1(n10091), .B2(n10107), .A(n10090), .ZN(P1_U3513) );
  MUX2_X1 U11214 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10092), .S(n10283), .Z(
        P1_U3512) );
  MUX2_X1 U11215 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10093), .S(n10283), .Z(
        P1_U3511) );
  INV_X1 U11216 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10095) );
  MUX2_X1 U11217 ( .A(n10095), .B(n10094), .S(n10283), .Z(n10096) );
  OAI21_X1 U11218 ( .B1(n10097), .B2(n10107), .A(n10096), .ZN(P1_U3510) );
  MUX2_X1 U11219 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10098), .S(n10283), .Z(
        P1_U3509) );
  INV_X1 U11220 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10100) );
  MUX2_X1 U11221 ( .A(n10100), .B(n10099), .S(n10283), .Z(n10101) );
  OAI21_X1 U11222 ( .B1(n10102), .B2(n10107), .A(n10101), .ZN(P1_U3507) );
  MUX2_X1 U11223 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10103), .S(n10283), .Z(
        P1_U3504) );
  INV_X1 U11224 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n10105) );
  MUX2_X1 U11225 ( .A(n10105), .B(n10104), .S(n10283), .Z(n10106) );
  OAI21_X1 U11226 ( .B1(n10108), .B2(n10107), .A(n10106), .ZN(P1_U3501) );
  MUX2_X1 U11227 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n10109), .S(n10283), .Z(
        P1_U3498) );
  MUX2_X1 U11228 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10110), .S(n10283), .Z(
        P1_U3495) );
  MUX2_X1 U11229 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10111), .S(n10283), .Z(
        P1_U3489) );
  MUX2_X1 U11230 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10112), .S(n10283), .Z(
        P1_U3486) );
  MUX2_X1 U11231 ( .A(P1_D_REG_1__SCAN_IN), .B(n10115), .S(n10235), .Z(
        P1_U3440) );
  MUX2_X1 U11232 ( .A(P1_D_REG_0__SCAN_IN), .B(n10116), .S(n10235), .Z(
        P1_U3439) );
  INV_X1 U11233 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10118) );
  NAND3_X1 U11234 ( .A1(n10118), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10120) );
  OAI22_X1 U11235 ( .A1(n10117), .A2(n10120), .B1(n10119), .B2(n10128), .ZN(
        n10121) );
  AOI21_X1 U11236 ( .B1(n10123), .B2(n10122), .A(n10121), .ZN(n10124) );
  INV_X1 U11237 ( .A(n10124), .ZN(P1_U3324) );
  INV_X1 U11238 ( .A(n7021), .ZN(n10126) );
  OAI222_X1 U11239 ( .A1(n10128), .A2(n10127), .B1(n10134), .B2(n10126), .C1(
        n4675), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U11240 ( .A1(n10131), .A2(P1_U3086), .B1(n10134), .B2(n10130), 
        .C1(n10129), .C2(n10128), .ZN(P1_U3329) );
  OAI222_X1 U11241 ( .A1(n10135), .A2(P1_U3086), .B1(n10134), .B2(n10133), 
        .C1(n10132), .C2(n10128), .ZN(P1_U3330) );
  INV_X1 U11242 ( .A(n10136), .ZN(n10137) );
  MUX2_X1 U11243 ( .A(n10137), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U11244 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11245 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U11246 ( .B1(n5846), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10138), .ZN(
        n10140) );
  XNOR2_X1 U11247 ( .A(n10140), .B(n10139), .ZN(n10144) );
  AOI22_X1 U11248 ( .A1(n10141), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10142) );
  OAI21_X1 U11249 ( .B1(n10144), .B2(n10143), .A(n10142), .ZN(P1_U3243) );
  INV_X1 U11250 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10157) );
  AOI211_X1 U11251 ( .C1(n10147), .C2(n10146), .A(n10206), .B(n10145), .ZN(
        n10152) );
  AOI211_X1 U11252 ( .C1(n10150), .C2(n10149), .A(n10158), .B(n10148), .ZN(
        n10151) );
  AOI211_X1 U11253 ( .C1(n10168), .C2(n10153), .A(n10152), .B(n10151), .ZN(
        n10156) );
  INV_X1 U11254 ( .A(n10154), .ZN(n10155) );
  OAI211_X1 U11255 ( .C1(n10220), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        P1_U3257) );
  AOI211_X1 U11256 ( .C1(n10161), .C2(n10160), .A(n10159), .B(n10158), .ZN(
        n10166) );
  AOI211_X1 U11257 ( .C1(n10164), .C2(n10163), .A(n10162), .B(n10206), .ZN(
        n10165) );
  AOI211_X1 U11258 ( .C1(n10168), .C2(n10167), .A(n10166), .B(n10165), .ZN(
        n10170) );
  OAI211_X1 U11259 ( .C1(n10171), .C2(n10220), .A(n10170), .B(n10169), .ZN(
        P1_U3258) );
  OAI21_X1 U11260 ( .B1(n10174), .B2(n10173), .A(n10172), .ZN(n10181) );
  NOR2_X1 U11261 ( .A1(n10215), .A2(n10175), .ZN(n10180) );
  AOI211_X1 U11262 ( .C1(n10178), .C2(n10177), .A(n10176), .B(n10206), .ZN(
        n10179) );
  AOI211_X1 U11263 ( .C1(n10211), .C2(n10181), .A(n10180), .B(n10179), .ZN(
        n10183) );
  OAI211_X1 U11264 ( .C1(n10220), .C2(n10184), .A(n10183), .B(n10182), .ZN(
        P1_U3259) );
  INV_X1 U11265 ( .A(n10185), .ZN(n10195) );
  INV_X1 U11266 ( .A(n10186), .ZN(n10187) );
  XNOR2_X1 U11267 ( .A(n10188), .B(n10187), .ZN(n10189) );
  OR2_X1 U11268 ( .A1(n10206), .A2(n10189), .ZN(n10194) );
  XNOR2_X1 U11269 ( .A(n10191), .B(n10190), .ZN(n10192) );
  NAND2_X1 U11270 ( .A1(n10211), .A2(n10192), .ZN(n10193) );
  OAI211_X1 U11271 ( .C1(n10215), .C2(n10195), .A(n10194), .B(n10193), .ZN(
        n10196) );
  INV_X1 U11272 ( .A(n10196), .ZN(n10198) );
  OAI211_X1 U11273 ( .C1(n10220), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        P1_U3260) );
  INV_X1 U11274 ( .A(n10200), .ZN(n10214) );
  NAND2_X1 U11275 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND2_X1 U11276 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  OR2_X1 U11277 ( .A1(n10206), .A2(n10205), .ZN(n10213) );
  NAND2_X1 U11278 ( .A1(n10208), .A2(n10207), .ZN(n10209) );
  NAND3_X1 U11279 ( .A1(n10211), .A2(n10210), .A3(n10209), .ZN(n10212) );
  OAI211_X1 U11280 ( .C1(n10215), .C2(n10214), .A(n10213), .B(n10212), .ZN(
        n10216) );
  INV_X1 U11281 ( .A(n10216), .ZN(n10218) );
  OAI211_X1 U11282 ( .C1(n10220), .C2(n10219), .A(n10218), .B(n10217), .ZN(
        P1_U3261) );
  OAI22_X1 U11283 ( .A1(n10224), .A2(n10223), .B1(n10222), .B2(n10221), .ZN(
        n10225) );
  AOI21_X1 U11284 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n4287), .A(n10225), .ZN(
        n10226) );
  OAI21_X1 U11285 ( .B1(n10228), .B2(n10227), .A(n10226), .ZN(n10229) );
  AOI21_X1 U11286 ( .B1(n10231), .B2(n10230), .A(n10229), .ZN(n10232) );
  OAI21_X1 U11287 ( .B1(n4287), .B2(n10233), .A(n10232), .ZN(P1_U3291) );
  AND2_X1 U11288 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10236), .ZN(P1_U3294) );
  AND2_X1 U11289 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10236), .ZN(P1_U3295) );
  AND2_X1 U11290 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10236), .ZN(P1_U3296) );
  AND2_X1 U11291 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10236), .ZN(P1_U3297) );
  AND2_X1 U11292 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10236), .ZN(P1_U3298) );
  AND2_X1 U11293 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10236), .ZN(P1_U3299) );
  AND2_X1 U11294 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10236), .ZN(P1_U3300) );
  AND2_X1 U11295 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10236), .ZN(P1_U3301) );
  AND2_X1 U11296 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10236), .ZN(P1_U3302) );
  AND2_X1 U11297 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10236), .ZN(P1_U3303) );
  AND2_X1 U11298 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10236), .ZN(P1_U3304) );
  AND2_X1 U11299 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10236), .ZN(P1_U3305) );
  AND2_X1 U11300 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10236), .ZN(P1_U3306) );
  AND2_X1 U11301 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10236), .ZN(P1_U3307) );
  AND2_X1 U11302 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10236), .ZN(P1_U3308) );
  AND2_X1 U11303 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10236), .ZN(P1_U3309) );
  AND2_X1 U11304 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10236), .ZN(P1_U3310) );
  AND2_X1 U11305 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10236), .ZN(P1_U3311) );
  AND2_X1 U11306 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10236), .ZN(P1_U3312) );
  AND2_X1 U11307 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10236), .ZN(P1_U3313) );
  AND2_X1 U11308 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10236), .ZN(P1_U3314) );
  NOR2_X1 U11309 ( .A1(n10235), .A2(n10234), .ZN(P1_U3315) );
  AND2_X1 U11310 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10236), .ZN(P1_U3316) );
  AND2_X1 U11311 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10236), .ZN(P1_U3317) );
  AND2_X1 U11312 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10236), .ZN(P1_U3318) );
  AND2_X1 U11313 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10236), .ZN(P1_U3319) );
  AND2_X1 U11314 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10236), .ZN(P1_U3320) );
  AND2_X1 U11315 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10236), .ZN(P1_U3321) );
  AND2_X1 U11316 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10236), .ZN(P1_U3322) );
  AND2_X1 U11317 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10236), .ZN(P1_U3323) );
  AOI22_X1 U11318 ( .A1(n10283), .A2(n10237), .B1(n5249), .B2(n10282), .ZN(
        P1_U3453) );
  INV_X1 U11319 ( .A(n10261), .ZN(n10274) );
  OAI21_X1 U11320 ( .B1(n10239), .B2(n10274), .A(n10238), .ZN(n10242) );
  INV_X1 U11321 ( .A(n10240), .ZN(n10241) );
  AOI211_X1 U11322 ( .C1(n10250), .C2(n10243), .A(n10242), .B(n10241), .ZN(
        n10284) );
  AOI22_X1 U11323 ( .A1(n10283), .A2(n10284), .B1(n5180), .B2(n10282), .ZN(
        P1_U3462) );
  OAI21_X1 U11324 ( .B1(n10245), .B2(n10274), .A(n10244), .ZN(n10248) );
  INV_X1 U11325 ( .A(n10246), .ZN(n10247) );
  AOI211_X1 U11326 ( .C1(n10250), .C2(n10249), .A(n10248), .B(n10247), .ZN(
        n10285) );
  INV_X1 U11327 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U11328 ( .A1(n10283), .A2(n10285), .B1(n10251), .B2(n10282), .ZN(
        P1_U3465) );
  AOI21_X1 U11329 ( .B1(n10261), .B2(n10253), .A(n10252), .ZN(n10254) );
  OAI211_X1 U11330 ( .C1(n10265), .C2(n10256), .A(n10255), .B(n10254), .ZN(
        n10257) );
  INV_X1 U11331 ( .A(n10257), .ZN(n10286) );
  INV_X1 U11332 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10258) );
  AOI22_X1 U11333 ( .A1(n10283), .A2(n10286), .B1(n10258), .B2(n10282), .ZN(
        P1_U3468) );
  AOI21_X1 U11334 ( .B1(n10261), .B2(n10260), .A(n10259), .ZN(n10262) );
  OAI211_X1 U11335 ( .C1(n10265), .C2(n10264), .A(n10263), .B(n10262), .ZN(
        n10266) );
  INV_X1 U11336 ( .A(n10266), .ZN(n10287) );
  INV_X1 U11337 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U11338 ( .A1(n10283), .A2(n10287), .B1(n10267), .B2(n10282), .ZN(
        P1_U3471) );
  INV_X1 U11339 ( .A(n10277), .ZN(n10272) );
  OAI21_X1 U11340 ( .B1(n4933), .B2(n10274), .A(n10268), .ZN(n10270) );
  AOI211_X1 U11341 ( .C1(n10272), .C2(n10271), .A(n10270), .B(n10269), .ZN(
        n10288) );
  AOI22_X1 U11342 ( .A1(n10283), .A2(n10288), .B1(n5335), .B2(n10282), .ZN(
        P1_U3474) );
  OAI21_X1 U11343 ( .B1(n10275), .B2(n10274), .A(n10273), .ZN(n10280) );
  AOI21_X1 U11344 ( .B1(n10278), .B2(n10277), .A(n10276), .ZN(n10279) );
  NOR3_X1 U11345 ( .A1(n10281), .A2(n10280), .A3(n10279), .ZN(n10290) );
  AOI22_X1 U11346 ( .A1(n10283), .A2(n10290), .B1(n5359), .B2(n10282), .ZN(
        P1_U3477) );
  AOI22_X1 U11347 ( .A1(n10291), .A2(n10284), .B1(n6448), .B2(n10289), .ZN(
        P1_U3525) );
  AOI22_X1 U11348 ( .A1(n10291), .A2(n10285), .B1(n6450), .B2(n10289), .ZN(
        P1_U3526) );
  AOI22_X1 U11349 ( .A1(n10291), .A2(n10286), .B1(n6451), .B2(n10289), .ZN(
        P1_U3527) );
  AOI22_X1 U11350 ( .A1(n10291), .A2(n10287), .B1(n6452), .B2(n10289), .ZN(
        P1_U3528) );
  AOI22_X1 U11351 ( .A1(n10291), .A2(n10288), .B1(n6453), .B2(n10289), .ZN(
        P1_U3529) );
  AOI22_X1 U11352 ( .A1(n10291), .A2(n10290), .B1(n5354), .B2(n10289), .ZN(
        P1_U3530) );
  AOI22_X1 U11353 ( .A1(n10301), .A2(n6738), .B1(n10292), .B2(n10298), .ZN(
        P2_U3393) );
  AOI22_X1 U11354 ( .A1(n10301), .A2(n6749), .B1(n10293), .B2(n10298), .ZN(
        P2_U3396) );
  AOI22_X1 U11355 ( .A1(n10301), .A2(n6761), .B1(n10294), .B2(n10298), .ZN(
        P2_U3399) );
  AOI22_X1 U11356 ( .A1(n10301), .A2(n6774), .B1(n10295), .B2(n10298), .ZN(
        P2_U3402) );
  INV_X1 U11357 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10297) );
  AOI22_X1 U11358 ( .A1(n10301), .A2(n10297), .B1(n10296), .B2(n10298), .ZN(
        P2_U3405) );
  INV_X1 U11359 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10300) );
  AOI22_X1 U11360 ( .A1(n10301), .A2(n10300), .B1(n10299), .B2(n10298), .ZN(
        P2_U3408) );
  OAI222_X1 U11361 ( .A1(n10306), .A2(n10305), .B1(n10306), .B2(n10304), .C1(
        n10303), .C2(n10302), .ZN(ADD_1068_U5) );
  AOI21_X1 U11362 ( .B1(n10309), .B2(n10308), .A(n10307), .ZN(ADD_1068_U46) );
  INV_X1 U11363 ( .A(n10312), .ZN(n10311) );
  OAI222_X1 U11364 ( .A1(n10314), .A2(n10313), .B1(n10314), .B2(n10312), .C1(
        n10311), .C2(n10310), .ZN(ADD_1068_U55) );
  OAI21_X1 U11365 ( .B1(n10317), .B2(n10316), .A(n10315), .ZN(ADD_1068_U56) );
  OAI21_X1 U11366 ( .B1(n10320), .B2(n10319), .A(n10318), .ZN(ADD_1068_U57) );
  OAI21_X1 U11367 ( .B1(n10323), .B2(n10322), .A(n10321), .ZN(ADD_1068_U58) );
  OAI21_X1 U11368 ( .B1(n10326), .B2(n10325), .A(n10324), .ZN(ADD_1068_U59) );
  OAI21_X1 U11369 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(ADD_1068_U60) );
  OAI21_X1 U11370 ( .B1(n10332), .B2(n10331), .A(n10330), .ZN(ADD_1068_U61) );
  OAI21_X1 U11371 ( .B1(n10335), .B2(n10334), .A(n10333), .ZN(ADD_1068_U62) );
  OAI21_X1 U11372 ( .B1(n10338), .B2(n10337), .A(n10336), .ZN(ADD_1068_U63) );
  OAI21_X1 U11373 ( .B1(n10341), .B2(n10340), .A(n10339), .ZN(ADD_1068_U50) );
  OAI21_X1 U11374 ( .B1(n10344), .B2(n10343), .A(n10342), .ZN(ADD_1068_U51) );
  OAI21_X1 U11375 ( .B1(n10347), .B2(n10346), .A(n10345), .ZN(ADD_1068_U47) );
  OAI21_X1 U11376 ( .B1(n10350), .B2(n10349), .A(n10348), .ZN(ADD_1068_U49) );
  OAI21_X1 U11377 ( .B1(n10353), .B2(n10352), .A(n10351), .ZN(ADD_1068_U48) );
  AOI21_X1 U11378 ( .B1(n10356), .B2(n10355), .A(n10354), .ZN(ADD_1068_U54) );
  AOI21_X1 U11379 ( .B1(n10359), .B2(n10358), .A(n10357), .ZN(ADD_1068_U53) );
  OAI21_X1 U11380 ( .B1(n10362), .B2(n10361), .A(n10360), .ZN(ADD_1068_U52) );
  NOR2_X1 U6984 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5172) );
  NOR2_X1 U6985 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5171) );
  NAND2_X1 U4882 ( .A1(n5190), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4807) );
  INV_X1 U7040 ( .A(n5330), .ZN(n5653) );
  BUF_X2 U4909 ( .A(n5035), .Z(n6735) );
  NAND2_X1 U4886 ( .A1(n7389), .A2(n7390), .ZN(n7687) );
  NOR2_X2 U4839 ( .A1(n7995), .A2(n10065), .ZN(n7994) );
  BUF_X2 U4802 ( .A(n6381), .Z(n6424) );
  CLKBUF_X1 U4811 ( .A(n9803), .Z(n4278) );
  AND2_X1 U4827 ( .A1(n4858), .A2(n4334), .ZN(n9091) );
  CLKBUF_X1 U4832 ( .A(n4581), .Z(n4573) );
  CLKBUF_X1 U4842 ( .A(n9206), .Z(n4280) );
  INV_X2 U4844 ( .A(n6419), .ZN(n4289) );
  NAND2_X2 U4900 ( .A1(n8384), .A2(n10125), .ZN(n5270) );
  OAI21_X1 U4901 ( .B1(n7156), .B2(P1_DATAO_REG_2__SCAN_IN), .A(n5199), .ZN(
        n5207) );
  INV_X2 U5017 ( .A(n5653), .ZN(n5889) );
  CLKBUF_X1 U5065 ( .A(n7078), .Z(n4302) );
  CLKBUF_X1 U6087 ( .A(n10125), .Z(n4675) );
  CLKBUF_X1 U6356 ( .A(n6165), .Z(n4590) );
  AND2_X1 U6504 ( .A1(n5140), .A2(n8733), .ZN(n10367) );
endmodule

