

module b22_C_SARLock_k_64_4 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6433, n6434, n6435, n6436, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037;

  NAND2_X1 U7182 ( .A1(n7080), .A2(n12833), .ZN(n13075) );
  NAND2_X1 U7183 ( .A1(n11451), .A2(n11450), .ZN(n13131) );
  NAND2_X1 U7184 ( .A1(n10386), .A2(n10385), .ZN(n10404) );
  OAI21_X1 U7185 ( .B1(n8224), .B2(n8223), .A(n6924), .ZN(n6923) );
  NOR2_X1 U7186 ( .A1(n14457), .A2(n14456), .ZN(n14455) );
  NAND2_X2 U7187 ( .A1(n9908), .A2(n9839), .ZN(n11823) );
  INV_X2 U7188 ( .A(n12183), .ZN(n12076) );
  BUF_X2 U7189 ( .A(n8601), .Z(n12043) );
  NOR2_X2 U7190 ( .A1(n13838), .A2(n9542), .ZN(n10390) );
  BUF_X2 U7191 ( .A(n8043), .Z(n8471) );
  INV_X1 U7192 ( .A(n10758), .ZN(n11434) );
  CLKBUF_X2 U7193 ( .A(n9511), .Z(n11607) );
  INV_X2 U7194 ( .A(n11869), .ZN(n9542) );
  AND2_X1 U7195 ( .A1(n9313), .A2(n13201), .ZN(n9354) );
  NAND2_X1 U7196 ( .A1(n6788), .A2(n7921), .ZN(n8034) );
  CLKBUF_X1 U7197 ( .A(n14052), .Z(n6433) );
  NOR2_X1 U7198 ( .A1(n10873), .A2(n14837), .ZN(n14052) );
  NAND2_X1 U7199 ( .A1(n9542), .A2(n10494), .ZN(n9838) );
  AOI21_X1 U7200 ( .B1(n8718), .B2(n6591), .A(n7595), .ZN(n11220) );
  NOR2_X1 U7201 ( .A1(n7651), .A2(n7612), .ZN(n7613) );
  NAND2_X1 U7202 ( .A1(n7016), .A2(n7015), .ZN(n11708) );
  INV_X1 U7203 ( .A(n9510), .ZN(n11724) );
  OR2_X1 U7204 ( .A1(n14516), .A2(n14515), .ZN(n7352) );
  INV_X1 U7205 ( .A(n11026), .ZN(n11433) );
  AOI21_X2 U7206 ( .B1(n11010), .B2(n12771), .A(n11009), .ZN(n11023) );
  NOR2_X1 U7207 ( .A1(n10985), .A2(n11661), .ZN(n11009) );
  INV_X1 U7208 ( .A(n11856), .ZN(n11813) );
  AND2_X1 U7209 ( .A1(n13537), .A2(n8488), .ZN(n13555) );
  CLKBUF_X2 U7210 ( .A(n8593), .Z(n12033) );
  OR2_X1 U7211 ( .A1(n8896), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8911) );
  OAI21_X1 U7212 ( .B1(n7003), .B2(n7002), .A(n6999), .ZN(n10187) );
  AND2_X1 U7214 ( .A1(n7428), .A2(n7427), .ZN(n12891) );
  AND2_X2 U7215 ( .A1(n13823), .A2(n13826), .ZN(n8012) );
  AOI21_X1 U7216 ( .B1(n11448), .B2(n8460), .A(n7594), .ZN(n13799) );
  OR2_X1 U7217 ( .A1(n8524), .A2(P1_IR_REG_26__SCAN_IN), .ZN(n8526) );
  NAND2_X1 U7218 ( .A1(n8533), .A2(n7729), .ZN(n12654) );
  CLKBUF_X2 U7219 ( .A(n7737), .Z(n12659) );
  AND2_X1 U7220 ( .A1(n10391), .A2(n10394), .ZN(n6434) );
  AND3_X1 U7221 ( .A1(n6539), .A2(n7588), .A3(n7613), .ZN(n6435) );
  INV_X1 U7222 ( .A(n11290), .ZN(n6448) );
  NOR3_X2 U7223 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .A3(
        P1_IR_REG_6__SCAN_IN), .ZN(n7920) );
  OAI21_X1 U7224 ( .B1(n13528), .B2(n7031), .A(n13676), .ZN(n13666) );
  NAND2_X2 U7225 ( .A1(n12675), .A2(n11712), .ZN(n12717) );
  XNOR2_X2 U7226 ( .A(n13778), .B(n13532), .ZN(n13638) );
  AOI21_X2 U7227 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n9623), .A(n9492), .ZN(
        n14457) );
  NAND2_X2 U7228 ( .A1(n9514), .A2(n9513), .ZN(n14579) );
  XNOR2_X2 U7229 ( .A(n6712), .B(n13538), .ZN(n13743) );
  XNOR2_X2 U7230 ( .A(n7731), .B(n7730), .ZN(n7737) );
  NOR2_X2 U7231 ( .A1(n8659), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8670) );
  XNOR2_X2 U7232 ( .A(n9695), .B(P2_IR_REG_16__SCAN_IN), .ZN(n14522) );
  OAI22_X2 U7233 ( .A1(n13602), .A2(n13603), .B1(n13534), .B2(n13533), .ZN(
        n13591) );
  NAND2_X2 U7234 ( .A1(n13622), .A2(n6967), .ZN(n13602) );
  AOI21_X2 U7235 ( .B1(n9401), .B2(P2_REG1_REG_2__SCAN_IN), .A(n9397), .ZN(
        n14448) );
  NAND2_X2 U7236 ( .A1(n9332), .A2(n12819), .ZN(n9575) );
  OAI21_X2 U7237 ( .B1(n10404), .B2(n10403), .A(n10405), .ZN(n10443) );
  AOI22_X2 U7238 ( .A1(n13032), .A2(n12838), .B1(n12837), .B2(n13141), .ZN(
        n13018) );
  NAND4_X2 U7239 ( .A1(n9336), .A2(n9335), .A3(n9334), .A4(n9333), .ZN(n11293)
         );
  AOI21_X2 U7240 ( .B1(n14463), .B2(P2_REG2_REG_5__SCAN_IN), .A(n14455), .ZN(
        n9494) );
  NAND2_X4 U7241 ( .A1(n8385), .A2(n8384), .ZN(n13778) );
  INV_X1 U7242 ( .A(n10577), .ZN(n6815) );
  XNOR2_X1 U7243 ( .A(n10577), .B(n13353), .ZN(n9707) );
  NAND2_X2 U7244 ( .A1(n6820), .A2(n7996), .ZN(n10577) );
  XNOR2_X2 U7245 ( .A(n7950), .B(P1_IR_REG_22__SCAN_IN), .ZN(n13838) );
  AOI21_X2 U7246 ( .B1(n12430), .B2(n12432), .A(n12058), .ZN(n12423) );
  NAND2_X2 U7247 ( .A1(n12440), .A2(n12151), .ZN(n12430) );
  INV_X1 U7248 ( .A(n11823), .ZN(n6436) );
  INV_X1 U7250 ( .A(n6450), .ZN(n6438) );
  INV_X1 U7251 ( .A(n6451), .ZN(n6439) );
  INV_X1 U7252 ( .A(n6451), .ZN(n6440) );
  INV_X1 U7253 ( .A(n6450), .ZN(n6441) );
  INV_X1 U7254 ( .A(n6440), .ZN(n6442) );
  INV_X1 U7255 ( .A(n6442), .ZN(n6443) );
  INV_X1 U7256 ( .A(n6442), .ZN(n6444) );
  INV_X1 U7257 ( .A(n6442), .ZN(n6445) );
  INV_X1 U7258 ( .A(n6442), .ZN(n6446) );
  INV_X1 U7259 ( .A(n6442), .ZN(n6447) );
  INV_X2 U7260 ( .A(n6448), .ZN(n6449) );
  INV_X1 U7261 ( .A(n6448), .ZN(n6450) );
  INV_X1 U7262 ( .A(n6448), .ZN(n6451) );
  INV_X1 U7263 ( .A(n11290), .ZN(n11301) );
  AOI21_X2 U7264 ( .B1(n10419), .B2(n12774), .A(n10418), .ZN(n10423) );
  AOI21_X2 U7265 ( .B1(n12888), .B2(n12889), .A(n6907), .ZN(n12885) );
  OAI22_X2 U7266 ( .A1(n12913), .A2(n12912), .B1(n12911), .B2(n12883), .ZN(
        n12888) );
  XNOR2_X2 U7267 ( .A(n7900), .B(SI_24_), .ZN(n8395) );
  OAI21_X2 U7268 ( .B1(n8383), .B2(n10645), .A(n7899), .ZN(n7900) );
  XNOR2_X2 U7269 ( .A(n7942), .B(n7940), .ZN(n13826) );
  OAI21_X2 U7270 ( .B1(n8395), .B2(n6868), .A(n7901), .ZN(n8413) );
  NAND2_X4 U7271 ( .A1(n11029), .A2(n11028), .ZN(n13156) );
  AOI21_X2 U7272 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9860), .A(n9685), .ZN(
        n9687) );
  NOR2_X2 U7273 ( .A1(n7868), .A2(n7262), .ZN(n7261) );
  XNOR2_X2 U7274 ( .A(n12805), .B(n12790), .ZN(n12792) );
  AOI21_X2 U7275 ( .B1(n14536), .B2(P2_REG2_REG_17__SCAN_IN), .A(n14526), .ZN(
        n12805) );
  XNOR2_X2 U7276 ( .A(n7369), .B(n9103), .ZN(n9129) );
  AND2_X2 U7277 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n7369) );
  AND2_X1 U7278 ( .A1(n13562), .A2(n13561), .ZN(n13744) );
  INV_X2 U7279 ( .A(n11605), .ZN(n13083) );
  OAI21_X1 U7280 ( .B1(n13309), .B2(n6736), .A(n6734), .ZN(n13293) );
  AND2_X1 U7281 ( .A1(n7972), .A2(n7971), .ZN(n13739) );
  OAI22_X1 U7282 ( .A1(n11406), .A2(n6780), .B1(n11407), .B2(n6466), .ZN(
        n11415) );
  NAND2_X1 U7283 ( .A1(n13223), .A2(n11750), .ZN(n11754) );
  NAND2_X1 U7284 ( .A1(n11046), .A2(n11045), .ZN(n12859) );
  NAND2_X1 U7285 ( .A1(n10944), .A2(n10943), .ZN(n11394) );
  OR2_X1 U7286 ( .A1(n10253), .A2(n6743), .ZN(n10255) );
  NOR2_X1 U7287 ( .A1(n9893), .A2(n6545), .ZN(n9905) );
  NAND2_X1 U7288 ( .A1(n12094), .A2(n12093), .ZN(n12088) );
  NAND2_X1 U7289 ( .A1(n12080), .A2(n12085), .ZN(n14759) );
  INV_X1 U7290 ( .A(n11325), .ZN(n14588) );
  INV_X1 U7291 ( .A(n10782), .ZN(n12278) );
  CLKBUF_X2 U7292 ( .A(n8106), .Z(n8271) );
  INV_X1 U7293 ( .A(n13352), .ZN(n10572) );
  INV_X1 U7294 ( .A(n9363), .ZN(n10046) );
  NAND4_X1 U7295 ( .A1(n8596), .A2(n8594), .A3(n8595), .A4(n8597), .ZN(n12279)
         );
  AND4_X2 U7296 ( .A1(n7989), .A2(n7987), .A3(n7986), .A4(n7988), .ZN(n7108)
         );
  INV_X4 U7297 ( .A(n14352), .ZN(n9843) );
  INV_X1 U7298 ( .A(n11293), .ZN(n10043) );
  INV_X4 U7299 ( .A(n11823), .ZN(n6452) );
  INV_X1 U7300 ( .A(n8005), .ZN(n6455) );
  INV_X4 U7301 ( .A(n11607), .ZN(n11584) );
  INV_X2 U7302 ( .A(n9247), .ZN(n8310) );
  NAND2_X1 U7303 ( .A1(n12646), .A2(n8537), .ZN(n8592) );
  BUF_X2 U7304 ( .A(n9353), .Z(n11590) );
  NAND2_X1 U7305 ( .A1(n8527), .A2(n8526), .ZN(n13835) );
  NAND2_X1 U7306 ( .A1(n8526), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7928) );
  OR2_X1 U7307 ( .A1(n7631), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n7642) );
  NOR2_X1 U7308 ( .A1(n8034), .A2(n7416), .ZN(n7121) );
  NOR2_X1 U7309 ( .A1(n8034), .A2(n7414), .ZN(n7413) );
  INV_X4 U7311 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7646) );
  AOI21_X1 U7312 ( .B1(n13576), .B2(n13575), .A(n13574), .ZN(n13753) );
  NAND2_X1 U7313 ( .A1(n7390), .A2(n13555), .ZN(n13554) );
  NAND2_X1 U7314 ( .A1(n13262), .A2(n11839), .ZN(n13318) );
  OR2_X1 U7315 ( .A1(n11510), .A2(n7520), .ZN(n7519) );
  XNOR2_X1 U7316 ( .A(n11884), .B(n11873), .ZN(n11991) );
  NAND2_X1 U7317 ( .A1(n13627), .A2(n7318), .ZN(n13767) );
  OR2_X1 U7318 ( .A1(n13649), .A2(n13648), .ZN(n13780) );
  NAND2_X1 U7319 ( .A1(n11972), .A2(n11971), .ZN(n11970) );
  NAND2_X1 U7320 ( .A1(n13624), .A2(n13623), .ZN(n13622) );
  AND2_X1 U7321 ( .A1(n8473), .A2(n8472), .ZN(n13736) );
  NOR2_X1 U7322 ( .A1(n12816), .A2(n14527), .ZN(n7368) );
  XNOR2_X1 U7323 ( .A(n13096), .B(n12769), .ZN(n12912) );
  AND2_X2 U7324 ( .A1(n12205), .A2(n12200), .ZN(n12300) );
  INV_X1 U7325 ( .A(n12310), .ZN(n12312) );
  INV_X1 U7326 ( .A(n13739), .ZN(n6453) );
  NAND2_X1 U7327 ( .A1(n11576), .A2(n11575), .ZN(n13088) );
  NAND2_X2 U7328 ( .A1(n11554), .A2(n11553), .ZN(n7078) );
  OR2_X1 U7329 ( .A1(n12552), .A2(n12316), .ZN(n12205) );
  CLKBUF_X1 U7330 ( .A(n12682), .Z(n6952) );
  XNOR2_X1 U7331 ( .A(n13631), .B(n6879), .ZN(n13623) );
  AOI21_X1 U7332 ( .B1(n7394), .B2(n7392), .A(n7402), .ZN(n7391) );
  NAND2_X1 U7333 ( .A1(n6711), .A2(n13508), .ZN(n13702) );
  NAND2_X1 U7334 ( .A1(n11249), .A2(n11248), .ZN(n12016) );
  NAND2_X1 U7335 ( .A1(n6823), .A2(n13786), .ZN(n13655) );
  OAI22_X1 U7336 ( .A1(n8905), .A2(n8906), .B1(P2_DATAO_REG_27__SCAN_IN), .B2(
        n13205), .ZN(n8919) );
  OAI21_X1 U7337 ( .B1(n11754), .B2(n6728), .A(n11764), .ZN(n6725) );
  NAND2_X1 U7338 ( .A1(n11502), .A2(n11501), .ZN(n13116) );
  NAND2_X1 U7339 ( .A1(n6667), .A2(n6921), .ZN(n8905) );
  AND2_X1 U7340 ( .A1(n7354), .A2(n7353), .ZN(n14529) );
  NAND2_X1 U7341 ( .A1(n8891), .A2(n8890), .ZN(n6667) );
  NOR2_X1 U7342 ( .A1(n6482), .A2(n13529), .ZN(n6824) );
  OAI21_X1 U7343 ( .B1(n11237), .B2(n6635), .A(n6633), .ZN(n11244) );
  NAND2_X1 U7344 ( .A1(n7312), .A2(n7311), .ZN(n14139) );
  AOI21_X1 U7345 ( .B1(n12482), .B2(n12136), .A(n12138), .ZN(n12475) );
  NOR2_X1 U7346 ( .A1(n7451), .A2(n12836), .ZN(n7447) );
  AND2_X1 U7347 ( .A1(n6642), .A2(n12135), .ZN(n12482) );
  AND2_X1 U7348 ( .A1(n12858), .A2(n6582), .ZN(n7454) );
  NAND2_X1 U7349 ( .A1(n7896), .A2(n7895), .ZN(n7898) );
  OR2_X1 U7350 ( .A1(n11385), .A2(n11384), .ZN(n7608) );
  NAND2_X1 U7351 ( .A1(n6643), .A2(n12126), .ZN(n11223) );
  NOR2_X1 U7352 ( .A1(n12787), .A2(n14490), .ZN(n12788) );
  OR2_X1 U7353 ( .A1(n6483), .A2(n10625), .ZN(n7099) );
  NAND2_X1 U7354 ( .A1(n11054), .A2(n12229), .ZN(n6643) );
  NAND2_X1 U7355 ( .A1(n11172), .A2(n11171), .ZN(n13151) );
  NAND2_X1 U7356 ( .A1(n6666), .A2(n8824), .ZN(n8833) );
  OAI21_X1 U7357 ( .B1(n6769), .B2(n6770), .A(n7537), .ZN(n11361) );
  AND2_X1 U7358 ( .A1(n7885), .A2(n6895), .ZN(n7273) );
  NOR2_X1 U7359 ( .A1(n11349), .A2(n6772), .ZN(n6769) );
  OAI21_X1 U7360 ( .B1(n8221), .B2(n7265), .A(n6850), .ZN(n7884) );
  NAND2_X1 U7361 ( .A1(n6691), .A2(n7328), .ZN(n8813) );
  NAND2_X1 U7362 ( .A1(n6434), .A2(n6822), .ZN(n10541) );
  NAND2_X1 U7363 ( .A1(n10179), .A2(n10178), .ZN(n11356) );
  OR2_X1 U7364 ( .A1(n11341), .A2(n11342), .ZN(n11343) );
  AND2_X1 U7365 ( .A1(n6656), .A2(n6655), .ZN(n10705) );
  NAND2_X1 U7366 ( .A1(n10087), .A2(n10086), .ZN(n14617) );
  NAND2_X1 U7367 ( .A1(n8081), .A2(n8080), .ZN(n10858) );
  OAI21_X1 U7368 ( .B1(n6776), .B2(n6775), .A(n6774), .ZN(n11334) );
  NAND2_X1 U7369 ( .A1(n6998), .A2(n6997), .ZN(n7476) );
  NAND2_X1 U7370 ( .A1(n10462), .A2(n12221), .ZN(n10461) );
  AND2_X1 U7371 ( .A1(n10121), .A2(n10147), .ZN(n11649) );
  XNOR2_X1 U7372 ( .A(n8568), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8733) );
  NOR2_X1 U7373 ( .A1(n9991), .A2(n7364), .ZN(n14468) );
  AND2_X1 U7374 ( .A1(n10127), .A2(n10051), .ZN(n11648) );
  NOR2_X1 U7375 ( .A1(n9687), .A2(n9686), .ZN(n9991) );
  NAND2_X1 U7376 ( .A1(n10580), .A2(n10367), .ZN(n10649) );
  INV_X4 U7377 ( .A(n11268), .ZN(n9067) );
  OR2_X2 U7378 ( .A1(n11824), .A2(n14091), .ZN(n11815) );
  AND4_X1 U7379 ( .A1(n8610), .A2(n8609), .A3(n8608), .A4(n8607), .ZN(n14761)
         );
  AND2_X1 U7380 ( .A1(n9843), .A2(n10114), .ZN(n14091) );
  CLKBUF_X3 U7381 ( .A(n8611), .Z(n12042) );
  NAND4_X1 U7382 ( .A1(n9359), .A2(n9358), .A3(n9357), .A4(n9356), .ZN(n12781)
         );
  INV_X1 U7383 ( .A(n8592), .ZN(n6458) );
  AND2_X1 U7384 ( .A1(n6641), .A2(n6640), .ZN(n14458) );
  INV_X1 U7385 ( .A(n8592), .ZN(n6457) );
  OR2_X1 U7386 ( .A1(n9488), .A2(n6500), .ZN(n6641) );
  NAND2_X4 U7387 ( .A1(n8934), .A2(n9154), .ZN(n8601) );
  NAND2_X2 U7388 ( .A1(n9544), .A2(n9838), .ZN(n11856) );
  INV_X2 U7389 ( .A(n13965), .ZN(n6454) );
  BUF_X2 U7390 ( .A(n9517), .Z(n11591) );
  NAND2_X1 U7391 ( .A1(n7724), .A2(n6880), .ZN(n6883) );
  INV_X1 U7392 ( .A(n12646), .ZN(n8538) );
  AND2_X1 U7393 ( .A1(n8536), .A2(n12639), .ZN(n8537) );
  NAND2_X1 U7394 ( .A1(n7069), .A2(n6890), .ZN(n12646) );
  BUF_X2 U7395 ( .A(n9355), .Z(n11612) );
  AND2_X1 U7396 ( .A1(n11671), .A2(n11680), .ZN(n14546) );
  CLKBUF_X1 U7397 ( .A(n10758), .Z(n11608) );
  OR2_X1 U7398 ( .A1(n14445), .A2(n14444), .ZN(n7358) );
  OR2_X1 U7399 ( .A1(n9330), .A2(n9331), .ZN(n14543) );
  NAND2_X1 U7400 ( .A1(n11026), .A2(n9154), .ZN(n9511) );
  NAND2_X1 U7401 ( .A1(n8516), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7950) );
  INV_X1 U7402 ( .A(n10389), .ZN(n10494) );
  AND2_X1 U7403 ( .A1(n11235), .A2(n13201), .ZN(n9355) );
  NAND2_X1 U7404 ( .A1(n6856), .A2(n6855), .ZN(n7982) );
  MUX2_X1 U7405 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7727), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7729) );
  NAND2_X1 U7406 ( .A1(n6639), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7731) );
  XNOR2_X1 U7407 ( .A(n7936), .B(n7935), .ZN(n13828) );
  NOR2_X1 U7408 ( .A1(n9400), .A2(n7359), .ZN(n14445) );
  XNOR2_X1 U7409 ( .A(n7941), .B(n6713), .ZN(n13823) );
  NAND2_X1 U7410 ( .A1(n7317), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U7411 ( .A1(n13817), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7941) );
  AND2_X1 U7412 ( .A1(n6435), .A2(n7649), .ZN(n7622) );
  XNOR2_X1 U7413 ( .A(n7619), .B(n7620), .ZN(n11282) );
  XNOR2_X2 U7414 ( .A(n9293), .B(P2_IR_REG_19__SCAN_IN), .ZN(n11680) );
  NAND3_X1 U7415 ( .A1(n9308), .A2(n9119), .A3(n9118), .ZN(n9126) );
  NOR2_X1 U7416 ( .A1(n7186), .A2(n6882), .ZN(n6881) );
  NOR2_X1 U7417 ( .A1(n9292), .A2(n7509), .ZN(n9289) );
  NAND2_X1 U7418 ( .A1(n9120), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9122) );
  AND2_X1 U7419 ( .A1(n7122), .A2(n7121), .ZN(n7951) );
  OR2_X1 U7420 ( .A1(n9110), .A2(n13197), .ZN(n9112) );
  NAND2_X1 U7421 ( .A1(n7071), .A2(n6476), .ZN(n9118) );
  INV_X1 U7422 ( .A(n6759), .ZN(n9292) );
  AND2_X1 U7423 ( .A1(n8670), .A2(n10033), .ZN(n8682) );
  NAND2_X2 U7424 ( .A1(n6866), .A2(n6864), .ZN(n7847) );
  INV_X1 U7425 ( .A(n7922), .ZN(n7122) );
  NOR2_X1 U7426 ( .A1(n7617), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n7588) );
  NOR2_X2 U7427 ( .A1(n7672), .A2(n7671), .ZN(n9216) );
  AND2_X1 U7428 ( .A1(n7649), .A2(n6581), .ZN(n7058) );
  INV_X1 U7429 ( .A(n9129), .ZN(n9301) );
  OR2_X1 U7430 ( .A1(n8649), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8659) );
  NAND2_X1 U7431 ( .A1(n6867), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6866) );
  AND2_X2 U7432 ( .A1(n9104), .A2(n9021), .ZN(n9162) );
  NAND3_X1 U7433 ( .A1(n13992), .A2(n7274), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n6867) );
  AND2_X1 U7434 ( .A1(n7616), .A2(n6884), .ZN(n7593) );
  AND3_X1 U7435 ( .A1(n7635), .A2(n7615), .A3(n7632), .ZN(n7592) );
  INV_X1 U7436 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9155) );
  INV_X1 U7437 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7700) );
  INV_X1 U7438 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n13992) );
  NOR2_X1 U7439 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7545) );
  INV_X1 U7440 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7650) );
  INV_X4 U7441 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7442 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9021) );
  INV_X1 U7443 ( .A(n13197), .ZN(n6456) );
  NOR2_X1 U7444 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n7370) );
  NOR2_X1 U7445 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n7371) );
  NOR2_X1 U7446 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n9019) );
  INV_X1 U7447 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7632) );
  INV_X1 U7448 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7635) );
  INV_X4 U7449 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  INV_X1 U7450 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9936) );
  INV_X1 U7451 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7660) );
  INV_X1 U7452 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7656) );
  INV_X1 U7453 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n7662) );
  NOR2_X1 U7454 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n9018) );
  OAI211_X1 U7455 ( .C1(n11026), .C2(n9352), .A(n9350), .B(n9351), .ZN(n9363)
         );
  XNOR2_X1 U7456 ( .A(n7970), .B(n7969), .ZN(n13200) );
  INV_X4 U7457 ( .A(n8027), .ZN(n8011) );
  NAND2_X1 U7458 ( .A1(n13823), .A2(n7959), .ZN(n8027) );
  AOI21_X2 U7459 ( .B1(n7259), .B2(n7260), .A(n7258), .ZN(n7257) );
  NAND2_X1 U7460 ( .A1(n9575), .A2(n11638), .ZN(n9510) );
  NOR2_X1 U7461 ( .A1(n11014), .A2(n14491), .ZN(n14490) );
  AND2_X1 U7462 ( .A1(n7997), .A2(n6821), .ZN(n6820) );
  OR2_X4 U7463 ( .A1(n14543), .A2(n11646), .ZN(n9339) );
  AOI21_X1 U7464 ( .B1(n9129), .B2(P2_REG1_REG_1__SCAN_IN), .A(n9139), .ZN(
        n9128) );
  NOR2_X2 U7465 ( .A1(n13051), .A2(n13141), .ZN(n7073) );
  NOR2_X2 U7466 ( .A1(n8754), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8767) );
  OR2_X2 U7467 ( .A1(n8752), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U7468 ( .A1(n9575), .A2(n11638), .ZN(n6459) );
  NOR2_X2 U7469 ( .A1(n10741), .A2(n13172), .ZN(n7081) );
  AOI21_X2 U7470 ( .B1(n14637), .B2(n7078), .A(n13092), .ZN(n13093) );
  NOR2_X2 U7471 ( .A1(n8911), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n14050) );
  NOR2_X1 U7472 ( .A1(n7193), .A2(n12870), .ZN(n7192) );
  INV_X1 U7473 ( .A(n7196), .ZN(n7193) );
  MUX2_X1 U7474 ( .A(n13528), .B(n13799), .S(n8106), .Z(n8340) );
  INV_X1 U7475 ( .A(n11446), .ZN(n6955) );
  OAI21_X1 U7476 ( .B1(n13745), .B2(n8017), .A(n6938), .ZN(n8463) );
  NAND2_X1 U7477 ( .A1(n13521), .A2(n8017), .ZN(n6938) );
  NAND2_X1 U7478 ( .A1(n6859), .A2(n6857), .ZN(n8462) );
  AND2_X1 U7479 ( .A1(n6863), .A2(n6858), .ZN(n6857) );
  NAND2_X1 U7480 ( .A1(n6861), .A2(n6862), .ZN(n6858) );
  OAI22_X1 U7481 ( .A1(n7447), .A2(n7443), .B1(n7455), .B2(n12862), .ZN(n7440)
         );
  NAND2_X1 U7482 ( .A1(n11754), .A2(n6727), .ZN(n6726) );
  AND2_X1 U7483 ( .A1(n11755), .A2(n13330), .ZN(n6727) );
  AND2_X1 U7484 ( .A1(n12254), .A2(n9042), .ZN(n9043) );
  AND2_X1 U7485 ( .A1(n6499), .A2(n7188), .ZN(n7185) );
  NOR2_X1 U7486 ( .A1(n10953), .A2(n7500), .ZN(n7012) );
  OR2_X1 U7487 ( .A1(n7078), .A2(n12849), .ZN(n12844) );
  AND2_X1 U7488 ( .A1(n7197), .A2(n12868), .ZN(n7196) );
  NAND2_X1 U7489 ( .A1(n12866), .A2(n7198), .ZN(n7197) );
  INV_X1 U7490 ( .A(n12865), .ZN(n7198) );
  OAI21_X1 U7491 ( .B1(n13018), .B2(n13017), .A(n6502), .ZN(n13004) );
  AOI21_X1 U7492 ( .B1(n12859), .B2(n7203), .A(n7202), .ZN(n13043) );
  NOR2_X1 U7493 ( .A1(n7205), .A2(n12862), .ZN(n7203) );
  NAND2_X1 U7494 ( .A1(n13293), .A2(n13292), .ZN(n7243) );
  NAND2_X1 U7495 ( .A1(n7222), .A2(n7220), .ZN(n13262) );
  AOI21_X1 U7496 ( .B1(n7223), .B2(n7225), .A(n7221), .ZN(n7220) );
  INV_X1 U7497 ( .A(n13264), .ZN(n7221) );
  INV_X1 U7498 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8199) );
  OR2_X1 U7499 ( .A1(n10820), .A2(n7133), .ZN(n7132) );
  NOR2_X1 U7500 ( .A1(n8209), .A2(n8207), .ZN(n7133) );
  AND3_X1 U7501 ( .A1(n8491), .A2(n8321), .A3(n13707), .ZN(n7111) );
  NAND2_X1 U7502 ( .A1(n11391), .A2(n6598), .ZN(n7536) );
  NAND2_X1 U7503 ( .A1(n6802), .A2(n8361), .ZN(n6801) );
  INV_X1 U7504 ( .A(n11413), .ZN(n6892) );
  NAND2_X1 U7505 ( .A1(n7524), .A2(n11509), .ZN(n7520) );
  AND2_X1 U7506 ( .A1(n7120), .A2(n8450), .ZN(n6988) );
  NAND2_X1 U7507 ( .A1(n14630), .A2(n9330), .ZN(n11290) );
  NOR2_X1 U7508 ( .A1(n13146), .A2(n7456), .ZN(n7455) );
  INV_X1 U7509 ( .A(n12863), .ZN(n7456) );
  NAND2_X1 U7510 ( .A1(n13096), .A2(n12883), .ZN(n7436) );
  AND2_X1 U7511 ( .A1(n7459), .A2(n7460), .ZN(n7449) );
  NAND2_X1 U7512 ( .A1(n7887), .A2(n9759), .ZN(n7890) );
  INV_X1 U7513 ( .A(n6851), .ZN(n6850) );
  OAI21_X1 U7514 ( .B1(n7265), .B2(n6982), .A(n7263), .ZN(n6851) );
  AOI21_X1 U7515 ( .B1(n7264), .B2(n7269), .A(n6608), .ZN(n7263) );
  INV_X1 U7516 ( .A(n7866), .ZN(n7262) );
  AND2_X1 U7517 ( .A1(n8988), .A2(n8926), .ZN(n12206) );
  OR2_X1 U7518 ( .A1(n12500), .A2(n12314), .ZN(n12193) );
  AND2_X1 U7519 ( .A1(n7572), .A2(n6567), .ZN(n7570) );
  AND2_X1 U7520 ( .A1(n12578), .A2(n12384), .ZN(n12168) );
  AND2_X1 U7521 ( .A1(n7577), .A2(n6568), .ZN(n7575) );
  OR2_X1 U7522 ( .A1(n12578), .A2(n12384), .ZN(n12176) );
  OAI21_X1 U7523 ( .B1(n11220), .B2(n7552), .A(n7550), .ZN(n12467) );
  INV_X1 U7524 ( .A(n7551), .ZN(n7550) );
  OAI21_X1 U7525 ( .B1(n6593), .B2(n7552), .A(n12464), .ZN(n7551) );
  INV_X1 U7526 ( .A(n7553), .ZN(n7552) );
  NAND2_X1 U7527 ( .A1(n7592), .A2(n7593), .ZN(n7617) );
  NAND2_X1 U7528 ( .A1(n8566), .A2(n8565), .ZN(n8568) );
  NAND2_X1 U7529 ( .A1(n8728), .A2(n8726), .ZN(n8566) );
  INV_X1 U7530 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7611) );
  AOI21_X1 U7531 ( .B1(n6686), .B2(n8557), .A(n6595), .ZN(n6684) );
  AND2_X1 U7532 ( .A1(n14536), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6652) );
  INV_X1 U7533 ( .A(n7459), .ZN(n7452) );
  INV_X1 U7534 ( .A(n7449), .ZN(n7446) );
  AOI21_X1 U7535 ( .B1(n10750), .B2(n10979), .A(n6506), .ZN(n7212) );
  NAND2_X1 U7536 ( .A1(n7190), .A2(n10219), .ZN(n10226) );
  AND2_X1 U7537 ( .A1(n9110), .A2(n9111), .ZN(n9034) );
  NAND2_X1 U7538 ( .A1(n10847), .A2(n10848), .ZN(n7237) );
  NAND2_X1 U7539 ( .A1(n8477), .A2(n9542), .ZN(n6790) );
  NAND2_X1 U7540 ( .A1(n13569), .A2(n13536), .ZN(n7390) );
  OR2_X1 U7541 ( .A1(n14116), .A2(n14086), .ZN(n13503) );
  XNOR2_X1 U7542 ( .A(n13349), .B(n10559), .ZN(n10384) );
  AND2_X1 U7543 ( .A1(n9247), .A2(n9299), .ZN(n8005) );
  OR2_X1 U7544 ( .A1(n13700), .A2(n13717), .ZN(n7032) );
  NOR2_X1 U7545 ( .A1(n10370), .A2(n14367), .ZN(n7296) );
  AOI21_X1 U7546 ( .B1(n6560), .B2(n10370), .A(n7295), .ZN(n7294) );
  NOR2_X1 U7547 ( .A1(n10368), .A2(n10652), .ZN(n7295) );
  OAI21_X1 U7548 ( .B1(n8427), .B2(n7282), .A(n7280), .ZN(n8459) );
  AOI21_X1 U7549 ( .B1(n7283), .B2(n7281), .A(n6621), .ZN(n7280) );
  INV_X1 U7550 ( .A(n7283), .ZN(n7282) );
  INV_X1 U7551 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8521) );
  AND3_X1 U7552 ( .A1(n7122), .A2(n6584), .A3(n7413), .ZN(n8522) );
  INV_X1 U7553 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n7253) );
  AND2_X1 U7554 ( .A1(n7371), .A2(n7370), .ZN(n7919) );
  INV_X1 U7555 ( .A(n8077), .ZN(n6870) );
  XNOR2_X1 U7556 ( .A(n7871), .B(SI_12_), .ZN(n8176) );
  INV_X1 U7557 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n7921) );
  INV_X1 U7558 ( .A(n8006), .ZN(n6788) );
  NAND2_X1 U7559 ( .A1(n6714), .A2(n7843), .ZN(n8003) );
  XNOR2_X1 U7560 ( .A(n13357), .B(P3_ADDR_REG_1__SCAN_IN), .ZN(n13887) );
  NOR2_X1 U7561 ( .A1(n13852), .A2(n13851), .ZN(n13881) );
  NAND2_X1 U7562 ( .A1(n11970), .A2(n6492), .ZN(n11925) );
  INV_X1 U7563 ( .A(n11882), .ZN(n7178) );
  INV_X1 U7564 ( .A(n12434), .ZN(n11964) );
  NAND2_X1 U7565 ( .A1(n11211), .A2(n11210), .ZN(n11238) );
  OR2_X1 U7566 ( .A1(n14042), .A2(n14041), .ZN(n7085) );
  OR2_X1 U7567 ( .A1(n12562), .A2(n12189), .ZN(n7596) );
  AOI22_X1 U7568 ( .A1(n12361), .A2(n12239), .B1(n12267), .B2(n12572), .ZN(
        n12346) );
  INV_X1 U7569 ( .A(n12422), .ZN(n8797) );
  AND3_X1 U7570 ( .A1(n8717), .A2(n8716), .A3(n8715), .ZN(n11212) );
  OAI21_X1 U7571 ( .B1(n14736), .B2(n8973), .A(n12123), .ZN(n11054) );
  NOR2_X1 U7572 ( .A1(n12300), .A2(n7547), .ZN(n7546) );
  INV_X1 U7573 ( .A(n8903), .ZN(n7547) );
  NOR2_X1 U7574 ( .A1(n12393), .A2(n7579), .ZN(n7578) );
  NOR2_X1 U7575 ( .A1(n6461), .A2(n8812), .ZN(n7579) );
  XNOR2_X1 U7576 ( .A(n12400), .B(n12269), .ZN(n12393) );
  OR2_X1 U7577 ( .A1(n12427), .A2(n11964), .ZN(n12063) );
  INV_X1 U7578 ( .A(n12468), .ZN(n7567) );
  AND2_X1 U7579 ( .A1(n9082), .A2(n12636), .ZN(n12253) );
  NAND2_X1 U7580 ( .A1(n12068), .A2(n12069), .ZN(n14837) );
  NAND2_X1 U7581 ( .A1(n7622), .A2(n6462), .ZN(n6639) );
  AOI21_X1 U7582 ( .B1(n8879), .B2(n8878), .A(n6990), .ZN(n8891) );
  AND2_X1 U7583 ( .A1(n11276), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6990) );
  AND2_X1 U7584 ( .A1(n8834), .A2(n7347), .ZN(n7344) );
  INV_X1 U7585 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7618) );
  INV_X1 U7586 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7187) );
  NAND2_X1 U7587 ( .A1(n6920), .A2(n6918), .ZN(n8781) );
  NAND2_X1 U7588 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n6919), .ZN(n6918) );
  OAI21_X1 U7589 ( .B1(n8656), .B2(n8554), .A(n8555), .ZN(n8666) );
  AND2_X1 U7590 ( .A1(n9183), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8554) );
  OR2_X1 U7591 ( .A1(n10949), .A2(n10948), .ZN(n7501) );
  NAND2_X1 U7592 ( .A1(n10755), .A2(n10756), .ZN(n7502) );
  NAND2_X1 U7593 ( .A1(n9804), .A2(n9803), .ZN(n9805) );
  AND2_X1 U7594 ( .A1(n9330), .A2(n9331), .ZN(n9326) );
  INV_X1 U7595 ( .A(n11591), .ZN(n11616) );
  AND2_X1 U7596 ( .A1(n14486), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7362) );
  XNOR2_X1 U7597 ( .A(n12797), .B(n14501), .ZN(n14504) );
  NAND2_X1 U7598 ( .A1(n12844), .A2(n11644), .ZN(n12889) );
  NAND2_X1 U7599 ( .A1(n7425), .A2(n7424), .ZN(n12974) );
  OR2_X1 U7600 ( .A1(n13126), .A2(n12840), .ZN(n7424) );
  AOI21_X1 U7601 ( .B1(n7192), .B2(n7199), .A(n6474), .ZN(n7191) );
  XNOR2_X1 U7602 ( .A(n13126), .B(n12840), .ZN(n12999) );
  AND2_X1 U7603 ( .A1(n6503), .A2(n12861), .ZN(n7204) );
  NAND2_X1 U7604 ( .A1(n7207), .A2(n12832), .ZN(n7206) );
  INV_X1 U7605 ( .A(n12859), .ZN(n7207) );
  NAND2_X1 U7606 ( .A1(n11436), .A2(n11435), .ZN(n13136) );
  AND2_X1 U7607 ( .A1(n7597), .A2(n9121), .ZN(n7475) );
  XNOR2_X1 U7608 ( .A(n9309), .B(P2_IR_REG_30__SCAN_IN), .ZN(n9313) );
  NAND2_X1 U7609 ( .A1(n7216), .A2(n6456), .ZN(n9309) );
  OR2_X1 U7610 ( .A1(n9393), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U7611 ( .A1(n10690), .A2(n10689), .ZN(n7238) );
  NOR2_X1 U7612 ( .A1(n7245), .A2(n9907), .ZN(n7249) );
  INV_X1 U7613 ( .A(n7251), .ZN(n7245) );
  AND2_X1 U7614 ( .A1(n7242), .A2(n13219), .ZN(n7241) );
  OR2_X1 U7615 ( .A1(n13319), .A2(n11847), .ZN(n7242) );
  AND2_X1 U7616 ( .A1(n7237), .A2(n7238), .ZN(n7234) );
  OR2_X1 U7617 ( .A1(n7235), .A2(n7233), .ZN(n7232) );
  INV_X1 U7618 ( .A(n7237), .ZN(n7233) );
  AND2_X1 U7619 ( .A1(n10849), .A2(n7236), .ZN(n7235) );
  NAND2_X1 U7620 ( .A1(n10691), .A2(n7238), .ZN(n7236) );
  NAND2_X1 U7621 ( .A1(n11756), .A2(n11755), .ZN(n11757) );
  OAI21_X1 U7622 ( .B1(n13253), .B2(n6722), .A(n6719), .ZN(n6723) );
  AOI21_X1 U7623 ( .B1(n13301), .B2(n6721), .A(n6720), .ZN(n6719) );
  INV_X1 U7624 ( .A(n13301), .ZN(n6722) );
  NAND2_X1 U7625 ( .A1(n9908), .A2(n9838), .ZN(n11824) );
  AND2_X1 U7626 ( .A1(n9247), .A2(n9154), .ZN(n8043) );
  NAND2_X1 U7627 ( .A1(n7219), .A2(n9239), .ZN(n9908) );
  AND2_X1 U7628 ( .A1(n9234), .A2(n9563), .ZN(n7219) );
  NAND2_X1 U7629 ( .A1(n7308), .A2(n6531), .ZN(n13558) );
  AND2_X1 U7630 ( .A1(n13536), .A2(n8489), .ZN(n13576) );
  OR2_X1 U7631 ( .A1(n13750), .A2(n13520), .ZN(n8489) );
  NAND2_X2 U7632 ( .A1(n8530), .A2(n13828), .ZN(n9247) );
  XNOR2_X1 U7633 ( .A(n13529), .B(n13678), .ZN(n13667) );
  OR2_X1 U7634 ( .A1(n13717), .A2(n13525), .ZN(n7410) );
  NAND2_X1 U7635 ( .A1(n10995), .A2(n10994), .ZN(n11146) );
  NOR2_X1 U7636 ( .A1(n7385), .A2(n10820), .ZN(n7380) );
  NAND2_X1 U7637 ( .A1(n13972), .A2(n13971), .ZN(n7312) );
  AND2_X1 U7638 ( .A1(n9246), .A2(n9543), .ZN(n14087) );
  AND2_X1 U7639 ( .A1(n9565), .A2(n9564), .ZN(n9852) );
  AND2_X1 U7640 ( .A1(n9245), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9243) );
  XNOR2_X1 U7641 ( .A(n8459), .B(n8458), .ZN(n11551) );
  NAND2_X1 U7642 ( .A1(n7266), .A2(n7267), .ZN(n8260) );
  OR2_X1 U7643 ( .A1(n7881), .A2(n7269), .ZN(n7266) );
  INV_X1 U7644 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8202) );
  NAND2_X1 U7645 ( .A1(n9053), .A2(n9052), .ZN(n10073) );
  AND2_X1 U7646 ( .A1(n12698), .A2(n12716), .ZN(n7481) );
  AND2_X1 U7647 ( .A1(n6846), .A2(n6845), .ZN(n14177) );
  INV_X1 U7648 ( .A(n14178), .ZN(n6845) );
  OR2_X1 U7649 ( .A1(n11283), .A2(n11638), .ZN(n6935) );
  NOR2_X1 U7650 ( .A1(n6449), .A2(n11284), .ZN(n6979) );
  AOI22_X1 U7651 ( .A1(n12782), .A2(n6451), .B1(n11301), .B2(n9363), .ZN(
        n11308) );
  AOI21_X1 U7652 ( .B1(n7116), .B2(n7114), .A(n7113), .ZN(n8058) );
  NOR2_X1 U7653 ( .A1(n8039), .A2(n8040), .ZN(n7113) );
  AOI21_X1 U7654 ( .B1(n8039), .B2(n8040), .A(n7115), .ZN(n7114) );
  INV_X1 U7655 ( .A(n8108), .ZN(n7128) );
  INV_X1 U7656 ( .A(n8107), .ZN(n7129) );
  NAND2_X1 U7657 ( .A1(n6549), .A2(n11328), .ZN(n6774) );
  NOR2_X1 U7658 ( .A1(n6549), .A2(n11328), .ZN(n6776) );
  NAND2_X1 U7659 ( .A1(n7528), .A2(n7532), .ZN(n7531) );
  INV_X1 U7660 ( .A(n11333), .ZN(n7532) );
  OAI22_X1 U7661 ( .A1(n8169), .A2(n7124), .B1(n8168), .B2(n7123), .ZN(n8184)
         );
  INV_X1 U7662 ( .A(n8167), .ZN(n7123) );
  NOR2_X1 U7663 ( .A1(n7125), .A2(n8167), .ZN(n7124) );
  NAND2_X1 U7664 ( .A1(n8184), .A2(n8185), .ZN(n8183) );
  MUX2_X1 U7665 ( .A(n8326), .B(n8325), .S(n13709), .Z(n8327) );
  NAND2_X1 U7666 ( .A1(n7130), .A2(n6805), .ZN(n6804) );
  NOR2_X1 U7667 ( .A1(n8240), .A2(n6527), .ZN(n6805) );
  AOI21_X1 U7668 ( .B1(n11397), .B2(n11396), .A(n11395), .ZN(n6957) );
  NAND2_X1 U7669 ( .A1(n7541), .A2(n7542), .ZN(n7540) );
  INV_X1 U7670 ( .A(n11401), .ZN(n7541) );
  MUX2_X1 U7671 ( .A(n13516), .B(n13778), .S(n8017), .Z(n8387) );
  INV_X1 U7672 ( .A(n8375), .ZN(n6994) );
  INV_X1 U7673 ( .A(n8402), .ZN(n6959) );
  INV_X1 U7674 ( .A(n8403), .ZN(n6962) );
  INV_X1 U7675 ( .A(n11429), .ZN(n7544) );
  AND2_X1 U7676 ( .A1(n6590), .A2(n6782), .ZN(n6781) );
  NAND2_X1 U7677 ( .A1(n6494), .A2(n6955), .ZN(n6782) );
  OAI211_X1 U7678 ( .C1(n12325), .C2(n12196), .A(n12312), .B(n12195), .ZN(
        n12201) );
  NOR2_X1 U7679 ( .A1(n6794), .A2(n8451), .ZN(n6792) );
  INV_X1 U7680 ( .A(n8463), .ZN(n7119) );
  INV_X1 U7681 ( .A(n8462), .ZN(n7118) );
  INV_X1 U7682 ( .A(n10032), .ZN(n7097) );
  NAND2_X1 U7683 ( .A1(n6563), .A2(n6470), .ZN(n7553) );
  INV_X1 U7684 ( .A(n12094), .ZN(n6651) );
  NAND2_X1 U7685 ( .A1(n11524), .A2(n11525), .ZN(n7523) );
  NAND2_X1 U7686 ( .A1(n7524), .A2(n7522), .ZN(n7521) );
  INV_X1 U7687 ( .A(n10235), .ZN(n7423) );
  OR2_X1 U7688 ( .A1(n13337), .A2(n13228), .ZN(n11147) );
  INV_X1 U7689 ( .A(n7273), .ZN(n6878) );
  NOR2_X1 U7690 ( .A1(n6603), .A2(n6983), .ZN(n6982) );
  INV_X1 U7691 ( .A(n7878), .ZN(n6983) );
  INV_X1 U7692 ( .A(n8159), .ZN(n7258) );
  INV_X1 U7693 ( .A(n8140), .ZN(n7867) );
  INV_X1 U7694 ( .A(n10837), .ZN(n7146) );
  INV_X1 U7695 ( .A(n11936), .ZN(n6634) );
  INV_X1 U7696 ( .A(n11241), .ZN(n6635) );
  INV_X1 U7697 ( .A(n7067), .ZN(n7063) );
  AND2_X1 U7698 ( .A1(n12240), .A2(n7340), .ZN(n7339) );
  NOR2_X1 U7699 ( .A1(n12310), .A2(n7341), .ZN(n7340) );
  AND2_X1 U7700 ( .A1(n12047), .A2(n12046), .ZN(n12215) );
  NAND2_X1 U7701 ( .A1(n7091), .A2(n7090), .ZN(n7089) );
  NAND2_X1 U7702 ( .A1(n7089), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7087) );
  NAND2_X1 U7703 ( .A1(n9927), .A2(n6520), .ZN(n7695) );
  OR2_X1 U7704 ( .A1(n9961), .A2(n7096), .ZN(n7094) );
  NAND2_X1 U7705 ( .A1(n7097), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7096) );
  OAI21_X1 U7706 ( .B1(n8701), .B2(n14944), .A(n14699), .ZN(n7754) );
  INV_X1 U7707 ( .A(n12432), .ZN(n7556) );
  NAND2_X1 U7708 ( .A1(n10461), .A2(n12087), .ZN(n10662) );
  NAND2_X1 U7709 ( .A1(n6644), .A2(n14775), .ZN(n9048) );
  INV_X1 U7710 ( .A(n12063), .ZN(n7057) );
  NAND2_X1 U7711 ( .A1(n12609), .A2(n12433), .ZN(n7565) );
  INV_X1 U7712 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n8570) );
  INV_X1 U7713 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n8567) );
  INV_X1 U7714 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7609) );
  NOR2_X1 U7715 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7610) );
  NAND2_X1 U7716 ( .A1(n6684), .A2(n6685), .ZN(n6682) );
  INV_X1 U7717 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8556) );
  AND2_X1 U7718 ( .A1(n7487), .A2(n7484), .ZN(n7483) );
  NAND2_X1 U7719 ( .A1(n7490), .A2(n12709), .ZN(n7484) );
  NAND2_X1 U7720 ( .A1(n13083), .A2(n12825), .ZN(n11635) );
  NAND2_X1 U7721 ( .A1(n7077), .A2(n12911), .ZN(n7076) );
  NOR2_X1 U7722 ( .A1(n7078), .A2(n13088), .ZN(n7077) );
  NAND2_X1 U7723 ( .A1(n7436), .A2(n6488), .ZN(n7432) );
  INV_X1 U7724 ( .A(n7191), .ZN(n6738) );
  NAND2_X1 U7725 ( .A1(n7444), .A2(n7457), .ZN(n7443) );
  INV_X1 U7726 ( .A(n7455), .ZN(n7444) );
  INV_X1 U7727 ( .A(n10979), .ZN(n7210) );
  NAND2_X1 U7728 ( .A1(n10984), .A2(n12772), .ZN(n7471) );
  NOR2_X1 U7729 ( .A1(n11659), .A2(n7473), .ZN(n7470) );
  NAND2_X1 U7730 ( .A1(n7466), .A2(n10317), .ZN(n7465) );
  NAND2_X1 U7731 ( .A1(n7463), .A2(n7467), .ZN(n7466) );
  INV_X1 U7732 ( .A(n10240), .ZN(n7467) );
  AND2_X1 U7733 ( .A1(n7422), .A2(n10237), .ZN(n7419) );
  OR2_X1 U7734 ( .A1(n11653), .A2(n7423), .ZN(n7422) );
  NAND2_X1 U7735 ( .A1(n11023), .A2(n7449), .ZN(n7448) );
  INV_X1 U7736 ( .A(n7451), .ZN(n7450) );
  INV_X1 U7737 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n9027) );
  NOR2_X1 U7738 ( .A1(n9264), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9391) );
  OR2_X1 U7739 ( .A1(n9220), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n9228) );
  NOR4_X1 U7740 ( .A1(n13587), .A2(n13628), .A3(n13638), .A4(n8502), .ZN(n8503) );
  NOR2_X1 U7741 ( .A1(n13667), .A2(n7316), .ZN(n7315) );
  INV_X1 U7742 ( .A(n13512), .ZN(n7316) );
  NAND2_X1 U7743 ( .A1(n13799), .A2(n7030), .ZN(n7029) );
  INV_X1 U7744 ( .A(n7032), .ZN(n7030) );
  INV_X1 U7745 ( .A(n13506), .ZN(n6707) );
  XNOR2_X1 U7746 ( .A(n13700), .B(n13709), .ZN(n8491) );
  NAND2_X1 U7747 ( .A1(n7027), .A2(n7026), .ZN(n11000) );
  INV_X1 U7748 ( .A(n10513), .ZN(n7305) );
  INV_X1 U7749 ( .A(n10508), .ZN(n7377) );
  NOR2_X1 U7750 ( .A1(n10511), .A2(n7379), .ZN(n7378) );
  INV_X1 U7751 ( .A(n10408), .ZN(n7379) );
  NOR2_X1 U7752 ( .A1(n11000), .A2(n13337), .ZN(n11159) );
  NAND2_X1 U7753 ( .A1(n8425), .A2(n12662), .ZN(n7286) );
  NOR2_X1 U7754 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n7926) );
  INV_X1 U7755 ( .A(n8396), .ZN(n6868) );
  OAI21_X1 U7756 ( .B1(n7886), .B2(n7272), .A(n7271), .ZN(n7894) );
  AOI21_X1 U7757 ( .B1(n6878), .B2(n6877), .A(n6876), .ZN(n7271) );
  INV_X1 U7758 ( .A(n7892), .ZN(n6876) );
  INV_X1 U7759 ( .A(n7272), .ZN(n6877) );
  AND2_X1 U7760 ( .A1(n7924), .A2(n7923), .ZN(n7925) );
  NOR2_X1 U7761 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n7924) );
  NOR2_X1 U7762 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n7923) );
  NAND2_X1 U7763 ( .A1(n7270), .A2(n7890), .ZN(n8353) );
  XNOR2_X1 U7764 ( .A(n8353), .B(SI_20_), .ZN(n8352) );
  AOI21_X1 U7765 ( .B1(n7852), .B2(n6732), .A(n6731), .ZN(n6730) );
  NOR2_X1 U7766 ( .A1(n7847), .A2(n7837), .ZN(n6873) );
  NAND2_X1 U7767 ( .A1(n7847), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n7838) );
  AOI21_X1 U7768 ( .B1(n7141), .B2(n7140), .A(n7139), .ZN(n13842) );
  AND2_X1 U7769 ( .A1(n14986), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7139) );
  INV_X1 U7770 ( .A(n6969), .ZN(n13845) );
  OAI21_X1 U7771 ( .B1(n13882), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n6495), .ZN(
        n6969) );
  XNOR2_X1 U7772 ( .A(n13845), .B(n6941), .ZN(n13899) );
  INV_X1 U7773 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14913) );
  AOI21_X1 U7774 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n13860), .A(n13859), .ZN(
        n13921) );
  NOR2_X1 U7775 ( .A1(n13876), .A2(n13875), .ZN(n13859) );
  INV_X1 U7776 ( .A(n12665), .ZN(n8943) );
  NAND2_X1 U7777 ( .A1(n10723), .A2(n9066), .ZN(n14671) );
  NOR2_X1 U7778 ( .A1(n11918), .A2(n7156), .ZN(n7155) );
  INV_X1 U7779 ( .A(n12008), .ZN(n7156) );
  OR2_X1 U7780 ( .A1(n11917), .A2(n12264), .ZN(n7153) );
  OR2_X1 U7781 ( .A1(n11918), .A2(n7159), .ZN(n7154) );
  NAND2_X1 U7782 ( .A1(n14671), .A2(n14670), .ZN(n14669) );
  INV_X1 U7783 ( .A(n11928), .ZN(n7179) );
  INV_X1 U7784 ( .A(n11264), .ZN(n7177) );
  INV_X1 U7785 ( .A(n7170), .ZN(n7167) );
  AND3_X1 U7786 ( .A1(n8604), .A2(n8603), .A3(n8602), .ZN(n10013) );
  AND2_X1 U7787 ( .A1(n7162), .A2(n11961), .ZN(n7161) );
  NAND2_X1 U7788 ( .A1(n7166), .A2(n7164), .ZN(n7162) );
  OR2_X1 U7789 ( .A1(n10725), .A2(n10726), .ZN(n10723) );
  NAND2_X1 U7790 ( .A1(n6885), .A2(n6604), .ZN(n7181) );
  AND4_X1 U7791 ( .A1(n8772), .A2(n8771), .A3(n8770), .A4(n8769), .ZN(n12018)
         );
  AND4_X1 U7792 ( .A1(n8675), .A2(n8674), .A3(n8673), .A4(n8672), .ZN(n9071)
         );
  AND4_X1 U7793 ( .A1(n8639), .A2(n8638), .A3(n8637), .A4(n8636), .ZN(n10728)
         );
  XNOR2_X1 U7794 ( .A(n7745), .B(n9667), .ZN(n9661) );
  XNOR2_X1 U7795 ( .A(n7752), .B(n14685), .ZN(n14683) );
  INV_X1 U7796 ( .A(n14718), .ZN(n8701) );
  OR2_X1 U7797 ( .A1(n10675), .A2(n7100), .ZN(n7098) );
  OR2_X1 U7798 ( .A1(n10625), .A2(n11057), .ZN(n7100) );
  INV_X1 U7799 ( .A(n7039), .ZN(n7037) );
  AOI21_X1 U7800 ( .B1(n6460), .B2(n7043), .A(n6544), .ZN(n7039) );
  AND2_X1 U7801 ( .A1(n12063), .A2(n12062), .ZN(n12422) );
  INV_X1 U7802 ( .A(n12271), .ZN(n12419) );
  OAI21_X1 U7803 ( .B1(n10933), .B2(n8971), .A(n8972), .ZN(n14736) );
  NAND2_X1 U7804 ( .A1(n8682), .A2(n9098), .ZN(n8693) );
  NAND2_X1 U7805 ( .A1(n10864), .A2(n8680), .ZN(n10865) );
  AND2_X1 U7806 ( .A1(n8692), .A2(n12119), .ZN(n12227) );
  OAI21_X1 U7807 ( .B1(n8646), .B2(n7586), .A(n7585), .ZN(n10825) );
  AOI21_X1 U7808 ( .B1(n12218), .B2(n7587), .A(n6472), .ZN(n7585) );
  INV_X1 U7809 ( .A(n7587), .ZN(n7586) );
  AND2_X1 U7810 ( .A1(n14748), .A2(n8648), .ZN(n7587) );
  NAND2_X1 U7811 ( .A1(n8646), .A2(n10773), .ZN(n10779) );
  NOR2_X1 U7812 ( .A1(n12281), .A2(n9952), .ZN(n14775) );
  INV_X1 U7813 ( .A(n10112), .ZN(n8994) );
  NAND2_X1 U7814 ( .A1(n7335), .A2(n6623), .ZN(n8988) );
  NAND2_X1 U7815 ( .A1(n8902), .A2(n12009), .ZN(n8903) );
  AOI21_X1 U7816 ( .B1(n12322), .B2(n8889), .A(n7603), .ZN(n12313) );
  INV_X1 U7817 ( .A(n12242), .ZN(n12335) );
  NAND2_X1 U7818 ( .A1(n7044), .A2(n12184), .ZN(n7041) );
  NAND2_X1 U7819 ( .A1(n12350), .A2(n6498), .ZN(n7044) );
  INV_X1 U7820 ( .A(n12239), .ZN(n12360) );
  OAI21_X2 U7821 ( .B1(n12369), .B2(n12168), .A(n12176), .ZN(n12359) );
  INV_X1 U7822 ( .A(n7575), .ZN(n7574) );
  AOI21_X1 U7823 ( .B1(n7575), .B2(n7573), .A(n6548), .ZN(n7572) );
  INV_X1 U7824 ( .A(n7578), .ZN(n7573) );
  AND2_X1 U7825 ( .A1(n12175), .A2(n12176), .ZN(n12371) );
  AOI21_X1 U7826 ( .B1(n7578), .B2(n6461), .A(n6558), .ZN(n7577) );
  NAND2_X1 U7827 ( .A1(n8936), .A2(n12076), .ZN(n14760) );
  AOI21_X1 U7828 ( .B1(n7055), .B2(n7054), .A(n12159), .ZN(n7053) );
  NOR2_X1 U7829 ( .A1(n12422), .A2(n7057), .ZN(n7054) );
  INV_X1 U7830 ( .A(n12423), .ZN(n7052) );
  AND2_X1 U7831 ( .A1(n12414), .A2(n8799), .ZN(n12405) );
  NAND2_X1 U7832 ( .A1(n12423), .A2(n12422), .ZN(n12525) );
  NAND2_X1 U7833 ( .A1(n7565), .A2(n7566), .ZN(n7560) );
  OR2_X1 U7834 ( .A1(n7561), .A2(n7559), .ZN(n7558) );
  INV_X1 U7835 ( .A(n7565), .ZN(n7559) );
  INV_X1 U7836 ( .A(n7562), .ZN(n7561) );
  OAI21_X1 U7837 ( .B1(n12454), .B2(n7563), .A(n8773), .ZN(n7562) );
  NAND2_X1 U7838 ( .A1(n12455), .A2(n12454), .ZN(n12453) );
  NAND2_X1 U7839 ( .A1(n11220), .A2(n12232), .ZN(n11219) );
  AND3_X1 U7840 ( .A1(n8935), .A2(n8934), .A3(n12076), .ZN(n14731) );
  INV_X1 U7841 ( .A(n14760), .ZN(n14730) );
  OAI22_X1 U7842 ( .A1(n12025), .A2(n6696), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(n14963), .ZN(n12041) );
  INV_X1 U7843 ( .A(n12026), .ZN(n6696) );
  NOR2_X1 U7844 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_30__SCAN_IN), .ZN(
        n6891) );
  INV_X1 U7845 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6657) );
  INV_X1 U7846 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U7847 ( .A1(n7349), .A2(n8866), .ZN(n8879) );
  INV_X1 U7848 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7620) );
  XNOR2_X1 U7849 ( .A(n8864), .B(n11514), .ZN(n8865) );
  NAND2_X1 U7850 ( .A1(n6619), .A2(n7347), .ZN(n7343) );
  INV_X1 U7851 ( .A(n7348), .ZN(n7345) );
  NAND2_X1 U7852 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n11871), .ZN(n7348) );
  INV_X1 U7853 ( .A(n7185), .ZN(n7183) );
  NAND2_X1 U7854 ( .A1(n8823), .A2(n10493), .ZN(n6666) );
  NAND2_X1 U7855 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7329), .ZN(n7328) );
  OAI21_X1 U7856 ( .B1(n8781), .B2(n6690), .A(n6688), .ZN(n6691) );
  INV_X1 U7857 ( .A(n6689), .ZN(n6688) );
  NOR2_X1 U7858 ( .A1(n7324), .A2(n10759), .ZN(n7322) );
  XNOR2_X1 U7859 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8699) );
  NAND2_X1 U7860 ( .A1(n8560), .A2(n8559), .ZN(n8700) );
  NOR2_X1 U7861 ( .A1(n7699), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n7705) );
  INV_X1 U7862 ( .A(n8557), .ZN(n6685) );
  NAND2_X1 U7863 ( .A1(n6668), .A2(n8553), .ZN(n8656) );
  NAND2_X1 U7864 ( .A1(n8642), .A2(n8640), .ZN(n6668) );
  INV_X1 U7865 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n8552) );
  INV_X1 U7866 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n6628) );
  NAND2_X1 U7867 ( .A1(n6670), .A2(n8546), .ZN(n8614) );
  XNOR2_X1 U7868 ( .A(n9037), .B(n9036), .ZN(n10910) );
  OR2_X1 U7869 ( .A1(n11722), .A2(n11723), .ZN(n7498) );
  NAND2_X1 U7870 ( .A1(n10754), .A2(n7503), .ZN(n7013) );
  INV_X1 U7871 ( .A(n10083), .ZN(n7008) );
  NOR2_X1 U7872 ( .A1(n7006), .A2(n7005), .ZN(n7004) );
  INV_X1 U7873 ( .A(n9976), .ZN(n7005) );
  NAND2_X1 U7874 ( .A1(n7485), .A2(n7486), .ZN(n7489) );
  INV_X1 U7875 ( .A(n9631), .ZN(n9629) );
  NOR2_X1 U7876 ( .A1(n11182), .A2(n11181), .ZN(n11420) );
  AOI21_X1 U7877 ( .B1(n7012), .B2(n7504), .A(n7010), .ZN(n7009) );
  INV_X1 U7878 ( .A(n11060), .ZN(n7010) );
  INV_X1 U7879 ( .A(n11637), .ZN(n7518) );
  OAI22_X1 U7880 ( .A1(n11681), .A2(n11674), .B1(n11673), .B2(n12819), .ZN(
        n11675) );
  AND4_X1 U7881 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n12881) );
  AND2_X1 U7882 ( .A1(n9313), .A2(n9312), .ZN(n9353) );
  AND2_X1 U7883 ( .A1(n11235), .A2(n9312), .ZN(n9517) );
  NOR2_X1 U7884 ( .A1(n14448), .A2(n14447), .ZN(n14446) );
  INV_X1 U7885 ( .A(n10530), .ZN(n6655) );
  INV_X1 U7886 ( .A(n10888), .ZN(n12796) );
  NOR2_X1 U7887 ( .A1(n14492), .A2(n7360), .ZN(n12797) );
  AND2_X1 U7888 ( .A1(n14497), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7360) );
  NOR2_X1 U7889 ( .A1(n14504), .A2(n14503), .ZN(n14502) );
  NAND2_X1 U7890 ( .A1(n6748), .A2(n6747), .ZN(n12937) );
  AND2_X1 U7891 ( .A1(n12938), .A2(n6504), .ZN(n6747) );
  NAND2_X1 U7892 ( .A1(n12968), .A2(n13110), .ZN(n12951) );
  NAND2_X1 U7893 ( .A1(n6897), .A2(n6896), .ZN(n12949) );
  OR2_X1 U7894 ( .A1(n13116), .A2(n12877), .ZN(n6896) );
  NAND2_X1 U7895 ( .A1(n12960), .A2(n6516), .ZN(n6897) );
  OR2_X1 U7896 ( .A1(n12949), .A2(n12950), .ZN(n6748) );
  XNOR2_X1 U7897 ( .A(n12879), .B(n12878), .ZN(n12950) );
  NOR2_X1 U7898 ( .A1(n12984), .A2(n12875), .ZN(n12960) );
  AND2_X1 U7899 ( .A1(n13121), .A2(n12874), .ZN(n12875) );
  NAND2_X1 U7900 ( .A1(n13041), .A2(n7192), .ZN(n6739) );
  NAND2_X1 U7901 ( .A1(n13043), .A2(n13042), .ZN(n13041) );
  AOI21_X1 U7902 ( .B1(n7447), .B2(n7446), .A(n7445), .ZN(n7437) );
  OR2_X1 U7903 ( .A1(n13156), .A2(n12856), .ZN(n12857) );
  OR2_X1 U7904 ( .A1(n11044), .A2(n6753), .ZN(n11046) );
  INV_X1 U7905 ( .A(n11043), .ZN(n6753) );
  OR2_X1 U7906 ( .A1(n11394), .A2(n11021), .ZN(n7460) );
  NAND2_X1 U7907 ( .A1(n10747), .A2(n10746), .ZN(n10749) );
  NAND2_X1 U7908 ( .A1(n7213), .A2(n11659), .ZN(n10980) );
  INV_X1 U7909 ( .A(n10749), .ZN(n7213) );
  NAND2_X1 U7910 ( .A1(n10423), .A2(n10440), .ZN(n10735) );
  XNOR2_X1 U7911 ( .A(n14638), .B(n10314), .ZN(n11657) );
  XNOR2_X1 U7912 ( .A(n11356), .B(n12775), .ZN(n7463) );
  NAND2_X1 U7913 ( .A1(n10255), .A2(n10240), .ZN(n10241) );
  NAND2_X1 U7914 ( .A1(n10230), .A2(n6528), .ZN(n10252) );
  NAND2_X1 U7915 ( .A1(n10207), .A2(n11653), .ZN(n10236) );
  NAND2_X1 U7916 ( .A1(n6716), .A2(n10138), .ZN(n10218) );
  NAND2_X1 U7917 ( .A1(n6749), .A2(n10046), .ZN(n10164) );
  AND2_X1 U7918 ( .A1(n10060), .A2(n10047), .ZN(n11647) );
  AOI211_X1 U7919 ( .C1(n13088), .C2(n12895), .A(n9339), .B(n12852), .ZN(
        n13087) );
  NAND2_X1 U7920 ( .A1(n11586), .A2(n11585), .ZN(n13096) );
  NAND2_X1 U7921 ( .A1(n13204), .A2(n11584), .ZN(n11586) );
  NAND2_X1 U7922 ( .A1(n11538), .A2(n11537), .ZN(n13100) );
  NAND2_X1 U7923 ( .A1(n11467), .A2(n11466), .ZN(n13126) );
  NAND2_X1 U7924 ( .A1(n10762), .A2(n10761), .ZN(n13167) );
  AND2_X1 U7925 ( .A1(n9271), .A2(n13207), .ZN(n14558) );
  NAND2_X1 U7926 ( .A1(n9034), .A2(n9036), .ZN(n9029) );
  OR2_X1 U7927 ( .A1(n9029), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n9032) );
  OAI21_X1 U7928 ( .B1(n9289), .B2(n7024), .A(n7022), .ZN(n9109) );
  NAND2_X1 U7929 ( .A1(n13197), .A2(n7023), .ZN(n7022) );
  NAND2_X1 U7930 ( .A1(n6456), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n7024) );
  OR2_X1 U7931 ( .A1(n9181), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n9827) );
  OR2_X1 U7932 ( .A1(n9719), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9693) );
  AND2_X1 U7933 ( .A1(n9162), .A2(n9155), .ZN(n9830) );
  NAND2_X1 U7934 ( .A1(n7244), .A2(n6529), .ZN(n13223) );
  NAND2_X1 U7935 ( .A1(n11739), .A2(n11738), .ZN(n7244) );
  AOI21_X1 U7936 ( .B1(n13286), .B2(n7224), .A(n11830), .ZN(n7223) );
  INV_X1 U7937 ( .A(n11822), .ZN(n7224) );
  INV_X1 U7938 ( .A(n13286), .ZN(n7225) );
  NAND2_X1 U7939 ( .A1(n11774), .A2(n13274), .ZN(n13276) );
  NAND2_X1 U7940 ( .A1(n7248), .A2(n7247), .ZN(n10301) );
  AOI21_X1 U7941 ( .B1(n7249), .B2(n9904), .A(n6561), .ZN(n7247) );
  NAND2_X1 U7942 ( .A1(n9905), .A2(n7249), .ZN(n7248) );
  AND2_X1 U7943 ( .A1(n6756), .A2(n10852), .ZN(n7229) );
  INV_X1 U7944 ( .A(n7234), .ZN(n7230) );
  INV_X1 U7945 ( .A(n7232), .ZN(n7231) );
  NOR2_X1 U7946 ( .A1(n8115), .A2(n9532), .ZN(n8134) );
  OAI211_X1 U7947 ( .C1(n11824), .C2(n10611), .A(n9842), .B(n9841), .ZN(n9880)
         );
  OR2_X1 U7948 ( .A1(n11823), .A2(n9840), .ZN(n9841) );
  INV_X1 U7949 ( .A(n11135), .ZN(n6746) );
  NAND2_X1 U7950 ( .A1(n7243), .A2(n6525), .ZN(n13253) );
  NAND2_X1 U7951 ( .A1(n11102), .A2(n11101), .ZN(n7226) );
  NAND2_X1 U7952 ( .A1(n10555), .A2(n10554), .ZN(n6757) );
  NAND2_X1 U7953 ( .A1(n8429), .A2(n8428), .ZN(n13491) );
  OAI21_X1 U7954 ( .B1(n8484), .B2(n8483), .A(n8482), .ZN(n8485) );
  AND2_X1 U7955 ( .A1(n8337), .A2(n8336), .ZN(n13528) );
  AND2_X1 U7956 ( .A1(n8219), .A2(n8218), .ZN(n13966) );
  AND4_X1 U7957 ( .A1(n8031), .A2(n8030), .A3(n8029), .A4(n8028), .ZN(n10370)
         );
  NAND2_X1 U7958 ( .A1(n7938), .A2(n7937), .ZN(n7958) );
  INV_X1 U7959 ( .A(n13555), .ZN(n13559) );
  NAND2_X1 U7960 ( .A1(n13582), .A2(n13520), .ZN(n7307) );
  OR2_X1 U7961 ( .A1(n7390), .A2(n13555), .ZN(n7389) );
  NAND2_X1 U7962 ( .A1(n13556), .A2(n14087), .ZN(n7387) );
  AND2_X1 U7963 ( .A1(n8453), .A2(n8439), .ZN(n13579) );
  NOR2_X1 U7964 ( .A1(n13576), .A2(n7310), .ZN(n7306) );
  NAND2_X1 U7965 ( .A1(n13535), .A2(n8490), .ZN(n13587) );
  OR2_X1 U7966 ( .A1(n13491), .A2(n15021), .ZN(n8490) );
  NAND2_X1 U7967 ( .A1(n13767), .A2(n6523), .ZN(n13588) );
  NAND2_X1 U7968 ( .A1(n13588), .A2(n13587), .ZN(n13586) );
  NAND2_X1 U7969 ( .A1(n13780), .A2(n7319), .ZN(n13627) );
  NOR2_X1 U7970 ( .A1(n13623), .A2(n7320), .ZN(n7319) );
  INV_X1 U7971 ( .A(n13517), .ZN(n7320) );
  NOR2_X1 U7972 ( .A1(n7399), .A2(n6465), .ZN(n7398) );
  INV_X1 U7973 ( .A(n13667), .ZN(n7399) );
  OR2_X1 U7974 ( .A1(n6564), .A2(n6465), .ZN(n7397) );
  INV_X1 U7975 ( .A(n13668), .ZN(n6823) );
  OR2_X1 U7976 ( .A1(n13683), .A2(n13684), .ZN(n13681) );
  INV_X1 U7977 ( .A(n7405), .ZN(n7404) );
  AOI21_X1 U7978 ( .B1(n7406), .B2(n13526), .A(n7409), .ZN(n7405) );
  AND2_X1 U7979 ( .A1(n13700), .A2(n13527), .ZN(n7409) );
  NOR2_X1 U7980 ( .A1(n13701), .A2(n7407), .ZN(n7406) );
  INV_X1 U7981 ( .A(n7410), .ZN(n7407) );
  INV_X1 U7982 ( .A(n8491), .ZN(n13701) );
  NAND2_X1 U7983 ( .A1(n8312), .A2(n8311), .ZN(n13717) );
  NAND2_X1 U7984 ( .A1(n11157), .A2(n6709), .ZN(n6708) );
  NOR2_X1 U7985 ( .A1(n13504), .A2(n6710), .ZN(n6709) );
  INV_X1 U7986 ( .A(n11156), .ZN(n6710) );
  NAND2_X1 U7987 ( .A1(n14139), .A2(n6524), .ZN(n11155) );
  NAND2_X1 U7988 ( .A1(n6698), .A2(n10818), .ZN(n13972) );
  NAND2_X1 U7989 ( .A1(n10409), .A2(n7378), .ZN(n10509) );
  INV_X1 U7990 ( .A(n10407), .ZN(n10448) );
  NAND2_X1 U7991 ( .A1(n10374), .A2(n10384), .ZN(n7299) );
  INV_X1 U7992 ( .A(n10384), .ZN(n14291) );
  AND3_X1 U7993 ( .A1(n8010), .A2(n8009), .A3(n8008), .ZN(n10367) );
  NAND2_X2 U7994 ( .A1(n8449), .A2(n8448), .ZN(n13750) );
  INV_X1 U7995 ( .A(n13522), .ZN(n14116) );
  NAND2_X1 U7996 ( .A1(n11159), .A2(n14128), .ZN(n14124) );
  NAND2_X1 U7997 ( .A1(n6752), .A2(n8414), .ZN(n8095) );
  INV_X1 U7998 ( .A(n9977), .ZN(n6752) );
  NAND2_X1 U7999 ( .A1(n9549), .A2(n9548), .ZN(n14373) );
  AND2_X1 U8000 ( .A1(n6819), .A2(n6818), .ZN(n6816) );
  NAND2_X1 U8001 ( .A1(n8043), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n6818) );
  OR2_X1 U8002 ( .A1(n14352), .A2(n10114), .ZN(n10362) );
  NAND2_X1 U8003 ( .A1(n9236), .A2(n9563), .ZN(n9566) );
  NAND2_X1 U8004 ( .A1(n7913), .A2(n7289), .ZN(n8468) );
  AND2_X1 U8005 ( .A1(n7912), .A2(n7291), .ZN(n7289) );
  XNOR2_X1 U8006 ( .A(n8518), .B(n8521), .ZN(n9245) );
  XNOR2_X1 U8007 ( .A(n7894), .B(n6953), .ZN(n7893) );
  AND2_X1 U8008 ( .A1(n7948), .A2(n7255), .ZN(n7254) );
  XNOR2_X1 U8009 ( .A(n8292), .B(n8291), .ZN(n11432) );
  OR2_X1 U8010 ( .A1(n8266), .A2(P1_IR_REG_17__SCAN_IN), .ZN(n8307) );
  OR2_X1 U8011 ( .A1(n8222), .A2(SI_14_), .ZN(n6924) );
  OR2_X1 U8012 ( .A1(n8178), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8179) );
  OR2_X1 U8013 ( .A1(n6989), .A2(n7260), .ZN(n7256) );
  NAND2_X1 U8014 ( .A1(n8077), .A2(n7863), .ZN(n6989) );
  NOR2_X1 U8015 ( .A1(n9671), .A2(P1_ADDR_REG_0__SCAN_IN), .ZN(n13889) );
  NAND2_X1 U8016 ( .A1(n13896), .A2(n13897), .ZN(n13901) );
  XNOR2_X1 U8017 ( .A(n13899), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n13900) );
  NAND2_X1 U8018 ( .A1(n7137), .A2(n13906), .ZN(n13908) );
  NAND2_X1 U8019 ( .A1(n13945), .A2(n13944), .ZN(n7137) );
  INV_X1 U8020 ( .A(n6844), .ZN(n13916) );
  OAI21_X1 U8021 ( .B1(n13946), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6508), .ZN(
        n6844) );
  OAI21_X1 U8022 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14698), .A(n13856), .ZN(
        n13878) );
  AOI21_X1 U8023 ( .B1(n13920), .B2(n13919), .A(n14172), .ZN(n13923) );
  OR2_X1 U8024 ( .A1(n14184), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n13930) );
  INV_X1 U8025 ( .A(n14185), .ZN(n13929) );
  NAND2_X1 U8026 ( .A1(n6831), .A2(n6830), .ZN(n13936) );
  NAND2_X1 U8027 ( .A1(n13984), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6830) );
  AND2_X1 U8028 ( .A1(n8856), .A2(n8855), .ZN(n12178) );
  AND2_X1 U8029 ( .A1(n11070), .A2(n11068), .ZN(n7182) );
  NAND2_X1 U8030 ( .A1(n7173), .A2(n6630), .ZN(n10455) );
  AOI21_X1 U8031 ( .B1(n7174), .B2(n10072), .A(n6538), .ZN(n7173) );
  NAND2_X1 U8032 ( .A1(n10073), .A2(n7174), .ZN(n6630) );
  AND3_X1 U8033 ( .A1(n8645), .A2(n8644), .A3(n8643), .ZN(n10775) );
  AOI21_X1 U8034 ( .B1(n9590), .B2(n12042), .A(n8776), .ZN(n11969) );
  AND3_X1 U8035 ( .A1(n8832), .A2(n8831), .A3(n8830), .ZN(n12396) );
  NAND2_X1 U8036 ( .A1(n11910), .A2(n11258), .ZN(n11972) );
  AND4_X1 U8037 ( .A1(n8725), .A2(n8724), .A3(n8723), .A4(n8722), .ZN(n11985)
         );
  NAND2_X1 U8038 ( .A1(n9092), .A2(n14785), .ZN(n14675) );
  INV_X1 U8039 ( .A(n14731), .ZN(n14762) );
  INV_X1 U8040 ( .A(n12068), .ZN(n12256) );
  NAND2_X1 U8041 ( .A1(n8843), .A2(n8842), .ZN(n12363) );
  OR2_X1 U8042 ( .A1(n8796), .A2(n8795), .ZN(n12434) );
  INV_X1 U8043 ( .A(n12018), .ZN(n12433) );
  AND4_X1 U8044 ( .A1(n8543), .A2(n8542), .A3(n8541), .A4(n8540), .ZN(n12468)
         );
  XNOR2_X1 U8045 ( .A(n7748), .B(n9964), .ZN(n9959) );
  NOR2_X1 U8046 ( .A1(n14024), .A2(n7722), .ZN(n14042) );
  NAND2_X1 U8047 ( .A1(n8816), .A2(n8815), .ZN(n12400) );
  NAND2_X1 U8048 ( .A1(n8788), .A2(n8787), .ZN(n12427) );
  XNOR2_X1 U8049 ( .A(n6653), .B(n12241), .ZN(n9014) );
  AOI21_X1 U8050 ( .B1(n12311), .B2(n7067), .A(n7064), .ZN(n6653) );
  INV_X1 U8051 ( .A(n8988), .ZN(n9013) );
  NAND2_X1 U8052 ( .A1(n8848), .A2(n8847), .ZN(n12572) );
  OR2_X1 U8053 ( .A1(n12043), .A2(n10645), .ZN(n8847) );
  NAND2_X1 U8054 ( .A1(n8836), .A2(n8835), .ZN(n12578) );
  INV_X1 U8055 ( .A(n12154), .ZN(n12609) );
  NAND2_X1 U8056 ( .A1(n12751), .A2(n6486), .ZN(n12669) );
  NAND2_X1 U8057 ( .A1(n10592), .A2(n10591), .ZN(n13172) );
  NAND2_X1 U8058 ( .A1(n12715), .A2(n11717), .ZN(n12699) );
  NAND2_X1 U8059 ( .A1(n12698), .A2(n11716), .ZN(n7480) );
  INV_X1 U8060 ( .A(n7489), .ZN(n12708) );
  NAND2_X1 U8061 ( .A1(n11410), .A2(n11409), .ZN(n13146) );
  NAND2_X1 U8062 ( .A1(n11711), .A2(n11710), .ZN(n11712) );
  NAND2_X1 U8063 ( .A1(n12717), .A2(n12716), .ZN(n12715) );
  NAND2_X1 U8064 ( .A1(n11419), .A2(n11418), .ZN(n13141) );
  NAND2_X1 U8065 ( .A1(n9307), .A2(n13071), .ZN(n12747) );
  INV_X1 U8066 ( .A(n12881), .ZN(n12882) );
  INV_X1 U8067 ( .A(n12701), .ZN(n12878) );
  OAI21_X1 U8068 ( .B1(n13008), .B2(n11459), .A(n11458), .ZN(n12869) );
  OAI21_X1 U8069 ( .B1(n13023), .B2(n11459), .A(n11443), .ZN(n12867) );
  INV_X1 U8070 ( .A(n14459), .ZN(n6640) );
  NOR2_X1 U8071 ( .A1(n14468), .A2(n14467), .ZN(n14466) );
  NOR2_X1 U8072 ( .A1(n14482), .A2(n14483), .ZN(n14481) );
  NOR2_X1 U8073 ( .A1(n14494), .A2(n14493), .ZN(n14492) );
  NAND2_X1 U8074 ( .A1(n14522), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7353) );
  NAND2_X1 U8075 ( .A1(n14522), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7351) );
  AOI21_X1 U8076 ( .B1(n14442), .B2(P2_ADDR_REG_19__SCAN_IN), .A(n12820), .ZN(
        n7367) );
  NAND2_X1 U8077 ( .A1(n12817), .A2(n12814), .ZN(n6665) );
  NAND2_X1 U8078 ( .A1(n13087), .A2(n13078), .ZN(n6944) );
  INV_X1 U8079 ( .A(n12887), .ZN(n7218) );
  AND2_X1 U8080 ( .A1(n7078), .A2(n12884), .ZN(n6907) );
  AND2_X1 U8081 ( .A1(n11489), .A2(n11488), .ZN(n12981) );
  AND2_X1 U8082 ( .A1(n9117), .A2(n7215), .ZN(n7214) );
  INV_X1 U8083 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7215) );
  OAI21_X1 U8084 ( .B1(n13318), .B2(n11847), .A(n7241), .ZN(n13217) );
  AOI21_X1 U8085 ( .B1(n13319), .B2(n11838), .A(n11847), .ZN(n6741) );
  NAND2_X1 U8086 ( .A1(n8214), .A2(n8213), .ZN(n14136) );
  NAND2_X1 U8087 ( .A1(n8146), .A2(n8145), .ZN(n10976) );
  NAND2_X1 U8088 ( .A1(n11551), .A2(n8460), .ZN(n6860) );
  NOR2_X1 U8089 ( .A1(n9885), .A2(n9884), .ZN(n9893) );
  NAND2_X1 U8090 ( .A1(n8360), .A2(n8359), .ZN(n13529) );
  NAND2_X1 U8091 ( .A1(n8251), .A2(n8250), .ZN(n14089) );
  AND2_X1 U8092 ( .A1(n8128), .A2(n8127), .ZN(n14412) );
  NAND2_X1 U8093 ( .A1(n8206), .A2(n8205), .ZN(n14145) );
  INV_X1 U8094 ( .A(n13491), .ZN(n13756) );
  INV_X1 U8095 ( .A(n14078), .ZN(n13320) );
  AND2_X1 U8096 ( .A1(n8515), .A2(n8514), .ZN(n6853) );
  INV_X1 U8097 ( .A(n8485), .ZN(n6798) );
  NAND2_X1 U8098 ( .A1(n8259), .A2(n8258), .ZN(n14086) );
  INV_X1 U8099 ( .A(n10114), .ZN(n13486) );
  NAND2_X1 U8100 ( .A1(n6496), .A2(n6473), .ZN(n13817) );
  NAND2_X1 U8101 ( .A1(n15036), .A2(n15037), .ZN(n13891) );
  INV_X1 U8102 ( .A(n7141), .ZN(n13886) );
  XNOR2_X1 U8103 ( .A(n13916), .B(n7143), .ZN(n13952) );
  INV_X1 U8104 ( .A(n13917), .ZN(n7143) );
  NAND2_X1 U8105 ( .A1(n13952), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7142) );
  AOI21_X1 U8106 ( .B1(n13926), .B2(n13925), .A(n14177), .ZN(n14182) );
  INV_X1 U8107 ( .A(n14181), .ZN(n6905) );
  NAND3_X1 U8108 ( .A1(n13930), .A2(n7136), .A3(n13929), .ZN(n7135) );
  INV_X1 U8109 ( .A(n13933), .ZN(n7136) );
  NAND2_X1 U8110 ( .A1(n7135), .A2(n14525), .ZN(n6832) );
  NOR2_X1 U8111 ( .A1(n14188), .A2(n6833), .ZN(n6829) );
  INV_X1 U8112 ( .A(n6832), .ZN(n6834) );
  AND2_X1 U8113 ( .A1(n13936), .A2(n13937), .ZN(n13986) );
  NOR2_X1 U8114 ( .A1(n11289), .A2(n11288), .ZN(n6980) );
  INV_X1 U8115 ( .A(n8023), .ZN(n7115) );
  OAI211_X1 U8116 ( .C1(n7129), .C2(n7128), .A(n8060), .B(n8059), .ZN(n6810)
         );
  AND2_X1 U8117 ( .A1(n8105), .A2(n10407), .ZN(n6809) );
  NAND2_X1 U8118 ( .A1(n7128), .A2(n7129), .ZN(n6808) );
  INV_X1 U8119 ( .A(n7530), .ZN(n7529) );
  AND2_X1 U8120 ( .A1(n7530), .A2(n11342), .ZN(n7526) );
  AND2_X1 U8121 ( .A1(n6773), .A2(n11348), .ZN(n6772) );
  INV_X1 U8122 ( .A(n6547), .ZN(n6773) );
  NAND2_X1 U8123 ( .A1(n6917), .A2(n6547), .ZN(n6771) );
  INV_X1 U8124 ( .A(n11353), .ZN(n7538) );
  INV_X1 U8125 ( .A(n8168), .ZN(n7125) );
  NAND2_X1 U8126 ( .A1(n12076), .A2(n12077), .ZN(n6645) );
  INV_X1 U8127 ( .A(n6644), .ZN(n6646) );
  NAND2_X1 U8128 ( .A1(n8209), .A2(n8207), .ZN(n7134) );
  INV_X1 U8129 ( .A(n7132), .ZN(n7131) );
  OAI21_X1 U8130 ( .B1(n6787), .B2(n6786), .A(n6551), .ZN(n11385) );
  OAI21_X1 U8131 ( .B1(n11371), .B2(n11370), .A(n6556), .ZN(n6787) );
  AOI21_X1 U8132 ( .B1(n11371), .B2(n11370), .A(n11369), .ZN(n6786) );
  INV_X1 U8133 ( .A(n8340), .ZN(n7112) );
  AND2_X1 U8134 ( .A1(n11407), .A2(n6466), .ZN(n6780) );
  NAND2_X1 U8135 ( .A1(n8386), .A2(n8388), .ZN(n7126) );
  NAND2_X1 U8136 ( .A1(n6961), .A2(n6960), .ZN(n8402) );
  NAND2_X1 U8137 ( .A1(n13607), .A2(n8271), .ZN(n6960) );
  NAND2_X1 U8138 ( .A1(n13772), .A2(n8399), .ZN(n6961) );
  NAND2_X1 U8139 ( .A1(n6813), .A2(n8416), .ZN(n6812) );
  NAND2_X1 U8140 ( .A1(n11463), .A2(n6513), .ZN(n7534) );
  OAI21_X1 U8141 ( .B1(n11447), .B2(n6783), .A(n6781), .ZN(n6784) );
  NOR2_X1 U8142 ( .A1(n6494), .A2(n6955), .ZN(n6783) );
  INV_X1 U8143 ( .A(n8461), .ZN(n6862) );
  AOI21_X1 U8144 ( .B1(n8461), .B2(n6455), .A(n8271), .ZN(n6861) );
  NAND2_X1 U8145 ( .A1(n13547), .A2(n8271), .ZN(n6863) );
  INV_X1 U8146 ( .A(n8261), .ZN(n7883) );
  NOR2_X1 U8147 ( .A1(n7511), .A2(n11498), .ZN(n6785) );
  NAND2_X1 U8148 ( .A1(n11526), .A2(n7525), .ZN(n7524) );
  INV_X1 U8149 ( .A(n11511), .ZN(n7522) );
  NAND2_X1 U8150 ( .A1(n12242), .A2(n12350), .ZN(n7341) );
  INV_X1 U8151 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7616) );
  INV_X1 U8152 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7615) );
  INV_X1 U8153 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n8564) );
  INV_X1 U8154 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8563) );
  AND2_X1 U8155 ( .A1(n12683), .A2(n6507), .ZN(n7487) );
  NAND2_X1 U8156 ( .A1(n12833), .A2(n12856), .ZN(n7459) );
  OR2_X1 U8157 ( .A1(n11755), .A2(n6729), .ZN(n6728) );
  INV_X1 U8158 ( .A(n13330), .ZN(n6729) );
  NAND3_X1 U8159 ( .A1(n7117), .A2(n6791), .A3(n6533), .ZN(n8466) );
  NAND2_X1 U8160 ( .A1(n9546), .A2(n9544), .ZN(n8477) );
  NOR2_X1 U8161 ( .A1(n13592), .A2(n13750), .ZN(n6826) );
  NOR2_X1 U8162 ( .A1(n7284), .A2(n7906), .ZN(n7283) );
  INV_X1 U8163 ( .A(n7286), .ZN(n7284) );
  INV_X1 U8164 ( .A(n6612), .ZN(n7281) );
  NAND2_X1 U8165 ( .A1(n6610), .A2(n7890), .ZN(n7272) );
  INV_X1 U8166 ( .A(n8291), .ZN(n6895) );
  INV_X1 U8167 ( .A(n7850), .ZN(n6732) );
  INV_X1 U8168 ( .A(n7853), .ZN(n6731) );
  NAND2_X1 U8169 ( .A1(n7847), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6986) );
  INV_X1 U8170 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7274) );
  INV_X1 U8171 ( .A(n6842), .ZN(n13844) );
  OAI21_X1 U8172 ( .B1(n13894), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n6464), .ZN(
        n6842) );
  INV_X1 U8173 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n13843) );
  NOR2_X1 U8174 ( .A1(n7093), .A2(n6552), .ZN(n7092) );
  INV_X1 U8175 ( .A(n7095), .ZN(n7093) );
  NAND2_X1 U8176 ( .A1(n10627), .A2(n6931), .ZN(n7757) );
  NAND2_X1 U8177 ( .A1(n10633), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6931) );
  NAND2_X1 U8178 ( .A1(n14004), .A2(n6933), .ZN(n7761) );
  OR2_X1 U8179 ( .A1(n13998), .A2(n12532), .ZN(n6933) );
  INV_X1 U8180 ( .A(n12266), .ZN(n12189) );
  NAND2_X1 U8181 ( .A1(n14758), .A2(n14759), .ZN(n7548) );
  NAND2_X1 U8182 ( .A1(n10665), .A2(n10469), .ZN(n12086) );
  AND3_X1 U8183 ( .A1(n8617), .A2(n8616), .A3(n8615), .ZN(n9054) );
  NAND2_X1 U8184 ( .A1(n10463), .A2(n10013), .ZN(n12080) );
  INV_X1 U8185 ( .A(n12200), .ZN(n7066) );
  INV_X1 U8186 ( .A(n7053), .ZN(n7049) );
  NAND2_X1 U8187 ( .A1(n7549), .A2(n7553), .ZN(n12465) );
  NAND2_X1 U8188 ( .A1(n11220), .A2(n6593), .ZN(n7549) );
  NAND2_X1 U8189 ( .A1(n6649), .A2(n6647), .ZN(n14743) );
  AOI21_X1 U8190 ( .B1(n12218), .B2(n6651), .A(n6648), .ZN(n6647) );
  INV_X1 U8191 ( .A(n12097), .ZN(n6648) );
  OR2_X1 U8192 ( .A1(n8946), .A2(P3_D_REG_0__SCAN_IN), .ZN(n7189) );
  INV_X1 U8193 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7730) );
  AOI21_X1 U8194 ( .B1(n7342), .B2(n6616), .A(n7350), .ZN(n8864) );
  AND2_X1 U8195 ( .A1(n11500), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7350) );
  INV_X1 U8196 ( .A(n8857), .ZN(n6695) );
  NAND2_X1 U8197 ( .A1(n11487), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U8198 ( .A1(n7327), .A2(n7325), .ZN(n8822) );
  NAND2_X1 U8199 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n7326), .ZN(n7325) );
  INV_X1 U8200 ( .A(n8783), .ZN(n6690) );
  OAI21_X1 U8201 ( .B1(n8782), .B2(n6690), .A(n8801), .ZN(n6689) );
  INV_X1 U8202 ( .A(n8571), .ZN(n6676) );
  NAND2_X1 U8203 ( .A1(n8746), .A2(n8760), .ZN(n6677) );
  INV_X1 U8204 ( .A(n8562), .ZN(n7334) );
  INV_X1 U8205 ( .A(n8559), .ZN(n6694) );
  OR2_X1 U8206 ( .A1(n7688), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n7693) );
  AOI21_X1 U8207 ( .B1(n7018), .B2(n7020), .A(n6512), .ZN(n7015) );
  AND2_X1 U8208 ( .A1(n6976), .A2(n6972), .ZN(n6971) );
  AND2_X1 U8209 ( .A1(n11555), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n11556) );
  NOR2_X1 U8210 ( .A1(n11394), .A2(n13167), .ZN(n6750) );
  NAND2_X1 U8211 ( .A1(n10271), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10425) );
  INV_X1 U8212 ( .A(n7432), .ZN(n7431) );
  NAND2_X1 U8213 ( .A1(n7434), .A2(n7436), .ZN(n7433) );
  AOI22_X1 U8214 ( .A1(n12974), .A2(n12982), .B1(n12981), .B2(n12874), .ZN(
        n12962) );
  NOR2_X1 U8215 ( .A1(n10327), .A2(n14638), .ZN(n10435) );
  INV_X1 U8216 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9036) );
  INV_X1 U8217 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9022) );
  INV_X1 U8218 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6760) );
  NOR2_X2 U8219 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9104) );
  INV_X1 U8220 ( .A(n7398), .ZN(n7392) );
  AND2_X1 U8221 ( .A1(n13778), .A2(n13532), .ZN(n7402) );
  NOR2_X1 U8222 ( .A1(n6485), .A2(n7383), .ZN(n7382) );
  INV_X1 U8223 ( .A(n10808), .ZN(n7383) );
  NOR2_X1 U8224 ( .A1(n13975), .A2(n6485), .ZN(n7385) );
  NAND2_X1 U8225 ( .A1(n10399), .A2(n10374), .ZN(n6704) );
  INV_X1 U8226 ( .A(n13349), .ZN(n10561) );
  NAND2_X1 U8227 ( .A1(n7294), .A2(n7296), .ZN(n7293) );
  NAND2_X1 U8228 ( .A1(n13354), .A2(n14351), .ZN(n9703) );
  NAND2_X1 U8229 ( .A1(n6826), .A2(n6825), .ZN(n13561) );
  INV_X1 U8230 ( .A(n6826), .ZN(n13577) );
  NAND2_X1 U8231 ( .A1(n10809), .A2(n10808), .ZN(n13976) );
  NAND2_X1 U8232 ( .A1(n13486), .A2(n7954), .ZN(n9546) );
  NAND2_X1 U8233 ( .A1(n6827), .A2(n14367), .ZN(n10650) );
  NAND2_X1 U8234 ( .A1(n8005), .A2(n7983), .ZN(n6819) );
  NAND2_X1 U8235 ( .A1(n6624), .A2(n7321), .ZN(n10614) );
  INV_X1 U8236 ( .A(n13835), .ZN(n9563) );
  OAI21_X1 U8237 ( .B1(n8459), .B2(n8458), .A(n7910), .ZN(n7970) );
  OR2_X1 U8238 ( .A1(n8305), .A2(n6875), .ZN(n7886) );
  INV_X1 U8239 ( .A(n8306), .ZN(n6875) );
  MUX2_X1 U8240 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n9154), .Z(n8306) );
  XNOR2_X1 U8241 ( .A(n7884), .B(SI_18_), .ZN(n8305) );
  AOI21_X1 U8242 ( .B1(n8246), .B2(n7268), .A(n6550), .ZN(n7267) );
  INV_X1 U8243 ( .A(n7880), .ZN(n7268) );
  INV_X1 U8244 ( .A(n8246), .ZN(n7269) );
  INV_X1 U8245 ( .A(n8210), .ZN(n8223) );
  XNOR2_X1 U8246 ( .A(n8221), .B(SI_14_), .ZN(n8220) );
  XNOR2_X1 U8247 ( .A(n7874), .B(SI_13_), .ZN(n8197) );
  INV_X1 U8248 ( .A(n7261), .ZN(n7260) );
  AOI21_X1 U8249 ( .B1(n7261), .B2(n7865), .A(n6555), .ZN(n7259) );
  NAND2_X1 U8250 ( .A1(n6854), .A2(SI_1_), .ZN(n6856) );
  INV_X1 U8251 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n13841) );
  XNOR2_X1 U8252 ( .A(n13844), .B(n13843), .ZN(n13882) );
  AOI21_X1 U8253 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n13855), .A(n13854), .ZN(
        n13914) );
  NOR2_X1 U8254 ( .A1(n13881), .A2(n13880), .ZN(n13854) );
  INV_X1 U8255 ( .A(n14188), .ZN(n6828) );
  OR2_X1 U8256 ( .A1(n12014), .A2(n12468), .ZN(n7170) );
  INV_X1 U8257 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n11963) );
  AOI21_X1 U8258 ( .B1(n11991), .B2(n12384), .A(n11265), .ZN(n11267) );
  XNOR2_X1 U8259 ( .A(n11268), .B(n10663), .ZN(n9060) );
  INV_X1 U8260 ( .A(n7145), .ZN(n7144) );
  OAI21_X1 U8261 ( .B1(n9069), .B2(n7146), .A(n9073), .ZN(n7145) );
  INV_X1 U8262 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8738) );
  NAND2_X1 U8263 ( .A1(n11244), .A2(n11243), .ZN(n11983) );
  AOI21_X1 U8264 ( .B1(n11241), .B2(n14729), .A(n6634), .ZN(n6633) );
  NAND2_X1 U8265 ( .A1(n11925), .A2(n11264), .ZN(n11884) );
  AND2_X1 U8266 ( .A1(n11246), .A2(n7600), .ZN(n7180) );
  NOR2_X1 U8267 ( .A1(n7336), .A2(n12244), .ZN(n12246) );
  NOR2_X1 U8268 ( .A1(n12053), .A2(n7338), .ZN(n7337) );
  NAND2_X1 U8269 ( .A1(n12211), .A2(n12243), .ZN(n12247) );
  AND4_X1 U8270 ( .A1(n8744), .A2(n8743), .A3(n8742), .A4(n8741), .ZN(n12469)
         );
  NAND2_X1 U8271 ( .A1(n6909), .A2(n6908), .ZN(n7775) );
  NAND2_X1 U8272 ( .A1(n12659), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n6908) );
  OR2_X1 U8273 ( .A1(n12659), .A2(n14790), .ZN(n6909) );
  OAI21_X1 U8274 ( .B1(n9216), .B2(P3_REG1_REG_2__SCAN_IN), .A(n6934), .ZN(
        n9730) );
  NAND2_X1 U8275 ( .A1(n9216), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n6934) );
  OR2_X1 U8276 ( .A1(n7681), .A2(n9207), .ZN(n7682) );
  INV_X1 U8277 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7035) );
  OR2_X1 U8278 ( .A1(n9658), .A2(n14904), .ZN(n9771) );
  AOI21_X1 U8279 ( .B1(n9661), .B2(P3_REG1_REG_3__SCAN_IN), .A(n6546), .ZN(
        n9763) );
  NAND2_X1 U8280 ( .A1(n7086), .A2(n9923), .ZN(n9925) );
  INV_X1 U8281 ( .A(n7087), .ZN(n7086) );
  NAND2_X1 U8282 ( .A1(n7089), .A2(n9923), .ZN(n9783) );
  NOR2_X1 U8283 ( .A1(n9762), .A2(n6930), .ZN(n7746) );
  NOR2_X1 U8284 ( .A1(n9776), .A2(n14856), .ZN(n6930) );
  NAND2_X1 U8285 ( .A1(n7088), .A2(n9922), .ZN(n9927) );
  NOR2_X1 U8286 ( .A1(n9961), .A2(n10830), .ZN(n9960) );
  NAND2_X1 U8287 ( .A1(n7094), .A2(n7095), .ZN(n10031) );
  NAND2_X1 U8288 ( .A1(n10028), .A2(n7751), .ZN(n7752) );
  AOI21_X1 U8289 ( .B1(n14712), .B2(n14711), .A(n14710), .ZN(n14715) );
  NAND2_X1 U8290 ( .A1(n10683), .A2(n7755), .ZN(n10628) );
  NAND2_X1 U8291 ( .A1(n10628), .A2(n10629), .ZN(n10627) );
  NOR2_X1 U8292 ( .A1(n10678), .A2(n10677), .ZN(n10676) );
  OR2_X1 U8293 ( .A1(n10675), .A2(n11057), .ZN(n7101) );
  AND2_X1 U8294 ( .A1(n7098), .A2(n6480), .ZN(n7716) );
  NOR3_X1 U8295 ( .A1(n10925), .A2(n10924), .A3(n10923), .ZN(n11087) );
  OR3_X1 U8296 ( .A1(n11087), .A2(n11086), .A3(n11085), .ZN(n11088) );
  NAND2_X1 U8297 ( .A1(n11079), .A2(n7823), .ZN(n7759) );
  NAND2_X1 U8298 ( .A1(n14005), .A2(n14006), .ZN(n14004) );
  OAI21_X1 U8299 ( .B1(n14003), .B2(n13999), .A(n14000), .ZN(n14019) );
  AOI21_X1 U8300 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n9388), .A(n14010), .ZN(
        n7721) );
  NOR2_X1 U8301 ( .A1(n14023), .A2(n14931), .ZN(n14024) );
  AND2_X1 U8302 ( .A1(n12193), .A2(n12194), .ZN(n12321) );
  INV_X1 U8303 ( .A(n8871), .ZN(n8872) );
  NOR2_X1 U8304 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8872), .ZN(n8883) );
  OR2_X1 U8305 ( .A1(n8837), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8849) );
  AND2_X1 U8306 ( .A1(n8817), .A2(n11973), .ZN(n8828) );
  NOR2_X1 U8307 ( .A1(n8805), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U8308 ( .A1(n8791), .A2(n11963), .ZN(n8792) );
  NAND2_X1 U8309 ( .A1(n7555), .A2(n7554), .ZN(n12416) );
  AOI21_X1 U8310 ( .B1(n6468), .B2(n7560), .A(n7564), .ZN(n7554) );
  AND2_X1 U8311 ( .A1(n8767), .A2(n8766), .ZN(n8791) );
  NOR2_X1 U8312 ( .A1(n8720), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8739) );
  AND4_X1 U8313 ( .A1(n8698), .A2(n8697), .A3(n8696), .A4(n8695), .ZN(n11051)
         );
  OR2_X1 U8314 ( .A1(n8693), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8707) );
  AOI21_X1 U8315 ( .B1(n7582), .B2(n7583), .A(n7581), .ZN(n7580) );
  INV_X1 U8316 ( .A(n12119), .ZN(n7581) );
  INV_X1 U8317 ( .A(n8680), .ZN(n7582) );
  NAND2_X1 U8318 ( .A1(n8970), .A2(n12114), .ZN(n10933) );
  AND2_X1 U8319 ( .A1(n12114), .A2(n12113), .ZN(n12222) );
  AND4_X1 U8320 ( .A1(n8654), .A2(n8653), .A3(n8652), .A4(n8651), .ZN(n10781)
         );
  NAND2_X1 U8321 ( .A1(n6650), .A2(n12094), .ZN(n10774) );
  NAND2_X1 U8322 ( .A1(n10662), .A2(n12219), .ZN(n6650) );
  AND4_X1 U8323 ( .A1(n8624), .A2(n8623), .A3(n8622), .A4(n8621), .ZN(n10782)
         );
  NAND2_X1 U8324 ( .A1(n7548), .A2(n8605), .ZN(n10466) );
  NAND2_X1 U8325 ( .A1(n7036), .A2(n12080), .ZN(n10462) );
  NAND2_X1 U8326 ( .A1(n8968), .A2(n14757), .ZN(n7036) );
  AND2_X1 U8327 ( .A1(n12086), .A2(n12087), .ZN(n12221) );
  AND4_X1 U8328 ( .A1(n8888), .A2(n8887), .A3(n8886), .A4(n8885), .ZN(n12314)
         );
  AOI21_X1 U8329 ( .B1(n7570), .B2(n7574), .A(n6559), .ZN(n7568) );
  INV_X1 U8330 ( .A(n12380), .ZN(n12378) );
  NAND2_X1 U8331 ( .A1(n6654), .A2(n7046), .ZN(n12379) );
  AOI21_X1 U8332 ( .B1(n7048), .B2(n7056), .A(n7047), .ZN(n7046) );
  NAND2_X1 U8333 ( .A1(n12423), .A2(n7048), .ZN(n6654) );
  INV_X1 U8334 ( .A(n12165), .ZN(n7047) );
  AND2_X1 U8335 ( .A1(n8765), .A2(n8764), .ZN(n12154) );
  NAND2_X1 U8336 ( .A1(n11223), .A2(n8975), .ZN(n6642) );
  OR2_X1 U8337 ( .A1(n14843), .A2(n14833), .ZN(n14848) );
  NAND2_X1 U8338 ( .A1(n7189), .A2(n8947), .ZN(n9040) );
  AND2_X1 U8339 ( .A1(n6697), .A2(n6627), .ZN(n12025) );
  NAND2_X1 U8340 ( .A1(n8919), .A2(n8920), .ZN(n6697) );
  XNOR2_X1 U8341 ( .A(n7735), .B(P3_IR_REG_21__SCAN_IN), .ZN(n9041) );
  XNOR2_X1 U8342 ( .A(n8822), .B(n11449), .ZN(n8823) );
  NOR2_X1 U8343 ( .A1(n6884), .A2(n7646), .ZN(n6880) );
  OAI21_X1 U8344 ( .B1(n6679), .B2(n6678), .A(n6673), .ZN(n8774) );
  INV_X1 U8345 ( .A(n6674), .ZN(n6673) );
  OAI21_X1 U8346 ( .B1(n8569), .B2(n6677), .A(n6675), .ZN(n6674) );
  AOI21_X1 U8347 ( .B1(n6676), .B2(n8760), .A(n6607), .ZN(n6675) );
  OAI21_X1 U8348 ( .B1(n8560), .B2(n7333), .A(n6692), .ZN(n8728) );
  AND2_X1 U8349 ( .A1(n7330), .A2(n6693), .ZN(n6692) );
  NAND2_X1 U8350 ( .A1(n7332), .A2(n6694), .ZN(n6693) );
  AOI21_X1 U8351 ( .B1(n7332), .B2(n7334), .A(n6609), .ZN(n7330) );
  NOR2_X1 U8352 ( .A1(n7709), .A2(n7708), .ZN(n14685) );
  INV_X1 U8353 ( .A(n6680), .ZN(n8689) );
  AOI21_X1 U8354 ( .B1(n8666), .B2(n6684), .A(n6681), .ZN(n6680) );
  NAND2_X1 U8355 ( .A1(n6682), .A2(n8558), .ZN(n6681) );
  XNOR2_X1 U8356 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8688) );
  OR2_X1 U8357 ( .A1(n7693), .A2(P3_IR_REG_7__SCAN_IN), .ZN(n7699) );
  NAND2_X1 U8358 ( .A1(n6669), .A2(n8551), .ZN(n8642) );
  XNOR2_X1 U8359 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8640) );
  XNOR2_X1 U8360 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8625) );
  NAND2_X1 U8361 ( .A1(n7668), .A2(n7545), .ZN(n7679) );
  XNOR2_X1 U8362 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8612) );
  NAND2_X1 U8363 ( .A1(n8545), .A2(n8544), .ZN(n8600) );
  XNOR2_X1 U8364 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8579) );
  AND2_X1 U8365 ( .A1(n9338), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8586) );
  NOR2_X1 U8366 ( .A1(n9808), .A2(n9807), .ZN(n9865) );
  INV_X1 U8367 ( .A(n12667), .ZN(n7497) );
  INV_X1 U8368 ( .A(n11727), .ZN(n7496) );
  OR2_X1 U8369 ( .A1(n9981), .A2(n9980), .ZN(n10097) );
  XNOR2_X1 U8370 ( .A(n6459), .B(n11294), .ZN(n9369) );
  INV_X1 U8371 ( .A(n7019), .ZN(n7018) );
  OAI21_X1 U8372 ( .B1(n7021), .B2(n7020), .A(n12692), .ZN(n7019) );
  INV_X1 U8373 ( .A(n12723), .ZN(n7020) );
  NOR2_X1 U8374 ( .A1(n12722), .A2(n11701), .ZN(n7021) );
  OR2_X1 U8375 ( .A1(n11032), .A2(n11031), .ZN(n11182) );
  INV_X1 U8376 ( .A(n9620), .ZN(n6997) );
  INV_X1 U8377 ( .A(n9621), .ZN(n6998) );
  INV_X1 U8378 ( .A(n10093), .ZN(n7002) );
  OAI21_X1 U8379 ( .B1(n7007), .B2(n7001), .A(n10185), .ZN(n7000) );
  AND2_X1 U8380 ( .A1(n11437), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n11452) );
  XNOR2_X1 U8381 ( .A(n13167), .B(n11724), .ZN(n10949) );
  OR2_X1 U8382 ( .A1(n10425), .A2(n10424), .ZN(n10598) );
  OR2_X1 U8383 ( .A1(n10598), .A2(n10768), .ZN(n10764) );
  NOR2_X1 U8384 ( .A1(n11490), .A2(n12736), .ZN(n11503) );
  NAND2_X1 U8385 ( .A1(n11468), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11490) );
  NOR2_X1 U8386 ( .A1(n10479), .A2(n7507), .ZN(n7506) );
  INV_X1 U8387 ( .A(n10266), .ZN(n7507) );
  NAND2_X1 U8388 ( .A1(n9805), .A2(n9806), .ZN(n9858) );
  NOR2_X1 U8389 ( .A1(n10764), .A2(n10763), .ZN(n10954) );
  INV_X1 U8390 ( .A(n11683), .ZN(n7516) );
  NAND2_X1 U8391 ( .A1(n11597), .A2(n11596), .ZN(n6981) );
  NOR2_X1 U8392 ( .A1(n11606), .A2(n7278), .ZN(n11624) );
  NAND2_X1 U8393 ( .A1(n11635), .A2(n7279), .ZN(n7278) );
  NAND2_X1 U8394 ( .A1(n12766), .A2(n6446), .ZN(n7279) );
  NAND2_X1 U8395 ( .A1(n11635), .A2(n11574), .ZN(n11642) );
  AND2_X1 U8396 ( .A1(n9326), .A2(n9318), .ZN(n12754) );
  AND4_X1 U8397 ( .A1(n11523), .A2(n11522), .A3(n11521), .A4(n11520), .ZN(
        n12701) );
  NAND2_X1 U8398 ( .A1(n9355), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9315) );
  OR2_X1 U8399 ( .A1(n10001), .A2(n7366), .ZN(n6659) );
  AND2_X1 U8400 ( .A1(n10002), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7366) );
  NOR2_X1 U8401 ( .A1(n14466), .A2(n7363), .ZN(n9995) );
  AND2_X1 U8402 ( .A1(n14474), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7363) );
  NAND2_X1 U8403 ( .A1(n9995), .A2(n9994), .ZN(n10521) );
  NOR2_X1 U8404 ( .A1(n10705), .A2(n7361), .ZN(n10707) );
  AND2_X1 U8405 ( .A1(n10706), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7361) );
  NOR2_X1 U8406 ( .A1(n12784), .A2(n6605), .ZN(n12785) );
  OR2_X1 U8407 ( .A1(n14519), .A2(n14518), .ZN(n7354) );
  XNOR2_X1 U8408 ( .A(n12810), .B(n12809), .ZN(n12800) );
  NOR2_X1 U8409 ( .A1(n12800), .A2(n12799), .ZN(n12811) );
  NOR2_X1 U8410 ( .A1(n7079), .A2(n7076), .ZN(n7075) );
  NOR2_X1 U8411 ( .A1(n12889), .A2(n7432), .ZN(n7430) );
  OR2_X1 U8412 ( .A1(n7433), .A2(n12889), .ZN(n7428) );
  AND2_X1 U8413 ( .A1(n11556), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n12853) );
  OR2_X1 U8414 ( .A1(n13105), .A2(n12880), .ZN(n7208) );
  NAND2_X1 U8415 ( .A1(n6740), .A2(n12873), .ZN(n12983) );
  NAND2_X1 U8416 ( .A1(n6739), .A2(n6737), .ZN(n6740) );
  NOR2_X1 U8417 ( .A1(n12871), .A2(n6738), .ZN(n6737) );
  AND2_X1 U8418 ( .A1(n13131), .A2(n12839), .ZN(n7426) );
  NOR2_X1 U8419 ( .A1(n13021), .A2(n13131), .ZN(n13007) );
  NAND2_X1 U8420 ( .A1(n7073), .A2(n7072), .ZN(n13021) );
  NAND2_X1 U8421 ( .A1(n7441), .A2(n7439), .ZN(n13032) );
  INV_X1 U8422 ( .A(n7440), .ZN(n7439) );
  NOR2_X1 U8423 ( .A1(n7446), .A2(n7443), .ZN(n7442) );
  NOR2_X2 U8424 ( .A1(n13075), .A2(n13151), .ZN(n13074) );
  INV_X1 U8425 ( .A(n7080), .ZN(n11040) );
  OAI21_X1 U8426 ( .B1(n10749), .B2(n7211), .A(n7209), .ZN(n11044) );
  AOI21_X1 U8427 ( .B1(n7212), .B2(n7210), .A(n6535), .ZN(n7209) );
  INV_X1 U8428 ( .A(n7212), .ZN(n7211) );
  NAND2_X1 U8429 ( .A1(n7469), .A2(n6521), .ZN(n10985) );
  NAND2_X1 U8430 ( .A1(n10423), .A2(n6517), .ZN(n7469) );
  INV_X1 U8431 ( .A(n7471), .ZN(n7468) );
  NOR2_X1 U8432 ( .A1(n10097), .A2(n10096), .ZN(n10191) );
  AND2_X1 U8433 ( .A1(n10191), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10271) );
  OAI21_X1 U8434 ( .B1(n10255), .B2(n10232), .A(n7464), .ZN(n10320) );
  INV_X1 U8435 ( .A(n7465), .ZN(n7464) );
  OAI21_X1 U8436 ( .B1(n10255), .B2(n7462), .A(n7461), .ZN(n10418) );
  NAND2_X1 U8437 ( .A1(n10252), .A2(n10231), .ZN(n10233) );
  NAND2_X1 U8438 ( .A1(n10233), .A2(n10232), .ZN(n10313) );
  OR2_X1 U8439 ( .A1(n10258), .A2(n11356), .ZN(n10327) );
  NAND2_X1 U8440 ( .A1(n10287), .A2(n10261), .ZN(n10258) );
  NAND2_X1 U8441 ( .A1(n7421), .A2(n7420), .ZN(n10253) );
  AOI21_X1 U8442 ( .B1(n7422), .B2(n6515), .A(n6471), .ZN(n7420) );
  NAND2_X1 U8443 ( .A1(n10207), .A2(n7419), .ZN(n7421) );
  AND2_X1 U8444 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9633) );
  AND2_X1 U8445 ( .A1(n10205), .A2(n10140), .ZN(n11650) );
  NAND2_X1 U8446 ( .A1(n6717), .A2(n10120), .ZN(n10136) );
  NAND2_X1 U8447 ( .A1(n6715), .A2(n10044), .ZN(n10166) );
  INV_X1 U8448 ( .A(n12981), .ZN(n13121) );
  NAND2_X1 U8449 ( .A1(n7448), .A2(n7450), .ZN(n13067) );
  OR2_X1 U8450 ( .A1(n14543), .A2(n11685), .ZN(n14627) );
  INV_X1 U8451 ( .A(n14627), .ZN(n14637) );
  AND2_X1 U8452 ( .A1(n9575), .A2(n14641), .ZN(n14583) );
  AND4_X1 U8453 ( .A1(n9113), .A2(n9114), .A3(n9115), .A4(n9116), .ZN(n7597)
         );
  NOR2_X1 U8454 ( .A1(n7509), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n7508) );
  INV_X1 U8455 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9111) );
  AND2_X1 U8456 ( .A1(n9394), .A2(n9502), .ZN(n10882) );
  OR2_X1 U8457 ( .A1(n9228), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9264) );
  INV_X1 U8458 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n9192) );
  NOR2_X1 U8459 ( .A1(n9827), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n9193) );
  INV_X1 U8460 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9338) );
  INV_X1 U8461 ( .A(n13319), .ZN(n6742) );
  INV_X1 U8462 ( .A(n8390), .ZN(n8377) );
  NAND2_X1 U8463 ( .A1(n9902), .A2(n7246), .ZN(n7251) );
  OR2_X1 U8464 ( .A1(n9905), .A2(n9904), .ZN(n7250) );
  INV_X1 U8465 ( .A(n11815), .ZN(n11858) );
  INV_X1 U8466 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8048) );
  OR2_X1 U8467 ( .A1(n8099), .A2(n8082), .ZN(n8115) );
  INV_X1 U8468 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9532) );
  OR2_X1 U8469 ( .A1(n8313), .A2(n7961), .ZN(n8330) );
  NAND2_X1 U8470 ( .A1(n7226), .A2(n6493), .ZN(n11136) );
  INV_X1 U8471 ( .A(n13343), .ZN(n13964) );
  XNOR2_X1 U8472 ( .A(n9878), .B(n11856), .ZN(n9892) );
  OAI21_X1 U8473 ( .B1(n14351), .B2(n11824), .A(n7107), .ZN(n9878) );
  NAND2_X1 U8474 ( .A1(n8005), .A2(n9347), .ZN(n6821) );
  NAND2_X1 U8475 ( .A1(n13309), .A2(n13310), .ZN(n13243) );
  OR2_X1 U8476 ( .A1(n8216), .A2(n8215), .ZN(n8232) );
  NAND2_X1 U8477 ( .A1(n6939), .A2(n6940), .ZN(n8510) );
  NAND2_X1 U8478 ( .A1(n7952), .A2(n8271), .ZN(n6940) );
  OR2_X1 U8479 ( .A1(n8092), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8124) );
  NAND2_X1 U8480 ( .A1(n13739), .A2(n7034), .ZN(n7033) );
  NOR2_X1 U8481 ( .A1(n13750), .A2(n13745), .ZN(n7034) );
  NAND2_X1 U8482 ( .A1(n13589), .A2(n13535), .ZN(n13570) );
  NAND2_X1 U8483 ( .A1(n13591), .A2(n13590), .ZN(n13589) );
  NAND2_X2 U8484 ( .A1(n6937), .A2(n8415), .ZN(n13763) );
  NAND2_X1 U8485 ( .A1(n13772), .A2(n6879), .ZN(n6967) );
  INV_X1 U8486 ( .A(n13623), .ZN(n13628) );
  AOI21_X1 U8487 ( .B1(n7315), .B2(n13684), .A(n6537), .ZN(n7313) );
  NAND2_X1 U8488 ( .A1(n6946), .A2(n6824), .ZN(n13668) );
  INV_X1 U8489 ( .A(n7029), .ZN(n6946) );
  NAND2_X1 U8490 ( .A1(n6708), .A2(n6706), .ZN(n6711) );
  NOR2_X1 U8491 ( .A1(n13509), .A2(n6707), .ZN(n6706) );
  NOR2_X1 U8492 ( .A1(n6482), .A2(n13717), .ZN(n13715) );
  NOR2_X1 U8493 ( .A1(n8232), .A2(n8231), .ZN(n8241) );
  INV_X1 U8494 ( .A(n7384), .ZN(n10993) );
  AOI21_X1 U8495 ( .B1(n13976), .B2(n13975), .A(n6485), .ZN(n7384) );
  NOR2_X1 U8496 ( .A1(n8170), .A2(n9606), .ZN(n8190) );
  NAND2_X1 U8497 ( .A1(n7301), .A2(n6699), .ZN(n10817) );
  NAND2_X1 U8498 ( .A1(n8181), .A2(n8180), .ZN(n11131) );
  INV_X1 U8499 ( .A(n7376), .ZN(n7375) );
  NAND2_X1 U8500 ( .A1(n10514), .A2(n14152), .ZN(n10799) );
  INV_X1 U8501 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n14989) );
  OR2_X1 U8502 ( .A1(n8153), .A2(n14989), .ZN(n8170) );
  INV_X1 U8503 ( .A(n14412), .ZN(n10545) );
  OR2_X1 U8504 ( .A1(n8097), .A2(n8096), .ZN(n8099) );
  NAND2_X1 U8505 ( .A1(n10611), .A2(n14351), .ZN(n10610) );
  AOI211_X1 U8506 ( .C1(n13561), .C2(n6453), .A(n13541), .B(n14352), .ZN(
        n13741) );
  NOR2_X1 U8507 ( .A1(n6482), .A2(n7032), .ZN(n13686) );
  OAI21_X1 U8508 ( .B1(n10369), .B2(n7296), .A(n7294), .ZN(n10495) );
  AND2_X1 U8509 ( .A1(n10390), .A2(n9713), .ZN(n14397) );
  AND2_X1 U8510 ( .A1(n10571), .A2(n14400), .ZN(n14368) );
  XNOR2_X1 U8511 ( .A(n7290), .B(n7917), .ZN(n11567) );
  NAND2_X1 U8512 ( .A1(n8468), .A2(n7915), .ZN(n7290) );
  NAND2_X1 U8513 ( .A1(n7970), .A2(n7969), .ZN(n7913) );
  INV_X1 U8514 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7929) );
  XNOR2_X1 U8515 ( .A(n8447), .B(n8446), .ZN(n13204) );
  NAND2_X1 U8516 ( .A1(n7415), .A2(n7122), .ZN(n8524) );
  NOR2_X1 U8517 ( .A1(n7411), .A2(n8034), .ZN(n7415) );
  XNOR2_X1 U8518 ( .A(n8358), .B(n8357), .ZN(n11464) );
  XNOR2_X1 U8519 ( .A(n8352), .B(n8338), .ZN(n11448) );
  XNOR2_X1 U8520 ( .A(n8247), .B(n8246), .ZN(n11168) );
  XNOR2_X1 U8521 ( .A(n8220), .B(n8210), .ZN(n10942) );
  XNOR2_X1 U8522 ( .A(n8142), .B(n8141), .ZN(n10268) );
  NAND2_X1 U8523 ( .A1(n8123), .A2(n7866), .ZN(n8142) );
  NAND2_X1 U8524 ( .A1(n8090), .A2(n8089), .ZN(n8091) );
  OR2_X1 U8525 ( .A1(n8078), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8092) );
  NAND2_X1 U8526 ( .A1(n6733), .A2(n7850), .ZN(n8041) );
  CLKBUF_X1 U8527 ( .A(n8034), .Z(n8044) );
  INV_X1 U8528 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6789) );
  OAI21_X1 U8529 ( .B1(n13887), .B2(n13888), .A(n6553), .ZN(n7141) );
  XNOR2_X1 U8530 ( .A(n13842), .B(n13841), .ZN(n13894) );
  XNOR2_X1 U8531 ( .A(n13882), .B(n6932), .ZN(n13884) );
  INV_X1 U8532 ( .A(n6847), .ZN(n13902) );
  OAI21_X1 U8533 ( .B1(n15026), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n6532), .ZN(
        n6847) );
  NOR2_X1 U8534 ( .A1(n13847), .A2(n13846), .ZN(n13905) );
  NOR2_X1 U8535 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n13899), .ZN(n13846) );
  INV_X1 U8536 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n13903) );
  INV_X1 U8537 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14911) );
  NAND2_X1 U8538 ( .A1(n13910), .A2(n13911), .ZN(n13912) );
  NAND2_X1 U8539 ( .A1(n15030), .A2(n15031), .ZN(n13910) );
  OAI21_X1 U8540 ( .B1(n13858), .B2(n14723), .A(n13857), .ZN(n13876) );
  OAI21_X1 U8541 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14913), .A(n13861), .ZN(
        n13873) );
  OAI21_X1 U8542 ( .B1(n14176), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6511), .ZN(
        n6846) );
  OAI22_X1 U8543 ( .A1(n14182), .A2(n6849), .B1(n14181), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n13928) );
  NOR2_X1 U8544 ( .A1(n6905), .A2(n14500), .ZN(n6849) );
  AND4_X1 U8545 ( .A1(n8916), .A2(n8915), .A3(n8914), .A4(n8913), .ZN(n12316)
         );
  NAND2_X1 U8546 ( .A1(n7181), .A2(n11246), .ZN(n11897) );
  INV_X1 U8547 ( .A(n12362), .ZN(n11906) );
  XNOR2_X1 U8548 ( .A(n11267), .B(n11266), .ZN(n11903) );
  AND2_X1 U8549 ( .A1(n11069), .A2(n11068), .ZN(n11071) );
  AND3_X1 U8550 ( .A1(n8704), .A2(n8703), .A3(n8702), .ZN(n14725) );
  NAND2_X1 U8551 ( .A1(n9056), .A2(n9055), .ZN(n10074) );
  INV_X1 U8552 ( .A(n10073), .ZN(n9056) );
  AND2_X1 U8553 ( .A1(n7149), .A2(n14668), .ZN(n7148) );
  OAI21_X1 U8554 ( .B1(n11920), .B2(n6487), .A(n7150), .ZN(n7149) );
  NAND2_X1 U8555 ( .A1(n7152), .A2(n6487), .ZN(n7151) );
  INV_X1 U8556 ( .A(n11920), .ZN(n7152) );
  AND4_X1 U8557 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n11072)
         );
  NAND2_X1 U8558 ( .A1(n14669), .A2(n9069), .ZN(n10838) );
  NAND2_X1 U8559 ( .A1(n10838), .A2(n10837), .ZN(n10836) );
  NAND2_X1 U8560 ( .A1(n7171), .A2(n9050), .ZN(n9947) );
  INV_X1 U8561 ( .A(n7172), .ZN(n7171) );
  NAND2_X1 U8562 ( .A1(n11970), .A2(n11261), .ZN(n11927) );
  NAND2_X1 U8563 ( .A1(n6632), .A2(n11241), .ZN(n11935) );
  NAND2_X1 U8564 ( .A1(n11237), .A2(n11236), .ZN(n6632) );
  AOI21_X1 U8565 ( .B1(n11970), .B2(n6501), .A(n7175), .ZN(n11944) );
  NAND2_X1 U8566 ( .A1(n7178), .A2(n7176), .ZN(n7175) );
  NAND2_X1 U8567 ( .A1(n11883), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U8568 ( .A1(n7168), .A2(n7170), .ZN(n11954) );
  NAND2_X1 U8569 ( .A1(n7169), .A2(n6592), .ZN(n7168) );
  NAND2_X1 U8570 ( .A1(n7160), .A2(n7164), .ZN(n11962) );
  NAND2_X1 U8571 ( .A1(n7169), .A2(n7165), .ZN(n7160) );
  NAND2_X1 U8572 ( .A1(n6636), .A2(n7161), .ZN(n11960) );
  NAND2_X1 U8573 ( .A1(n12016), .A2(n7164), .ZN(n6636) );
  NAND2_X1 U8574 ( .A1(n6965), .A2(n6617), .ZN(n11273) );
  AND2_X1 U8575 ( .A1(n10074), .A2(n9059), .ZN(n10350) );
  NAND2_X1 U8576 ( .A1(n10074), .A2(n7174), .ZN(n10349) );
  INV_X1 U8577 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9098) );
  OR2_X1 U8578 ( .A1(n9097), .A2(n9096), .ZN(n14666) );
  XNOR2_X1 U8579 ( .A(n11238), .B(n11239), .ZN(n11237) );
  INV_X1 U8580 ( .A(n7161), .ZN(n6638) );
  AOI21_X1 U8581 ( .B1(n7163), .B2(n7161), .A(n6599), .ZN(n6637) );
  NAND2_X1 U8582 ( .A1(n9063), .A2(n9062), .ZN(n10725) );
  NAND2_X1 U8583 ( .A1(n10455), .A2(n10454), .ZN(n9063) );
  NAND2_X1 U8584 ( .A1(n8881), .A2(n8880), .ZN(n12500) );
  OR2_X1 U8585 ( .A1(n8601), .A2(n12662), .ZN(n8880) );
  NAND2_X1 U8586 ( .A1(n9944), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14678) );
  INV_X1 U8587 ( .A(n11051), .ZN(n12274) );
  INV_X1 U8588 ( .A(n11072), .ZN(n14732) );
  INV_X1 U8589 ( .A(n9071), .ZN(n12275) );
  INV_X1 U8590 ( .A(n10781), .ZN(n12276) );
  INV_X1 U8591 ( .A(n14761), .ZN(n10665) );
  NAND4_X1 U8592 ( .A1(n8585), .A2(n8584), .A3(n8583), .A4(n8582), .ZN(n12281)
         );
  OAI21_X1 U8593 ( .B1(n7672), .B2(n7106), .A(n7105), .ZN(n9727) );
  OR2_X1 U8594 ( .A1(n7671), .A2(n14774), .ZN(n7106) );
  OAI21_X1 U8595 ( .B1(n7672), .B2(n7671), .A(n14774), .ZN(n7105) );
  NAND2_X1 U8596 ( .A1(n9744), .A2(n7676), .ZN(n9726) );
  OAI22_X1 U8597 ( .A1(n9959), .A2(n7750), .B1(n8667), .B2(n7749), .ZN(n10030)
         );
  NAND2_X1 U8598 ( .A1(n7098), .A2(n7099), .ZN(n10624) );
  AND2_X1 U8599 ( .A1(n7101), .A2(n6483), .ZN(n10626) );
  XNOR2_X1 U8600 ( .A(n7716), .B(n8734), .ZN(n10917) );
  XNOR2_X1 U8601 ( .A(n7719), .B(n9259), .ZN(n12283) );
  XNOR2_X1 U8602 ( .A(n7759), .B(n12292), .ZN(n12285) );
  NOR2_X1 U8603 ( .A1(n12283), .A2(n12459), .ZN(n12282) );
  OAI21_X1 U8604 ( .B1(n12283), .B2(n7103), .A(n7102), .ZN(n14010) );
  NAND2_X1 U8605 ( .A1(n7104), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7103) );
  NAND2_X1 U8606 ( .A1(n7720), .A2(n7104), .ZN(n7102) );
  INV_X1 U8607 ( .A(n14009), .ZN(n7104) );
  INV_X1 U8608 ( .A(n7085), .ZN(n14043) );
  INV_X1 U8609 ( .A(n7773), .ZN(n7082) );
  NAND2_X1 U8610 ( .A1(n7085), .A2(n7084), .ZN(n7083) );
  NAND2_X1 U8611 ( .A1(n13951), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7084) );
  AND2_X1 U8612 ( .A1(n7764), .A2(n7738), .ZN(n14040) );
  XNOR2_X1 U8613 ( .A(n6928), .B(n7763), .ZN(n7771) );
  NAND2_X1 U8614 ( .A1(n14030), .A2(n6929), .ZN(n6928) );
  NAND2_X1 U8615 ( .A1(n13951), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6929) );
  OR2_X1 U8616 ( .A1(n8601), .A2(n12658), .ZN(n8894) );
  NAND2_X1 U8617 ( .A1(n8870), .A2(n8869), .ZN(n12343) );
  OR2_X1 U8618 ( .A1(n8601), .A2(n11097), .ZN(n8869) );
  AND2_X1 U8619 ( .A1(n7045), .A2(n6498), .ZN(n12351) );
  NAND2_X1 U8620 ( .A1(n12359), .A2(n12360), .ZN(n7045) );
  NAND2_X1 U8621 ( .A1(n8827), .A2(n8826), .ZN(n12388) );
  NAND2_X1 U8622 ( .A1(n10865), .A2(n7583), .ZN(n10934) );
  AND2_X1 U8623 ( .A1(n10865), .A2(n8681), .ZN(n10935) );
  NAND2_X1 U8624 ( .A1(n10779), .A2(n7587), .ZN(n14747) );
  NAND2_X1 U8625 ( .A1(n12253), .A2(n8966), .ZN(n14785) );
  NOR2_X1 U8626 ( .A1(n12055), .A2(n8994), .ZN(n14769) );
  AND2_X1 U8627 ( .A1(n8987), .A2(n14785), .ZN(n14793) );
  INV_X2 U8628 ( .A(n14793), .ZN(n14791) );
  OR2_X1 U8629 ( .A1(n8601), .A2(n12653), .ZN(n8909) );
  NAND2_X1 U8630 ( .A1(n8904), .A2(n8903), .ZN(n12301) );
  AOI21_X1 U8631 ( .B1(n12311), .B2(n12312), .A(n8980), .ZN(n12299) );
  INV_X1 U8632 ( .A(n12497), .ZN(n8902) );
  NAND2_X1 U8633 ( .A1(n7040), .A2(n7041), .ZN(n12333) );
  NAND2_X1 U8634 ( .A1(n12359), .A2(n7042), .ZN(n7040) );
  NAND2_X1 U8635 ( .A1(n7571), .A2(n7572), .ZN(n12370) );
  OR2_X1 U8636 ( .A1(n12405), .A2(n7574), .ZN(n7571) );
  INV_X1 U8637 ( .A(n12388), .ZN(n12583) );
  NAND2_X1 U8638 ( .A1(n7577), .A2(n7576), .ZN(n12381) );
  NAND2_X1 U8639 ( .A1(n12405), .A2(n7578), .ZN(n7576) );
  AOI21_X1 U8640 ( .B1(n12405), .B2(n8812), .A(n6461), .ZN(n12394) );
  NAND2_X1 U8641 ( .A1(n7050), .A2(n7053), .ZN(n12392) );
  NAND2_X1 U8642 ( .A1(n7052), .A2(n7051), .ZN(n7050) );
  NAND2_X1 U8643 ( .A1(n8804), .A2(n8803), .ZN(n12593) );
  NAND2_X1 U8644 ( .A1(n12525), .A2(n12063), .ZN(n12403) );
  NAND2_X1 U8645 ( .A1(n7557), .A2(n7558), .ZN(n12431) );
  OR2_X1 U8646 ( .A1(n12455), .A2(n7560), .ZN(n7557) );
  NAND2_X1 U8647 ( .A1(n12453), .A2(n7566), .ZN(n12444) );
  NAND2_X1 U8648 ( .A1(n8737), .A2(n8736), .ZN(n12634) );
  AND2_X1 U8649 ( .A1(n11219), .A2(n8732), .ZN(n12483) );
  NAND2_X1 U8650 ( .A1(n14851), .A2(n14821), .ZN(n12635) );
  NAND2_X1 U8651 ( .A1(n14851), .A2(n14848), .ZN(n12622) );
  AND2_X1 U8652 ( .A1(n8945), .A2(n8944), .ZN(n12637) );
  AND2_X1 U8653 ( .A1(n9081), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12636) );
  OR3_X1 U8654 ( .A1(n8535), .A2(n7646), .A3(n7070), .ZN(n7069) );
  AOI21_X1 U8655 ( .B1(n8535), .B2(n7070), .A(n6891), .ZN(n6890) );
  INV_X1 U8656 ( .A(n8537), .ZN(n12648) );
  NAND2_X1 U8657 ( .A1(n6435), .A2(n7058), .ZN(n7728) );
  INV_X1 U8658 ( .A(SI_26_), .ZN(n12662) );
  XNOR2_X1 U8659 ( .A(n6631), .B(n7059), .ZN(n12665) );
  NAND2_X1 U8660 ( .A1(n7726), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6631) );
  NAND2_X1 U8661 ( .A1(n7622), .A2(n7623), .ZN(n7726) );
  OAI21_X1 U8662 ( .B1(n6481), .B2(n7184), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7619) );
  NAND2_X1 U8663 ( .A1(n7185), .A2(n7628), .ZN(n7184) );
  NAND2_X1 U8664 ( .A1(n7342), .A2(n7343), .ZN(n8858) );
  NAND2_X1 U8665 ( .A1(n7346), .A2(n7348), .ZN(n8846) );
  NAND2_X1 U8666 ( .A1(n8833), .A2(n8834), .ZN(n7346) );
  NAND2_X1 U8667 ( .A1(n7186), .A2(n6499), .ZN(n7732) );
  INV_X1 U8668 ( .A(n9041), .ZN(n12069) );
  NAND2_X1 U8669 ( .A1(n8929), .A2(n6484), .ZN(n10112) );
  INV_X1 U8670 ( .A(SI_20_), .ZN(n10110) );
  NAND2_X1 U8671 ( .A1(n6687), .A2(n8783), .ZN(n8800) );
  NAND2_X1 U8672 ( .A1(n8781), .A2(n8782), .ZN(n6687) );
  AND2_X1 U8673 ( .A1(P3_U3151), .A2(n9154), .ZN(n13947) );
  INV_X1 U8674 ( .A(SI_16_), .ZN(n9387) );
  INV_X1 U8675 ( .A(SI_15_), .ZN(n9260) );
  NAND2_X1 U8676 ( .A1(n6679), .A2(n6671), .ZN(n8761) );
  INV_X1 U8677 ( .A(n6672), .ZN(n6671) );
  OAI21_X1 U8678 ( .B1(n8569), .B2(n7324), .A(n8571), .ZN(n6672) );
  NAND2_X1 U8679 ( .A1(n7323), .A2(n8569), .ZN(n8747) );
  NAND2_X1 U8680 ( .A1(n8733), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7323) );
  OR2_X1 U8681 ( .A1(n7648), .A2(n7647), .ZN(n11084) );
  INV_X1 U8682 ( .A(SI_12_), .ZN(n9198) );
  NAND2_X1 U8683 ( .A1(n7331), .A2(n8562), .ZN(n8714) );
  NAND2_X1 U8684 ( .A1(n8700), .A2(n8699), .ZN(n7331) );
  INV_X1 U8685 ( .A(SI_10_), .ZN(n9203) );
  NAND2_X1 U8686 ( .A1(n7665), .A2(n7664), .ZN(n14718) );
  INV_X1 U8687 ( .A(n14685), .ZN(n9178) );
  INV_X1 U8688 ( .A(n6683), .ZN(n8676) );
  AOI21_X1 U8689 ( .B1(n8666), .B2(n8665), .A(n6685), .ZN(n6683) );
  NAND2_X1 U8690 ( .A1(n7675), .A2(n7674), .ZN(n9752) );
  OR2_X1 U8691 ( .A1(n9296), .A2(n9038), .ZN(n9125) );
  OAI21_X1 U8692 ( .B1(n9970), .B2(n9971), .A(n9976), .ZN(n10084) );
  OR2_X1 U8693 ( .A1(n10945), .A2(n10946), .ZN(n10947) );
  NAND2_X1 U8694 ( .A1(n7013), .A2(n7499), .ZN(n10952) );
  NAND2_X1 U8695 ( .A1(n10267), .A2(n10266), .ZN(n10478) );
  AND2_X1 U8696 ( .A1(n7488), .A2(n6507), .ZN(n12684) );
  NAND2_X1 U8697 ( .A1(n7489), .A2(n7490), .ZN(n7488) );
  INV_X1 U8698 ( .A(n7493), .ZN(n7492) );
  OAI21_X1 U8699 ( .B1(n6486), .B2(n7495), .A(n7494), .ZN(n7493) );
  NAND2_X1 U8700 ( .A1(n11731), .A2(n7496), .ZN(n7494) );
  OR2_X1 U8701 ( .A1(n11731), .A2(n7496), .ZN(n7495) );
  NAND2_X1 U8702 ( .A1(n11551), .A2(n11584), .ZN(n11554) );
  NAND2_X1 U8703 ( .A1(n10094), .A2(n10093), .ZN(n10186) );
  NAND2_X1 U8704 ( .A1(n7003), .A2(n6615), .ZN(n10094) );
  XNOR2_X1 U8705 ( .A(n9370), .B(n9369), .ZN(n9343) );
  NAND2_X1 U8706 ( .A1(n9342), .A2(n9343), .ZN(n9373) );
  NAND2_X1 U8707 ( .A1(n7014), .A2(n7018), .ZN(n12691) );
  OR2_X1 U8708 ( .A1(n6952), .A2(n7020), .ZN(n7014) );
  NAND2_X1 U8709 ( .A1(n7017), .A2(n12723), .ZN(n12693) );
  NAND2_X1 U8710 ( .A1(n6952), .A2(n7021), .ZN(n7017) );
  NOR2_X1 U8711 ( .A1(n11691), .A2(n11690), .ZN(n12710) );
  NAND2_X1 U8712 ( .A1(n7476), .A2(n9619), .ZN(n9632) );
  INV_X1 U8713 ( .A(n11284), .ZN(n14545) );
  NAND2_X1 U8714 ( .A1(n6952), .A2(n11702), .ZN(n12726) );
  OAI21_X1 U8715 ( .B1(n10754), .B2(n10755), .A(n10756), .ZN(n10951) );
  OR2_X1 U8716 ( .A1(n9329), .A2(n11639), .ZN(n12744) );
  INV_X1 U8717 ( .A(n12744), .ZN(n12757) );
  NOR2_X1 U8718 ( .A1(n12708), .A2(n11695), .ZN(n12741) );
  NOR2_X1 U8719 ( .A1(n7478), .A2(n11720), .ZN(n7477) );
  INV_X1 U8720 ( .A(n7480), .ZN(n7478) );
  NAND2_X1 U8721 ( .A1(n9515), .A2(P2_STATE_REG_SCAN_IN), .ZN(n12742) );
  AND2_X1 U8722 ( .A1(n6767), .A2(n7513), .ZN(n6766) );
  NOR2_X1 U8723 ( .A1(n6477), .A2(n11687), .ZN(n7513) );
  NAND2_X1 U8724 ( .A1(n11628), .A2(n11633), .ZN(n6767) );
  NOR2_X1 U8725 ( .A1(n6534), .A2(n6765), .ZN(n6764) );
  INV_X1 U8726 ( .A(n11633), .ZN(n6765) );
  NAND2_X1 U8727 ( .A1(n7515), .A2(n11684), .ZN(n7514) );
  OAI21_X1 U8728 ( .B1(n13054), .B2(n11459), .A(n11188), .ZN(n12863) );
  NAND4_X1 U8729 ( .A1(n9322), .A2(n9321), .A3(n9320), .A4(n9319), .ZN(n12782)
         );
  NAND2_X1 U8730 ( .A1(n9355), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9321) );
  NAND2_X1 U8731 ( .A1(n9517), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9320) );
  AND2_X1 U8732 ( .A1(n9401), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7359) );
  INV_X1 U8733 ( .A(n7358), .ZN(n14443) );
  NOR2_X1 U8734 ( .A1(n14446), .A2(n6497), .ZN(n9399) );
  NOR2_X1 U8735 ( .A1(n9399), .A2(n9398), .ZN(n9488) );
  NOR2_X1 U8736 ( .A1(n9403), .A2(n9402), .ZN(n9492) );
  AND2_X1 U8737 ( .A1(n7358), .A2(n7357), .ZN(n9403) );
  NAND2_X1 U8738 ( .A1(n14451), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7357) );
  INV_X1 U8739 ( .A(n6641), .ZN(n14460) );
  NOR2_X1 U8740 ( .A1(n14458), .A2(n6594), .ZN(n9491) );
  NOR2_X1 U8741 ( .A1(n9681), .A2(n6911), .ZN(n9684) );
  AND2_X1 U8742 ( .A1(n9860), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6911) );
  NOR2_X1 U8743 ( .A1(n9684), .A2(n9683), .ZN(n10001) );
  AND2_X1 U8744 ( .A1(n10002), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7364) );
  AND2_X1 U8745 ( .A1(n6659), .A2(n6658), .ZN(n14469) );
  INV_X1 U8746 ( .A(n14470), .ZN(n6658) );
  INV_X1 U8747 ( .A(n6659), .ZN(n14471) );
  NOR2_X1 U8748 ( .A1(n14469), .A2(n7365), .ZN(n10006) );
  AND2_X1 U8749 ( .A1(n14474), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7365) );
  NOR2_X1 U8750 ( .A1(n14478), .A2(n7356), .ZN(n10522) );
  AND2_X1 U8751 ( .A1(n14486), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7356) );
  NAND2_X1 U8752 ( .A1(n10522), .A2(n10523), .ZN(n10701) );
  INV_X1 U8753 ( .A(n6656), .ZN(n10531) );
  NAND2_X1 U8754 ( .A1(n10701), .A2(n7355), .ZN(n10702) );
  OR2_X1 U8755 ( .A1(n10706), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7355) );
  NAND2_X1 U8756 ( .A1(n10702), .A2(n10703), .ZN(n10881) );
  XNOR2_X1 U8757 ( .A(n12785), .B(n12786), .ZN(n14491) );
  NOR2_X1 U8758 ( .A1(n12795), .A2(n6606), .ZN(n14494) );
  INV_X1 U8759 ( .A(n7354), .ZN(n14517) );
  NOR2_X1 U8760 ( .A1(n14502), .A2(n12798), .ZN(n14516) );
  INV_X1 U8761 ( .A(n7352), .ZN(n14514) );
  NOR2_X1 U8762 ( .A1(n14533), .A2(n14532), .ZN(n14530) );
  INV_X1 U8763 ( .A(n12814), .ZN(n14531) );
  NAND2_X1 U8764 ( .A1(n9130), .A2(n12822), .ZN(n14527) );
  NOR2_X1 U8765 ( .A1(n9134), .A2(P2_U3088), .ZN(n14442) );
  INV_X1 U8766 ( .A(n13096), .ZN(n12911) );
  OAI21_X1 U8767 ( .B1(n12917), .B2(n12926), .A(n6488), .ZN(n12903) );
  INV_X1 U8768 ( .A(n13100), .ZN(n12924) );
  AND2_X1 U8769 ( .A1(n6748), .A2(n6504), .ZN(n12939) );
  AND2_X2 U8770 ( .A1(n11516), .A2(n11515), .ZN(n13110) );
  INV_X1 U8771 ( .A(n6748), .ZN(n12948) );
  NAND2_X1 U8772 ( .A1(n6739), .A2(n7191), .ZN(n13000) );
  NAND2_X1 U8773 ( .A1(n7194), .A2(n7196), .ZN(n13013) );
  NAND2_X1 U8774 ( .A1(n7195), .A2(n12866), .ZN(n7194) );
  INV_X1 U8775 ( .A(n13041), .ZN(n7195) );
  NAND2_X1 U8776 ( .A1(n13041), .A2(n12865), .ZN(n13027) );
  NAND2_X1 U8777 ( .A1(n7200), .A2(n7204), .ZN(n13059) );
  NAND2_X1 U8778 ( .A1(n12859), .A2(n7201), .ZN(n7200) );
  OAI21_X1 U8779 ( .B1(n11023), .B2(n7438), .A(n7437), .ZN(n13048) );
  INV_X1 U8780 ( .A(n7447), .ZN(n7438) );
  NAND2_X1 U8781 ( .A1(n7206), .A2(n7201), .ZN(n13065) );
  NAND2_X1 U8782 ( .A1(n7206), .A2(n12857), .ZN(n13063) );
  NAND2_X1 U8783 ( .A1(n7453), .A2(n7460), .ZN(n12834) );
  OR2_X1 U8784 ( .A1(n11023), .A2(n11022), .ZN(n7453) );
  NAND2_X1 U8785 ( .A1(n10980), .A2(n10979), .ZN(n11008) );
  NAND2_X1 U8786 ( .A1(n10735), .A2(n7472), .ZN(n10737) );
  NAND2_X1 U8787 ( .A1(n10422), .A2(n10421), .ZN(n11374) );
  NAND2_X1 U8788 ( .A1(n10241), .A2(n7463), .ZN(n10318) );
  NAND2_X1 U8789 ( .A1(n10230), .A2(n10229), .ZN(n10250) );
  NAND2_X1 U8790 ( .A1(n10236), .A2(n10235), .ZN(n10283) );
  NAND2_X1 U8791 ( .A1(n9862), .A2(n9861), .ZN(n14601) );
  NAND2_X1 U8792 ( .A1(n14554), .A2(n10056), .ZN(n13076) );
  OR2_X1 U8793 ( .A1(n9511), .A2(n9348), .ZN(n9351) );
  OR2_X1 U8794 ( .A1(n10758), .A2(n9349), .ZN(n9350) );
  NAND2_X1 U8795 ( .A1(n14566), .A2(n9306), .ZN(n13071) );
  AND2_X1 U8796 ( .A1(n14554), .A2(n12819), .ZN(n13078) );
  INV_X2 U8797 ( .A(n14661), .ZN(n14663) );
  INV_X2 U8798 ( .A(n14646), .ZN(n14648) );
  AND2_X1 U8799 ( .A1(n9304), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14566) );
  NAND2_X1 U8800 ( .A1(n7216), .A2(n9311), .ZN(n13201) );
  MUX2_X1 U8801 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9310), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n9311) );
  XNOR2_X1 U8802 ( .A(n9028), .B(P2_IR_REG_26__SCAN_IN), .ZN(n13207) );
  AND2_X1 U8803 ( .A1(n9031), .A2(n9032), .ZN(n11118) );
  INV_X1 U8804 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11500) );
  INV_X1 U8805 ( .A(n7893), .ZN(n8371) );
  INV_X1 U8806 ( .A(n9330), .ZN(n11672) );
  NAND2_X1 U8807 ( .A1(n6992), .A2(n6991), .ZN(n9291) );
  NAND2_X1 U8808 ( .A1(n7510), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6991) );
  INV_X1 U8809 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9834) );
  AND2_X1 U8810 ( .A1(n9833), .A2(n10068), .ZN(n14536) );
  INV_X1 U8811 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n11025) );
  INV_X1 U8812 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9395) );
  INV_X1 U8813 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9267) );
  INV_X1 U8814 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9183) );
  OAI21_X1 U8815 ( .B1(n6596), .B2(n10691), .A(n7238), .ZN(n10850) );
  NAND2_X1 U8816 ( .A1(n7244), .A2(n11742), .ZN(n13225) );
  AND4_X1 U8817 ( .A1(n8120), .A2(n8119), .A3(n8118), .A4(n8117), .ZN(n10974)
         );
  NAND2_X1 U8818 ( .A1(n13243), .A2(n11784), .ZN(n13247) );
  AOI21_X1 U8819 ( .B1(n7241), .B2(n11847), .A(n11855), .ZN(n7240) );
  NAND2_X1 U8820 ( .A1(n7228), .A2(n7232), .ZN(n10851) );
  NAND2_X1 U8821 ( .A1(n6596), .A2(n7234), .ZN(n7228) );
  XNOR2_X1 U8822 ( .A(n9892), .B(n9891), .ZN(n9885) );
  INV_X1 U8823 ( .A(n9880), .ZN(n9881) );
  INV_X1 U8824 ( .A(n14351), .ZN(n10619) );
  NAND2_X1 U8825 ( .A1(n7243), .A2(n11794), .ZN(n13255) );
  NAND2_X1 U8826 ( .A1(n11136), .A2(n11135), .ZN(n11199) );
  OAI21_X1 U8827 ( .B1(n13236), .B2(n7225), .A(n7223), .ZN(n13263) );
  NAND2_X1 U8828 ( .A1(n13331), .A2(n13330), .ZN(n7227) );
  NOR2_X1 U8829 ( .A1(n10339), .A2(n10303), .ZN(n10552) );
  NAND2_X1 U8830 ( .A1(n13285), .A2(n13286), .ZN(n13284) );
  NAND2_X1 U8831 ( .A1(n13236), .A2(n11822), .ZN(n13285) );
  NAND2_X1 U8832 ( .A1(n7229), .A2(n7231), .ZN(n6754) );
  AOI21_X1 U8833 ( .B1(n11784), .B2(n6735), .A(n6554), .ZN(n6734) );
  INV_X1 U8834 ( .A(n11784), .ZN(n6736) );
  INV_X1 U8835 ( .A(n13310), .ZN(n6735) );
  INV_X1 U8836 ( .A(n6745), .ZN(n6744) );
  OAI21_X1 U8837 ( .B1(n6493), .B2(n6746), .A(n11198), .ZN(n6745) );
  NAND2_X1 U8838 ( .A1(n13253), .A2(n13300), .ZN(n6718) );
  NOR2_X1 U8839 ( .A1(n13334), .A2(n13963), .ZN(n14073) );
  OR2_X1 U8840 ( .A1(n9837), .A2(n9848), .ZN(n13334) );
  XNOR2_X1 U8841 ( .A(n11754), .B(n11755), .ZN(n13331) );
  NAND2_X1 U8842 ( .A1(n8230), .A2(n8229), .ZN(n13337) );
  AND2_X1 U8843 ( .A1(n9854), .A2(n14397), .ZN(n14075) );
  INV_X1 U8844 ( .A(n13528), .ZN(n13256) );
  OR2_X2 U8845 ( .A1(n9908), .A2(n9244), .ZN(n15020) );
  OR2_X1 U8846 ( .A1(n13824), .A2(n6455), .ZN(n8473) );
  INV_X1 U8847 ( .A(n13538), .ZN(n13539) );
  NAND2_X1 U8848 ( .A1(n13558), .A2(n6522), .ZN(n6712) );
  AND2_X1 U8849 ( .A1(n7308), .A2(n7307), .ZN(n13560) );
  NAND2_X1 U8850 ( .A1(n7388), .A2(n7387), .ZN(n7386) );
  NAND2_X1 U8851 ( .A1(n13557), .A2(n6454), .ZN(n7388) );
  NAND2_X1 U8852 ( .A1(n13586), .A2(n7309), .ZN(n13575) );
  AND2_X1 U8853 ( .A1(n13518), .A2(n13627), .ZN(n13604) );
  AND2_X1 U8854 ( .A1(n13603), .A2(n13518), .ZN(n7318) );
  NAND2_X1 U8855 ( .A1(n7396), .A2(n7397), .ZN(n13639) );
  AND2_X1 U8856 ( .A1(n7396), .A2(n7394), .ZN(n13637) );
  NAND2_X1 U8857 ( .A1(n7398), .A2(n13666), .ZN(n7396) );
  AND2_X1 U8858 ( .A1(n7400), .A2(n7403), .ZN(n13652) );
  NAND2_X1 U8859 ( .A1(n13666), .A2(n13667), .ZN(n7400) );
  NAND2_X1 U8860 ( .A1(n13681), .A2(n13512), .ZN(n13665) );
  NAND2_X1 U8861 ( .A1(n7408), .A2(n7410), .ZN(n13694) );
  AND2_X1 U8862 ( .A1(n7408), .A2(n7406), .ZN(n13693) );
  OR2_X1 U8863 ( .A1(n6489), .A2(n13526), .ZN(n7408) );
  NAND2_X1 U8864 ( .A1(n11432), .A2(n8460), .ZN(n8294) );
  NAND2_X1 U8865 ( .A1(n6708), .A2(n13506), .ZN(n13706) );
  AND2_X1 U8866 ( .A1(n8269), .A2(n8268), .ZN(n13522) );
  NAND2_X1 U8867 ( .A1(n11157), .A2(n11156), .ZN(n13505) );
  AND2_X1 U8868 ( .A1(n10820), .A2(n10819), .ZN(n7311) );
  AND2_X1 U8869 ( .A1(n14313), .A2(n9843), .ZN(n13725) );
  INV_X1 U8870 ( .A(n7027), .ZN(n10813) );
  NAND2_X1 U8871 ( .A1(n7312), .A2(n10819), .ZN(n10821) );
  NAND2_X1 U8872 ( .A1(n10509), .A2(n10508), .ZN(n10791) );
  NAND2_X1 U8873 ( .A1(n7302), .A2(n10513), .ZN(n10795) );
  NAND2_X1 U8874 ( .A1(n10512), .A2(n10511), .ZN(n7302) );
  INV_X1 U8875 ( .A(n14313), .ZN(n13720) );
  OAI21_X1 U8876 ( .B1(n14290), .B2(n7300), .A(n6467), .ZN(n6703) );
  OR2_X1 U8877 ( .A1(n14322), .A2(n14094), .ZN(n14298) );
  NAND2_X1 U8878 ( .A1(n7298), .A2(n10374), .ZN(n10398) );
  NAND2_X1 U8879 ( .A1(n14290), .A2(n14291), .ZN(n7298) );
  NAND2_X1 U8880 ( .A1(n10369), .A2(n10368), .ZN(n10646) );
  NAND2_X1 U8881 ( .A1(n10576), .A2(n10366), .ZN(n14308) );
  NOR2_X1 U8882 ( .A1(n14322), .A2(n14379), .ZN(n13977) );
  OR2_X1 U8883 ( .A1(n9837), .A2(n9569), .ZN(n14438) );
  AND2_X2 U8884 ( .A1(n9651), .A2(n9650), .ZN(n14425) );
  XNOR2_X1 U8885 ( .A(n8529), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9239) );
  OAI21_X1 U8886 ( .B1(n8528), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8529) );
  INV_X1 U8887 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6713) );
  NAND2_X1 U8888 ( .A1(n6496), .A2(n7951), .ZN(n7317) );
  NAND2_X1 U8889 ( .A1(n7951), .A2(n7934), .ZN(n7939) );
  INV_X1 U8890 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n11276) );
  NAND2_X1 U8891 ( .A1(n8528), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U8892 ( .A1(n7252), .A2(n7254), .ZN(n8516) );
  INV_X1 U8893 ( .A(n7947), .ZN(n7252) );
  OAI211_X1 U8894 ( .C1(n7951), .C2(n6807), .A(n7947), .B(n6806), .ZN(n10114)
         );
  NAND2_X1 U8895 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n6807) );
  NAND2_X1 U8896 ( .A1(n7931), .A2(n13816), .ZN(n6806) );
  INV_X1 U8897 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9793) );
  INV_X1 U8898 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9900) );
  AND2_X1 U8899 ( .A1(n8204), .A2(n8211), .ZN(n14190) );
  OR2_X1 U8900 ( .A1(n6989), .A2(n8121), .ZN(n8122) );
  INV_X1 U8901 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n9219) );
  INV_X1 U8902 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9191) );
  OAI21_X1 U8903 ( .B1(n8089), .B2(n8090), .A(n8091), .ZN(n9977) );
  INV_X1 U8904 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9186) );
  NAND2_X1 U8905 ( .A1(n7374), .A2(n7373), .ZN(n7372) );
  INV_X1 U8906 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n7837) );
  NAND2_X1 U8907 ( .A1(n9154), .A2(P1_U3086), .ZN(n13833) );
  XNOR2_X1 U8908 ( .A(n13890), .B(n6985), .ZN(n15036) );
  AOI21_X1 U8909 ( .B1(n14965), .B2(n13893), .A(n13940), .ZN(n15034) );
  XNOR2_X1 U8910 ( .A(n13900), .B(n13901), .ZN(n15026) );
  XNOR2_X1 U8911 ( .A(n13902), .B(n7138), .ZN(n13945) );
  INV_X1 U8912 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7138) );
  XNOR2_X1 U8913 ( .A(n13908), .B(n13909), .ZN(n15030) );
  XNOR2_X1 U8914 ( .A(n13912), .B(n13913), .ZN(n13946) );
  NAND2_X1 U8915 ( .A1(n6837), .A2(n6836), .ZN(n14174) );
  NAND2_X1 U8916 ( .A1(n6839), .A2(n6840), .ZN(n6836) );
  OAI21_X1 U8917 ( .B1(n13918), .B2(n6841), .A(n14489), .ZN(n6840) );
  XNOR2_X1 U8918 ( .A(n13923), .B(n13924), .ZN(n14176) );
  INV_X1 U8919 ( .A(n6846), .ZN(n14179) );
  NOR2_X1 U8920 ( .A1(n13928), .A2(n13927), .ZN(n14184) );
  AND2_X1 U8921 ( .A1(n13928), .A2(n13927), .ZN(n14185) );
  OAI22_X1 U8922 ( .A1(n9014), .A2(n12540), .B1(n9013), .B2(n12548), .ZN(n9001) );
  NAND2_X1 U8923 ( .A1(n7479), .A2(n7480), .ZN(n12706) );
  AOI21_X1 U8924 ( .B1(n6662), .B2(n12819), .A(n6661), .ZN(n6660) );
  OAI21_X1 U8925 ( .B1(n7368), .B2(n6664), .A(n11680), .ZN(n6663) );
  INV_X1 U8926 ( .A(n7367), .ZN(n6661) );
  NAND2_X1 U8927 ( .A1(n6944), .A2(n7218), .ZN(n6943) );
  INV_X1 U8928 ( .A(n6903), .ZN(n6902) );
  OAI21_X1 U8929 ( .B1(n13582), .B2(n13329), .A(n13222), .ZN(n6903) );
  NAND2_X1 U8930 ( .A1(n8486), .A2(n6514), .ZN(n6852) );
  OR2_X1 U8931 ( .A1(n6798), .A2(n6797), .ZN(n6796) );
  INV_X1 U8932 ( .A(n6799), .ZN(n6795) );
  NAND2_X1 U8933 ( .A1(n7142), .A2(n13918), .ZN(n13954) );
  INV_X1 U8934 ( .A(n14182), .ZN(n6848) );
  INV_X1 U8935 ( .A(n7135), .ZN(n14187) );
  NOR2_X1 U8936 ( .A1(n6834), .A2(n14188), .ZN(n13983) );
  NAND2_X1 U8937 ( .A1(n6829), .A2(n6832), .ZN(n13982) );
  OR2_X1 U8938 ( .A1(n13986), .A2(n13987), .ZN(n6947) );
  NOR2_X1 U8939 ( .A1(n13988), .A2(n13987), .ZN(n13997) );
  AND2_X1 U8940 ( .A1(n7041), .A2(n12242), .ZN(n6460) );
  NAND2_X1 U8941 ( .A1(n6565), .A2(n11251), .ZN(n7164) );
  NAND4_X1 U8942 ( .A1(n9317), .A2(n9316), .A3(n9315), .A4(n9314), .ZN(n11289)
         );
  AND2_X1 U8943 ( .A1(n12411), .A2(n12270), .ZN(n6461) );
  AND2_X1 U8944 ( .A1(n7623), .A2(n7059), .ZN(n6462) );
  NAND2_X1 U8945 ( .A1(n10082), .A2(n10081), .ZN(n6463) );
  INV_X1 U8946 ( .A(n11348), .ZN(n6917) );
  INV_X1 U8947 ( .A(n6481), .ZN(n7186) );
  AND3_X2 U8948 ( .A1(n8038), .A2(n8037), .A3(n8036), .ZN(n14367) );
  NAND2_X1 U8949 ( .A1(n9576), .A2(n10058), .ZN(n7418) );
  OR2_X1 U8950 ( .A1(n13842), .A2(n13841), .ZN(n6464) );
  NAND2_X1 U8951 ( .A1(n11569), .A2(n11568), .ZN(n11605) );
  INV_X1 U8952 ( .A(n8508), .ZN(n6887) );
  INV_X1 U8953 ( .A(n12862), .ZN(n13058) );
  AND2_X1 U8954 ( .A1(n13661), .A2(n13530), .ZN(n6465) );
  AND2_X1 U8955 ( .A1(n11405), .A2(n11404), .ZN(n6466) );
  AND2_X1 U8956 ( .A1(n10397), .A2(n7299), .ZN(n6467) );
  INV_X2 U8957 ( .A(n11824), .ZN(n9889) );
  AND2_X1 U8958 ( .A1(n7556), .A2(n7558), .ZN(n6468) );
  AND3_X1 U8959 ( .A1(n6954), .A2(n6574), .A3(n6887), .ZN(n6469) );
  NAND2_X1 U8960 ( .A1(n12634), .A2(n12469), .ZN(n6470) );
  AND2_X1 U8961 ( .A1(n11347), .A2(n10238), .ZN(n6471) );
  AND2_X1 U8962 ( .A1(n12276), .A2(n14820), .ZN(n6472) );
  INV_X1 U8963 ( .A(n11525), .ZN(n7525) );
  AND3_X1 U8964 ( .A1(n7122), .A2(n7121), .A3(n7940), .ZN(n6473) );
  AND2_X1 U8965 ( .A1(n13131), .A2(n12869), .ZN(n6474) );
  OR2_X1 U8966 ( .A1(n11415), .A2(n11414), .ZN(n6475) );
  INV_X1 U8967 ( .A(n7043), .ZN(n7042) );
  NAND2_X1 U8968 ( .A1(n12184), .A2(n12360), .ZN(n7043) );
  XNOR2_X1 U8969 ( .A(n7946), .B(P1_IR_REG_20__SCAN_IN), .ZN(n10389) );
  AND2_X1 U8970 ( .A1(n6456), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6476) );
  NAND2_X1 U8971 ( .A1(n11637), .A2(n7516), .ZN(n6477) );
  INV_X1 U8972 ( .A(n7164), .ZN(n7163) );
  OR2_X1 U8973 ( .A1(n12593), .A2(n12270), .ZN(n12217) );
  OR2_X1 U8974 ( .A1(n13984), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n6478) );
  AND2_X1 U8975 ( .A1(n12924), .A2(n12881), .ZN(n6479) );
  AND2_X1 U8976 ( .A1(n7099), .A2(n6620), .ZN(n6480) );
  INV_X1 U8977 ( .A(n9239), .ZN(n9233) );
  AND2_X1 U8978 ( .A1(n11147), .A2(n8492), .ZN(n11145) );
  INV_X1 U8979 ( .A(n11145), .ZN(n6901) );
  INV_X1 U8980 ( .A(n13300), .ZN(n6721) );
  INV_X1 U8981 ( .A(n7028), .ZN(n13685) );
  NOR2_X1 U8982 ( .A1(n6482), .A2(n7029), .ZN(n7028) );
  INV_X1 U8983 ( .A(n10858), .ZN(n6822) );
  NAND2_X1 U8984 ( .A1(n7659), .A2(n7658), .ZN(n10633) );
  INV_X1 U8985 ( .A(n14029), .ZN(n13951) );
  INV_X1 U8986 ( .A(n9339), .ZN(n11713) );
  NAND3_X1 U8987 ( .A1(n7649), .A2(n7613), .A3(n7588), .ZN(n6481) );
  INV_X1 U8988 ( .A(n8606), .ZN(n8851) );
  INV_X1 U8989 ( .A(n8243), .ZN(n8317) );
  NAND2_X1 U8990 ( .A1(n8895), .A2(n8894), .ZN(n12497) );
  OR2_X1 U8991 ( .A1(n14124), .A2(n14116), .ZN(n6482) );
  INV_X1 U8992 ( .A(n8719), .ZN(n8821) );
  INV_X1 U8993 ( .A(n8012), .ZN(n8334) );
  NAND2_X1 U8994 ( .A1(n8294), .A2(n8293), .ZN(n13700) );
  NAND2_X1 U8995 ( .A1(n8166), .A2(n8165), .ZN(n11100) );
  OR2_X1 U8996 ( .A1(n7714), .A2(n10682), .ZN(n6483) );
  AND2_X1 U8997 ( .A1(n6759), .A2(n7508), .ZN(n9110) );
  OR2_X1 U8998 ( .A1(n6481), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n6484) );
  INV_X1 U8999 ( .A(n13984), .ZN(n6833) );
  INV_X1 U9000 ( .A(n7079), .ZN(n13086) );
  NAND2_X1 U9001 ( .A1(n11610), .A2(n11609), .ZN(n7079) );
  NOR2_X1 U9002 ( .A1(n14145), .A2(n11200), .ZN(n6485) );
  AND2_X1 U9003 ( .A1(n7497), .A2(n7498), .ZN(n6486) );
  INV_X1 U9004 ( .A(n13772), .ZN(n13631) );
  AND2_X2 U9005 ( .A1(n8398), .A2(n8397), .ZN(n13772) );
  NAND2_X1 U9006 ( .A1(n8910), .A2(n8909), .ZN(n12552) );
  AND2_X1 U9007 ( .A1(n7154), .A2(n7153), .ZN(n6487) );
  OR2_X1 U9008 ( .A1(n12924), .A2(n12882), .ZN(n6488) );
  NAND2_X1 U9009 ( .A1(n6723), .A2(n13235), .ZN(n13236) );
  NAND2_X1 U9010 ( .A1(n6779), .A2(n6777), .ZN(n11284) );
  INV_X1 U9011 ( .A(n11273), .ZN(n12569) );
  INV_X1 U9012 ( .A(n11654), .ZN(n6743) );
  AND2_X2 U9013 ( .A1(n13524), .A2(n13523), .ZN(n6489) );
  XOR2_X1 U9014 ( .A(n12981), .B(n11729), .Z(n6490) );
  XNOR2_X1 U9015 ( .A(n9112), .B(n9111), .ZN(n9294) );
  AND2_X1 U9016 ( .A1(n6718), .A2(n13301), .ZN(n6491) );
  INV_X1 U9017 ( .A(n7321), .ZN(n10613) );
  NAND2_X1 U9018 ( .A1(n9703), .A2(n9705), .ZN(n7321) );
  XNOR2_X1 U9019 ( .A(n13151), .B(n12860), .ZN(n13066) );
  AND2_X1 U9020 ( .A1(n7179), .A2(n11261), .ZN(n6492) );
  OR2_X1 U9021 ( .A1(n7690), .A2(n7689), .ZN(n9788) );
  NAND2_X1 U9022 ( .A1(n8574), .A2(n8573), .ZN(n12616) );
  AND2_X1 U9023 ( .A1(n11109), .A2(n11107), .ZN(n6493) );
  INV_X1 U9024 ( .A(n7500), .ZN(n7499) );
  OAI21_X1 U9025 ( .B1(n10950), .B2(n7502), .A(n7501), .ZN(n7500) );
  AND2_X1 U9026 ( .A1(n11445), .A2(n11444), .ZN(n6494) );
  INV_X1 U9027 ( .A(n7265), .ZN(n7264) );
  NAND2_X1 U9028 ( .A1(n7267), .A2(n6540), .ZN(n7265) );
  OR2_X1 U9029 ( .A1(n13844), .A2(n13843), .ZN(n6495) );
  AND2_X1 U9030 ( .A1(n7934), .A2(n7935), .ZN(n6496) );
  XNOR2_X1 U9031 ( .A(n7949), .B(n7948), .ZN(n11869) );
  NAND2_X1 U9032 ( .A1(n13586), .A2(n7306), .ZN(n7308) );
  AND2_X1 U9033 ( .A1(n14451), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6497) );
  OR2_X1 U9034 ( .A1(n12572), .A2(n12178), .ZN(n6498) );
  AND2_X1 U9035 ( .A1(n7618), .A2(n7187), .ZN(n6499) );
  NOR2_X1 U9036 ( .A1(n12203), .A2(n12206), .ZN(n12241) );
  INV_X1 U9037 ( .A(n13136), .ZN(n7072) );
  INV_X1 U9038 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14986) );
  AOI21_X1 U9039 ( .B1(n7067), .B2(n8980), .A(n7066), .ZN(n7065) );
  INV_X1 U9040 ( .A(n7065), .ZN(n7064) );
  INV_X2 U9041 ( .A(n7847), .ZN(n9299) );
  AND2_X1 U9042 ( .A1(n9623), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6500) );
  AND2_X1 U9043 ( .A1(n11883), .A2(n6492), .ZN(n6501) );
  OR2_X1 U9044 ( .A1(n7072), .A2(n12867), .ZN(n6502) );
  XNOR2_X1 U9045 ( .A(n13088), .B(n11643), .ZN(n12886) );
  INV_X1 U9046 ( .A(n12886), .ZN(n6976) );
  OR2_X1 U9047 ( .A1(n7205), .A2(n12832), .ZN(n6503) );
  NAND2_X1 U9048 ( .A1(n12879), .A2(n12878), .ZN(n6504) );
  OR2_X1 U9049 ( .A1(n6481), .A2(n7183), .ZN(n6505) );
  INV_X1 U9050 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9159) );
  AND2_X1 U9051 ( .A1(n13167), .A2(n12771), .ZN(n6506) );
  NAND2_X1 U9052 ( .A1(n11698), .A2(n11697), .ZN(n6507) );
  OR2_X1 U9053 ( .A1(n13913), .A2(n13912), .ZN(n6508) );
  AND2_X1 U9054 ( .A1(n11920), .A2(n7155), .ZN(n6509) );
  AND2_X1 U9055 ( .A1(n13839), .A2(n9247), .ZN(n13661) );
  INV_X1 U9056 ( .A(n13661), .ZN(n13786) );
  AND3_X1 U9057 ( .A1(n12201), .A2(n12200), .A3(n12199), .ZN(n6510) );
  INV_X1 U9058 ( .A(n12709), .ZN(n7486) );
  OR2_X1 U9059 ( .A1(n13923), .A2(n13924), .ZN(n6511) );
  INV_X1 U9060 ( .A(n13745), .ZN(n6825) );
  AND2_X1 U9061 ( .A1(n11705), .A2(n11707), .ZN(n6512) );
  AND2_X1 U9062 ( .A1(n11461), .A2(n11460), .ZN(n6513) );
  AND2_X1 U9063 ( .A1(n8487), .A2(n8520), .ZN(n6514) );
  INV_X1 U9064 ( .A(n6455), .ZN(n8414) );
  AND2_X1 U9065 ( .A1(n10237), .A2(n7423), .ZN(n6515) );
  INV_X1 U9066 ( .A(n10374), .ZN(n7300) );
  OR2_X1 U9067 ( .A1(n12970), .A2(n12876), .ZN(n6516) );
  AND2_X1 U9068 ( .A1(n7471), .A2(n10440), .ZN(n6517) );
  AND2_X1 U9069 ( .A1(n13780), .A2(n13517), .ZN(n6518) );
  OR2_X1 U9070 ( .A1(n9247), .A2(n7985), .ZN(n6519) );
  OR2_X1 U9071 ( .A1(n7797), .A2(n7692), .ZN(n6520) );
  OR2_X1 U9072 ( .A1(n7470), .A2(n7468), .ZN(n6521) );
  OR2_X1 U9073 ( .A1(n6825), .A2(n13521), .ZN(n6522) );
  INV_X1 U9074 ( .A(n6751), .ZN(n12978) );
  NOR2_X1 U9075 ( .A1(n12993), .A2(n13121), .ZN(n6751) );
  NOR2_X1 U9076 ( .A1(n12391), .A2(n7049), .ZN(n7048) );
  OR2_X1 U9077 ( .A1(n13534), .A2(n13519), .ZN(n6523) );
  AND2_X1 U9078 ( .A1(n6901), .A2(n10999), .ZN(n6524) );
  AND2_X1 U9079 ( .A1(n11801), .A2(n11794), .ZN(n6525) );
  NOR2_X1 U9080 ( .A1(n12282), .A2(n7720), .ZN(n6526) );
  NOR2_X1 U9081 ( .A1(n7132), .A2(n7134), .ZN(n6527) );
  INV_X1 U9082 ( .A(n12866), .ZN(n7199) );
  INV_X1 U9083 ( .A(n7473), .ZN(n7472) );
  INV_X1 U9084 ( .A(n7504), .ZN(n7503) );
  OR2_X1 U9085 ( .A1(n10950), .A2(n7505), .ZN(n7504) );
  AND2_X1 U9086 ( .A1(n6743), .A2(n10229), .ZN(n6528) );
  AND2_X1 U9087 ( .A1(n11749), .A2(n11742), .ZN(n6529) );
  AND2_X1 U9088 ( .A1(n7433), .A2(n7429), .ZN(n6530) );
  INV_X1 U9089 ( .A(n7310), .ZN(n7309) );
  AND2_X1 U9090 ( .A1(n8978), .A2(n12184), .ZN(n12350) );
  INV_X1 U9091 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n9337) );
  INV_X1 U9092 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7628) );
  AND2_X1 U9093 ( .A1(n13559), .A2(n7307), .ZN(n6531) );
  OR2_X1 U9094 ( .A1(n13901), .A2(n13900), .ZN(n6532) );
  NAND2_X1 U9095 ( .A1(n7119), .A2(n7118), .ZN(n6533) );
  NAND2_X1 U9096 ( .A1(n11675), .A2(n11684), .ZN(n6534) );
  NOR2_X1 U9097 ( .A1(n13167), .A2(n12771), .ZN(n6535) );
  AND2_X1 U9098 ( .A1(n7040), .A2(n6460), .ZN(n6536) );
  AND2_X1 U9099 ( .A1(n12097), .A2(n12101), .ZN(n12218) );
  NOR2_X1 U9100 ( .A1(n13529), .A2(n13678), .ZN(n6537) );
  INV_X1 U9101 ( .A(n7457), .ZN(n7445) );
  NAND2_X1 U9102 ( .A1(n7458), .A2(n12860), .ZN(n7457) );
  AND2_X1 U9103 ( .A1(n9060), .A2(n10782), .ZN(n6538) );
  AND4_X1 U9104 ( .A1(n7621), .A2(n7620), .A3(n7188), .A4(n7628), .ZN(n6539)
         );
  OR2_X1 U9105 ( .A1(n7883), .A2(SI_17_), .ZN(n6540) );
  OR2_X1 U9106 ( .A1(n8386), .A2(n8388), .ZN(n6541) );
  NOR2_X1 U9107 ( .A1(n8510), .A2(n8509), .ZN(n6542) );
  NAND3_X1 U9108 ( .A1(n7122), .A2(n7413), .A3(n7255), .ZN(n6543) );
  AND2_X1 U9109 ( .A1(n12343), .A2(n12189), .ZN(n6544) );
  AND2_X1 U9110 ( .A1(n9894), .A2(n9895), .ZN(n6545) );
  AND2_X1 U9111 ( .A1(n7745), .A2(n9207), .ZN(n6546) );
  AND2_X1 U9112 ( .A1(n11346), .A2(n11345), .ZN(n6547) );
  NOR2_X1 U9113 ( .A1(n12388), .A2(n12268), .ZN(n6548) );
  NAND2_X1 U9114 ( .A1(n9027), .A2(n7510), .ZN(n7509) );
  AND2_X1 U9115 ( .A1(n7397), .A2(n7395), .ZN(n7394) );
  AND2_X1 U9116 ( .A1(n11324), .A2(n11323), .ZN(n6549) );
  INV_X1 U9117 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7023) );
  AND2_X1 U9118 ( .A1(n7882), .A2(n9387), .ZN(n6550) );
  OR2_X1 U9119 ( .A1(n11379), .A2(n11378), .ZN(n6551) );
  AND2_X1 U9120 ( .A1(n10034), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6552) );
  INV_X1 U9121 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7614) );
  INV_X1 U9122 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n7070) );
  NAND2_X1 U9123 ( .A1(n13357), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n6553) );
  INV_X1 U9124 ( .A(n7584), .ZN(n7583) );
  NAND2_X1 U9125 ( .A1(n12227), .A2(n8681), .ZN(n7584) );
  AND2_X1 U9126 ( .A1(n11788), .A2(n11787), .ZN(n6554) );
  AND2_X1 U9127 ( .A1(n7867), .A2(n9203), .ZN(n6555) );
  OR2_X1 U9128 ( .A1(n11377), .A2(n7533), .ZN(n6556) );
  NOR3_X1 U9129 ( .A1(n8277), .A2(n8276), .A3(n8285), .ZN(n6557) );
  NOR2_X1 U9130 ( .A1(n12588), .A2(n12383), .ZN(n6558) );
  NOR2_X1 U9131 ( .A1(n8844), .A2(n12384), .ZN(n6559) );
  AND2_X1 U9132 ( .A1(n9013), .A2(n12262), .ZN(n12203) );
  NAND2_X1 U9133 ( .A1(n10368), .A2(n10652), .ZN(n6560) );
  AND2_X1 U9134 ( .A1(n10299), .A2(n10298), .ZN(n6561) );
  NAND2_X1 U9135 ( .A1(n11352), .A2(n11353), .ZN(n6562) );
  NAND2_X1 U9136 ( .A1(n8745), .A2(n8732), .ZN(n6563) );
  INV_X1 U9137 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7510) );
  AND2_X1 U9138 ( .A1(n13531), .A2(n7403), .ZN(n6564) );
  INV_X1 U9139 ( .A(n6839), .ZN(n6838) );
  NAND2_X1 U9140 ( .A1(n13918), .A2(n6841), .ZN(n6839) );
  OR2_X1 U9141 ( .A1(n11252), .A2(n7167), .ZN(n6565) );
  AND2_X1 U9142 ( .A1(n7830), .A2(n14029), .ZN(n6566) );
  INV_X1 U9143 ( .A(n13953), .ZN(n6841) );
  OR2_X1 U9144 ( .A1(n12578), .A2(n12363), .ZN(n6567) );
  OR2_X1 U9145 ( .A1(n12583), .A2(n12396), .ZN(n6568) );
  AND2_X1 U9146 ( .A1(n6486), .A2(n11731), .ZN(n6569) );
  OR2_X1 U9147 ( .A1(n11429), .A2(n11431), .ZN(n6570) );
  OR2_X1 U9148 ( .A1(n11391), .A2(n6598), .ZN(n6571) );
  OR2_X1 U9149 ( .A1(n12998), .A2(n12872), .ZN(n6572) );
  NOR2_X1 U9150 ( .A1(n11100), .A2(n13344), .ZN(n6573) );
  XOR2_X1 U9151 ( .A(n13736), .B(n13543), .Z(n6574) );
  NOR2_X1 U9152 ( .A1(n13741), .A2(n13740), .ZN(n6575) );
  AND2_X1 U9153 ( .A1(n6542), .A2(n8520), .ZN(n6576) );
  AND2_X1 U9154 ( .A1(n12300), .A2(n7339), .ZN(n6577) );
  AND2_X1 U9155 ( .A1(n9126), .A2(n9337), .ZN(n6578) );
  NAND2_X1 U9156 ( .A1(n13146), .A2(n12863), .ZN(n6579) );
  NAND2_X1 U9157 ( .A1(n13100), .A2(n12882), .ZN(n6580) );
  AND2_X1 U9158 ( .A1(n6462), .A2(n7730), .ZN(n6581) );
  NAND2_X1 U9159 ( .A1(n11022), .A2(n7460), .ZN(n6582) );
  OR2_X1 U9160 ( .A1(n7544), .A2(n11430), .ZN(n6583) );
  AND2_X1 U9161 ( .A1(n7254), .A2(n7253), .ZN(n6584) );
  AND2_X1 U9162 ( .A1(n13934), .A2(n13933), .ZN(n14188) );
  NAND2_X1 U9163 ( .A1(n11400), .A2(n11401), .ZN(n6585) );
  AND2_X1 U9164 ( .A1(n7838), .A2(n9173), .ZN(n6586) );
  AND2_X1 U9165 ( .A1(n10371), .A2(n7293), .ZN(n6587) );
  INV_X1 U9166 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9117) );
  AND2_X1 U9167 ( .A1(n12740), .A2(n11694), .ZN(n7490) );
  INV_X1 U9168 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9121) );
  INV_X1 U9169 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n6884) );
  NAND4_X1 U9170 ( .A1(n11642), .A2(n11627), .A3(n11626), .A4(n11625), .ZN(
        n6588) );
  AND2_X1 U9171 ( .A1(n6848), .A2(n6905), .ZN(n6589) );
  OR2_X1 U9172 ( .A1(n11463), .A2(n6513), .ZN(n6590) );
  INV_X1 U9173 ( .A(n6463), .ZN(n7006) );
  INV_X1 U9174 ( .A(n10399), .ZN(n7297) );
  INV_X1 U9175 ( .A(n7159), .ZN(n7158) );
  NAND2_X1 U9176 ( .A1(n11887), .A2(n12314), .ZN(n7159) );
  INV_X1 U9177 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n7931) );
  INV_X1 U9178 ( .A(n8362), .ZN(n6802) );
  MUX2_X1 U9179 ( .A(n13533), .B(n13763), .S(n8479), .Z(n8417) );
  INV_X1 U9180 ( .A(n8417), .ZN(n6813) );
  INV_X1 U9181 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n7374) );
  INV_X1 U9182 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n7255) );
  INV_X1 U9183 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7188) );
  AND2_X1 U9184 ( .A1(n7613), .A2(n7649), .ZN(n7644) );
  INV_X1 U9185 ( .A(n13607), .ZN(n6879) );
  NAND2_X1 U9186 ( .A1(n14729), .A2(n11212), .ZN(n6591) );
  NAND2_X1 U9187 ( .A1(n12014), .A2(n12468), .ZN(n6592) );
  AND2_X1 U9188 ( .A1(n6470), .A2(n12232), .ZN(n6593) );
  INV_X1 U9189 ( .A(n8420), .ZN(n8298) );
  OAI21_X1 U9190 ( .B1(n6596), .B2(n7231), .A(n7229), .ZN(n10899) );
  AND2_X1 U9191 ( .A1(n14463), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6594) );
  XNOR2_X1 U9192 ( .A(n8523), .B(P1_IR_REG_24__SCAN_IN), .ZN(n9234) );
  OAI21_X1 U9193 ( .B1(n7226), .B2(n6746), .A(n6744), .ZN(n11739) );
  NAND2_X1 U9194 ( .A1(n11155), .A2(n11154), .ZN(n14098) );
  XOR2_X1 U9195 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .Z(n6595) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7326) );
  INV_X1 U9197 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n7059) );
  AND2_X1 U9198 ( .A1(n6758), .A2(n6757), .ZN(n6596) );
  INV_X1 U9199 ( .A(n14729), .ZN(n11236) );
  XNOR2_X1 U9200 ( .A(n7683), .B(P3_IR_REG_4__SCAN_IN), .ZN(n9776) );
  INV_X1 U9201 ( .A(n13234), .ZN(n6720) );
  NAND2_X1 U9202 ( .A1(n7227), .A2(n11757), .ZN(n14070) );
  AND3_X1 U9203 ( .A1(n14567), .A2(n11647), .A3(n7417), .ZN(n6597) );
  AND2_X1 U9204 ( .A1(n10779), .A2(n8648), .ZN(n14746) );
  INV_X1 U9205 ( .A(n8665), .ZN(n6686) );
  XNOR2_X1 U9206 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8665) );
  AND2_X1 U9207 ( .A1(n11388), .A2(n11387), .ZN(n6598) );
  AND2_X1 U9208 ( .A1(n11253), .A2(n12271), .ZN(n6599) );
  AND2_X1 U9209 ( .A1(n7012), .A2(n7013), .ZN(n6600) );
  INV_X1 U9210 ( .A(n8746), .ZN(n7324) );
  INV_X1 U9211 ( .A(n7073), .ZN(n13036) );
  AND2_X1 U9212 ( .A1(n14139), .A2(n10999), .ZN(n6601) );
  NOR2_X1 U9213 ( .A1(n11969), .A2(n12419), .ZN(n7564) );
  AND2_X1 U9214 ( .A1(n10735), .A2(n7470), .ZN(n6602) );
  AND2_X1 U9215 ( .A1(n8223), .A2(SI_14_), .ZN(n6603) );
  NAND2_X1 U9216 ( .A1(n11981), .A2(n12469), .ZN(n6604) );
  INV_X1 U9217 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6941) );
  INV_X1 U9218 ( .A(n7056), .ZN(n7051) );
  OR2_X1 U9219 ( .A1(n12216), .A2(n7057), .ZN(n7056) );
  INV_X1 U9220 ( .A(n7566), .ZN(n7563) );
  NAND2_X1 U9221 ( .A1(n12616), .A2(n7567), .ZN(n7566) );
  AND2_X1 U9222 ( .A1(n12796), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n6605) );
  AND2_X1 U9223 ( .A1(n12796), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6606) );
  AND2_X1 U9224 ( .A1(n12593), .A2(n12270), .ZN(n12216) );
  INV_X1 U9225 ( .A(n12216), .ZN(n7055) );
  INV_X1 U9226 ( .A(n7333), .ZN(n7332) );
  OAI21_X1 U9227 ( .B1(n8699), .B2(n7334), .A(n8713), .ZN(n7333) );
  INV_X1 U9228 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10759) );
  AND2_X1 U9229 ( .A1(n9900), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6607) );
  AND2_X1 U9230 ( .A1(n7883), .A2(SI_17_), .ZN(n6608) );
  AND2_X1 U9231 ( .A1(n8563), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6609) );
  AND2_X1 U9232 ( .A1(n7591), .A2(n7606), .ZN(n6610) );
  INV_X1 U9233 ( .A(n7166), .ZN(n7165) );
  NAND2_X1 U9234 ( .A1(n11251), .A2(n6592), .ZN(n7166) );
  NAND2_X1 U9235 ( .A1(n9291), .A2(n9290), .ZN(n11671) );
  INV_X1 U9236 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6919) );
  AND2_X1 U9237 ( .A1(n14546), .A2(n9294), .ZN(n14630) );
  INV_X1 U9238 ( .A(n8760), .ZN(n6678) );
  AND2_X1 U9239 ( .A1(n7081), .A2(n11010), .ZN(n6611) );
  INV_X1 U9240 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11465) );
  OR2_X1 U9241 ( .A1(n8425), .A2(n12662), .ZN(n6612) );
  NAND2_X1 U9242 ( .A1(n6703), .A2(n10399), .ZN(n10447) );
  INV_X1 U9243 ( .A(n14136), .ZN(n7026) );
  INV_X1 U9244 ( .A(n10756), .ZN(n7505) );
  INV_X1 U9245 ( .A(n13151), .ZN(n7458) );
  NAND2_X1 U9246 ( .A1(n7226), .A2(n11107), .ZN(n11108) );
  INV_X1 U9247 ( .A(n6455), .ZN(n8460) );
  NAND2_X1 U9248 ( .A1(n12836), .A2(n12857), .ZN(n7205) );
  INV_X1 U9249 ( .A(n7205), .ZN(n7201) );
  INV_X1 U9250 ( .A(n7081), .ZN(n10981) );
  NOR2_X1 U9251 ( .A1(n9960), .A2(n7698), .ZN(n6613) );
  AND2_X1 U9252 ( .A1(n7250), .A2(n7249), .ZN(n6614) );
  OR2_X1 U9253 ( .A1(n7007), .A2(n7006), .ZN(n6615) );
  AND2_X1 U9254 ( .A1(n7343), .A2(n6695), .ZN(n6616) );
  OR2_X1 U9255 ( .A1(n8601), .A2(n11281), .ZN(n6617) );
  AND2_X1 U9256 ( .A1(n10409), .A2(n10408), .ZN(n6618) );
  OR2_X1 U9257 ( .A1(n8845), .A2(n7345), .ZN(n6619) );
  NAND2_X1 U9258 ( .A1(n10633), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6620) );
  AND2_X1 U9259 ( .A1(n8444), .A2(SI_27_), .ZN(n6621) );
  INV_X1 U9260 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10070) );
  INV_X1 U9261 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n11169) );
  INV_X1 U9262 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10113) );
  AND2_X1 U9263 ( .A1(n6838), .A2(n7142), .ZN(n6622) );
  INV_X1 U9264 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6922) );
  INV_X1 U9265 ( .A(n12749), .ZN(n12763) );
  INV_X1 U9266 ( .A(n14376), .ZN(n7025) );
  INV_X1 U9267 ( .A(n11680), .ZN(n12819) );
  OR2_X1 U9268 ( .A1(n12043), .A2(n12650), .ZN(n6623) );
  INV_X1 U9269 ( .A(n8106), .ZN(n8399) );
  OR2_X1 U9270 ( .A1(n10611), .A2(n9840), .ZN(n6624) );
  NAND2_X1 U9271 ( .A1(n10042), .A2(n11284), .ZN(n10163) );
  INV_X1 U9272 ( .A(n10163), .ZN(n6749) );
  INV_X1 U9273 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n13834) );
  AND2_X1 U9274 ( .A1(n9050), .A2(n9046), .ZN(n6625) );
  INV_X1 U9275 ( .A(SI_22_), .ZN(n6953) );
  AND2_X1 U9276 ( .A1(n9299), .A2(P2_U3088), .ZN(n6626) );
  NAND2_X1 U9277 ( .A1(n13830), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6627) );
  INV_X1 U9278 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6985) );
  INV_X1 U9279 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7275) );
  INV_X1 U9280 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6987) );
  INV_X1 U9281 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7329) );
  INV_X1 U9282 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n6932) );
  AND3_X2 U9283 ( .A1(n7545), .A2(n7668), .A3(n6628), .ZN(n7649) );
  NAND2_X4 U9284 ( .A1(n9043), .A2(n6629), .ZN(n11268) );
  NAND3_X1 U9285 ( .A1(n7189), .A2(n9039), .A3(n8947), .ZN(n6629) );
  AND2_X1 U9286 ( .A1(n10351), .A2(n9059), .ZN(n7174) );
  OAI21_X2 U9287 ( .B1(n12016), .B2(n6638), .A(n6637), .ZN(n11999) );
  NAND2_X1 U9288 ( .A1(n11999), .A2(n11998), .ZN(n11997) );
  NAND2_X1 U9289 ( .A1(n9045), .A2(n14796), .ZN(n6644) );
  NAND2_X1 U9290 ( .A1(n6644), .A2(n12077), .ZN(n9945) );
  NAND2_X1 U9291 ( .A1(n6644), .A2(n12072), .ZN(n12073) );
  OAI21_X1 U9292 ( .B1(n6646), .B2(n12076), .A(n6645), .ZN(n12078) );
  NAND3_X1 U9293 ( .A1(n10662), .A2(n12218), .A3(n12219), .ZN(n6649) );
  NOR2_X1 U9294 ( .A1(n14530), .A2(n6652), .ZN(n12810) );
  OAI21_X2 U9295 ( .B1(n12379), .B2(n12170), .A(n12164), .ZN(n12369) );
  OR2_X2 U9296 ( .A1(n14481), .A2(n7362), .ZN(n6656) );
  NAND3_X1 U9297 ( .A1(n6435), .A2(n7058), .A3(n6657), .ZN(n8533) );
  NAND2_X1 U9298 ( .A1(n6663), .A2(n6660), .ZN(P2_U3233) );
  OAI22_X1 U9299 ( .A1(n12817), .A2(n14531), .B1(n14527), .B2(n12818), .ZN(
        n6662) );
  NAND2_X1 U9300 ( .A1(n6665), .A2(n12815), .ZN(n6664) );
  NAND2_X1 U9301 ( .A1(n8627), .A2(n8625), .ZN(n6669) );
  NAND2_X1 U9302 ( .A1(n8614), .A2(n8612), .ZN(n8549) );
  NAND2_X1 U9303 ( .A1(n8600), .A2(n8598), .ZN(n6670) );
  NAND2_X1 U9304 ( .A1(n8733), .A2(n7322), .ZN(n6679) );
  NAND2_X1 U9305 ( .A1(n10817), .A2(n10816), .ZN(n6698) );
  NAND2_X1 U9306 ( .A1(n10512), .A2(n7303), .ZN(n6699) );
  OAI21_X1 U9307 ( .B1(n14290), .B2(n6704), .A(n10448), .ZN(n6701) );
  NAND2_X1 U9308 ( .A1(n6702), .A2(n6700), .ZN(n6705) );
  INV_X1 U9309 ( .A(n6701), .ZN(n6700) );
  OR2_X1 U9310 ( .A1(n6467), .A2(n7297), .ZN(n6702) );
  NAND2_X1 U9311 ( .A1(n6705), .A2(n10400), .ZN(n10540) );
  NAND2_X1 U9312 ( .A1(n13702), .A2(n13701), .ZN(n13511) );
  INV_X1 U9313 ( .A(n13823), .ZN(n7960) );
  NAND2_X1 U9314 ( .A1(n7994), .A2(n7842), .ZN(n6714) );
  OAI21_X2 U9315 ( .B1(n7982), .B2(n7981), .A(n6856), .ZN(n7994) );
  NAND2_X1 U9316 ( .A1(n7840), .A2(SI_0_), .ZN(n7981) );
  NAND2_X1 U9317 ( .A1(n11645), .A2(n7418), .ZN(n6715) );
  OR2_X1 U9318 ( .A1(n7418), .A2(n9577), .ZN(n10059) );
  NAND2_X1 U9319 ( .A1(n10136), .A2(n10135), .ZN(n6716) );
  NAND2_X1 U9320 ( .A1(n10116), .A2(n10117), .ZN(n6717) );
  NAND3_X1 U9321 ( .A1(n11757), .A2(n6726), .A3(n6724), .ZN(n13272) );
  INV_X1 U9322 ( .A(n6725), .ZN(n6724) );
  NAND2_X1 U9323 ( .A1(n13272), .A2(n13273), .ZN(n11774) );
  OAI21_X2 U9324 ( .B1(n6733), .B2(n8042), .A(n6730), .ZN(n8068) );
  NAND2_X1 U9325 ( .A1(n8033), .A2(n7849), .ZN(n6733) );
  OAI21_X1 U9326 ( .B1(n13262), .B2(n6742), .A(n6741), .ZN(n13218) );
  NAND2_X1 U9327 ( .A1(n13318), .A2(n13319), .ZN(n13317) );
  INV_X2 U9328 ( .A(n11294), .ZN(n10042) );
  NAND2_X2 U9329 ( .A1(n6950), .A2(n9303), .ZN(n11294) );
  AND2_X2 U9330 ( .A1(n7081), .A2(n6750), .ZN(n7080) );
  NOR2_X2 U9331 ( .A1(n12951), .A2(n13105), .ZN(n7602) );
  NOR2_X2 U9332 ( .A1(n12978), .A2(n13116), .ZN(n12968) );
  NAND2_X1 U9333 ( .A1(n7857), .A2(n7856), .ZN(n8090) );
  AND2_X2 U9334 ( .A1(n10289), .A2(n14610), .ZN(n10287) );
  NAND3_X1 U9335 ( .A1(n6755), .A2(n10898), .A3(n6754), .ZN(n10967) );
  NAND3_X1 U9336 ( .A1(n6758), .A2(n7229), .A3(n6757), .ZN(n6755) );
  NAND2_X1 U9337 ( .A1(n7232), .A2(n7230), .ZN(n6756) );
  INV_X1 U9338 ( .A(n10551), .ZN(n6758) );
  NAND2_X1 U9339 ( .A1(n6759), .A2(n7597), .ZN(n9120) );
  AND4_X4 U9340 ( .A1(n9825), .A2(n7474), .A3(n9824), .A4(n9162), .ZN(n6759)
         );
  NAND2_X1 U9341 ( .A1(n6759), .A2(n9027), .ZN(n9287) );
  NAND2_X1 U9342 ( .A1(n6759), .A2(n7475), .ZN(n7071) );
  NAND3_X1 U9343 ( .A1(n6759), .A2(n7475), .A3(n9117), .ZN(n9308) );
  NAND3_X1 U9344 ( .A1(n6759), .A2(n7475), .A3(n7214), .ZN(n7216) );
  NAND3_X1 U9345 ( .A1(n9022), .A2(n9159), .A3(n6760), .ZN(n9829) );
  MUX2_X1 U9346 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9828), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n9833) );
  NAND3_X1 U9347 ( .A1(n6763), .A2(n6761), .A3(n6768), .ZN(P2_U3328) );
  NAND2_X1 U9348 ( .A1(n6762), .A2(n6766), .ZN(n6761) );
  NAND2_X1 U9349 ( .A1(n7287), .A2(n11633), .ZN(n6762) );
  OAI21_X1 U9350 ( .B1(n7287), .B2(n11628), .A(n6764), .ZN(n6763) );
  AND2_X1 U9351 ( .A1(n7514), .A2(n11688), .ZN(n6768) );
  NAND2_X1 U9352 ( .A1(n6562), .A2(n6771), .ZN(n6770) );
  NAND2_X1 U9353 ( .A1(n11322), .A2(n11321), .ZN(n6775) );
  NAND2_X1 U9354 ( .A1(n9154), .A2(SI_0_), .ZN(n6778) );
  NAND2_X2 U9355 ( .A1(n13206), .A2(n9126), .ZN(n11026) );
  NAND2_X1 U9356 ( .A1(n13206), .A2(n6578), .ZN(n6779) );
  NAND2_X1 U9357 ( .A1(n11026), .A2(n13215), .ZN(n6777) );
  XNOR2_X1 U9358 ( .A(n6778), .B(n9338), .ZN(n13215) );
  NAND2_X1 U9359 ( .A1(n11415), .A2(n11414), .ZN(n6893) );
  NAND2_X1 U9360 ( .A1(n6784), .A2(n7534), .ZN(n11480) );
  OAI22_X2 U9361 ( .A1(n7512), .A2(n6785), .B1(n11497), .B2(n11496), .ZN(
        n11510) );
  INV_X1 U9362 ( .A(n11510), .ZN(n11508) );
  NAND3_X1 U9363 ( .A1(n6789), .A2(n7373), .A3(n7374), .ZN(n8006) );
  OAI21_X2 U9364 ( .B1(n8477), .B2(n10389), .A(n6790), .ZN(n8106) );
  INV_X1 U9365 ( .A(n8106), .ZN(n8017) );
  INV_X1 U9366 ( .A(n8452), .ZN(n6793) );
  NAND2_X1 U9367 ( .A1(n8466), .A2(n8465), .ZN(n6996) );
  NAND2_X1 U9368 ( .A1(n6793), .A2(n6792), .ZN(n6791) );
  INV_X1 U9369 ( .A(n7120), .ZN(n6794) );
  NAND3_X1 U9370 ( .A1(n6852), .A2(n6796), .A3(n6795), .ZN(P1_U3242) );
  NAND2_X1 U9371 ( .A1(n8485), .A2(n6966), .ZN(n8486) );
  NAND2_X1 U9372 ( .A1(n6966), .A2(n6576), .ZN(n6797) );
  OAI21_X1 U9373 ( .B1(n6853), .B2(n10913), .A(n8532), .ZN(n6799) );
  NAND3_X1 U9374 ( .A1(n8343), .A2(n8342), .A3(n8361), .ZN(n6800) );
  NAND3_X1 U9375 ( .A1(n6803), .A2(n6801), .A3(n6800), .ZN(n8376) );
  NAND3_X1 U9376 ( .A1(n8343), .A2(n8342), .A3(n6802), .ZN(n6803) );
  NAND3_X1 U9377 ( .A1(n6804), .A2(n8239), .A3(n7111), .ZN(n7109) );
  NAND3_X1 U9378 ( .A1(n6810), .A2(n6809), .A3(n6808), .ZN(n7127) );
  NAND3_X1 U9379 ( .A1(n6814), .A2(n6812), .A3(n6811), .ZN(n8432) );
  NAND3_X1 U9380 ( .A1(n8405), .A2(n8416), .A3(n8404), .ZN(n6811) );
  NAND3_X1 U9381 ( .A1(n8405), .A2(n8404), .A3(n6813), .ZN(n6814) );
  AND3_X1 U9382 ( .A1(n10611), .A2(n14351), .A3(n6815), .ZN(n10580) );
  AND2_X2 U9383 ( .A1(n6816), .A2(n6519), .ZN(n14351) );
  INV_X1 U9384 ( .A(n13724), .ZN(n10611) );
  OAI21_X1 U9385 ( .B1(n9247), .B2(n7373), .A(n6817), .ZN(n13724) );
  NAND2_X1 U9386 ( .A1(n9247), .A2(n13840), .ZN(n6817) );
  AND2_X2 U9387 ( .A1(n10542), .A2(n14418), .ZN(n10514) );
  NOR2_X2 U9388 ( .A1(n10545), .A2(n10541), .ZN(n10542) );
  NAND3_X1 U9389 ( .A1(n6827), .A2(n14367), .A3(n7025), .ZN(n14300) );
  INV_X1 U9390 ( .A(n10649), .ZN(n6827) );
  NAND3_X1 U9391 ( .A1(n6828), .A2(n6832), .A3(n6478), .ZN(n6831) );
  INV_X1 U9392 ( .A(n7142), .ZN(n6835) );
  OAI21_X1 U9393 ( .B1(n6840), .B2(n13953), .A(n6835), .ZN(n6837) );
  INV_X1 U9394 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6843) );
  NAND2_X1 U9395 ( .A1(n8068), .A2(n7855), .ZN(n7857) );
  NAND2_X1 U9396 ( .A1(n8221), .A2(n6982), .ZN(n7881) );
  NAND2_X1 U9397 ( .A1(n7839), .A2(n7838), .ZN(n6854) );
  NAND2_X1 U9398 ( .A1(n6586), .A2(n7839), .ZN(n6855) );
  NAND2_X1 U9399 ( .A1(n11551), .A2(n6861), .ZN(n6859) );
  NAND2_X2 U9400 ( .A1(n6860), .A2(n8461), .ZN(n13745) );
  NAND2_X1 U9401 ( .A1(n6865), .A2(n7275), .ZN(n6864) );
  NAND3_X1 U9402 ( .A1(n7277), .A2(n7276), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n6865) );
  OAI211_X2 U9403 ( .C1(n6870), .C2(n6869), .A(n7870), .B(n6872), .ZN(n8177)
         );
  NAND2_X1 U9404 ( .A1(n7257), .A2(n7863), .ZN(n6869) );
  NAND2_X1 U9405 ( .A1(n7257), .A2(n6871), .ZN(n6872) );
  INV_X1 U9406 ( .A(n7259), .ZN(n6871) );
  NAND2_X1 U9407 ( .A1(n6942), .A2(n7846), .ZN(n8033) );
  INV_X1 U9408 ( .A(n6873), .ZN(n7839) );
  NAND2_X1 U9409 ( .A1(n7873), .A2(n7872), .ZN(n8198) );
  NAND2_X1 U9410 ( .A1(n8075), .A2(n8074), .ZN(n8077) );
  NAND2_X1 U9411 ( .A1(n8091), .A2(n7860), .ZN(n8075) );
  NAND2_X1 U9412 ( .A1(n6874), .A2(n7126), .ZN(n8403) );
  NAND3_X1 U9413 ( .A1(n6899), .A2(n6541), .A3(n6898), .ZN(n6874) );
  MUX2_X1 U9414 ( .A(n8511), .B(n8512), .S(n8510), .Z(n8513) );
  NAND2_X1 U9415 ( .A1(n7172), .A2(n9050), .ZN(n10011) );
  INV_X1 U9416 ( .A(n11983), .ZN(n6885) );
  OAI21_X2 U9417 ( .B1(n14669), .B2(n7146), .A(n7144), .ZN(n9077) );
  NAND2_X2 U9418 ( .A1(n6883), .A2(n6881), .ZN(n12055) );
  NOR2_X1 U9419 ( .A1(P3_IR_REG_19__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n6882) );
  NOR2_X2 U9420 ( .A1(n7642), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n7638) );
  NAND2_X1 U9421 ( .A1(n9075), .A2(n9074), .ZN(n11069) );
  NAND2_X1 U9422 ( .A1(n7644), .A2(n7614), .ZN(n7631) );
  NAND2_X1 U9423 ( .A1(n7062), .A2(n12311), .ZN(n7060) );
  AOI21_X2 U9424 ( .B1(n7065), .B2(n7063), .A(n12203), .ZN(n7062) );
  NAND2_X1 U9425 ( .A1(n8549), .A2(n8548), .ZN(n8627) );
  NAND2_X1 U9426 ( .A1(n6886), .A2(n7589), .ZN(n12056) );
  NAND3_X1 U9427 ( .A1(n7060), .A2(n7061), .A3(n7598), .ZN(n6886) );
  XNOR2_X1 U9428 ( .A(n8919), .B(n8908), .ZN(n12651) );
  INV_X1 U9429 ( .A(n7958), .ZN(n13733) );
  INV_X1 U9430 ( .A(n11604), .ZN(n11599) );
  NAND2_X1 U9431 ( .A1(n7884), .A2(SI_18_), .ZN(n7885) );
  AOI21_X2 U9432 ( .B1(n6888), .B2(n14373), .A(n7386), .ZN(n13747) );
  NAND2_X1 U9433 ( .A1(n7389), .A2(n13554), .ZN(n6888) );
  NAND2_X1 U9434 ( .A1(n6889), .A2(n8339), .ZN(n8343) );
  NAND3_X1 U9435 ( .A1(n7112), .A2(n7110), .A3(n7109), .ZN(n6889) );
  NAND2_X1 U9436 ( .A1(n14743), .A2(n14742), .ZN(n14745) );
  NAND2_X1 U9437 ( .A1(n12441), .A2(n12443), .ZN(n12440) );
  AOI21_X1 U9438 ( .B1(n12475), .B2(n12145), .A(n8976), .ZN(n12452) );
  OAI21_X2 U9439 ( .B1(n12326), .B2(n8979), .A(n12194), .ZN(n12311) );
  NOR2_X2 U9440 ( .A1(n8538), .A2(n8537), .ZN(n8593) );
  NAND2_X1 U9441 ( .A1(n12926), .A2(n6488), .ZN(n7435) );
  NAND2_X1 U9442 ( .A1(n8198), .A2(n8197), .ZN(n7876) );
  NAND2_X1 U9443 ( .A1(n6893), .A2(n6892), .ZN(n11416) );
  NAND2_X1 U9444 ( .A1(n7535), .A2(n7536), .ZN(n11397) );
  NAND2_X1 U9445 ( .A1(n11485), .A2(n11484), .ZN(n7512) );
  NAND2_X1 U9446 ( .A1(n11366), .A2(n11365), .ZN(n11371) );
  OAI211_X1 U9447 ( .C1(n11512), .C2(n7521), .A(n7523), .B(n7519), .ZN(n11536)
         );
  OAI21_X1 U9448 ( .B1(n6957), .B2(n6956), .A(n7540), .ZN(n11406) );
  NAND2_X1 U9449 ( .A1(n6894), .A2(n11311), .ZN(n11317) );
  NAND3_X1 U9450 ( .A1(n6914), .A2(n11306), .A3(n6913), .ZN(n6894) );
  NAND2_X1 U9451 ( .A1(n7718), .A2(n7824), .ZN(n7719) );
  NAND2_X1 U9452 ( .A1(n7696), .A2(n7697), .ZN(n9961) );
  NAND2_X1 U9453 ( .A1(n12668), .A2(n12667), .ZN(n6936) );
  XNOR2_X1 U9454 ( .A(n11708), .B(n6490), .ZN(n12734) );
  XNOR2_X1 U9455 ( .A(n7083), .B(n7082), .ZN(n7739) );
  NOR2_X2 U9456 ( .A1(n12732), .A2(n7605), .ZN(n11709) );
  NAND2_X1 U9457 ( .A1(n12241), .A2(n6577), .ZN(n7338) );
  NAND2_X1 U9458 ( .A1(n12243), .A2(n7337), .ZN(n7336) );
  OAI22_X1 U9459 ( .A1(n12250), .A2(n12249), .B1(n12248), .B2(n14780), .ZN(
        n12251) );
  XNOR2_X1 U9460 ( .A(n12025), .B(n12026), .ZN(n12647) );
  NAND2_X1 U9461 ( .A1(n12647), .A2(n8611), .ZN(n7335) );
  NAND2_X1 U9462 ( .A1(n8774), .A2(n8775), .ZN(n6920) );
  NAND2_X1 U9463 ( .A1(n8865), .A2(n11122), .ZN(n7349) );
  AOI21_X1 U9464 ( .B1(n7038), .B2(n6460), .A(n7037), .ZN(n12326) );
  INV_X1 U9465 ( .A(n7076), .ZN(n7074) );
  INV_X1 U9466 ( .A(n7078), .ZN(n12899) );
  NAND2_X1 U9467 ( .A1(n8437), .A2(n8436), .ZN(n8452) );
  NAND2_X1 U9468 ( .A1(n8327), .A2(n8328), .ZN(n6900) );
  AOI21_X1 U9469 ( .B1(n7111), .B2(n6557), .A(n6900), .ZN(n7110) );
  NOR2_X2 U9470 ( .A1(n11670), .A2(n6970), .ZN(n11681) );
  OAI21_X1 U9471 ( .B1(n7204), .B2(n12862), .A(n6579), .ZN(n7202) );
  NOR2_X1 U9472 ( .A1(n12983), .A2(n12982), .ZN(n12984) );
  OAI21_X1 U9473 ( .B1(n8466), .B2(n8465), .A(n8464), .ZN(n8467) );
  INV_X1 U9474 ( .A(n13799), .ZN(n7031) );
  NAND2_X1 U9475 ( .A1(n8484), .A2(n8483), .ZN(n6966) );
  NAND2_X1 U9476 ( .A1(n6995), .A2(n6994), .ZN(n6898) );
  NAND2_X1 U9477 ( .A1(n8374), .A2(n8373), .ZN(n6899) );
  NAND2_X1 U9478 ( .A1(n6989), .A2(n8121), .ZN(n8123) );
  INV_X1 U9479 ( .A(n7304), .ZN(n7303) );
  AOI21_X1 U9480 ( .B1(n7303), .B2(n7305), .A(n6573), .ZN(n7301) );
  NAND2_X1 U9481 ( .A1(n7256), .A2(n7259), .ZN(n8160) );
  OAI21_X1 U9482 ( .B1(n10511), .B2(n7305), .A(n10794), .ZN(n7304) );
  NAND2_X1 U9483 ( .A1(n7314), .A2(n7313), .ZN(n13653) );
  NAND2_X1 U9484 ( .A1(n6904), .A2(n6902), .ZN(P1_U3214) );
  NAND2_X1 U9485 ( .A1(n6910), .A2(n13320), .ZN(n6904) );
  INV_X1 U9486 ( .A(n9903), .ZN(n7246) );
  NOR2_X1 U9487 ( .A1(n13538), .A2(n6906), .ZN(n6954) );
  NAND4_X1 U9488 ( .A1(n8503), .A2(n13576), .A3(n13555), .A4(n13601), .ZN(
        n6906) );
  NOR2_X1 U9489 ( .A1(n14033), .A2(n6566), .ZN(n7831) );
  OR2_X1 U9490 ( .A1(n7833), .A2(n14036), .ZN(n7834) );
  OAI21_X1 U9491 ( .B1(n13218), .B2(n13219), .A(n13217), .ZN(n6910) );
  NOR2_X1 U9492 ( .A1(n12811), .A2(n12812), .ZN(n12813) );
  NAND2_X1 U9493 ( .A1(n10707), .A2(n10708), .ZN(n10878) );
  NAND2_X1 U9494 ( .A1(n10006), .A2(n10005), .ZN(n10527) );
  NAND3_X1 U9495 ( .A1(n6916), .A2(n6588), .A3(n6912), .ZN(n7287) );
  OR2_X1 U9496 ( .A1(n11623), .A2(n11624), .ZN(n6912) );
  NAND2_X1 U9497 ( .A1(n8468), .A2(n6984), .ZN(n13824) );
  INV_X1 U9498 ( .A(n7394), .ZN(n7393) );
  INV_X1 U9499 ( .A(n7401), .ZN(n13624) );
  INV_X1 U9500 ( .A(n8513), .ZN(n8514) );
  NAND2_X1 U9501 ( .A1(n13742), .A2(n14373), .ZN(n6948) );
  OAI21_X1 U9502 ( .B1(n13666), .B2(n7393), .A(n7391), .ZN(n7401) );
  NAND2_X1 U9503 ( .A1(n7953), .A2(n8017), .ZN(n6939) );
  NAND2_X1 U9504 ( .A1(n7288), .A2(n11599), .ZN(n6916) );
  NAND2_X1 U9505 ( .A1(n11305), .A2(n11304), .ZN(n6913) );
  NAND2_X1 U9506 ( .A1(n11298), .A2(n11297), .ZN(n6914) );
  NAND2_X1 U9507 ( .A1(n6915), .A2(n6988), .ZN(n7117) );
  NAND2_X1 U9508 ( .A1(n8452), .A2(n8451), .ZN(n6915) );
  NAND2_X1 U9509 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n6922), .ZN(n6921) );
  NOR2_X1 U9510 ( .A1(n12312), .A2(n8980), .ZN(n7068) );
  NAND2_X1 U9511 ( .A1(n7062), .A2(n7064), .ZN(n7061) );
  XNOR2_X1 U9512 ( .A(n6923), .B(n8226), .ZN(n11024) );
  OAI21_X1 U9513 ( .B1(n12925), .B2(n6479), .A(n6580), .ZN(n6993) );
  XNOR2_X1 U9514 ( .A(n12885), .B(n6976), .ZN(n13091) );
  XNOR2_X2 U9515 ( .A(n13156), .B(n11030), .ZN(n12832) );
  NAND2_X1 U9516 ( .A1(n6927), .A2(n6925), .ZN(n12208) );
  AOI21_X1 U9517 ( .B1(n6510), .B2(n12076), .A(n6926), .ZN(n6925) );
  NAND2_X1 U9518 ( .A1(n12204), .A2(n12205), .ZN(n6926) );
  OR2_X1 U9519 ( .A1(n12202), .A2(n12076), .ZN(n6927) );
  NAND2_X1 U9520 ( .A1(n11279), .A2(n12042), .ZN(n6965) );
  NOR2_X2 U9521 ( .A1(n9829), .A2(n9024), .ZN(n7474) );
  NAND2_X1 U9522 ( .A1(n10218), .A2(n10217), .ZN(n7190) );
  INV_X1 U9523 ( .A(n13885), .ZN(n7140) );
  NAND2_X1 U9524 ( .A1(n14016), .A2(n7762), .ZN(n14031) );
  NAND2_X1 U9525 ( .A1(n14017), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n14016) );
  NAND2_X1 U9526 ( .A1(n10918), .A2(n7758), .ZN(n11080) );
  NAND2_X1 U9527 ( .A1(n6935), .A2(n11284), .ZN(n11288) );
  NAND3_X1 U9528 ( .A1(n6936), .A2(n12669), .A3(n12763), .ZN(n12673) );
  OAI21_X2 U9529 ( .B1(n10754), .B2(n7011), .A(n7009), .ZN(n11175) );
  NAND2_X1 U9530 ( .A1(n11300), .A2(n11299), .ZN(n11307) );
  NAND2_X1 U9531 ( .A1(n7482), .A2(n7483), .ZN(n12682) );
  NAND2_X1 U9532 ( .A1(n9288), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n6992) );
  NAND2_X1 U9533 ( .A1(n12674), .A2(n12676), .ZN(n12675) );
  NAND2_X1 U9534 ( .A1(n8076), .A2(n8077), .ZN(n10085) );
  NAND2_X1 U9535 ( .A1(n6977), .A2(n6971), .ZN(n6970) );
  NAND2_X1 U9536 ( .A1(n11527), .A2(n8414), .ZN(n6937) );
  OAI211_X1 U9537 ( .C1(n13743), .C2(n14368), .A(n6948), .B(n6575), .ZN(n13806) );
  NAND2_X1 U9538 ( .A1(n6962), .A2(n6959), .ZN(n8404) );
  XNOR2_X2 U9539 ( .A(n8383), .B(SI_23_), .ZN(n11499) );
  OAI211_X1 U9540 ( .C1(n13091), .C2(n14583), .A(n13090), .B(n13089), .ZN(
        n13178) );
  INV_X1 U9541 ( .A(n13110), .ZN(n12879) );
  NAND2_X1 U9542 ( .A1(n7893), .A2(n11277), .ZN(n7896) );
  NAND2_X1 U9543 ( .A1(n12912), .A2(n7435), .ZN(n7434) );
  INV_X1 U9544 ( .A(n6993), .ZN(n12913) );
  OAI21_X2 U9545 ( .B1(n8413), .B2(n8412), .A(n7905), .ZN(n8427) );
  NAND2_X1 U9546 ( .A1(n11343), .A2(n11344), .ZN(n11349) );
  INV_X1 U9547 ( .A(n11669), .ZN(n6977) );
  INV_X1 U9548 ( .A(n6951), .ZN(n6950) );
  AOI21_X1 U9549 ( .B1(n13004), .B2(n13012), .A(n7426), .ZN(n12989) );
  OAI22_X2 U9550 ( .A1(n12944), .A2(n12842), .B1(n13110), .B2(n12878), .ZN(
        n12931) );
  NAND2_X1 U9551 ( .A1(n8003), .A2(n7845), .ZN(n6942) );
  NAND3_X1 U9552 ( .A1(n7427), .A2(n7428), .A3(n12844), .ZN(n12845) );
  NAND2_X1 U9553 ( .A1(n12989), .A2(n6572), .ZN(n7425) );
  AOI22_X2 U9554 ( .A1(n12962), .A2(n12841), .B1(n12876), .B2(n13116), .ZN(
        n12944) );
  AOI22_X2 U9555 ( .A1(n12931), .A2(n12930), .B1(n12843), .B2(n13105), .ZN(
        n12917) );
  AOI21_X1 U9556 ( .B1(n6945), .B2(n14554), .A(n6943), .ZN(n7217) );
  INV_X1 U9557 ( .A(n13090), .ZN(n6945) );
  AOI21_X2 U9558 ( .B1(n14397), .B2(n13745), .A(n13744), .ZN(n13746) );
  OR2_X2 U9559 ( .A1(n13763), .A2(n13629), .ZN(n13606) );
  NAND2_X1 U9560 ( .A1(n12303), .A2(n8918), .ZN(n8927) );
  NAND2_X1 U9561 ( .A1(n7569), .A2(n7568), .ZN(n12361) );
  NAND2_X1 U9562 ( .A1(n13570), .A2(n13576), .ZN(n13569) );
  XNOR2_X1 U9563 ( .A(n6947), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND2_X1 U9564 ( .A1(n6949), .A2(n12242), .ZN(n12191) );
  NAND2_X1 U9565 ( .A1(n6963), .A2(n12187), .ZN(n6949) );
  NAND2_X1 U9566 ( .A1(n7881), .A2(n7880), .ZN(n8247) );
  AND2_X2 U9567 ( .A1(n7602), .A2(n12924), .ZN(n12921) );
  OAI22_X1 U9568 ( .A1(n9511), .A2(n9302), .B1(n11026), .B2(n9301), .ZN(n6951)
         );
  NAND2_X1 U9569 ( .A1(n10124), .A2(n14588), .ZN(n10143) );
  NAND2_X1 U9570 ( .A1(n13007), .A2(n12998), .ZN(n12993) );
  NAND2_X1 U9571 ( .A1(n12908), .A2(n12899), .ZN(n12895) );
  XNOR2_X1 U9572 ( .A(n11709), .B(n11710), .ZN(n12674) );
  INV_X1 U9573 ( .A(n7012), .ZN(n7011) );
  NAND2_X2 U9574 ( .A1(n12753), .A2(n12752), .ZN(n12751) );
  NAND2_X1 U9575 ( .A1(n11302), .A2(n11303), .ZN(n11298) );
  NAND2_X1 U9576 ( .A1(n11292), .A2(n11291), .ZN(n11302) );
  NOR2_X1 U9577 ( .A1(n11508), .A2(n11509), .ZN(n11512) );
  OAI21_X1 U9578 ( .B1(n11397), .B2(n11396), .A(n6585), .ZN(n6956) );
  AOI21_X1 U9579 ( .B1(n6958), .B2(n6981), .A(n11598), .ZN(n7288) );
  NAND2_X1 U9580 ( .A1(n11480), .A2(n11481), .ZN(n11479) );
  NAND2_X1 U9581 ( .A1(n11317), .A2(n11318), .ZN(n11316) );
  NAND2_X1 U9582 ( .A1(n11550), .A2(n11549), .ZN(n6958) );
  INV_X1 U9583 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7277) );
  INV_X1 U9584 ( .A(n8376), .ZN(n6995) );
  XNOR2_X1 U9585 ( .A(n13884), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15025) );
  NAND2_X1 U9586 ( .A1(n6964), .A2(n12350), .ZN(n6963) );
  INV_X1 U9587 ( .A(n12188), .ZN(n6964) );
  NAND2_X1 U9588 ( .A1(n8462), .A2(n8463), .ZN(n7120) );
  NAND2_X1 U9589 ( .A1(n6968), .A2(n11153), .ZN(n13524) );
  INV_X1 U9590 ( .A(n11152), .ZN(n6968) );
  NAND2_X1 U9591 ( .A1(n13677), .A2(n13684), .ZN(n13676) );
  OAI21_X1 U9592 ( .B1(n10409), .B2(n7377), .A(n7375), .ZN(n10793) );
  OAI21_X1 U9593 ( .B1(n7378), .B2(n7377), .A(n10790), .ZN(n7376) );
  NOR2_X1 U9594 ( .A1(n13936), .A2(n13937), .ZN(n13987) );
  NAND2_X1 U9595 ( .A1(n12937), .A2(n7208), .ZN(n12925) );
  NAND2_X1 U9596 ( .A1(n10050), .A2(n10049), .ZN(n10117) );
  NAND3_X1 U9597 ( .A1(n11416), .A2(n6570), .A3(n6475), .ZN(n7543) );
  NAND3_X1 U9598 ( .A1(n11386), .A2(n7608), .A3(n6571), .ZN(n7535) );
  NAND2_X1 U9599 ( .A1(n8506), .A2(n8505), .ZN(n8515) );
  NAND2_X1 U9600 ( .A1(n11287), .A2(n6978), .ZN(n11303) );
  INV_X1 U9601 ( .A(n11303), .ZN(n11304) );
  NAND2_X1 U9602 ( .A1(n11682), .A2(n7517), .ZN(n7515) );
  NOR2_X1 U9603 ( .A1(n12889), .A2(n6973), .ZN(n6972) );
  NAND2_X1 U9604 ( .A1(n6975), .A2(n6974), .ZN(n6973) );
  NOR2_X1 U9605 ( .A1(n11668), .A2(n12938), .ZN(n6974) );
  INV_X1 U9606 ( .A(n12926), .ZN(n6975) );
  NOR2_X1 U9607 ( .A1(n6980), .A2(n6979), .ZN(n6978) );
  NAND2_X1 U9608 ( .A1(n8470), .A2(n8469), .ZN(n6984) );
  NOR2_X1 U9609 ( .A1(n13986), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n13988) );
  NAND2_X1 U9610 ( .A1(n15025), .A2(n15024), .ZN(n13896) );
  OAI21_X1 U9611 ( .B1(n7847), .B2(n6987), .A(n6986), .ZN(n7841) );
  XNOR2_X2 U9612 ( .A(n7898), .B(n7897), .ZN(n8383) );
  INV_X1 U9613 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7276) );
  NAND2_X1 U9614 ( .A1(n7285), .A2(n7286), .ZN(n8447) );
  OAI21_X1 U9615 ( .B1(n13091), .B2(n13081), .A(n7217), .ZN(P2_U3236) );
  NAND2_X1 U9616 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  NAND3_X1 U9617 ( .A1(n7835), .A2(n7834), .A3(n7836), .ZN(P3_U3201) );
  NAND2_X1 U9618 ( .A1(n8833), .A2(n7344), .ZN(n7342) );
  NAND2_X1 U9619 ( .A1(n8813), .A2(n8814), .ZN(n7327) );
  OAI21_X1 U9620 ( .B1(n11334), .B2(n7529), .A(n7531), .ZN(n11341) );
  AOI21_X1 U9621 ( .B1(n11385), .B2(n11384), .A(n11382), .ZN(n11383) );
  NAND2_X2 U9622 ( .A1(n7876), .A2(n7875), .ZN(n8221) );
  NAND2_X1 U9623 ( .A1(n8467), .A2(n6996), .ZN(n8484) );
  NAND3_X1 U9624 ( .A1(n7476), .A2(n9629), .A3(n9619), .ZN(n9804) );
  NAND2_X1 U9625 ( .A1(n10093), .A2(n6463), .ZN(n7001) );
  INV_X1 U9626 ( .A(n7000), .ZN(n6999) );
  NAND2_X1 U9627 ( .A1(n9970), .A2(n7004), .ZN(n7003) );
  AOI21_X1 U9628 ( .B1(n9971), .B2(n9976), .A(n7008), .ZN(n7007) );
  NAND2_X1 U9629 ( .A1(n12682), .A2(n7018), .ZN(n7016) );
  INV_X4 U9630 ( .A(n9299), .ZN(n9154) );
  MUX2_X1 U9631 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n9299), .Z(n7854) );
  MUX2_X1 U9632 ( .A(n9721), .B(n8570), .S(n9299), .Z(n8210) );
  MUX2_X1 U9633 ( .A(n11025), .B(n9900), .S(n9299), .Z(n8225) );
  MUX2_X1 U9634 ( .A(n10759), .B(n8567), .S(n9299), .Z(n7874) );
  MUX2_X1 U9635 ( .A(n9834), .B(n9793), .S(n9299), .Z(n8261) );
  NAND2_X1 U9636 ( .A1(n7893), .A2(n9299), .ZN(n8372) );
  NOR2_X2 U9637 ( .A1(n13973), .A2(n14145), .ZN(n7027) );
  NOR2_X2 U9638 ( .A1(n13592), .A2(n7033), .ZN(n13541) );
  NAND2_X1 U9639 ( .A1(n7668), .A2(n7035), .ZN(n7670) );
  NAND2_X1 U9640 ( .A1(n14767), .A2(n12279), .ZN(n12085) );
  INV_X2 U9641 ( .A(n12279), .ZN(n10463) );
  INV_X1 U9642 ( .A(n12359), .ZN(n7038) );
  NOR2_X2 U9643 ( .A1(n8917), .A2(n7068), .ZN(n7067) );
  NOR2_X2 U9644 ( .A1(n10213), .A2(n14601), .ZN(n10289) );
  OR2_X2 U9645 ( .A1(n10143), .A2(n11331), .ZN(n10213) );
  NOR2_X2 U9646 ( .A1(n10164), .A2(n14579), .ZN(n10124) );
  AND2_X1 U9647 ( .A1(n12921), .A2(n7074), .ZN(n12852) );
  AND2_X1 U9648 ( .A1(n12921), .A2(n12911), .ZN(n12908) );
  NAND2_X1 U9649 ( .A1(n12921), .A2(n7075), .ZN(n12828) );
  NOR2_X4 U9650 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7668) );
  INV_X1 U9651 ( .A(n7691), .ZN(n7091) );
  NAND2_X1 U9652 ( .A1(n7087), .A2(n9923), .ZN(n7088) );
  INV_X1 U9653 ( .A(n9788), .ZN(n7090) );
  NAND2_X1 U9654 ( .A1(n7698), .A2(n7097), .ZN(n7095) );
  NAND2_X1 U9655 ( .A1(n7094), .A2(n7092), .ZN(n7711) );
  INV_X1 U9656 ( .A(n7101), .ZN(n10674) );
  NAND2_X1 U9657 ( .A1(n9726), .A2(n9727), .ZN(n9725) );
  NAND2_X1 U9658 ( .A1(n9725), .A2(n7677), .ZN(n7681) );
  INV_X2 U9659 ( .A(n7108), .ZN(n13354) );
  NAND2_X1 U9660 ( .A1(n10619), .A2(n7108), .ZN(n9705) );
  NAND2_X1 U9661 ( .A1(n7108), .A2(n14351), .ZN(n9698) );
  AND2_X1 U9662 ( .A1(n13354), .A2(n6454), .ZN(n13726) );
  NAND2_X1 U9663 ( .A1(n13354), .A2(n6436), .ZN(n7107) );
  OAI22_X1 U9664 ( .A1(n11815), .A2(n7108), .B1(n14351), .B2(n11823), .ZN(
        n9891) );
  OAI22_X1 U9665 ( .A1(n10572), .A2(n13965), .B1(n7108), .B2(n13963), .ZN(
        n10573) );
  XNOR2_X1 U9666 ( .A(n14353), .B(n7108), .ZN(n10612) );
  NAND2_X1 U9667 ( .A1(n7109), .A2(n7110), .ZN(n8341) );
  NAND3_X1 U9668 ( .A1(n8021), .A2(n10375), .A3(n8020), .ZN(n7116) );
  NAND2_X1 U9669 ( .A1(n7127), .A2(n8114), .ZN(n8131) );
  NAND3_X1 U9670 ( .A1(n8189), .A2(n8188), .A3(n7131), .ZN(n7130) );
  NAND2_X1 U9671 ( .A1(n13930), .A2(n13929), .ZN(n13934) );
  INV_X1 U9672 ( .A(n9077), .ZN(n9075) );
  NAND2_X1 U9673 ( .A1(n12007), .A2(n6509), .ZN(n7147) );
  OAI211_X1 U9674 ( .C1(n12007), .C2(n7151), .A(n7148), .B(n7147), .ZN(n7157)
         );
  AOI21_X1 U9675 ( .B1(n12007), .B2(n12008), .A(n7158), .ZN(n11919) );
  OAI21_X1 U9676 ( .B1(n11920), .B2(n7155), .A(n6487), .ZN(n7150) );
  NAND2_X1 U9677 ( .A1(n7157), .A2(n11924), .ZN(P3_U3160) );
  INV_X1 U9678 ( .A(n12016), .ZN(n7169) );
  NAND2_X1 U9679 ( .A1(n10010), .A2(n10011), .ZN(n9053) );
  NAND2_X1 U9680 ( .A1(n9049), .A2(n9046), .ZN(n7172) );
  NAND2_X1 U9681 ( .A1(n7181), .A2(n7180), .ZN(n11249) );
  NAND2_X1 U9682 ( .A1(n11069), .A2(n7182), .ZN(n11211) );
  NAND2_X1 U9683 ( .A1(n13236), .A2(n7223), .ZN(n7222) );
  NAND2_X1 U9684 ( .A1(n7239), .A2(n7240), .ZN(n11862) );
  NAND2_X1 U9685 ( .A1(n13318), .A2(n7241), .ZN(n7239) );
  XNOR2_X1 U9686 ( .A(n10301), .B(n10302), .ZN(n10340) );
  NAND2_X1 U9687 ( .A1(n7250), .A2(n7251), .ZN(n9906) );
  NAND2_X1 U9688 ( .A1(n7122), .A2(n7413), .ZN(n7947) );
  NAND2_X1 U9689 ( .A1(n7886), .A2(n7273), .ZN(n7270) );
  NAND2_X1 U9690 ( .A1(n7886), .A2(n7885), .ZN(n8292) );
  NAND2_X1 U9691 ( .A1(n8427), .A2(n6612), .ZN(n7285) );
  NAND2_X1 U9692 ( .A1(n7913), .A2(n7912), .ZN(n8470) );
  INV_X1 U9693 ( .A(n8469), .ZN(n7291) );
  OAI22_X1 U9694 ( .A1(n11903), .A2(n12267), .B1(n11266), .B2(n11267), .ZN(
        n11270) );
  NAND2_X1 U9695 ( .A1(n6587), .A2(n7292), .ZN(n10373) );
  NAND2_X1 U9696 ( .A1(n10369), .A2(n7294), .ZN(n7292) );
  INV_X1 U9697 ( .A(n7308), .ZN(n13574) );
  NOR2_X1 U9698 ( .A1(n15021), .A2(n13756), .ZN(n7310) );
  NAND2_X1 U9699 ( .A1(n13683), .A2(n7315), .ZN(n7314) );
  NAND2_X1 U9700 ( .A1(n13653), .A2(n13654), .ZN(n13515) );
  NAND2_X1 U9701 ( .A1(n10614), .A2(n9698), .ZN(n10570) );
  AND2_X2 U9702 ( .A1(n7352), .A2(n7351), .ZN(n14533) );
  NOR2_X2 U9703 ( .A1(n14529), .A2(n14528), .ZN(n14526) );
  NOR2_X2 U9704 ( .A1(n14505), .A2(n12789), .ZN(n14519) );
  NAND2_X1 U9705 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(n7372), .ZN(n7995) );
  NAND2_X1 U9706 ( .A1(n10809), .A2(n7382), .ZN(n7381) );
  NAND2_X1 U9707 ( .A1(n7381), .A2(n7380), .ZN(n10995) );
  INV_X1 U9708 ( .A(n13638), .ZN(n7395) );
  NAND2_X1 U9709 ( .A1(n13793), .A2(n13678), .ZN(n7403) );
  AOI21_X2 U9710 ( .B1(n10443), .B2(n10407), .A(n10406), .ZN(n10537) );
  AOI21_X2 U9711 ( .B1(n6489), .B2(n7406), .A(n7404), .ZN(n13677) );
  INV_X1 U9712 ( .A(n7933), .ZN(n7412) );
  INV_X1 U9713 ( .A(n7925), .ZN(n7416) );
  NAND2_X1 U9714 ( .A1(n7925), .A2(n7931), .ZN(n7414) );
  NAND3_X1 U9715 ( .A1(n7412), .A2(n7925), .A3(n7931), .ZN(n7411) );
  NOR2_X1 U9716 ( .A1(n7922), .A2(n8034), .ZN(n8227) );
  OAI21_X2 U9717 ( .B1(n10497), .B2(n10383), .A(n10382), .ZN(n14292) );
  OAI21_X2 U9718 ( .B1(n10648), .B2(n10379), .A(n10380), .ZN(n10497) );
  NAND2_X1 U9719 ( .A1(n10378), .A2(n10377), .ZN(n10648) );
  NOR2_X1 U9720 ( .A1(n7418), .A2(n11671), .ZN(n7417) );
  XNOR2_X1 U9721 ( .A(n9577), .B(n7418), .ZN(n9580) );
  XNOR2_X1 U9722 ( .A(n7418), .B(n10045), .ZN(n10162) );
  NAND2_X1 U9723 ( .A1(n12917), .A2(n7430), .ZN(n7427) );
  NAND2_X1 U9724 ( .A1(n12917), .A2(n7431), .ZN(n7429) );
  NAND2_X1 U9725 ( .A1(n11023), .A2(n7442), .ZN(n7441) );
  NOR2_X2 U9726 ( .A1(n7454), .A2(n7452), .ZN(n7451) );
  NAND2_X1 U9727 ( .A1(n7465), .A2(n10319), .ZN(n7461) );
  NAND2_X1 U9728 ( .A1(n7463), .A2(n10319), .ZN(n7462) );
  NOR2_X1 U9729 ( .A1(n10736), .A2(n12773), .ZN(n7473) );
  AND2_X1 U9731 ( .A1(n9025), .A2(n9026), .ZN(n9824) );
  NAND2_X1 U9732 ( .A1(n12717), .A2(n7481), .ZN(n7479) );
  AND2_X2 U9733 ( .A1(n7479), .A2(n7477), .ZN(n12753) );
  INV_X1 U9734 ( .A(n12710), .ZN(n7485) );
  NAND2_X1 U9735 ( .A1(n12710), .A2(n7490), .ZN(n7482) );
  NAND2_X1 U9736 ( .A1(n12751), .A2(n6569), .ZN(n7491) );
  OAI211_X1 U9737 ( .C1(n12751), .C2(n7495), .A(n7491), .B(n7492), .ZN(n11737)
         );
  NAND2_X1 U9738 ( .A1(n12751), .A2(n7498), .ZN(n12668) );
  NAND2_X1 U9739 ( .A1(n10187), .A2(n10188), .ZN(n10267) );
  NAND2_X1 U9740 ( .A1(n10267), .A2(n7506), .ZN(n10485) );
  NAND2_X1 U9741 ( .A1(n9858), .A2(n9857), .ZN(n9970) );
  INV_X1 U9742 ( .A(n11496), .ZN(n7511) );
  NAND2_X1 U9743 ( .A1(n11675), .A2(n7518), .ZN(n7517) );
  NAND2_X1 U9744 ( .A1(n11536), .A2(n11535), .ZN(n11549) );
  NAND2_X1 U9745 ( .A1(n7527), .A2(n7526), .ZN(n11340) );
  NAND2_X1 U9746 ( .A1(n11332), .A2(n11333), .ZN(n7530) );
  NAND2_X1 U9747 ( .A1(n11334), .A2(n7531), .ZN(n7527) );
  INV_X1 U9748 ( .A(n11332), .ZN(n7528) );
  INV_X1 U9749 ( .A(n11378), .ZN(n7533) );
  NAND2_X1 U9750 ( .A1(n7539), .A2(n7538), .ZN(n7537) );
  INV_X1 U9751 ( .A(n11352), .ZN(n7539) );
  INV_X1 U9752 ( .A(n11400), .ZN(n7542) );
  NAND2_X1 U9753 ( .A1(n7543), .A2(n6583), .ZN(n11447) );
  NAND2_X1 U9754 ( .A1(n8904), .A2(n7546), .ZN(n12303) );
  NAND3_X1 U9755 ( .A1(n7548), .A2(n8605), .A3(n8618), .ZN(n10464) );
  NAND2_X1 U9756 ( .A1(n12455), .A2(n6468), .ZN(n7555) );
  NAND2_X1 U9757 ( .A1(n12405), .A2(n7570), .ZN(n7569) );
  OAI21_X2 U9758 ( .B1(n10864), .B2(n7584), .A(n7580), .ZN(n14728) );
  NAND2_X1 U9759 ( .A1(n7734), .A2(n6505), .ZN(n12068) );
  OAI21_X1 U9760 ( .B1(n14084), .B2(n14099), .A(n11151), .ZN(n11152) );
  CLKBUF_X1 U9761 ( .A(n9126), .Z(n9323) );
  NAND2_X1 U9762 ( .A1(n9517), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U9763 ( .A1(n8798), .A2(n8797), .ZN(n12414) );
  INV_X1 U9764 ( .A(n12414), .ZN(n12415) );
  INV_X1 U9765 ( .A(n11361), .ZN(n11364) );
  INV_X1 U9766 ( .A(n14763), .ZN(n9045) );
  INV_X1 U9767 ( .A(n11480), .ZN(n11483) );
  OAI21_X1 U9768 ( .B1(n11536), .B2(n11535), .A(n11534), .ZN(n11550) );
  AND2_X1 U9769 ( .A1(n12243), .A2(n12054), .ZN(n7589) );
  NOR3_X1 U9770 ( .A1(n12908), .A2(n12907), .A3(n9339), .ZN(n7590) );
  OR2_X1 U9771 ( .A1(n8351), .A2(SI_20_), .ZN(n7591) );
  INV_X1 U9772 ( .A(n12300), .ZN(n8917) );
  AND4_X1 U9773 ( .A1(n8901), .A2(n8900), .A3(n8899), .A4(n8898), .ZN(n12009)
         );
  AND2_X1 U9774 ( .A1(n8471), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n7594) );
  INV_X1 U9775 ( .A(n14015), .ZN(n9591) );
  AND2_X1 U9776 ( .A1(n11236), .A2(n8974), .ZN(n7595) );
  INV_X1 U9777 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11449) );
  INV_X1 U9778 ( .A(n12214), .ZN(n12053) );
  INV_X1 U9779 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n13816) );
  AND2_X1 U9780 ( .A1(n12215), .A2(n12048), .ZN(n7598) );
  INV_X1 U9781 ( .A(n10913), .ZN(n8520) );
  INV_X2 U9782 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13197) );
  INV_X1 U9783 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7948) );
  NOR2_X1 U9784 ( .A1(n8682), .A2(n8671), .ZN(n7599) );
  NAND2_X1 U9785 ( .A1(n11895), .A2(n12272), .ZN(n7600) );
  OR2_X1 U9786 ( .A1(n8849), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7601) );
  INV_X1 U9787 ( .A(n9354), .ZN(n11573) );
  INV_X1 U9788 ( .A(n11877), .ZN(n11266) );
  AND2_X1 U9789 ( .A1(n12321), .A2(n12500), .ZN(n7603) );
  NOR3_X1 U9790 ( .A1(n12921), .A2(n12920), .A3(n9339), .ZN(n7604) );
  NAND2_X2 U9791 ( .A1(n10055), .A2(n13071), .ZN(n14554) );
  CLKBUF_X2 U9792 ( .A(P2_U3947), .Z(n12783) );
  AND2_X1 U9793 ( .A1(n11708), .A2(n6490), .ZN(n7605) );
  OR2_X1 U9794 ( .A1(n8356), .A2(SI_21_), .ZN(n7606) );
  NOR3_X1 U9795 ( .A1(n13641), .A2(n13640), .A3(n14352), .ZN(n7607) );
  INV_X1 U9796 ( .A(n9313), .ZN(n11235) );
  AND2_X1 U9797 ( .A1(n13546), .A2(n14093), .ZN(n14315) );
  INV_X1 U9798 ( .A(n11302), .ZN(n11305) );
  INV_X1 U9799 ( .A(n11318), .ZN(n11319) );
  MUX2_X1 U9800 ( .A(n9703), .B(n9705), .S(n8399), .Z(n7991) );
  INV_X1 U9801 ( .A(n11362), .ZN(n11363) );
  OR2_X1 U9802 ( .A1(n8058), .A2(n8057), .ZN(n8059) );
  INV_X1 U9803 ( .A(n11377), .ZN(n11379) );
  INV_X1 U9804 ( .A(n11430), .ZN(n11431) );
  INV_X1 U9805 ( .A(n11481), .ZN(n11482) );
  AOI22_X1 U9806 ( .A1(n13116), .A2(n6449), .B1(n6443), .B2(n12877), .ZN(
        n11511) );
  INV_X1 U9807 ( .A(n11524), .ZN(n11526) );
  INV_X1 U9808 ( .A(n12051), .ZN(n12052) );
  NAND2_X1 U9809 ( .A1(n12053), .A2(n12052), .ZN(n12054) );
  INV_X1 U9810 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n9023) );
  INV_X1 U9811 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7930) );
  OR2_X1 U9812 ( .A1(n7695), .A2(n9964), .ZN(n7696) );
  INV_X1 U9813 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10424) );
  XNOR2_X1 U9814 ( .A(n9331), .B(n11638), .ZN(n9332) );
  NOR2_X1 U9815 ( .A1(n14300), .A2(n10559), .ZN(n10391) );
  NOR2_X1 U9816 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8161) );
  NOR2_X1 U9817 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(n7601), .ZN(n8871) );
  OR2_X1 U9818 ( .A1(n8707), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8720) );
  OAI21_X1 U9819 ( .B1(n7711), .B2(n9178), .A(n7710), .ZN(n14681) );
  OR2_X1 U9820 ( .A1(n8792), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8805) );
  AND2_X1 U9821 ( .A1(n12634), .A2(n11980), .ZN(n12138) );
  OR2_X1 U9822 ( .A1(n12634), .A2(n11980), .ZN(n12136) );
  INV_X1 U9823 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n8561) );
  INV_X1 U9824 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9980) );
  BUF_X1 U9825 ( .A(n9510), .Z(n11729) );
  INV_X1 U9826 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n11181) );
  INV_X1 U9827 ( .A(n13201), .ZN(n9312) );
  INV_X1 U9828 ( .A(n11671), .ZN(n11646) );
  INV_X1 U9829 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n8215) );
  INV_X1 U9830 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n8096) );
  OR2_X1 U9831 ( .A1(n8330), .A2(n8329), .ZN(n8344) );
  INV_X1 U9832 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8231) );
  INV_X1 U9833 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9606) );
  NAND2_X1 U9834 ( .A1(n13838), .A2(n9542), .ZN(n9846) );
  INV_X1 U9835 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7940) );
  NOR2_X1 U9836 ( .A1(n13907), .A2(n14911), .ZN(n13851) );
  OAI21_X1 U9837 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14916), .A(n13863), .ZN(
        n13870) );
  AND2_X1 U9838 ( .A1(n8943), .A2(n7625), .ZN(n7626) );
  INV_X1 U9839 ( .A(n10072), .ZN(n9055) );
  INV_X1 U9840 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n10033) );
  NAND2_X1 U9841 ( .A1(n12281), .A2(n10023), .ZN(n14776) );
  INV_X1 U9842 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8633) );
  OR2_X1 U9843 ( .A1(n8606), .A2(n11888), .ZN(n8898) );
  INV_X1 U9844 ( .A(n12321), .ZN(n12325) );
  NAND2_X1 U9845 ( .A1(n8828), .A2(n11929), .ZN(n8837) );
  AND2_X1 U9846 ( .A1(n12126), .A2(n12130), .ZN(n12229) );
  INV_X1 U9847 ( .A(n12637), .ZN(n9004) );
  INV_X1 U9848 ( .A(n12363), .ZN(n12384) );
  AND2_X1 U9849 ( .A1(n9006), .A2(n12212), .ZN(n12418) );
  NAND2_X1 U9850 ( .A1(n8942), .A2(n8943), .ZN(n8946) );
  INV_X1 U9851 ( .A(n11556), .ZN(n11589) );
  NAND2_X1 U9852 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(n11518), .ZN(n11543) );
  INV_X1 U9853 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10768) );
  AND2_X1 U9854 ( .A1(n11559), .A2(n11558), .ZN(n11732) );
  AND2_X1 U9855 ( .A1(n11452), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11468) );
  AND2_X1 U9856 ( .A1(n11420), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11437) );
  INV_X1 U9857 ( .A(n12824), .ZN(n12756) );
  NAND2_X1 U9858 ( .A1(n9330), .A2(n11671), .ZN(n11638) );
  INV_X1 U9859 ( .A(n11374), .ZN(n10736) );
  OAI21_X1 U9860 ( .B1(n9032), .B2(P2_IR_REG_25__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U9861 ( .A1(n10965), .A2(n10964), .ZN(n10966) );
  INV_X1 U9862 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n8082) );
  AND2_X1 U9863 ( .A1(n10301), .A2(n10302), .ZN(n10303) );
  INV_X1 U9864 ( .A(n8407), .ZN(n8389) );
  AND2_X1 U9865 ( .A1(n13234), .A2(n11810), .ZN(n13301) );
  NAND2_X1 U9866 ( .A1(n8252), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8313) );
  NOR2_X1 U9867 ( .A1(n8344), .A2(n13257), .ZN(n8363) );
  INV_X1 U9868 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n13877) );
  INV_X1 U9869 ( .A(n13601), .ZN(n13603) );
  INV_X1 U9870 ( .A(n13342), .ZN(n11200) );
  INV_X1 U9871 ( .A(n9846), .ZN(n9246) );
  INV_X1 U9872 ( .A(n9852), .ZN(n10361) );
  AND2_X1 U9873 ( .A1(n8022), .A2(n10377), .ZN(n10375) );
  OR2_X1 U9874 ( .A1(n14322), .A2(n10365), .ZN(n10576) );
  INV_X1 U9875 ( .A(n11149), .ZN(n14099) );
  INV_X1 U9876 ( .A(n10790), .ZN(n10794) );
  INV_X1 U9877 ( .A(n10410), .ZN(n10511) );
  AND2_X1 U9878 ( .A1(n9568), .A2(n9567), .ZN(n10359) );
  OAI22_X1 U9879 ( .A1(n13905), .A2(n13849), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n13848), .ZN(n13850) );
  AOI22_X1 U9880 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14206), .B1(n13873), 
        .B2(n13862), .ZN(n13871) );
  NAND2_X1 U9881 ( .A1(n7627), .A2(n7626), .ZN(n9082) );
  OR2_X1 U9882 ( .A1(n12253), .A2(n7725), .ZN(n7767) );
  INV_X1 U9883 ( .A(n14666), .ZN(n12019) );
  INV_X1 U9884 ( .A(n14678), .ZN(n11977) );
  INV_X1 U9885 ( .A(n12023), .ZN(n14668) );
  OR2_X1 U9886 ( .A1(n8606), .A2(n8921), .ZN(n12037) );
  AND3_X1 U9887 ( .A1(n8811), .A2(n8810), .A3(n8809), .ZN(n12420) );
  INV_X1 U9888 ( .A(n12469), .ZN(n11980) );
  NOR2_X1 U9889 ( .A1(n7717), .A2(n10916), .ZN(n11078) );
  XNOR2_X1 U9890 ( .A(n7721), .B(n14015), .ZN(n14023) );
  AND2_X1 U9891 ( .A1(n7764), .A2(n12659), .ZN(n14703) );
  INV_X1 U9892 ( .A(n12418), .ZN(n14778) );
  OR2_X1 U9893 ( .A1(n14793), .A2(n14783), .ZN(n8986) );
  INV_X1 U9894 ( .A(n14785), .ZN(n14772) );
  INV_X1 U9895 ( .A(n12548), .ZN(n12536) );
  AND2_X1 U9896 ( .A1(n8960), .A2(n8959), .ZN(n8999) );
  AND2_X1 U9897 ( .A1(n14049), .A2(n14048), .ZN(n14056) );
  AND2_X1 U9898 ( .A1(n12060), .A2(n8977), .ZN(n12432) );
  INV_X1 U9899 ( .A(n14837), .ZN(n14821) );
  NAND2_X1 U9900 ( .A1(n8985), .A2(n8984), .ZN(n14843) );
  AND2_X1 U9901 ( .A1(n14769), .A2(n12068), .ZN(n14833) );
  XNOR2_X1 U9902 ( .A(n7629), .B(n7628), .ZN(n9081) );
  AND2_X1 U9903 ( .A1(n7637), .A2(n7724), .ZN(n14029) );
  INV_X1 U9904 ( .A(n12657), .ZN(n13948) );
  AND2_X1 U9905 ( .A1(n11589), .A2(n11588), .ZN(n12909) );
  INV_X1 U9906 ( .A(n12742), .ZN(n12758) );
  AND4_X1 U9907 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n12883) );
  AND4_X1 U9908 ( .A1(n11494), .A2(n11493), .A3(n11492), .A4(n11491), .ZN(
        n11495) );
  INV_X1 U9909 ( .A(n11590), .ZN(n11459) );
  AND2_X1 U9910 ( .A1(n13206), .A2(n9130), .ZN(n12814) );
  INV_X1 U9911 ( .A(n12815), .ZN(n14537) );
  AND2_X1 U9912 ( .A1(n9134), .A2(n13202), .ZN(n9130) );
  INV_X1 U9913 ( .A(n9339), .ZN(n12952) );
  INV_X1 U9914 ( .A(n14562), .ZN(n9585) );
  AND2_X1 U9915 ( .A1(n9154), .A2(P2_U3088), .ZN(n10909) );
  AND2_X1 U9916 ( .A1(n8241), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8252) );
  NOR2_X1 U9917 ( .A1(n10357), .A2(n10361), .ZN(n9850) );
  INV_X1 U9918 ( .A(n13608), .ZN(n15021) );
  AND4_X1 U9919 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n13607)
         );
  INV_X1 U9920 ( .A(n14284), .ZN(n14226) );
  OR2_X1 U9921 ( .A1(n10364), .A2(n8520), .ZN(n9252) );
  XNOR2_X1 U9922 ( .A(n13540), .B(n13539), .ZN(n13742) );
  INV_X1 U9923 ( .A(n14298), .ZN(n14310) );
  INV_X1 U9924 ( .A(n14397), .ZN(n14417) );
  INV_X1 U9925 ( .A(n14373), .ZN(n14379) );
  INV_X1 U9926 ( .A(n14368), .ZN(n14421) );
  NOR2_X1 U9927 ( .A1(n9852), .A2(n9649), .ZN(n9651) );
  AND2_X1 U9928 ( .A1(n9908), .A2(n9243), .ZN(n10364) );
  INV_X1 U9929 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n7935) );
  AND2_X1 U9930 ( .A1(n8126), .A2(n8143), .ZN(n9471) );
  AND2_X1 U9931 ( .A1(n7768), .A2(n7767), .ZN(n14664) );
  INV_X1 U9932 ( .A(n12400), .ZN(n12588) );
  NAND2_X1 U9933 ( .A1(n9079), .A2(n12253), .ZN(n12023) );
  INV_X1 U9934 ( .A(n12009), .ZN(n12264) );
  INV_X1 U9935 ( .A(n12420), .ZN(n12270) );
  INV_X1 U9936 ( .A(n11985), .ZN(n12273) );
  INV_X1 U9937 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14698) );
  INV_X1 U9938 ( .A(n14040), .ZN(n14708) );
  AND2_X1 U9939 ( .A1(n14787), .A2(n8986), .ZN(n12493) );
  OR2_X1 U9940 ( .A1(n14793), .A2(n14770), .ZN(n14787) );
  NAND2_X1 U9941 ( .A1(n14868), .A2(n14848), .ZN(n12540) );
  NAND2_X1 U9942 ( .A1(n14868), .A2(n14821), .ZN(n12548) );
  AND2_X2 U9943 ( .A1(n8999), .A2(n8998), .ZN(n14868) );
  INV_X1 U9944 ( .A(n12427), .ZN(n12600) );
  INV_X1 U9945 ( .A(n14851), .ZN(n14849) );
  AND2_X2 U9946 ( .A1(n9010), .A2(n12253), .ZN(n14851) );
  NAND2_X1 U9947 ( .A1(n8946), .A2(n12636), .ZN(n9262) );
  XNOR2_X1 U9948 ( .A(n7624), .B(n7623), .ZN(n11098) );
  INV_X1 U9949 ( .A(SI_19_), .ZN(n9759) );
  INV_X1 U9950 ( .A(SI_13_), .ZN(n9223) );
  INV_X1 U9951 ( .A(n13948), .ZN(n12664) );
  INV_X1 U9952 ( .A(n13126), .ZN(n12998) );
  INV_X1 U9953 ( .A(n12747), .ZN(n12761) );
  OR2_X1 U9954 ( .A1(n9329), .A2(n9328), .ZN(n12749) );
  INV_X1 U9955 ( .A(n12883), .ZN(n12769) );
  INV_X1 U9956 ( .A(n11495), .ZN(n12874) );
  INV_X1 U9957 ( .A(n14442), .ZN(n14540) );
  OR2_X1 U9958 ( .A1(n9586), .A2(n14562), .ZN(n14661) );
  AND3_X1 U9959 ( .A1(n14635), .A2(n14634), .A3(n14633), .ZN(n14660) );
  OR2_X1 U9960 ( .A1(n9586), .A2(n9585), .ZN(n14646) );
  NOR2_X1 U9961 ( .A1(n14563), .A2(n14558), .ZN(n14559) );
  INV_X1 U9962 ( .A(n14559), .ZN(n14560) );
  INV_X1 U9963 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14963) );
  INV_X1 U9964 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11487) );
  INV_X1 U9965 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9721) );
  INV_X1 U9966 ( .A(n13750), .ZN(n13582) );
  INV_X1 U9967 ( .A(n13763), .ZN(n13534) );
  INV_X1 U9968 ( .A(n14075), .ZN(n13329) );
  NAND2_X1 U9969 ( .A1(n9850), .A2(n9849), .ZN(n14078) );
  OAI21_X1 U9970 ( .B1(n13669), .B2(n8298), .A(n8350), .ZN(n13678) );
  INV_X1 U9971 ( .A(n10974), .ZN(n13346) );
  NAND2_X1 U9972 ( .A1(n9423), .A2(n8530), .ZN(n14284) );
  INV_X1 U9973 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14916) );
  NAND2_X1 U9974 ( .A1(n9252), .A2(n9250), .ZN(n14288) );
  INV_X1 U9975 ( .A(n13977), .ZN(n13705) );
  NAND2_X1 U9976 ( .A1(n10364), .A2(n10363), .ZN(n14093) );
  INV_X1 U9977 ( .A(n14308), .ZN(n13675) );
  INV_X2 U9978 ( .A(n14438), .ZN(n14441) );
  AND3_X1 U9979 ( .A1(n14142), .A2(n14141), .A3(n14140), .ZN(n14167) );
  INV_X1 U9980 ( .A(n14425), .ZN(n14423) );
  AND2_X2 U9981 ( .A1(n9566), .A2(n10364), .ZN(n14350) );
  AND2_X2 U9982 ( .A1(n7630), .A2(n12636), .ZN(P3_U3897) );
  OR4_X1 U9983 ( .A1(n9102), .A2(n9101), .A3(n9100), .A4(n9099), .ZN(P3_U3171)
         );
  NOR2_X1 U9984 ( .A1(n9125), .A2(P2_U3088), .ZN(P2_U3947) );
  NAND4_X1 U9985 ( .A1(n7610), .A2(n7700), .A3(n7662), .A4(n7609), .ZN(n7651)
         );
  NAND4_X1 U9986 ( .A1(n7656), .A2(n7660), .A3(n7650), .A4(n7611), .ZN(n7612)
         );
  INV_X1 U9987 ( .A(n11282), .ZN(n7627) );
  NOR2_X1 U9988 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7621) );
  OR2_X1 U9989 ( .A1(n7622), .A2(n7646), .ZN(n7624) );
  INV_X1 U9990 ( .A(n11098), .ZN(n7625) );
  INV_X1 U9991 ( .A(n9082), .ZN(n7630) );
  NAND2_X1 U9992 ( .A1(n6505), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9993 ( .A1(n7638), .A2(n7632), .ZN(n7634) );
  NAND2_X1 U9994 ( .A1(n7634), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7633) );
  MUX2_X1 U9995 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7633), .S(
        P3_IR_REG_18__SCAN_IN), .Z(n7637) );
  INV_X1 U9996 ( .A(n7634), .ZN(n7636) );
  NAND2_X1 U9997 ( .A1(n7636), .A2(n7635), .ZN(n7724) );
  OR2_X1 U9998 ( .A1(n7638), .A2(n7646), .ZN(n7639) );
  XNOR2_X1 U9999 ( .A(n7639), .B(P3_IR_REG_17__SCAN_IN), .ZN(n14015) );
  NAND2_X1 U10000 ( .A1(n7642), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7640) );
  XNOR2_X1 U10001 ( .A(n7640), .B(P3_IR_REG_16__SCAN_IN), .ZN(n13998) );
  INV_X1 U10002 ( .A(n13998), .ZN(n9388) );
  NAND2_X1 U10003 ( .A1(n7631), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7641) );
  MUX2_X1 U10004 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7641), .S(
        P3_IR_REG_15__SCAN_IN), .Z(n7643) );
  NAND2_X1 U10005 ( .A1(n7643), .A2(n7642), .ZN(n9259) );
  NOR2_X1 U10006 ( .A1(n7644), .A2(n7646), .ZN(n7645) );
  MUX2_X1 U10007 ( .A(n7646), .B(n7645), .S(P3_IR_REG_14__SCAN_IN), .Z(n7648)
         );
  INV_X1 U10008 ( .A(n7631), .ZN(n7647) );
  NAND2_X1 U10009 ( .A1(n11084), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7824) );
  NAND2_X1 U10010 ( .A1(n7649), .A2(n7650), .ZN(n7688) );
  OR2_X1 U10011 ( .A1(n7688), .A2(n7651), .ZN(n7664) );
  NOR2_X1 U10012 ( .A1(n7664), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n7655) );
  NAND2_X1 U10013 ( .A1(n7655), .A2(n7656), .ZN(n7658) );
  NAND2_X1 U10014 ( .A1(n7658), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7652) );
  MUX2_X1 U10015 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7652), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7654) );
  INV_X1 U10016 ( .A(n7644), .ZN(n7653) );
  NAND2_X1 U10017 ( .A1(n7654), .A2(n7653), .ZN(n10922) );
  INV_X1 U10018 ( .A(n10922), .ZN(n8734) );
  OR2_X1 U10019 ( .A1(n7655), .A2(n7646), .ZN(n7657) );
  MUX2_X1 U10020 ( .A(n7657), .B(P3_IR_REG_31__SCAN_IN), .S(n7656), .Z(n7659)
         );
  NAND2_X1 U10021 ( .A1(n7664), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7661) );
  XNOR2_X1 U10022 ( .A(n7661), .B(n7660), .ZN(n9174) );
  INV_X1 U10023 ( .A(n9174), .ZN(n10682) );
  NAND2_X1 U10024 ( .A1(n7705), .A2(n7662), .ZN(n7707) );
  NAND2_X1 U10025 ( .A1(n7707), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7663) );
  MUX2_X1 U10026 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7663), .S(
        P3_IR_REG_10__SCAN_IN), .Z(n7665) );
  NAND2_X1 U10027 ( .A1(n7688), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7667) );
  INV_X1 U10028 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7666) );
  XNOR2_X1 U10029 ( .A(n7667), .B(n7666), .ZN(n9931) );
  INV_X1 U10030 ( .A(n9931), .ZN(n7797) );
  INV_X1 U10031 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n7692) );
  INV_X1 U10032 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n14774) );
  NOR2_X1 U10033 ( .A1(n7668), .A2(n7646), .ZN(n7669) );
  MUX2_X1 U10034 ( .A(n7646), .B(n7669), .S(P3_IR_REG_2__SCAN_IN), .Z(n7672)
         );
  INV_X1 U10035 ( .A(n7670), .ZN(n7671) );
  NAND2_X1 U10036 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n7673) );
  MUX2_X1 U10037 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7673), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n7675) );
  INV_X1 U10038 ( .A(n7668), .ZN(n7674) );
  INV_X1 U10039 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10022) );
  NOR2_X1 U10040 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10022), .ZN(n9675) );
  NAND2_X1 U10041 ( .A1(n7668), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7676) );
  OAI21_X1 U10042 ( .B1(n9752), .B2(n9675), .A(n7676), .ZN(n9742) );
  INV_X1 U10043 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n14790) );
  OR2_X1 U10044 ( .A1(n9742), .A2(n14790), .ZN(n9744) );
  OR2_X1 U10045 ( .A1(n9216), .A2(n14774), .ZN(n7677) );
  NAND2_X1 U10046 ( .A1(n7670), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7678) );
  MUX2_X1 U10047 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7678), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n7680) );
  AND2_X1 U10048 ( .A1(n7680), .A2(n7679), .ZN(n9667) );
  INV_X1 U10049 ( .A(n9667), .ZN(n9207) );
  NAND2_X1 U10050 ( .A1(n7681), .A2(n9207), .ZN(n9769) );
  NAND2_X1 U10051 ( .A1(n9769), .A2(n7682), .ZN(n9658) );
  INV_X1 U10052 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U10053 ( .A1(n9771), .A2(n9769), .ZN(n7684) );
  NAND2_X1 U10054 ( .A1(n7679), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7683) );
  XNOR2_X1 U10055 ( .A(n9776), .B(P3_REG2_REG_4__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U10056 ( .A1(n7684), .A2(n9768), .ZN(n9773) );
  INV_X1 U10057 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n7685) );
  OR2_X1 U10058 ( .A1(n9776), .A2(n7685), .ZN(n7686) );
  NAND2_X1 U10059 ( .A1(n9773), .A2(n7686), .ZN(n7691) );
  NOR2_X1 U10060 ( .A1(n7649), .A2(n7646), .ZN(n7687) );
  MUX2_X1 U10061 ( .A(n7646), .B(n7687), .S(P3_IR_REG_5__SCAN_IN), .Z(n7690)
         );
  INV_X1 U10062 ( .A(n7688), .ZN(n7689) );
  NAND2_X1 U10063 ( .A1(n7691), .A2(n9788), .ZN(n9923) );
  INV_X1 U10064 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9782) );
  MUX2_X1 U10065 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n7692), .S(n9931), .Z(n9922)
         );
  NAND2_X1 U10066 ( .A1(n7693), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7694) );
  XNOR2_X1 U10067 ( .A(n7694), .B(P3_IR_REG_7__SCAN_IN), .ZN(n8667) );
  INV_X1 U10068 ( .A(n8667), .ZN(n9964) );
  NAND2_X1 U10069 ( .A1(n7695), .A2(n9964), .ZN(n7697) );
  INV_X1 U10070 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n10830) );
  INV_X1 U10071 ( .A(n7697), .ZN(n7698) );
  NAND2_X1 U10072 ( .A1(n7699), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7701) );
  MUX2_X1 U10073 ( .A(n7701), .B(P3_IR_REG_31__SCAN_IN), .S(n7700), .Z(n7703)
         );
  INV_X1 U10074 ( .A(n7705), .ZN(n7702) );
  NAND2_X1 U10075 ( .A1(n7703), .A2(n7702), .ZN(n10034) );
  INV_X1 U10076 ( .A(n10034), .ZN(n7806) );
  INV_X1 U10077 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n7704) );
  AOI22_X1 U10078 ( .A1(n7806), .A2(P3_REG2_REG_8__SCAN_IN), .B1(n7704), .B2(
        n10034), .ZN(n10032) );
  NOR2_X1 U10079 ( .A1(n7705), .A2(n7646), .ZN(n7706) );
  MUX2_X1 U10080 ( .A(n7646), .B(n7706), .S(P3_IR_REG_9__SCAN_IN), .Z(n7709)
         );
  INV_X1 U10081 ( .A(n7707), .ZN(n7708) );
  NAND2_X1 U10082 ( .A1(n7711), .A2(n9178), .ZN(n7710) );
  INV_X1 U10083 ( .A(n7710), .ZN(n7712) );
  INV_X1 U10084 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n14976) );
  NOR2_X1 U10085 ( .A1(n14976), .A2(n14681), .ZN(n14680) );
  NOR2_X1 U10086 ( .A1(n7712), .A2(n14680), .ZN(n14707) );
  INV_X1 U10087 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n7713) );
  AOI22_X1 U10088 ( .A1(n8701), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n7713), .B2(
        n14718), .ZN(n14706) );
  NOR2_X1 U10089 ( .A1(n14707), .A2(n14706), .ZN(n14705) );
  AOI21_X1 U10090 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14718), .A(n14705), 
        .ZN(n7714) );
  INV_X1 U10091 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11057) );
  XOR2_X1 U10092 ( .A(n9174), .B(n7714), .Z(n10675) );
  INV_X1 U10093 ( .A(n10633), .ZN(n7819) );
  INV_X1 U10094 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n7715) );
  AOI22_X1 U10095 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n7819), .B1(n10633), 
        .B2(n7715), .ZN(n10625) );
  NOR2_X1 U10096 ( .A1(n8734), .A2(n7716), .ZN(n7717) );
  INV_X1 U10097 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n14910) );
  NOR2_X1 U10098 ( .A1(n14910), .A2(n10917), .ZN(n10916) );
  OAI21_X1 U10099 ( .B1(n11084), .B2(P3_REG2_REG_14__SCAN_IN), .A(n7824), .ZN(
        n11077) );
  NOR2_X1 U10100 ( .A1(n11078), .A2(n11077), .ZN(n11076) );
  INV_X1 U10101 ( .A(n11076), .ZN(n7718) );
  AND2_X1 U10102 ( .A1(n9259), .A2(n7719), .ZN(n7720) );
  INV_X1 U10103 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12459) );
  INV_X1 U10104 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U10105 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n13998), .B1(n9388), 
        .B2(n12447), .ZN(n14009) );
  NOR2_X1 U10106 ( .A1(n14015), .A2(n7721), .ZN(n7722) );
  INV_X1 U10107 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14931) );
  INV_X1 U10108 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n7723) );
  AOI22_X1 U10109 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n14029), .B1(n13951), 
        .B2(n7723), .ZN(n14041) );
  XNOR2_X1 U10110 ( .A(n12055), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n7773) );
  OR2_X1 U10111 ( .A1(n9081), .A2(P3_U3151), .ZN(n12259) );
  INV_X1 U10112 ( .A(n12259), .ZN(n7725) );
  NAND2_X1 U10113 ( .A1(n7728), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7727) );
  NAND2_X4 U10114 ( .A1(n12654), .A2(n7737), .ZN(n8934) );
  NAND2_X1 U10115 ( .A1(n7732), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7733) );
  MUX2_X1 U10116 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7733), .S(
        P3_IR_REG_22__SCAN_IN), .Z(n7734) );
  NAND2_X1 U10117 ( .A1(n6484), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7735) );
  NAND2_X1 U10118 ( .A1(n12256), .A2(n9041), .ZN(n12183) );
  NAND2_X1 U10119 ( .A1(n12076), .A2(n9081), .ZN(n7736) );
  AND2_X1 U10120 ( .A1(n8934), .A2(n7736), .ZN(n7766) );
  AND2_X1 U10121 ( .A1(n7767), .A2(n7766), .ZN(n7764) );
  OR2_X1 U10122 ( .A1(n12654), .A2(n12659), .ZN(n8935) );
  INV_X1 U10123 ( .A(n8935), .ZN(n7738) );
  NAND2_X1 U10124 ( .A1(n7739), .A2(n14040), .ZN(n7836) );
  INV_X1 U10125 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U10126 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n13951), .B1(n14029), 
        .B2(n12527), .ZN(n14032) );
  INV_X1 U10127 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U10128 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n9388), .B1(n13998), 
        .B2(n12532), .ZN(n14006) );
  NAND2_X1 U10129 ( .A1(n11084), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7823) );
  INV_X1 U10130 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n7756) );
  AOI22_X1 U10131 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n10633), .B1(n7819), 
        .B2(n7756), .ZN(n10629) );
  INV_X1 U10132 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n14944) );
  AOI22_X1 U10133 ( .A1(n8701), .A2(n14944), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n14718), .ZN(n14701) );
  NAND2_X1 U10134 ( .A1(n10034), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7751) );
  INV_X1 U10135 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n14862) );
  AOI22_X1 U10136 ( .A1(n7806), .A2(n14862), .B1(P3_REG1_REG_8__SCAN_IN), .B2(
        n10034), .ZN(n10029) );
  INV_X1 U10137 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n14859) );
  INV_X1 U10138 ( .A(n9776), .ZN(n9210) );
  INV_X1 U10139 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n7740) );
  INV_X1 U10140 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U10141 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n7741), .ZN(n9672) );
  INV_X1 U10142 ( .A(n9672), .ZN(n7743) );
  OR2_X1 U10143 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n9672), .ZN(n7742) );
  OAI21_X1 U10144 ( .B1(n9752), .B2(n7743), .A(n7742), .ZN(n9746) );
  INV_X1 U10145 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n9745) );
  OR2_X1 U10146 ( .A1(n9746), .A2(n9745), .ZN(n9748) );
  OAI21_X1 U10147 ( .B1(P3_IR_REG_1__SCAN_IN), .B2(n9672), .A(n9748), .ZN(
        n9729) );
  NAND2_X1 U10148 ( .A1(n9730), .A2(n9729), .ZN(n9728) );
  OR2_X1 U10149 ( .A1(n9216), .A2(n7740), .ZN(n7744) );
  NAND2_X1 U10150 ( .A1(n9728), .A2(n7744), .ZN(n7745) );
  INV_X1 U10151 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n14856) );
  MUX2_X1 U10152 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n14856), .S(n9776), .Z(n9764) );
  NOR2_X1 U10153 ( .A1(n9763), .A2(n9764), .ZN(n9762) );
  XNOR2_X1 U10154 ( .A(n7746), .B(n7090), .ZN(n9781) );
  INV_X1 U10155 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n7747) );
  OAI22_X1 U10156 ( .A1(n9781), .A2(n7747), .B1(n7090), .B2(n7746), .ZN(n9920)
         );
  MUX2_X1 U10157 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n14859), .S(n9931), .Z(n9921) );
  NAND2_X1 U10158 ( .A1(n9920), .A2(n9921), .ZN(n9919) );
  OAI21_X1 U10159 ( .B1(n7797), .B2(n14859), .A(n9919), .ZN(n7748) );
  INV_X1 U10160 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n7750) );
  INV_X1 U10161 ( .A(n7748), .ZN(n7749) );
  NAND2_X1 U10162 ( .A1(n9178), .A2(n7752), .ZN(n7753) );
  NAND2_X1 U10163 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n14683), .ZN(n14682) );
  NAND2_X1 U10164 ( .A1(n7753), .A2(n14682), .ZN(n14700) );
  NAND2_X1 U10165 ( .A1(n14701), .A2(n14700), .ZN(n14699) );
  NAND2_X1 U10166 ( .A1(n9174), .A2(n7754), .ZN(n7755) );
  XNOR2_X1 U10167 ( .A(n7754), .B(n10682), .ZN(n10684) );
  NAND2_X1 U10168 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n10684), .ZN(n10683) );
  NAND2_X1 U10169 ( .A1(n10922), .A2(n7757), .ZN(n7758) );
  XNOR2_X1 U10170 ( .A(n8734), .B(n7757), .ZN(n10919) );
  NAND2_X1 U10171 ( .A1(P3_REG1_REG_13__SCAN_IN), .A2(n10919), .ZN(n10918) );
  OAI21_X1 U10172 ( .B1(n11084), .B2(P3_REG1_REG_14__SCAN_IN), .A(n7823), .ZN(
        n7822) );
  INV_X1 U10173 ( .A(n7822), .ZN(n11081) );
  NAND2_X1 U10174 ( .A1(n11080), .A2(n11081), .ZN(n11079) );
  NAND2_X1 U10175 ( .A1(n9259), .A2(n7759), .ZN(n7760) );
  NAND2_X1 U10176 ( .A1(P3_REG1_REG_15__SCAN_IN), .A2(n12285), .ZN(n12284) );
  NAND2_X1 U10177 ( .A1(n7760), .A2(n12284), .ZN(n14005) );
  NAND2_X1 U10178 ( .A1(n9591), .A2(n7761), .ZN(n7762) );
  XNOR2_X1 U10179 ( .A(n14015), .B(n7761), .ZN(n14017) );
  NAND2_X1 U10180 ( .A1(n14032), .A2(n14031), .ZN(n14030) );
  XNOR2_X1 U10181 ( .A(n12055), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n7772) );
  INV_X1 U10182 ( .A(n7772), .ZN(n7763) );
  INV_X1 U10183 ( .A(P3_U3897), .ZN(n12280) );
  INV_X1 U10184 ( .A(n7764), .ZN(n7765) );
  MUX2_X1 U10185 ( .A(n12280), .B(n7765), .S(n12654), .Z(n14719) );
  NAND2_X1 U10186 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n11913)
         );
  INV_X1 U10187 ( .A(n7766), .ZN(n7768) );
  NAND2_X1 U10188 ( .A1(n14664), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7769) );
  OAI211_X1 U10189 ( .C1(n14719), .C2(n12055), .A(n11913), .B(n7769), .ZN(
        n7770) );
  AOI21_X1 U10190 ( .B1(n7771), .B2(n14703), .A(n7770), .ZN(n7835) );
  MUX2_X1 U10191 ( .A(n7773), .B(n7772), .S(n12659), .Z(n7832) );
  MUX2_X1 U10192 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12659), .Z(n7829) );
  INV_X1 U10193 ( .A(n9752), .ZN(n7776) );
  XNOR2_X1 U10194 ( .A(n7775), .B(n7776), .ZN(n9741) );
  INV_X1 U10195 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n7774) );
  MUX2_X1 U10196 ( .A(n10022), .B(n7774), .S(n12659), .Z(n9676) );
  AND2_X1 U10197 ( .A1(n9676), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n9670) );
  NAND2_X1 U10198 ( .A1(n9741), .A2(n9670), .ZN(n7779) );
  INV_X1 U10199 ( .A(n7775), .ZN(n7777) );
  NAND2_X1 U10200 ( .A1(n7777), .A2(n7776), .ZN(n7778) );
  NAND2_X1 U10201 ( .A1(n7779), .A2(n7778), .ZN(n9723) );
  MUX2_X1 U10202 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12659), .Z(n7780) );
  XNOR2_X1 U10203 ( .A(n7780), .B(n9216), .ZN(n9724) );
  NAND2_X1 U10204 ( .A1(n9723), .A2(n9724), .ZN(n7783) );
  INV_X1 U10205 ( .A(n7780), .ZN(n7781) );
  NAND2_X1 U10206 ( .A1(n7781), .A2(n9216), .ZN(n7782) );
  NAND2_X1 U10207 ( .A1(n7783), .A2(n7782), .ZN(n9656) );
  MUX2_X1 U10208 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12659), .Z(n7784) );
  XNOR2_X1 U10209 ( .A(n7784), .B(n9667), .ZN(n9657) );
  NAND2_X1 U10210 ( .A1(n9656), .A2(n9657), .ZN(n7787) );
  INV_X1 U10211 ( .A(n7784), .ZN(n7785) );
  NAND2_X1 U10212 ( .A1(n7785), .A2(n9667), .ZN(n7786) );
  NAND2_X1 U10213 ( .A1(n7787), .A2(n7786), .ZN(n9760) );
  MUX2_X1 U10214 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12659), .Z(n7788) );
  XNOR2_X1 U10215 ( .A(n7788), .B(n9776), .ZN(n9761) );
  NAND2_X1 U10216 ( .A1(n9760), .A2(n9761), .ZN(n7791) );
  INV_X1 U10217 ( .A(n7788), .ZN(n7789) );
  NAND2_X1 U10218 ( .A1(n7789), .A2(n9776), .ZN(n7790) );
  NAND2_X1 U10219 ( .A1(n7791), .A2(n7790), .ZN(n9779) );
  MUX2_X1 U10220 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12659), .Z(n7792) );
  XNOR2_X1 U10221 ( .A(n7792), .B(n7090), .ZN(n9780) );
  NAND2_X1 U10222 ( .A1(n9779), .A2(n9780), .ZN(n7795) );
  INV_X1 U10223 ( .A(n7792), .ZN(n7793) );
  NAND2_X1 U10224 ( .A1(n7793), .A2(n7090), .ZN(n7794) );
  NAND2_X1 U10225 ( .A1(n7795), .A2(n7794), .ZN(n9917) );
  MUX2_X1 U10226 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12659), .Z(n7796) );
  XNOR2_X1 U10227 ( .A(n7796), .B(n7797), .ZN(n9918) );
  NAND2_X1 U10228 ( .A1(n9917), .A2(n9918), .ZN(n7800) );
  INV_X1 U10229 ( .A(n7796), .ZN(n7798) );
  NAND2_X1 U10230 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  NAND2_X1 U10231 ( .A1(n7800), .A2(n7799), .ZN(n9957) );
  MUX2_X1 U10232 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12659), .Z(n7801) );
  XNOR2_X1 U10233 ( .A(n7801), .B(n8667), .ZN(n9958) );
  NAND2_X1 U10234 ( .A1(n9957), .A2(n9958), .ZN(n7804) );
  INV_X1 U10235 ( .A(n7801), .ZN(n7802) );
  NAND2_X1 U10236 ( .A1(n7802), .A2(n8667), .ZN(n7803) );
  NAND2_X1 U10237 ( .A1(n7804), .A2(n7803), .ZN(n10026) );
  MUX2_X1 U10238 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12659), .Z(n7805) );
  XNOR2_X1 U10239 ( .A(n7805), .B(n7806), .ZN(n10027) );
  NAND2_X1 U10240 ( .A1(n10026), .A2(n10027), .ZN(n7809) );
  INV_X1 U10241 ( .A(n7805), .ZN(n7807) );
  NAND2_X1 U10242 ( .A1(n7807), .A2(n7806), .ZN(n7808) );
  NAND2_X1 U10243 ( .A1(n7809), .A2(n7808), .ZN(n14688) );
  MUX2_X1 U10244 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12659), .Z(n7810) );
  NAND2_X1 U10245 ( .A1(n7810), .A2(n9178), .ZN(n14687) );
  NAND2_X1 U10246 ( .A1(n14688), .A2(n14687), .ZN(n14712) );
  INV_X1 U10247 ( .A(n7810), .ZN(n7811) );
  NAND2_X1 U10248 ( .A1(n7811), .A2(n14685), .ZN(n14711) );
  MUX2_X1 U10249 ( .A(n7713), .B(n14944), .S(n12659), .Z(n7812) );
  NAND2_X1 U10250 ( .A1(n7812), .A2(n8701), .ZN(n7815) );
  INV_X1 U10251 ( .A(n7812), .ZN(n7813) );
  NAND2_X1 U10252 ( .A1(n7813), .A2(n14718), .ZN(n7814) );
  NAND2_X1 U10253 ( .A1(n7815), .A2(n7814), .ZN(n14710) );
  INV_X1 U10254 ( .A(n7815), .ZN(n7816) );
  NOR2_X1 U10255 ( .A1(n14715), .A2(n7816), .ZN(n10678) );
  MUX2_X1 U10256 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12659), .Z(n7817) );
  XNOR2_X1 U10257 ( .A(n7817), .B(n9174), .ZN(n10677) );
  NOR2_X1 U10258 ( .A1(n7817), .A2(n9174), .ZN(n10637) );
  MUX2_X1 U10259 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12659), .Z(n7818) );
  XNOR2_X1 U10260 ( .A(n7818), .B(n10633), .ZN(n10636) );
  NOR3_X1 U10261 ( .A1(n10676), .A2(n10637), .A3(n10636), .ZN(n10925) );
  INV_X1 U10262 ( .A(n7818), .ZN(n7820) );
  NOR2_X1 U10263 ( .A1(n7820), .A2(n7819), .ZN(n10924) );
  MUX2_X1 U10264 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12659), .Z(n7821) );
  XNOR2_X1 U10265 ( .A(n7821), .B(n10922), .ZN(n10923) );
  NOR2_X1 U10266 ( .A1(n7821), .A2(n10922), .ZN(n11086) );
  MUX2_X1 U10267 ( .A(n11077), .B(n7822), .S(n12659), .Z(n11085) );
  MUX2_X1 U10268 ( .A(n7824), .B(n7823), .S(n12659), .Z(n7825) );
  NAND2_X1 U10269 ( .A1(n11088), .A2(n7825), .ZN(n7826) );
  INV_X1 U10270 ( .A(n7826), .ZN(n7827) );
  INV_X1 U10271 ( .A(n9259), .ZN(n12292) );
  XNOR2_X1 U10272 ( .A(n7826), .B(n9259), .ZN(n12288) );
  MUX2_X1 U10273 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12659), .Z(n12287) );
  NOR2_X1 U10274 ( .A1(n12288), .A2(n12287), .ZN(n12286) );
  AOI21_X1 U10275 ( .B1(n7827), .B2(n12292), .A(n12286), .ZN(n14003) );
  MUX2_X1 U10276 ( .A(n12447), .B(n12532), .S(n12659), .Z(n7828) );
  NOR2_X1 U10277 ( .A1(n7828), .A2(n13998), .ZN(n13999) );
  NAND2_X1 U10278 ( .A1(n7828), .A2(n13998), .ZN(n14000) );
  XNOR2_X1 U10279 ( .A(n7829), .B(n9591), .ZN(n14020) );
  NOR2_X1 U10280 ( .A1(n14019), .A2(n14020), .ZN(n14018) );
  AOI21_X1 U10281 ( .B1(n7829), .B2(n9591), .A(n14018), .ZN(n7830) );
  XNOR2_X1 U10282 ( .A(n7830), .B(n14029), .ZN(n14034) );
  MUX2_X1 U10283 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n12659), .Z(n14035) );
  NOR2_X1 U10284 ( .A1(n14034), .A2(n14035), .ZN(n14033) );
  XOR2_X1 U10285 ( .A(n7832), .B(n7831), .Z(n7833) );
  NAND2_X1 U10286 ( .A1(P3_U3897), .A2(n12654), .ZN(n14036) );
  INV_X1 U10287 ( .A(SI_1_), .ZN(n9173) );
  MUX2_X1 U10288 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(P1_DATAO_REG_0__SCAN_IN), 
        .S(n7847), .Z(n7840) );
  NAND2_X1 U10289 ( .A1(n7841), .A2(SI_2_), .ZN(n7843) );
  OAI21_X1 U10290 ( .B1(n7841), .B2(SI_2_), .A(n7843), .ZN(n7993) );
  INV_X1 U10291 ( .A(n7993), .ZN(n7842) );
  MUX2_X1 U10292 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n7847), .Z(n7844) );
  NAND2_X1 U10293 ( .A1(n7844), .A2(SI_3_), .ZN(n7846) );
  OAI21_X1 U10294 ( .B1(n7844), .B2(SI_3_), .A(n7846), .ZN(n8004) );
  INV_X1 U10295 ( .A(n8004), .ZN(n7845) );
  MUX2_X1 U10296 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n7847), .Z(n7848) );
  NAND2_X1 U10297 ( .A1(n7848), .A2(SI_4_), .ZN(n7850) );
  OAI21_X1 U10298 ( .B1(n7848), .B2(SI_4_), .A(n7850), .ZN(n8032) );
  INV_X1 U10299 ( .A(n8032), .ZN(n7849) );
  MUX2_X1 U10300 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n7847), .Z(n7851) );
  NAND2_X1 U10301 ( .A1(n7851), .A2(SI_5_), .ZN(n7853) );
  OAI21_X1 U10302 ( .B1(n7851), .B2(SI_5_), .A(n7853), .ZN(n8042) );
  INV_X1 U10303 ( .A(n8042), .ZN(n7852) );
  NAND2_X1 U10304 ( .A1(n7854), .A2(SI_6_), .ZN(n7856) );
  OAI21_X1 U10305 ( .B1(n7854), .B2(SI_6_), .A(n7856), .ZN(n8067) );
  INV_X1 U10306 ( .A(n8067), .ZN(n7855) );
  MUX2_X1 U10307 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9154), .Z(n7858) );
  NAND2_X1 U10308 ( .A1(n7858), .A2(SI_7_), .ZN(n7860) );
  OAI21_X1 U10309 ( .B1(n7858), .B2(SI_7_), .A(n7860), .ZN(n7859) );
  INV_X1 U10310 ( .A(n7859), .ZN(n8089) );
  MUX2_X1 U10311 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9154), .Z(n7861) );
  NAND2_X1 U10312 ( .A1(n7861), .A2(SI_8_), .ZN(n7863) );
  OAI21_X1 U10313 ( .B1(n7861), .B2(SI_8_), .A(n7863), .ZN(n7862) );
  INV_X1 U10314 ( .A(n7862), .ZN(n8074) );
  MUX2_X1 U10315 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9154), .Z(n7864) );
  NAND2_X1 U10316 ( .A1(n7864), .A2(SI_9_), .ZN(n7866) );
  OAI21_X1 U10317 ( .B1(n7864), .B2(SI_9_), .A(n7866), .ZN(n7865) );
  INV_X1 U10318 ( .A(n7865), .ZN(n8121) );
  MUX2_X1 U10319 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9154), .Z(n8140) );
  NOR2_X1 U10320 ( .A1(n7867), .A2(n9203), .ZN(n7868) );
  MUX2_X1 U10321 ( .A(n8563), .B(n9267), .S(n9154), .Z(n7869) );
  XNOR2_X1 U10322 ( .A(n7869), .B(SI_11_), .ZN(n8159) );
  INV_X1 U10323 ( .A(SI_11_), .ZN(n9175) );
  NAND2_X1 U10324 ( .A1(n7869), .A2(n9175), .ZN(n7870) );
  MUX2_X1 U10325 ( .A(n8564), .B(n9395), .S(n9154), .Z(n7871) );
  NAND2_X1 U10326 ( .A1(n8177), .A2(n8176), .ZN(n7873) );
  NAND2_X1 U10327 ( .A1(n7871), .A2(n9198), .ZN(n7872) );
  NAND2_X1 U10328 ( .A1(n7874), .A2(n9223), .ZN(n7875) );
  INV_X1 U10329 ( .A(n8225), .ZN(n7877) );
  NAND2_X1 U10330 ( .A1(n7877), .A2(SI_15_), .ZN(n7878) );
  NOR2_X1 U10331 ( .A1(n8223), .A2(SI_14_), .ZN(n7879) );
  AOI22_X1 U10332 ( .A1(n7879), .A2(n7878), .B1(n8225), .B2(n9260), .ZN(n7880)
         );
  MUX2_X1 U10333 ( .A(n6919), .B(n11169), .S(n9154), .Z(n7882) );
  XNOR2_X1 U10334 ( .A(n7882), .B(SI_16_), .ZN(n8246) );
  MUX2_X1 U10335 ( .A(n7326), .B(n10113), .S(n9154), .Z(n7887) );
  INV_X1 U10336 ( .A(n7887), .ZN(n7888) );
  NAND2_X1 U10337 ( .A1(n7888), .A2(SI_19_), .ZN(n7889) );
  NAND2_X1 U10338 ( .A1(n7890), .A2(n7889), .ZN(n8291) );
  INV_X1 U10339 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10493) );
  MUX2_X1 U10340 ( .A(n10493), .B(n11449), .S(n9154), .Z(n8338) );
  INV_X1 U10341 ( .A(n8338), .ZN(n8351) );
  MUX2_X1 U10342 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9154), .Z(n8356) );
  NOR2_X1 U10343 ( .A1(n8338), .A2(n10110), .ZN(n7891) );
  AOI22_X1 U10344 ( .A1(n7891), .A2(n7606), .B1(n8356), .B2(SI_21_), .ZN(n7892) );
  MUX2_X1 U10345 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n9154), .Z(n11277) );
  NAND2_X1 U10346 ( .A1(n7894), .A2(SI_22_), .ZN(n7895) );
  MUX2_X1 U10347 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9154), .Z(n7897) );
  NAND2_X1 U10348 ( .A1(n7898), .A2(n7897), .ZN(n7899) );
  MUX2_X1 U10349 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n9154), .Z(n8396) );
  NAND2_X1 U10350 ( .A1(n7900), .A2(SI_24_), .ZN(n7901) );
  INV_X1 U10351 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13211) );
  MUX2_X1 U10352 ( .A(n11276), .B(n13211), .S(n9154), .Z(n7902) );
  INV_X1 U10353 ( .A(SI_25_), .ZN(n11097) );
  NAND2_X1 U10354 ( .A1(n7902), .A2(n11097), .ZN(n7905) );
  INV_X1 U10355 ( .A(n7902), .ZN(n7903) );
  NAND2_X1 U10356 ( .A1(n7903), .A2(SI_25_), .ZN(n7904) );
  NAND2_X1 U10357 ( .A1(n7905), .A2(n7904), .ZN(n8412) );
  MUX2_X1 U10358 ( .A(n13834), .B(n6922), .S(n9154), .Z(n8425) );
  MUX2_X1 U10359 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9154), .Z(n8444) );
  NOR2_X1 U10360 ( .A1(n8444), .A2(SI_27_), .ZN(n7906) );
  INV_X1 U10361 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n13830) );
  INV_X1 U10362 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11552) );
  MUX2_X1 U10363 ( .A(n13830), .B(n11552), .S(n9154), .Z(n7907) );
  INV_X1 U10364 ( .A(SI_28_), .ZN(n12653) );
  NAND2_X1 U10365 ( .A1(n7907), .A2(n12653), .ZN(n7910) );
  INV_X1 U10366 ( .A(n7907), .ZN(n7908) );
  NAND2_X1 U10367 ( .A1(n7908), .A2(SI_28_), .ZN(n7909) );
  NAND2_X1 U10368 ( .A1(n7910), .A2(n7909), .ZN(n8458) );
  INV_X1 U10369 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13825) );
  MUX2_X1 U10370 ( .A(n13825), .B(n14963), .S(n9154), .Z(n7911) );
  XNOR2_X1 U10371 ( .A(n7911), .B(SI_29_), .ZN(n7969) );
  INV_X1 U10372 ( .A(SI_29_), .ZN(n12650) );
  NAND2_X1 U10373 ( .A1(n7911), .A2(n12650), .ZN(n7912) );
  MUX2_X1 U10374 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9154), .Z(n7914) );
  NAND2_X1 U10375 ( .A1(n7914), .A2(SI_30_), .ZN(n7915) );
  OAI21_X1 U10376 ( .B1(n7914), .B2(SI_30_), .A(n7915), .ZN(n8469) );
  MUX2_X1 U10377 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9154), .Z(n7916) );
  XNOR2_X1 U10378 ( .A(n7916), .B(SI_31_), .ZN(n7917) );
  NOR2_X1 U10379 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n7918) );
  NAND4_X1 U10380 ( .A1(n7920), .A2(n7919), .A3(n8161), .A4(n7918), .ZN(n7922)
         );
  NOR2_X1 U10381 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n7927) );
  NAND4_X1 U10382 ( .A1(n7927), .A2(n7926), .A3(n8521), .A4(n7255), .ZN(n7933)
         );
  XNOR2_X2 U10383 ( .A(n7928), .B(n7929), .ZN(n8530) );
  NAND3_X1 U10384 ( .A1(n7931), .A2(n7930), .A3(n7929), .ZN(n7932) );
  NOR2_X1 U10385 ( .A1(n7933), .A2(n7932), .ZN(n7934) );
  NAND2_X1 U10386 ( .A1(n7939), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7936) );
  NAND2_X1 U10387 ( .A1(n11567), .A2(n8460), .ZN(n7938) );
  NAND2_X1 U10388 ( .A1(n8471), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7937) );
  INV_X1 U10389 ( .A(n13826), .ZN(n7959) );
  INV_X1 U10390 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n7945) );
  AND2_X2 U10391 ( .A1(n7960), .A2(n13826), .ZN(n8243) );
  NAND2_X1 U10392 ( .A1(n8243), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n7944) );
  NAND2_X1 U10393 ( .A1(n8012), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n7943) );
  OAI211_X1 U10394 ( .C1(n8027), .C2(n7945), .A(n7944), .B(n7943), .ZN(n13494)
         );
  NOR2_X1 U10395 ( .A1(n13733), .A2(n13494), .ZN(n7953) );
  INV_X1 U10396 ( .A(n13494), .ZN(n7957) );
  NOR2_X1 U10397 ( .A1(n7958), .A2(n7957), .ZN(n7952) );
  NAND2_X1 U10398 ( .A1(n7947), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7946) );
  NAND2_X1 U10399 ( .A1(n6543), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7949) );
  NAND2_X1 U10400 ( .A1(n13838), .A2(n10114), .ZN(n9544) );
  INV_X1 U10401 ( .A(n13838), .ZN(n7954) );
  NAND2_X1 U10402 ( .A1(n7954), .A2(n10494), .ZN(n7955) );
  NAND2_X1 U10403 ( .A1(n9846), .A2(n7955), .ZN(n7956) );
  OR2_X1 U10404 ( .A1(n9838), .A2(n10114), .ZN(n10365) );
  NAND2_X1 U10405 ( .A1(n7956), .A2(n10365), .ZN(n8507) );
  NAND2_X1 U10406 ( .A1(n11869), .A2(n10389), .ZN(n8504) );
  NAND2_X1 U10407 ( .A1(n8507), .A2(n8504), .ZN(n8509) );
  XNOR2_X1 U10408 ( .A(n7958), .B(n7957), .ZN(n8508) );
  NOR2_X1 U10409 ( .A1(n8508), .A2(n8507), .ZN(n8487) );
  NAND2_X1 U10410 ( .A1(n8012), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U10411 ( .A1(n8243), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n7967) );
  AND2_X2 U10412 ( .A1(n7960), .A2(n7959), .ZN(n8420) );
  NAND2_X1 U10413 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n8049) );
  NOR2_X1 U10414 ( .A1(n8049), .A2(n8048), .ZN(n8061) );
  NAND2_X1 U10415 ( .A1(n8061), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8097) );
  NAND2_X1 U10416 ( .A1(n8134), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8153) );
  NAND2_X1 U10417 ( .A1(n8190), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8216) );
  NAND2_X1 U10418 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n7961) );
  INV_X1 U10419 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8329) );
  INV_X1 U10420 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n13257) );
  NAND2_X1 U10421 ( .A1(n8363), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8378) );
  INV_X1 U10422 ( .A(n8378), .ZN(n7962) );
  NAND2_X1 U10423 ( .A1(n7962), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n8390) );
  NAND2_X1 U10424 ( .A1(n8377), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8407) );
  NAND2_X1 U10425 ( .A1(n8389), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8418) );
  INV_X1 U10426 ( .A(n8418), .ZN(n8406) );
  NAND2_X1 U10427 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n8406), .ZN(n8438) );
  INV_X1 U10428 ( .A(n8438), .ZN(n7963) );
  NAND2_X1 U10429 ( .A1(n7963), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8453) );
  INV_X1 U10430 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7964) );
  NOR2_X1 U10431 ( .A1(n8453), .A2(n7964), .ZN(n13544) );
  NAND2_X1 U10432 ( .A1(n8420), .A2(n13544), .ZN(n7966) );
  NAND2_X1 U10433 ( .A1(n8011), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7965) );
  AND4_X1 U10434 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n11865)
         );
  NAND2_X1 U10435 ( .A1(n13200), .A2(n8414), .ZN(n7972) );
  NAND2_X1 U10436 ( .A1(n8471), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7971) );
  INV_X1 U10437 ( .A(n8106), .ZN(n8479) );
  MUX2_X1 U10438 ( .A(n11865), .B(n13739), .S(n8479), .Z(n8465) );
  NAND2_X1 U10439 ( .A1(n8243), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n7976) );
  NAND2_X1 U10440 ( .A1(n8012), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n7975) );
  NAND2_X1 U10441 ( .A1(n8011), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10442 ( .A1(n8420), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n7973) );
  AND4_X2 U10443 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n9840)
         );
  INV_X1 U10444 ( .A(SI_0_), .ZN(n7977) );
  NOR2_X1 U10445 ( .A1(n9154), .A2(n7977), .ZN(n7978) );
  INV_X1 U10446 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8587) );
  XNOR2_X1 U10447 ( .A(n7978), .B(n8587), .ZN(n13840) );
  NAND2_X1 U10448 ( .A1(n9840), .A2(n13724), .ZN(n8494) );
  NAND2_X1 U10449 ( .A1(n8494), .A2(n9838), .ZN(n7979) );
  INV_X1 U10450 ( .A(n9840), .ZN(n13355) );
  NAND2_X1 U10451 ( .A1(n10611), .A2(n13355), .ZN(n8493) );
  NAND2_X1 U10452 ( .A1(n7979), .A2(n8493), .ZN(n7980) );
  INV_X1 U10453 ( .A(n8494), .ZN(n9704) );
  MUX2_X1 U10454 ( .A(n7980), .B(n9704), .S(n8399), .Z(n7990) );
  XNOR2_X1 U10455 ( .A(n7982), .B(n7981), .ZN(n9302) );
  INV_X1 U10456 ( .A(n9302), .ZN(n7983) );
  NAND2_X1 U10457 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n7984) );
  XNOR2_X1 U10458 ( .A(n7984), .B(P1_IR_REG_1__SCAN_IN), .ZN(n13359) );
  INV_X1 U10459 ( .A(n13359), .ZN(n7985) );
  NAND2_X1 U10460 ( .A1(n8420), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n7989) );
  NAND2_X1 U10461 ( .A1(n8011), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n7988) );
  NAND2_X1 U10462 ( .A1(n8012), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n7987) );
  NAND2_X1 U10463 ( .A1(n8243), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7986) );
  NAND2_X1 U10464 ( .A1(n7990), .A2(n10613), .ZN(n7992) );
  NAND2_X1 U10465 ( .A1(n7992), .A2(n7991), .ZN(n8002) );
  XNOR2_X1 U10466 ( .A(n7994), .B(n7993), .ZN(n9347) );
  NAND2_X1 U10467 ( .A1(n8043), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7997) );
  XNOR2_X1 U10468 ( .A(n7995), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13376) );
  NAND2_X1 U10469 ( .A1(n8310), .A2(n13376), .ZN(n7996) );
  NAND2_X1 U10470 ( .A1(n8420), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n8001) );
  NAND2_X1 U10471 ( .A1(n8243), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8000) );
  NAND2_X1 U10472 ( .A1(n8011), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U10473 ( .A1(n8012), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n7998) );
  NAND4_X1 U10474 ( .A1(n8001), .A2(n8000), .A3(n7999), .A4(n7998), .ZN(n13353) );
  NAND2_X1 U10475 ( .A1(n8002), .A2(n9707), .ZN(n8021) );
  XNOR2_X1 U10476 ( .A(n8003), .B(n8004), .ZN(n9512) );
  NAND2_X1 U10477 ( .A1(n8005), .A2(n9512), .ZN(n8010) );
  NAND2_X1 U10478 ( .A1(n8043), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8009) );
  NAND2_X1 U10479 ( .A1(n8006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8007) );
  XNOR2_X1 U10480 ( .A(n8007), .B(P1_IR_REG_3__SCAN_IN), .ZN(n13388) );
  NAND2_X1 U10481 ( .A1(n8310), .A2(n13388), .ZN(n8008) );
  INV_X1 U10482 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8025) );
  NAND2_X1 U10483 ( .A1(n8420), .A2(n8025), .ZN(n8016) );
  NAND2_X1 U10484 ( .A1(n8243), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8015) );
  NAND2_X1 U10485 ( .A1(n8011), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10486 ( .A1(n8012), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8013) );
  NAND4_X1 U10487 ( .A1(n8016), .A2(n8015), .A3(n8014), .A4(n8013), .ZN(n13352) );
  NAND2_X1 U10488 ( .A1(n10367), .A2(n13352), .ZN(n8022) );
  INV_X1 U10489 ( .A(n10367), .ZN(n14309) );
  NAND2_X1 U10490 ( .A1(n10572), .A2(n14309), .ZN(n10377) );
  NAND2_X1 U10491 ( .A1(n8479), .A2(n10577), .ZN(n8019) );
  NAND2_X1 U10492 ( .A1(n6815), .A2(n8271), .ZN(n8018) );
  MUX2_X1 U10493 ( .A(n8019), .B(n8018), .S(n13353), .Z(n8020) );
  MUX2_X1 U10494 ( .A(n10377), .B(n8022), .S(n8399), .Z(n8023) );
  NAND2_X1 U10495 ( .A1(n8012), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8031) );
  NAND2_X1 U10496 ( .A1(n8243), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8030) );
  INV_X1 U10497 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n8024) );
  NAND2_X1 U10498 ( .A1(n8025), .A2(n8024), .ZN(n8026) );
  AND2_X1 U10499 ( .A1(n8026), .A2(n8049), .ZN(n10654) );
  NAND2_X1 U10500 ( .A1(n8420), .A2(n10654), .ZN(n8029) );
  NAND2_X1 U10501 ( .A1(n8011), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n8028) );
  XNOR2_X1 U10502 ( .A(n8033), .B(n8032), .ZN(n9622) );
  NAND2_X1 U10503 ( .A1(n9622), .A2(n8414), .ZN(n8038) );
  NAND2_X1 U10504 ( .A1(n8471), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8037) );
  NAND2_X1 U10505 ( .A1(n8044), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8035) );
  XNOR2_X1 U10506 ( .A(n8035), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13400) );
  NAND2_X1 U10507 ( .A1(n8310), .A2(n13400), .ZN(n8036) );
  MUX2_X1 U10508 ( .A(n10370), .B(n14367), .S(n8399), .Z(n8040) );
  INV_X1 U10509 ( .A(n14367), .ZN(n10652) );
  INV_X1 U10510 ( .A(n10370), .ZN(n13351) );
  MUX2_X1 U10511 ( .A(n10652), .B(n13351), .S(n8399), .Z(n8039) );
  XNOR2_X1 U10512 ( .A(n8041), .B(n8042), .ZN(n9795) );
  NAND2_X1 U10513 ( .A1(n9795), .A2(n8460), .ZN(n8047) );
  NOR2_X1 U10514 ( .A1(n8044), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n8070) );
  OR2_X1 U10515 ( .A1(n8070), .A2(n13816), .ZN(n8045) );
  XNOR2_X1 U10516 ( .A(n8045), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9449) );
  AOI22_X1 U10517 ( .A1(n8471), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n8310), .B2(
        n9449), .ZN(n8046) );
  NAND2_X1 U10518 ( .A1(n8047), .A2(n8046), .ZN(n14376) );
  NAND2_X1 U10519 ( .A1(n8243), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8054) );
  NAND2_X1 U10520 ( .A1(n8012), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8053) );
  AND2_X1 U10521 ( .A1(n8049), .A2(n8048), .ZN(n8050) );
  NOR2_X1 U10522 ( .A1(n8061), .A2(n8050), .ZN(n10498) );
  NAND2_X1 U10523 ( .A1(n8420), .A2(n10498), .ZN(n8052) );
  NAND2_X1 U10524 ( .A1(n8011), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n8051) );
  NAND4_X1 U10525 ( .A1(n8054), .A2(n8053), .A3(n8052), .A4(n8051), .ZN(n13350) );
  MUX2_X1 U10526 ( .A(n14376), .B(n13350), .S(n8399), .Z(n8057) );
  NAND2_X1 U10527 ( .A1(n8058), .A2(n8057), .ZN(n8056) );
  MUX2_X1 U10528 ( .A(n13350), .B(n14376), .S(n8399), .Z(n8055) );
  NAND2_X1 U10529 ( .A1(n8056), .A2(n8055), .ZN(n8060) );
  NAND2_X1 U10530 ( .A1(n8243), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n8066) );
  NAND2_X1 U10531 ( .A1(n8011), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n8065) );
  OR2_X1 U10532 ( .A1(n8061), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n8062) );
  AND2_X1 U10533 ( .A1(n8097), .A2(n8062), .ZN(n14296) );
  NAND2_X1 U10534 ( .A1(n8420), .A2(n14296), .ZN(n8064) );
  NAND2_X1 U10535 ( .A1(n8012), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n8063) );
  NAND4_X1 U10536 ( .A1(n8066), .A2(n8065), .A3(n8064), .A4(n8063), .ZN(n13349) );
  XNOR2_X1 U10537 ( .A(n8068), .B(n8067), .ZN(n9859) );
  NAND2_X1 U10538 ( .A1(n9859), .A2(n8414), .ZN(n8073) );
  INV_X1 U10539 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8069) );
  NAND2_X1 U10540 ( .A1(n8070), .A2(n8069), .ZN(n8078) );
  NAND2_X1 U10541 ( .A1(n8078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8071) );
  XNOR2_X1 U10542 ( .A(n8071), .B(P1_IR_REG_6__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U10543 ( .A1(n8471), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8310), .B2(
        n13413), .ZN(n8072) );
  NAND2_X1 U10544 ( .A1(n8073), .A2(n8072), .ZN(n10559) );
  MUX2_X1 U10545 ( .A(n13349), .B(n10559), .S(n8017), .Z(n8108) );
  OR2_X1 U10546 ( .A1(n8075), .A2(n8074), .ZN(n8076) );
  OR2_X1 U10547 ( .A1(n10085), .A2(n6455), .ZN(n8081) );
  NAND2_X1 U10548 ( .A1(n8124), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8079) );
  XNOR2_X1 U10549 ( .A(n8079), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9467) );
  AOI22_X1 U10550 ( .A1(n8471), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8310), .B2(
        n9467), .ZN(n8080) );
  NAND2_X1 U10551 ( .A1(n8243), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n8088) );
  NAND2_X1 U10552 ( .A1(n8012), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n8087) );
  NAND2_X1 U10553 ( .A1(n8099), .A2(n8082), .ZN(n8083) );
  NAND2_X1 U10554 ( .A1(n8115), .A2(n8083), .ZN(n10861) );
  INV_X1 U10555 ( .A(n10861), .ZN(n8084) );
  NAND2_X1 U10556 ( .A1(n8420), .A2(n8084), .ZN(n8086) );
  NAND2_X1 U10557 ( .A1(n8011), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n8085) );
  NAND4_X1 U10558 ( .A1(n8088), .A2(n8087), .A3(n8086), .A4(n8085), .ZN(n13347) );
  XNOR2_X1 U10559 ( .A(n10858), .B(n13347), .ZN(n10407) );
  NAND2_X1 U10560 ( .A1(n8092), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8093) );
  XNOR2_X1 U10561 ( .A(n8093), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U10562 ( .A1(n8471), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8310), .B2(
        n13425), .ZN(n8094) );
  NAND2_X1 U10563 ( .A1(n8095), .A2(n8094), .ZN(n14396) );
  NAND2_X1 U10564 ( .A1(n8243), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8103) );
  NAND2_X1 U10565 ( .A1(n8011), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n8102) );
  NAND2_X1 U10566 ( .A1(n8097), .A2(n8096), .ZN(n8098) );
  AND2_X1 U10567 ( .A1(n8099), .A2(n8098), .ZN(n10698) );
  NAND2_X1 U10568 ( .A1(n8420), .A2(n10698), .ZN(n8101) );
  NAND2_X1 U10569 ( .A1(n8012), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n8100) );
  NAND4_X1 U10570 ( .A1(n8103), .A2(n8102), .A3(n8101), .A4(n8100), .ZN(n13348) );
  MUX2_X1 U10571 ( .A(n14396), .B(n13348), .S(n8271), .Z(n8104) );
  INV_X1 U10572 ( .A(n8104), .ZN(n8110) );
  MUX2_X1 U10573 ( .A(n14396), .B(n13348), .S(n8017), .Z(n8109) );
  NAND2_X1 U10574 ( .A1(n8110), .A2(n8109), .ZN(n8105) );
  INV_X1 U10575 ( .A(n10559), .ZN(n14387) );
  MUX2_X1 U10576 ( .A(n10561), .B(n14387), .S(n8271), .Z(n8107) );
  NOR2_X1 U10577 ( .A1(n8110), .A2(n8109), .ZN(n8113) );
  NAND2_X1 U10578 ( .A1(n10858), .A2(n13347), .ZN(n8112) );
  MUX2_X1 U10579 ( .A(n13347), .B(n10858), .S(n8017), .Z(n8111) );
  AOI22_X1 U10580 ( .A1(n8113), .A2(n10407), .B1(n8112), .B2(n8111), .ZN(n8114) );
  NAND2_X1 U10581 ( .A1(n8012), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n8120) );
  NAND2_X1 U10582 ( .A1(n8243), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n8119) );
  AND2_X1 U10583 ( .A1(n8115), .A2(n9532), .ZN(n8116) );
  NOR2_X1 U10584 ( .A1(n8134), .A2(n8116), .ZN(n10906) );
  NAND2_X1 U10585 ( .A1(n8420), .A2(n10906), .ZN(n8118) );
  NAND2_X1 U10586 ( .A1(n8011), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n8117) );
  NAND2_X1 U10587 ( .A1(n8123), .A2(n8122), .ZN(n10177) );
  OR2_X1 U10588 ( .A1(n10177), .A2(n6455), .ZN(n8128) );
  OAI21_X1 U10589 ( .B1(n8124), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8163) );
  INV_X1 U10590 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8125) );
  OR2_X1 U10591 ( .A1(n8163), .A2(n8125), .ZN(n8126) );
  NAND2_X1 U10592 ( .A1(n8163), .A2(n8125), .ZN(n8143) );
  AOI22_X1 U10593 ( .A1(n8471), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8310), .B2(
        n9471), .ZN(n8127) );
  MUX2_X1 U10594 ( .A(n10974), .B(n14412), .S(n8271), .Z(n8130) );
  MUX2_X1 U10595 ( .A(n13346), .B(n10545), .S(n8017), .Z(n8129) );
  OAI21_X1 U10596 ( .B1(n8131), .B2(n8130), .A(n8129), .ZN(n8133) );
  NAND2_X1 U10597 ( .A1(n8131), .A2(n8130), .ZN(n8132) );
  NAND2_X1 U10598 ( .A1(n8133), .A2(n8132), .ZN(n8150) );
  NAND2_X1 U10599 ( .A1(n8243), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n8139) );
  NAND2_X1 U10600 ( .A1(n8011), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n8138) );
  OR2_X1 U10601 ( .A1(n8134), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n8135) );
  AND2_X1 U10602 ( .A1(n8135), .A2(n8153), .ZN(n10971) );
  NAND2_X1 U10603 ( .A1(n8420), .A2(n10971), .ZN(n8137) );
  NAND2_X1 U10604 ( .A1(n8012), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n8136) );
  NAND4_X1 U10605 ( .A1(n8139), .A2(n8138), .A3(n8137), .A4(n8136), .ZN(n13345) );
  XNOR2_X1 U10606 ( .A(n8140), .B(SI_10_), .ZN(n8141) );
  NAND2_X1 U10607 ( .A1(n10268), .A2(n8414), .ZN(n8146) );
  NAND2_X1 U10608 ( .A1(n8143), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8144) );
  XNOR2_X1 U10609 ( .A(n8144), .B(P1_IR_REG_10__SCAN_IN), .ZN(n13440) );
  AOI22_X1 U10610 ( .A1(n8471), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n13440), 
        .B2(n8310), .ZN(n8145) );
  MUX2_X1 U10611 ( .A(n13345), .B(n10976), .S(n8017), .Z(n8149) );
  NAND2_X1 U10612 ( .A1(n8150), .A2(n8149), .ZN(n8148) );
  MUX2_X1 U10613 ( .A(n13345), .B(n10976), .S(n8271), .Z(n8147) );
  NAND2_X1 U10614 ( .A1(n8148), .A2(n8147), .ZN(n8152) );
  OR2_X1 U10615 ( .A1(n8150), .A2(n8149), .ZN(n8151) );
  NAND2_X1 U10616 ( .A1(n8152), .A2(n8151), .ZN(n8169) );
  NAND2_X1 U10617 ( .A1(n8153), .A2(n14989), .ZN(n8154) );
  AND2_X1 U10618 ( .A1(n8170), .A2(n8154), .ZN(n11115) );
  NAND2_X1 U10619 ( .A1(n8420), .A2(n11115), .ZN(n8158) );
  NAND2_X1 U10620 ( .A1(n8243), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8157) );
  NAND2_X1 U10621 ( .A1(n8011), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U10622 ( .A1(n8012), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n8155) );
  NAND4_X1 U10623 ( .A1(n8158), .A2(n8157), .A3(n8156), .A4(n8155), .ZN(n13344) );
  XNOR2_X1 U10624 ( .A(n8160), .B(n8159), .ZN(n10420) );
  NAND2_X1 U10625 ( .A1(n10420), .A2(n8460), .ZN(n8166) );
  OR2_X1 U10626 ( .A1(n8161), .A2(n13816), .ZN(n8162) );
  NAND2_X1 U10627 ( .A1(n8163), .A2(n8162), .ZN(n8178) );
  INV_X1 U10628 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8164) );
  XNOR2_X1 U10629 ( .A(n8178), .B(n8164), .ZN(n9601) );
  AOI22_X1 U10630 ( .A1(n8471), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8310), 
        .B2(n9601), .ZN(n8165) );
  MUX2_X1 U10631 ( .A(n13344), .B(n11100), .S(n8271), .Z(n8168) );
  MUX2_X1 U10632 ( .A(n13344), .B(n11100), .S(n8017), .Z(n8167) );
  NAND2_X1 U10633 ( .A1(n8012), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U10634 ( .A1(n8243), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n8174) );
  AND2_X1 U10635 ( .A1(n8170), .A2(n9606), .ZN(n8171) );
  NOR2_X1 U10636 ( .A1(n8190), .A2(n8171), .ZN(n11142) );
  NAND2_X1 U10637 ( .A1(n8420), .A2(n11142), .ZN(n8173) );
  NAND2_X1 U10638 ( .A1(n8011), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n8172) );
  NAND4_X1 U10639 ( .A1(n8175), .A2(n8174), .A3(n8173), .A4(n8172), .ZN(n13343) );
  XNOR2_X1 U10640 ( .A(n8177), .B(n8176), .ZN(n10590) );
  NAND2_X1 U10641 ( .A1(n10590), .A2(n8414), .ZN(n8181) );
  NAND2_X1 U10642 ( .A1(n8179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U10643 ( .A(n8200), .B(P1_IR_REG_12__SCAN_IN), .ZN(n13451) );
  AOI22_X1 U10644 ( .A1(n13451), .A2(n8310), .B1(n8471), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n8180) );
  MUX2_X1 U10645 ( .A(n13343), .B(n11131), .S(n8017), .Z(n8185) );
  MUX2_X1 U10646 ( .A(n13343), .B(n11131), .S(n8271), .Z(n8182) );
  NAND2_X1 U10647 ( .A1(n8183), .A2(n8182), .ZN(n8189) );
  INV_X1 U10648 ( .A(n8184), .ZN(n8187) );
  INV_X1 U10649 ( .A(n8185), .ZN(n8186) );
  NAND2_X1 U10650 ( .A1(n8187), .A2(n8186), .ZN(n8188) );
  OR2_X1 U10651 ( .A1(n8190), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n8191) );
  NAND2_X1 U10652 ( .A1(n8216), .A2(n8191), .ZN(n13981) );
  INV_X1 U10653 ( .A(n13981), .ZN(n8192) );
  NAND2_X1 U10654 ( .A1(n8192), .A2(n8420), .ZN(n8196) );
  NAND2_X1 U10655 ( .A1(n8243), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10656 ( .A1(n8011), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8194) );
  NAND2_X1 U10657 ( .A1(n8012), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8193) );
  NAND4_X1 U10658 ( .A1(n8196), .A2(n8195), .A3(n8194), .A4(n8193), .ZN(n13342) );
  XNOR2_X1 U10659 ( .A(n8198), .B(n8197), .ZN(n10757) );
  NAND2_X1 U10660 ( .A1(n10757), .A2(n8414), .ZN(n8206) );
  AOI21_X1 U10661 ( .B1(n8200), .B2(n8199), .A(n13816), .ZN(n8201) );
  NAND2_X1 U10662 ( .A1(n8201), .A2(P1_IR_REG_13__SCAN_IN), .ZN(n8204) );
  INV_X1 U10663 ( .A(n8201), .ZN(n8203) );
  NAND2_X1 U10664 ( .A1(n8203), .A2(n8202), .ZN(n8211) );
  AOI22_X1 U10665 ( .A1(n14190), .A2(n8310), .B1(n8471), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n8205) );
  MUX2_X1 U10666 ( .A(n13342), .B(n14145), .S(n8271), .Z(n8208) );
  MUX2_X1 U10667 ( .A(n13342), .B(n14145), .S(n8017), .Z(n8207) );
  INV_X1 U10668 ( .A(n8208), .ZN(n8209) );
  NAND2_X1 U10669 ( .A1(n10942), .A2(n8460), .ZN(n8214) );
  NAND2_X1 U10670 ( .A1(n8211), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8212) );
  XNOR2_X1 U10671 ( .A(n8212), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14211) );
  AOI22_X1 U10672 ( .A1(n14211), .A2(n8310), .B1(n8471), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n8213) );
  NAND2_X1 U10673 ( .A1(n8216), .A2(n8215), .ZN(n8217) );
  AND2_X1 U10674 ( .A1(n8232), .A2(n8217), .ZN(n13230) );
  AOI22_X1 U10675 ( .A1(n13230), .A2(n8420), .B1(n8011), .B2(
        P1_REG1_REG_14__SCAN_IN), .ZN(n8219) );
  AOI22_X1 U10676 ( .A1(n8243), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8012), .B2(
        P1_REG0_REG_14__SCAN_IN), .ZN(n8218) );
  XNOR2_X1 U10677 ( .A(n14136), .B(n13966), .ZN(n10820) );
  INV_X1 U10678 ( .A(n8220), .ZN(n8224) );
  INV_X1 U10679 ( .A(n8221), .ZN(n8222) );
  XNOR2_X1 U10680 ( .A(n8225), .B(SI_15_), .ZN(n8226) );
  NAND2_X1 U10681 ( .A1(n11024), .A2(n8414), .ZN(n8230) );
  OR2_X1 U10682 ( .A1(n8227), .A2(n13816), .ZN(n8228) );
  INV_X1 U10683 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8248) );
  XNOR2_X1 U10684 ( .A(n8228), .B(n8248), .ZN(n14230) );
  INV_X1 U10685 ( .A(n14230), .ZN(n13473) );
  AOI22_X1 U10686 ( .A1(n8471), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8310), 
        .B2(n13473), .ZN(n8229) );
  AND2_X1 U10687 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  OR2_X1 U10688 ( .A1(n8233), .A2(n8241), .ZN(n13332) );
  AOI22_X1 U10689 ( .A1(n8243), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8012), .B2(
        P1_REG0_REG_15__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10690 ( .A1(n8011), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n8234) );
  OAI211_X1 U10691 ( .C1(n13332), .C2(n8298), .A(n8235), .B(n8234), .ZN(n14088) );
  INV_X1 U10692 ( .A(n14088), .ZN(n13228) );
  NAND2_X1 U10693 ( .A1(n13337), .A2(n13228), .ZN(n8492) );
  NAND2_X1 U10694 ( .A1(n14136), .A2(n13966), .ZN(n8236) );
  NAND2_X1 U10695 ( .A1(n8492), .A2(n8236), .ZN(n8238) );
  OR2_X1 U10696 ( .A1(n14136), .A2(n13966), .ZN(n10994) );
  NAND2_X1 U10697 ( .A1(n11147), .A2(n10994), .ZN(n8237) );
  MUX2_X1 U10698 ( .A(n8238), .B(n8237), .S(n8271), .Z(n8240) );
  MUX2_X1 U10699 ( .A(n8492), .B(n11147), .S(n8017), .Z(n8239) );
  NOR2_X1 U10700 ( .A1(n8241), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8242) );
  OR2_X1 U10701 ( .A1(n8252), .A2(n8242), .ZN(n14092) );
  AOI22_X1 U10702 ( .A1(n8011), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8243), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n8245) );
  NAND2_X1 U10703 ( .A1(n8012), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8244) );
  OAI211_X1 U10704 ( .C1(n14092), .C2(n8298), .A(n8245), .B(n8244), .ZN(n13340) );
  NAND2_X1 U10705 ( .A1(n11168), .A2(n8460), .ZN(n8251) );
  AND2_X1 U10706 ( .A1(n8227), .A2(n8248), .ZN(n8264) );
  OR2_X1 U10707 ( .A1(n8264), .A2(n13816), .ZN(n8249) );
  XNOR2_X1 U10708 ( .A(n8249), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14239) );
  AOI22_X1 U10709 ( .A1(n8471), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8310), 
        .B2(n14239), .ZN(n8250) );
  MUX2_X1 U10710 ( .A(n13340), .B(n14089), .S(n8271), .Z(n8286) );
  OR2_X1 U10711 ( .A1(n8252), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8253) );
  AND2_X1 U10712 ( .A1(n8313), .A2(n8253), .ZN(n13281) );
  NAND2_X1 U10713 ( .A1(n13281), .A2(n8420), .ZN(n8259) );
  INV_X1 U10714 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U10715 ( .A1(n8012), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U10716 ( .A1(n8011), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8254) );
  OAI211_X1 U10717 ( .C1(n8317), .C2(n8256), .A(n8255), .B(n8254), .ZN(n8257)
         );
  INV_X1 U10718 ( .A(n8257), .ZN(n8258) );
  NAND2_X1 U10719 ( .A1(n8286), .A2(n14086), .ZN(n8270) );
  OR2_X1 U10720 ( .A1(n13340), .A2(n8399), .ZN(n8273) );
  XNOR2_X1 U10721 ( .A(n8261), .B(SI_17_), .ZN(n8262) );
  XNOR2_X1 U10722 ( .A(n8260), .B(n8262), .ZN(n11408) );
  NAND2_X1 U10723 ( .A1(n11408), .A2(n8460), .ZN(n8269) );
  INV_X1 U10724 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U10725 ( .A1(n8264), .A2(n8263), .ZN(n8266) );
  NAND2_X1 U10726 ( .A1(n8266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8265) );
  MUX2_X1 U10727 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8265), .S(
        P1_IR_REG_17__SCAN_IN), .Z(n8267) );
  AND2_X1 U10728 ( .A1(n8267), .A2(n8307), .ZN(n14258) );
  AOI22_X1 U10729 ( .A1(n8471), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8310), 
        .B2(n14258), .ZN(n8268) );
  AOI21_X1 U10730 ( .B1(n8270), .B2(n8273), .A(n13522), .ZN(n8277) );
  INV_X1 U10731 ( .A(n14086), .ZN(n11765) );
  NAND2_X1 U10732 ( .A1(n8286), .A2(n11765), .ZN(n8272) );
  OR2_X1 U10733 ( .A1(n14089), .A2(n8271), .ZN(n8278) );
  AOI21_X1 U10734 ( .B1(n8272), .B2(n8278), .A(n14116), .ZN(n8276) );
  NAND2_X1 U10735 ( .A1(n14086), .A2(n8479), .ZN(n8279) );
  OR2_X1 U10736 ( .A1(n14089), .A2(n8279), .ZN(n8275) );
  INV_X1 U10737 ( .A(n8273), .ZN(n8282) );
  NAND2_X1 U10738 ( .A1(n8282), .A2(n11765), .ZN(n8274) );
  NAND2_X1 U10739 ( .A1(n8275), .A2(n8274), .ZN(n8285) );
  INV_X1 U10740 ( .A(n8278), .ZN(n8281) );
  INV_X1 U10741 ( .A(n8279), .ZN(n8280) );
  AOI21_X1 U10742 ( .B1(n8286), .B2(n8281), .A(n8280), .ZN(n8289) );
  NAND2_X1 U10743 ( .A1(n8286), .A2(n8282), .ZN(n8283) );
  OAI21_X1 U10744 ( .B1(n8479), .B2(n14086), .A(n8283), .ZN(n8284) );
  NAND2_X1 U10745 ( .A1(n8284), .A2(n14116), .ZN(n8288) );
  NAND2_X1 U10746 ( .A1(n8286), .A2(n8285), .ZN(n8287) );
  OAI211_X1 U10747 ( .C1(n8289), .C2(n14116), .A(n8288), .B(n8287), .ZN(n8290)
         );
  INV_X1 U10748 ( .A(n8290), .ZN(n8321) );
  AOI22_X1 U10749 ( .A1(n8471), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n13486), 
        .B2(n8310), .ZN(n8293) );
  INV_X1 U10750 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8296) );
  INV_X1 U10751 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8295) );
  OAI21_X1 U10752 ( .B1(n8313), .B2(n8296), .A(n8295), .ZN(n8297) );
  NAND2_X1 U10753 ( .A1(n8297), .A2(n8330), .ZN(n13695) );
  OR2_X1 U10754 ( .A1(n13695), .A2(n8298), .ZN(n8304) );
  INV_X1 U10755 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n8301) );
  NAND2_X1 U10756 ( .A1(n8012), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8300) );
  NAND2_X1 U10757 ( .A1(n8011), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8299) );
  OAI211_X1 U10758 ( .C1(n8317), .C2(n8301), .A(n8300), .B(n8299), .ZN(n8302)
         );
  INV_X1 U10759 ( .A(n8302), .ZN(n8303) );
  NAND2_X1 U10760 ( .A1(n8304), .A2(n8303), .ZN(n13709) );
  XNOR2_X1 U10761 ( .A(n8305), .B(n8306), .ZN(n11417) );
  NAND2_X1 U10762 ( .A1(n11417), .A2(n8460), .ZN(n8312) );
  NAND2_X1 U10763 ( .A1(n8307), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8309) );
  INV_X1 U10764 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n8308) );
  XNOR2_X1 U10765 ( .A(n8309), .B(n8308), .ZN(n13479) );
  INV_X1 U10766 ( .A(n13479), .ZN(n14275) );
  AOI22_X1 U10767 ( .A1(n8471), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8310), 
        .B2(n14275), .ZN(n8311) );
  XNOR2_X1 U10768 ( .A(n8313), .B(P1_REG3_REG_18__SCAN_IN), .ZN(n13716) );
  NAND2_X1 U10769 ( .A1(n13716), .A2(n8420), .ZN(n8320) );
  INV_X1 U10770 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10771 ( .A1(n8012), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10772 ( .A1(n8011), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8314) );
  OAI211_X1 U10773 ( .C1(n8317), .C2(n8316), .A(n8315), .B(n8314), .ZN(n8318)
         );
  INV_X1 U10774 ( .A(n8318), .ZN(n8319) );
  NAND2_X1 U10775 ( .A1(n8320), .A2(n8319), .ZN(n13507) );
  XNOR2_X1 U10776 ( .A(n13717), .B(n13507), .ZN(n13707) );
  INV_X1 U10777 ( .A(n13507), .ZN(n13525) );
  NAND3_X1 U10778 ( .A1(n13717), .A2(n13525), .A3(n8399), .ZN(n8323) );
  OR3_X1 U10779 ( .A1(n13717), .A2(n13525), .A3(n8479), .ZN(n8322) );
  NAND2_X1 U10780 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND2_X1 U10781 ( .A1(n8491), .A2(n8324), .ZN(n8328) );
  NAND2_X1 U10782 ( .A1(n13700), .A2(n8479), .ZN(n8326) );
  OR2_X1 U10783 ( .A1(n13700), .A2(n8399), .ZN(n8325) );
  NAND2_X1 U10784 ( .A1(n8330), .A2(n8329), .ZN(n8331) );
  NAND2_X1 U10785 ( .A1(n8344), .A2(n8331), .ZN(n13296) );
  INV_X1 U10786 ( .A(n13296), .ZN(n13687) );
  NAND2_X1 U10787 ( .A1(n13687), .A2(n8420), .ZN(n8337) );
  INV_X1 U10788 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n15000) );
  NAND2_X1 U10789 ( .A1(n8243), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8333) );
  NAND2_X1 U10790 ( .A1(n8011), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n8332) );
  OAI211_X1 U10791 ( .C1(n15000), .C2(n8334), .A(n8333), .B(n8332), .ZN(n8335)
         );
  INV_X1 U10792 ( .A(n8335), .ZN(n8336) );
  MUX2_X1 U10793 ( .A(n13256), .B(n7031), .S(n8017), .Z(n8339) );
  NAND2_X1 U10794 ( .A1(n8341), .A2(n8340), .ZN(n8342) );
  AND2_X1 U10795 ( .A1(n8344), .A2(n13257), .ZN(n8345) );
  OR2_X1 U10796 ( .A1(n8345), .A2(n8363), .ZN(n13669) );
  INV_X1 U10797 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10798 ( .A1(n8243), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U10799 ( .A1(n8012), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8346) );
  OAI211_X1 U10800 ( .C1(n8027), .C2(n8348), .A(n8347), .B(n8346), .ZN(n8349)
         );
  INV_X1 U10801 ( .A(n8349), .ZN(n8350) );
  NAND2_X1 U10802 ( .A1(n8352), .A2(n8351), .ZN(n8355) );
  OR2_X1 U10803 ( .A1(n8353), .A2(n10110), .ZN(n8354) );
  NAND2_X1 U10804 ( .A1(n8355), .A2(n8354), .ZN(n8358) );
  XNOR2_X1 U10805 ( .A(n8356), .B(SI_21_), .ZN(n8357) );
  NAND2_X1 U10806 ( .A1(n11464), .A2(n8414), .ZN(n8360) );
  NAND2_X1 U10807 ( .A1(n8471), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8359) );
  MUX2_X1 U10808 ( .A(n13678), .B(n13529), .S(n8017), .Z(n8362) );
  MUX2_X1 U10809 ( .A(n13678), .B(n13529), .S(n8106), .Z(n8361) );
  OR2_X1 U10810 ( .A1(n8363), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n8364) );
  AND2_X1 U10811 ( .A1(n8364), .A2(n8378), .ZN(n13657) );
  NAND2_X1 U10812 ( .A1(n13657), .A2(n8420), .ZN(n8370) );
  INV_X1 U10813 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U10814 ( .A1(n8012), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8366) );
  NAND2_X1 U10815 ( .A1(n8243), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n8365) );
  OAI211_X1 U10816 ( .C1(n8367), .C2(n8027), .A(n8366), .B(n8365), .ZN(n8368)
         );
  INV_X1 U10817 ( .A(n8368), .ZN(n8369) );
  NAND2_X1 U10818 ( .A1(n8370), .A2(n8369), .ZN(n13513) );
  XNOR2_X1 U10819 ( .A(n8372), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n13839) );
  MUX2_X1 U10820 ( .A(n13513), .B(n13661), .S(n8106), .Z(n8375) );
  NAND2_X1 U10821 ( .A1(n8376), .A2(n8375), .ZN(n8374) );
  MUX2_X1 U10822 ( .A(n13513), .B(n13661), .S(n8017), .Z(n8373) );
  NAND2_X1 U10823 ( .A1(n8012), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n8382) );
  NAND2_X1 U10824 ( .A1(n8243), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n8381) );
  INV_X1 U10825 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13239) );
  AOI21_X1 U10826 ( .B1(n13239), .B2(n8378), .A(n8377), .ZN(n13643) );
  NAND2_X1 U10827 ( .A1(n8420), .A2(n13643), .ZN(n8380) );
  NAND2_X1 U10828 ( .A1(n8011), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n8379) );
  NAND4_X1 U10829 ( .A1(n8382), .A2(n8381), .A3(n8380), .A4(n8379), .ZN(n13516) );
  NAND2_X1 U10830 ( .A1(n11499), .A2(n8460), .ZN(n8385) );
  NAND2_X1 U10831 ( .A1(n8471), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n8384) );
  MUX2_X1 U10832 ( .A(n13516), .B(n13778), .S(n8271), .Z(n8386) );
  INV_X1 U10833 ( .A(n8387), .ZN(n8388) );
  NAND2_X1 U10834 ( .A1(n8243), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10835 ( .A1(n8012), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n8393) );
  INV_X1 U10836 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n13288) );
  AOI21_X1 U10837 ( .B1(n13288), .B2(n8390), .A(n8389), .ZN(n13630) );
  NAND2_X1 U10838 ( .A1(n8420), .A2(n13630), .ZN(n8392) );
  NAND2_X1 U10839 ( .A1(n8011), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8391) );
  XNOR2_X1 U10840 ( .A(n8395), .B(n8396), .ZN(n11513) );
  NAND2_X1 U10841 ( .A1(n11513), .A2(n8460), .ZN(n8398) );
  NAND2_X1 U10842 ( .A1(n8471), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10843 ( .A1(n8403), .A2(n8402), .ZN(n8401) );
  MUX2_X1 U10844 ( .A(n13607), .B(n13772), .S(n8271), .Z(n8400) );
  NAND2_X1 U10845 ( .A1(n8401), .A2(n8400), .ZN(n8405) );
  NAND2_X1 U10846 ( .A1(n8243), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n8411) );
  NAND2_X1 U10847 ( .A1(n8011), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8410) );
  INV_X1 U10848 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n13266) );
  AOI21_X1 U10849 ( .B1(n13266), .B2(n8407), .A(n8406), .ZN(n13611) );
  NAND2_X1 U10850 ( .A1(n8420), .A2(n13611), .ZN(n8409) );
  NAND2_X1 U10851 ( .A1(n8012), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8408) );
  NAND4_X1 U10852 ( .A1(n8411), .A2(n8410), .A3(n8409), .A4(n8408), .ZN(n13533) );
  XNOR2_X1 U10853 ( .A(n8413), .B(n8412), .ZN(n11527) );
  NAND2_X1 U10854 ( .A1(n8471), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8415) );
  MUX2_X1 U10855 ( .A(n13533), .B(n13763), .S(n8271), .Z(n8416) );
  NAND2_X1 U10856 ( .A1(n8012), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8424) );
  NAND2_X1 U10857 ( .A1(n8243), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n8423) );
  INV_X1 U10858 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U10859 ( .A1(n13324), .A2(n8418), .ZN(n8419) );
  AND2_X1 U10860 ( .A1(n8419), .A2(n8438), .ZN(n13594) );
  NAND2_X1 U10861 ( .A1(n8420), .A2(n13594), .ZN(n8422) );
  NAND2_X1 U10862 ( .A1(n8011), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8421) );
  NAND4_X1 U10863 ( .A1(n8424), .A2(n8423), .A3(n8422), .A4(n8421), .ZN(n13608) );
  XNOR2_X1 U10864 ( .A(n8425), .B(SI_26_), .ZN(n8426) );
  XNOR2_X1 U10865 ( .A(n8427), .B(n8426), .ZN(n13208) );
  NAND2_X1 U10866 ( .A1(n13208), .A2(n8460), .ZN(n8429) );
  NAND2_X1 U10867 ( .A1(n8471), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8428) );
  MUX2_X1 U10868 ( .A(n13608), .B(n13491), .S(n8271), .Z(n8433) );
  NAND2_X1 U10869 ( .A1(n8432), .A2(n8433), .ZN(n8431) );
  MUX2_X1 U10870 ( .A(n13608), .B(n13491), .S(n8479), .Z(n8430) );
  NAND2_X1 U10871 ( .A1(n8431), .A2(n8430), .ZN(n8437) );
  INV_X1 U10872 ( .A(n8432), .ZN(n8435) );
  INV_X1 U10873 ( .A(n8433), .ZN(n8434) );
  NAND2_X1 U10874 ( .A1(n8435), .A2(n8434), .ZN(n8436) );
  NAND2_X1 U10875 ( .A1(n8012), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n8443) );
  NAND2_X1 U10876 ( .A1(n8243), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n8442) );
  INV_X1 U10877 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n13220) );
  NAND2_X1 U10878 ( .A1(n8438), .A2(n13220), .ZN(n8439) );
  NAND2_X1 U10879 ( .A1(n8420), .A2(n13579), .ZN(n8441) );
  NAND2_X1 U10880 ( .A1(n8011), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8440) );
  NAND4_X1 U10881 ( .A1(n8443), .A2(n8442), .A3(n8441), .A4(n8440), .ZN(n13556) );
  INV_X1 U10882 ( .A(n8444), .ZN(n8445) );
  XNOR2_X1 U10883 ( .A(n8445), .B(SI_27_), .ZN(n8446) );
  NAND2_X1 U10884 ( .A1(n13204), .A2(n8460), .ZN(n8449) );
  NAND2_X1 U10885 ( .A1(n8471), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8448) );
  MUX2_X1 U10886 ( .A(n13556), .B(n13750), .S(n8479), .Z(n8451) );
  MUX2_X1 U10887 ( .A(n13556), .B(n13750), .S(n8271), .Z(n8450) );
  NAND2_X1 U10888 ( .A1(n8012), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10889 ( .A1(n8243), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n8456) );
  XNOR2_X1 U10890 ( .A(n8453), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13563) );
  NAND2_X1 U10891 ( .A1(n8420), .A2(n13563), .ZN(n8455) );
  NAND2_X1 U10892 ( .A1(n8011), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n8454) );
  NAND4_X1 U10893 ( .A1(n8457), .A2(n8456), .A3(n8455), .A4(n8454), .ZN(n13547) );
  NAND2_X1 U10894 ( .A1(n8471), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8461) );
  INV_X1 U10895 ( .A(n11865), .ZN(n13557) );
  MUX2_X1 U10896 ( .A(n13557), .B(n6453), .S(n8271), .Z(n8464) );
  NAND2_X1 U10897 ( .A1(n8471), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U10898 ( .A1(n8011), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n8476) );
  NAND2_X1 U10899 ( .A1(n8243), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10900 ( .A1(n8012), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8474) );
  AND3_X1 U10901 ( .A1(n8476), .A2(n8475), .A3(n8474), .ZN(n8480) );
  AOI22_X1 U10902 ( .A1(n8479), .A2(n13494), .B1(n11869), .B2(n8477), .ZN(
        n8478) );
  OAI22_X1 U10903 ( .A1(n13736), .A2(n8479), .B1(n8480), .B2(n8478), .ZN(n8483) );
  INV_X1 U10904 ( .A(n8480), .ZN(n13543) );
  OAI21_X1 U10905 ( .B1(n13494), .B2(n10494), .A(n13543), .ZN(n8481) );
  MUX2_X1 U10906 ( .A(n13736), .B(n8481), .S(n8106), .Z(n8482) );
  XOR2_X1 U10907 ( .A(n13557), .B(n6453), .Z(n13538) );
  INV_X1 U10908 ( .A(n13547), .ZN(n13521) );
  NAND2_X1 U10909 ( .A1(n13745), .A2(n13521), .ZN(n13537) );
  OR2_X1 U10910 ( .A1(n13745), .A2(n13521), .ZN(n8488) );
  INV_X1 U10911 ( .A(n13556), .ZN(n13520) );
  NAND2_X1 U10912 ( .A1(n13750), .A2(n13520), .ZN(n13536) );
  NAND2_X1 U10913 ( .A1(n13491), .A2(n15021), .ZN(n13535) );
  INV_X1 U10914 ( .A(n13516), .ZN(n13532) );
  INV_X1 U10915 ( .A(n13513), .ZN(n13530) );
  XNOR2_X1 U10916 ( .A(n13786), .B(n13530), .ZN(n13531) );
  INV_X1 U10917 ( .A(n13707), .ZN(n13526) );
  XNOR2_X1 U10918 ( .A(n14145), .B(n11200), .ZN(n13971) );
  XNOR2_X1 U10919 ( .A(n11131), .B(n13964), .ZN(n10816) );
  XNOR2_X1 U10920 ( .A(n11100), .B(n13344), .ZN(n10790) );
  XNOR2_X1 U10921 ( .A(n14396), .B(n13348), .ZN(n10387) );
  INV_X1 U10922 ( .A(n9707), .ZN(n10569) );
  INV_X1 U10923 ( .A(n10375), .ZN(n9700) );
  NAND2_X1 U10924 ( .A1(n8494), .A2(n8493), .ZN(n13723) );
  NOR4_X1 U10925 ( .A1(n10569), .A2(n9700), .A3(n7321), .A4(n13723), .ZN(n8495) );
  XNOR2_X1 U10926 ( .A(n14376), .B(n13350), .ZN(n10496) );
  XNOR2_X1 U10927 ( .A(n10652), .B(n13351), .ZN(n10647) );
  NAND4_X1 U10928 ( .A1(n10387), .A2(n8495), .A3(n10496), .A4(n10647), .ZN(
        n8496) );
  NOR3_X1 U10929 ( .A1(n8496), .A2(n14291), .A3(n10448), .ZN(n8497) );
  XNOR2_X1 U10930 ( .A(n10976), .B(n13345), .ZN(n10410) );
  XNOR2_X1 U10931 ( .A(n10545), .B(n13346), .ZN(n10536) );
  NAND4_X1 U10932 ( .A1(n10410), .A2(n8497), .A3(n10790), .A4(n10536), .ZN(
        n8498) );
  NOR3_X1 U10933 ( .A1(n13971), .A2(n10816), .A3(n8498), .ZN(n8499) );
  NAND2_X1 U10934 ( .A1(n14116), .A2(n14086), .ZN(n13506) );
  NAND2_X1 U10935 ( .A1(n13503), .A2(n13506), .ZN(n11153) );
  XNOR2_X1 U10936 ( .A(n14089), .B(n13340), .ZN(n11149) );
  NAND4_X1 U10937 ( .A1(n11145), .A2(n8499), .A3(n11153), .A4(n11149), .ZN(
        n8500) );
  NOR4_X1 U10938 ( .A1(n13701), .A2(n13526), .A3(n10820), .A4(n8500), .ZN(
        n8501) );
  XNOR2_X1 U10939 ( .A(n7031), .B(n13256), .ZN(n13684) );
  NAND4_X1 U10940 ( .A1(n13531), .A2(n8501), .A3(n13684), .A4(n13667), .ZN(
        n8502) );
  XNOR2_X1 U10941 ( .A(n13763), .B(n13533), .ZN(n13601) );
  XNOR2_X1 U10942 ( .A(n6469), .B(n10114), .ZN(n8506) );
  INV_X1 U10943 ( .A(n8504), .ZN(n8505) );
  INV_X1 U10944 ( .A(n8507), .ZN(n8512) );
  NOR2_X1 U10945 ( .A1(n6887), .A2(n8509), .ZN(n8511) );
  INV_X1 U10946 ( .A(n8522), .ZN(n8517) );
  NAND2_X1 U10947 ( .A1(n8517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8518) );
  INV_X1 U10948 ( .A(n9245), .ZN(n8519) );
  NAND2_X1 U10949 ( .A1(n8519), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10913) );
  NAND2_X1 U10950 ( .A1(n8522), .A2(n8521), .ZN(n8528) );
  NAND2_X1 U10951 ( .A1(n8524), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8525) );
  MUX2_X1 U10952 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8525), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8527) );
  INV_X1 U10953 ( .A(n13828), .ZN(n9543) );
  INV_X1 U10954 ( .A(n8530), .ZN(n13492) );
  NAND2_X1 U10955 ( .A1(n10494), .A2(n10114), .ZN(n9713) );
  NAND2_X1 U10956 ( .A1(n9246), .A2(n9713), .ZN(n10358) );
  NAND4_X1 U10957 ( .A1(n10364), .A2(n14087), .A3(n13492), .A4(n10358), .ZN(
        n8531) );
  OAI211_X1 U10958 ( .C1(n13838), .C2(n10913), .A(n8531), .B(P1_B_REG_SCAN_IN), 
        .ZN(n8532) );
  NOR2_X2 U10959 ( .A1(n8533), .A2(P3_IR_REG_29__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U10960 ( .A1(n8533), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8534) );
  MUX2_X1 U10961 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8534), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8536) );
  INV_X1 U10962 ( .A(n8535), .ZN(n12639) );
  NAND2_X1 U10963 ( .A1(n12033), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8543) );
  NAND2_X1 U10964 ( .A1(n6458), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8542) );
  AND2_X2 U10965 ( .A1(n8538), .A2(n12648), .ZN(n8719) );
  NAND2_X1 U10966 ( .A1(n8922), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8541) );
  NAND2_X2 U10967 ( .A1(n8538), .A2(n8537), .ZN(n8606) );
  NOR2_X2 U10968 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8634) );
  NAND2_X1 U10969 ( .A1(n8634), .A2(n8633), .ZN(n8649) );
  NAND2_X1 U10970 ( .A1(n8739), .A2(n8738), .ZN(n8752) );
  AND2_X1 U10971 ( .A1(n8754), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8539) );
  NOR2_X1 U10972 ( .A1(n8767), .A2(n8539), .ZN(n12460) );
  OR2_X1 U10973 ( .A1(n8606), .A2(n12460), .ZN(n8540) );
  NAND2_X1 U10974 ( .A1(n8579), .A2(n8586), .ZN(n8545) );
  INV_X1 U10975 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9300) );
  NAND2_X1 U10976 ( .A1(n9300), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8544) );
  XNOR2_X1 U10977 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8598) );
  INV_X1 U10978 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9349) );
  NAND2_X1 U10979 ( .A1(n9349), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8546) );
  INV_X1 U10980 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8547) );
  NAND2_X1 U10981 ( .A1(n8547), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8548) );
  INV_X1 U10982 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n8550) );
  NAND2_X1 U10983 ( .A1(n8550), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10984 ( .A1(n8552), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8553) );
  NAND2_X1 U10985 ( .A1(n9186), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8555) );
  NAND2_X1 U10986 ( .A1(n8556), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8557) );
  NAND2_X1 U10987 ( .A1(n9191), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8558) );
  NAND2_X1 U10988 ( .A1(n8689), .A2(n8688), .ZN(n8560) );
  NAND2_X1 U10989 ( .A1(n9219), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8559) );
  NAND2_X1 U10990 ( .A1(n8561), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8562) );
  XNOR2_X1 U10991 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8713) );
  XNOR2_X1 U10992 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n8726) );
  NAND2_X1 U10993 ( .A1(n8564), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8565) );
  NAND2_X1 U10994 ( .A1(n8568), .A2(n8567), .ZN(n8569) );
  XNOR2_X1 U10995 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8746) );
  NAND2_X1 U10996 ( .A1(n8570), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U10997 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8760) );
  XNOR2_X1 U10998 ( .A(n8761), .B(n6678), .ZN(n9258) );
  AND2_X2 U10999 ( .A1(n8934), .A2(n9299), .ZN(n8611) );
  NAND2_X1 U11000 ( .A1(n9258), .A2(n12042), .ZN(n8574) );
  OAI22_X1 U11001 ( .A1(n8601), .A2(n9260), .B1(n8934), .B2(n9259), .ZN(n8572)
         );
  INV_X1 U11002 ( .A(n8572), .ZN(n8573) );
  NAND2_X1 U11003 ( .A1(n6457), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8578) );
  NAND2_X1 U11004 ( .A1(n8719), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U11005 ( .A1(n8593), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8576) );
  INV_X1 U11006 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n14786) );
  OR2_X1 U11007 ( .A1(n8606), .A2(n14786), .ZN(n8575) );
  AND4_X2 U11008 ( .A1(n8578), .A2(n8577), .A3(n8576), .A4(n8575), .ZN(n14763)
         );
  XNOR2_X1 U11009 ( .A(n8579), .B(n8586), .ZN(n9171) );
  NAND2_X1 U11010 ( .A1(n8611), .A2(n9171), .ZN(n8581) );
  OR2_X1 U11011 ( .A1(n8934), .A2(n9752), .ZN(n8580) );
  OAI211_X1 U11012 ( .C1(n8601), .C2(n9173), .A(n8581), .B(n8580), .ZN(n14781)
         );
  INV_X1 U11013 ( .A(n14781), .ZN(n14796) );
  NAND2_X1 U11014 ( .A1(n14763), .A2(n14781), .ZN(n12077) );
  NAND2_X1 U11015 ( .A1(n6458), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8585) );
  INV_X1 U11016 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9956) );
  OR2_X1 U11017 ( .A1(n8606), .A2(n9956), .ZN(n8584) );
  NAND2_X1 U11018 ( .A1(n8719), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8583) );
  NAND2_X1 U11019 ( .A1(n8593), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8582) );
  INV_X1 U11020 ( .A(n8586), .ZN(n8589) );
  NAND2_X1 U11021 ( .A1(n8587), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8588) );
  NAND2_X1 U11022 ( .A1(n8589), .A2(n8588), .ZN(n8590) );
  MUX2_X1 U11023 ( .A(n8590), .B(SI_0_), .S(n9154), .Z(n12666) );
  MUX2_X1 U11024 ( .A(P3_IR_REG_0__SCAN_IN), .B(n12666), .S(n8934), .Z(n10023)
         );
  NAND2_X1 U11025 ( .A1(n9945), .A2(n14776), .ZN(n8591) );
  NAND2_X1 U11026 ( .A1(n14763), .A2(n14796), .ZN(n9044) );
  NAND2_X1 U11027 ( .A1(n8591), .A2(n9044), .ZN(n14758) );
  NAND2_X1 U11028 ( .A1(n6457), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8597) );
  NAND2_X1 U11029 ( .A1(n8719), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8596) );
  NAND2_X1 U11030 ( .A1(n8593), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8595) );
  INV_X1 U11031 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10019) );
  OR2_X1 U11032 ( .A1(n8606), .A2(n10019), .ZN(n8594) );
  INV_X1 U11033 ( .A(n8598), .ZN(n8599) );
  XNOR2_X1 U11034 ( .A(n8600), .B(n8599), .ZN(n9218) );
  NAND2_X1 U11035 ( .A1(n8611), .A2(n9218), .ZN(n8604) );
  OR2_X1 U11036 ( .A1(n8601), .A2(SI_2_), .ZN(n8603) );
  OR2_X1 U11037 ( .A1(n8934), .A2(n9216), .ZN(n8602) );
  INV_X1 U11038 ( .A(n10013), .ZN(n14767) );
  NAND2_X1 U11039 ( .A1(n10463), .A2(n14767), .ZN(n8605) );
  NAND2_X1 U11040 ( .A1(n6458), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8610) );
  NAND2_X1 U11041 ( .A1(n8719), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8609) );
  NAND2_X1 U11042 ( .A1(n8593), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8608) );
  OR2_X1 U11043 ( .A1(n8606), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8607) );
  INV_X1 U11044 ( .A(n8612), .ZN(n8613) );
  XNOR2_X1 U11045 ( .A(n8614), .B(n8613), .ZN(n9206) );
  NAND2_X1 U11046 ( .A1(n12042), .A2(n9206), .ZN(n8617) );
  OR2_X1 U11047 ( .A1(n8601), .A2(SI_3_), .ZN(n8616) );
  OR2_X1 U11048 ( .A1(n8934), .A2(n9667), .ZN(n8615) );
  INV_X1 U11049 ( .A(n9054), .ZN(n10469) );
  NAND2_X1 U11050 ( .A1(n14761), .A2(n9054), .ZN(n12087) );
  INV_X1 U11051 ( .A(n12221), .ZN(n8618) );
  NAND2_X1 U11052 ( .A1(n10665), .A2(n9054), .ZN(n8619) );
  NAND2_X1 U11053 ( .A1(n10464), .A2(n8619), .ZN(n10667) );
  NAND2_X1 U11054 ( .A1(n6458), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8624) );
  INV_X2 U11055 ( .A(n8821), .ZN(n8922) );
  NAND2_X1 U11056 ( .A1(n8922), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8623) );
  NAND2_X1 U11057 ( .A1(n8593), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8622) );
  AND2_X1 U11058 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8620) );
  NOR2_X1 U11059 ( .A1(n8634), .A2(n8620), .ZN(n10664) );
  OR2_X1 U11060 ( .A1(n8606), .A2(n10664), .ZN(n8621) );
  INV_X1 U11061 ( .A(n8625), .ZN(n8626) );
  XNOR2_X1 U11062 ( .A(n8627), .B(n8626), .ZN(n9209) );
  NAND2_X1 U11063 ( .A1(n12042), .A2(n9209), .ZN(n8630) );
  OR2_X1 U11064 ( .A1(n12043), .A2(SI_4_), .ZN(n8629) );
  OR2_X1 U11065 ( .A1(n8934), .A2(n9776), .ZN(n8628) );
  AND3_X2 U11066 ( .A1(n8630), .A2(n8629), .A3(n8628), .ZN(n10663) );
  NAND2_X1 U11067 ( .A1(n10782), .A2(n10663), .ZN(n12094) );
  INV_X1 U11068 ( .A(n10663), .ZN(n8631) );
  NAND2_X1 U11069 ( .A1(n12278), .A2(n8631), .ZN(n12093) );
  NAND2_X1 U11070 ( .A1(n10667), .A2(n12088), .ZN(n10666) );
  NAND2_X1 U11071 ( .A1(n12278), .A2(n10663), .ZN(n8632) );
  NAND2_X1 U11072 ( .A1(n10666), .A2(n8632), .ZN(n10777) );
  INV_X1 U11073 ( .A(n10777), .ZN(n8646) );
  NAND2_X1 U11074 ( .A1(n12033), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8639) );
  NAND2_X1 U11075 ( .A1(n6458), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8638) );
  NAND2_X1 U11076 ( .A1(n8719), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8637) );
  OR2_X1 U11077 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  AND2_X1 U11078 ( .A1(n8649), .A2(n8635), .ZN(n10776) );
  OR2_X1 U11079 ( .A1(n8606), .A2(n10776), .ZN(n8636) );
  INV_X1 U11080 ( .A(n8640), .ZN(n8641) );
  XNOR2_X1 U11081 ( .A(n8642), .B(n8641), .ZN(n9212) );
  NAND2_X1 U11082 ( .A1(n12042), .A2(n9212), .ZN(n8645) );
  OR2_X1 U11083 ( .A1(n12043), .A2(SI_5_), .ZN(n8644) );
  OR2_X1 U11084 ( .A1(n8934), .A2(n7090), .ZN(n8643) );
  NAND2_X1 U11085 ( .A1(n10728), .A2(n10775), .ZN(n12097) );
  INV_X1 U11086 ( .A(n10728), .ZN(n12277) );
  INV_X1 U11087 ( .A(n10775), .ZN(n8647) );
  NAND2_X1 U11088 ( .A1(n12277), .A2(n8647), .ZN(n12101) );
  NAND2_X1 U11089 ( .A1(n10728), .A2(n8647), .ZN(n8648) );
  NAND2_X1 U11090 ( .A1(n6458), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8654) );
  NAND2_X1 U11091 ( .A1(n8719), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8653) );
  NAND2_X1 U11092 ( .A1(n12033), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8652) );
  NAND2_X1 U11093 ( .A1(n8649), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8650) );
  AND2_X1 U11094 ( .A1(n8659), .A2(n8650), .ZN(n14756) );
  OR2_X1 U11095 ( .A1(n8606), .A2(n14756), .ZN(n8651) );
  INV_X1 U11096 ( .A(SI_6_), .ZN(n9214) );
  XNOR2_X1 U11097 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8655) );
  XNOR2_X1 U11098 ( .A(n8656), .B(n8655), .ZN(n9213) );
  NAND2_X1 U11099 ( .A1(n12042), .A2(n9213), .ZN(n8658) );
  OR2_X1 U11100 ( .A1(n8934), .A2(n9931), .ZN(n8657) );
  OAI211_X1 U11101 ( .C1(n12043), .C2(n9214), .A(n8658), .B(n8657), .ZN(n14820) );
  NAND2_X1 U11102 ( .A1(n10781), .A2(n14820), .ZN(n12106) );
  INV_X1 U11103 ( .A(n14820), .ZN(n9064) );
  NAND2_X1 U11104 ( .A1(n12276), .A2(n9064), .ZN(n12103) );
  NAND2_X1 U11105 ( .A1(n12106), .A2(n12103), .ZN(n14748) );
  NAND2_X1 U11106 ( .A1(n6457), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8664) );
  AND2_X1 U11107 ( .A1(n8659), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8660) );
  NOR2_X1 U11108 ( .A1(n8670), .A2(n8660), .ZN(n14679) );
  OR2_X1 U11109 ( .A1(n8606), .A2(n14679), .ZN(n8663) );
  NAND2_X1 U11110 ( .A1(n12033), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8662) );
  NAND2_X1 U11111 ( .A1(n8922), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8661) );
  NAND4_X1 U11112 ( .A1(n8664), .A2(n8663), .A3(n8662), .A4(n8661), .ZN(n12107) );
  XNOR2_X1 U11113 ( .A(n8666), .B(n8665), .ZN(n9167) );
  NAND2_X1 U11114 ( .A1(n12042), .A2(n9167), .ZN(n8669) );
  OR2_X1 U11115 ( .A1(n8934), .A2(n8667), .ZN(n8668) );
  OAI211_X1 U11116 ( .C1(n12043), .C2(SI_7_), .A(n8669), .B(n8668), .ZN(n14826) );
  XNOR2_X1 U11117 ( .A(n12107), .B(n14826), .ZN(n12226) );
  NAND2_X1 U11118 ( .A1(n10825), .A2(n12226), .ZN(n10864) );
  INV_X1 U11119 ( .A(n14826), .ZN(n14676) );
  NAND2_X1 U11120 ( .A1(n12107), .A2(n14676), .ZN(n10863) );
  NAND2_X1 U11121 ( .A1(n12033), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8675) );
  NAND2_X1 U11122 ( .A1(n6458), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8674) );
  NAND2_X1 U11123 ( .A1(n8922), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8673) );
  NOR2_X1 U11124 ( .A1(n8670), .A2(n10033), .ZN(n8671) );
  OR2_X1 U11125 ( .A1(n8606), .A2(n7599), .ZN(n8672) );
  INV_X1 U11126 ( .A(SI_8_), .ZN(n9201) );
  XNOR2_X1 U11127 ( .A(n8676), .B(n6595), .ZN(n9200) );
  NAND2_X1 U11128 ( .A1(n12042), .A2(n9200), .ZN(n8678) );
  OR2_X1 U11129 ( .A1(n8934), .A2(n10034), .ZN(n8677) );
  OAI211_X1 U11130 ( .C1(n12043), .C2(n9201), .A(n8678), .B(n8677), .ZN(n10871) );
  NAND2_X1 U11131 ( .A1(n9071), .A2(n10871), .ZN(n12114) );
  INV_X1 U11132 ( .A(n10871), .ZN(n9070) );
  NAND2_X1 U11133 ( .A1(n12275), .A2(n9070), .ZN(n12113) );
  INV_X1 U11134 ( .A(n12222), .ZN(n8679) );
  AND2_X1 U11135 ( .A1(n10863), .A2(n8679), .ZN(n8680) );
  NAND2_X1 U11136 ( .A1(n9071), .A2(n9070), .ZN(n8681) );
  NAND2_X1 U11137 ( .A1(n6458), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8687) );
  NAND2_X1 U11138 ( .A1(n8719), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8686) );
  NAND2_X1 U11139 ( .A1(n12033), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8685) );
  OR2_X1 U11140 ( .A1(n8682), .A2(n9098), .ZN(n8683) );
  AND2_X1 U11141 ( .A1(n8693), .A2(n8683), .ZN(n10938) );
  OR2_X1 U11142 ( .A1(n8606), .A2(n10938), .ZN(n8684) );
  XNOR2_X1 U11143 ( .A(n8689), .B(n8688), .ZN(n9180) );
  NAND2_X1 U11144 ( .A1(n12042), .A2(n9180), .ZN(n8691) );
  OR2_X1 U11145 ( .A1(n8934), .A2(n14685), .ZN(n8690) );
  OAI211_X1 U11146 ( .C1(n12043), .C2(SI_9_), .A(n8691), .B(n8690), .ZN(n14836) );
  NAND2_X1 U11147 ( .A1(n11072), .A2(n14836), .ZN(n8692) );
  INV_X1 U11148 ( .A(n14836), .ZN(n12118) );
  NAND2_X1 U11149 ( .A1(n14732), .A2(n12118), .ZN(n12119) );
  NAND2_X1 U11150 ( .A1(n6457), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8698) );
  NAND2_X1 U11151 ( .A1(n8719), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8697) );
  NAND2_X1 U11152 ( .A1(n12033), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8696) );
  NAND2_X1 U11153 ( .A1(n8693), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8694) );
  AND2_X1 U11154 ( .A1(n8707), .A2(n8694), .ZN(n14741) );
  OR2_X1 U11155 ( .A1(n8606), .A2(n14741), .ZN(n8695) );
  XNOR2_X1 U11156 ( .A(n8700), .B(n8699), .ZN(n9204) );
  NAND2_X1 U11157 ( .A1(n12042), .A2(n9204), .ZN(n8704) );
  OR2_X1 U11158 ( .A1(n8934), .A2(n8701), .ZN(n8703) );
  OR2_X1 U11159 ( .A1(n12043), .A2(SI_10_), .ZN(n8702) );
  NAND2_X1 U11160 ( .A1(n11051), .A2(n14725), .ZN(n12123) );
  INV_X1 U11161 ( .A(n14725), .ZN(n8705) );
  NAND2_X1 U11162 ( .A1(n12274), .A2(n8705), .ZN(n12124) );
  NAND2_X1 U11163 ( .A1(n12123), .A2(n12124), .ZN(n14735) );
  NAND2_X1 U11164 ( .A1(n14728), .A2(n14735), .ZN(n14727) );
  NAND2_X1 U11165 ( .A1(n12274), .A2(n14725), .ZN(n8706) );
  NAND2_X1 U11166 ( .A1(n14727), .A2(n8706), .ZN(n11050) );
  INV_X1 U11167 ( .A(n11050), .ZN(n8718) );
  NAND2_X1 U11168 ( .A1(n12033), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11169 ( .A1(n8707), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8708) );
  AND2_X1 U11170 ( .A1(n8720), .A2(n8708), .ZN(n11055) );
  OR2_X1 U11171 ( .A1(n8606), .A2(n11055), .ZN(n8711) );
  NAND2_X1 U11172 ( .A1(n6457), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8710) );
  NAND2_X1 U11173 ( .A1(n8719), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8709) );
  NAND4_X1 U11174 ( .A1(n8712), .A2(n8711), .A3(n8710), .A4(n8709), .ZN(n14729) );
  XNOR2_X1 U11175 ( .A(n8714), .B(n8713), .ZN(n9176) );
  NAND2_X1 U11176 ( .A1(n12042), .A2(n9176), .ZN(n8717) );
  OR2_X1 U11177 ( .A1(n12043), .A2(SI_11_), .ZN(n8716) );
  OR2_X1 U11178 ( .A1(n8934), .A2(n10682), .ZN(n8715) );
  INV_X1 U11179 ( .A(n11212), .ZN(n8974) );
  NAND2_X1 U11180 ( .A1(n12033), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U11181 ( .A1(n6458), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U11182 ( .A1(n8719), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8723) );
  AND2_X1 U11183 ( .A1(n8720), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8721) );
  NOR2_X1 U11184 ( .A1(n8739), .A2(n8721), .ZN(n11937) );
  OR2_X1 U11185 ( .A1(n8606), .A2(n11937), .ZN(n8722) );
  INV_X1 U11186 ( .A(n8726), .ZN(n8727) );
  XNOR2_X1 U11187 ( .A(n8728), .B(n8727), .ZN(n9197) );
  NAND2_X1 U11188 ( .A1(n9197), .A2(n12042), .ZN(n8731) );
  OAI22_X1 U11189 ( .A1(n8601), .A2(n9198), .B1(n8934), .B2(n10633), .ZN(n8729) );
  INV_X1 U11190 ( .A(n8729), .ZN(n8730) );
  NAND2_X1 U11191 ( .A1(n8731), .A2(n8730), .ZN(n11941) );
  NAND2_X1 U11192 ( .A1(n11985), .A2(n11941), .ZN(n12135) );
  INV_X1 U11193 ( .A(n11941), .ZN(n11226) );
  NAND2_X1 U11194 ( .A1(n12273), .A2(n11226), .ZN(n12132) );
  NAND2_X1 U11195 ( .A1(n12135), .A2(n12132), .ZN(n12232) );
  NAND2_X1 U11196 ( .A1(n12273), .A2(n11941), .ZN(n8732) );
  XNOR2_X1 U11197 ( .A(n8733), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n9224) );
  NAND2_X1 U11198 ( .A1(n9224), .A2(n12042), .ZN(n8737) );
  OAI22_X1 U11199 ( .A1(n12043), .A2(SI_13_), .B1(n8734), .B2(n8934), .ZN(
        n8735) );
  INV_X1 U11200 ( .A(n8735), .ZN(n8736) );
  NAND2_X1 U11201 ( .A1(n12033), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8744) );
  NAND2_X1 U11202 ( .A1(n6458), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U11203 ( .A1(n8922), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8742) );
  OR2_X1 U11204 ( .A1(n8739), .A2(n8738), .ZN(n8740) );
  AND2_X1 U11205 ( .A1(n8740), .A2(n8752), .ZN(n12487) );
  OR2_X1 U11206 ( .A1(n8606), .A2(n12487), .ZN(n8741) );
  OR2_X1 U11207 ( .A1(n12634), .A2(n12469), .ZN(n8745) );
  XNOR2_X1 U11208 ( .A(n8747), .B(n8746), .ZN(n9227) );
  NAND2_X1 U11209 ( .A1(n9227), .A2(n12042), .ZN(n8751) );
  INV_X1 U11210 ( .A(n11084), .ZN(n8748) );
  OAI22_X1 U11211 ( .A1(n8601), .A2(SI_14_), .B1(n8748), .B2(n8934), .ZN(n8749) );
  INV_X1 U11212 ( .A(n8749), .ZN(n8750) );
  NAND2_X1 U11213 ( .A1(n8751), .A2(n8750), .ZN(n12623) );
  NAND2_X1 U11214 ( .A1(n12033), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8758) );
  NAND2_X1 U11215 ( .A1(n8752), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8753) );
  AND2_X1 U11216 ( .A1(n8754), .A2(n8753), .ZN(n12478) );
  OR2_X1 U11217 ( .A1(n8606), .A2(n12478), .ZN(n8757) );
  NAND2_X1 U11218 ( .A1(n6457), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8756) );
  NAND2_X1 U11219 ( .A1(n8922), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8755) );
  NAND4_X1 U11220 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n12272) );
  OR2_X1 U11221 ( .A1(n12623), .A2(n12272), .ZN(n12152) );
  NAND2_X1 U11222 ( .A1(n12623), .A2(n12272), .ZN(n12145) );
  NAND2_X1 U11223 ( .A1(n12152), .A2(n12145), .ZN(n12464) );
  INV_X1 U11224 ( .A(n12272), .ZN(n11894) );
  OR2_X1 U11225 ( .A1(n12623), .A2(n11894), .ZN(n8759) );
  NAND2_X1 U11226 ( .A1(n12467), .A2(n8759), .ZN(n12455) );
  XNOR2_X1 U11227 ( .A(n12616), .B(n12468), .ZN(n12454) );
  XNOR2_X1 U11228 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n8775) );
  INV_X1 U11229 ( .A(n8775), .ZN(n8762) );
  XNOR2_X1 U11230 ( .A(n8774), .B(n8762), .ZN(n9386) );
  NAND2_X1 U11231 ( .A1(n9386), .A2(n12042), .ZN(n8765) );
  OAI22_X1 U11232 ( .A1(n8601), .A2(n9387), .B1(n8934), .B2(n9388), .ZN(n8763)
         );
  INV_X1 U11233 ( .A(n8763), .ZN(n8764) );
  NAND2_X1 U11234 ( .A1(n12033), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U11235 ( .A1(n6458), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8771) );
  NAND2_X1 U11236 ( .A1(n8922), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8770) );
  INV_X1 U11237 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8766) );
  NOR2_X1 U11238 ( .A1(n8767), .A2(n8766), .ZN(n8768) );
  OR2_X1 U11239 ( .A1(n8791), .A2(n8768), .ZN(n12448) );
  INV_X1 U11240 ( .A(n12448), .ZN(n11956) );
  OR2_X1 U11241 ( .A1(n8606), .A2(n11956), .ZN(n8769) );
  NAND2_X1 U11242 ( .A1(n12154), .A2(n12018), .ZN(n8773) );
  AOI22_X1 U11243 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n9834), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9793), .ZN(n8782) );
  XOR2_X1 U11244 ( .A(n8781), .B(n8782), .Z(n9590) );
  INV_X1 U11245 ( .A(SI_17_), .ZN(n9592) );
  OAI22_X1 U11246 ( .A1(n8601), .A2(n9592), .B1(n8934), .B2(n9591), .ZN(n8776)
         );
  NAND2_X1 U11247 ( .A1(n12033), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8780) );
  XNOR2_X1 U11248 ( .A(n8791), .B(P3_REG3_REG_17__SCAN_IN), .ZN(n12436) );
  OR2_X1 U11249 ( .A1(n8606), .A2(n12436), .ZN(n8779) );
  NAND2_X1 U11250 ( .A1(n6457), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8778) );
  NAND2_X1 U11251 ( .A1(n8922), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8777) );
  NAND4_X1 U11252 ( .A1(n8780), .A2(n8779), .A3(n8778), .A4(n8777), .ZN(n12271) );
  NAND2_X1 U11253 ( .A1(n11969), .A2(n12271), .ZN(n12060) );
  INV_X1 U11254 ( .A(n11969), .ZN(n12603) );
  NAND2_X1 U11255 ( .A1(n12603), .A2(n12419), .ZN(n8977) );
  INV_X1 U11256 ( .A(n12416), .ZN(n8798) );
  NAND2_X1 U11257 ( .A1(n9793), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8783) );
  XNOR2_X1 U11258 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .ZN(n8801) );
  INV_X1 U11259 ( .A(n8801), .ZN(n8784) );
  XNOR2_X1 U11260 ( .A(n8800), .B(n8784), .ZN(n13949) );
  NAND2_X1 U11261 ( .A1(n13949), .A2(n12042), .ZN(n8788) );
  INV_X1 U11262 ( .A(SI_18_), .ZN(n8785) );
  OAI22_X1 U11263 ( .A1(n12043), .A2(n8785), .B1(n8934), .B2(n13951), .ZN(
        n8786) );
  INV_X1 U11264 ( .A(n8786), .ZN(n8787) );
  NAND2_X1 U11265 ( .A1(n12033), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8790) );
  NAND2_X1 U11266 ( .A1(n6458), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8789) );
  NAND2_X1 U11267 ( .A1(n8790), .A2(n8789), .ZN(n8796) );
  NAND2_X1 U11268 ( .A1(n8792), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8793) );
  AND2_X1 U11269 ( .A1(n8805), .A2(n8793), .ZN(n12421) );
  NAND2_X1 U11270 ( .A1(n8922), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8794) );
  OAI21_X1 U11271 ( .B1(n12421), .B2(n8606), .A(n8794), .ZN(n8795) );
  NAND2_X1 U11272 ( .A1(n12427), .A2(n11964), .ZN(n12062) );
  NAND2_X1 U11273 ( .A1(n12600), .A2(n11964), .ZN(n8799) );
  AOI22_X1 U11274 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10113), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n7326), .ZN(n8814) );
  XNOR2_X1 U11275 ( .A(n8813), .B(n8814), .ZN(n9758) );
  NAND2_X1 U11276 ( .A1(n9758), .A2(n12042), .ZN(n8804) );
  INV_X1 U11277 ( .A(n12055), .ZN(n12245) );
  OAI22_X1 U11278 ( .A1(n12043), .A2(SI_19_), .B1(n12245), .B2(n8934), .ZN(
        n8802) );
  INV_X1 U11279 ( .A(n8802), .ZN(n8803) );
  AND2_X1 U11280 ( .A1(n8805), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8806) );
  OR2_X1 U11281 ( .A1(n8806), .A2(n8817), .ZN(n12410) );
  NAND2_X1 U11282 ( .A1(n12410), .A2(n8851), .ZN(n8811) );
  NAND2_X1 U11283 ( .A1(n12033), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8808) );
  NAND2_X1 U11284 ( .A1(n6458), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n8807) );
  AND2_X1 U11285 ( .A1(n8808), .A2(n8807), .ZN(n8810) );
  NAND2_X1 U11286 ( .A1(n8922), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8809) );
  NAND2_X1 U11287 ( .A1(n12593), .A2(n12420), .ZN(n8812) );
  INV_X1 U11288 ( .A(n12593), .ZN(n12411) );
  XNOR2_X1 U11289 ( .A(n8823), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U11290 ( .A1(n10109), .A2(n12042), .ZN(n8816) );
  OR2_X1 U11291 ( .A1(n8601), .A2(n10110), .ZN(n8815) );
  INV_X1 U11292 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12398) );
  INV_X1 U11293 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n11973) );
  NOR2_X1 U11294 ( .A1(n8817), .A2(n11973), .ZN(n8818) );
  OR2_X1 U11295 ( .A1(n8828), .A2(n8818), .ZN(n12399) );
  NAND2_X1 U11296 ( .A1(n12399), .A2(n8851), .ZN(n8820) );
  AOI22_X1 U11297 ( .A1(n6457), .A2(P3_REG1_REG_20__SCAN_IN), .B1(n12033), 
        .B2(P3_REG0_REG_20__SCAN_IN), .ZN(n8819) );
  OAI211_X1 U11298 ( .C1(n8821), .C2(n12398), .A(n8820), .B(n8819), .ZN(n12269) );
  INV_X1 U11299 ( .A(n12269), .ZN(n12383) );
  NAND2_X1 U11300 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8822), .ZN(n8824) );
  INV_X1 U11301 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U11302 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11465), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n11871), .ZN(n8834) );
  INV_X1 U11303 ( .A(n8834), .ZN(n8825) );
  XNOR2_X1 U11304 ( .A(n8833), .B(n8825), .ZN(n10222) );
  NAND2_X1 U11305 ( .A1(n10222), .A2(n12042), .ZN(n8827) );
  INV_X1 U11306 ( .A(SI_21_), .ZN(n10224) );
  OR2_X1 U11307 ( .A1(n12043), .A2(n10224), .ZN(n8826) );
  INV_X1 U11308 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n11929) );
  OR2_X1 U11309 ( .A1(n8828), .A2(n11929), .ZN(n8829) );
  NAND2_X1 U11310 ( .A1(n8837), .A2(n8829), .ZN(n12387) );
  NAND2_X1 U11311 ( .A1(n12387), .A2(n8851), .ZN(n8832) );
  AOI22_X1 U11312 ( .A1(n6457), .A2(P3_REG1_REG_21__SCAN_IN), .B1(n8593), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8831) );
  NAND2_X1 U11313 ( .A1(n8922), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8830) );
  INV_X1 U11314 ( .A(n12396), .ZN(n12268) );
  INV_X1 U11315 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U11316 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11487), .B2(n14899), .ZN(n8845) );
  XNOR2_X1 U11317 ( .A(n8846), .B(n8845), .ZN(n10347) );
  NAND2_X1 U11318 ( .A1(n10347), .A2(n12042), .ZN(n8836) );
  OR2_X1 U11319 ( .A1(n8601), .A2(n6953), .ZN(n8835) );
  NAND2_X1 U11320 ( .A1(n8837), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8838) );
  NAND2_X1 U11321 ( .A1(n8849), .A2(n8838), .ZN(n12375) );
  NAND2_X1 U11322 ( .A1(n12375), .A2(n8851), .ZN(n8843) );
  NAND2_X1 U11323 ( .A1(n8922), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8841) );
  NAND2_X1 U11324 ( .A1(n12033), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8840) );
  NAND2_X1 U11325 ( .A1(n6458), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8839) );
  AND3_X1 U11326 ( .A1(n8841), .A2(n8840), .A3(n8839), .ZN(n8842) );
  INV_X1 U11327 ( .A(n12578), .ZN(n8844) );
  INV_X1 U11328 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10915) );
  AOI22_X1 U11329 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11500), .B2(n10915), .ZN(n8857) );
  XNOR2_X1 U11330 ( .A(n8858), .B(n8857), .ZN(n10643) );
  NAND2_X1 U11331 ( .A1(n10643), .A2(n12042), .ZN(n8848) );
  INV_X1 U11332 ( .A(SI_23_), .ZN(n10645) );
  NAND2_X1 U11333 ( .A1(n8849), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U11334 ( .A1(n8850), .A2(n7601), .ZN(n12366) );
  NAND2_X1 U11335 ( .A1(n12366), .A2(n8851), .ZN(n8856) );
  NAND2_X1 U11336 ( .A1(n8922), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U11337 ( .A1(n6458), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U11338 ( .A1(n12033), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8852) );
  AND3_X1 U11339 ( .A1(n8854), .A2(n8853), .A3(n8852), .ZN(n8855) );
  XNOR2_X1 U11340 ( .A(n12572), .B(n12178), .ZN(n12239) );
  INV_X1 U11341 ( .A(n12178), .ZN(n12267) );
  INV_X1 U11342 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11122) );
  XOR2_X1 U11343 ( .A(n11122), .B(n8865), .Z(n11279) );
  INV_X1 U11344 ( .A(SI_24_), .ZN(n11281) );
  NAND2_X1 U11345 ( .A1(n12033), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8862) );
  AOI21_X1 U11346 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(n7601), .A(n8871), .ZN(
        n12352) );
  OR2_X1 U11347 ( .A1(n8606), .A2(n12352), .ZN(n8861) );
  NAND2_X1 U11348 ( .A1(n6458), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U11349 ( .A1(n8922), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8859) );
  NAND4_X1 U11350 ( .A1(n8862), .A2(n8861), .A3(n8860), .A4(n8859), .ZN(n12362) );
  NAND2_X1 U11351 ( .A1(n11273), .A2(n12362), .ZN(n8863) );
  AOI22_X1 U11352 ( .A1(n12346), .A2(n8863), .B1(n11906), .B2(n12569), .ZN(
        n12336) );
  NAND2_X1 U11353 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8864), .ZN(n8866) );
  AOI22_X1 U11354 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13211), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n11276), .ZN(n8867) );
  INV_X1 U11355 ( .A(n8867), .ZN(n8868) );
  XNOR2_X1 U11356 ( .A(n8879), .B(n8868), .ZN(n11095) );
  NAND2_X1 U11357 ( .A1(n11095), .A2(n12042), .ZN(n8870) );
  NAND2_X1 U11358 ( .A1(n6457), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8877) );
  AND2_X1 U11359 ( .A1(P3_REG3_REG_25__SCAN_IN), .A2(n8872), .ZN(n8873) );
  NOR2_X1 U11360 ( .A1(n8883), .A2(n8873), .ZN(n12341) );
  OR2_X1 U11361 ( .A1(n8606), .A2(n12341), .ZN(n8876) );
  NAND2_X1 U11362 ( .A1(n8922), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U11363 ( .A1(n12033), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8874) );
  NAND4_X1 U11364 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n12266) );
  XNOR2_X1 U11365 ( .A(n12343), .B(n12266), .ZN(n12242) );
  NAND2_X1 U11366 ( .A1(n12336), .A2(n12335), .ZN(n12334) );
  INV_X1 U11367 ( .A(n12343), .ZN(n12562) );
  NAND2_X1 U11368 ( .A1(n12334), .A2(n7596), .ZN(n12322) );
  NAND2_X1 U11369 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13211), .ZN(n8878) );
  AOI22_X1 U11370 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n13834), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n6922), .ZN(n8890) );
  XNOR2_X1 U11371 ( .A(n8891), .B(n8890), .ZN(n12660) );
  NAND2_X1 U11372 ( .A1(n12660), .A2(n8611), .ZN(n8881) );
  INV_X1 U11373 ( .A(n12500), .ZN(n12330) );
  NAND2_X1 U11374 ( .A1(n12033), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8888) );
  NAND2_X1 U11375 ( .A1(n6457), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8887) );
  NAND2_X1 U11376 ( .A1(n8922), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8886) );
  INV_X1 U11377 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n8882) );
  OR2_X1 U11378 ( .A1(n8883), .A2(n8882), .ZN(n8884) );
  NAND2_X1 U11379 ( .A1(n8883), .A2(n8882), .ZN(n8896) );
  AND2_X1 U11380 ( .A1(n8884), .A2(n8896), .ZN(n12327) );
  OR2_X1 U11381 ( .A1(n8606), .A2(n12327), .ZN(n8885) );
  NAND2_X1 U11382 ( .A1(n12330), .A2(n12314), .ZN(n8889) );
  NAND2_X1 U11383 ( .A1(n12500), .A2(n12314), .ZN(n12194) );
  INV_X1 U11384 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13205) );
  INV_X1 U11385 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n13831) );
  AOI22_X1 U11386 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(
        P1_DATAO_REG_27__SCAN_IN), .B1(n13205), .B2(n13831), .ZN(n8892) );
  INV_X1 U11387 ( .A(n8892), .ZN(n8893) );
  XNOR2_X1 U11388 ( .A(n8905), .B(n8893), .ZN(n12655) );
  NAND2_X1 U11389 ( .A1(n12655), .A2(n12042), .ZN(n8895) );
  INV_X1 U11390 ( .A(SI_27_), .ZN(n12658) );
  NAND2_X1 U11391 ( .A1(n12033), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8901) );
  NAND2_X1 U11392 ( .A1(n6458), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8900) );
  NAND2_X1 U11393 ( .A1(n8719), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11394 ( .A1(n8896), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8897) );
  AND2_X1 U11395 ( .A1(n8911), .A2(n8897), .ZN(n11888) );
  OR2_X1 U11396 ( .A1(n12497), .A2(n12009), .ZN(n12197) );
  NAND2_X1 U11397 ( .A1(n12497), .A2(n12009), .ZN(n12199) );
  NAND2_X2 U11398 ( .A1(n12197), .A2(n12199), .ZN(n12310) );
  NAND2_X1 U11399 ( .A1(n12313), .A2(n12310), .ZN(n8904) );
  NOR2_X1 U11400 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n13831), .ZN(n8906) );
  AOI22_X1 U11401 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n11552), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n13830), .ZN(n8907) );
  INV_X1 U11402 ( .A(n8907), .ZN(n8908) );
  NAND2_X1 U11403 ( .A1(n12651), .A2(n12042), .ZN(n8910) );
  NAND2_X1 U11404 ( .A1(n8593), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11405 ( .A1(n6457), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U11406 ( .A1(n8719), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8914) );
  AND2_X1 U11407 ( .A1(n8911), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8912) );
  NOR2_X1 U11408 ( .A1(n14050), .A2(n8912), .ZN(n12306) );
  OR2_X1 U11409 ( .A1(n8606), .A2(n12306), .ZN(n8913) );
  NAND2_X1 U11410 ( .A1(n12552), .A2(n12316), .ZN(n12200) );
  INV_X1 U11411 ( .A(n12316), .ZN(n12263) );
  NAND2_X1 U11412 ( .A1(n12552), .A2(n12263), .ZN(n8918) );
  NAND2_X1 U11413 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n11552), .ZN(n8920) );
  OAI22_X1 U11414 ( .A1(n14963), .A2(n13825), .B1(P2_DATAO_REG_29__SCAN_IN), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12026) );
  INV_X1 U11415 ( .A(n14050), .ZN(n8921) );
  NAND2_X1 U11416 ( .A1(n6458), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8925) );
  NAND2_X1 U11417 ( .A1(n8922), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11418 ( .A1(n12033), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8923) );
  NAND4_X1 U11419 ( .A1(n12037), .A2(n8925), .A3(n8924), .A4(n8923), .ZN(
        n12262) );
  INV_X1 U11420 ( .A(n12262), .ZN(n8926) );
  XNOR2_X1 U11421 ( .A(n8927), .B(n12241), .ZN(n8930) );
  NAND2_X1 U11422 ( .A1(n12245), .A2(n12256), .ZN(n9006) );
  NAND2_X1 U11423 ( .A1(n6481), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8928) );
  MUX2_X1 U11424 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8928), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8929) );
  NAND2_X1 U11425 ( .A1(n9041), .A2(n8994), .ZN(n12212) );
  NAND2_X1 U11426 ( .A1(n8930), .A2(n14778), .ZN(n8940) );
  NAND2_X1 U11427 ( .A1(n6458), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8933) );
  NAND2_X1 U11428 ( .A1(n8719), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8932) );
  NAND2_X1 U11429 ( .A1(n8593), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8931) );
  NAND4_X1 U11430 ( .A1(n12037), .A2(n8933), .A3(n8932), .A4(n8931), .ZN(
        n12261) );
  NAND2_X1 U11431 ( .A1(n8935), .A2(n8934), .ZN(n8936) );
  INV_X1 U11432 ( .A(P3_B_REG_SCAN_IN), .ZN(n8937) );
  NOR2_X1 U11433 ( .A1(n12654), .A2(n8937), .ZN(n8938) );
  NOR2_X1 U11434 ( .A1(n14760), .A2(n8938), .ZN(n14048) );
  AOI22_X1 U11435 ( .A1(n14731), .A2(n12263), .B1(n12261), .B2(n14048), .ZN(
        n8939) );
  NAND2_X1 U11436 ( .A1(n8940), .A2(n8939), .ZN(n9011) );
  XNOR2_X1 U11437 ( .A(n11282), .B(P3_B_REG_SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11438 ( .A1(n8941), .A2(n11098), .ZN(n8942) );
  OR2_X1 U11439 ( .A1(n8946), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8945) );
  NAND2_X1 U11440 ( .A1(n12665), .A2(n11098), .ZN(n8944) );
  NAND2_X1 U11441 ( .A1(n11282), .A2(n12665), .ZN(n8947) );
  XNOR2_X1 U11442 ( .A(n12637), .B(n9040), .ZN(n8960) );
  NOR2_X1 U11443 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .ZN(
        n8951) );
  NOR4_X1 U11444 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_17__SCAN_IN), .A4(P3_D_REG_25__SCAN_IN), .ZN(n8950) );
  NOR4_X1 U11445 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_29__SCAN_IN), .A3(
        P3_D_REG_10__SCAN_IN), .A4(P3_D_REG_31__SCAN_IN), .ZN(n8949) );
  NOR4_X1 U11446 ( .A1(P3_D_REG_20__SCAN_IN), .A2(P3_D_REG_19__SCAN_IN), .A3(
        P3_D_REG_18__SCAN_IN), .A4(P3_D_REG_27__SCAN_IN), .ZN(n8948) );
  NAND4_X1 U11447 ( .A1(n8951), .A2(n8950), .A3(n8949), .A4(n8948), .ZN(n8957)
         );
  NOR4_X1 U11448 ( .A1(P3_D_REG_26__SCAN_IN), .A2(P3_D_REG_9__SCAN_IN), .A3(
        P3_D_REG_16__SCAN_IN), .A4(P3_D_REG_15__SCAN_IN), .ZN(n8955) );
  NOR4_X1 U11449 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_21__SCAN_IN), .A4(P3_D_REG_11__SCAN_IN), .ZN(n8954) );
  NOR4_X1 U11450 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8953) );
  NOR4_X1 U11451 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8952) );
  NAND4_X1 U11452 ( .A1(n8955), .A2(n8954), .A3(n8953), .A4(n8952), .ZN(n8956)
         );
  NOR2_X1 U11453 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  OR2_X1 U11454 ( .A1(n8946), .A2(n8958), .ZN(n9005) );
  AND2_X1 U11455 ( .A1(n9005), .A2(n12253), .ZN(n8959) );
  NOR2_X1 U11456 ( .A1(n12068), .A2(n10112), .ZN(n8961) );
  NAND2_X1 U11457 ( .A1(n8961), .A2(n12055), .ZN(n8984) );
  NAND2_X1 U11458 ( .A1(n8984), .A2(n12183), .ZN(n8962) );
  NAND2_X2 U11459 ( .A1(n12055), .A2(n10112), .ZN(n12254) );
  NAND2_X1 U11460 ( .A1(n12254), .A2(n12076), .ZN(n9083) );
  AND2_X1 U11461 ( .A1(n8962), .A2(n9083), .ZN(n8997) );
  NAND2_X1 U11462 ( .A1(n12637), .A2(n8962), .ZN(n8963) );
  OAI21_X1 U11463 ( .B1(n12637), .B2(n8997), .A(n8963), .ZN(n8964) );
  INV_X1 U11464 ( .A(n8964), .ZN(n8965) );
  NAND2_X1 U11465 ( .A1(n8999), .A2(n8965), .ZN(n8987) );
  AND2_X1 U11466 ( .A1(n14769), .A2(n14821), .ZN(n8966) );
  MUX2_X1 U11467 ( .A(P3_REG2_REG_29__SCAN_IN), .B(n9011), .S(n14791), .Z(
        n8967) );
  INV_X1 U11468 ( .A(n8967), .ZN(n8992) );
  INV_X1 U11469 ( .A(n10023), .ZN(n9952) );
  NAND2_X1 U11470 ( .A1(n9048), .A2(n12077), .ZN(n14757) );
  INV_X1 U11471 ( .A(n14759), .ZN(n8968) );
  INV_X1 U11472 ( .A(n12088), .ZN(n12219) );
  INV_X1 U11473 ( .A(n14748), .ZN(n14742) );
  NAND2_X1 U11474 ( .A1(n14745), .A2(n12106), .ZN(n10824) );
  INV_X1 U11475 ( .A(n12226), .ZN(n12105) );
  NAND2_X1 U11476 ( .A1(n10824), .A2(n12105), .ZN(n8969) );
  INV_X1 U11477 ( .A(n12107), .ZN(n10839) );
  NAND2_X1 U11478 ( .A1(n10839), .A2(n14676), .ZN(n12109) );
  NAND2_X1 U11479 ( .A1(n8969), .A2(n12109), .ZN(n10862) );
  NAND2_X1 U11480 ( .A1(n10862), .A2(n12222), .ZN(n8970) );
  NOR2_X1 U11481 ( .A1(n14732), .A2(n14836), .ZN(n8971) );
  NAND2_X1 U11482 ( .A1(n14732), .A2(n14836), .ZN(n8972) );
  INV_X1 U11483 ( .A(n12124), .ZN(n8973) );
  NAND2_X1 U11484 ( .A1(n11236), .A2(n11212), .ZN(n12126) );
  NAND2_X1 U11485 ( .A1(n14729), .A2(n8974), .ZN(n12130) );
  INV_X1 U11486 ( .A(n12232), .ZN(n8975) );
  INV_X1 U11487 ( .A(n12152), .ZN(n8976) );
  NAND2_X1 U11488 ( .A1(n12616), .A2(n12468), .ZN(n12150) );
  OAI21_X1 U11489 ( .B1(n12452), .B2(n12454), .A(n12150), .ZN(n12441) );
  XNOR2_X1 U11490 ( .A(n12609), .B(n12433), .ZN(n12443) );
  NAND2_X1 U11491 ( .A1(n12609), .A2(n12018), .ZN(n12151) );
  INV_X1 U11492 ( .A(n8977), .ZN(n12058) );
  INV_X1 U11493 ( .A(n12393), .ZN(n12391) );
  NAND2_X1 U11494 ( .A1(n12588), .A2(n12269), .ZN(n12165) );
  NOR2_X1 U11495 ( .A1(n12388), .A2(n12396), .ZN(n12170) );
  NAND2_X1 U11496 ( .A1(n12388), .A2(n12396), .ZN(n12164) );
  NAND2_X1 U11497 ( .A1(n12569), .A2(n12362), .ZN(n8978) );
  NAND2_X1 U11498 ( .A1(n11273), .A2(n11906), .ZN(n12184) );
  INV_X1 U11499 ( .A(n12193), .ZN(n8979) );
  INV_X1 U11500 ( .A(n12199), .ZN(n8980) );
  NAND2_X1 U11501 ( .A1(n14769), .A2(n9041), .ZN(n14770) );
  INV_X1 U11502 ( .A(n12254), .ZN(n9095) );
  NOR2_X1 U11503 ( .A1(n9041), .A2(n8994), .ZN(n8981) );
  XNOR2_X1 U11504 ( .A(n8981), .B(n12068), .ZN(n8983) );
  NAND2_X1 U11505 ( .A1(n12055), .A2(n12069), .ZN(n8982) );
  NAND2_X1 U11506 ( .A1(n8983), .A2(n8982), .ZN(n9085) );
  NAND3_X1 U11507 ( .A1(n9095), .A2(n9085), .A3(n14837), .ZN(n8985) );
  INV_X1 U11508 ( .A(n14843), .ZN(n14783) );
  OR2_X1 U11509 ( .A1(n8987), .A2(n14769), .ZN(n10873) );
  AOI22_X1 U11510 ( .A1(n8988), .A2(n6433), .B1(n14772), .B2(n14050), .ZN(
        n8989) );
  OAI21_X1 U11511 ( .B1(n9014), .B2(n12493), .A(n8989), .ZN(n8990) );
  INV_X1 U11512 ( .A(n8990), .ZN(n8991) );
  NAND2_X1 U11513 ( .A1(n8992), .A2(n8991), .ZN(P3_U3204) );
  NAND2_X1 U11514 ( .A1(n12055), .A2(n12256), .ZN(n8993) );
  OAI21_X1 U11515 ( .B1(n14837), .B2(n8994), .A(n8993), .ZN(n8995) );
  AOI21_X1 U11516 ( .B1(n8995), .B2(n12254), .A(n12076), .ZN(n8996) );
  MUX2_X1 U11517 ( .A(n8997), .B(n8996), .S(n9004), .Z(n8998) );
  MUX2_X1 U11518 ( .A(P3_REG1_REG_29__SCAN_IN), .B(n9011), .S(n14868), .Z(
        n9000) );
  INV_X1 U11519 ( .A(n9000), .ZN(n9003) );
  INV_X1 U11520 ( .A(n9001), .ZN(n9002) );
  NAND2_X1 U11521 ( .A1(n9003), .A2(n9002), .ZN(P3_U3488) );
  NAND3_X1 U11522 ( .A1(n9004), .A2(n9040), .A3(n9005), .ZN(n9097) );
  INV_X1 U11523 ( .A(n9085), .ZN(n9009) );
  INV_X1 U11524 ( .A(n9040), .ZN(n9241) );
  NAND3_X1 U11525 ( .A1(n9241), .A2(n12637), .A3(n9005), .ZN(n9091) );
  INV_X1 U11526 ( .A(n9006), .ZN(n9007) );
  NOR2_X1 U11527 ( .A1(n9041), .A2(n10112), .ZN(n9039) );
  NAND2_X1 U11528 ( .A1(n9007), .A2(n9039), .ZN(n9086) );
  NAND2_X1 U11529 ( .A1(n9095), .A2(n12076), .ZN(n9940) );
  AND2_X1 U11530 ( .A1(n9086), .A2(n9940), .ZN(n9008) );
  OAI22_X1 U11531 ( .A1(n9097), .A2(n9009), .B1(n9091), .B2(n9008), .ZN(n9010)
         );
  MUX2_X1 U11532 ( .A(P3_REG0_REG_29__SCAN_IN), .B(n9011), .S(n14851), .Z(
        n9012) );
  INV_X1 U11533 ( .A(n9012), .ZN(n9017) );
  OAI22_X1 U11534 ( .A1(n9014), .A2(n12622), .B1(n9013), .B2(n12635), .ZN(
        n9015) );
  INV_X1 U11535 ( .A(n9015), .ZN(n9016) );
  NAND2_X1 U11536 ( .A1(n9017), .A2(n9016), .ZN(P3_U3456) );
  NOR2_X1 U11537 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n9020) );
  NAND2_X1 U11538 ( .A1(n9155), .A2(n9023), .ZN(n9024) );
  NOR2_X1 U11539 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n9026) );
  NOR2_X1 U11540 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n9025) );
  NAND2_X1 U11541 ( .A1(n9029), .A2(n6456), .ZN(n9030) );
  MUX2_X1 U11542 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9030), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n9031) );
  NAND2_X1 U11543 ( .A1(n9032), .A2(n6456), .ZN(n9033) );
  XNOR2_X1 U11544 ( .A(n9033), .B(P2_IR_REG_25__SCAN_IN), .ZN(n9274) );
  NAND3_X1 U11545 ( .A1(n13207), .A2(n11118), .A3(n9274), .ZN(n9296) );
  INV_X1 U11546 ( .A(n9034), .ZN(n9035) );
  NAND2_X1 U11547 ( .A1(n9035), .A2(n6456), .ZN(n9037) );
  INV_X1 U11548 ( .A(n10910), .ZN(n9038) );
  INV_X1 U11549 ( .A(n9039), .ZN(n12249) );
  NAND2_X1 U11550 ( .A1(n9041), .A2(n10112), .ZN(n9042) );
  MUX2_X1 U11551 ( .A(n9044), .B(n12077), .S(n11268), .Z(n9050) );
  NAND3_X1 U11552 ( .A1(n9045), .A2(n9067), .A3(n14781), .ZN(n9046) );
  NAND2_X1 U11553 ( .A1(n14776), .A2(n9067), .ZN(n9047) );
  NAND2_X1 U11554 ( .A1(n9048), .A2(n9047), .ZN(n9049) );
  XNOR2_X1 U11555 ( .A(n11268), .B(n10013), .ZN(n9051) );
  XNOR2_X1 U11556 ( .A(n9051), .B(n12279), .ZN(n10010) );
  NAND2_X1 U11557 ( .A1(n9051), .A2(n10463), .ZN(n9052) );
  XNOR2_X1 U11558 ( .A(n11268), .B(n9054), .ZN(n9057) );
  XNOR2_X1 U11559 ( .A(n9057), .B(n14761), .ZN(n10072) );
  INV_X1 U11560 ( .A(n9057), .ZN(n9058) );
  NAND2_X1 U11561 ( .A1(n9058), .A2(n10665), .ZN(n9059) );
  XNOR2_X1 U11562 ( .A(n9060), .B(n12278), .ZN(n10351) );
  XNOR2_X1 U11563 ( .A(n11268), .B(n10775), .ZN(n9061) );
  XNOR2_X1 U11564 ( .A(n9061), .B(n12277), .ZN(n10454) );
  NAND2_X1 U11565 ( .A1(n9061), .A2(n10728), .ZN(n9062) );
  XNOR2_X1 U11566 ( .A(n11268), .B(n9064), .ZN(n9065) );
  XNOR2_X1 U11567 ( .A(n9065), .B(n12276), .ZN(n10726) );
  NAND2_X1 U11568 ( .A1(n9065), .A2(n12276), .ZN(n9066) );
  XNOR2_X1 U11569 ( .A(n12226), .B(n9067), .ZN(n14670) );
  INV_X1 U11570 ( .A(n14670), .ZN(n9068) );
  NAND2_X1 U11571 ( .A1(n9068), .A2(n12107), .ZN(n9069) );
  XNOR2_X1 U11572 ( .A(n11268), .B(n9070), .ZN(n9072) );
  XNOR2_X1 U11573 ( .A(n9072), .B(n9071), .ZN(n10837) );
  NAND2_X1 U11574 ( .A1(n9072), .A2(n12275), .ZN(n9073) );
  XNOR2_X1 U11575 ( .A(n11268), .B(n12118), .ZN(n11067) );
  XNOR2_X1 U11576 ( .A(n11067), .B(n11072), .ZN(n9076) );
  INV_X1 U11577 ( .A(n9076), .ZN(n9074) );
  NAND2_X1 U11578 ( .A1(n9077), .A2(n9076), .ZN(n9080) );
  NAND2_X1 U11579 ( .A1(n9085), .A2(n14837), .ZN(n9078) );
  OAI22_X1 U11580 ( .A1(n9097), .A2(n9086), .B1(n9091), .B2(n9078), .ZN(n9079)
         );
  AOI21_X1 U11581 ( .B1(n11069), .B2(n9080), .A(n12023), .ZN(n9102) );
  NAND3_X1 U11582 ( .A1(n9083), .A2(n9082), .A3(n9081), .ZN(n9084) );
  AOI21_X1 U11583 ( .B1(n9091), .B2(n9085), .A(n9084), .ZN(n9089) );
  NAND2_X1 U11584 ( .A1(n9086), .A2(n12183), .ZN(n9087) );
  NAND2_X1 U11585 ( .A1(n9097), .A2(n9087), .ZN(n9088) );
  NAND2_X1 U11586 ( .A1(n9089), .A2(n9088), .ZN(n9944) );
  NOR2_X1 U11587 ( .A1(n14678), .A2(n10938), .ZN(n9101) );
  NAND2_X1 U11588 ( .A1(n12253), .A2(n14821), .ZN(n9090) );
  OR2_X1 U11589 ( .A1(n9091), .A2(n9090), .ZN(n9092) );
  AND2_X1 U11590 ( .A1(n14675), .A2(n12118), .ZN(n9100) );
  NAND2_X1 U11591 ( .A1(n12275), .A2(n14731), .ZN(n9094) );
  NAND2_X1 U11592 ( .A1(n12274), .A2(n14730), .ZN(n9093) );
  AND2_X1 U11593 ( .A1(n9094), .A2(n9093), .ZN(n10936) );
  NAND2_X1 U11594 ( .A1(n12253), .A2(n9095), .ZN(n9096) );
  OAI22_X1 U11595 ( .A1(n10936), .A2(n14666), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9098), .ZN(n9099) );
  INV_X2 U11596 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U11597 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n9103) );
  XOR2_X1 U11598 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9301), .Z(n9140) );
  INV_X1 U11599 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14649) );
  NOR3_X1 U11600 ( .A1(n9140), .A2(n14649), .A3(n9337), .ZN(n9139) );
  NOR2_X1 U11601 ( .A1(n9104), .A2(n13197), .ZN(n9105) );
  MUX2_X1 U11602 ( .A(n13197), .B(n9105), .S(P2_IR_REG_2__SCAN_IN), .Z(n9106)
         );
  INV_X1 U11603 ( .A(n9106), .ZN(n9108) );
  INV_X1 U11604 ( .A(n9162), .ZN(n9107) );
  NAND2_X1 U11605 ( .A1(n9108), .A2(n9107), .ZN(n9352) );
  XOR2_X1 U11606 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n9352), .Z(n9127) );
  NOR2_X1 U11607 ( .A1(n9128), .A2(n9127), .ZN(n9397) );
  NOR2_X2 U11608 ( .A1(n9109), .A2(n9110), .ZN(n9330) );
  NAND2_X1 U11609 ( .A1(n9326), .A2(n10910), .ZN(n9123) );
  NOR2_X1 U11610 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), 
        .ZN(n9116) );
  NOR2_X1 U11611 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n9115) );
  NOR2_X1 U11612 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), 
        .ZN(n9114) );
  NOR2_X1 U11613 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), 
        .ZN(n9113) );
  NAND2_X1 U11614 ( .A1(n13197), .A2(n9117), .ZN(n9119) );
  XNOR2_X2 U11615 ( .A(n9122), .B(n9121), .ZN(n13206) );
  NAND2_X1 U11616 ( .A1(n9123), .A2(n11026), .ZN(n9124) );
  NAND2_X1 U11617 ( .A1(n9125), .A2(n9124), .ZN(n9134) );
  NOR2_X1 U11618 ( .A1(n9323), .A2(P2_U3088), .ZN(n13202) );
  AOI211_X1 U11619 ( .C1(n9128), .C2(n9127), .A(n9397), .B(n14531), .ZN(n9138)
         );
  XNOR2_X1 U11620 ( .A(n9129), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n9143) );
  INV_X1 U11621 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14556) );
  NOR3_X1 U11622 ( .A1(n9143), .A2(n14556), .A3(n9337), .ZN(n9142) );
  AOI21_X1 U11623 ( .B1(n9129), .B2(P2_REG2_REG_1__SCAN_IN), .A(n9142), .ZN(
        n9132) );
  INV_X1 U11624 ( .A(n9352), .ZN(n9401) );
  XNOR2_X1 U11625 ( .A(n9401), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n9131) );
  NOR2_X1 U11626 ( .A1(n9132), .A2(n9131), .ZN(n9400) );
  INV_X1 U11627 ( .A(n13206), .ZN(n12822) );
  AOI211_X1 U11628 ( .C1(n9132), .C2(n9131), .A(n9400), .B(n14527), .ZN(n9137)
         );
  NOR2_X1 U11629 ( .A1(n14540), .A2(n14965), .ZN(n9136) );
  AND2_X1 U11630 ( .A1(n9323), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9133) );
  NAND2_X1 U11631 ( .A1(n9134), .A2(n9133), .ZN(n12815) );
  INV_X1 U11632 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10172) );
  OAI22_X1 U11633 ( .A1(n12815), .A2(n9352), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10172), .ZN(n9135) );
  OR4_X1 U11634 ( .A1(n9138), .A2(n9137), .A3(n9136), .A4(n9135), .ZN(P2_U3216) );
  NAND2_X1 U11635 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n9141) );
  AOI211_X1 U11636 ( .C1(n9141), .C2(n9140), .A(n9139), .B(n14531), .ZN(n9148)
         );
  NAND2_X1 U11637 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n9144) );
  AOI211_X1 U11638 ( .C1(n9144), .C2(n9143), .A(n9142), .B(n14527), .ZN(n9147)
         );
  NOR2_X1 U11639 ( .A1(n14540), .A2(n6985), .ZN(n9146) );
  INV_X1 U11640 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n10156) );
  OAI22_X1 U11641 ( .A1(n12815), .A2(n9301), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10156), .ZN(n9145) );
  OR4_X1 U11642 ( .A1(n9148), .A2(n9147), .A3(n9146), .A4(n9145), .ZN(P2_U3215) );
  AND2_X1 U11643 ( .A1(n9299), .A2(P1_U3086), .ZN(n10912) );
  INV_X2 U11644 ( .A(n10912), .ZN(n13837) );
  INV_X1 U11645 ( .A(n13376), .ZN(n9149) );
  OAI222_X1 U11646 ( .A1(n13833), .A2(n6987), .B1(n13837), .B2(n9348), .C1(
        P1_U3086), .C2(n9149), .ZN(P1_U3353) );
  INV_X1 U11647 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9151) );
  INV_X1 U11648 ( .A(n9512), .ZN(n9165) );
  INV_X1 U11649 ( .A(n13388), .ZN(n9150) );
  OAI222_X1 U11650 ( .A1(n13833), .A2(n9151), .B1(n13837), .B2(n9165), .C1(
        P1_U3086), .C2(n9150), .ZN(P1_U3352) );
  INV_X1 U11651 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9153) );
  INV_X1 U11652 ( .A(n9622), .ZN(n9158) );
  INV_X1 U11653 ( .A(n13400), .ZN(n9152) );
  OAI222_X1 U11654 ( .A1(n13833), .A2(n9153), .B1(n13837), .B2(n9158), .C1(
        P1_U3086), .C2(n9152), .ZN(P1_U3351) );
  INV_X2 U11655 ( .A(n10909), .ZN(n13213) );
  OR2_X1 U11656 ( .A1(n9830), .A2(n13197), .ZN(n9156) );
  XNOR2_X1 U11657 ( .A(n9156), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9623) );
  AOI22_X1 U11658 ( .A1(n9623), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n6626), .ZN(n9157) );
  OAI21_X1 U11659 ( .B1(n9158), .B2(n13213), .A(n9157), .ZN(P2_U3323) );
  INV_X1 U11660 ( .A(n9795), .ZN(n9169) );
  NAND2_X1 U11661 ( .A1(n9830), .A2(n9159), .ZN(n9181) );
  NAND2_X1 U11662 ( .A1(n9181), .A2(n6456), .ZN(n9160) );
  XNOR2_X1 U11663 ( .A(n9160), .B(P2_IR_REG_5__SCAN_IN), .ZN(n14463) );
  AOI22_X1 U11664 ( .A1(n14463), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n6626), .ZN(n9161) );
  OAI21_X1 U11665 ( .B1(n9169), .B2(n13213), .A(n9161), .ZN(P2_U3322) );
  OR2_X1 U11666 ( .A1(n9162), .A2(n13197), .ZN(n9163) );
  XNOR2_X1 U11667 ( .A(n9163), .B(P2_IR_REG_3__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U11668 ( .A1(n14451), .A2(P2_STATE_REG_SCAN_IN), .B1(n6626), .B2(
        P1_DATAO_REG_3__SCAN_IN), .ZN(n9164) );
  OAI21_X1 U11669 ( .B1(n9165), .B2(n13213), .A(n9164), .ZN(P2_U3324) );
  INV_X2 U11670 ( .A(n6626), .ZN(n13210) );
  OAI222_X1 U11671 ( .A1(P2_U3088), .A2(n9301), .B1(n13213), .B2(n9302), .C1(
        n9300), .C2(n13210), .ZN(P2_U3326) );
  OAI222_X1 U11672 ( .A1(n9352), .A2(P2_U3088), .B1(n13213), .B2(n9348), .C1(
        n9349), .C2(n13210), .ZN(P2_U3325) );
  NAND2_X1 U11673 ( .A1(n9299), .A2(P3_U3151), .ZN(n12657) );
  INV_X2 U11674 ( .A(n13947), .ZN(n12661) );
  INV_X1 U11675 ( .A(SI_7_), .ZN(n9166) );
  OAI222_X1 U11676 ( .A1(n12657), .A2(n9167), .B1(n12661), .B2(n9166), .C1(
        n9964), .C2(P3_U3151), .ZN(P3_U3288) );
  INV_X1 U11677 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9170) );
  INV_X1 U11678 ( .A(n9449), .ZN(n9168) );
  OAI222_X1 U11679 ( .A1(n13833), .A2(n9170), .B1(n13837), .B2(n9169), .C1(
        P1_U3086), .C2(n9168), .ZN(P1_U3350) );
  INV_X1 U11680 ( .A(n9171), .ZN(n9172) );
  OAI222_X1 U11681 ( .A1(P3_U3151), .A2(n9752), .B1(n12661), .B2(n9173), .C1(
        n12657), .C2(n9172), .ZN(P3_U3294) );
  OAI222_X1 U11682 ( .A1(n13833), .A2(n7837), .B1(n7985), .B2(P1_U3086), .C1(
        n13837), .C2(n9302), .ZN(P1_U3354) );
  OAI222_X1 U11683 ( .A1(n12657), .A2(n9176), .B1(n12661), .B2(n9175), .C1(
        n9174), .C2(P3_U3151), .ZN(P3_U3284) );
  INV_X1 U11684 ( .A(n13833), .ZN(n13819) );
  AOI22_X1 U11685 ( .A1(n13425), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n13819), .ZN(n9177) );
  OAI21_X1 U11686 ( .B1(n9977), .B2(n13837), .A(n9177), .ZN(P1_U3348) );
  INV_X1 U11687 ( .A(SI_9_), .ZN(n9179) );
  OAI222_X1 U11688 ( .A1(n12657), .A2(n9180), .B1(n12661), .B2(n9179), .C1(
        n9178), .C2(P3_U3151), .ZN(P3_U3286) );
  NAND2_X1 U11689 ( .A1(n9827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9182) );
  XNOR2_X1 U11690 ( .A(n9182), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9860) );
  INV_X1 U11691 ( .A(n9860), .ZN(n9496) );
  INV_X1 U11692 ( .A(n9859), .ZN(n9185) );
  OAI222_X1 U11693 ( .A1(n9496), .A2(P2_U3088), .B1(n13213), .B2(n9185), .C1(
        n9183), .C2(n13210), .ZN(P2_U3321) );
  INV_X1 U11694 ( .A(n13413), .ZN(n9184) );
  OAI222_X1 U11695 ( .A1(n13833), .A2(n9186), .B1(n13837), .B2(n9185), .C1(
        P1_U3086), .C2(n9184), .ZN(P1_U3349) );
  INV_X1 U11696 ( .A(n9193), .ZN(n9187) );
  NAND2_X1 U11697 ( .A1(n9187), .A2(n6456), .ZN(n9188) );
  XNOR2_X1 U11698 ( .A(n9188), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10002) );
  INV_X1 U11699 ( .A(n10002), .ZN(n9190) );
  INV_X1 U11700 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9189) );
  OAI222_X1 U11701 ( .A1(P2_U3088), .A2(n9190), .B1(n13213), .B2(n9977), .C1(
        n9189), .C2(n13210), .ZN(P2_U3320) );
  INV_X1 U11702 ( .A(n9467), .ZN(n9456) );
  OAI222_X1 U11703 ( .A1(n13837), .A2(n10085), .B1(n9456), .B2(P1_U3086), .C1(
        n9191), .C2(n13833), .ZN(P1_U3347) );
  NAND2_X1 U11704 ( .A1(n9193), .A2(n9192), .ZN(n9220) );
  NAND2_X1 U11705 ( .A1(n9220), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9194) );
  XNOR2_X1 U11706 ( .A(n9194), .B(P2_IR_REG_8__SCAN_IN), .ZN(n14474) );
  INV_X1 U11707 ( .A(n14474), .ZN(n9196) );
  INV_X1 U11708 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9195) );
  OAI222_X1 U11709 ( .A1(P2_U3088), .A2(n9196), .B1(n13213), .B2(n10085), .C1(
        n9195), .C2(n13210), .ZN(P2_U3319) );
  INV_X1 U11710 ( .A(n9197), .ZN(n9199) );
  OAI222_X1 U11711 ( .A1(n12664), .A2(n9199), .B1(n10633), .B2(P3_U3151), .C1(
        n9198), .C2(n12661), .ZN(P3_U3283) );
  INV_X1 U11712 ( .A(n9200), .ZN(n9202) );
  OAI222_X1 U11713 ( .A1(n12664), .A2(n9202), .B1(n12661), .B2(n9201), .C1(
        n10034), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U11714 ( .A1(n12664), .A2(n9204), .B1(n12661), .B2(n9203), .C1(
        n14718), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U11715 ( .A(SI_3_), .ZN(n9205) );
  OAI222_X1 U11716 ( .A1(n9207), .A2(P3_U3151), .B1(n12664), .B2(n9206), .C1(
        n9205), .C2(n12661), .ZN(P3_U3292) );
  INV_X1 U11717 ( .A(SI_4_), .ZN(n9208) );
  OAI222_X1 U11718 ( .A1(n9210), .A2(P3_U3151), .B1(n12664), .B2(n9209), .C1(
        n9208), .C2(n12661), .ZN(P3_U3291) );
  INV_X1 U11719 ( .A(SI_5_), .ZN(n9211) );
  OAI222_X1 U11720 ( .A1(n9788), .A2(P3_U3151), .B1(n12664), .B2(n9212), .C1(
        n9211), .C2(n12661), .ZN(P3_U3290) );
  INV_X1 U11721 ( .A(n9213), .ZN(n9215) );
  OAI222_X1 U11722 ( .A1(n9931), .A2(P3_U3151), .B1(n12664), .B2(n9215), .C1(
        n9214), .C2(n12661), .ZN(P3_U3289) );
  INV_X1 U11723 ( .A(n9216), .ZN(n9734) );
  INV_X1 U11724 ( .A(SI_2_), .ZN(n9217) );
  OAI222_X1 U11725 ( .A1(n9734), .A2(P3_U3151), .B1(n12664), .B2(n9218), .C1(
        n9217), .C2(n12661), .ZN(P3_U3293) );
  INV_X1 U11726 ( .A(n9471), .ZN(n9538) );
  OAI222_X1 U11727 ( .A1(n13837), .A2(n10177), .B1(n9538), .B2(P1_U3086), .C1(
        n9219), .C2(n13833), .ZN(P1_U3346) );
  NAND2_X1 U11728 ( .A1(n9228), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9221) );
  XNOR2_X1 U11729 ( .A(n9221), .B(P2_IR_REG_9__SCAN_IN), .ZN(n10528) );
  INV_X1 U11730 ( .A(n10528), .ZN(n9997) );
  INV_X1 U11731 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9222) );
  OAI222_X1 U11732 ( .A1(P2_U3088), .A2(n9997), .B1(n13213), .B2(n10177), .C1(
        n9222), .C2(n13210), .ZN(P2_U3318) );
  OAI222_X1 U11733 ( .A1(n12657), .A2(n9224), .B1(n12661), .B2(n9223), .C1(
        n10922), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U11734 ( .A(n10268), .ZN(n9231) );
  AOI22_X1 U11735 ( .A1(n13440), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n13819), .ZN(n9225) );
  OAI21_X1 U11736 ( .B1(n9231), .B2(n13837), .A(n9225), .ZN(P1_U3345) );
  INV_X1 U11737 ( .A(SI_14_), .ZN(n9226) );
  OAI222_X1 U11738 ( .A1(n12657), .A2(n9227), .B1(n12661), .B2(n9226), .C1(
        n11084), .C2(P3_U3151), .ZN(P3_U3281) );
  NAND2_X1 U11739 ( .A1(n9264), .A2(n6456), .ZN(n9229) );
  XNOR2_X1 U11740 ( .A(n9229), .B(P2_IR_REG_10__SCAN_IN), .ZN(n14486) );
  INV_X1 U11741 ( .A(n14486), .ZN(n9232) );
  INV_X1 U11742 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9230) );
  OAI222_X1 U11743 ( .A1(n9232), .A2(P2_U3088), .B1(n13213), .B2(n9231), .C1(
        n9230), .C2(n13210), .ZN(P2_U3317) );
  NAND2_X1 U11744 ( .A1(n9233), .A2(P1_B_REG_SCAN_IN), .ZN(n9235) );
  MUX2_X1 U11745 ( .A(n9235), .B(P1_B_REG_SCAN_IN), .S(n9234), .Z(n9236) );
  NAND2_X1 U11746 ( .A1(n9243), .A2(n13835), .ZN(n9238) );
  OAI22_X1 U11747 ( .A1(n14350), .A2(P1_D_REG_0__SCAN_IN), .B1(n9234), .B2(
        n9238), .ZN(n9237) );
  INV_X1 U11748 ( .A(n9237), .ZN(P1_U3445) );
  OAI22_X1 U11749 ( .A1(n14350), .A2(P1_D_REG_1__SCAN_IN), .B1(n9239), .B2(
        n9238), .ZN(n9240) );
  INV_X1 U11750 ( .A(n9240), .ZN(P1_U3446) );
  INV_X1 U11751 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U11752 ( .A1(n9241), .A2(n12636), .ZN(n9242) );
  OAI21_X1 U11753 ( .B1(n12636), .B2(n14896), .A(n9242), .ZN(P3_U3376) );
  INV_X1 U11754 ( .A(n9243), .ZN(n9244) );
  INV_X1 U11755 ( .A(n15020), .ZN(P1_U4016) );
  NAND2_X1 U11756 ( .A1(n9246), .A2(n9245), .ZN(n9248) );
  NAND2_X1 U11757 ( .A1(n9248), .A2(n9247), .ZN(n9250) );
  INV_X1 U11758 ( .A(n14288), .ZN(n9607) );
  NOR2_X1 U11759 ( .A1(n9607), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11760 ( .A(n10420), .ZN(n9268) );
  AOI22_X1 U11761 ( .A1(n9601), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n13819), .ZN(n9249) );
  OAI21_X1 U11762 ( .B1(n9268), .B2(n13837), .A(n9249), .ZN(P1_U3344) );
  AND2_X1 U11763 ( .A1(n9262), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11764 ( .A1(n9262), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U11765 ( .A1(n9262), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11766 ( .A1(n9262), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11767 ( .A1(n9262), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11768 ( .A1(n9262), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11769 ( .A1(n9262), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11770 ( .A1(n9262), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11771 ( .A1(n9262), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11772 ( .A1(n9262), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11773 ( .A1(n9262), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11774 ( .A1(n9262), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11775 ( .A1(n9262), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11776 ( .A1(n9262), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11777 ( .A1(n9262), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U11778 ( .A1(n9262), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11779 ( .A1(n9262), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11780 ( .A1(n9262), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11781 ( .A1(n9262), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11782 ( .A1(n9262), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11783 ( .A1(n9262), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11784 ( .A1(n9262), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U11785 ( .A1(n9262), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11786 ( .A1(n9262), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U11787 ( .A1(n9262), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11788 ( .A1(n9262), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11789 ( .A1(n9262), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11790 ( .A1(n9262), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  INV_X1 U11791 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9257) );
  INV_X1 U11792 ( .A(n9250), .ZN(n9251) );
  NAND2_X1 U11793 ( .A1(n9252), .A2(n9251), .ZN(n9437) );
  INV_X1 U11794 ( .A(n9437), .ZN(n9423) );
  INV_X1 U11795 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9253) );
  OAI21_X1 U11796 ( .B1(n8530), .B2(P1_REG2_REG_0__SCAN_IN), .A(n9543), .ZN(
        n13371) );
  AOI21_X1 U11797 ( .B1(n8530), .B2(n9253), .A(n13371), .ZN(n9254) );
  XNOR2_X1 U11798 ( .A(n9254), .B(n7373), .ZN(n9255) );
  AOI22_X1 U11799 ( .A1(n9423), .A2(n9255), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n9256) );
  OAI21_X1 U11800 ( .B1(n14288), .B2(n9257), .A(n9256), .ZN(P1_U3243) );
  INV_X1 U11801 ( .A(n9258), .ZN(n9261) );
  OAI222_X1 U11802 ( .A1(n12664), .A2(n9261), .B1(n12661), .B2(n9260), .C1(
        n9259), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U11803 ( .A(n9262), .ZN(n9263) );
  INV_X1 U11804 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n14898) );
  NOR2_X1 U11805 ( .A1(n9263), .A2(n14898), .ZN(P3_U3243) );
  INV_X1 U11806 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n14928) );
  NOR2_X1 U11807 ( .A1(n9263), .A2(n14928), .ZN(P3_U3242) );
  INV_X1 U11808 ( .A(n9391), .ZN(n9265) );
  NAND2_X1 U11809 ( .A1(n9265), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9266) );
  XNOR2_X1 U11810 ( .A(n9266), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10706) );
  INV_X1 U11811 ( .A(n10706), .ZN(n10526) );
  OAI222_X1 U11812 ( .A1(P2_U3088), .A2(n10526), .B1(n13213), .B2(n9268), .C1(
        n9267), .C2(n13210), .ZN(P2_U3316) );
  INV_X1 U11813 ( .A(P2_B_REG_SCAN_IN), .ZN(n9269) );
  XNOR2_X1 U11814 ( .A(n11118), .B(n9269), .ZN(n9270) );
  INV_X1 U11815 ( .A(n9274), .ZN(n13214) );
  NAND2_X1 U11816 ( .A1(n9270), .A2(n13214), .ZN(n9271) );
  INV_X1 U11817 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U11818 ( .A1(n14558), .A2(n14561), .ZN(n9273) );
  OR2_X1 U11819 ( .A1(n11118), .A2(n13207), .ZN(n9272) );
  NAND2_X1 U11820 ( .A1(n9273), .A2(n9272), .ZN(n14562) );
  INV_X1 U11821 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14564) );
  NAND2_X1 U11822 ( .A1(n14558), .A2(n14564), .ZN(n9276) );
  OR2_X1 U11823 ( .A1(n13207), .A2(n9274), .ZN(n9275) );
  NAND2_X1 U11824 ( .A1(n9276), .A2(n9275), .ZN(n14565) );
  INV_X1 U11825 ( .A(n14565), .ZN(n10052) );
  NOR4_X1 U11826 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_8__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n9285) );
  OR4_X1 U11827 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_11__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n9282) );
  NOR4_X1 U11828 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9280) );
  NOR4_X1 U11829 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9279) );
  NOR4_X1 U11830 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9278) );
  NOR4_X1 U11831 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9277) );
  NAND4_X1 U11832 ( .A1(n9280), .A2(n9279), .A3(n9278), .A4(n9277), .ZN(n9281)
         );
  NOR4_X1 U11833 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9282), .A4(n9281), .ZN(n9284) );
  NOR4_X1 U11834 ( .A1(P2_D_REG_3__SCAN_IN), .A2(P2_D_REG_4__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9283) );
  NAND3_X1 U11835 ( .A1(n9285), .A2(n9284), .A3(n9283), .ZN(n9286) );
  NAND2_X1 U11836 ( .A1(n14558), .A2(n9286), .ZN(n9572) );
  NAND3_X1 U11837 ( .A1(n9585), .A2(n10052), .A3(n9572), .ZN(n9295) );
  NAND2_X1 U11838 ( .A1(n9287), .A2(n6456), .ZN(n9288) );
  INV_X1 U11839 ( .A(n9289), .ZN(n9290) );
  NAND2_X1 U11840 ( .A1(n9292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U11841 ( .A1(n14630), .A2(n11672), .ZN(n9573) );
  NAND2_X1 U11842 ( .A1(n9295), .A2(n9573), .ZN(n9298) );
  AND2_X1 U11843 ( .A1(n9296), .A2(n10910), .ZN(n9304) );
  NAND2_X1 U11844 ( .A1(n11671), .A2(n12819), .ZN(n11639) );
  NAND2_X1 U11845 ( .A1(n9326), .A2(n11639), .ZN(n9571) );
  AND2_X1 U11846 ( .A1(n9304), .A2(n9571), .ZN(n9297) );
  NAND2_X1 U11847 ( .A1(n9298), .A2(n9297), .ZN(n9515) );
  NOR2_X1 U11848 ( .A1(n9515), .A2(P2_U3088), .ZN(n9487) );
  OR2_X1 U11850 ( .A1(n10758), .A2(n9300), .ZN(n9303) );
  NAND4_X1 U11851 ( .A1(n9585), .A2(n10052), .A3(n14566), .A4(n9572), .ZN(
        n9329) );
  INV_X1 U11852 ( .A(n9329), .ZN(n9305) );
  NOR2_X1 U11853 ( .A1(n14543), .A2(n11671), .ZN(n10056) );
  NAND2_X1 U11854 ( .A1(n9305), .A2(n10056), .ZN(n9307) );
  INV_X1 U11855 ( .A(n9573), .ZN(n9306) );
  NAND2_X1 U11856 ( .A1(n9308), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9310) );
  NAND2_X1 U11857 ( .A1(n9354), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11858 ( .A1(n9353), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n9314) );
  INV_X1 U11859 ( .A(n11289), .ZN(n9481) );
  INV_X1 U11860 ( .A(n9323), .ZN(n9318) );
  NAND2_X1 U11861 ( .A1(n11289), .A2(n12754), .ZN(n9325) );
  NAND2_X1 U11862 ( .A1(n9354), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9322) );
  NAND2_X1 U11863 ( .A1(n9353), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n9319) );
  AND2_X2 U11864 ( .A1(n9326), .A2(n9323), .ZN(n12824) );
  NAND2_X1 U11865 ( .A1(n12782), .A2(n12824), .ZN(n9324) );
  NAND2_X1 U11866 ( .A1(n9325), .A2(n9324), .ZN(n9579) );
  AOI22_X1 U11867 ( .A1(n11294), .A2(n12747), .B1(n12757), .B2(n9579), .ZN(
        n9346) );
  INV_X1 U11868 ( .A(n11639), .ZN(n11685) );
  INV_X1 U11869 ( .A(n9326), .ZN(n9327) );
  NAND2_X1 U11870 ( .A1(n14627), .A2(n9327), .ZN(n9328) );
  INV_X1 U11871 ( .A(n9294), .ZN(n9331) );
  NAND2_X1 U11872 ( .A1(n9354), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11873 ( .A1(n9517), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9335) );
  NAND2_X1 U11874 ( .A1(n9353), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n9334) );
  NAND2_X1 U11875 ( .A1(n9355), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U11876 ( .A1(n11293), .A2(n9339), .ZN(n9370) );
  NAND2_X1 U11877 ( .A1(n9481), .A2(n14545), .ZN(n9577) );
  NAND2_X1 U11878 ( .A1(n11713), .A2(n14545), .ZN(n9340) );
  NAND2_X1 U11879 ( .A1(n9577), .A2(n9340), .ZN(n9482) );
  AND2_X1 U11880 ( .A1(n6459), .A2(n11284), .ZN(n9341) );
  OR2_X1 U11881 ( .A1(n9482), .A2(n9341), .ZN(n9342) );
  OAI21_X1 U11882 ( .B1(n9343), .B2(n9342), .A(n9373), .ZN(n9344) );
  NAND2_X1 U11883 ( .A1(n12763), .A2(n9344), .ZN(n9345) );
  OAI211_X1 U11884 ( .C1(n9487), .C2(n10156), .A(n9346), .B(n9345), .ZN(
        P2_U3194) );
  INV_X1 U11885 ( .A(n9347), .ZN(n9348) );
  INV_X1 U11886 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10063) );
  NAND2_X1 U11887 ( .A1(n11590), .A2(n10063), .ZN(n9359) );
  NAND2_X1 U11888 ( .A1(n9354), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9358) );
  NAND2_X1 U11889 ( .A1(n9517), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9357) );
  NAND2_X1 U11890 ( .A1(n9355), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11891 ( .A1(n12781), .A2(n12824), .ZN(n9361) );
  NAND2_X1 U11892 ( .A1(n11293), .A2(n12754), .ZN(n9360) );
  AND2_X1 U11893 ( .A1(n9361), .A2(n9360), .ZN(n10170) );
  INV_X1 U11894 ( .A(n10170), .ZN(n9362) );
  AOI22_X1 U11895 ( .A1(n9363), .A2(n12747), .B1(n12757), .B2(n9362), .ZN(
        n9378) );
  XNOR2_X1 U11896 ( .A(n9510), .B(n10046), .ZN(n9364) );
  NAND2_X1 U11897 ( .A1(n12782), .A2(n9339), .ZN(n9365) );
  NAND2_X1 U11898 ( .A1(n9364), .A2(n9365), .ZN(n9508) );
  INV_X1 U11899 ( .A(n9364), .ZN(n9367) );
  INV_X1 U11900 ( .A(n9365), .ZN(n9366) );
  NAND2_X1 U11901 ( .A1(n9367), .A2(n9366), .ZN(n9368) );
  AND2_X1 U11902 ( .A1(n9508), .A2(n9368), .ZN(n9375) );
  INV_X1 U11903 ( .A(n9369), .ZN(n9371) );
  NAND2_X1 U11904 ( .A1(n9371), .A2(n9370), .ZN(n9372) );
  NAND2_X1 U11905 ( .A1(n9373), .A2(n9372), .ZN(n9374) );
  NAND2_X1 U11906 ( .A1(n9374), .A2(n9375), .ZN(n9509) );
  OAI21_X1 U11907 ( .B1(n9375), .B2(n9374), .A(n9509), .ZN(n9376) );
  NAND2_X1 U11908 ( .A1(n9376), .A2(n12763), .ZN(n9377) );
  OAI211_X1 U11909 ( .C1(n9487), .C2(n10172), .A(n9378), .B(n9377), .ZN(
        P2_U3209) );
  INV_X1 U11910 ( .A(n10590), .ZN(n9396) );
  AOI22_X1 U11911 ( .A1(n13451), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n13819), .ZN(n9379) );
  OAI21_X1 U11912 ( .B1(n9396), .B2(n13837), .A(n9379), .ZN(P1_U3343) );
  INV_X1 U11913 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14957) );
  INV_X1 U11914 ( .A(n14527), .ZN(n9999) );
  AOI22_X1 U11915 ( .A1(n9999), .A2(P2_REG2_REG_0__SCAN_IN), .B1(n12814), .B2(
        P2_REG1_REG_0__SCAN_IN), .ZN(n9382) );
  NOR2_X1 U11916 ( .A1(n14527), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9380) );
  AOI211_X1 U11917 ( .C1(n12814), .C2(n14649), .A(n14537), .B(n9380), .ZN(
        n9381) );
  MUX2_X1 U11918 ( .A(n9382), .B(n9381), .S(P2_IR_REG_0__SCAN_IN), .Z(n9384)
         );
  NAND2_X1 U11919 ( .A1(n14442), .A2(P2_ADDR_REG_0__SCAN_IN), .ZN(n9383) );
  OAI211_X1 U11920 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n14957), .A(n9384), .B(
        n9383), .ZN(P2_U3214) );
  NAND2_X1 U11921 ( .A1(n13256), .A2(P1_U4016), .ZN(n9385) );
  OAI21_X1 U11922 ( .B1(n11449), .B2(P1_U4016), .A(n9385), .ZN(P1_U3580) );
  INV_X1 U11923 ( .A(n9386), .ZN(n9389) );
  OAI222_X1 U11924 ( .A1(n12657), .A2(n9389), .B1(n9388), .B2(P3_U3151), .C1(
        n9387), .C2(n12661), .ZN(P3_U3279) );
  INV_X1 U11925 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11926 ( .A1(n9391), .A2(n9390), .ZN(n9393) );
  NAND2_X1 U11927 ( .A1(n9393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9392) );
  MUX2_X1 U11928 ( .A(n6456), .B(n9392), .S(P2_IR_REG_12__SCAN_IN), .Z(n9394)
         );
  INV_X1 U11929 ( .A(n10882), .ZN(n10711) );
  OAI222_X1 U11930 ( .A1(P2_U3088), .A2(n10711), .B1(n13213), .B2(n9396), .C1(
        n9395), .C2(n13210), .ZN(P2_U3315) );
  XNOR2_X1 U11931 ( .A(n14451), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n14447) );
  XNOR2_X1 U11932 ( .A(n9623), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n9398) );
  AOI211_X1 U11933 ( .C1(n9399), .C2(n9398), .A(n14531), .B(n9488), .ZN(n9407)
         );
  XNOR2_X1 U11934 ( .A(n14451), .B(P2_REG2_REG_3__SCAN_IN), .ZN(n14444) );
  XNOR2_X1 U11935 ( .A(n9623), .B(P2_REG2_REG_4__SCAN_IN), .ZN(n9402) );
  AOI211_X1 U11936 ( .C1(n9403), .C2(n9402), .A(n14527), .B(n9492), .ZN(n9406)
         );
  INV_X1 U11937 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n13883) );
  NAND2_X1 U11938 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n9641) );
  NAND2_X1 U11939 ( .A1(n14537), .A2(n9623), .ZN(n9404) );
  OAI211_X1 U11940 ( .C1(n14540), .C2(n13883), .A(n9641), .B(n9404), .ZN(n9405) );
  OR3_X1 U11941 ( .A1(n9407), .A2(n9406), .A3(n9405), .ZN(P2_U3218) );
  NAND2_X1 U11942 ( .A1(n12280), .A2(P3_DATAO_REG_15__SCAN_IN), .ZN(n9408) );
  OAI21_X1 U11943 ( .B1(n12468), .B2(n12280), .A(n9408), .ZN(P3_U3506) );
  INV_X1 U11944 ( .A(n10757), .ZN(n9506) );
  AOI22_X1 U11945 ( .A1(n14190), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n13819), .ZN(n9409) );
  OAI21_X1 U11946 ( .B1(n9506), .B2(n13837), .A(n9409), .ZN(P1_U3342) );
  INV_X1 U11947 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n14435) );
  MUX2_X1 U11948 ( .A(n14435), .B(P1_REG1_REG_8__SCAN_IN), .S(n9467), .Z(n9422) );
  INV_X1 U11949 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n14427) );
  MUX2_X1 U11950 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n14427), .S(n13376), .Z(
        n13382) );
  INV_X1 U11951 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9410) );
  XNOR2_X1 U11952 ( .A(n13359), .B(n9410), .ZN(n13362) );
  AND2_X1 U11953 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13361) );
  NAND2_X1 U11954 ( .A1(n13362), .A2(n13361), .ZN(n13360) );
  NAND2_X1 U11955 ( .A1(n13359), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11956 ( .A1(n13360), .A2(n9411), .ZN(n13381) );
  NAND2_X1 U11957 ( .A1(n13382), .A2(n13381), .ZN(n13380) );
  NAND2_X1 U11958 ( .A1(n13376), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U11959 ( .A1(n13380), .A2(n9412), .ZN(n13390) );
  INV_X1 U11960 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9823) );
  MUX2_X1 U11961 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9823), .S(n13388), .Z(
        n13391) );
  NAND2_X1 U11962 ( .A1(n13390), .A2(n13391), .ZN(n13389) );
  NAND2_X1 U11963 ( .A1(n13388), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9413) );
  NAND2_X1 U11964 ( .A1(n13389), .A2(n9413), .ZN(n13402) );
  INV_X1 U11965 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14429) );
  MUX2_X1 U11966 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n14429), .S(n13400), .Z(
        n13403) );
  NAND2_X1 U11967 ( .A1(n13402), .A2(n13403), .ZN(n13401) );
  NAND2_X1 U11968 ( .A1(n13400), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n9414) );
  NAND2_X1 U11969 ( .A1(n13401), .A2(n9414), .ZN(n9445) );
  XNOR2_X1 U11970 ( .A(n9449), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9446) );
  OR2_X1 U11971 ( .A1(n9445), .A2(n9446), .ZN(n9443) );
  OR2_X1 U11972 ( .A1(n9449), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n9415) );
  AND2_X1 U11973 ( .A1(n9443), .A2(n9415), .ZN(n13415) );
  INV_X1 U11974 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9416) );
  XNOR2_X1 U11975 ( .A(n13413), .B(n9416), .ZN(n13416) );
  NAND2_X1 U11976 ( .A1(n13415), .A2(n13416), .ZN(n13414) );
  NAND2_X1 U11977 ( .A1(n13413), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9417) );
  NAND2_X1 U11978 ( .A1(n13414), .A2(n9417), .ZN(n13427) );
  INV_X1 U11979 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9418) );
  XNOR2_X1 U11980 ( .A(n13425), .B(n9418), .ZN(n13428) );
  NAND2_X1 U11981 ( .A1(n13427), .A2(n13428), .ZN(n13426) );
  NAND2_X1 U11982 ( .A1(n13425), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n9419) );
  NAND2_X1 U11983 ( .A1(n13426), .A2(n9419), .ZN(n9421) );
  OR2_X1 U11984 ( .A1(n9421), .A2(n9422), .ZN(n9458) );
  INV_X1 U11985 ( .A(n9458), .ZN(n9420) );
  AOI21_X1 U11986 ( .B1(n9422), .B2(n9421), .A(n9420), .ZN(n9442) );
  NOR2_X2 U11987 ( .A1(n9437), .A2(n9543), .ZN(n14276) );
  INV_X1 U11988 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n13853) );
  NAND2_X1 U11989 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10855) );
  OAI21_X1 U11990 ( .B1(n14288), .B2(n13853), .A(n10855), .ZN(n9424) );
  AOI21_X1 U11991 ( .B1(n14276), .B2(n9467), .A(n9424), .ZN(n9441) );
  INV_X1 U11992 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10449) );
  XNOR2_X1 U11993 ( .A(n9467), .B(n10449), .ZN(n9439) );
  INV_X1 U11994 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10583) );
  MUX2_X1 U11995 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10583), .S(n13376), .Z(
        n13379) );
  INV_X1 U11996 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9425) );
  XNOR2_X1 U11997 ( .A(n13359), .B(n9425), .ZN(n13364) );
  AND2_X1 U11998 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13368) );
  NAND2_X1 U11999 ( .A1(n13364), .A2(n13368), .ZN(n13363) );
  NAND2_X1 U12000 ( .A1(n13359), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n9426) );
  NAND2_X1 U12001 ( .A1(n13363), .A2(n9426), .ZN(n13378) );
  NAND2_X1 U12002 ( .A1(n13379), .A2(n13378), .ZN(n13377) );
  NAND2_X1 U12003 ( .A1(n13376), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9427) );
  NAND2_X1 U12004 ( .A1(n13377), .A2(n9427), .ZN(n13393) );
  INV_X1 U12005 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n14314) );
  MUX2_X1 U12006 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n14314), .S(n13388), .Z(
        n13394) );
  NAND2_X1 U12007 ( .A1(n13393), .A2(n13394), .ZN(n13392) );
  NAND2_X1 U12008 ( .A1(n13388), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n9428) );
  NAND2_X1 U12009 ( .A1(n13392), .A2(n9428), .ZN(n13405) );
  INV_X1 U12010 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10659) );
  MUX2_X1 U12011 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n10659), .S(n13400), .Z(
        n13406) );
  NAND2_X1 U12012 ( .A1(n13405), .A2(n13406), .ZN(n13404) );
  NAND2_X1 U12013 ( .A1(n13400), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9429) );
  NAND2_X1 U12014 ( .A1(n13404), .A2(n9429), .ZN(n9451) );
  INV_X1 U12015 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9430) );
  XNOR2_X1 U12016 ( .A(n9449), .B(n9430), .ZN(n9452) );
  NAND2_X1 U12017 ( .A1(n9451), .A2(n9452), .ZN(n9450) );
  NAND2_X1 U12018 ( .A1(n9449), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n9431) );
  NAND2_X1 U12019 ( .A1(n9450), .A2(n9431), .ZN(n13418) );
  INV_X1 U12020 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n9432) );
  XNOR2_X1 U12021 ( .A(n13413), .B(n9432), .ZN(n13419) );
  NAND2_X1 U12022 ( .A1(n13418), .A2(n13419), .ZN(n13417) );
  NAND2_X1 U12023 ( .A1(n13413), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9433) );
  NAND2_X1 U12024 ( .A1(n13417), .A2(n9433), .ZN(n13430) );
  INV_X1 U12025 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9434) );
  XNOR2_X1 U12026 ( .A(n13425), .B(n9434), .ZN(n13431) );
  NAND2_X1 U12027 ( .A1(n13430), .A2(n13431), .ZN(n13429) );
  NAND2_X1 U12028 ( .A1(n13425), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9435) );
  NAND2_X1 U12029 ( .A1(n13429), .A2(n9435), .ZN(n9438) );
  NAND2_X1 U12030 ( .A1(n13492), .A2(n9543), .ZN(n9436) );
  NOR2_X2 U12031 ( .A1(n9437), .A2(n9436), .ZN(n14280) );
  NAND2_X1 U12032 ( .A1(n9438), .A2(n9439), .ZN(n9469) );
  OAI211_X1 U12033 ( .C1(n9439), .C2(n9438), .A(n14280), .B(n9469), .ZN(n9440)
         );
  OAI211_X1 U12034 ( .C1(n9442), .C2(n14284), .A(n9441), .B(n9440), .ZN(
        P1_U3251) );
  INV_X1 U12035 ( .A(n9443), .ZN(n9444) );
  AOI21_X1 U12036 ( .B1(n9446), .B2(n9445), .A(n9444), .ZN(n9455) );
  INV_X1 U12037 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U12038 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9447) );
  OAI21_X1 U12039 ( .B1(n14288), .B2(n13898), .A(n9447), .ZN(n9448) );
  AOI21_X1 U12040 ( .B1(n14276), .B2(n9449), .A(n9448), .ZN(n9454) );
  OAI211_X1 U12041 ( .C1(n9452), .C2(n9451), .A(n14280), .B(n9450), .ZN(n9453)
         );
  OAI211_X1 U12042 ( .C1(n9455), .C2(n14284), .A(n9454), .B(n9453), .ZN(
        P1_U3248) );
  INV_X1 U12043 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14155) );
  MUX2_X1 U12044 ( .A(n14155), .B(P1_REG1_REG_11__SCAN_IN), .S(n9601), .Z(
        n9464) );
  NAND2_X1 U12045 ( .A1(n9456), .A2(n14435), .ZN(n9457) );
  NAND2_X1 U12046 ( .A1(n9458), .A2(n9457), .ZN(n9530) );
  INV_X1 U12047 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9459) );
  MUX2_X1 U12048 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9459), .S(n9471), .Z(n9531)
         );
  NAND2_X1 U12049 ( .A1(n9530), .A2(n9531), .ZN(n9529) );
  NAND2_X1 U12050 ( .A1(n9538), .A2(n9459), .ZN(n9460) );
  AND2_X1 U12051 ( .A1(n9529), .A2(n9460), .ZN(n13437) );
  INV_X1 U12052 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14439) );
  MUX2_X1 U12053 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n14439), .S(n13440), .Z(
        n13436) );
  NAND2_X1 U12054 ( .A1(n13437), .A2(n13436), .ZN(n13435) );
  NAND2_X1 U12055 ( .A1(n13440), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9461) );
  NAND2_X1 U12056 ( .A1(n13435), .A2(n9461), .ZN(n9463) );
  OR2_X1 U12057 ( .A1(n9463), .A2(n9464), .ZN(n9603) );
  INV_X1 U12058 ( .A(n9603), .ZN(n9462) );
  AOI21_X1 U12059 ( .B1(n9464), .B2(n9463), .A(n9462), .ZN(n9480) );
  INV_X1 U12060 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9465) );
  NAND2_X1 U12061 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n11111)
         );
  OAI21_X1 U12062 ( .B1(n14288), .B2(n9465), .A(n11111), .ZN(n9466) );
  AOI21_X1 U12063 ( .B1(n14276), .B2(n9601), .A(n9466), .ZN(n9479) );
  NAND2_X1 U12064 ( .A1(n9467), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9468) );
  NAND2_X1 U12065 ( .A1(n9469), .A2(n9468), .ZN(n9534) );
  INV_X1 U12066 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9470) );
  MUX2_X1 U12067 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n9470), .S(n9471), .Z(n9535)
         );
  NAND2_X1 U12068 ( .A1(n9534), .A2(n9535), .ZN(n9533) );
  NAND2_X1 U12069 ( .A1(n9471), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9472) );
  NAND2_X1 U12070 ( .A1(n9533), .A2(n9472), .ZN(n13442) );
  INV_X1 U12071 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9473) );
  XNOR2_X1 U12072 ( .A(n13440), .B(n9473), .ZN(n13443) );
  NAND2_X1 U12073 ( .A1(n13442), .A2(n13443), .ZN(n13441) );
  NAND2_X1 U12074 ( .A1(n13440), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9474) );
  NAND2_X1 U12075 ( .A1(n13441), .A2(n9474), .ZN(n9477) );
  INV_X1 U12076 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9475) );
  XNOR2_X1 U12077 ( .A(n9601), .B(n9475), .ZN(n9476) );
  NAND2_X1 U12078 ( .A1(n9477), .A2(n9476), .ZN(n9596) );
  OAI211_X1 U12079 ( .C1(n9477), .C2(n9476), .A(n9596), .B(n14280), .ZN(n9478)
         );
  OAI211_X1 U12080 ( .C1(n9480), .C2(n14284), .A(n9479), .B(n9478), .ZN(
        P1_U3254) );
  NAND2_X1 U12081 ( .A1(n11293), .A2(n12824), .ZN(n14550) );
  NOR3_X1 U12082 ( .A1(n9481), .A2(n14545), .A3(n12952), .ZN(n9483) );
  OAI21_X1 U12083 ( .B1(n9483), .B2(n9482), .A(n12763), .ZN(n9484) );
  OAI21_X1 U12084 ( .B1(n14550), .B2(n12744), .A(n9484), .ZN(n9485) );
  AOI21_X1 U12085 ( .B1(n14545), .B2(n12747), .A(n9485), .ZN(n9486) );
  OAI21_X1 U12086 ( .B1(n9487), .B2(n14957), .A(n9486), .ZN(P2_U3204) );
  XNOR2_X1 U12087 ( .A(n14463), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n14459) );
  INV_X1 U12088 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9489) );
  MUX2_X1 U12089 ( .A(n9489), .B(P2_REG1_REG_6__SCAN_IN), .S(n9860), .Z(n9490)
         );
  NOR2_X1 U12090 ( .A1(n9491), .A2(n9490), .ZN(n9681) );
  AOI211_X1 U12091 ( .C1(n9491), .C2(n9490), .A(n14531), .B(n9681), .ZN(n9499)
         );
  XNOR2_X1 U12092 ( .A(n14463), .B(P2_REG2_REG_5__SCAN_IN), .ZN(n14456) );
  XNOR2_X1 U12093 ( .A(n9860), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n9493) );
  NOR2_X1 U12094 ( .A1(n9494), .A2(n9493), .ZN(n9685) );
  AOI211_X1 U12095 ( .C1(n9494), .C2(n9493), .A(n14527), .B(n9685), .ZN(n9498)
         );
  NAND2_X1 U12096 ( .A1(n14442), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9495) );
  NAND2_X1 U12097 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9873) );
  OAI211_X1 U12098 ( .C1(n12815), .C2(n9496), .A(n9495), .B(n9873), .ZN(n9497)
         );
  OR3_X1 U12099 ( .A1(n9499), .A2(n9498), .A3(n9497), .ZN(P2_U3220) );
  INV_X1 U12100 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n14901) );
  NAND2_X1 U12101 ( .A1(n12107), .A2(P3_U3897), .ZN(n9500) );
  OAI21_X1 U12102 ( .B1(P3_U3897), .B2(n14901), .A(n9500), .ZN(P3_U3498) );
  NAND2_X1 U12103 ( .A1(n9502), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U12104 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9501), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n9505) );
  INV_X1 U12105 ( .A(n9502), .ZN(n9504) );
  INV_X1 U12106 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U12107 ( .A1(n9504), .A2(n9503), .ZN(n9719) );
  NAND2_X1 U12108 ( .A1(n9505), .A2(n9719), .ZN(n10888) );
  OAI222_X1 U12109 ( .A1(P2_U3088), .A2(n10888), .B1(n13213), .B2(n9506), .C1(
        n10759), .C2(n13210), .ZN(P2_U3314) );
  INV_X1 U12110 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n15007) );
  NAND2_X1 U12111 ( .A1(n10665), .A2(P3_U3897), .ZN(n9507) );
  OAI21_X1 U12112 ( .B1(P3_U3897), .B2(n15007), .A(n9507), .ZN(P3_U3494) );
  NAND2_X1 U12113 ( .A1(n9509), .A2(n9508), .ZN(n9621) );
  AOI22_X1 U12114 ( .A1(n11434), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n11433), 
        .B2(n14451), .ZN(n9514) );
  NAND2_X1 U12115 ( .A1(n9512), .A2(n11584), .ZN(n9513) );
  INV_X1 U12116 ( .A(n14579), .ZN(n10118) );
  XNOR2_X1 U12117 ( .A(n9510), .B(n10118), .ZN(n9615) );
  NAND2_X1 U12118 ( .A1(n12781), .A2(n9339), .ZN(n9616) );
  XNOR2_X1 U12119 ( .A(n9615), .B(n9616), .ZN(n9620) );
  XNOR2_X1 U12120 ( .A(n9621), .B(n9620), .ZN(n9527) );
  NAND2_X1 U12121 ( .A1(n9354), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9521) );
  NOR2_X1 U12122 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9516) );
  NOR2_X1 U12123 ( .A1(n9633), .A2(n9516), .ZN(n9643) );
  NAND2_X1 U12124 ( .A1(n11590), .A2(n9643), .ZN(n9520) );
  NAND2_X1 U12125 ( .A1(n11591), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9519) );
  NAND2_X1 U12126 ( .A1(n9355), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9518) );
  NAND4_X1 U12127 ( .A1(n9521), .A2(n9520), .A3(n9519), .A4(n9518), .ZN(n12780) );
  NAND2_X1 U12128 ( .A1(n12780), .A2(n12824), .ZN(n9523) );
  NAND2_X1 U12129 ( .A1(n12782), .A2(n12754), .ZN(n9522) );
  NAND2_X1 U12130 ( .A1(n9523), .A2(n9522), .ZN(n14578) );
  AOI22_X1 U12131 ( .A1(n12757), .A2(n14578), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9524) );
  OAI21_X1 U12132 ( .B1(n12761), .B2(n10118), .A(n9524), .ZN(n9525) );
  AOI21_X1 U12133 ( .B1(n12758), .B2(n10063), .A(n9525), .ZN(n9526) );
  OAI21_X1 U12134 ( .B1(n9527), .B2(n12749), .A(n9526), .ZN(P2_U3190) );
  INV_X1 U12135 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n14939) );
  NAND2_X1 U12136 ( .A1(n11980), .A2(P3_U3897), .ZN(n9528) );
  OAI21_X1 U12137 ( .B1(P3_U3897), .B2(n14939), .A(n9528), .ZN(P3_U3504) );
  OAI21_X1 U12138 ( .B1(n9531), .B2(n9530), .A(n9529), .ZN(n9540) );
  INV_X1 U12139 ( .A(n14276), .ZN(n14231) );
  NOR2_X1 U12140 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9532), .ZN(n10902) );
  AOI21_X1 U12141 ( .B1(n9607), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n10902), .ZN(
        n9537) );
  OAI211_X1 U12142 ( .C1(n9535), .C2(n9534), .A(n14280), .B(n9533), .ZN(n9536)
         );
  OAI211_X1 U12143 ( .C1(n14231), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9539)
         );
  AOI21_X1 U12144 ( .B1(n14226), .B2(n9540), .A(n9539), .ZN(n9541) );
  INV_X1 U12145 ( .A(n9541), .ZN(P1_U3252) );
  OR2_X1 U12146 ( .A1(n9846), .A2(n9543), .ZN(n13965) );
  INV_X1 U12147 ( .A(n9838), .ZN(n9839) );
  AOI21_X1 U12148 ( .B1(n9839), .B2(n13838), .A(n13486), .ZN(n9545) );
  NAND2_X1 U12149 ( .A1(n9545), .A2(n11856), .ZN(n10571) );
  INV_X1 U12150 ( .A(n9546), .ZN(n9547) );
  NAND2_X1 U12151 ( .A1(n9547), .A2(n10494), .ZN(n14400) );
  NAND2_X1 U12152 ( .A1(n13838), .A2(n13486), .ZN(n9549) );
  OR2_X1 U12153 ( .A1(n11869), .A2(n10494), .ZN(n9548) );
  INV_X1 U12154 ( .A(n13723), .ZN(n9550) );
  AOI21_X1 U12155 ( .B1(n14368), .B2(n14379), .A(n9550), .ZN(n9551) );
  AOI211_X1 U12156 ( .C1(n10390), .C2(n13724), .A(n13726), .B(n9551), .ZN(
        n9652) );
  NOR4_X1 U12157 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_17__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n9555) );
  NOR4_X1 U12158 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n9554) );
  NOR4_X1 U12159 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9553) );
  NOR4_X1 U12160 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9552) );
  NAND4_X1 U12161 ( .A1(n9555), .A2(n9554), .A3(n9553), .A4(n9552), .ZN(n9561)
         );
  NOR2_X1 U12162 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .ZN(
        n9559) );
  NOR4_X1 U12163 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n9558) );
  NOR4_X1 U12164 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n9557) );
  NOR4_X1 U12165 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n9556) );
  NAND4_X1 U12166 ( .A1(n9559), .A2(n9558), .A3(n9557), .A4(n9556), .ZN(n9560)
         );
  NOR2_X1 U12167 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  OR2_X1 U12168 ( .A1(n9566), .A2(n9562), .ZN(n9851) );
  NAND2_X1 U12169 ( .A1(n9851), .A2(n10364), .ZN(n10357) );
  OR2_X1 U12170 ( .A1(n9566), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9565) );
  OR2_X1 U12171 ( .A1(n9234), .A2(n9563), .ZN(n9564) );
  NAND2_X1 U12172 ( .A1(n9850), .A2(n10358), .ZN(n9837) );
  OR2_X1 U12173 ( .A1(n9566), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U12174 ( .A1(n9233), .A2(n13835), .ZN(n9567) );
  INV_X1 U12175 ( .A(n10359), .ZN(n9848) );
  NAND2_X2 U12176 ( .A1(n10390), .A2(n10494), .ZN(n14352) );
  NAND2_X1 U12177 ( .A1(n9848), .A2(n10362), .ZN(n9569) );
  NAND2_X1 U12178 ( .A1(n14438), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9570) );
  OAI21_X1 U12179 ( .B1(n9652), .B2(n14438), .A(n9570), .ZN(P1_U3528) );
  NAND3_X1 U12180 ( .A1(n14566), .A2(n9572), .A3(n9571), .ZN(n10053) );
  NAND2_X1 U12181 ( .A1(n14565), .A2(n9573), .ZN(n9574) );
  OR2_X1 U12182 ( .A1(n10053), .A2(n9574), .ZN(n9586) );
  INV_X1 U12183 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9584) );
  INV_X1 U12184 ( .A(n14630), .ZN(n14641) );
  NAND2_X1 U12185 ( .A1(n10043), .A2(n11294), .ZN(n10058) );
  NAND2_X1 U12186 ( .A1(n11293), .A2(n10042), .ZN(n9576) );
  NAND2_X1 U12187 ( .A1(n11289), .A2(n14545), .ZN(n11645) );
  NAND2_X1 U12188 ( .A1(n9330), .A2(n11646), .ZN(n9578) );
  NAND2_X1 U12189 ( .A1(n9331), .A2(n11680), .ZN(n11611) );
  NAND2_X2 U12190 ( .A1(n9578), .A2(n11611), .ZN(n14548) );
  AOI21_X1 U12191 ( .B1(n9580), .B2(n14548), .A(n9579), .ZN(n10157) );
  NAND2_X1 U12192 ( .A1(n14545), .A2(n11294), .ZN(n9581) );
  AND3_X1 U12193 ( .A1(n10163), .A2(n12952), .A3(n9581), .ZN(n10159) );
  AOI21_X1 U12194 ( .B1(n14637), .B2(n11294), .A(n10159), .ZN(n9582) );
  OAI211_X1 U12195 ( .C1(n14583), .C2(n10162), .A(n10157), .B(n9582), .ZN(
        n9587) );
  NAND2_X1 U12196 ( .A1(n14663), .A2(n9587), .ZN(n9583) );
  OAI21_X1 U12197 ( .B1(n14663), .B2(n9584), .A(n9583), .ZN(P2_U3500) );
  INV_X1 U12198 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9589) );
  NAND2_X1 U12199 ( .A1(n14648), .A2(n9587), .ZN(n9588) );
  OAI21_X1 U12200 ( .B1(n14648), .B2(n9589), .A(n9588), .ZN(P2_U3433) );
  INV_X1 U12201 ( .A(n9590), .ZN(n9593) );
  OAI222_X1 U12202 ( .A1(n12657), .A2(n9593), .B1(n12661), .B2(n9592), .C1(
        n9591), .C2(P3_U3151), .ZN(P3_U3278) );
  NAND2_X1 U12203 ( .A1(n13451), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9594) );
  OR2_X1 U12204 ( .A1(n13451), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n13469) );
  NAND2_X1 U12205 ( .A1(n9594), .A2(n13469), .ZN(n9599) );
  NAND2_X1 U12206 ( .A1(n9601), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9595) );
  NAND2_X1 U12207 ( .A1(n9596), .A2(n9595), .ZN(n9598) );
  OR2_X1 U12208 ( .A1(n9598), .A2(n9599), .ZN(n13470) );
  INV_X1 U12209 ( .A(n13470), .ZN(n9597) );
  AOI21_X1 U12210 ( .B1(n9599), .B2(n9598), .A(n9597), .ZN(n9614) );
  INV_X1 U12211 ( .A(n14280), .ZN(n9613) );
  INV_X1 U12212 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9600) );
  MUX2_X1 U12213 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9600), .S(n13451), .Z(
        n9605) );
  OR2_X1 U12214 ( .A1(n9601), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U12215 ( .A1(n9603), .A2(n9602), .ZN(n9604) );
  NAND2_X1 U12216 ( .A1(n9604), .A2(n9605), .ZN(n13453) );
  OAI21_X1 U12217 ( .B1(n9605), .B2(n9604), .A(n13453), .ZN(n9611) );
  INV_X1 U12218 ( .A(n13451), .ZN(n9609) );
  NOR2_X1 U12219 ( .A1(n9606), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11138) );
  AOI21_X1 U12220 ( .B1(n9607), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n11138), .ZN(
        n9608) );
  OAI21_X1 U12221 ( .B1(n14231), .B2(n9609), .A(n9608), .ZN(n9610) );
  AOI21_X1 U12222 ( .B1(n9611), .B2(n14226), .A(n9610), .ZN(n9612) );
  OAI21_X1 U12223 ( .B1(n9614), .B2(n9613), .A(n9612), .ZN(P1_U3255) );
  INV_X1 U12224 ( .A(n9615), .ZN(n9618) );
  INV_X1 U12225 ( .A(n9616), .ZN(n9617) );
  NAND2_X1 U12226 ( .A1(n9618), .A2(n9617), .ZN(n9619) );
  NAND2_X1 U12227 ( .A1(n9622), .A2(n11584), .ZN(n9625) );
  AOI22_X1 U12228 ( .A1(n11434), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n11433), 
        .B2(n9623), .ZN(n9624) );
  NAND2_X1 U12229 ( .A1(n9625), .A2(n9624), .ZN(n11325) );
  XNOR2_X1 U12230 ( .A(n9510), .B(n11325), .ZN(n9627) );
  AND2_X1 U12231 ( .A1(n12780), .A2(n9339), .ZN(n9626) );
  OR2_X1 U12232 ( .A1(n9627), .A2(n9626), .ZN(n9803) );
  NAND2_X1 U12233 ( .A1(n9627), .A2(n9626), .ZN(n9628) );
  NAND2_X1 U12234 ( .A1(n9803), .A2(n9628), .ZN(n9631) );
  INV_X1 U12235 ( .A(n9804), .ZN(n9630) );
  AOI21_X1 U12236 ( .B1(n9632), .B2(n9631), .A(n9630), .ZN(n9647) );
  NAND2_X1 U12237 ( .A1(n9354), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9638) );
  NAND2_X1 U12238 ( .A1(n9633), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9808) );
  OAI21_X1 U12239 ( .B1(n9633), .B2(P2_REG3_REG_5__SCAN_IN), .A(n9808), .ZN(
        n10141) );
  INV_X1 U12240 ( .A(n10141), .ZN(n9634) );
  NAND2_X1 U12241 ( .A1(n11590), .A2(n9634), .ZN(n9637) );
  NAND2_X1 U12242 ( .A1(n11591), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12243 ( .A1(n11612), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9635) );
  NAND4_X1 U12244 ( .A1(n9638), .A2(n9637), .A3(n9636), .A4(n9635), .ZN(n12779) );
  NAND2_X1 U12245 ( .A1(n12779), .A2(n12824), .ZN(n9640) );
  NAND2_X1 U12246 ( .A1(n12781), .A2(n12754), .ZN(n9639) );
  NAND2_X1 U12247 ( .A1(n9640), .A2(n9639), .ZN(n10130) );
  INV_X1 U12248 ( .A(n10130), .ZN(n9642) );
  OAI21_X1 U12249 ( .B1(n12744), .B2(n9642), .A(n9641), .ZN(n9645) );
  INV_X1 U12250 ( .A(n9643), .ZN(n10122) );
  NOR2_X1 U12251 ( .A1(n12742), .A2(n10122), .ZN(n9644) );
  AOI211_X1 U12252 ( .C1(n11325), .C2(n12747), .A(n9645), .B(n9644), .ZN(n9646) );
  OAI21_X1 U12253 ( .B1(n9647), .B2(n12749), .A(n9646), .ZN(P2_U3202) );
  INV_X1 U12254 ( .A(n11168), .ZN(n9696) );
  AOI22_X1 U12255 ( .A1(n14239), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n13819), .ZN(n9648) );
  OAI21_X1 U12256 ( .B1(n9696), .B2(n13837), .A(n9648), .ZN(P1_U3339) );
  NAND2_X1 U12257 ( .A1(n10362), .A2(n10358), .ZN(n9649) );
  NOR2_X1 U12258 ( .A1(n10359), .A2(n10357), .ZN(n9650) );
  INV_X1 U12259 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9654) );
  OR2_X1 U12260 ( .A1(n9652), .A2(n14423), .ZN(n9653) );
  OAI21_X1 U12261 ( .B1(n14425), .B2(n9654), .A(n9653), .ZN(P1_U3459) );
  INV_X1 U12262 ( .A(n10942), .ZN(n9722) );
  AOI22_X1 U12263 ( .A1(n14211), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n13819), .ZN(n9655) );
  OAI21_X1 U12264 ( .B1(n9722), .B2(n13837), .A(n9655), .ZN(P1_U3341) );
  XOR2_X1 U12265 ( .A(n9657), .B(n9656), .Z(n9669) );
  INV_X1 U12266 ( .A(n14719), .ZN(n14686) );
  AOI22_X1 U12267 ( .A1(n14664), .A2(P3_ADDR_REG_3__SCAN_IN), .B1(
        P3_REG3_REG_3__SCAN_IN), .B2(P3_U3151), .ZN(n9665) );
  NAND2_X1 U12268 ( .A1(n9658), .A2(n14904), .ZN(n9659) );
  NAND2_X1 U12269 ( .A1(n9771), .A2(n9659), .ZN(n9660) );
  NAND2_X1 U12270 ( .A1(n14040), .A2(n9660), .ZN(n9664) );
  XNOR2_X1 U12271 ( .A(n9661), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12272 ( .A1(n14703), .A2(n9662), .ZN(n9663) );
  NAND3_X1 U12273 ( .A1(n9665), .A2(n9664), .A3(n9663), .ZN(n9666) );
  AOI21_X1 U12274 ( .B1(n14686), .B2(n9667), .A(n9666), .ZN(n9668) );
  OAI21_X1 U12275 ( .B1(n9669), .B2(n14036), .A(n9668), .ZN(P3_U3185) );
  INV_X1 U12276 ( .A(n14036), .ZN(n14713) );
  NOR3_X1 U12277 ( .A1(n14040), .A2(n14703), .A3(n14713), .ZN(n9680) );
  INV_X1 U12278 ( .A(n9670), .ZN(n9740) );
  INV_X1 U12279 ( .A(n14664), .ZN(n14724) );
  INV_X1 U12280 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n9671) );
  OAI22_X1 U12281 ( .A1(n14724), .A2(n9671), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9956), .ZN(n9674) );
  INV_X1 U12282 ( .A(n14703), .ZN(n9767) );
  NOR2_X1 U12283 ( .A1(n9767), .A2(n9672), .ZN(n9673) );
  AOI211_X1 U12284 ( .C1(n9675), .C2(n14040), .A(n9674), .B(n9673), .ZN(n9679)
         );
  OR2_X1 U12285 ( .A1(n9676), .A2(n14036), .ZN(n9677) );
  MUX2_X1 U12286 ( .A(n9677), .B(n14719), .S(P3_IR_REG_0__SCAN_IN), .Z(n9678)
         );
  OAI211_X1 U12287 ( .C1(n9680), .C2(n9740), .A(n9679), .B(n9678), .ZN(
        P3_U3182) );
  INV_X1 U12288 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9682) );
  MUX2_X1 U12289 ( .A(n9682), .B(P2_REG1_REG_7__SCAN_IN), .S(n10002), .Z(n9683) );
  AOI211_X1 U12290 ( .C1(n9684), .C2(n9683), .A(n14531), .B(n10001), .ZN(n9692) );
  XNOR2_X1 U12291 ( .A(n10002), .B(P2_REG2_REG_7__SCAN_IN), .ZN(n9686) );
  AOI211_X1 U12292 ( .C1(n9687), .C2(n9686), .A(n14527), .B(n9991), .ZN(n9691)
         );
  INV_X1 U12293 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13909) );
  NAND2_X1 U12294 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n9689) );
  NAND2_X1 U12295 ( .A1(n14537), .A2(n10002), .ZN(n9688) );
  OAI211_X1 U12296 ( .C1(n14540), .C2(n13909), .A(n9689), .B(n9688), .ZN(n9690) );
  OR3_X1 U12297 ( .A1(n9692), .A2(n9691), .A3(n9690), .ZN(P2_U3221) );
  NAND2_X1 U12298 ( .A1(n9693), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9937) );
  NAND2_X1 U12299 ( .A1(n9937), .A2(n9936), .ZN(n9694) );
  NAND2_X1 U12300 ( .A1(n9694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9695) );
  INV_X1 U12301 ( .A(n14522), .ZN(n9697) );
  OAI222_X1 U12302 ( .A1(P2_U3088), .A2(n9697), .B1(n13213), .B2(n9696), .C1(
        n11169), .C2(n13210), .ZN(P2_U3311) );
  INV_X1 U12303 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9718) );
  NAND2_X1 U12304 ( .A1(n10570), .A2(n10569), .ZN(n10568) );
  INV_X1 U12305 ( .A(n13353), .ZN(n10615) );
  NAND2_X1 U12306 ( .A1(n6815), .A2(n10615), .ZN(n9699) );
  NAND2_X1 U12307 ( .A1(n10568), .A2(n9699), .ZN(n9701) );
  NAND2_X1 U12308 ( .A1(n9701), .A2(n9700), .ZN(n10369) );
  OR2_X1 U12309 ( .A1(n9701), .A2(n9700), .ZN(n9702) );
  NAND2_X1 U12310 ( .A1(n10369), .A2(n9702), .ZN(n14307) );
  INV_X1 U12311 ( .A(n14307), .ZN(n9716) );
  NAND2_X1 U12312 ( .A1(n9704), .A2(n9703), .ZN(n9706) );
  NAND2_X1 U12313 ( .A1(n9706), .A2(n9705), .ZN(n10567) );
  NAND2_X1 U12314 ( .A1(n10567), .A2(n9707), .ZN(n9709) );
  NAND2_X1 U12315 ( .A1(n10615), .A2(n10577), .ZN(n9708) );
  NAND2_X1 U12316 ( .A1(n9709), .A2(n9708), .ZN(n10376) );
  XNOR2_X1 U12317 ( .A(n10376), .B(n10375), .ZN(n9712) );
  OR2_X1 U12318 ( .A1(n10370), .A2(n13965), .ZN(n9711) );
  NAND2_X1 U12319 ( .A1(n13353), .A2(n14087), .ZN(n9710) );
  NAND2_X1 U12320 ( .A1(n9711), .A2(n9710), .ZN(n9912) );
  AOI21_X1 U12321 ( .B1(n9712), .B2(n14373), .A(n9912), .ZN(n14321) );
  OR2_X1 U12322 ( .A1(n10580), .A2(n10367), .ZN(n9714) );
  AND3_X1 U12323 ( .A1(n10649), .A2(n9843), .A3(n9714), .ZN(n14312) );
  AOI21_X1 U12324 ( .B1(n14397), .B2(n14309), .A(n14312), .ZN(n9715) );
  OAI211_X1 U12325 ( .C1(n9716), .C2(n14368), .A(n14321), .B(n9715), .ZN(n9821) );
  NAND2_X1 U12326 ( .A1(n9821), .A2(n14425), .ZN(n9717) );
  OAI21_X1 U12327 ( .B1(n14425), .B2(n9718), .A(n9717), .ZN(P1_U3468) );
  NAND2_X1 U12328 ( .A1(n9719), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9720) );
  XNOR2_X1 U12329 ( .A(n9720), .B(P2_IR_REG_14__SCAN_IN), .ZN(n14497) );
  INV_X1 U12330 ( .A(n14497), .ZN(n12786) );
  OAI222_X1 U12331 ( .A1(P2_U3088), .A2(n12786), .B1(n13213), .B2(n9722), .C1(
        n9721), .C2(n13210), .ZN(P2_U3313) );
  XOR2_X1 U12332 ( .A(n9724), .B(n9723), .Z(n9739) );
  OAI21_X1 U12333 ( .B1(n9727), .B2(n9726), .A(n9725), .ZN(n9737) );
  OAI21_X1 U12334 ( .B1(n9730), .B2(n9729), .A(n9728), .ZN(n9731) );
  NAND2_X1 U12335 ( .A1(n14703), .A2(n9731), .ZN(n9733) );
  NAND2_X1 U12336 ( .A1(n14664), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n9732) );
  OAI211_X1 U12337 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10019), .A(n9733), .B(
        n9732), .ZN(n9736) );
  NOR2_X1 U12338 ( .A1(n14719), .A2(n9734), .ZN(n9735) );
  AOI211_X1 U12339 ( .C1(n14040), .C2(n9737), .A(n9736), .B(n9735), .ZN(n9738)
         );
  OAI21_X1 U12340 ( .B1(n9739), .B2(n14036), .A(n9738), .ZN(P3_U3184) );
  XNOR2_X1 U12341 ( .A(n9741), .B(n9740), .ZN(n9757) );
  NAND2_X1 U12342 ( .A1(n9742), .A2(n14790), .ZN(n9743) );
  NAND2_X1 U12343 ( .A1(n9744), .A2(n9743), .ZN(n9755) );
  NAND2_X1 U12344 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  NAND2_X1 U12345 ( .A1(n9748), .A2(n9747), .ZN(n9749) );
  NAND2_X1 U12346 ( .A1(n14703), .A2(n9749), .ZN(n9751) );
  NAND2_X1 U12347 ( .A1(n14664), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n9750) );
  OAI211_X1 U12348 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n14786), .A(n9751), .B(
        n9750), .ZN(n9754) );
  NOR2_X1 U12349 ( .A1(n14719), .A2(n9752), .ZN(n9753) );
  AOI211_X1 U12350 ( .C1(n14040), .C2(n9755), .A(n9754), .B(n9753), .ZN(n9756)
         );
  OAI21_X1 U12351 ( .B1(n14036), .B2(n9757), .A(n9756), .ZN(P3_U3183) );
  OAI222_X1 U12352 ( .A1(P3_U3151), .A2(n12055), .B1(n12661), .B2(n9759), .C1(
        n12657), .C2(n9758), .ZN(P3_U3276) );
  XOR2_X1 U12353 ( .A(n9761), .B(n9760), .Z(n9778) );
  AOI21_X1 U12354 ( .B1(n9764), .B2(n9763), .A(n9762), .ZN(n9766) );
  AND2_X1 U12355 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10354) );
  AOI21_X1 U12356 ( .B1(n14664), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10354), .ZN(
        n9765) );
  OAI21_X1 U12357 ( .B1(n9767), .B2(n9766), .A(n9765), .ZN(n9775) );
  INV_X1 U12358 ( .A(n9768), .ZN(n9770) );
  NAND3_X1 U12359 ( .A1(n9771), .A2(n9770), .A3(n9769), .ZN(n9772) );
  AOI21_X1 U12360 ( .B1(n9773), .B2(n9772), .A(n14708), .ZN(n9774) );
  AOI211_X1 U12361 ( .C1(n14686), .C2(n9776), .A(n9775), .B(n9774), .ZN(n9777)
         );
  OAI21_X1 U12362 ( .B1(n9778), .B2(n14036), .A(n9777), .ZN(P3_U3186) );
  XOR2_X1 U12363 ( .A(n9780), .B(n9779), .Z(n9792) );
  XOR2_X1 U12364 ( .A(P3_REG1_REG_5__SCAN_IN), .B(n9781), .Z(n9790) );
  AND2_X1 U12365 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10458) );
  AOI21_X1 U12366 ( .B1(n14664), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10458), .ZN(
        n9787) );
  NAND2_X1 U12367 ( .A1(n9783), .A2(n9782), .ZN(n9784) );
  NAND2_X1 U12368 ( .A1(n9925), .A2(n9784), .ZN(n9785) );
  NAND2_X1 U12369 ( .A1(n14040), .A2(n9785), .ZN(n9786) );
  OAI211_X1 U12370 ( .C1(n14719), .C2(n9788), .A(n9787), .B(n9786), .ZN(n9789)
         );
  AOI21_X1 U12371 ( .B1(n14703), .B2(n9790), .A(n9789), .ZN(n9791) );
  OAI21_X1 U12372 ( .B1(n9792), .B2(n14036), .A(n9791), .ZN(P3_U3187) );
  INV_X1 U12373 ( .A(n11408), .ZN(n9835) );
  INV_X1 U12374 ( .A(n14258), .ZN(n9794) );
  OAI222_X1 U12375 ( .A1(n13837), .A2(n9835), .B1(n9794), .B2(P1_U3086), .C1(
        n9793), .C2(n13833), .ZN(P1_U3338) );
  NAND2_X1 U12376 ( .A1(n9795), .A2(n11584), .ZN(n9797) );
  AOI22_X1 U12377 ( .A1(n11434), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n11433), 
        .B2(n14463), .ZN(n9796) );
  NAND2_X1 U12378 ( .A1(n9797), .A2(n9796), .ZN(n11331) );
  XNOR2_X1 U12379 ( .A(n11331), .B(n11724), .ZN(n9798) );
  NAND2_X1 U12380 ( .A1(n12779), .A2(n9339), .ZN(n9799) );
  NAND2_X1 U12381 ( .A1(n9798), .A2(n9799), .ZN(n9857) );
  INV_X1 U12382 ( .A(n9798), .ZN(n9801) );
  INV_X1 U12383 ( .A(n9799), .ZN(n9800) );
  NAND2_X1 U12384 ( .A1(n9801), .A2(n9800), .ZN(n9802) );
  AND2_X1 U12385 ( .A1(n9857), .A2(n9802), .ZN(n9806) );
  OAI21_X1 U12386 ( .B1(n9806), .B2(n9805), .A(n9858), .ZN(n9819) );
  NOR2_X1 U12387 ( .A1(n12742), .A2(n10141), .ZN(n9818) );
  NAND2_X1 U12388 ( .A1(n11591), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U12389 ( .A1(n9354), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9812) );
  INV_X1 U12390 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n9807) );
  AND2_X1 U12391 ( .A1(n9808), .A2(n9807), .ZN(n9809) );
  NOR2_X1 U12392 ( .A1(n9865), .A2(n9809), .ZN(n9863) );
  NAND2_X1 U12393 ( .A1(n11590), .A2(n9863), .ZN(n9811) );
  NAND2_X1 U12394 ( .A1(n11612), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9810) );
  NAND4_X1 U12395 ( .A1(n9813), .A2(n9812), .A3(n9811), .A4(n9810), .ZN(n12778) );
  NAND2_X1 U12396 ( .A1(n12778), .A2(n12824), .ZN(n9815) );
  NAND2_X1 U12397 ( .A1(n12780), .A2(n12754), .ZN(n9814) );
  AND2_X1 U12398 ( .A1(n9815), .A2(n9814), .ZN(n10152) );
  NAND2_X1 U12399 ( .A1(n12747), .A2(n11331), .ZN(n9816) );
  NAND2_X1 U12400 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14464) );
  OAI211_X1 U12401 ( .C1(n10152), .C2(n12744), .A(n9816), .B(n14464), .ZN(
        n9817) );
  AOI211_X1 U12402 ( .C1(n9819), .C2(n12763), .A(n9818), .B(n9817), .ZN(n9820)
         );
  INV_X1 U12403 ( .A(n9820), .ZN(P2_U3199) );
  NAND2_X1 U12404 ( .A1(n9821), .A2(n14441), .ZN(n9822) );
  OAI21_X1 U12405 ( .B1(n14441), .B2(n9823), .A(n9822), .ZN(P1_U3531) );
  AND2_X1 U12406 ( .A1(n9825), .A2(n9824), .ZN(n9832) );
  INV_X1 U12407 ( .A(n9832), .ZN(n9826) );
  OAI21_X1 U12408 ( .B1(n9827), .B2(n9826), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9828) );
  INV_X1 U12409 ( .A(n9829), .ZN(n9831) );
  NAND3_X1 U12410 ( .A1(n9832), .A2(n9831), .A3(n9830), .ZN(n10068) );
  INV_X1 U12411 ( .A(n14536), .ZN(n9836) );
  OAI222_X1 U12412 ( .A1(P2_U3088), .A2(n9836), .B1(n13213), .B2(n9835), .C1(
        n9834), .C2(n13210), .ZN(P2_U3310) );
  INV_X1 U12413 ( .A(n13334), .ZN(n10337) );
  NAND2_X1 U12414 ( .A1(n10337), .A2(n6454), .ZN(n13313) );
  INV_X1 U12415 ( .A(n13313), .ZN(n14074) );
  INV_X1 U12416 ( .A(n9908), .ZN(n9844) );
  NAND2_X1 U12417 ( .A1(n9844), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n9842) );
  AOI22_X1 U12418 ( .A1(n6452), .A2(n13724), .B1(n9844), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n9845) );
  OAI21_X1 U12419 ( .B1(n11815), .B2(n9840), .A(n9845), .ZN(n9879) );
  XOR2_X1 U12420 ( .A(n9880), .B(n9879), .Z(n13370) );
  NAND2_X1 U12421 ( .A1(n14417), .A2(n9846), .ZN(n9847) );
  NOR2_X1 U12422 ( .A1(n9848), .A2(n9847), .ZN(n9849) );
  AOI22_X1 U12423 ( .A1(n14074), .A2(n13354), .B1(n13370), .B2(n13320), .ZN(
        n9856) );
  NAND3_X1 U12424 ( .A1(n9852), .A2(n10359), .A3(n9851), .ZN(n9853) );
  NAND2_X1 U12425 ( .A1(n9853), .A2(n10362), .ZN(n9909) );
  AND2_X1 U12426 ( .A1(n9909), .A2(n10364), .ZN(n9854) );
  NAND2_X1 U12427 ( .A1(n9854), .A2(n10358), .ZN(n9896) );
  AOI22_X1 U12428 ( .A1(n14075), .A2(n13724), .B1(n9896), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n9855) );
  NAND2_X1 U12429 ( .A1(n9856), .A2(n9855), .ZN(P1_U3232) );
  NAND2_X1 U12430 ( .A1(n9859), .A2(n11584), .ZN(n9862) );
  AOI22_X1 U12431 ( .A1(n11434), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n11433), 
        .B2(n9860), .ZN(n9861) );
  XNOR2_X1 U12432 ( .A(n14601), .B(n11724), .ZN(n9972) );
  NAND2_X1 U12433 ( .A1(n12778), .A2(n9339), .ZN(n9973) );
  XNOR2_X1 U12434 ( .A(n9972), .B(n9973), .ZN(n9971) );
  XNOR2_X1 U12435 ( .A(n9970), .B(n9971), .ZN(n9877) );
  INV_X1 U12436 ( .A(n9863), .ZN(n10210) );
  NAND2_X1 U12437 ( .A1(n9864), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12438 ( .A1(n9865), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9981) );
  OR2_X1 U12439 ( .A1(n9865), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9866) );
  AND2_X1 U12440 ( .A1(n9981), .A2(n9866), .ZN(n10290) );
  NAND2_X1 U12441 ( .A1(n11590), .A2(n10290), .ZN(n9869) );
  NAND2_X1 U12442 ( .A1(n11591), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9868) );
  NAND2_X1 U12443 ( .A1(n11612), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9867) );
  NAND4_X1 U12444 ( .A1(n9870), .A2(n9869), .A3(n9868), .A4(n9867), .ZN(n12777) );
  NAND2_X1 U12445 ( .A1(n12777), .A2(n12824), .ZN(n9872) );
  NAND2_X1 U12446 ( .A1(n12779), .A2(n12754), .ZN(n9871) );
  NAND2_X1 U12447 ( .A1(n9872), .A2(n9871), .ZN(n10208) );
  NAND2_X1 U12448 ( .A1(n12757), .A2(n10208), .ZN(n9874) );
  OAI211_X1 U12449 ( .C1(n12742), .C2(n10210), .A(n9874), .B(n9873), .ZN(n9875) );
  AOI21_X1 U12450 ( .B1(n14601), .B2(n12747), .A(n9875), .ZN(n9876) );
  OAI21_X1 U12451 ( .B1(n9877), .B2(n12749), .A(n9876), .ZN(P2_U3211) );
  NAND2_X1 U12452 ( .A1(n9879), .A2(n9880), .ZN(n9883) );
  NAND2_X1 U12453 ( .A1(n9881), .A2(n11813), .ZN(n9882) );
  NAND2_X1 U12454 ( .A1(n9883), .A2(n9882), .ZN(n9884) );
  AOI21_X1 U12455 ( .B1(n9885), .B2(n9884), .A(n9893), .ZN(n9888) );
  INV_X1 U12456 ( .A(n14087), .ZN(n13963) );
  AOI22_X1 U12457 ( .A1(n14074), .A2(n13353), .B1(n14073), .B2(n13355), .ZN(
        n9887) );
  AOI22_X1 U12458 ( .A1(n14075), .A2(n10619), .B1(n9896), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n9886) );
  OAI211_X1 U12459 ( .C1(n9888), .C2(n14078), .A(n9887), .B(n9886), .ZN(
        P1_U3222) );
  OAI22_X1 U12460 ( .A1(n11815), .A2(n10615), .B1(n6815), .B2(n11823), .ZN(
        n9903) );
  AOI22_X1 U12461 ( .A1(n6452), .A2(n13353), .B1(n9889), .B2(n10577), .ZN(
        n9890) );
  XNOR2_X1 U12462 ( .A(n9890), .B(n11856), .ZN(n9902) );
  XOR2_X1 U12463 ( .A(n9903), .B(n9902), .Z(n9904) );
  INV_X1 U12464 ( .A(n9891), .ZN(n9895) );
  INV_X1 U12465 ( .A(n9892), .ZN(n9894) );
  XOR2_X1 U12466 ( .A(n9904), .B(n9905), .Z(n9899) );
  AOI22_X1 U12467 ( .A1(n14074), .A2(n13352), .B1(n14073), .B2(n13354), .ZN(
        n9898) );
  AOI22_X1 U12468 ( .A1(n14075), .A2(n10577), .B1(n9896), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n9897) );
  OAI211_X1 U12469 ( .C1(n9899), .C2(n14078), .A(n9898), .B(n9897), .ZN(
        P1_U3237) );
  INV_X1 U12470 ( .A(n11024), .ZN(n9938) );
  OAI222_X1 U12471 ( .A1(n13837), .A2(n9938), .B1(n14230), .B2(P1_U3086), .C1(
        n9900), .C2(n13833), .ZN(P1_U3340) );
  OAI22_X1 U12472 ( .A1(n10572), .A2(n11823), .B1(n11824), .B2(n10367), .ZN(
        n9901) );
  XNOR2_X1 U12473 ( .A(n9901), .B(n11856), .ZN(n10299) );
  OAI22_X1 U12474 ( .A1(n11815), .A2(n10572), .B1(n10367), .B2(n11823), .ZN(
        n10298) );
  XNOR2_X1 U12475 ( .A(n10299), .B(n10298), .ZN(n9907) );
  AOI211_X1 U12476 ( .C1(n9907), .C2(n9906), .A(n14078), .B(n6614), .ZN(n9916)
         );
  NAND3_X1 U12477 ( .A1(n9909), .A2(n9908), .A3(n10358), .ZN(n9910) );
  NAND2_X1 U12478 ( .A1(n9910), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9911) );
  AND2_X1 U12479 ( .A1(n9911), .A2(n10913), .ZN(n14083) );
  AOI22_X1 U12480 ( .A1(n10337), .A2(n9912), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n9914) );
  NAND2_X1 U12481 ( .A1(n14075), .A2(n14309), .ZN(n9913) );
  OAI211_X1 U12482 ( .C1(n14083), .C2(P1_REG3_REG_3__SCAN_IN), .A(n9914), .B(
        n9913), .ZN(n9915) );
  OR2_X1 U12483 ( .A1(n9916), .A2(n9915), .ZN(P1_U3218) );
  XOR2_X1 U12484 ( .A(n9918), .B(n9917), .Z(n9935) );
  OAI21_X1 U12485 ( .B1(n9921), .B2(n9920), .A(n9919), .ZN(n9933) );
  AND2_X1 U12486 ( .A1(P3_U3151), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n10729) );
  AOI21_X1 U12487 ( .B1(n14664), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10729), .ZN(
        n9930) );
  INV_X1 U12488 ( .A(n9922), .ZN(n9924) );
  NAND3_X1 U12489 ( .A1(n9925), .A2(n9924), .A3(n9923), .ZN(n9926) );
  NAND2_X1 U12490 ( .A1(n9927), .A2(n9926), .ZN(n9928) );
  NAND2_X1 U12491 ( .A1(n14040), .A2(n9928), .ZN(n9929) );
  OAI211_X1 U12492 ( .C1(n14719), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9932)
         );
  AOI21_X1 U12493 ( .B1(n14703), .B2(n9933), .A(n9932), .ZN(n9934) );
  OAI21_X1 U12494 ( .B1(n9935), .B2(n14036), .A(n9934), .ZN(P3_U3188) );
  XNOR2_X1 U12495 ( .A(n9937), .B(n9936), .ZN(n14501) );
  OAI222_X1 U12496 ( .A1(P2_U3088), .A2(n14501), .B1(n13213), .B2(n9938), .C1(
        n11025), .C2(n13210), .ZN(P2_U3312) );
  INV_X1 U12497 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n14924) );
  NAND2_X1 U12498 ( .A1(n12281), .A2(n9952), .ZN(n12072) );
  INV_X1 U12499 ( .A(n12072), .ZN(n9939) );
  NOR2_X1 U12500 ( .A1(n14775), .A2(n9939), .ZN(n12220) );
  INV_X1 U12501 ( .A(n9940), .ZN(n9941) );
  NOR3_X1 U12502 ( .A1(n12220), .A2(n14821), .A3(n9941), .ZN(n9942) );
  AOI21_X1 U12503 ( .B1(n14730), .B2(n9045), .A(n9942), .ZN(n10021) );
  OAI21_X1 U12504 ( .B1(n9952), .B2(n14837), .A(n10021), .ZN(n12549) );
  NAND2_X1 U12505 ( .A1(n12549), .A2(n14851), .ZN(n9943) );
  OAI21_X1 U12506 ( .B1(n14851), .B2(n14924), .A(n9943), .ZN(P3_U3390) );
  NOR2_X1 U12507 ( .A1(n9944), .A2(P3_U3151), .ZN(n10020) );
  INV_X1 U12508 ( .A(n14775), .ZN(n12070) );
  NAND3_X1 U12509 ( .A1(n12070), .A2(n9945), .A3(n11268), .ZN(n9946) );
  OAI211_X1 U12510 ( .C1(n6625), .C2(n14776), .A(n9947), .B(n9946), .ZN(n9948)
         );
  NAND2_X1 U12511 ( .A1(n9948), .A2(n14668), .ZN(n9951) );
  NAND2_X1 U12512 ( .A1(n12281), .A2(n14731), .ZN(n9949) );
  OAI21_X1 U12513 ( .B1(n10463), .B2(n14760), .A(n9949), .ZN(n14777) );
  AOI22_X1 U12514 ( .A1(n12019), .A2(n14777), .B1(n14675), .B2(n14781), .ZN(
        n9950) );
  OAI211_X1 U12515 ( .C1(n10020), .C2(n14786), .A(n9951), .B(n9950), .ZN(
        P3_U3162) );
  INV_X1 U12516 ( .A(n12220), .ZN(n9954) );
  NAND2_X1 U12517 ( .A1(n12019), .A2(n14730), .ZN(n12000) );
  INV_X1 U12518 ( .A(n14675), .ZN(n12006) );
  OAI22_X1 U12519 ( .A1(n12000), .A2(n14763), .B1(n12006), .B2(n9952), .ZN(
        n9953) );
  AOI21_X1 U12520 ( .B1(n14668), .B2(n9954), .A(n9953), .ZN(n9955) );
  OAI21_X1 U12521 ( .B1(n10020), .B2(n9956), .A(n9955), .ZN(P3_U3172) );
  XOR2_X1 U12522 ( .A(n9958), .B(n9957), .Z(n9969) );
  XOR2_X1 U12523 ( .A(P3_REG1_REG_7__SCAN_IN), .B(n9959), .Z(n9967) );
  AOI21_X1 U12524 ( .B1(n10830), .B2(n9961), .A(n9960), .ZN(n9962) );
  NOR2_X1 U12525 ( .A1(n9962), .A2(n14708), .ZN(n9966) );
  NAND2_X1 U12526 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n14665) );
  NAND2_X1 U12527 ( .A1(n14664), .A2(P3_ADDR_REG_7__SCAN_IN), .ZN(n9963) );
  OAI211_X1 U12528 ( .C1(n14719), .C2(n9964), .A(n14665), .B(n9963), .ZN(n9965) );
  AOI211_X1 U12529 ( .C1(n9967), .C2(n14703), .A(n9966), .B(n9965), .ZN(n9968)
         );
  OAI21_X1 U12530 ( .B1(n9969), .B2(n14036), .A(n9968), .ZN(P3_U3189) );
  INV_X1 U12531 ( .A(n9972), .ZN(n9975) );
  INV_X1 U12532 ( .A(n9973), .ZN(n9974) );
  NAND2_X1 U12533 ( .A1(n9975), .A2(n9974), .ZN(n9976) );
  OR2_X1 U12534 ( .A1(n9977), .A2(n11607), .ZN(n9979) );
  AOI22_X1 U12535 ( .A1(n11434), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n11433), 
        .B2(n10002), .ZN(n9978) );
  NAND2_X1 U12536 ( .A1(n9979), .A2(n9978), .ZN(n11347) );
  XNOR2_X1 U12537 ( .A(n11347), .B(n9510), .ZN(n10082) );
  NAND2_X1 U12538 ( .A1(n12777), .A2(n9339), .ZN(n10080) );
  XNOR2_X1 U12539 ( .A(n10082), .B(n10080), .ZN(n10083) );
  XNOR2_X1 U12540 ( .A(n10084), .B(n10083), .ZN(n9990) );
  INV_X1 U12541 ( .A(n11347), .ZN(n14610) );
  NAND2_X1 U12542 ( .A1(n9864), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9986) );
  NAND2_X1 U12543 ( .A1(n11591), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12544 ( .A1(n9981), .A2(n9980), .ZN(n9982) );
  AND2_X1 U12545 ( .A1(n10097), .A2(n9982), .ZN(n10259) );
  NAND2_X1 U12546 ( .A1(n11590), .A2(n10259), .ZN(n9984) );
  NAND2_X1 U12547 ( .A1(n11612), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9983) );
  NAND4_X1 U12548 ( .A1(n9986), .A2(n9985), .A3(n9984), .A4(n9983), .ZN(n12776) );
  INV_X1 U12549 ( .A(n12776), .ZN(n10239) );
  INV_X1 U12550 ( .A(n12778), .ZN(n11338) );
  INV_X1 U12551 ( .A(n12754), .ZN(n12848) );
  OAI22_X1 U12552 ( .A1(n10239), .A2(n12756), .B1(n11338), .B2(n12848), .ZN(
        n10284) );
  AOI22_X1 U12553 ( .A1(n12757), .A2(n10284), .B1(P2_REG3_REG_7__SCAN_IN), 
        .B2(P2_U3088), .ZN(n9987) );
  OAI21_X1 U12554 ( .B1(n12761), .B2(n14610), .A(n9987), .ZN(n9988) );
  AOI21_X1 U12555 ( .B1(n10290), .B2(n12758), .A(n9988), .ZN(n9989) );
  OAI21_X1 U12556 ( .B1(n9990), .B2(n12749), .A(n9989), .ZN(P2_U3185) );
  XNOR2_X1 U12557 ( .A(n14474), .B(P2_REG2_REG_8__SCAN_IN), .ZN(n14467) );
  INV_X1 U12558 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9992) );
  MUX2_X1 U12559 ( .A(n9992), .B(P2_REG2_REG_9__SCAN_IN), .S(n10528), .Z(n9993) );
  INV_X1 U12560 ( .A(n9993), .ZN(n9994) );
  OAI21_X1 U12561 ( .B1(n9995), .B2(n9994), .A(n10521), .ZN(n10000) );
  NAND2_X1 U12562 ( .A1(n14442), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n9996) );
  NAND2_X1 U12563 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3088), .ZN(n10200) );
  OAI211_X1 U12564 ( .C1(n12815), .C2(n9997), .A(n9996), .B(n10200), .ZN(n9998) );
  AOI21_X1 U12565 ( .B1(n10000), .B2(n9999), .A(n9998), .ZN(n10009) );
  INV_X1 U12566 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10003) );
  MUX2_X1 U12567 ( .A(n10003), .B(P2_REG1_REG_8__SCAN_IN), .S(n14474), .Z(
        n14470) );
  INV_X1 U12568 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10004) );
  MUX2_X1 U12569 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10004), .S(n10528), .Z(
        n10005) );
  OAI21_X1 U12570 ( .B1(n10006), .B2(n10005), .A(n10527), .ZN(n10007) );
  NAND2_X1 U12571 ( .A1(n10007), .A2(n12814), .ZN(n10008) );
  NAND2_X1 U12572 ( .A1(n10009), .A2(n10008), .ZN(P2_U3223) );
  XNOR2_X1 U12573 ( .A(n10011), .B(n10010), .ZN(n10012) );
  NAND2_X1 U12574 ( .A1(n10012), .A2(n14668), .ZN(n10018) );
  NOR2_X1 U12575 ( .A1(n14666), .A2(n14762), .ZN(n12003) );
  NAND2_X1 U12576 ( .A1(n12003), .A2(n9045), .ZN(n10015) );
  NAND2_X1 U12577 ( .A1(n14675), .A2(n10013), .ZN(n10014) );
  OAI211_X1 U12578 ( .C1(n12000), .C2(n14761), .A(n10015), .B(n10014), .ZN(
        n10016) );
  INV_X1 U12579 ( .A(n10016), .ZN(n10017) );
  OAI211_X1 U12580 ( .C1(n10020), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        P3_U3177) );
  MUX2_X1 U12581 ( .A(n10022), .B(n10021), .S(n14791), .Z(n10025) );
  AOI22_X1 U12582 ( .A1(n6433), .A2(n10023), .B1(P3_REG3_REG_0__SCAN_IN), .B2(
        n14772), .ZN(n10024) );
  NAND2_X1 U12583 ( .A1(n10025), .A2(n10024), .ZN(P3_U3233) );
  XOR2_X1 U12584 ( .A(n10026), .B(n10027), .Z(n10041) );
  OAI21_X1 U12585 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(n10039) );
  AOI21_X1 U12586 ( .B1(n6613), .B2(n10032), .A(n10031), .ZN(n10037) );
  NOR2_X1 U12587 ( .A1(n10033), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10841) );
  NOR2_X1 U12588 ( .A1(n14719), .A2(n10034), .ZN(n10035) );
  AOI211_X1 U12589 ( .C1(n14664), .C2(P3_ADDR_REG_8__SCAN_IN), .A(n10841), .B(
        n10035), .ZN(n10036) );
  OAI21_X1 U12590 ( .B1(n10037), .B2(n14708), .A(n10036), .ZN(n10038) );
  AOI21_X1 U12591 ( .B1(n10039), .B2(n14703), .A(n10038), .ZN(n10040) );
  OAI21_X1 U12592 ( .B1(n10041), .B2(n14036), .A(n10040), .ZN(P3_U3190) );
  INV_X1 U12593 ( .A(n11645), .ZN(n10045) );
  NAND2_X1 U12594 ( .A1(n10043), .A2(n10042), .ZN(n10044) );
  INV_X1 U12595 ( .A(n12782), .ZN(n10048) );
  NAND2_X1 U12596 ( .A1(n10048), .A2(n9363), .ZN(n10060) );
  NAND2_X1 U12597 ( .A1(n12782), .A2(n10046), .ZN(n10047) );
  INV_X1 U12598 ( .A(n11647), .ZN(n10165) );
  NAND2_X1 U12599 ( .A1(n10166), .A2(n10165), .ZN(n10050) );
  NAND2_X1 U12600 ( .A1(n10048), .A2(n10046), .ZN(n10049) );
  INV_X1 U12601 ( .A(n12781), .ZN(n10119) );
  NAND2_X1 U12602 ( .A1(n10119), .A2(n14579), .ZN(n10127) );
  NAND2_X1 U12603 ( .A1(n12781), .A2(n10118), .ZN(n10051) );
  XNOR2_X1 U12604 ( .A(n11648), .B(n10117), .ZN(n14582) );
  INV_X1 U12605 ( .A(n9575), .ZN(n14549) );
  NAND2_X1 U12606 ( .A1(n10052), .A2(n14562), .ZN(n10054) );
  OR2_X1 U12607 ( .A1(n10054), .A2(n10053), .ZN(n10055) );
  OAI211_X2 U12608 ( .C1(n11680), .C2(n14549), .A(n14554), .B(n11729), .ZN(
        n13081) );
  AOI211_X1 U12609 ( .C1(n14579), .C2(n10164), .A(n9339), .B(n10124), .ZN(
        n14577) );
  INV_X1 U12610 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10057) );
  OAI22_X1 U12611 ( .A1(n13076), .A2(n10118), .B1(n10057), .B2(n14554), .ZN(
        n10066) );
  NAND2_X1 U12612 ( .A1(n10059), .A2(n10058), .ZN(n10168) );
  NAND2_X1 U12613 ( .A1(n10168), .A2(n11647), .ZN(n10167) );
  NAND2_X1 U12614 ( .A1(n10167), .A2(n10060), .ZN(n10061) );
  NAND2_X1 U12615 ( .A1(n10061), .A2(n11648), .ZN(n10128) );
  OAI21_X1 U12616 ( .B1(n11648), .B2(n10061), .A(n10128), .ZN(n10062) );
  NAND2_X1 U12617 ( .A1(n10062), .A2(n14548), .ZN(n14580) );
  INV_X1 U12618 ( .A(n13071), .ZN(n14553) );
  AOI21_X1 U12619 ( .B1(n14553), .B2(n10063), .A(n14578), .ZN(n10064) );
  AOI21_X1 U12620 ( .B1(n14580), .B2(n10064), .A(n14557), .ZN(n10065) );
  AOI211_X1 U12621 ( .C1(n13078), .C2(n14577), .A(n10066), .B(n10065), .ZN(
        n10067) );
  OAI21_X1 U12622 ( .B1(n14582), .B2(n13081), .A(n10067), .ZN(P2_U3262) );
  NAND2_X1 U12623 ( .A1(n10068), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n10069) );
  XNOR2_X1 U12624 ( .A(n10069), .B(n9023), .ZN(n12809) );
  INV_X1 U12625 ( .A(n11417), .ZN(n10071) );
  OAI222_X1 U12626 ( .A1(n12809), .A2(P2_U3088), .B1(n13213), .B2(n10071), 
        .C1(n10070), .C2(n13210), .ZN(P2_U3309) );
  OAI222_X1 U12627 ( .A1(n13833), .A2(n7329), .B1(n13837), .B2(n10071), .C1(
        P1_U3086), .C2(n13479), .ZN(P1_U3337) );
  AOI21_X1 U12628 ( .B1(n10073), .B2(n10072), .A(n12023), .ZN(n10075) );
  NAND2_X1 U12629 ( .A1(n10075), .A2(n10074), .ZN(n10079) );
  INV_X1 U12630 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10470) );
  OAI22_X1 U12631 ( .A1(n12006), .A2(n10469), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10470), .ZN(n10077) );
  INV_X1 U12632 ( .A(n12003), .ZN(n11974) );
  OAI22_X1 U12633 ( .A1(n11974), .A2(n10463), .B1(n10782), .B2(n12000), .ZN(
        n10076) );
  AOI211_X1 U12634 ( .C1(n11977), .C2(n10470), .A(n10077), .B(n10076), .ZN(
        n10078) );
  NAND2_X1 U12635 ( .A1(n10079), .A2(n10078), .ZN(P3_U3158) );
  INV_X1 U12636 ( .A(n10080), .ZN(n10081) );
  OR2_X1 U12637 ( .A1(n10085), .A2(n11607), .ZN(n10087) );
  AOI22_X1 U12638 ( .A1(n11434), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n11433), 
        .B2(n14474), .ZN(n10086) );
  XNOR2_X1 U12639 ( .A(n14617), .B(n11724), .ZN(n10088) );
  NAND2_X1 U12640 ( .A1(n12776), .A2(n9339), .ZN(n10089) );
  NAND2_X1 U12641 ( .A1(n10088), .A2(n10089), .ZN(n10185) );
  INV_X1 U12642 ( .A(n10088), .ZN(n10091) );
  INV_X1 U12643 ( .A(n10089), .ZN(n10090) );
  NAND2_X1 U12644 ( .A1(n10091), .A2(n10090), .ZN(n10092) );
  AND2_X1 U12645 ( .A1(n10185), .A2(n10092), .ZN(n10093) );
  OAI21_X1 U12646 ( .B1(n10094), .B2(n10093), .A(n10186), .ZN(n10095) );
  NAND2_X1 U12647 ( .A1(n10095), .A2(n12763), .ZN(n10108) );
  NAND2_X1 U12648 ( .A1(n11591), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10102) );
  NAND2_X1 U12649 ( .A1(n9864), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n10101) );
  INV_X1 U12650 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10096) );
  AND2_X1 U12651 ( .A1(n10097), .A2(n10096), .ZN(n10098) );
  NOR2_X1 U12652 ( .A1(n10191), .A2(n10098), .ZN(n10190) );
  NAND2_X1 U12653 ( .A1(n11590), .A2(n10190), .ZN(n10100) );
  NAND2_X1 U12654 ( .A1(n11612), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n10099) );
  NAND4_X1 U12655 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n12775) );
  NAND2_X1 U12656 ( .A1(n12775), .A2(n12824), .ZN(n10104) );
  NAND2_X1 U12657 ( .A1(n12777), .A2(n12754), .ZN(n10103) );
  AND2_X1 U12658 ( .A1(n10104), .A2(n10103), .ZN(n10256) );
  NAND2_X1 U12659 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n14475) );
  OAI21_X1 U12660 ( .B1(n12744), .B2(n10256), .A(n14475), .ZN(n10106) );
  INV_X1 U12661 ( .A(n14617), .ZN(n10261) );
  NOR2_X1 U12662 ( .A1(n12761), .A2(n10261), .ZN(n10105) );
  AOI211_X1 U12663 ( .C1(n12758), .C2(n10259), .A(n10106), .B(n10105), .ZN(
        n10107) );
  NAND2_X1 U12664 ( .A1(n10108), .A2(n10107), .ZN(P2_U3193) );
  INV_X1 U12665 ( .A(n10109), .ZN(n10111) );
  OAI222_X1 U12666 ( .A1(n10112), .A2(P3_U3151), .B1(n12664), .B2(n10111), 
        .C1(n10110), .C2(n12661), .ZN(P3_U3275) );
  INV_X1 U12667 ( .A(n11432), .ZN(n10115) );
  OAI222_X1 U12668 ( .A1(n12819), .A2(P2_U3088), .B1(n13213), .B2(n10115), 
        .C1(n10113), .C2(n13210), .ZN(P2_U3308) );
  OAI222_X1 U12669 ( .A1(n13833), .A2(n7326), .B1(n13837), .B2(n10115), .C1(
        P1_U3086), .C2(n10114), .ZN(P1_U3336) );
  INV_X1 U12670 ( .A(n11648), .ZN(n10116) );
  NAND2_X1 U12671 ( .A1(n10119), .A2(n10118), .ZN(n10120) );
  NAND2_X1 U12672 ( .A1(n14588), .A2(n12780), .ZN(n10121) );
  INV_X1 U12673 ( .A(n12780), .ZN(n10137) );
  NAND2_X1 U12674 ( .A1(n10137), .A2(n11325), .ZN(n10147) );
  XNOR2_X1 U12675 ( .A(n10136), .B(n11649), .ZN(n14586) );
  NOR2_X1 U12676 ( .A1(n11638), .A2(n12819), .ZN(n14542) );
  NAND2_X1 U12677 ( .A1(n14554), .A2(n14542), .ZN(n10155) );
  INV_X1 U12678 ( .A(n13076), .ZN(n11017) );
  INV_X1 U12679 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10123) );
  OAI22_X1 U12680 ( .A1(n14554), .A2(n10123), .B1(n10122), .B2(n13071), .ZN(
        n10126) );
  INV_X1 U12681 ( .A(n13078), .ZN(n12953) );
  OAI211_X1 U12682 ( .C1(n10124), .C2(n14588), .A(n10143), .B(n12952), .ZN(
        n14587) );
  NOR2_X1 U12683 ( .A1(n12953), .A2(n14587), .ZN(n10125) );
  AOI211_X1 U12684 ( .C1(n11017), .C2(n11325), .A(n10126), .B(n10125), .ZN(
        n10134) );
  NAND2_X1 U12685 ( .A1(n10128), .A2(n10127), .ZN(n10129) );
  NAND2_X1 U12686 ( .A1(n10129), .A2(n11649), .ZN(n10148) );
  OAI21_X1 U12687 ( .B1(n11649), .B2(n10129), .A(n10148), .ZN(n10131) );
  AOI21_X1 U12688 ( .B1(n10131), .B2(n14548), .A(n10130), .ZN(n10132) );
  OAI21_X1 U12689 ( .B1(n14586), .B2(n9575), .A(n10132), .ZN(n14589) );
  NAND2_X1 U12690 ( .A1(n14589), .A2(n14554), .ZN(n10133) );
  OAI211_X1 U12691 ( .C1(n14586), .C2(n10155), .A(n10134), .B(n10133), .ZN(
        P2_U3261) );
  INV_X1 U12692 ( .A(n11649), .ZN(n10135) );
  NAND2_X1 U12693 ( .A1(n14588), .A2(n10137), .ZN(n10138) );
  INV_X1 U12694 ( .A(n12779), .ZN(n10139) );
  NAND2_X1 U12695 ( .A1(n11331), .A2(n10139), .ZN(n10205) );
  OR2_X1 U12696 ( .A1(n11331), .A2(n10139), .ZN(n10140) );
  XNOR2_X1 U12697 ( .A(n10218), .B(n11650), .ZN(n14593) );
  INV_X1 U12698 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10142) );
  OAI22_X1 U12699 ( .A1(n14554), .A2(n10142), .B1(n10141), .B2(n13071), .ZN(
        n10146) );
  INV_X1 U12700 ( .A(n10143), .ZN(n10144) );
  INV_X1 U12701 ( .A(n11331), .ZN(n14595) );
  OAI211_X1 U12702 ( .C1(n10144), .C2(n14595), .A(n12952), .B(n10213), .ZN(
        n14594) );
  NOR2_X1 U12703 ( .A1(n12953), .A2(n14594), .ZN(n10145) );
  AOI211_X1 U12704 ( .C1(n11017), .C2(n11331), .A(n10146), .B(n10145), .ZN(
        n10154) );
  NAND2_X1 U12705 ( .A1(n10148), .A2(n10147), .ZN(n10149) );
  NAND2_X1 U12706 ( .A1(n10149), .A2(n11650), .ZN(n10206) );
  OAI21_X1 U12707 ( .B1(n11650), .B2(n10149), .A(n10206), .ZN(n10150) );
  NAND2_X1 U12708 ( .A1(n10150), .A2(n14548), .ZN(n10151) );
  OAI211_X1 U12709 ( .C1(n14593), .C2(n9575), .A(n10152), .B(n10151), .ZN(
        n14596) );
  NAND2_X1 U12710 ( .A1(n14596), .A2(n14554), .ZN(n10153) );
  OAI211_X1 U12711 ( .C1(n14593), .C2(n10155), .A(n10154), .B(n10153), .ZN(
        P2_U3260) );
  INV_X2 U12712 ( .A(n14554), .ZN(n14557) );
  OAI22_X1 U12713 ( .A1(n14557), .A2(n10157), .B1(n10156), .B2(n13071), .ZN(
        n10158) );
  AOI21_X1 U12714 ( .B1(P2_REG2_REG_1__SCAN_IN), .B2(n14557), .A(n10158), .ZN(
        n10161) );
  AOI22_X1 U12715 ( .A1(n11017), .A2(n11294), .B1(n13078), .B2(n10159), .ZN(
        n10160) );
  OAI211_X1 U12716 ( .C1(n10162), .C2(n13081), .A(n10161), .B(n10160), .ZN(
        P2_U3264) );
  OAI211_X1 U12717 ( .C1(n6749), .C2(n10046), .A(n12952), .B(n10164), .ZN(
        n14572) );
  INV_X1 U12718 ( .A(n13081), .ZN(n10296) );
  XNOR2_X1 U12719 ( .A(n10166), .B(n10165), .ZN(n14575) );
  AOI22_X1 U12720 ( .A1(n10296), .A2(n14575), .B1(n11017), .B2(n9363), .ZN(
        n10176) );
  OAI21_X1 U12721 ( .B1(n11647), .B2(n10168), .A(n10167), .ZN(n10169) );
  NAND2_X1 U12722 ( .A1(n10169), .A2(n14548), .ZN(n10171) );
  NAND2_X1 U12723 ( .A1(n10171), .A2(n10170), .ZN(n14573) );
  INV_X1 U12724 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n10173) );
  OAI22_X1 U12725 ( .A1(n14554), .A2(n10173), .B1(n10172), .B2(n13071), .ZN(
        n10174) );
  AOI21_X1 U12726 ( .B1(n14554), .B2(n14573), .A(n10174), .ZN(n10175) );
  OAI211_X1 U12727 ( .C1(n12953), .C2(n14572), .A(n10176), .B(n10175), .ZN(
        P2_U3263) );
  OR2_X1 U12728 ( .A1(n10177), .A2(n11607), .ZN(n10179) );
  AOI22_X1 U12729 ( .A1(n11434), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10528), 
        .B2(n11433), .ZN(n10178) );
  XNOR2_X1 U12730 ( .A(n11356), .B(n11724), .ZN(n10180) );
  NAND2_X1 U12731 ( .A1(n12775), .A2(n9339), .ZN(n10181) );
  NAND2_X1 U12732 ( .A1(n10180), .A2(n10181), .ZN(n10266) );
  INV_X1 U12733 ( .A(n10180), .ZN(n10183) );
  INV_X1 U12734 ( .A(n10181), .ZN(n10182) );
  NAND2_X1 U12735 ( .A1(n10183), .A2(n10182), .ZN(n10184) );
  AND2_X1 U12736 ( .A1(n10266), .A2(n10184), .ZN(n10188) );
  OAI21_X1 U12737 ( .B1(n10188), .B2(n10187), .A(n10267), .ZN(n10189) );
  NAND2_X1 U12738 ( .A1(n10189), .A2(n12763), .ZN(n10204) );
  INV_X1 U12739 ( .A(n10190), .ZN(n10246) );
  NAND2_X1 U12740 ( .A1(n9864), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10197) );
  NAND2_X1 U12741 ( .A1(n11591), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U12742 ( .A1(n10191), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10192) );
  OR2_X1 U12743 ( .A1(n10271), .A2(n10192), .ZN(n10325) );
  INV_X1 U12744 ( .A(n10325), .ZN(n10193) );
  NAND2_X1 U12745 ( .A1(n11590), .A2(n10193), .ZN(n10195) );
  NAND2_X1 U12746 ( .A1(n11612), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n10194) );
  NAND4_X1 U12747 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n12774) );
  NAND2_X1 U12748 ( .A1(n12774), .A2(n12824), .ZN(n10199) );
  NAND2_X1 U12749 ( .A1(n12776), .A2(n12754), .ZN(n10198) );
  NAND2_X1 U12750 ( .A1(n10199), .A2(n10198), .ZN(n10242) );
  NAND2_X1 U12751 ( .A1(n12757), .A2(n10242), .ZN(n10201) );
  OAI211_X1 U12752 ( .C1(n12742), .C2(n10246), .A(n10201), .B(n10200), .ZN(
        n10202) );
  AOI21_X1 U12753 ( .B1(n11356), .B2(n12747), .A(n10202), .ZN(n10203) );
  NAND2_X1 U12754 ( .A1(n10204), .A2(n10203), .ZN(P2_U3203) );
  NAND2_X1 U12755 ( .A1(n10206), .A2(n10205), .ZN(n10207) );
  XNOR2_X1 U12756 ( .A(n14601), .B(n12778), .ZN(n11653) );
  OAI21_X1 U12757 ( .B1(n10207), .B2(n11653), .A(n10236), .ZN(n10209) );
  AOI21_X1 U12758 ( .B1(n10209), .B2(n14548), .A(n10208), .ZN(n14603) );
  INV_X1 U12759 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10211) );
  OAI22_X1 U12760 ( .A1(n14554), .A2(n10211), .B1(n10210), .B2(n13071), .ZN(
        n10216) );
  NAND2_X1 U12761 ( .A1(n10213), .A2(n14601), .ZN(n10212) );
  NAND2_X1 U12762 ( .A1(n10212), .A2(n12952), .ZN(n10214) );
  OR2_X1 U12763 ( .A1(n10214), .A2(n10289), .ZN(n14602) );
  NOR2_X1 U12764 ( .A1(n12953), .A2(n14602), .ZN(n10215) );
  AOI211_X1 U12765 ( .C1(n11017), .C2(n14601), .A(n10216), .B(n10215), .ZN(
        n10221) );
  INV_X1 U12766 ( .A(n11650), .ZN(n10217) );
  OR2_X1 U12767 ( .A1(n11331), .A2(n12779), .ZN(n10219) );
  XNOR2_X1 U12768 ( .A(n10226), .B(n11653), .ZN(n14600) );
  INV_X1 U12769 ( .A(n14600), .ZN(n14607) );
  NAND2_X1 U12770 ( .A1(n14607), .A2(n10296), .ZN(n10220) );
  OAI211_X1 U12771 ( .C1(n14603), .C2(n14557), .A(n10221), .B(n10220), .ZN(
        P2_U3259) );
  INV_X1 U12772 ( .A(n10222), .ZN(n10223) );
  OAI222_X1 U12773 ( .A1(P3_U3151), .A2(n12069), .B1(n12661), .B2(n10224), 
        .C1(n12664), .C2(n10223), .ZN(P3_U3274) );
  INV_X1 U12774 ( .A(n10296), .ZN(n10334) );
  INV_X1 U12775 ( .A(n11653), .ZN(n10225) );
  NAND2_X1 U12776 ( .A1(n10226), .A2(n10225), .ZN(n10228) );
  OR2_X1 U12777 ( .A1(n14601), .A2(n12778), .ZN(n10227) );
  NAND2_X1 U12778 ( .A1(n10228), .A2(n10227), .ZN(n10286) );
  INV_X1 U12779 ( .A(n12777), .ZN(n10238) );
  XNOR2_X1 U12780 ( .A(n11347), .B(n10238), .ZN(n11652) );
  NAND2_X1 U12781 ( .A1(n10286), .A2(n11652), .ZN(n10230) );
  OR2_X1 U12782 ( .A1(n11347), .A2(n12777), .ZN(n10229) );
  XNOR2_X1 U12783 ( .A(n14617), .B(n12776), .ZN(n11654) );
  NAND2_X1 U12784 ( .A1(n14617), .A2(n12776), .ZN(n10231) );
  INV_X1 U12785 ( .A(n7463), .ZN(n10232) );
  OR2_X1 U12786 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U12787 ( .A1(n10313), .A2(n10234), .ZN(n14632) );
  NAND2_X1 U12788 ( .A1(n14601), .A2(n11338), .ZN(n10235) );
  OR2_X1 U12789 ( .A1(n11347), .A2(n10238), .ZN(n10237) );
  OR2_X1 U12790 ( .A1(n14617), .A2(n10239), .ZN(n10240) );
  OAI211_X1 U12791 ( .C1(n10241), .C2(n7463), .A(n10318), .B(n14548), .ZN(
        n10244) );
  INV_X1 U12792 ( .A(n10242), .ZN(n10243) );
  AND2_X1 U12793 ( .A1(n10244), .A2(n10243), .ZN(n14635) );
  MUX2_X1 U12794 ( .A(n9992), .B(n14635), .S(n14554), .Z(n10249) );
  AOI21_X1 U12795 ( .B1(n10258), .B2(n11356), .A(n9339), .ZN(n10245) );
  AND2_X1 U12796 ( .A1(n10245), .A2(n10327), .ZN(n14625) );
  INV_X1 U12797 ( .A(n11356), .ZN(n14628) );
  OAI22_X1 U12798 ( .A1(n13076), .A2(n14628), .B1(n10246), .B2(n13071), .ZN(
        n10247) );
  AOI21_X1 U12799 ( .B1(n14625), .B2(n13078), .A(n10247), .ZN(n10248) );
  OAI211_X1 U12800 ( .C1(n10334), .C2(n14632), .A(n10249), .B(n10248), .ZN(
        P2_U3256) );
  NAND2_X1 U12801 ( .A1(n10250), .A2(n11654), .ZN(n10251) );
  NAND2_X1 U12802 ( .A1(n10252), .A2(n10251), .ZN(n14620) );
  NAND2_X1 U12803 ( .A1(n10253), .A2(n6743), .ZN(n10254) );
  NAND3_X1 U12804 ( .A1(n10255), .A2(n14548), .A3(n10254), .ZN(n10257) );
  NAND2_X1 U12805 ( .A1(n10257), .A2(n10256), .ZN(n14623) );
  NAND2_X1 U12806 ( .A1(n14623), .A2(n14554), .ZN(n10265) );
  OAI211_X1 U12807 ( .C1(n10287), .C2(n10261), .A(n12952), .B(n10258), .ZN(
        n14618) );
  INV_X1 U12808 ( .A(n14618), .ZN(n10263) );
  AOI22_X1 U12809 ( .A1(n14557), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10259), 
        .B2(n14553), .ZN(n10260) );
  OAI21_X1 U12810 ( .B1(n10261), .B2(n13076), .A(n10260), .ZN(n10262) );
  AOI21_X1 U12811 ( .B1(n10263), .B2(n13078), .A(n10262), .ZN(n10264) );
  OAI211_X1 U12812 ( .C1(n10334), .C2(n14620), .A(n10265), .B(n10264), .ZN(
        P2_U3257) );
  NAND2_X1 U12813 ( .A1(n10268), .A2(n11584), .ZN(n10270) );
  AOI22_X1 U12814 ( .A1(n14486), .A2(n11433), .B1(n11434), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n10269) );
  NAND2_X2 U12815 ( .A1(n10270), .A2(n10269), .ZN(n14638) );
  XNOR2_X1 U12816 ( .A(n14638), .B(n11724), .ZN(n10480) );
  NAND2_X1 U12817 ( .A1(n12774), .A2(n9339), .ZN(n10481) );
  XNOR2_X1 U12818 ( .A(n10480), .B(n10481), .ZN(n10479) );
  XNOR2_X1 U12819 ( .A(n10478), .B(n10479), .ZN(n10282) );
  NAND2_X1 U12820 ( .A1(n11591), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10276) );
  NAND2_X1 U12821 ( .A1(n9864), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10275) );
  OR2_X1 U12822 ( .A1(n10271), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10272) );
  AND2_X1 U12823 ( .A1(n10425), .A2(n10272), .ZN(n10434) );
  NAND2_X1 U12824 ( .A1(n11590), .A2(n10434), .ZN(n10274) );
  NAND2_X1 U12825 ( .A1(n11612), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10273) );
  NAND4_X1 U12826 ( .A1(n10276), .A2(n10275), .A3(n10274), .A4(n10273), .ZN(
        n12773) );
  NAND2_X1 U12827 ( .A1(n12773), .A2(n12824), .ZN(n10278) );
  NAND2_X1 U12828 ( .A1(n12775), .A2(n12754), .ZN(n10277) );
  NAND2_X1 U12829 ( .A1(n10278), .A2(n10277), .ZN(n10322) );
  NAND2_X1 U12830 ( .A1(n12757), .A2(n10322), .ZN(n10279) );
  NAND2_X1 U12831 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n14487)
         );
  OAI211_X1 U12832 ( .C1(n12742), .C2(n10325), .A(n10279), .B(n14487), .ZN(
        n10280) );
  AOI21_X1 U12833 ( .B1(n14638), .B2(n12747), .A(n10280), .ZN(n10281) );
  OAI21_X1 U12834 ( .B1(n10282), .B2(n12749), .A(n10281), .ZN(P2_U3189) );
  XOR2_X1 U12835 ( .A(n11652), .B(n10283), .Z(n10285) );
  AOI21_X1 U12836 ( .B1(n10285), .B2(n14548), .A(n10284), .ZN(n14611) );
  XNOR2_X1 U12837 ( .A(n10286), .B(n11652), .ZN(n14615) );
  INV_X1 U12838 ( .A(n10287), .ZN(n10288) );
  OAI211_X1 U12839 ( .C1(n14610), .C2(n10289), .A(n10288), .B(n12952), .ZN(
        n14609) );
  INV_X1 U12840 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10292) );
  INV_X1 U12841 ( .A(n10290), .ZN(n10291) );
  OAI22_X1 U12842 ( .A1(n14554), .A2(n10292), .B1(n10291), .B2(n13071), .ZN(
        n10293) );
  AOI21_X1 U12843 ( .B1(n11017), .B2(n11347), .A(n10293), .ZN(n10294) );
  OAI21_X1 U12844 ( .B1(n14609), .B2(n12953), .A(n10294), .ZN(n10295) );
  AOI21_X1 U12845 ( .B1(n14615), .B2(n10296), .A(n10295), .ZN(n10297) );
  OAI21_X1 U12846 ( .B1(n14611), .B2(n14557), .A(n10297), .ZN(P2_U3258) );
  OAI22_X1 U12847 ( .A1(n11815), .A2(n10370), .B1(n14367), .B2(n11823), .ZN(
        n10302) );
  OAI22_X1 U12848 ( .A1(n14367), .A2(n11824), .B1(n11823), .B2(n10370), .ZN(
        n10300) );
  XOR2_X1 U12849 ( .A(n11856), .B(n10300), .Z(n10341) );
  NOR2_X1 U12850 ( .A1(n10340), .A2(n10341), .ZN(n10339) );
  AOI22_X1 U12851 ( .A1(n9889), .A2(n14376), .B1(n6452), .B2(n13350), .ZN(
        n10304) );
  XNOR2_X1 U12852 ( .A(n10304), .B(n11856), .ZN(n10550) );
  AOI22_X1 U12853 ( .A1(n11858), .A2(n13350), .B1(n6452), .B2(n14376), .ZN(
        n10553) );
  XNOR2_X1 U12854 ( .A(n10550), .B(n10553), .ZN(n10305) );
  XNOR2_X1 U12855 ( .A(n10552), .B(n10305), .ZN(n10311) );
  INV_X1 U12856 ( .A(n14083), .ZN(n13326) );
  OR2_X1 U12857 ( .A1(n10370), .A2(n13963), .ZN(n10307) );
  NAND2_X1 U12858 ( .A1(n13349), .A2(n6454), .ZN(n10306) );
  NAND2_X1 U12859 ( .A1(n10307), .A2(n10306), .ZN(n14375) );
  AOI22_X1 U12860 ( .A1(n10337), .A2(n14375), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10308) );
  OAI21_X1 U12861 ( .B1(n13329), .B2(n7025), .A(n10308), .ZN(n10309) );
  AOI21_X1 U12862 ( .B1(n10498), .B2(n13326), .A(n10309), .ZN(n10310) );
  OAI21_X1 U12863 ( .B1(n10311), .B2(n14078), .A(n10310), .ZN(P1_U3227) );
  NAND2_X1 U12864 ( .A1(n11356), .A2(n12775), .ZN(n10312) );
  NAND2_X1 U12865 ( .A1(n10313), .A2(n10312), .ZN(n10315) );
  INV_X1 U12866 ( .A(n12774), .ZN(n10314) );
  NAND2_X1 U12867 ( .A1(n10315), .A2(n11657), .ZN(n10439) );
  OR2_X1 U12868 ( .A1(n10315), .A2(n11657), .ZN(n10316) );
  NAND2_X1 U12869 ( .A1(n10439), .A2(n10316), .ZN(n14642) );
  INV_X1 U12870 ( .A(n12775), .ZN(n11358) );
  OR2_X1 U12871 ( .A1(n11356), .A2(n11358), .ZN(n10317) );
  INV_X1 U12872 ( .A(n11657), .ZN(n10319) );
  NOR2_X1 U12873 ( .A1(n10320), .A2(n10319), .ZN(n10321) );
  INV_X1 U12874 ( .A(n14548), .ZN(n12946) );
  OR3_X1 U12875 ( .A1(n10418), .A2(n10321), .A3(n12946), .ZN(n10324) );
  INV_X1 U12876 ( .A(n10322), .ZN(n10323) );
  NAND2_X1 U12877 ( .A1(n10324), .A2(n10323), .ZN(n14645) );
  NAND2_X1 U12878 ( .A1(n14645), .A2(n14554), .ZN(n10333) );
  INV_X1 U12879 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10326) );
  OAI22_X1 U12880 ( .A1(n14554), .A2(n10326), .B1(n10325), .B2(n13071), .ZN(
        n10331) );
  NAND2_X1 U12881 ( .A1(n14638), .A2(n10327), .ZN(n10328) );
  NAND2_X1 U12882 ( .A1(n10328), .A2(n12952), .ZN(n10329) );
  OR2_X1 U12883 ( .A1(n10435), .A2(n10329), .ZN(n14639) );
  NOR2_X1 U12884 ( .A1(n14639), .A2(n12953), .ZN(n10330) );
  AOI211_X1 U12885 ( .C1(n11017), .C2(n14638), .A(n10331), .B(n10330), .ZN(
        n10332) );
  OAI211_X1 U12886 ( .C1(n10334), .C2(n14642), .A(n10333), .B(n10332), .ZN(
        P2_U3255) );
  NAND2_X1 U12887 ( .A1(n13352), .A2(n14087), .ZN(n10336) );
  NAND2_X1 U12888 ( .A1(n13350), .A2(n6454), .ZN(n10335) );
  NAND2_X1 U12889 ( .A1(n10336), .A2(n10335), .ZN(n10653) );
  NAND2_X1 U12890 ( .A1(n10337), .A2(n10653), .ZN(n10338) );
  NAND2_X1 U12891 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n13398) );
  OAI211_X1 U12892 ( .C1(n13329), .C2(n14367), .A(n10338), .B(n13398), .ZN(
        n10343) );
  AOI211_X1 U12893 ( .C1(n10341), .C2(n10340), .A(n14078), .B(n10339), .ZN(
        n10342) );
  AOI211_X1 U12894 ( .C1(n10654), .C2(n13326), .A(n10343), .B(n10342), .ZN(
        n10344) );
  INV_X1 U12895 ( .A(n10344), .ZN(P1_U3230) );
  NOR2_X1 U12896 ( .A1(n12661), .A2(SI_22_), .ZN(n10345) );
  AOI21_X1 U12897 ( .B1(n12068), .B2(P3_STATE_REG_SCAN_IN), .A(n10345), .ZN(
        n10346) );
  OAI21_X1 U12898 ( .B1(n10347), .B2(n12664), .A(n10346), .ZN(n10348) );
  INV_X1 U12899 ( .A(n10348), .ZN(P3_U3273) );
  OAI21_X1 U12900 ( .B1(n10351), .B2(n10350), .A(n10349), .ZN(n10352) );
  NAND2_X1 U12901 ( .A1(n10352), .A2(n14668), .ZN(n10356) );
  OAI22_X1 U12902 ( .A1(n11974), .A2(n14761), .B1(n10728), .B2(n12000), .ZN(
        n10353) );
  AOI211_X1 U12903 ( .C1(n10663), .C2(n14675), .A(n10354), .B(n10353), .ZN(
        n10355) );
  OAI211_X1 U12904 ( .C1(n10664), .C2(n14678), .A(n10356), .B(n10355), .ZN(
        P3_U3170) );
  INV_X1 U12905 ( .A(n10357), .ZN(n10360) );
  NAND4_X1 U12906 ( .A1(n10361), .A2(n10360), .A3(n10359), .A4(n10358), .ZN(
        n13546) );
  INV_X1 U12907 ( .A(n10362), .ZN(n10363) );
  INV_X2 U12908 ( .A(n13970), .ZN(n14322) );
  OR2_X1 U12909 ( .A1(n14322), .A2(n10571), .ZN(n10366) );
  NAND2_X1 U12910 ( .A1(n10367), .A2(n10572), .ZN(n10368) );
  INV_X1 U12911 ( .A(n10496), .ZN(n10371) );
  OR2_X1 U12912 ( .A1(n14376), .A2(n13350), .ZN(n10372) );
  NAND2_X1 U12913 ( .A1(n10373), .A2(n10372), .ZN(n14290) );
  OR2_X1 U12914 ( .A1(n10559), .A2(n13349), .ZN(n10374) );
  XNOR2_X1 U12915 ( .A(n10398), .B(n10387), .ZN(n14399) );
  NAND2_X1 U12916 ( .A1(n10376), .A2(n10375), .ZN(n10378) );
  NOR2_X1 U12917 ( .A1(n13351), .A2(n14367), .ZN(n10379) );
  NAND2_X1 U12918 ( .A1(n13351), .A2(n14367), .ZN(n10380) );
  INV_X1 U12919 ( .A(n13350), .ZN(n10381) );
  NOR2_X1 U12920 ( .A1(n14376), .A2(n10381), .ZN(n10383) );
  NAND2_X1 U12921 ( .A1(n14376), .A2(n10381), .ZN(n10382) );
  NAND2_X1 U12922 ( .A1(n14292), .A2(n10384), .ZN(n10386) );
  NAND2_X1 U12923 ( .A1(n10559), .A2(n10561), .ZN(n10385) );
  INV_X1 U12924 ( .A(n10387), .ZN(n10397) );
  XNOR2_X1 U12925 ( .A(n10404), .B(n10397), .ZN(n10388) );
  AOI22_X1 U12926 ( .A1(n14087), .A2(n13349), .B1(n13347), .B2(n6454), .ZN(
        n10696) );
  OAI21_X1 U12927 ( .B1(n10388), .B2(n14379), .A(n10696), .ZN(n14394) );
  INV_X1 U12928 ( .A(n14396), .ZN(n10394) );
  NAND2_X1 U12929 ( .A1(n10390), .A2(n10389), .ZN(n14094) );
  INV_X1 U12930 ( .A(n10391), .ZN(n14301) );
  AOI211_X1 U12931 ( .C1(n14396), .C2(n14301), .A(n14352), .B(n6434), .ZN(
        n14395) );
  NOR2_X2 U12932 ( .A1(n13546), .A2(n13486), .ZN(n14313) );
  NAND2_X1 U12933 ( .A1(n14395), .A2(n14313), .ZN(n10393) );
  INV_X1 U12934 ( .A(n14093), .ZN(n14311) );
  AOI22_X1 U12935 ( .A1(n14315), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n10698), 
        .B2(n14311), .ZN(n10392) );
  OAI211_X1 U12936 ( .C1(n10394), .C2(n14298), .A(n10393), .B(n10392), .ZN(
        n10395) );
  AOI21_X1 U12937 ( .B1(n13970), .B2(n14394), .A(n10395), .ZN(n10396) );
  OAI21_X1 U12938 ( .B1(n13675), .B2(n14399), .A(n10396), .ZN(P1_U3286) );
  OR2_X1 U12939 ( .A1(n14396), .A2(n13348), .ZN(n10399) );
  OR2_X1 U12940 ( .A1(n10858), .A2(n13347), .ZN(n10400) );
  INV_X1 U12941 ( .A(n10536), .ZN(n10539) );
  NAND2_X1 U12942 ( .A1(n10540), .A2(n10539), .ZN(n10402) );
  NAND2_X1 U12943 ( .A1(n14412), .A2(n10974), .ZN(n10401) );
  NAND2_X1 U12944 ( .A1(n10402), .A2(n10401), .ZN(n10512) );
  XNOR2_X1 U12945 ( .A(n10512), .B(n10511), .ZN(n14422) );
  INV_X1 U12946 ( .A(n14422), .ZN(n10417) );
  INV_X1 U12947 ( .A(n13348), .ZN(n10692) );
  AND2_X1 U12948 ( .A1(n14396), .A2(n10692), .ZN(n10403) );
  OR2_X1 U12949 ( .A1(n14396), .A2(n10692), .ZN(n10405) );
  INV_X1 U12950 ( .A(n13347), .ZN(n10904) );
  NOR2_X1 U12951 ( .A1(n10858), .A2(n10904), .ZN(n10406) );
  NAND2_X1 U12952 ( .A1(n10537), .A2(n10536), .ZN(n10409) );
  OR2_X1 U12953 ( .A1(n14412), .A2(n13346), .ZN(n10408) );
  OAI211_X1 U12954 ( .C1(n6618), .C2(n10410), .A(n14373), .B(n10509), .ZN(
        n10411) );
  OAI21_X1 U12955 ( .B1(n10974), .B2(n13963), .A(n10411), .ZN(n14419) );
  INV_X1 U12956 ( .A(n14315), .ZN(n13970) );
  INV_X1 U12957 ( .A(n10976), .ZN(n14418) );
  INV_X1 U12958 ( .A(n10514), .ZN(n10412) );
  OAI211_X1 U12959 ( .C1(n14418), .C2(n10542), .A(n10412), .B(n9843), .ZN(
        n14416) );
  NAND2_X1 U12960 ( .A1(n13344), .A2(n6454), .ZN(n14415) );
  AOI21_X1 U12961 ( .B1(n14416), .B2(n14415), .A(n13720), .ZN(n10415) );
  AOI22_X1 U12962 ( .A1(n14322), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n10971), 
        .B2(n14311), .ZN(n10413) );
  OAI21_X1 U12963 ( .B1(n14418), .B2(n14298), .A(n10413), .ZN(n10414) );
  AOI211_X1 U12964 ( .C1(n14419), .C2(n13970), .A(n10415), .B(n10414), .ZN(
        n10416) );
  OAI21_X1 U12965 ( .B1(n13675), .B2(n10417), .A(n10416), .ZN(P1_U3283) );
  INV_X1 U12966 ( .A(n14638), .ZN(n10419) );
  NAND2_X1 U12967 ( .A1(n10420), .A2(n11584), .ZN(n10422) );
  AOI22_X1 U12968 ( .A1(n10706), .A2(n11433), .B1(n11434), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n10421) );
  INV_X1 U12969 ( .A(n12773), .ZN(n11376) );
  XNOR2_X1 U12970 ( .A(n11374), .B(n11376), .ZN(n11658) );
  INV_X1 U12971 ( .A(n11658), .ZN(n10440) );
  OAI21_X1 U12972 ( .B1(n10423), .B2(n10440), .A(n10735), .ZN(n10433) );
  NAND2_X1 U12973 ( .A1(n9864), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10430) );
  NAND2_X1 U12974 ( .A1(n10425), .A2(n10424), .ZN(n10426) );
  AND2_X1 U12975 ( .A1(n10598), .A2(n10426), .ZN(n10742) );
  NAND2_X1 U12976 ( .A1(n11590), .A2(n10742), .ZN(n10429) );
  NAND2_X1 U12977 ( .A1(n11591), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U12978 ( .A1(n11612), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10427) );
  NAND4_X1 U12979 ( .A1(n10430), .A2(n10429), .A3(n10428), .A4(n10427), .ZN(
        n12772) );
  NAND2_X1 U12980 ( .A1(n12772), .A2(n12824), .ZN(n10432) );
  NAND2_X1 U12981 ( .A1(n12774), .A2(n12754), .ZN(n10431) );
  NAND2_X1 U12982 ( .A1(n10432), .A2(n10431), .ZN(n10487) );
  AOI21_X1 U12983 ( .B1(n10433), .B2(n14548), .A(n10487), .ZN(n10717) );
  INV_X1 U12984 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10520) );
  INV_X1 U12985 ( .A(n10434), .ZN(n10489) );
  OAI22_X1 U12986 ( .A1(n14554), .A2(n10520), .B1(n10489), .B2(n13071), .ZN(
        n10437) );
  NAND2_X1 U12987 ( .A1(n10736), .A2(n10435), .ZN(n10741) );
  OAI211_X1 U12988 ( .C1(n10736), .C2(n10435), .A(n10741), .B(n12952), .ZN(
        n10716) );
  NOR2_X1 U12989 ( .A1(n10716), .A2(n12953), .ZN(n10436) );
  AOI211_X1 U12990 ( .C1(n11017), .C2(n11374), .A(n10437), .B(n10436), .ZN(
        n10442) );
  NAND2_X1 U12991 ( .A1(n14638), .A2(n12774), .ZN(n10438) );
  NAND2_X1 U12992 ( .A1(n10439), .A2(n10438), .ZN(n10745) );
  XNOR2_X1 U12993 ( .A(n10745), .B(n10440), .ZN(n10719) );
  NAND2_X1 U12994 ( .A1(n10719), .A2(n10296), .ZN(n10441) );
  OAI211_X1 U12995 ( .C1(n10717), .C2(n14557), .A(n10442), .B(n10441), .ZN(
        P2_U3254) );
  XNOR2_X1 U12996 ( .A(n10443), .B(n10448), .ZN(n10446) );
  OR2_X1 U12997 ( .A1(n10974), .A2(n13965), .ZN(n10445) );
  NAND2_X1 U12998 ( .A1(n13348), .A2(n14087), .ZN(n10444) );
  NAND2_X1 U12999 ( .A1(n10445), .A2(n10444), .ZN(n10854) );
  AOI21_X1 U13000 ( .B1(n10446), .B2(n14373), .A(n10854), .ZN(n14406) );
  XNOR2_X1 U13001 ( .A(n10447), .B(n10448), .ZN(n14408) );
  NAND2_X1 U13002 ( .A1(n14408), .A2(n14308), .ZN(n10453) );
  OAI22_X1 U13003 ( .A1(n13970), .A2(n10449), .B1(n10861), .B2(n14093), .ZN(
        n10451) );
  OAI211_X1 U13004 ( .C1(n6434), .C2(n6822), .A(n9843), .B(n10541), .ZN(n14405) );
  NOR2_X1 U13005 ( .A1(n14405), .A2(n13720), .ZN(n10450) );
  AOI211_X1 U13006 ( .C1(n14310), .C2(n10858), .A(n10451), .B(n10450), .ZN(
        n10452) );
  OAI211_X1 U13007 ( .C1(n14322), .C2(n14406), .A(n10453), .B(n10452), .ZN(
        P1_U3285) );
  XNOR2_X1 U13008 ( .A(n10455), .B(n10454), .ZN(n10456) );
  NAND2_X1 U13009 ( .A1(n10456), .A2(n14668), .ZN(n10460) );
  OAI22_X1 U13010 ( .A1(n11974), .A2(n10782), .B1(n10781), .B2(n12000), .ZN(
        n10457) );
  AOI211_X1 U13011 ( .C1(n10775), .C2(n14675), .A(n10458), .B(n10457), .ZN(
        n10459) );
  OAI211_X1 U13012 ( .C1(n10776), .C2(n14678), .A(n10460), .B(n10459), .ZN(
        P3_U3167) );
  OAI21_X1 U13013 ( .B1(n10462), .B2(n12221), .A(n10461), .ZN(n14808) );
  INV_X1 U13014 ( .A(n14808), .ZN(n10473) );
  OAI22_X1 U13015 ( .A1(n10463), .A2(n14762), .B1(n10782), .B2(n14760), .ZN(
        n10468) );
  INV_X1 U13016 ( .A(n10464), .ZN(n10465) );
  AOI211_X1 U13017 ( .C1(n12221), .C2(n10466), .A(n12418), .B(n10465), .ZN(
        n10467) );
  AOI211_X1 U13018 ( .C1(n14843), .C2(n14808), .A(n10468), .B(n10467), .ZN(
        n14805) );
  MUX2_X1 U13019 ( .A(n14904), .B(n14805), .S(n14791), .Z(n10472) );
  INV_X1 U13020 ( .A(n10873), .ZN(n14726) );
  NOR2_X1 U13021 ( .A1(n10469), .A2(n14837), .ZN(n14807) );
  AOI22_X1 U13022 ( .A1(n14726), .A2(n14807), .B1(n14772), .B2(n10470), .ZN(
        n10471) );
  OAI211_X1 U13023 ( .C1(n10473), .C2(n14787), .A(n10472), .B(n10471), .ZN(
        P3_U3230) );
  XNOR2_X1 U13024 ( .A(n11374), .B(n11724), .ZN(n10477) );
  INV_X1 U13025 ( .A(n10477), .ZN(n10475) );
  NAND2_X1 U13026 ( .A1(n12773), .A2(n9339), .ZN(n10476) );
  INV_X1 U13027 ( .A(n10476), .ZN(n10474) );
  NAND2_X1 U13028 ( .A1(n10475), .A2(n10474), .ZN(n10588) );
  NAND2_X1 U13029 ( .A1(n10477), .A2(n10476), .ZN(n10586) );
  NAND2_X1 U13030 ( .A1(n10588), .A2(n10586), .ZN(n10486) );
  INV_X1 U13031 ( .A(n10480), .ZN(n10483) );
  INV_X1 U13032 ( .A(n10481), .ZN(n10482) );
  NAND2_X1 U13033 ( .A1(n10483), .A2(n10482), .ZN(n10484) );
  NAND2_X1 U13034 ( .A1(n10485), .A2(n10484), .ZN(n10587) );
  XOR2_X1 U13035 ( .A(n10486), .B(n10587), .Z(n10492) );
  NAND2_X1 U13036 ( .A1(n12757), .A2(n10487), .ZN(n10488) );
  NAND2_X1 U13037 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n10525)
         );
  OAI211_X1 U13038 ( .C1(n12742), .C2(n10489), .A(n10488), .B(n10525), .ZN(
        n10490) );
  AOI21_X1 U13039 ( .B1(n11374), .B2(n12747), .A(n10490), .ZN(n10491) );
  OAI21_X1 U13040 ( .B1(n10492), .B2(n12749), .A(n10491), .ZN(P2_U3208) );
  INV_X1 U13041 ( .A(n11448), .ZN(n10519) );
  OAI222_X1 U13042 ( .A1(n13837), .A2(n10519), .B1(n10494), .B2(P1_U3086), 
        .C1(n10493), .C2(n13833), .ZN(P1_U3335) );
  XNOR2_X1 U13043 ( .A(n10495), .B(n10496), .ZN(n14381) );
  INV_X1 U13044 ( .A(n14381), .ZN(n14384) );
  XNOR2_X1 U13045 ( .A(n10497), .B(n10496), .ZN(n14380) );
  INV_X1 U13046 ( .A(n14375), .ZN(n10500) );
  INV_X1 U13047 ( .A(n10498), .ZN(n10499) );
  OAI22_X1 U13048 ( .A1(n14322), .A2(n10500), .B1(n10499), .B2(n14093), .ZN(
        n10501) );
  AOI21_X1 U13049 ( .B1(n14310), .B2(n14376), .A(n10501), .ZN(n10505) );
  AOI21_X1 U13050 ( .B1(n10650), .B2(n14376), .A(n14352), .ZN(n10502) );
  NAND2_X1 U13051 ( .A1(n10502), .A2(n14300), .ZN(n14377) );
  INV_X1 U13052 ( .A(n14377), .ZN(n10503) );
  AOI22_X1 U13053 ( .A1(n14313), .A2(n10503), .B1(n14315), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n10504) );
  OAI211_X1 U13054 ( .C1(n13705), .C2(n14380), .A(n10505), .B(n10504), .ZN(
        n10506) );
  AOI21_X1 U13055 ( .B1(n14384), .B2(n14308), .A(n10506), .ZN(n10507) );
  INV_X1 U13056 ( .A(n10507), .ZN(P1_U3288) );
  INV_X1 U13057 ( .A(n13345), .ZN(n10968) );
  OR2_X1 U13058 ( .A1(n10976), .A2(n10968), .ZN(n10508) );
  XNOR2_X1 U13059 ( .A(n10791), .B(n10794), .ZN(n10510) );
  AOI222_X1 U13060 ( .A1(n13345), .A2(n14087), .B1(n13343), .B2(n6454), .C1(
        n14373), .C2(n10510), .ZN(n14151) );
  OR2_X1 U13061 ( .A1(n10976), .A2(n13345), .ZN(n10513) );
  XNOR2_X1 U13062 ( .A(n10795), .B(n10794), .ZN(n14154) );
  INV_X1 U13063 ( .A(n11100), .ZN(n14152) );
  OAI211_X1 U13064 ( .C1(n10514), .C2(n14152), .A(n9843), .B(n10799), .ZN(
        n14150) );
  AOI22_X1 U13065 ( .A1(n14315), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11115), 
        .B2(n14311), .ZN(n10516) );
  NAND2_X1 U13066 ( .A1(n11100), .A2(n14310), .ZN(n10515) );
  OAI211_X1 U13067 ( .C1(n14150), .C2(n13720), .A(n10516), .B(n10515), .ZN(
        n10517) );
  AOI21_X1 U13068 ( .B1(n14154), .B2(n14308), .A(n10517), .ZN(n10518) );
  OAI21_X1 U13069 ( .B1(n14151), .B2(n14322), .A(n10518), .ZN(P1_U3282) );
  OAI222_X1 U13070 ( .A1(n11671), .A2(P2_U3088), .B1(n13210), .B2(n11449), 
        .C1(n10519), .C2(n13213), .ZN(P2_U3307) );
  XNOR2_X1 U13071 ( .A(n10706), .B(n10520), .ZN(n10523) );
  OAI21_X1 U13072 ( .B1(P2_REG2_REG_9__SCAN_IN), .B2(n10528), .A(n10521), .ZN(
        n14479) );
  XNOR2_X1 U13073 ( .A(n14486), .B(P2_REG2_REG_10__SCAN_IN), .ZN(n14480) );
  NOR2_X1 U13074 ( .A1(n14479), .A2(n14480), .ZN(n14478) );
  OAI21_X1 U13075 ( .B1(n10523), .B2(n10522), .A(n10701), .ZN(n10524) );
  INV_X1 U13076 ( .A(n10524), .ZN(n10535) );
  OAI21_X1 U13077 ( .B1(n12815), .B2(n10526), .A(n10525), .ZN(n10533) );
  OAI21_X1 U13078 ( .B1(P2_REG1_REG_9__SCAN_IN), .B2(n10528), .A(n10527), .ZN(
        n14482) );
  INV_X1 U13079 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10529) );
  MUX2_X1 U13080 ( .A(n10529), .B(P2_REG1_REG_10__SCAN_IN), .S(n14486), .Z(
        n14483) );
  XNOR2_X1 U13081 ( .A(n10706), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n10530) );
  AOI211_X1 U13082 ( .C1(n10531), .C2(n10530), .A(n14531), .B(n10705), .ZN(
        n10532) );
  AOI211_X1 U13083 ( .C1(n14442), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n10533), 
        .B(n10532), .ZN(n10534) );
  OAI21_X1 U13084 ( .B1(n10535), .B2(n14527), .A(n10534), .ZN(P2_U3225) );
  XNOR2_X1 U13085 ( .A(n10537), .B(n10536), .ZN(n10538) );
  AOI222_X1 U13086 ( .A1(n13347), .A2(n14087), .B1(n13345), .B2(n6454), .C1(
        n14373), .C2(n10538), .ZN(n14411) );
  MUX2_X1 U13087 ( .A(n9470), .B(n14411), .S(n13970), .Z(n10549) );
  XNOR2_X1 U13088 ( .A(n10540), .B(n10539), .ZN(n14414) );
  INV_X1 U13089 ( .A(n10541), .ZN(n10544) );
  INV_X1 U13090 ( .A(n10542), .ZN(n10543) );
  OAI211_X1 U13091 ( .C1(n14412), .C2(n10544), .A(n10543), .B(n9843), .ZN(
        n14410) );
  AOI22_X1 U13092 ( .A1(n14310), .A2(n10545), .B1(n14311), .B2(n10906), .ZN(
        n10546) );
  OAI21_X1 U13093 ( .B1(n14410), .B2(n13720), .A(n10546), .ZN(n10547) );
  AOI21_X1 U13094 ( .B1(n14414), .B2(n14308), .A(n10547), .ZN(n10548) );
  NAND2_X1 U13095 ( .A1(n10549), .A2(n10548), .ZN(P1_U3284) );
  AOI21_X1 U13096 ( .B1(n10552), .B2(n10553), .A(n10550), .ZN(n10551) );
  INV_X1 U13097 ( .A(n10552), .ZN(n10555) );
  INV_X1 U13098 ( .A(n10553), .ZN(n10554) );
  NAND2_X1 U13099 ( .A1(n10559), .A2(n9889), .ZN(n10557) );
  NAND2_X1 U13100 ( .A1(n6452), .A2(n13349), .ZN(n10556) );
  NAND2_X1 U13101 ( .A1(n10557), .A2(n10556), .ZN(n10558) );
  XNOR2_X1 U13102 ( .A(n10558), .B(n11856), .ZN(n10690) );
  NAND2_X1 U13103 ( .A1(n10559), .A2(n6452), .ZN(n10560) );
  OAI21_X1 U13104 ( .B1(n10561), .B2(n11815), .A(n10560), .ZN(n10689) );
  XNOR2_X1 U13105 ( .A(n10690), .B(n10689), .ZN(n10691) );
  XNOR2_X1 U13106 ( .A(n6596), .B(n10691), .ZN(n10566) );
  AOI22_X1 U13107 ( .A1(n14087), .A2(n13350), .B1(n13348), .B2(n6454), .ZN(
        n14293) );
  INV_X1 U13108 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10562) );
  OAI22_X1 U13109 ( .A1(n13334), .A2(n14293), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10562), .ZN(n10564) );
  NOR2_X1 U13110 ( .A1(n13329), .A2(n14387), .ZN(n10563) );
  AOI211_X1 U13111 ( .C1(n14296), .C2(n13326), .A(n10564), .B(n10563), .ZN(
        n10565) );
  OAI21_X1 U13112 ( .B1(n10566), .B2(n14078), .A(n10565), .ZN(P1_U3239) );
  XNOR2_X1 U13113 ( .A(n10567), .B(n10569), .ZN(n10575) );
  OAI21_X1 U13114 ( .B1(n10570), .B2(n10569), .A(n10568), .ZN(n14362) );
  INV_X1 U13115 ( .A(n10571), .ZN(n14403) );
  AOI21_X1 U13116 ( .B1(n14362), .B2(n14403), .A(n10573), .ZN(n10574) );
  OAI21_X1 U13117 ( .B1(n14379), .B2(n10575), .A(n10574), .ZN(n14360) );
  INV_X1 U13118 ( .A(n10576), .ZN(n14304) );
  AOI22_X1 U13119 ( .A1(n14304), .A2(n14362), .B1(n14310), .B2(n10577), .ZN(
        n10582) );
  NAND2_X1 U13120 ( .A1(n10610), .A2(n10577), .ZN(n10578) );
  NAND2_X1 U13121 ( .A1(n10578), .A2(n9843), .ZN(n10579) );
  NOR2_X1 U13122 ( .A1(n10580), .A2(n10579), .ZN(n14358) );
  AOI22_X1 U13123 ( .A1(n14313), .A2(n14358), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14311), .ZN(n10581) );
  OAI211_X1 U13124 ( .C1(n10583), .C2(n13970), .A(n10582), .B(n10581), .ZN(
        n10584) );
  AOI21_X1 U13125 ( .B1(n13970), .B2(n14360), .A(n10584), .ZN(n10585) );
  INV_X1 U13126 ( .A(n10585), .ZN(P1_U3291) );
  NAND2_X1 U13127 ( .A1(n10587), .A2(n10586), .ZN(n10589) );
  NAND2_X1 U13128 ( .A1(n10589), .A2(n10588), .ZN(n10754) );
  NAND2_X1 U13129 ( .A1(n10590), .A2(n11584), .ZN(n10592) );
  AOI22_X1 U13130 ( .A1(n10882), .A2(n11433), .B1(n11434), .B2(
        P1_DATAO_REG_12__SCAN_IN), .ZN(n10591) );
  XNOR2_X1 U13131 ( .A(n13172), .B(n11729), .ZN(n10596) );
  INV_X1 U13132 ( .A(n10596), .ZN(n10594) );
  AND2_X1 U13133 ( .A1(n12772), .A2(n9339), .ZN(n10595) );
  INV_X1 U13134 ( .A(n10595), .ZN(n10593) );
  NAND2_X1 U13135 ( .A1(n10594), .A2(n10593), .ZN(n10756) );
  AND2_X1 U13136 ( .A1(n10596), .A2(n10595), .ZN(n10755) );
  NOR2_X1 U13137 ( .A1(n7505), .A2(n10755), .ZN(n10597) );
  XNOR2_X1 U13138 ( .A(n10754), .B(n10597), .ZN(n10609) );
  NAND2_X1 U13139 ( .A1(n11591), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13140 ( .A1(n9864), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10602) );
  NAND2_X1 U13141 ( .A1(n10598), .A2(n10768), .ZN(n10599) );
  AND2_X1 U13142 ( .A1(n10764), .A2(n10599), .ZN(n10982) );
  NAND2_X1 U13143 ( .A1(n11590), .A2(n10982), .ZN(n10601) );
  NAND2_X1 U13144 ( .A1(n11612), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10600) );
  NAND4_X1 U13145 ( .A1(n10603), .A2(n10602), .A3(n10601), .A4(n10600), .ZN(
        n12771) );
  NAND2_X1 U13146 ( .A1(n12771), .A2(n12824), .ZN(n10605) );
  NAND2_X1 U13147 ( .A1(n12773), .A2(n12754), .ZN(n10604) );
  AND2_X1 U13148 ( .A1(n10605), .A2(n10604), .ZN(n10738) );
  NAND2_X1 U13149 ( .A1(n12758), .A2(n10742), .ZN(n10606) );
  NAND2_X1 U13150 ( .A1(P2_U3088), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n10709)
         );
  OAI211_X1 U13151 ( .C1(n10738), .C2(n12744), .A(n10606), .B(n10709), .ZN(
        n10607) );
  AOI21_X1 U13152 ( .B1(n13172), .B2(n12747), .A(n10607), .ZN(n10608) );
  OAI21_X1 U13153 ( .B1(n10609), .B2(n12749), .A(n10608), .ZN(P2_U3196) );
  OAI21_X1 U13154 ( .B1(n14351), .B2(n10611), .A(n10610), .ZN(n14353) );
  MUX2_X1 U13155 ( .A(n10613), .B(n10612), .S(n9840), .Z(n10618) );
  OAI21_X1 U13156 ( .B1(n7321), .B2(n6624), .A(n10614), .ZN(n14356) );
  OAI22_X1 U13157 ( .A1(n10615), .A2(n13965), .B1(n9840), .B2(n13963), .ZN(
        n10616) );
  AOI21_X1 U13158 ( .B1(n14356), .B2(n14403), .A(n10616), .ZN(n10617) );
  OAI21_X1 U13159 ( .B1(n14379), .B2(n10618), .A(n10617), .ZN(n14354) );
  INV_X1 U13160 ( .A(n13725), .ZN(n13618) );
  AOI22_X1 U13161 ( .A1(n14304), .A2(n14356), .B1(n14310), .B2(n10619), .ZN(
        n10621) );
  AOI22_X1 U13162 ( .A1(n14315), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n14311), .ZN(n10620) );
  OAI211_X1 U13163 ( .C1(n13618), .C2(n14353), .A(n10621), .B(n10620), .ZN(
        n10622) );
  AOI21_X1 U13164 ( .B1(n13970), .B2(n14354), .A(n10622), .ZN(n10623) );
  INV_X1 U13165 ( .A(n10623), .ZN(P1_U3292) );
  AOI21_X1 U13166 ( .B1(n10626), .B2(n10625), .A(n10624), .ZN(n10642) );
  OAI21_X1 U13167 ( .B1(n10629), .B2(n10628), .A(n10627), .ZN(n10635) );
  INV_X1 U13168 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n10630) );
  NOR2_X1 U13169 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10630), .ZN(n10631) );
  AOI21_X1 U13170 ( .B1(n14664), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n10631), 
        .ZN(n10632) );
  OAI21_X1 U13171 ( .B1(n14719), .B2(n10633), .A(n10632), .ZN(n10634) );
  AOI21_X1 U13172 ( .B1(n10635), .B2(n14703), .A(n10634), .ZN(n10641) );
  INV_X1 U13173 ( .A(n10925), .ZN(n10639) );
  OAI21_X1 U13174 ( .B1(n10676), .B2(n10637), .A(n10636), .ZN(n10638) );
  NAND3_X1 U13175 ( .A1(n10639), .A2(n14713), .A3(n10638), .ZN(n10640) );
  OAI211_X1 U13176 ( .C1(n10642), .C2(n14708), .A(n10641), .B(n10640), .ZN(
        P3_U3194) );
  NAND2_X1 U13177 ( .A1(n10643), .A2(n13948), .ZN(n10644) );
  OAI211_X1 U13178 ( .C1(n10645), .C2(n12661), .A(n10644), .B(n12259), .ZN(
        P3_U3272) );
  XNOR2_X1 U13179 ( .A(n10646), .B(n10647), .ZN(n14369) );
  XNOR2_X1 U13180 ( .A(n10648), .B(n10647), .ZN(n14372) );
  AOI21_X1 U13181 ( .B1(n10649), .B2(n10652), .A(n14352), .ZN(n10651) );
  AND2_X1 U13182 ( .A1(n10651), .A2(n10650), .ZN(n14364) );
  AOI22_X1 U13183 ( .A1(n14364), .A2(n14313), .B1(n14310), .B2(n10652), .ZN(
        n10658) );
  INV_X1 U13184 ( .A(n10653), .ZN(n14365) );
  INV_X1 U13185 ( .A(n10654), .ZN(n10655) );
  OAI22_X1 U13186 ( .A1(n14315), .A2(n14365), .B1(n10655), .B2(n14093), .ZN(
        n10656) );
  INV_X1 U13187 ( .A(n10656), .ZN(n10657) );
  OAI211_X1 U13188 ( .C1(n10659), .C2(n13970), .A(n10658), .B(n10657), .ZN(
        n10660) );
  AOI21_X1 U13189 ( .B1(n13977), .B2(n14372), .A(n10660), .ZN(n10661) );
  OAI21_X1 U13190 ( .B1(n13675), .B2(n14369), .A(n10661), .ZN(P1_U3289) );
  XNOR2_X1 U13191 ( .A(n10662), .B(n12088), .ZN(n10670) );
  INV_X1 U13192 ( .A(n10670), .ZN(n14813) );
  INV_X1 U13193 ( .A(n14787), .ZN(n10832) );
  NAND2_X1 U13194 ( .A1(n10663), .A2(n14821), .ZN(n14810) );
  OAI22_X1 U13195 ( .A1(n10873), .A2(n14810), .B1(n10664), .B2(n14785), .ZN(
        n10672) );
  AOI22_X1 U13196 ( .A1(n14730), .A2(n12277), .B1(n10665), .B2(n14731), .ZN(
        n10669) );
  OAI211_X1 U13197 ( .C1(n10667), .C2(n12088), .A(n10666), .B(n14778), .ZN(
        n10668) );
  OAI211_X1 U13198 ( .C1(n10670), .C2(n14783), .A(n10669), .B(n10668), .ZN(
        n14811) );
  MUX2_X1 U13199 ( .A(n14811), .B(P3_REG2_REG_4__SCAN_IN), .S(n14793), .Z(
        n10671) );
  AOI211_X1 U13200 ( .C1(n14813), .C2(n10832), .A(n10672), .B(n10671), .ZN(
        n10673) );
  INV_X1 U13201 ( .A(n10673), .ZN(P3_U3229) );
  AOI21_X1 U13202 ( .B1(n11057), .B2(n10675), .A(n10674), .ZN(n10688) );
  INV_X1 U13203 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n13860) );
  NAND2_X1 U13204 ( .A1(P3_REG3_REG_11__SCAN_IN), .A2(P3_U3151), .ZN(n11213)
         );
  OAI21_X1 U13205 ( .B1(n14724), .B2(n13860), .A(n11213), .ZN(n10681) );
  AOI21_X1 U13206 ( .B1(n10678), .B2(n10677), .A(n10676), .ZN(n10679) );
  NOR2_X1 U13207 ( .A1(n10679), .A2(n14036), .ZN(n10680) );
  AOI211_X1 U13208 ( .C1(n14686), .C2(n10682), .A(n10681), .B(n10680), .ZN(
        n10687) );
  OAI21_X1 U13209 ( .B1(n10684), .B2(P3_REG1_REG_11__SCAN_IN), .A(n10683), 
        .ZN(n10685) );
  NAND2_X1 U13210 ( .A1(n10685), .A2(n14703), .ZN(n10686) );
  OAI211_X1 U13211 ( .C1(n10688), .C2(n14708), .A(n10687), .B(n10686), .ZN(
        P3_U3193) );
  NOR2_X1 U13212 ( .A1(n11815), .A2(n10692), .ZN(n10693) );
  AOI21_X1 U13213 ( .B1(n14396), .B2(n6452), .A(n10693), .ZN(n10845) );
  AOI22_X1 U13214 ( .A1(n14396), .A2(n9889), .B1(n6452), .B2(n13348), .ZN(
        n10694) );
  XNOR2_X1 U13215 ( .A(n10694), .B(n11856), .ZN(n10846) );
  XOR2_X1 U13216 ( .A(n10845), .B(n10846), .Z(n10849) );
  XNOR2_X1 U13217 ( .A(n10850), .B(n10849), .ZN(n10700) );
  NAND2_X1 U13218 ( .A1(n14075), .A2(n14396), .ZN(n10695) );
  NAND2_X1 U13219 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n13423) );
  OAI211_X1 U13220 ( .C1(n10696), .C2(n13334), .A(n10695), .B(n13423), .ZN(
        n10697) );
  AOI21_X1 U13221 ( .B1(n10698), .B2(n13326), .A(n10697), .ZN(n10699) );
  OAI21_X1 U13222 ( .B1(n10700), .B2(n14078), .A(n10699), .ZN(P1_U3213) );
  XOR2_X1 U13223 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n10882), .Z(n10703) );
  OAI21_X1 U13224 ( .B1(n10703), .B2(n10702), .A(n10881), .ZN(n10704) );
  INV_X1 U13225 ( .A(n10704), .ZN(n10715) );
  XOR2_X1 U13226 ( .A(n10882), .B(P2_REG1_REG_12__SCAN_IN), .Z(n10708) );
  OAI21_X1 U13227 ( .B1(n10708), .B2(n10707), .A(n10878), .ZN(n10713) );
  NAND2_X1 U13228 ( .A1(n14442), .A2(P2_ADDR_REG_12__SCAN_IN), .ZN(n10710) );
  OAI211_X1 U13229 ( .C1(n12815), .C2(n10711), .A(n10710), .B(n10709), .ZN(
        n10712) );
  AOI21_X1 U13230 ( .B1(n10713), .B2(n12814), .A(n10712), .ZN(n10714) );
  OAI21_X1 U13231 ( .B1(n10715), .B2(n14527), .A(n10714), .ZN(P2_U3226) );
  INV_X1 U13232 ( .A(n14583), .ZN(n14614) );
  OAI211_X1 U13233 ( .C1(n10736), .C2(n14627), .A(n10717), .B(n10716), .ZN(
        n10718) );
  AOI21_X1 U13234 ( .B1(n14614), .B2(n10719), .A(n10718), .ZN(n10722) );
  NAND2_X1 U13235 ( .A1(n14661), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n10720) );
  OAI21_X1 U13236 ( .B1(n10722), .B2(n14661), .A(n10720), .ZN(P2_U3510) );
  NAND2_X1 U13237 ( .A1(n14646), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n10721) );
  OAI21_X1 U13238 ( .B1(n10722), .B2(n14646), .A(n10721), .ZN(P2_U3463) );
  INV_X1 U13239 ( .A(n10723), .ZN(n10724) );
  AOI211_X1 U13240 ( .C1(n10726), .C2(n10725), .A(n12023), .B(n10724), .ZN(
        n10733) );
  NAND2_X1 U13241 ( .A1(n12107), .A2(n14730), .ZN(n10727) );
  OAI21_X1 U13242 ( .B1(n10728), .B2(n14762), .A(n10727), .ZN(n14751) );
  AOI21_X1 U13243 ( .B1(n12019), .B2(n14751), .A(n10729), .ZN(n10731) );
  NAND2_X1 U13244 ( .A1(n14675), .A2(n14820), .ZN(n10730) );
  OAI211_X1 U13245 ( .C1(n14678), .C2(n14756), .A(n10731), .B(n10730), .ZN(
        n10732) );
  OR2_X1 U13246 ( .A1(n10733), .A2(n10732), .ZN(P3_U3179) );
  INV_X1 U13247 ( .A(n12772), .ZN(n10734) );
  XNOR2_X1 U13248 ( .A(n13172), .B(n10734), .ZN(n11659) );
  AOI211_X1 U13249 ( .C1(n11659), .C2(n10737), .A(n12946), .B(n6602), .ZN(
        n10740) );
  INV_X1 U13250 ( .A(n10738), .ZN(n10739) );
  NOR2_X1 U13251 ( .A1(n10740), .A2(n10739), .ZN(n13174) );
  AOI211_X1 U13252 ( .C1(n13172), .C2(n10741), .A(n9339), .B(n7081), .ZN(
        n13171) );
  INV_X1 U13253 ( .A(n13172), .ZN(n10984) );
  AOI22_X1 U13254 ( .A1(n14557), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n10742), 
        .B2(n14553), .ZN(n10743) );
  OAI21_X1 U13255 ( .B1(n10984), .B2(n13076), .A(n10743), .ZN(n10752) );
  INV_X1 U13256 ( .A(n11659), .ZN(n10750) );
  OR2_X1 U13257 ( .A1(n11374), .A2(n12773), .ZN(n10744) );
  NAND2_X1 U13258 ( .A1(n10745), .A2(n10744), .ZN(n10747) );
  NAND2_X1 U13259 ( .A1(n11374), .A2(n12773), .ZN(n10746) );
  INV_X1 U13260 ( .A(n10980), .ZN(n10748) );
  AOI21_X1 U13261 ( .B1(n10750), .B2(n10749), .A(n10748), .ZN(n13175) );
  NOR2_X1 U13262 ( .A1(n13175), .A2(n13081), .ZN(n10751) );
  AOI211_X1 U13263 ( .C1(n13171), .C2(n13078), .A(n10752), .B(n10751), .ZN(
        n10753) );
  OAI21_X1 U13264 ( .B1(n13174), .B2(n14557), .A(n10753), .ZN(P2_U3253) );
  NAND2_X1 U13265 ( .A1(n10757), .A2(n11584), .ZN(n10762) );
  OAI22_X1 U13266 ( .A1(n10888), .A2(n11026), .B1(n11608), .B2(n10759), .ZN(
        n10760) );
  INV_X1 U13267 ( .A(n10760), .ZN(n10761) );
  NAND2_X1 U13268 ( .A1(n12771), .A2(n9339), .ZN(n10948) );
  XNOR2_X1 U13269 ( .A(n10949), .B(n10948), .ZN(n10950) );
  XNOR2_X1 U13270 ( .A(n10951), .B(n10950), .ZN(n10772) );
  INV_X1 U13271 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10763) );
  AND2_X1 U13272 ( .A1(n10764), .A2(n10763), .ZN(n10765) );
  OR2_X1 U13273 ( .A1(n10765), .A2(n10954), .ZN(n11013) );
  AOI22_X1 U13274 ( .A1(n11591), .A2(P2_REG1_REG_14__SCAN_IN), .B1(n9864), 
        .B2(P2_REG2_REG_14__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13275 ( .A1(n11612), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10766) );
  OAI211_X1 U13276 ( .C1(n11013), .C2(n11459), .A(n10767), .B(n10766), .ZN(
        n12770) );
  AOI22_X1 U13277 ( .A1(n12770), .A2(n12824), .B1(n12754), .B2(n12772), .ZN(
        n10986) );
  OAI22_X1 U13278 ( .A1(n12744), .A2(n10986), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10768), .ZN(n10770) );
  INV_X1 U13279 ( .A(n13167), .ZN(n11010) );
  NOR2_X1 U13280 ( .A1(n11010), .A2(n12761), .ZN(n10769) );
  AOI211_X1 U13281 ( .C1(n12758), .C2(n10982), .A(n10770), .B(n10769), .ZN(
        n10771) );
  OAI21_X1 U13282 ( .B1(n10772), .B2(n12749), .A(n10771), .ZN(P2_U3206) );
  INV_X1 U13283 ( .A(n12218), .ZN(n10773) );
  XNOR2_X1 U13284 ( .A(n10774), .B(n10773), .ZN(n10786) );
  INV_X1 U13285 ( .A(n10786), .ZN(n14818) );
  NAND2_X1 U13286 ( .A1(n10775), .A2(n14821), .ZN(n14815) );
  OAI22_X1 U13287 ( .A1(n10873), .A2(n14815), .B1(n10776), .B2(n14785), .ZN(
        n10788) );
  NAND2_X1 U13288 ( .A1(n10777), .A2(n12218), .ZN(n10778) );
  NAND2_X1 U13289 ( .A1(n10779), .A2(n10778), .ZN(n10780) );
  NAND2_X1 U13290 ( .A1(n10780), .A2(n14778), .ZN(n10785) );
  OAI22_X1 U13291 ( .A1(n10782), .A2(n14762), .B1(n10781), .B2(n14760), .ZN(
        n10783) );
  INV_X1 U13292 ( .A(n10783), .ZN(n10784) );
  OAI211_X1 U13293 ( .C1(n10786), .C2(n14783), .A(n10785), .B(n10784), .ZN(
        n14816) );
  MUX2_X1 U13294 ( .A(n14816), .B(P3_REG2_REG_5__SCAN_IN), .S(n14793), .Z(
        n10787) );
  AOI211_X1 U13295 ( .C1(n14818), .C2(n10832), .A(n10788), .B(n10787), .ZN(
        n10789) );
  INV_X1 U13296 ( .A(n10789), .ZN(P3_U3228) );
  INV_X1 U13297 ( .A(n13344), .ZN(n11140) );
  OR2_X1 U13298 ( .A1(n11100), .A2(n11140), .ZN(n10792) );
  NAND2_X1 U13299 ( .A1(n10793), .A2(n10792), .ZN(n10807) );
  INV_X1 U13300 ( .A(n10816), .ZN(n10806) );
  XNOR2_X1 U13301 ( .A(n10807), .B(n10806), .ZN(n10798) );
  XNOR2_X1 U13302 ( .A(n10817), .B(n10816), .ZN(n13960) );
  NAND2_X1 U13303 ( .A1(n13960), .A2(n14403), .ZN(n10797) );
  AOI22_X1 U13304 ( .A1(n14087), .A2(n13344), .B1(n13342), .B2(n6454), .ZN(
        n10796) );
  OAI211_X1 U13305 ( .C1(n14379), .C2(n10798), .A(n10797), .B(n10796), .ZN(
        n13958) );
  INV_X1 U13306 ( .A(n13958), .ZN(n10805) );
  INV_X1 U13307 ( .A(n10799), .ZN(n10800) );
  INV_X1 U13308 ( .A(n11131), .ZN(n13957) );
  OR2_X2 U13309 ( .A1(n10799), .A2(n11131), .ZN(n13973) );
  OAI211_X1 U13310 ( .C1(n10800), .C2(n13957), .A(n9843), .B(n13973), .ZN(
        n13956) );
  AOI22_X1 U13311 ( .A1(n14322), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11142), 
        .B2(n14311), .ZN(n10802) );
  NAND2_X1 U13312 ( .A1(n11131), .A2(n14310), .ZN(n10801) );
  OAI211_X1 U13313 ( .C1(n13956), .C2(n13720), .A(n10802), .B(n10801), .ZN(
        n10803) );
  AOI21_X1 U13314 ( .B1(n13960), .B2(n14304), .A(n10803), .ZN(n10804) );
  OAI21_X1 U13315 ( .B1(n10805), .B2(n14322), .A(n10804), .ZN(P1_U3281) );
  NAND2_X1 U13316 ( .A1(n10807), .A2(n10806), .ZN(n10809) );
  OR2_X1 U13317 ( .A1(n11131), .A2(n13964), .ZN(n10808) );
  INV_X1 U13318 ( .A(n13971), .ZN(n13975) );
  XNOR2_X1 U13319 ( .A(n10993), .B(n10820), .ZN(n10812) );
  NAND2_X1 U13320 ( .A1(n14088), .A2(n6454), .ZN(n10810) );
  OAI21_X1 U13321 ( .B1(n11200), .B2(n13963), .A(n10810), .ZN(n10811) );
  AOI21_X1 U13322 ( .B1(n10812), .B2(n14373), .A(n10811), .ZN(n14142) );
  INV_X1 U13323 ( .A(n11000), .ZN(n11001) );
  AOI21_X1 U13324 ( .B1(n14136), .B2(n10813), .A(n11001), .ZN(n14137) );
  AOI22_X1 U13325 ( .A1(n14315), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n13230), 
        .B2(n14311), .ZN(n10814) );
  OAI21_X1 U13326 ( .B1(n7026), .B2(n14298), .A(n10814), .ZN(n10815) );
  AOI21_X1 U13327 ( .B1(n14137), .B2(n13725), .A(n10815), .ZN(n10823) );
  OR2_X1 U13328 ( .A1(n11131), .A2(n13343), .ZN(n10818) );
  OR2_X1 U13329 ( .A1(n14145), .A2(n13342), .ZN(n10819) );
  INV_X1 U13330 ( .A(n10820), .ZN(n10992) );
  NAND2_X1 U13331 ( .A1(n10821), .A2(n10992), .ZN(n14138) );
  NAND3_X1 U13332 ( .A1(n14139), .A2(n14138), .A3(n14308), .ZN(n10822) );
  OAI211_X1 U13333 ( .C1(n14142), .C2(n14315), .A(n10823), .B(n10822), .ZN(
        P1_U3279) );
  INV_X1 U13334 ( .A(n14679), .ZN(n10829) );
  XNOR2_X1 U13335 ( .A(n10824), .B(n12226), .ZN(n14827) );
  OAI211_X1 U13336 ( .C1(n10825), .C2(n12226), .A(n10864), .B(n14778), .ZN(
        n10828) );
  NAND2_X1 U13337 ( .A1(n12276), .A2(n14731), .ZN(n10827) );
  NAND2_X1 U13338 ( .A1(n12275), .A2(n14730), .ZN(n10826) );
  AND2_X1 U13339 ( .A1(n10827), .A2(n10826), .ZN(n14667) );
  OAI211_X1 U13340 ( .C1(n14783), .C2(n14827), .A(n10828), .B(n14667), .ZN(
        n14829) );
  AOI21_X1 U13341 ( .B1(n14772), .B2(n10829), .A(n14829), .ZN(n10835) );
  INV_X1 U13342 ( .A(n14827), .ZN(n10833) );
  INV_X1 U13343 ( .A(n6433), .ZN(n12355) );
  OAI22_X1 U13344 ( .A1(n12355), .A2(n14826), .B1(n10830), .B2(n14791), .ZN(
        n10831) );
  AOI21_X1 U13345 ( .B1(n10833), .B2(n10832), .A(n10831), .ZN(n10834) );
  OAI21_X1 U13346 ( .B1(n10835), .B2(n14793), .A(n10834), .ZN(P3_U3226) );
  OAI211_X1 U13347 ( .C1(n10838), .C2(n10837), .A(n10836), .B(n14668), .ZN(
        n10843) );
  OAI22_X1 U13348 ( .A1(n11974), .A2(n10839), .B1(n11072), .B2(n12000), .ZN(
        n10840) );
  AOI211_X1 U13349 ( .C1(n10871), .C2(n14675), .A(n10841), .B(n10840), .ZN(
        n10842) );
  OAI211_X1 U13350 ( .C1(n7599), .C2(n14678), .A(n10843), .B(n10842), .ZN(
        P3_U3161) );
  AOI22_X1 U13351 ( .A1(n10858), .A2(n6452), .B1(n11858), .B2(n13347), .ZN(
        n10892) );
  AOI22_X1 U13352 ( .A1(n10858), .A2(n9889), .B1(n6452), .B2(n13347), .ZN(
        n10844) );
  XNOR2_X1 U13353 ( .A(n10844), .B(n11856), .ZN(n10893) );
  XOR2_X1 U13354 ( .A(n10892), .B(n10893), .Z(n10852) );
  INV_X1 U13355 ( .A(n10845), .ZN(n10848) );
  INV_X1 U13356 ( .A(n10846), .ZN(n10847) );
  OAI21_X1 U13357 ( .B1(n10852), .B2(n10851), .A(n10899), .ZN(n10853) );
  NAND2_X1 U13358 ( .A1(n10853), .A2(n13320), .ZN(n10860) );
  INV_X1 U13359 ( .A(n10854), .ZN(n10856) );
  OAI21_X1 U13360 ( .B1(n13334), .B2(n10856), .A(n10855), .ZN(n10857) );
  AOI21_X1 U13361 ( .B1(n14075), .B2(n10858), .A(n10857), .ZN(n10859) );
  OAI211_X1 U13362 ( .C1(n14083), .C2(n10861), .A(n10860), .B(n10859), .ZN(
        P1_U3221) );
  XNOR2_X1 U13363 ( .A(n10862), .B(n12222), .ZN(n14834) );
  INV_X1 U13364 ( .A(n14834), .ZN(n10877) );
  NAND2_X1 U13365 ( .A1(n10864), .A2(n10863), .ZN(n10867) );
  INV_X1 U13366 ( .A(n10865), .ZN(n10866) );
  AOI21_X1 U13367 ( .B1(n12222), .B2(n10867), .A(n10866), .ZN(n10870) );
  AOI22_X1 U13368 ( .A1(n14732), .A2(n14730), .B1(n14731), .B2(n12107), .ZN(
        n10869) );
  NAND2_X1 U13369 ( .A1(n14834), .A2(n14843), .ZN(n10868) );
  OAI211_X1 U13370 ( .C1(n10870), .C2(n12418), .A(n10869), .B(n10868), .ZN(
        n14831) );
  NAND2_X1 U13371 ( .A1(n14831), .A2(n14791), .ZN(n10876) );
  AND2_X1 U13372 ( .A1(n10871), .A2(n14821), .ZN(n14832) );
  INV_X1 U13373 ( .A(n14832), .ZN(n10872) );
  OAI22_X1 U13374 ( .A1(n10873), .A2(n10872), .B1(n7599), .B2(n14785), .ZN(
        n10874) );
  AOI21_X1 U13375 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14793), .A(n10874), .ZN(
        n10875) );
  OAI211_X1 U13376 ( .C1(n10877), .C2(n14787), .A(n10876), .B(n10875), .ZN(
        P3_U3225) );
  XNOR2_X1 U13377 ( .A(n12796), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n10880) );
  OAI21_X1 U13378 ( .B1(n10882), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10878), 
        .ZN(n10879) );
  NOR2_X1 U13379 ( .A1(n10879), .A2(n10880), .ZN(n12795) );
  AOI211_X1 U13380 ( .C1(n10880), .C2(n10879), .A(n14531), .B(n12795), .ZN(
        n10891) );
  OAI21_X1 U13381 ( .B1(n10882), .B2(P2_REG2_REG_12__SCAN_IN), .A(n10881), 
        .ZN(n10885) );
  NAND2_X1 U13382 ( .A1(n12796), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10883) );
  OAI21_X1 U13383 ( .B1(n12796), .B2(P2_REG2_REG_13__SCAN_IN), .A(n10883), 
        .ZN(n10884) );
  NOR2_X1 U13384 ( .A1(n10885), .A2(n10884), .ZN(n12784) );
  AOI211_X1 U13385 ( .C1(n10885), .C2(n10884), .A(n14527), .B(n12784), .ZN(
        n10890) );
  NAND2_X1 U13386 ( .A1(n14442), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n10887) );
  NAND2_X1 U13387 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n10886)
         );
  OAI211_X1 U13388 ( .C1(n12815), .C2(n10888), .A(n10887), .B(n10886), .ZN(
        n10889) );
  OR3_X1 U13389 ( .A1(n10891), .A2(n10890), .A3(n10889), .ZN(P2_U3227) );
  NAND2_X1 U13390 ( .A1(n10893), .A2(n10892), .ZN(n10897) );
  AND2_X1 U13391 ( .A1(n10899), .A2(n10897), .ZN(n10901) );
  OAI22_X1 U13392 ( .A1(n14412), .A2(n11824), .B1(n10974), .B2(n11823), .ZN(
        n10894) );
  XNOR2_X1 U13393 ( .A(n10894), .B(n11813), .ZN(n10963) );
  OR2_X1 U13394 ( .A1(n14412), .A2(n11823), .ZN(n10896) );
  NAND2_X1 U13395 ( .A1(n11858), .A2(n13346), .ZN(n10895) );
  NAND2_X1 U13396 ( .A1(n10896), .A2(n10895), .ZN(n10964) );
  XNOR2_X1 U13397 ( .A(n10963), .B(n10964), .ZN(n10900) );
  AND2_X1 U13398 ( .A1(n10900), .A2(n10897), .ZN(n10898) );
  OAI211_X1 U13399 ( .C1(n10901), .C2(n10900), .A(n13320), .B(n10967), .ZN(
        n10908) );
  INV_X1 U13400 ( .A(n14073), .ZN(n13267) );
  AOI21_X1 U13401 ( .B1(n14074), .B2(n13345), .A(n10902), .ZN(n10903) );
  OAI21_X1 U13402 ( .B1(n10904), .B2(n13267), .A(n10903), .ZN(n10905) );
  AOI21_X1 U13403 ( .B1(n10906), .B2(n13326), .A(n10905), .ZN(n10907) );
  OAI211_X1 U13404 ( .C1(n14412), .C2(n13329), .A(n10908), .B(n10907), .ZN(
        P1_U3231) );
  NAND2_X1 U13405 ( .A1(n11499), .A2(n10909), .ZN(n10911) );
  NOR2_X1 U13406 ( .A1(n10910), .A2(P2_U3088), .ZN(n11684) );
  INV_X1 U13407 ( .A(n11684), .ZN(n11687) );
  OAI211_X1 U13408 ( .C1(n11500), .C2(n13210), .A(n10911), .B(n11687), .ZN(
        P2_U3304) );
  NAND2_X1 U13409 ( .A1(n11499), .A2(n10912), .ZN(n10914) );
  OAI211_X1 U13410 ( .C1(n10915), .C2(n13833), .A(n10914), .B(n10913), .ZN(
        P1_U3332) );
  AOI21_X1 U13411 ( .B1(n14910), .B2(n10917), .A(n10916), .ZN(n10932) );
  OAI21_X1 U13412 ( .B1(P3_REG1_REG_13__SCAN_IN), .B2(n10919), .A(n10918), 
        .ZN(n10930) );
  AND2_X1 U13413 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n10920) );
  AOI21_X1 U13414 ( .B1(n14664), .B2(P3_ADDR_REG_13__SCAN_IN), .A(n10920), 
        .ZN(n10921) );
  OAI21_X1 U13415 ( .B1(n14719), .B2(n10922), .A(n10921), .ZN(n10929) );
  INV_X1 U13416 ( .A(n11087), .ZN(n10927) );
  OAI21_X1 U13417 ( .B1(n10925), .B2(n10924), .A(n10923), .ZN(n10926) );
  AOI21_X1 U13418 ( .B1(n10927), .B2(n10926), .A(n14036), .ZN(n10928) );
  AOI211_X1 U13419 ( .C1(n10930), .C2(n14703), .A(n10929), .B(n10928), .ZN(
        n10931) );
  OAI21_X1 U13420 ( .B1(n10932), .B2(n14708), .A(n10931), .ZN(P3_U3195) );
  XNOR2_X1 U13421 ( .A(n10933), .B(n12227), .ZN(n14839) );
  OAI211_X1 U13422 ( .C1(n10935), .C2(n12227), .A(n10934), .B(n14778), .ZN(
        n10937) );
  NAND2_X1 U13423 ( .A1(n10937), .A2(n10936), .ZN(n14840) );
  NAND2_X1 U13424 ( .A1(n14840), .A2(n14791), .ZN(n10941) );
  OAI22_X1 U13425 ( .A1(n14791), .A2(n14976), .B1(n10938), .B2(n14785), .ZN(
        n10939) );
  AOI21_X1 U13426 ( .B1(n12118), .B2(n6433), .A(n10939), .ZN(n10940) );
  OAI211_X1 U13427 ( .C1(n12493), .C2(n14839), .A(n10941), .B(n10940), .ZN(
        P3_U3224) );
  NAND2_X1 U13428 ( .A1(n10942), .A2(n11584), .ZN(n10944) );
  AOI22_X1 U13429 ( .A1(n14497), .A2(n11433), .B1(n11434), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n10943) );
  XNOR2_X1 U13430 ( .A(n11394), .B(n11724), .ZN(n10945) );
  NAND2_X1 U13431 ( .A1(n12770), .A2(n9339), .ZN(n10946) );
  NAND2_X1 U13432 ( .A1(n10945), .A2(n10946), .ZN(n11060) );
  NAND2_X1 U13433 ( .A1(n11060), .A2(n10947), .ZN(n10953) );
  AOI21_X1 U13434 ( .B1(n10953), .B2(n10952), .A(n6600), .ZN(n10962) );
  NOR2_X1 U13435 ( .A1(n12742), .A2(n11013), .ZN(n10960) );
  NAND2_X1 U13436 ( .A1(n10954), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n11032) );
  OR2_X1 U13437 ( .A1(n10954), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10955) );
  NAND2_X1 U13438 ( .A1(n11032), .A2(n10955), .ZN(n11063) );
  AOI22_X1 U13439 ( .A1(n11591), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n9864), 
        .B2(P2_REG2_REG_15__SCAN_IN), .ZN(n10957) );
  NAND2_X1 U13440 ( .A1(n11612), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10956) );
  OAI211_X1 U13441 ( .C1(n11063), .C2(n11459), .A(n10957), .B(n10956), .ZN(
        n12856) );
  AND2_X1 U13442 ( .A1(n12771), .A2(n12754), .ZN(n10958) );
  AOI21_X1 U13443 ( .B1(n12856), .B2(n12824), .A(n10958), .ZN(n11011) );
  NAND2_X1 U13444 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14498)
         );
  OAI21_X1 U13445 ( .B1(n12744), .B2(n11011), .A(n14498), .ZN(n10959) );
  AOI211_X1 U13446 ( .C1(n11394), .C2(n12747), .A(n10960), .B(n10959), .ZN(
        n10961) );
  OAI21_X1 U13447 ( .B1(n10962), .B2(n12749), .A(n10961), .ZN(P2_U3187) );
  INV_X1 U13448 ( .A(n10963), .ZN(n10965) );
  NAND2_X1 U13449 ( .A1(n10967), .A2(n10966), .ZN(n11102) );
  NOR2_X1 U13450 ( .A1(n11815), .A2(n10968), .ZN(n10969) );
  AOI21_X1 U13451 ( .B1(n10976), .B2(n6452), .A(n10969), .ZN(n11104) );
  AOI22_X1 U13452 ( .A1(n10976), .A2(n9889), .B1(n6452), .B2(n13345), .ZN(
        n10970) );
  XNOR2_X1 U13453 ( .A(n10970), .B(n11856), .ZN(n11103) );
  XOR2_X1 U13454 ( .A(n11104), .B(n11103), .Z(n11101) );
  XNOR2_X1 U13455 ( .A(n11102), .B(n11101), .ZN(n10978) );
  AOI22_X1 U13456 ( .A1(n14074), .A2(n13344), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10973) );
  NAND2_X1 U13457 ( .A1(n13326), .A2(n10971), .ZN(n10972) );
  OAI211_X1 U13458 ( .C1(n10974), .C2(n13267), .A(n10973), .B(n10972), .ZN(
        n10975) );
  AOI21_X1 U13459 ( .B1(n14075), .B2(n10976), .A(n10975), .ZN(n10977) );
  OAI21_X1 U13460 ( .B1(n10978), .B2(n14078), .A(n10977), .ZN(P1_U3217) );
  INV_X1 U13461 ( .A(n12771), .ZN(n11390) );
  XNOR2_X1 U13462 ( .A(n13167), .B(n11390), .ZN(n11661) );
  OR2_X1 U13463 ( .A1(n13172), .A2(n12772), .ZN(n10979) );
  XOR2_X1 U13464 ( .A(n11661), .B(n11008), .Z(n13170) );
  AOI211_X1 U13465 ( .C1(n13167), .C2(n10981), .A(n9339), .B(n6611), .ZN(
        n13166) );
  AOI22_X1 U13466 ( .A1(n14557), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10982), 
        .B2(n14553), .ZN(n10983) );
  OAI21_X1 U13467 ( .B1(n11010), .B2(n13076), .A(n10983), .ZN(n10990) );
  AOI211_X1 U13468 ( .C1(n11661), .C2(n10985), .A(n12946), .B(n11009), .ZN(
        n10988) );
  INV_X1 U13469 ( .A(n10986), .ZN(n10987) );
  NOR2_X1 U13470 ( .A1(n10988), .A2(n10987), .ZN(n13169) );
  NOR2_X1 U13471 ( .A1(n13169), .A2(n14557), .ZN(n10989) );
  AOI211_X1 U13472 ( .C1(n13166), .C2(n13078), .A(n10990), .B(n10989), .ZN(
        n10991) );
  OAI21_X1 U13473 ( .B1(n13081), .B2(n13170), .A(n10991), .ZN(P2_U3252) );
  XNOR2_X1 U13474 ( .A(n11146), .B(n6901), .ZN(n10996) );
  NAND2_X1 U13475 ( .A1(n10996), .A2(n14373), .ZN(n10998) );
  NOR2_X1 U13476 ( .A1(n13966), .A2(n13963), .ZN(n10997) );
  AOI21_X1 U13477 ( .B1(n13340), .B2(n6454), .A(n10997), .ZN(n13333) );
  NAND2_X1 U13478 ( .A1(n10998), .A2(n13333), .ZN(n14133) );
  INV_X1 U13479 ( .A(n14133), .ZN(n11007) );
  INV_X1 U13480 ( .A(n13966), .ZN(n13341) );
  NAND2_X1 U13481 ( .A1(n14136), .A2(n13341), .ZN(n10999) );
  OAI21_X1 U13482 ( .B1(n6601), .B2(n6901), .A(n11155), .ZN(n14135) );
  INV_X1 U13483 ( .A(n13337), .ZN(n14132) );
  INV_X1 U13484 ( .A(n11159), .ZN(n14090) );
  OAI211_X1 U13485 ( .C1(n14132), .C2(n11001), .A(n14090), .B(n9843), .ZN(
        n14131) );
  INV_X1 U13486 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11002) );
  OAI22_X1 U13487 ( .A1(n13970), .A2(n11002), .B1(n13332), .B2(n14093), .ZN(
        n11003) );
  AOI21_X1 U13488 ( .B1(n13337), .B2(n14310), .A(n11003), .ZN(n11004) );
  OAI21_X1 U13489 ( .B1(n14131), .B2(n13720), .A(n11004), .ZN(n11005) );
  AOI21_X1 U13490 ( .B1(n14135), .B2(n14308), .A(n11005), .ZN(n11006) );
  OAI21_X1 U13491 ( .B1(n14322), .B2(n11007), .A(n11006), .ZN(P1_U3278) );
  OR2_X1 U13492 ( .A1(n11394), .A2(n12770), .ZN(n11043) );
  NAND2_X1 U13493 ( .A1(n11394), .A2(n12770), .ZN(n11045) );
  NAND2_X1 U13494 ( .A1(n11043), .A2(n11045), .ZN(n11662) );
  XOR2_X1 U13495 ( .A(n11044), .B(n11662), .Z(n13164) );
  INV_X1 U13496 ( .A(n13164), .ZN(n11020) );
  XOR2_X1 U13497 ( .A(n11662), .B(n11023), .Z(n11012) );
  OAI21_X1 U13498 ( .B1(n11012), .B2(n12946), .A(n11011), .ZN(n13162) );
  NAND2_X1 U13499 ( .A1(n13162), .A2(n14554), .ZN(n11019) );
  INV_X1 U13500 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n11014) );
  OAI22_X1 U13501 ( .A1(n14554), .A2(n11014), .B1(n11013), .B2(n13071), .ZN(
        n11016) );
  INV_X1 U13502 ( .A(n11394), .ZN(n13161) );
  OAI211_X1 U13503 ( .C1(n13161), .C2(n6611), .A(n11040), .B(n12952), .ZN(
        n13160) );
  NOR2_X1 U13504 ( .A1(n13160), .A2(n12953), .ZN(n11015) );
  AOI211_X1 U13505 ( .C1(n11017), .C2(n11394), .A(n11016), .B(n11015), .ZN(
        n11018) );
  OAI211_X1 U13506 ( .C1(n11020), .C2(n13081), .A(n11019), .B(n11018), .ZN(
        P2_U3251) );
  NOR2_X1 U13507 ( .A1(n13161), .A2(n12770), .ZN(n11022) );
  INV_X1 U13508 ( .A(n12770), .ZN(n11021) );
  NAND2_X1 U13509 ( .A1(n11024), .A2(n11584), .ZN(n11029) );
  OAI22_X1 U13510 ( .A1(n14501), .A2(n11026), .B1(n11608), .B2(n11025), .ZN(
        n11027) );
  INV_X1 U13511 ( .A(n11027), .ZN(n11028) );
  INV_X1 U13512 ( .A(n12856), .ZN(n11030) );
  XNOR2_X1 U13513 ( .A(n12834), .B(n12832), .ZN(n11038) );
  INV_X1 U13514 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n11031) );
  NAND2_X1 U13515 ( .A1(n11032), .A2(n11031), .ZN(n11033) );
  NAND2_X1 U13516 ( .A1(n11182), .A2(n11033), .ZN(n13072) );
  AOI22_X1 U13517 ( .A1(n11591), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n9864), 
        .B2(P2_REG2_REG_16__SCAN_IN), .ZN(n11035) );
  NAND2_X1 U13518 ( .A1(n11612), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n11034) );
  OAI211_X1 U13519 ( .C1(n13072), .C2(n11459), .A(n11035), .B(n11034), .ZN(
        n12860) );
  NAND2_X1 U13520 ( .A1(n12860), .A2(n12824), .ZN(n11037) );
  NAND2_X1 U13521 ( .A1(n12770), .A2(n12754), .ZN(n11036) );
  NAND2_X1 U13522 ( .A1(n11037), .A2(n11036), .ZN(n11061) );
  AOI21_X1 U13523 ( .B1(n11038), .B2(n14548), .A(n11061), .ZN(n13158) );
  INV_X1 U13524 ( .A(n13075), .ZN(n11039) );
  AOI211_X1 U13525 ( .C1(n13156), .C2(n11040), .A(n9339), .B(n11039), .ZN(
        n13155) );
  INV_X1 U13526 ( .A(n13156), .ZN(n12833) );
  INV_X1 U13527 ( .A(n11063), .ZN(n11041) );
  AOI22_X1 U13528 ( .A1(n14557), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n11041), 
        .B2(n14553), .ZN(n11042) );
  OAI21_X1 U13529 ( .B1(n12833), .B2(n13076), .A(n11042), .ZN(n11048) );
  XNOR2_X1 U13530 ( .A(n12859), .B(n12832), .ZN(n13159) );
  NOR2_X1 U13531 ( .A1(n13159), .A2(n13081), .ZN(n11047) );
  AOI211_X1 U13532 ( .C1(n13155), .C2(n13078), .A(n11048), .B(n11047), .ZN(
        n11049) );
  OAI21_X1 U13533 ( .B1(n13158), .B2(n14557), .A(n11049), .ZN(P2_U3250) );
  XNOR2_X1 U13534 ( .A(n11050), .B(n12229), .ZN(n11053) );
  OAI22_X1 U13535 ( .A1(n11985), .A2(n14760), .B1(n11051), .B2(n14762), .ZN(
        n11052) );
  AOI21_X1 U13536 ( .B1(n11053), .B2(n14778), .A(n11052), .ZN(n14062) );
  XNOR2_X1 U13537 ( .A(n11054), .B(n12229), .ZN(n14060) );
  INV_X1 U13538 ( .A(n12493), .ZN(n14737) );
  AND2_X1 U13539 ( .A1(n11212), .A2(n14821), .ZN(n14059) );
  INV_X1 U13540 ( .A(n11055), .ZN(n11216) );
  AOI22_X1 U13541 ( .A1(n14726), .A2(n14059), .B1(n14772), .B2(n11216), .ZN(
        n11056) );
  OAI21_X1 U13542 ( .B1(n11057), .B2(n14791), .A(n11056), .ZN(n11058) );
  AOI21_X1 U13543 ( .B1(n14060), .B2(n14737), .A(n11058), .ZN(n11059) );
  OAI21_X1 U13544 ( .B1(n14062), .B2(n14793), .A(n11059), .ZN(P3_U3222) );
  XOR2_X1 U13545 ( .A(n11729), .B(n13156), .Z(n11176) );
  XNOR2_X1 U13546 ( .A(n11175), .B(n11176), .ZN(n11178) );
  NAND2_X1 U13547 ( .A1(n12856), .A2(n9339), .ZN(n11177) );
  XNOR2_X1 U13548 ( .A(n11178), .B(n11177), .ZN(n11066) );
  AOI22_X1 U13549 ( .A1(n12757), .A2(n11061), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11062) );
  OAI21_X1 U13550 ( .B1(n11063), .B2(n12742), .A(n11062), .ZN(n11064) );
  AOI21_X1 U13551 ( .B1(n13156), .B2(n12747), .A(n11064), .ZN(n11065) );
  OAI21_X1 U13552 ( .B1(n11066), .B2(n12749), .A(n11065), .ZN(P2_U3213) );
  NAND2_X1 U13553 ( .A1(n11067), .A2(n11072), .ZN(n11068) );
  XNOR2_X1 U13554 ( .A(n11268), .B(n14725), .ZN(n11208) );
  XNOR2_X1 U13555 ( .A(n11208), .B(n12274), .ZN(n11070) );
  OAI211_X1 U13556 ( .C1(n11071), .C2(n11070), .A(n11211), .B(n14668), .ZN(
        n11075) );
  AND2_X1 U13557 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n14702) );
  OAI22_X1 U13558 ( .A1(n11974), .A2(n11072), .B1(n11236), .B2(n12000), .ZN(
        n11073) );
  AOI211_X1 U13559 ( .C1(n14725), .C2(n14675), .A(n14702), .B(n11073), .ZN(
        n11074) );
  OAI211_X1 U13560 ( .C1(n14741), .C2(n14678), .A(n11075), .B(n11074), .ZN(
        P3_U3157) );
  AOI21_X1 U13561 ( .B1(n11078), .B2(n11077), .A(n11076), .ZN(n11094) );
  OAI21_X1 U13562 ( .B1(n11081), .B2(n11080), .A(n11079), .ZN(n11092) );
  NAND2_X1 U13563 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n11083)
         );
  NAND2_X1 U13564 ( .A1(n14664), .A2(P3_ADDR_REG_14__SCAN_IN), .ZN(n11082) );
  OAI211_X1 U13565 ( .C1(n14719), .C2(n11084), .A(n11083), .B(n11082), .ZN(
        n11091) );
  OAI21_X1 U13566 ( .B1(n11087), .B2(n11086), .A(n11085), .ZN(n11089) );
  AND3_X1 U13567 ( .A1(n11089), .A2(n14713), .A3(n11088), .ZN(n11090) );
  AOI211_X1 U13568 ( .C1(n14703), .C2(n11092), .A(n11091), .B(n11090), .ZN(
        n11093) );
  OAI21_X1 U13569 ( .B1(n11094), .B2(n14708), .A(n11093), .ZN(P3_U3196) );
  INV_X1 U13570 ( .A(n11095), .ZN(n11096) );
  OAI222_X1 U13571 ( .A1(n11098), .A2(P3_U3151), .B1(n12661), .B2(n11097), 
        .C1(n12664), .C2(n11096), .ZN(P3_U3270) );
  AOI22_X1 U13572 ( .A1(n11100), .A2(n9889), .B1(n6452), .B2(n13344), .ZN(
        n11099) );
  XNOR2_X1 U13573 ( .A(n11099), .B(n11856), .ZN(n11123) );
  AOI22_X1 U13574 ( .A1(n11100), .A2(n6452), .B1(n11858), .B2(n13344), .ZN(
        n11124) );
  XNOR2_X1 U13575 ( .A(n11123), .B(n11124), .ZN(n11110) );
  INV_X1 U13576 ( .A(n11103), .ZN(n11106) );
  INV_X1 U13577 ( .A(n11104), .ZN(n11105) );
  NAND2_X1 U13578 ( .A1(n11106), .A2(n11105), .ZN(n11107) );
  INV_X1 U13579 ( .A(n11110), .ZN(n11109) );
  INV_X1 U13580 ( .A(n11136), .ZN(n11132) );
  AOI21_X1 U13581 ( .B1(n11110), .B2(n11108), .A(n11132), .ZN(n11117) );
  NAND2_X1 U13582 ( .A1(n14073), .A2(n13345), .ZN(n11112) );
  OAI211_X1 U13583 ( .C1(n13964), .C2(n13313), .A(n11112), .B(n11111), .ZN(
        n11114) );
  NOR2_X1 U13584 ( .A1(n14152), .A2(n13329), .ZN(n11113) );
  AOI211_X1 U13585 ( .C1(n11115), .C2(n13326), .A(n11114), .B(n11113), .ZN(
        n11116) );
  OAI21_X1 U13586 ( .B1(n11117), .B2(n14078), .A(n11116), .ZN(P1_U3236) );
  INV_X1 U13587 ( .A(n11118), .ZN(n11119) );
  INV_X1 U13588 ( .A(n11513), .ZN(n11121) );
  INV_X1 U13589 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11514) );
  OAI222_X1 U13590 ( .A1(n11119), .A2(P2_U3088), .B1(n13213), .B2(n11121), 
        .C1(n11514), .C2(n13210), .ZN(P2_U3303) );
  INV_X1 U13591 ( .A(n9234), .ZN(n11120) );
  OAI222_X1 U13592 ( .A1(n13833), .A2(n11122), .B1(n13837), .B2(n11121), .C1(
        n11120), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U13593 ( .A(n11123), .ZN(n11126) );
  INV_X1 U13594 ( .A(n11124), .ZN(n11125) );
  NOR2_X1 U13595 ( .A1(n11126), .A2(n11125), .ZN(n11134) );
  NAND2_X1 U13596 ( .A1(n11131), .A2(n9889), .ZN(n11128) );
  NAND2_X1 U13597 ( .A1(n6452), .A2(n13343), .ZN(n11127) );
  NAND2_X1 U13598 ( .A1(n11128), .A2(n11127), .ZN(n11129) );
  XNOR2_X1 U13599 ( .A(n11129), .B(n11813), .ZN(n11194) );
  NOR2_X1 U13600 ( .A1(n11815), .A2(n13964), .ZN(n11130) );
  AOI21_X1 U13601 ( .B1(n11131), .B2(n6452), .A(n11130), .ZN(n11195) );
  XNOR2_X1 U13602 ( .A(n11194), .B(n11195), .ZN(n11133) );
  OAI21_X1 U13603 ( .B1(n11132), .B2(n11134), .A(n11133), .ZN(n11137) );
  NOR2_X1 U13604 ( .A1(n11134), .A2(n11133), .ZN(n11135) );
  NAND3_X1 U13605 ( .A1(n11137), .A2(n13320), .A3(n11199), .ZN(n11144) );
  AOI21_X1 U13606 ( .B1(n14074), .B2(n13342), .A(n11138), .ZN(n11139) );
  OAI21_X1 U13607 ( .B1(n11140), .B2(n13267), .A(n11139), .ZN(n11141) );
  AOI21_X1 U13608 ( .B1(n11142), .B2(n13326), .A(n11141), .ZN(n11143) );
  OAI211_X1 U13609 ( .C1(n13957), .C2(n13329), .A(n11144), .B(n11143), .ZN(
        P1_U3224) );
  NAND2_X1 U13610 ( .A1(n11146), .A2(n11145), .ZN(n11148) );
  NAND2_X1 U13611 ( .A1(n11148), .A2(n11147), .ZN(n14084) );
  INV_X1 U13612 ( .A(n13340), .ZN(n11150) );
  NAND2_X1 U13613 ( .A1(n14089), .A2(n11150), .ZN(n11151) );
  INV_X1 U13614 ( .A(n11153), .ZN(n11158) );
  OAI21_X1 U13615 ( .B1(n6968), .B2(n11153), .A(n13524), .ZN(n14120) );
  OR2_X1 U13616 ( .A1(n13337), .A2(n14088), .ZN(n11154) );
  NAND2_X1 U13617 ( .A1(n14098), .A2(n14099), .ZN(n11157) );
  OR2_X1 U13618 ( .A1(n14089), .A2(n13340), .ZN(n11156) );
  XNOR2_X1 U13619 ( .A(n13505), .B(n11158), .ZN(n14123) );
  NAND2_X1 U13620 ( .A1(n14123), .A2(n14308), .ZN(n11167) );
  INV_X1 U13621 ( .A(n14089), .ZN(n14128) );
  INV_X1 U13622 ( .A(n14124), .ZN(n11160) );
  OAI21_X1 U13623 ( .B1(n11160), .B2(n13522), .A(n6482), .ZN(n14119) );
  INV_X1 U13624 ( .A(n14119), .ZN(n11165) );
  AOI22_X1 U13625 ( .A1(n13507), .A2(n6454), .B1(n14087), .B2(n13340), .ZN(
        n14118) );
  INV_X1 U13626 ( .A(n13281), .ZN(n11161) );
  OAI22_X1 U13627 ( .A1(n14322), .A2(n14118), .B1(n11161), .B2(n14093), .ZN(
        n11162) );
  AOI21_X1 U13628 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14322), .A(n11162), 
        .ZN(n11163) );
  OAI21_X1 U13629 ( .B1(n13522), .B2(n14298), .A(n11163), .ZN(n11164) );
  AOI21_X1 U13630 ( .B1(n11165), .B2(n13725), .A(n11164), .ZN(n11166) );
  OAI211_X1 U13631 ( .C1(n14120), .C2(n13705), .A(n11167), .B(n11166), .ZN(
        P1_U3276) );
  NAND2_X1 U13632 ( .A1(n11168), .A2(n11584), .ZN(n11172) );
  NOR2_X1 U13633 ( .A1(n11608), .A2(n11169), .ZN(n11170) );
  AOI21_X1 U13634 ( .B1(n14522), .B2(n11433), .A(n11170), .ZN(n11171) );
  XNOR2_X1 U13635 ( .A(n13151), .B(n11724), .ZN(n11174) );
  NAND2_X1 U13636 ( .A1(n12860), .A2(n9339), .ZN(n11173) );
  NAND2_X1 U13637 ( .A1(n11174), .A2(n11173), .ZN(n11689) );
  OAI21_X1 U13638 ( .B1(n11174), .B2(n11173), .A(n11689), .ZN(n11180) );
  OAI22_X1 U13639 ( .A1(n11178), .A2(n11177), .B1(n11176), .B2(n11175), .ZN(
        n11179) );
  NOR2_X1 U13640 ( .A1(n11179), .A2(n11180), .ZN(n11691) );
  AOI21_X1 U13641 ( .B1(n11180), .B2(n11179), .A(n11691), .ZN(n11193) );
  NOR2_X1 U13642 ( .A1(n12742), .A2(n13072), .ZN(n11191) );
  AND2_X1 U13643 ( .A1(n11182), .A2(n11181), .ZN(n11183) );
  OR2_X1 U13644 ( .A1(n11183), .A2(n11420), .ZN(n13054) );
  INV_X1 U13645 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n11186) );
  NAND2_X1 U13646 ( .A1(n11612), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U13647 ( .A1(n9864), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n11184) );
  OAI211_X1 U13648 ( .C1(n11616), .C2(n11186), .A(n11185), .B(n11184), .ZN(
        n11187) );
  INV_X1 U13649 ( .A(n11187), .ZN(n11188) );
  AND2_X1 U13650 ( .A1(n12856), .A2(n12754), .ZN(n11189) );
  AOI21_X1 U13651 ( .B1(n12863), .B2(n12824), .A(n11189), .ZN(n13068) );
  NAND2_X1 U13652 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n14523)
         );
  OAI21_X1 U13653 ( .B1(n12744), .B2(n13068), .A(n14523), .ZN(n11190) );
  AOI211_X1 U13654 ( .C1(n13151), .C2(n12747), .A(n11191), .B(n11190), .ZN(
        n11192) );
  OAI21_X1 U13655 ( .B1(n11193), .B2(n12749), .A(n11192), .ZN(P2_U3198) );
  INV_X1 U13656 ( .A(n11194), .ZN(n11197) );
  INV_X1 U13657 ( .A(n11195), .ZN(n11196) );
  NAND2_X1 U13658 ( .A1(n11197), .A2(n11196), .ZN(n11198) );
  NOR2_X1 U13659 ( .A1(n11815), .A2(n11200), .ZN(n11201) );
  AOI21_X1 U13660 ( .B1(n14145), .B2(n6452), .A(n11201), .ZN(n11740) );
  AOI22_X1 U13661 ( .A1(n14145), .A2(n9889), .B1(n6452), .B2(n13342), .ZN(
        n11202) );
  XNOR2_X1 U13662 ( .A(n11202), .B(n11856), .ZN(n11741) );
  XOR2_X1 U13663 ( .A(n11740), .B(n11741), .Z(n11738) );
  XNOR2_X1 U13664 ( .A(n11739), .B(n11738), .ZN(n11207) );
  NAND2_X1 U13665 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14204)
         );
  OAI21_X1 U13666 ( .B1(n13313), .B2(n13966), .A(n14204), .ZN(n11203) );
  AOI21_X1 U13667 ( .B1(n14073), .B2(n13343), .A(n11203), .ZN(n11204) );
  OAI21_X1 U13668 ( .B1(n14083), .B2(n13981), .A(n11204), .ZN(n11205) );
  AOI21_X1 U13669 ( .B1(n14075), .B2(n14145), .A(n11205), .ZN(n11206) );
  OAI21_X1 U13670 ( .B1(n11207), .B2(n14078), .A(n11206), .ZN(P1_U3234) );
  INV_X1 U13671 ( .A(n11208), .ZN(n11209) );
  NAND2_X1 U13672 ( .A1(n11209), .A2(n12274), .ZN(n11210) );
  XNOR2_X1 U13673 ( .A(n11268), .B(n11212), .ZN(n11239) );
  XNOR2_X1 U13674 ( .A(n11237), .B(n14729), .ZN(n11218) );
  AOI22_X1 U13675 ( .A1(n12003), .A2(n12274), .B1(n11212), .B2(n14675), .ZN(
        n11214) );
  OAI211_X1 U13676 ( .C1(n11985), .C2(n12000), .A(n11214), .B(n11213), .ZN(
        n11215) );
  AOI21_X1 U13677 ( .B1(n11977), .B2(n11216), .A(n11215), .ZN(n11217) );
  OAI21_X1 U13678 ( .B1(n11218), .B2(n12023), .A(n11217), .ZN(P3_U3176) );
  OAI211_X1 U13679 ( .C1(n11220), .C2(n12232), .A(n11219), .B(n14778), .ZN(
        n11222) );
  AOI22_X1 U13680 ( .A1(n11980), .A2(n14730), .B1(n14731), .B2(n14729), .ZN(
        n11221) );
  NAND2_X1 U13681 ( .A1(n11222), .A2(n11221), .ZN(n11229) );
  MUX2_X1 U13682 ( .A(n11229), .B(P3_REG0_REG_12__SCAN_IN), .S(n14849), .Z(
        n11225) );
  XNOR2_X1 U13683 ( .A(n11223), .B(n12232), .ZN(n11234) );
  OAI22_X1 U13684 ( .A1(n11234), .A2(n12622), .B1(n11226), .B2(n12635), .ZN(
        n11224) );
  OR2_X1 U13685 ( .A1(n11225), .A2(n11224), .ZN(P3_U3426) );
  MUX2_X1 U13686 ( .A(P3_REG1_REG_12__SCAN_IN), .B(n11229), .S(n14868), .Z(
        n11228) );
  OAI22_X1 U13687 ( .A1(n11234), .A2(n12540), .B1(n11226), .B2(n12548), .ZN(
        n11227) );
  OR2_X1 U13688 ( .A1(n11228), .A2(n11227), .ZN(P3_U3471) );
  INV_X1 U13689 ( .A(n11229), .ZN(n11230) );
  MUX2_X1 U13690 ( .A(n11230), .B(n7715), .S(n14793), .Z(n11233) );
  INV_X1 U13691 ( .A(n11937), .ZN(n11231) );
  AOI22_X1 U13692 ( .A1(n6433), .A2(n11941), .B1(n14772), .B2(n11231), .ZN(
        n11232) );
  OAI211_X1 U13693 ( .C1(n12493), .C2(n11234), .A(n11233), .B(n11232), .ZN(
        P3_U3221) );
  INV_X1 U13694 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n12038) );
  OAI222_X1 U13695 ( .A1(P2_U3088), .A2(n11235), .B1(n13213), .B2(n13824), 
        .C1(n12038), .C2(n13210), .ZN(P2_U3297) );
  INV_X1 U13696 ( .A(n11464), .ZN(n11870) );
  OAI222_X1 U13697 ( .A1(n11672), .A2(P2_U3088), .B1(n13213), .B2(n11870), 
        .C1(n11465), .C2(n13210), .ZN(P2_U3306) );
  INV_X1 U13698 ( .A(n11238), .ZN(n11240) );
  NAND2_X1 U13699 ( .A1(n11240), .A2(n11239), .ZN(n11241) );
  XNOR2_X1 U13700 ( .A(n11268), .B(n11941), .ZN(n11242) );
  XNOR2_X1 U13701 ( .A(n11242), .B(n12273), .ZN(n11936) );
  NAND2_X1 U13702 ( .A1(n11242), .A2(n11985), .ZN(n11243) );
  XNOR2_X1 U13703 ( .A(n12634), .B(n9067), .ZN(n11981) );
  INV_X1 U13704 ( .A(n11981), .ZN(n11245) );
  NAND2_X1 U13705 ( .A1(n11245), .A2(n11980), .ZN(n11246) );
  XNOR2_X1 U13706 ( .A(n12623), .B(n11268), .ZN(n11895) );
  INV_X1 U13707 ( .A(n11895), .ZN(n11247) );
  NAND2_X1 U13708 ( .A1(n11247), .A2(n11894), .ZN(n11248) );
  XNOR2_X1 U13709 ( .A(n12616), .B(n11268), .ZN(n12014) );
  XNOR2_X1 U13710 ( .A(n12154), .B(n11268), .ZN(n11952) );
  AND2_X1 U13711 ( .A1(n11952), .A2(n12433), .ZN(n11252) );
  INV_X1 U13712 ( .A(n11952), .ZN(n11250) );
  NAND2_X1 U13713 ( .A1(n11250), .A2(n12018), .ZN(n11251) );
  XNOR2_X1 U13714 ( .A(n11969), .B(n11268), .ZN(n11253) );
  XNOR2_X1 U13715 ( .A(n11253), .B(n12419), .ZN(n11961) );
  XNOR2_X1 U13716 ( .A(n12427), .B(n11268), .ZN(n11254) );
  XNOR2_X1 U13717 ( .A(n11254), .B(n12434), .ZN(n11998) );
  INV_X1 U13718 ( .A(n11254), .ZN(n11255) );
  NAND2_X1 U13719 ( .A1(n11255), .A2(n12434), .ZN(n11256) );
  NAND2_X1 U13720 ( .A1(n11997), .A2(n11256), .ZN(n11912) );
  XNOR2_X1 U13721 ( .A(n12593), .B(n11268), .ZN(n11257) );
  XNOR2_X1 U13722 ( .A(n11257), .B(n12420), .ZN(n11911) );
  NAND2_X1 U13723 ( .A1(n11912), .A2(n11911), .ZN(n11910) );
  NAND2_X1 U13724 ( .A1(n11257), .A2(n12270), .ZN(n11258) );
  XNOR2_X1 U13725 ( .A(n12400), .B(n11268), .ZN(n11259) );
  XNOR2_X1 U13726 ( .A(n11259), .B(n12269), .ZN(n11971) );
  INV_X1 U13727 ( .A(n11259), .ZN(n11260) );
  NAND2_X1 U13728 ( .A1(n11260), .A2(n12269), .ZN(n11261) );
  XNOR2_X1 U13729 ( .A(n12583), .B(n11268), .ZN(n11262) );
  XNOR2_X1 U13730 ( .A(n11262), .B(n12268), .ZN(n11928) );
  INV_X1 U13731 ( .A(n11262), .ZN(n11263) );
  NAND2_X1 U13732 ( .A1(n11263), .A2(n12396), .ZN(n11264) );
  XNOR2_X1 U13733 ( .A(n12578), .B(n9067), .ZN(n11873) );
  INV_X1 U13734 ( .A(n11873), .ZN(n11875) );
  AND2_X1 U13735 ( .A1(n11884), .A2(n11875), .ZN(n11265) );
  XNOR2_X1 U13736 ( .A(n12572), .B(n11268), .ZN(n11877) );
  XNOR2_X1 U13737 ( .A(n12569), .B(n11268), .ZN(n11881) );
  XNOR2_X1 U13738 ( .A(n11881), .B(n12362), .ZN(n11269) );
  XNOR2_X1 U13739 ( .A(n11270), .B(n11269), .ZN(n11275) );
  OAI22_X1 U13740 ( .A1(n12178), .A2(n14762), .B1(n12189), .B2(n14760), .ZN(
        n12347) );
  AOI22_X1 U13741 ( .A1(n12347), .A2(n12019), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11271) );
  OAI21_X1 U13742 ( .B1(n12352), .B2(n14678), .A(n11271), .ZN(n11272) );
  AOI21_X1 U13743 ( .B1(n11273), .B2(n14675), .A(n11272), .ZN(n11274) );
  OAI21_X1 U13744 ( .B1(n11275), .B2(n12023), .A(n11274), .ZN(P3_U3169) );
  INV_X1 U13745 ( .A(n11527), .ZN(n13212) );
  OAI222_X1 U13746 ( .A1(n13833), .A2(n11276), .B1(n13837), .B2(n13212), .C1(
        n9233), .C2(P1_U3086), .ZN(P1_U3330) );
  XNOR2_X1 U13747 ( .A(n8371), .B(n11277), .ZN(n11486) );
  INV_X1 U13748 ( .A(n11486), .ZN(n11278) );
  OAI222_X1 U13749 ( .A1(n13210), .A2(n11487), .B1(n13213), .B2(n11278), .C1(
        P2_U3088), .C2(n9294), .ZN(P2_U3305) );
  INV_X1 U13750 ( .A(n11279), .ZN(n11280) );
  OAI222_X1 U13751 ( .A1(n11282), .A2(P3_U3151), .B1(n12661), .B2(n11281), 
        .C1(n12657), .C2(n11280), .ZN(P3_U3271) );
  NOR2_X1 U13752 ( .A1(n9331), .A2(n12819), .ZN(n11283) );
  NOR2_X1 U13753 ( .A1(n11284), .A2(n11638), .ZN(n11285) );
  NOR2_X1 U13754 ( .A1(n11301), .A2(n11285), .ZN(n11286) );
  NAND2_X1 U13755 ( .A1(n11289), .A2(n11286), .ZN(n11287) );
  NAND2_X1 U13756 ( .A1(n11301), .A2(n11294), .ZN(n11292) );
  NAND2_X1 U13757 ( .A1(n11293), .A2(n6450), .ZN(n11291) );
  NAND2_X1 U13758 ( .A1(n11293), .A2(n6441), .ZN(n11296) );
  NAND2_X1 U13759 ( .A1(n6449), .A2(n11294), .ZN(n11295) );
  NAND2_X1 U13760 ( .A1(n11296), .A2(n11295), .ZN(n11297) );
  NAND2_X1 U13761 ( .A1(n6439), .A2(n12782), .ZN(n11300) );
  NAND2_X1 U13762 ( .A1(n6451), .A2(n9363), .ZN(n11299) );
  NAND2_X1 U13763 ( .A1(n11307), .A2(n11308), .ZN(n11306) );
  INV_X1 U13764 ( .A(n11307), .ZN(n11310) );
  INV_X1 U13765 ( .A(n11308), .ZN(n11309) );
  NAND2_X1 U13766 ( .A1(n11310), .A2(n11309), .ZN(n11311) );
  NAND2_X1 U13767 ( .A1(n12781), .A2(n6451), .ZN(n11313) );
  NAND2_X1 U13768 ( .A1(n14579), .A2(n6438), .ZN(n11312) );
  NAND2_X1 U13769 ( .A1(n11313), .A2(n11312), .ZN(n11318) );
  AOI22_X1 U13770 ( .A1(n12781), .A2(n6441), .B1(n14579), .B2(n6450), .ZN(
        n11314) );
  INV_X1 U13771 ( .A(n11314), .ZN(n11315) );
  NAND2_X1 U13772 ( .A1(n11316), .A2(n11315), .ZN(n11322) );
  INV_X1 U13773 ( .A(n11317), .ZN(n11320) );
  NAND2_X1 U13774 ( .A1(n11320), .A2(n11319), .ZN(n11321) );
  NAND2_X1 U13775 ( .A1(n11325), .A2(n6451), .ZN(n11324) );
  NAND2_X1 U13776 ( .A1(n12780), .A2(n6440), .ZN(n11323) );
  NAND2_X1 U13777 ( .A1(n11325), .A2(n6439), .ZN(n11327) );
  NAND2_X1 U13778 ( .A1(n12780), .A2(n6449), .ZN(n11326) );
  NAND2_X1 U13779 ( .A1(n11327), .A2(n11326), .ZN(n11328) );
  NAND2_X1 U13780 ( .A1(n11331), .A2(n6438), .ZN(n11330) );
  NAND2_X1 U13781 ( .A1(n12779), .A2(n6451), .ZN(n11329) );
  NAND2_X1 U13782 ( .A1(n11330), .A2(n11329), .ZN(n11333) );
  AOI22_X1 U13783 ( .A1(n11331), .A2(n6450), .B1(n6440), .B2(n12779), .ZN(
        n11332) );
  NAND2_X1 U13784 ( .A1(n14601), .A2(n6442), .ZN(n11336) );
  NAND2_X1 U13785 ( .A1(n12778), .A2(n6444), .ZN(n11335) );
  NAND2_X1 U13786 ( .A1(n11336), .A2(n11335), .ZN(n11342) );
  NAND2_X1 U13787 ( .A1(n14601), .A2(n6440), .ZN(n11337) );
  OAI21_X1 U13788 ( .B1(n6441), .B2(n11338), .A(n11337), .ZN(n11339) );
  NAND2_X1 U13789 ( .A1(n11340), .A2(n11339), .ZN(n11344) );
  NAND2_X1 U13790 ( .A1(n11347), .A2(n6439), .ZN(n11346) );
  NAND2_X1 U13791 ( .A1(n12777), .A2(n6450), .ZN(n11345) );
  AOI22_X1 U13792 ( .A1(n11347), .A2(n6449), .B1(n6438), .B2(n12777), .ZN(
        n11348) );
  NAND2_X1 U13793 ( .A1(n14617), .A2(n6442), .ZN(n11351) );
  NAND2_X1 U13794 ( .A1(n12776), .A2(n6443), .ZN(n11350) );
  NAND2_X1 U13795 ( .A1(n11351), .A2(n11350), .ZN(n11353) );
  AOI22_X1 U13796 ( .A1(n14617), .A2(n6444), .B1(n6451), .B2(n12776), .ZN(
        n11352) );
  NAND2_X1 U13797 ( .A1(n11356), .A2(n6446), .ZN(n11355) );
  NAND2_X1 U13798 ( .A1(n12775), .A2(n6450), .ZN(n11354) );
  NAND2_X1 U13799 ( .A1(n11355), .A2(n11354), .ZN(n11362) );
  NAND2_X1 U13800 ( .A1(n11361), .A2(n11362), .ZN(n11360) );
  NAND2_X1 U13801 ( .A1(n11356), .A2(n6442), .ZN(n11357) );
  OAI21_X1 U13802 ( .B1(n11358), .B2(n6450), .A(n11357), .ZN(n11359) );
  NAND2_X1 U13803 ( .A1(n11360), .A2(n11359), .ZN(n11366) );
  NAND2_X1 U13804 ( .A1(n11364), .A2(n11363), .ZN(n11365) );
  NAND2_X1 U13805 ( .A1(n14638), .A2(n6442), .ZN(n11368) );
  NAND2_X1 U13806 ( .A1(n12774), .A2(n6447), .ZN(n11367) );
  NAND2_X1 U13807 ( .A1(n11368), .A2(n11367), .ZN(n11370) );
  AOI22_X1 U13808 ( .A1(n14638), .A2(n6447), .B1(n6451), .B2(n12774), .ZN(
        n11369) );
  NAND2_X1 U13809 ( .A1(n11374), .A2(n6445), .ZN(n11373) );
  NAND2_X1 U13810 ( .A1(n12773), .A2(n6449), .ZN(n11372) );
  NAND2_X1 U13811 ( .A1(n11373), .A2(n11372), .ZN(n11378) );
  NAND2_X1 U13812 ( .A1(n11374), .A2(n6451), .ZN(n11375) );
  OAI21_X1 U13813 ( .B1(n11376), .B2(n6449), .A(n11375), .ZN(n11377) );
  NAND2_X1 U13814 ( .A1(n13172), .A2(n6451), .ZN(n11381) );
  NAND2_X1 U13815 ( .A1(n12772), .A2(n6447), .ZN(n11380) );
  NAND2_X1 U13816 ( .A1(n11381), .A2(n11380), .ZN(n11384) );
  AOI22_X1 U13817 ( .A1(n13172), .A2(n6447), .B1(n6442), .B2(n12772), .ZN(
        n11382) );
  INV_X1 U13818 ( .A(n11383), .ZN(n11386) );
  NAND2_X1 U13819 ( .A1(n13167), .A2(n6447), .ZN(n11388) );
  NAND2_X1 U13820 ( .A1(n12771), .A2(n6449), .ZN(n11387) );
  NAND2_X1 U13821 ( .A1(n13167), .A2(n6450), .ZN(n11389) );
  OAI21_X1 U13822 ( .B1(n11390), .B2(n6449), .A(n11389), .ZN(n11391) );
  NAND2_X1 U13823 ( .A1(n11394), .A2(n6449), .ZN(n11393) );
  NAND2_X1 U13824 ( .A1(n12770), .A2(n6447), .ZN(n11392) );
  NAND2_X1 U13825 ( .A1(n11393), .A2(n11392), .ZN(n11396) );
  AOI22_X1 U13826 ( .A1(n11394), .A2(n6446), .B1(n6442), .B2(n12770), .ZN(
        n11395) );
  NAND2_X1 U13827 ( .A1(n13156), .A2(n6447), .ZN(n11399) );
  NAND2_X1 U13828 ( .A1(n12856), .A2(n6450), .ZN(n11398) );
  NAND2_X1 U13829 ( .A1(n11399), .A2(n11398), .ZN(n11401) );
  AOI22_X1 U13830 ( .A1(n13156), .A2(n6451), .B1(n6447), .B2(n12856), .ZN(
        n11400) );
  NAND2_X1 U13831 ( .A1(n13151), .A2(n6451), .ZN(n11403) );
  NAND2_X1 U13832 ( .A1(n12860), .A2(n6447), .ZN(n11402) );
  NAND2_X1 U13833 ( .A1(n11403), .A2(n11402), .ZN(n11407) );
  NAND2_X1 U13834 ( .A1(n13151), .A2(n6445), .ZN(n11405) );
  NAND2_X1 U13835 ( .A1(n12860), .A2(n6450), .ZN(n11404) );
  NAND2_X1 U13836 ( .A1(n11408), .A2(n11584), .ZN(n11410) );
  AOI22_X1 U13837 ( .A1(n11434), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n11433), 
        .B2(n14536), .ZN(n11409) );
  NAND2_X1 U13838 ( .A1(n13146), .A2(n6446), .ZN(n11412) );
  NAND2_X1 U13839 ( .A1(n12863), .A2(n6449), .ZN(n11411) );
  NAND2_X1 U13840 ( .A1(n11412), .A2(n11411), .ZN(n11414) );
  AOI22_X1 U13841 ( .A1(n13146), .A2(n6451), .B1(n6445), .B2(n12863), .ZN(
        n11413) );
  NAND2_X1 U13842 ( .A1(n11417), .A2(n11584), .ZN(n11419) );
  INV_X1 U13843 ( .A(n12809), .ZN(n12790) );
  AOI22_X1 U13844 ( .A1(n11434), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n11433), 
        .B2(n12790), .ZN(n11418) );
  NAND2_X1 U13845 ( .A1(n13141), .A2(n6442), .ZN(n11427) );
  NOR2_X1 U13846 ( .A1(n11420), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11421) );
  OR2_X1 U13847 ( .A1(n11437), .A2(n11421), .ZN(n13037) );
  INV_X1 U13848 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n12799) );
  NAND2_X1 U13849 ( .A1(n11612), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n11423) );
  NAND2_X1 U13850 ( .A1(n9864), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n11422) );
  OAI211_X1 U13851 ( .C1(n11616), .C2(n12799), .A(n11423), .B(n11422), .ZN(
        n11424) );
  INV_X1 U13852 ( .A(n11424), .ZN(n11425) );
  OAI21_X1 U13853 ( .B1(n13037), .B2(n11459), .A(n11425), .ZN(n12864) );
  NAND2_X1 U13854 ( .A1(n12864), .A2(n6446), .ZN(n11426) );
  NAND2_X1 U13855 ( .A1(n11427), .A2(n11426), .ZN(n11430) );
  INV_X1 U13856 ( .A(n12864), .ZN(n12837) );
  NAND2_X1 U13857 ( .A1(n13141), .A2(n6445), .ZN(n11428) );
  OAI21_X1 U13858 ( .B1(n6447), .B2(n12837), .A(n11428), .ZN(n11429) );
  NAND2_X1 U13859 ( .A1(n11432), .A2(n11584), .ZN(n11436) );
  AOI22_X1 U13860 ( .A1(n11434), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n11680), 
        .B2(n11433), .ZN(n11435) );
  NAND2_X1 U13861 ( .A1(n13136), .A2(n6446), .ZN(n11445) );
  NOR2_X1 U13862 ( .A1(n11437), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n11438) );
  OR2_X1 U13863 ( .A1(n11452), .A2(n11438), .ZN(n13023) );
  INV_X1 U13864 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U13865 ( .A1(n11612), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11440) );
  NAND2_X1 U13866 ( .A1(n9864), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n11439) );
  OAI211_X1 U13867 ( .C1(n11616), .C2(n11441), .A(n11440), .B(n11439), .ZN(
        n11442) );
  INV_X1 U13868 ( .A(n11442), .ZN(n11443) );
  NAND2_X1 U13869 ( .A1(n12867), .A2(n6442), .ZN(n11444) );
  AOI22_X1 U13870 ( .A1(n13136), .A2(n6449), .B1(n6447), .B2(n12867), .ZN(
        n11446) );
  NAND2_X1 U13871 ( .A1(n11448), .A2(n11584), .ZN(n11451) );
  OR2_X1 U13872 ( .A1(n11608), .A2(n11449), .ZN(n11450) );
  NAND2_X1 U13873 ( .A1(n13131), .A2(n6450), .ZN(n11461) );
  NOR2_X1 U13874 ( .A1(n11452), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n11453) );
  OR2_X1 U13875 ( .A1(n11468), .A2(n11453), .ZN(n13008) );
  INV_X1 U13876 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n11456) );
  NAND2_X1 U13877 ( .A1(n11612), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n11455) );
  NAND2_X1 U13878 ( .A1(n9864), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11454) );
  OAI211_X1 U13879 ( .C1(n11616), .C2(n11456), .A(n11455), .B(n11454), .ZN(
        n11457) );
  INV_X1 U13880 ( .A(n11457), .ZN(n11458) );
  NAND2_X1 U13881 ( .A1(n12869), .A2(n6446), .ZN(n11460) );
  INV_X1 U13882 ( .A(n12869), .ZN(n12839) );
  NAND2_X1 U13883 ( .A1(n13131), .A2(n6447), .ZN(n11462) );
  OAI21_X1 U13884 ( .B1(n6445), .B2(n12839), .A(n11462), .ZN(n11463) );
  NAND2_X1 U13885 ( .A1(n11464), .A2(n11584), .ZN(n11467) );
  OR2_X1 U13886 ( .A1(n11608), .A2(n11465), .ZN(n11466) );
  NAND2_X1 U13887 ( .A1(n13126), .A2(n6447), .ZN(n11476) );
  OR2_X1 U13888 ( .A1(n11468), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11469) );
  AND2_X1 U13889 ( .A1(n11469), .A2(n11490), .ZN(n12996) );
  NAND2_X1 U13890 ( .A1(n12996), .A2(n11590), .ZN(n11474) );
  INV_X1 U13891 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n14959) );
  NAND2_X1 U13892 ( .A1(n11612), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n11471) );
  NAND2_X1 U13893 ( .A1(n9864), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11470) );
  OAI211_X1 U13894 ( .C1(n11616), .C2(n14959), .A(n11471), .B(n11470), .ZN(
        n11472) );
  INV_X1 U13895 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U13896 ( .A1(n11474), .A2(n11473), .ZN(n12872) );
  NAND2_X1 U13897 ( .A1(n12872), .A2(n6442), .ZN(n11475) );
  NAND2_X1 U13898 ( .A1(n11476), .A2(n11475), .ZN(n11481) );
  AOI22_X1 U13899 ( .A1(n13126), .A2(n6449), .B1(n6445), .B2(n12872), .ZN(
        n11477) );
  INV_X1 U13900 ( .A(n11477), .ZN(n11478) );
  NAND2_X1 U13901 ( .A1(n11479), .A2(n11478), .ZN(n11485) );
  NAND2_X1 U13902 ( .A1(n11483), .A2(n11482), .ZN(n11484) );
  NAND2_X1 U13903 ( .A1(n11486), .A2(n11584), .ZN(n11489) );
  OR2_X1 U13904 ( .A1(n11608), .A2(n11487), .ZN(n11488) );
  NAND2_X1 U13905 ( .A1(n9864), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11494) );
  NAND2_X1 U13906 ( .A1(n11591), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n11493) );
  INV_X1 U13907 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12736) );
  AOI21_X1 U13908 ( .B1(n12736), .B2(n11490), .A(n11503), .ZN(n12979) );
  NAND2_X1 U13909 ( .A1(n11590), .A2(n12979), .ZN(n11492) );
  NAND2_X1 U13910 ( .A1(n11612), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n11491) );
  OAI22_X1 U13911 ( .A1(n12981), .A2(n6447), .B1(n11495), .B2(n6450), .ZN(
        n11497) );
  INV_X1 U13912 ( .A(n11497), .ZN(n11498) );
  AOI22_X1 U13913 ( .A1(n13121), .A2(n6438), .B1(n6451), .B2(n12874), .ZN(
        n11496) );
  NAND2_X1 U13914 ( .A1(n11499), .A2(n11584), .ZN(n11502) );
  OR2_X1 U13915 ( .A1(n11608), .A2(n11500), .ZN(n11501) );
  NAND2_X1 U13916 ( .A1(n9864), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11507) );
  NAND2_X1 U13917 ( .A1(n11591), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U13918 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(n11503), .ZN(n11517) );
  OAI21_X1 U13919 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(n11503), .A(n11517), 
        .ZN(n12966) );
  INV_X1 U13920 ( .A(n12966), .ZN(n12679) );
  NAND2_X1 U13921 ( .A1(n11590), .A2(n12679), .ZN(n11505) );
  NAND2_X1 U13922 ( .A1(n11612), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n11504) );
  NAND4_X1 U13923 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n12877) );
  AOI22_X1 U13924 ( .A1(n13116), .A2(n6441), .B1(n6442), .B2(n12877), .ZN(
        n11509) );
  NAND2_X1 U13925 ( .A1(n11513), .A2(n11584), .ZN(n11516) );
  OR2_X1 U13926 ( .A1(n11608), .A2(n11514), .ZN(n11515) );
  NAND2_X1 U13927 ( .A1(n9864), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n11523) );
  NAND2_X1 U13928 ( .A1(n11612), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11522) );
  INV_X1 U13929 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12718) );
  NAND2_X1 U13930 ( .A1(n12718), .A2(n11517), .ZN(n11519) );
  INV_X1 U13931 ( .A(n11517), .ZN(n11518) );
  AND2_X1 U13932 ( .A1(n11519), .A2(n11543), .ZN(n12954) );
  NAND2_X1 U13933 ( .A1(n11590), .A2(n12954), .ZN(n11521) );
  NAND2_X1 U13934 ( .A1(n11591), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11520) );
  OAI22_X1 U13935 ( .A1(n13110), .A2(n6439), .B1(n12701), .B2(n6450), .ZN(
        n11525) );
  AOI22_X1 U13936 ( .A1(n12879), .A2(n6440), .B1(n6451), .B2(n12878), .ZN(
        n11524) );
  NAND2_X1 U13937 ( .A1(n11527), .A2(n11584), .ZN(n11529) );
  OR2_X1 U13938 ( .A1(n11608), .A2(n13211), .ZN(n11528) );
  NAND2_X2 U13939 ( .A1(n11529), .A2(n11528), .ZN(n13105) );
  NAND2_X1 U13940 ( .A1(n9864), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U13941 ( .A1(n11591), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11532) );
  XNOR2_X1 U13942 ( .A(n11543), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n12934) );
  NAND2_X1 U13943 ( .A1(n11590), .A2(n12934), .ZN(n11531) );
  NAND2_X1 U13944 ( .A1(n11612), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U13945 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n12880) );
  AOI22_X1 U13946 ( .A1(n13105), .A2(n6447), .B1(n6450), .B2(n12880), .ZN(
        n11535) );
  INV_X1 U13947 ( .A(n13105), .ZN(n12936) );
  INV_X1 U13948 ( .A(n12880), .ZN(n12843) );
  OAI22_X1 U13949 ( .A1(n12936), .A2(n6447), .B1(n12843), .B2(n6442), .ZN(
        n11534) );
  NAND2_X1 U13950 ( .A1(n13208), .A2(n11584), .ZN(n11538) );
  OR2_X1 U13951 ( .A1(n11608), .A2(n6922), .ZN(n11537) );
  NAND2_X1 U13952 ( .A1(n11591), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U13953 ( .A1(n9864), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11547) );
  INV_X1 U13954 ( .A(n11543), .ZN(n11540) );
  AND2_X1 U13955 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n11539) );
  NAND2_X1 U13956 ( .A1(n11540), .A2(n11539), .ZN(n11587) );
  INV_X1 U13957 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n11542) );
  INV_X1 U13958 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n11541) );
  OAI21_X1 U13959 ( .B1(n11543), .B2(n11542), .A(n11541), .ZN(n11544) );
  AND2_X1 U13960 ( .A1(n11587), .A2(n11544), .ZN(n12922) );
  NAND2_X1 U13961 ( .A1(n11590), .A2(n12922), .ZN(n11546) );
  NAND2_X1 U13962 ( .A1(n11612), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n11545) );
  AOI22_X1 U13963 ( .A1(n13100), .A2(n6442), .B1(n6445), .B2(n12882), .ZN(
        n11597) );
  OAI22_X1 U13964 ( .A1(n12924), .A2(n6451), .B1(n6447), .B2(n12881), .ZN(
        n11596) );
  OR2_X1 U13965 ( .A1(n11608), .A2(n11552), .ZN(n11553) );
  NAND2_X1 U13966 ( .A1(n11591), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n11563) );
  NAND2_X1 U13967 ( .A1(n9864), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n11562) );
  INV_X1 U13968 ( .A(n11587), .ZN(n11555) );
  INV_X1 U13969 ( .A(n12853), .ZN(n11559) );
  INV_X1 U13970 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11557) );
  NAND2_X1 U13971 ( .A1(n11589), .A2(n11557), .ZN(n11558) );
  NAND2_X1 U13972 ( .A1(n11590), .A2(n11732), .ZN(n11561) );
  NAND2_X1 U13973 ( .A1(n11612), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U13974 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n12884) );
  AND2_X1 U13975 ( .A1(n12884), .A2(n6444), .ZN(n11564) );
  AOI21_X1 U13976 ( .B1(n7078), .B2(n6449), .A(n11564), .ZN(n11627) );
  NAND2_X1 U13977 ( .A1(n7078), .A2(n6445), .ZN(n11566) );
  NAND2_X1 U13978 ( .A1(n12884), .A2(n6449), .ZN(n11565) );
  NAND2_X1 U13979 ( .A1(n11566), .A2(n11565), .ZN(n11625) );
  NAND2_X1 U13980 ( .A1(n11567), .A2(n11584), .ZN(n11569) );
  INV_X1 U13981 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12029) );
  OR2_X1 U13982 ( .A1(n11608), .A2(n12029), .ZN(n11568) );
  INV_X1 U13983 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n11572) );
  NAND2_X1 U13984 ( .A1(n11591), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n11571) );
  NAND2_X1 U13985 ( .A1(n11612), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n11570) );
  OAI211_X1 U13986 ( .C1(n11573), .C2(n11572), .A(n11571), .B(n11570), .ZN(
        n12766) );
  NAND2_X1 U13987 ( .A1(n11605), .A2(n12766), .ZN(n11574) );
  NAND2_X1 U13988 ( .A1(n13200), .A2(n11584), .ZN(n11576) );
  OR2_X1 U13989 ( .A1(n11608), .A2(n14963), .ZN(n11575) );
  NAND2_X1 U13990 ( .A1(n9864), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11580) );
  NAND2_X1 U13991 ( .A1(n11590), .A2(n12853), .ZN(n11579) );
  NAND2_X1 U13992 ( .A1(n11591), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11578) );
  NAND2_X1 U13993 ( .A1(n11612), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n11577) );
  NAND4_X1 U13994 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n12768) );
  AND2_X1 U13995 ( .A1(n12768), .A2(n6450), .ZN(n11581) );
  AOI21_X1 U13996 ( .B1(n13088), .B2(n6445), .A(n11581), .ZN(n11620) );
  NAND2_X1 U13997 ( .A1(n13088), .A2(n6451), .ZN(n11583) );
  NAND2_X1 U13998 ( .A1(n12768), .A2(n6446), .ZN(n11582) );
  NAND2_X1 U13999 ( .A1(n11583), .A2(n11582), .ZN(n11619) );
  NAND2_X1 U14000 ( .A1(n11620), .A2(n11619), .ZN(n11626) );
  OAI211_X1 U14001 ( .C1(n11627), .C2(n11625), .A(n11642), .B(n11626), .ZN(
        n11604) );
  OR2_X1 U14002 ( .A1(n11608), .A2(n13205), .ZN(n11585) );
  NAND2_X1 U14003 ( .A1(n9864), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n11595) );
  NAND2_X1 U14004 ( .A1(n11612), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n11594) );
  INV_X1 U14005 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12670) );
  NAND2_X1 U14006 ( .A1(n11587), .A2(n12670), .ZN(n11588) );
  NAND2_X1 U14007 ( .A1(n11590), .A2(n12909), .ZN(n11593) );
  NAND2_X1 U14008 ( .A1(n11591), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11592) );
  OAI22_X1 U14009 ( .A1(n12911), .A2(n6450), .B1(n6446), .B2(n12883), .ZN(
        n11600) );
  AOI22_X1 U14010 ( .A1(n13096), .A2(n6442), .B1(n6447), .B2(n12769), .ZN(
        n11601) );
  OAI22_X1 U14011 ( .A1(n11600), .A2(n11601), .B1(n11597), .B2(n11596), .ZN(
        n11598) );
  INV_X1 U14012 ( .A(n11600), .ZN(n11603) );
  INV_X1 U14013 ( .A(n11601), .ZN(n11602) );
  NOR3_X1 U14014 ( .A1(n11604), .A2(n11603), .A3(n11602), .ZN(n11628) );
  NOR2_X1 U14015 ( .A1(n13083), .A2(n6445), .ZN(n11606) );
  OR2_X1 U14016 ( .A1(n13824), .A2(n11607), .ZN(n11610) );
  OR2_X1 U14017 ( .A1(n11608), .A2(n12038), .ZN(n11609) );
  INV_X1 U14018 ( .A(n12766), .ZN(n12825) );
  NOR2_X1 U14019 ( .A1(n12825), .A2(n6445), .ZN(n11634) );
  OAI211_X1 U14020 ( .C1(n11611), .C2(n11646), .A(n9330), .B(n11639), .ZN(
        n11617) );
  INV_X1 U14021 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U14022 ( .A1(n9864), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11614) );
  NAND2_X1 U14023 ( .A1(n11612), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11613) );
  OAI211_X1 U14024 ( .C1(n11616), .C2(n11615), .A(n11614), .B(n11613), .ZN(
        n12767) );
  OAI21_X1 U14025 ( .B1(n11634), .B2(n11617), .A(n12767), .ZN(n11618) );
  OAI21_X1 U14026 ( .B1(n13086), .B2(n6449), .A(n11618), .ZN(n11630) );
  AOI22_X1 U14027 ( .A1(n7079), .A2(n6451), .B1(n6446), .B2(n12767), .ZN(
        n11629) );
  INV_X1 U14028 ( .A(n11619), .ZN(n11622) );
  INV_X1 U14029 ( .A(n11620), .ZN(n11621) );
  AOI22_X1 U14030 ( .A1(n11630), .A2(n11629), .B1(n11622), .B2(n11621), .ZN(
        n11623) );
  INV_X1 U14031 ( .A(n11629), .ZN(n11632) );
  INV_X1 U14032 ( .A(n11630), .ZN(n11631) );
  NAND2_X1 U14033 ( .A1(n11632), .A2(n11631), .ZN(n11633) );
  INV_X1 U14034 ( .A(n11634), .ZN(n11636) );
  OAI211_X1 U14035 ( .C1(n13083), .C2(n6450), .A(n11636), .B(n11635), .ZN(
        n11637) );
  INV_X1 U14036 ( .A(n11638), .ZN(n11641) );
  OAI21_X1 U14037 ( .B1(n11672), .B2(n11680), .A(n11639), .ZN(n11640) );
  AOI21_X1 U14038 ( .B1(n11641), .B2(n9294), .A(n11640), .ZN(n11683) );
  INV_X1 U14039 ( .A(n11642), .ZN(n11670) );
  INV_X1 U14040 ( .A(n12768), .ZN(n11643) );
  INV_X1 U14041 ( .A(n12884), .ZN(n12849) );
  NAND2_X1 U14042 ( .A1(n7078), .A2(n12849), .ZN(n11644) );
  XNOR2_X1 U14043 ( .A(n13105), .B(n12843), .ZN(n12938) );
  XNOR2_X1 U14044 ( .A(n13100), .B(n12881), .ZN(n12926) );
  INV_X1 U14045 ( .A(n12872), .ZN(n12840) );
  XNOR2_X1 U14046 ( .A(n13131), .B(n12869), .ZN(n13012) );
  XNOR2_X1 U14047 ( .A(n13146), .B(n12863), .ZN(n12862) );
  OAI21_X1 U14048 ( .B1(n11289), .B2(n14545), .A(n11645), .ZN(n14567) );
  NAND4_X1 U14049 ( .A1(n6597), .A2(n11650), .A3(n11649), .A4(n11648), .ZN(
        n11651) );
  NOR2_X1 U14050 ( .A1(n11652), .A2(n11651), .ZN(n11655) );
  NAND4_X1 U14051 ( .A1(n7463), .A2(n11655), .A3(n11654), .A4(n11653), .ZN(
        n11656) );
  OR4_X1 U14052 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n11660) );
  NOR2_X1 U14053 ( .A1(n11661), .A2(n11660), .ZN(n11663) );
  NAND4_X1 U14054 ( .A1(n12862), .A2(n11663), .A3(n13066), .A4(n11662), .ZN(
        n11664) );
  NOR2_X1 U14055 ( .A1(n11664), .A2(n12832), .ZN(n11665) );
  XNOR2_X1 U14056 ( .A(n13136), .B(n12867), .ZN(n13026) );
  XNOR2_X1 U14057 ( .A(n13141), .B(n12864), .ZN(n13031) );
  NAND4_X1 U14058 ( .A1(n13012), .A2(n11665), .A3(n13026), .A4(n13031), .ZN(
        n11666) );
  NOR2_X1 U14059 ( .A1(n12999), .A2(n11666), .ZN(n11667) );
  XNOR2_X1 U14060 ( .A(n13116), .B(n12877), .ZN(n12961) );
  XNOR2_X1 U14061 ( .A(n13121), .B(n12874), .ZN(n12982) );
  NAND4_X1 U14062 ( .A1(n12950), .A2(n11667), .A3(n12961), .A4(n12982), .ZN(
        n11668) );
  INV_X1 U14063 ( .A(n12767), .ZN(n12847) );
  OAI21_X1 U14064 ( .B1(n7079), .B2(n12847), .A(n12912), .ZN(n11669) );
  NAND2_X1 U14065 ( .A1(n11672), .A2(n11680), .ZN(n11674) );
  MUX2_X1 U14066 ( .A(n11672), .B(n9294), .S(n11671), .Z(n11673) );
  NAND2_X1 U14067 ( .A1(n7079), .A2(n12847), .ZN(n11676) );
  NAND3_X1 U14068 ( .A1(n11681), .A2(n11680), .A3(n11676), .ZN(n11679) );
  INV_X1 U14069 ( .A(n11676), .ZN(n11677) );
  AOI211_X1 U14070 ( .C1(n11677), .C2(n12819), .A(n9330), .B(n14546), .ZN(
        n11678) );
  OAI211_X1 U14071 ( .C1(n11681), .C2(n11680), .A(n11679), .B(n11678), .ZN(
        n11682) );
  NAND4_X1 U14072 ( .A1(n14566), .A2(n12754), .A3(n12822), .A4(n11685), .ZN(
        n11686) );
  OAI211_X1 U14073 ( .C1(n9331), .C2(n11687), .A(n11686), .B(P2_B_REG_SCAN_IN), 
        .ZN(n11688) );
  NAND2_X1 U14074 ( .A1(n12882), .A2(n9339), .ZN(n11721) );
  INV_X1 U14075 ( .A(n11721), .ZN(n11723) );
  XNOR2_X1 U14076 ( .A(n13100), .B(n11729), .ZN(n11722) );
  INV_X1 U14077 ( .A(n11689), .ZN(n11690) );
  XNOR2_X1 U14078 ( .A(n13146), .B(n11724), .ZN(n11693) );
  NAND2_X1 U14079 ( .A1(n12863), .A2(n9339), .ZN(n11692) );
  NAND2_X1 U14080 ( .A1(n11693), .A2(n11692), .ZN(n11694) );
  OAI21_X1 U14081 ( .B1(n11693), .B2(n11692), .A(n11694), .ZN(n12709) );
  INV_X1 U14082 ( .A(n11694), .ZN(n11695) );
  XNOR2_X1 U14083 ( .A(n13141), .B(n11729), .ZN(n11698) );
  NAND2_X1 U14084 ( .A1(n12864), .A2(n9339), .ZN(n11696) );
  XNOR2_X1 U14085 ( .A(n11698), .B(n11696), .ZN(n12740) );
  INV_X1 U14086 ( .A(n11696), .ZN(n11697) );
  AND2_X1 U14087 ( .A1(n12867), .A2(n9339), .ZN(n11700) );
  XNOR2_X1 U14088 ( .A(n13136), .B(n11729), .ZN(n11699) );
  NOR2_X1 U14089 ( .A1(n11699), .A2(n11700), .ZN(n11701) );
  AOI21_X1 U14090 ( .B1(n11700), .B2(n11699), .A(n11701), .ZN(n12683) );
  INV_X1 U14091 ( .A(n11701), .ZN(n11702) );
  XNOR2_X1 U14092 ( .A(n13131), .B(n11729), .ZN(n11704) );
  AND2_X1 U14093 ( .A1(n12869), .A2(n9339), .ZN(n11703) );
  NOR2_X1 U14094 ( .A1(n11704), .A2(n11703), .ZN(n12722) );
  NAND2_X1 U14095 ( .A1(n11704), .A2(n11703), .ZN(n12723) );
  XNOR2_X1 U14096 ( .A(n13126), .B(n11729), .ZN(n11705) );
  NAND2_X1 U14097 ( .A1(n12872), .A2(n9339), .ZN(n11706) );
  XNOR2_X1 U14098 ( .A(n11705), .B(n11706), .ZN(n12692) );
  INV_X1 U14099 ( .A(n11706), .ZN(n11707) );
  NAND2_X1 U14100 ( .A1(n12874), .A2(n9339), .ZN(n12733) );
  NOR2_X1 U14101 ( .A1(n12734), .A2(n12733), .ZN(n12732) );
  XNOR2_X1 U14102 ( .A(n13116), .B(n11729), .ZN(n11710) );
  INV_X1 U14103 ( .A(n12877), .ZN(n12876) );
  NOR2_X1 U14104 ( .A1(n12876), .A2(n12952), .ZN(n12676) );
  INV_X1 U14105 ( .A(n11709), .ZN(n11711) );
  XNOR2_X1 U14106 ( .A(n13110), .B(n11729), .ZN(n11715) );
  OR2_X1 U14107 ( .A1(n12701), .A2(n11713), .ZN(n11714) );
  NOR2_X1 U14108 ( .A1(n11715), .A2(n11714), .ZN(n11716) );
  AOI21_X1 U14109 ( .B1(n11715), .B2(n11714), .A(n11716), .ZN(n12716) );
  INV_X1 U14110 ( .A(n11716), .ZN(n11717) );
  XNOR2_X1 U14111 ( .A(n13105), .B(n11724), .ZN(n11719) );
  NAND2_X1 U14112 ( .A1(n12880), .A2(n9339), .ZN(n11718) );
  NOR2_X1 U14113 ( .A1(n11719), .A2(n11718), .ZN(n11720) );
  AOI21_X1 U14114 ( .B1(n11719), .B2(n11718), .A(n11720), .ZN(n12698) );
  XNOR2_X1 U14115 ( .A(n11722), .B(n11721), .ZN(n12752) );
  XNOR2_X1 U14116 ( .A(n12911), .B(n11724), .ZN(n11726) );
  NOR2_X1 U14117 ( .A1(n12883), .A2(n12952), .ZN(n11725) );
  NAND2_X1 U14118 ( .A1(n11726), .A2(n11725), .ZN(n11727) );
  OAI21_X1 U14119 ( .B1(n11726), .B2(n11725), .A(n11727), .ZN(n12667) );
  NAND2_X1 U14120 ( .A1(n12884), .A2(n9339), .ZN(n11728) );
  XNOR2_X1 U14121 ( .A(n11729), .B(n11728), .ZN(n11730) );
  XNOR2_X1 U14122 ( .A(n7078), .B(n11730), .ZN(n11731) );
  INV_X1 U14123 ( .A(n11732), .ZN(n12893) );
  NAND2_X1 U14124 ( .A1(n12768), .A2(n12824), .ZN(n11733) );
  OAI21_X1 U14125 ( .B1(n12883), .B2(n12848), .A(n11733), .ZN(n12890) );
  AOI22_X1 U14126 ( .A1(n12757), .A2(n12890), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11734) );
  OAI21_X1 U14127 ( .B1(n12893), .B2(n12742), .A(n11734), .ZN(n11735) );
  AOI21_X1 U14128 ( .B1(n7078), .B2(n12747), .A(n11735), .ZN(n11736) );
  OAI21_X1 U14129 ( .B1(n11737), .B2(n12749), .A(n11736), .ZN(P2_U3192) );
  OR2_X1 U14130 ( .A1(n11741), .A2(n11740), .ZN(n11742) );
  NAND2_X1 U14131 ( .A1(n14136), .A2(n9889), .ZN(n11744) );
  NAND2_X1 U14132 ( .A1(n6452), .A2(n13341), .ZN(n11743) );
  NAND2_X1 U14133 ( .A1(n11744), .A2(n11743), .ZN(n11745) );
  XNOR2_X1 U14134 ( .A(n11745), .B(n11813), .ZN(n11748) );
  NOR2_X1 U14135 ( .A1(n11815), .A2(n13966), .ZN(n11746) );
  AOI21_X1 U14136 ( .B1(n14136), .B2(n6452), .A(n11746), .ZN(n11747) );
  NAND2_X1 U14137 ( .A1(n11748), .A2(n11747), .ZN(n11750) );
  OAI21_X1 U14138 ( .B1(n11748), .B2(n11747), .A(n11750), .ZN(n13226) );
  INV_X1 U14139 ( .A(n13226), .ZN(n11749) );
  NAND2_X1 U14140 ( .A1(n13337), .A2(n9889), .ZN(n11752) );
  NAND2_X1 U14141 ( .A1(n6452), .A2(n14088), .ZN(n11751) );
  NAND2_X1 U14142 ( .A1(n11752), .A2(n11751), .ZN(n11753) );
  XNOR2_X1 U14143 ( .A(n11753), .B(n11856), .ZN(n11755) );
  OAI22_X1 U14144 ( .A1(n14132), .A2(n11823), .B1(n13228), .B2(n11815), .ZN(
        n13330) );
  INV_X1 U14145 ( .A(n11754), .ZN(n11756) );
  NAND2_X1 U14146 ( .A1(n14089), .A2(n9889), .ZN(n11759) );
  NAND2_X1 U14147 ( .A1(n13340), .A2(n6452), .ZN(n11758) );
  NAND2_X1 U14148 ( .A1(n11759), .A2(n11758), .ZN(n11760) );
  XNOR2_X1 U14149 ( .A(n11760), .B(n11813), .ZN(n11763) );
  AND2_X1 U14150 ( .A1(n11858), .A2(n13340), .ZN(n11761) );
  AOI21_X1 U14151 ( .B1(n14089), .B2(n6452), .A(n11761), .ZN(n11762) );
  NAND2_X1 U14152 ( .A1(n11763), .A2(n11762), .ZN(n13273) );
  OAI21_X1 U14153 ( .B1(n11763), .B2(n11762), .A(n13273), .ZN(n14072) );
  INV_X1 U14154 ( .A(n14072), .ZN(n11764) );
  OAI22_X1 U14155 ( .A1(n13522), .A2(n11824), .B1(n11765), .B2(n11823), .ZN(
        n11766) );
  XNOR2_X1 U14156 ( .A(n11766), .B(n11813), .ZN(n11769) );
  OR2_X1 U14157 ( .A1(n13522), .A2(n11823), .ZN(n11768) );
  NAND2_X1 U14158 ( .A1(n14086), .A2(n11858), .ZN(n11767) );
  AND2_X1 U14159 ( .A1(n11768), .A2(n11767), .ZN(n11770) );
  NAND2_X1 U14160 ( .A1(n11769), .A2(n11770), .ZN(n11775) );
  INV_X1 U14161 ( .A(n11769), .ZN(n11772) );
  INV_X1 U14162 ( .A(n11770), .ZN(n11771) );
  NAND2_X1 U14163 ( .A1(n11772), .A2(n11771), .ZN(n11773) );
  AND2_X1 U14164 ( .A1(n11775), .A2(n11773), .ZN(n13274) );
  NAND2_X1 U14165 ( .A1(n13276), .A2(n11775), .ZN(n13309) );
  NAND2_X1 U14166 ( .A1(n13717), .A2(n9889), .ZN(n11777) );
  NAND2_X1 U14167 ( .A1(n13507), .A2(n6452), .ZN(n11776) );
  NAND2_X1 U14168 ( .A1(n11777), .A2(n11776), .ZN(n11778) );
  XNOR2_X1 U14169 ( .A(n11778), .B(n11856), .ZN(n11783) );
  AOI22_X1 U14170 ( .A1(n13717), .A2(n6452), .B1(n11858), .B2(n13507), .ZN(
        n11781) );
  XNOR2_X1 U14171 ( .A(n11783), .B(n11781), .ZN(n13310) );
  AOI22_X1 U14172 ( .A1(n13700), .A2(n9889), .B1(n6452), .B2(n13709), .ZN(
        n11779) );
  XNOR2_X1 U14173 ( .A(n11779), .B(n11856), .ZN(n11785) );
  AND2_X1 U14174 ( .A1(n13709), .A2(n11858), .ZN(n11780) );
  AOI21_X1 U14175 ( .B1(n13700), .B2(n6452), .A(n11780), .ZN(n11786) );
  XNOR2_X1 U14176 ( .A(n11785), .B(n11786), .ZN(n13244) );
  INV_X1 U14177 ( .A(n11781), .ZN(n11782) );
  NOR2_X1 U14178 ( .A1(n11783), .A2(n11782), .ZN(n13245) );
  NOR2_X1 U14179 ( .A1(n13244), .A2(n13245), .ZN(n11784) );
  INV_X1 U14180 ( .A(n11785), .ZN(n11788) );
  INV_X1 U14181 ( .A(n11786), .ZN(n11787) );
  OR2_X1 U14182 ( .A1(n13799), .A2(n11823), .ZN(n11790) );
  NAND2_X1 U14183 ( .A1(n13256), .A2(n11858), .ZN(n11789) );
  NAND2_X1 U14184 ( .A1(n11790), .A2(n11789), .ZN(n11792) );
  OAI22_X1 U14185 ( .A1(n13799), .A2(n11824), .B1(n13528), .B2(n11823), .ZN(
        n11791) );
  XNOR2_X1 U14186 ( .A(n11791), .B(n11856), .ZN(n11793) );
  XOR2_X1 U14187 ( .A(n11792), .B(n11793), .Z(n13292) );
  NAND2_X1 U14188 ( .A1(n11793), .A2(n11792), .ZN(n11794) );
  NAND2_X1 U14189 ( .A1(n13529), .A2(n9889), .ZN(n11796) );
  NAND2_X1 U14190 ( .A1(n13678), .A2(n6452), .ZN(n11795) );
  NAND2_X1 U14191 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  XNOR2_X1 U14192 ( .A(n11797), .B(n11813), .ZN(n11800) );
  AND2_X1 U14193 ( .A1(n13678), .A2(n11858), .ZN(n11798) );
  AOI21_X1 U14194 ( .B1(n13529), .B2(n6452), .A(n11798), .ZN(n11799) );
  NAND2_X1 U14195 ( .A1(n11800), .A2(n11799), .ZN(n13300) );
  OAI21_X1 U14196 ( .B1(n11800), .B2(n11799), .A(n13300), .ZN(n13254) );
  INV_X1 U14197 ( .A(n13254), .ZN(n11801) );
  NAND2_X1 U14198 ( .A1(n13661), .A2(n9889), .ZN(n11803) );
  NAND2_X1 U14199 ( .A1(n13513), .A2(n6452), .ZN(n11802) );
  NAND2_X1 U14200 ( .A1(n11803), .A2(n11802), .ZN(n11804) );
  XNOR2_X1 U14201 ( .A(n11804), .B(n11813), .ZN(n11806) );
  AND2_X1 U14202 ( .A1(n13513), .A2(n11858), .ZN(n11805) );
  AOI21_X1 U14203 ( .B1(n13661), .B2(n6452), .A(n11805), .ZN(n11807) );
  NAND2_X1 U14204 ( .A1(n11806), .A2(n11807), .ZN(n13234) );
  INV_X1 U14205 ( .A(n11806), .ZN(n11809) );
  INV_X1 U14206 ( .A(n11807), .ZN(n11808) );
  NAND2_X1 U14207 ( .A1(n11809), .A2(n11808), .ZN(n11810) );
  NAND2_X1 U14208 ( .A1(n13778), .A2(n9889), .ZN(n11812) );
  NAND2_X1 U14209 ( .A1(n6452), .A2(n13516), .ZN(n11811) );
  NAND2_X1 U14210 ( .A1(n11812), .A2(n11811), .ZN(n11814) );
  XNOR2_X1 U14211 ( .A(n11814), .B(n11813), .ZN(n11817) );
  NOR2_X1 U14212 ( .A1(n11815), .A2(n13532), .ZN(n11816) );
  AOI21_X1 U14213 ( .B1(n13778), .B2(n6436), .A(n11816), .ZN(n11818) );
  NAND2_X1 U14214 ( .A1(n11817), .A2(n11818), .ZN(n11822) );
  INV_X1 U14215 ( .A(n11817), .ZN(n11820) );
  INV_X1 U14216 ( .A(n11818), .ZN(n11819) );
  NAND2_X1 U14217 ( .A1(n11820), .A2(n11819), .ZN(n11821) );
  AND2_X1 U14218 ( .A1(n11822), .A2(n11821), .ZN(n13235) );
  OAI22_X1 U14219 ( .A1(n13772), .A2(n11824), .B1(n13607), .B2(n11823), .ZN(
        n11825) );
  XNOR2_X1 U14220 ( .A(n11825), .B(n11856), .ZN(n11829) );
  OR2_X1 U14221 ( .A1(n13772), .A2(n11823), .ZN(n11827) );
  NAND2_X1 U14222 ( .A1(n11858), .A2(n6879), .ZN(n11826) );
  NAND2_X1 U14223 ( .A1(n11827), .A2(n11826), .ZN(n11828) );
  NOR2_X1 U14224 ( .A1(n11829), .A2(n11828), .ZN(n11830) );
  AOI21_X1 U14225 ( .B1(n11829), .B2(n11828), .A(n11830), .ZN(n13286) );
  NAND2_X1 U14226 ( .A1(n13763), .A2(n9889), .ZN(n11832) );
  NAND2_X1 U14227 ( .A1(n6436), .A2(n13533), .ZN(n11831) );
  NAND2_X1 U14228 ( .A1(n11832), .A2(n11831), .ZN(n11833) );
  XNOR2_X1 U14229 ( .A(n11833), .B(n11856), .ZN(n11837) );
  NAND2_X1 U14230 ( .A1(n13763), .A2(n6452), .ZN(n11835) );
  NAND2_X1 U14231 ( .A1(n11858), .A2(n13533), .ZN(n11834) );
  NAND2_X1 U14232 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  NOR2_X1 U14233 ( .A1(n11837), .A2(n11836), .ZN(n11838) );
  AOI21_X1 U14234 ( .B1(n11837), .B2(n11836), .A(n11838), .ZN(n13264) );
  INV_X1 U14235 ( .A(n11838), .ZN(n11839) );
  NAND2_X1 U14236 ( .A1(n13491), .A2(n9889), .ZN(n11841) );
  NAND2_X1 U14237 ( .A1(n6452), .A2(n13608), .ZN(n11840) );
  NAND2_X1 U14238 ( .A1(n11841), .A2(n11840), .ZN(n11842) );
  XNOR2_X1 U14239 ( .A(n11842), .B(n11856), .ZN(n11846) );
  NAND2_X1 U14240 ( .A1(n13491), .A2(n6452), .ZN(n11844) );
  NAND2_X1 U14241 ( .A1(n11858), .A2(n13608), .ZN(n11843) );
  NAND2_X1 U14242 ( .A1(n11844), .A2(n11843), .ZN(n11845) );
  NOR2_X1 U14243 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  AOI21_X1 U14244 ( .B1(n11846), .B2(n11845), .A(n11847), .ZN(n13319) );
  NAND2_X1 U14245 ( .A1(n13750), .A2(n9889), .ZN(n11849) );
  NAND2_X1 U14246 ( .A1(n6452), .A2(n13556), .ZN(n11848) );
  NAND2_X1 U14247 ( .A1(n11849), .A2(n11848), .ZN(n11850) );
  XNOR2_X1 U14248 ( .A(n11850), .B(n11856), .ZN(n11854) );
  NAND2_X1 U14249 ( .A1(n13750), .A2(n6452), .ZN(n11852) );
  NAND2_X1 U14250 ( .A1(n11858), .A2(n13556), .ZN(n11851) );
  NAND2_X1 U14251 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  NOR2_X1 U14252 ( .A1(n11854), .A2(n11853), .ZN(n11855) );
  AOI21_X1 U14253 ( .B1(n11854), .B2(n11853), .A(n11855), .ZN(n13219) );
  AOI22_X1 U14254 ( .A1(n13745), .A2(n9889), .B1(n6452), .B2(n13547), .ZN(
        n11857) );
  XNOR2_X1 U14255 ( .A(n11857), .B(n11856), .ZN(n11860) );
  AOI22_X1 U14256 ( .A1(n13745), .A2(n6436), .B1(n11858), .B2(n13547), .ZN(
        n11859) );
  XNOR2_X1 U14257 ( .A(n11860), .B(n11859), .ZN(n11861) );
  XNOR2_X1 U14258 ( .A(n11862), .B(n11861), .ZN(n11868) );
  AOI22_X1 U14259 ( .A1(n14073), .A2(n13556), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11864) );
  NAND2_X1 U14260 ( .A1(n13326), .A2(n13563), .ZN(n11863) );
  OAI211_X1 U14261 ( .C1(n11865), .C2(n13313), .A(n11864), .B(n11863), .ZN(
        n11866) );
  AOI21_X1 U14262 ( .B1(n13745), .B2(n14075), .A(n11866), .ZN(n11867) );
  OAI21_X1 U14263 ( .B1(n11868), .B2(n14078), .A(n11867), .ZN(P1_U3220) );
  OAI222_X1 U14264 ( .A1(n13833), .A2(n11871), .B1(n13837), .B2(n11870), .C1(
        P1_U3086), .C2(n11869), .ZN(P1_U3334) );
  XNOR2_X1 U14265 ( .A(n12497), .B(n9067), .ZN(n11917) );
  XNOR2_X1 U14266 ( .A(n11917), .B(n12264), .ZN(n11918) );
  INV_X1 U14267 ( .A(n11881), .ZN(n11872) );
  OAI22_X1 U14268 ( .A1(n11872), .A2(n11906), .B1(n12178), .B2(n11877), .ZN(
        n11874) );
  AOI21_X1 U14269 ( .B1(n11873), .B2(n12363), .A(n11874), .ZN(n11883) );
  AOI21_X1 U14270 ( .B1(n11877), .B2(n12178), .A(n11906), .ZN(n11880) );
  INV_X1 U14271 ( .A(n11874), .ZN(n11876) );
  NAND3_X1 U14272 ( .A1(n11876), .A2(n12384), .A3(n11875), .ZN(n11879) );
  NAND3_X1 U14273 ( .A1(n11877), .A2(n12178), .A3(n11906), .ZN(n11878) );
  OAI211_X1 U14274 ( .C1(n11881), .C2(n11880), .A(n11879), .B(n11878), .ZN(
        n11882) );
  XNOR2_X1 U14275 ( .A(n12343), .B(n9067), .ZN(n11885) );
  XNOR2_X1 U14276 ( .A(n11885), .B(n12266), .ZN(n11945) );
  OAI22_X1 U14277 ( .A1(n11944), .A2(n11945), .B1(n11885), .B2(n12266), .ZN(
        n12007) );
  XNOR2_X1 U14278 ( .A(n12500), .B(n9067), .ZN(n11886) );
  XNOR2_X1 U14279 ( .A(n11886), .B(n12314), .ZN(n12008) );
  INV_X1 U14280 ( .A(n11886), .ZN(n11887) );
  XOR2_X1 U14281 ( .A(n11918), .B(n11919), .Z(n11893) );
  INV_X1 U14282 ( .A(n12314), .ZN(n12265) );
  AOI22_X1 U14283 ( .A1(n12003), .A2(n12265), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11890) );
  INV_X1 U14284 ( .A(n11888), .ZN(n12318) );
  NAND2_X1 U14285 ( .A1(n11977), .A2(n12318), .ZN(n11889) );
  OAI211_X1 U14286 ( .C1(n12316), .C2(n12000), .A(n11890), .B(n11889), .ZN(
        n11891) );
  AOI21_X1 U14287 ( .B1(n12497), .B2(n14675), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14288 ( .B1(n11893), .B2(n12023), .A(n11892), .ZN(P3_U3154) );
  XNOR2_X1 U14289 ( .A(n11895), .B(n11894), .ZN(n11896) );
  XNOR2_X1 U14290 ( .A(n11897), .B(n11896), .ZN(n11902) );
  INV_X1 U14291 ( .A(n12623), .ZN(n12476) );
  NOR2_X1 U14292 ( .A1(n14678), .A2(n12478), .ZN(n11900) );
  AOI22_X1 U14293 ( .A1(n12003), .A2(n11980), .B1(P3_REG3_REG_14__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11898) );
  OAI21_X1 U14294 ( .B1(n12468), .B2(n12000), .A(n11898), .ZN(n11899) );
  AOI211_X1 U14295 ( .C1(n12476), .C2(n14675), .A(n11900), .B(n11899), .ZN(
        n11901) );
  OAI21_X1 U14296 ( .B1(n11902), .B2(n12023), .A(n11901), .ZN(P3_U3155) );
  XNOR2_X1 U14297 ( .A(n11903), .B(n12178), .ZN(n11909) );
  AOI22_X1 U14298 ( .A1(n12003), .A2(n12363), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11905) );
  NAND2_X1 U14299 ( .A1(n11977), .A2(n12366), .ZN(n11904) );
  OAI211_X1 U14300 ( .C1(n11906), .C2(n12000), .A(n11905), .B(n11904), .ZN(
        n11907) );
  AOI21_X1 U14301 ( .B1(n12572), .B2(n14675), .A(n11907), .ZN(n11908) );
  OAI21_X1 U14302 ( .B1(n11909), .B2(n12023), .A(n11908), .ZN(P3_U3156) );
  OAI211_X1 U14303 ( .C1(n11912), .C2(n11911), .A(n11910), .B(n14668), .ZN(
        n11916) );
  AOI22_X1 U14304 ( .A1(n12269), .A2(n14730), .B1(n14731), .B2(n12434), .ZN(
        n12406) );
  OAI21_X1 U14305 ( .B1(n12406), .B2(n14666), .A(n11913), .ZN(n11914) );
  AOI21_X1 U14306 ( .B1(n11977), .B2(n12410), .A(n11914), .ZN(n11915) );
  OAI211_X1 U14307 ( .C1(n12006), .C2(n12593), .A(n11916), .B(n11915), .ZN(
        P3_U3159) );
  XNOR2_X1 U14308 ( .A(n12300), .B(n9067), .ZN(n11920) );
  NAND2_X1 U14309 ( .A1(n12262), .A2(n14730), .ZN(n11921) );
  OAI21_X1 U14310 ( .B1(n12009), .B2(n14762), .A(n11921), .ZN(n12302) );
  AOI22_X1 U14311 ( .A1(n12019), .A2(n12302), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11922) );
  OAI21_X1 U14312 ( .B1(n14678), .B2(n12306), .A(n11922), .ZN(n11923) );
  AOI21_X1 U14313 ( .B1(n12552), .B2(n14675), .A(n11923), .ZN(n11924) );
  INV_X1 U14314 ( .A(n11925), .ZN(n11926) );
  AOI21_X1 U14315 ( .B1(n11928), .B2(n11927), .A(n11926), .ZN(n11934) );
  OAI22_X1 U14316 ( .A1(n12384), .A2(n12000), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11929), .ZN(n11931) );
  NOR2_X1 U14317 ( .A1(n11974), .A2(n12383), .ZN(n11930) );
  AOI211_X1 U14318 ( .C1(n11977), .C2(n12387), .A(n11931), .B(n11930), .ZN(
        n11933) );
  NAND2_X1 U14319 ( .A1(n12388), .A2(n14675), .ZN(n11932) );
  OAI211_X1 U14320 ( .C1(n11934), .C2(n12023), .A(n11933), .B(n11932), .ZN(
        P3_U3163) );
  XOR2_X1 U14321 ( .A(n11935), .B(n11936), .Z(n11943) );
  NOR2_X1 U14322 ( .A1(n14678), .A2(n11937), .ZN(n11940) );
  AOI22_X1 U14323 ( .A1(n12003), .A2(n14729), .B1(P3_REG3_REG_12__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11938) );
  OAI21_X1 U14324 ( .B1(n12469), .B2(n12000), .A(n11938), .ZN(n11939) );
  AOI211_X1 U14325 ( .C1(n11941), .C2(n14675), .A(n11940), .B(n11939), .ZN(
        n11942) );
  OAI21_X1 U14326 ( .B1(n11943), .B2(n12023), .A(n11942), .ZN(P3_U3164) );
  XOR2_X1 U14327 ( .A(n11945), .B(n11944), .Z(n11951) );
  AND2_X1 U14328 ( .A1(n12362), .A2(n14731), .ZN(n11946) );
  AOI21_X1 U14329 ( .B1(n12265), .B2(n14730), .A(n11946), .ZN(n12337) );
  INV_X1 U14330 ( .A(n12337), .ZN(n11947) );
  AOI22_X1 U14331 ( .A1(n11947), .A2(n12019), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11948) );
  OAI21_X1 U14332 ( .B1(n12341), .B2(n14678), .A(n11948), .ZN(n11949) );
  AOI21_X1 U14333 ( .B1(n12343), .B2(n14675), .A(n11949), .ZN(n11950) );
  OAI21_X1 U14334 ( .B1(n11951), .B2(n12023), .A(n11950), .ZN(P3_U3165) );
  XNOR2_X1 U14335 ( .A(n11952), .B(n12018), .ZN(n11953) );
  XNOR2_X1 U14336 ( .A(n11954), .B(n11953), .ZN(n11959) );
  OAI22_X1 U14337 ( .A1(n12419), .A2(n14760), .B1(n12468), .B2(n14762), .ZN(
        n12445) );
  NAND2_X1 U14338 ( .A1(n12445), .A2(n12019), .ZN(n11955) );
  NAND2_X1 U14339 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14012)
         );
  OAI211_X1 U14340 ( .C1(n14678), .C2(n11956), .A(n11955), .B(n14012), .ZN(
        n11957) );
  AOI21_X1 U14341 ( .B1(n12609), .B2(n14675), .A(n11957), .ZN(n11958) );
  OAI21_X1 U14342 ( .B1(n11959), .B2(n12023), .A(n11958), .ZN(P3_U3166) );
  OAI211_X1 U14343 ( .C1(n11962), .C2(n11961), .A(n11960), .B(n14668), .ZN(
        n11968) );
  NOR2_X1 U14344 ( .A1(n14678), .A2(n12436), .ZN(n11966) );
  OAI22_X1 U14345 ( .A1(n12000), .A2(n11964), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11963), .ZN(n11965) );
  AOI211_X1 U14346 ( .C1(n12003), .C2(n12433), .A(n11966), .B(n11965), .ZN(
        n11967) );
  OAI211_X1 U14347 ( .C1(n11969), .C2(n12006), .A(n11968), .B(n11967), .ZN(
        P3_U3168) );
  OAI211_X1 U14348 ( .C1(n11972), .C2(n11971), .A(n11970), .B(n14668), .ZN(
        n11979) );
  OAI22_X1 U14349 ( .A1(n12000), .A2(n12396), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11973), .ZN(n11976) );
  NOR2_X1 U14350 ( .A1(n11974), .A2(n12420), .ZN(n11975) );
  AOI211_X1 U14351 ( .C1(n11977), .C2(n12399), .A(n11976), .B(n11975), .ZN(
        n11978) );
  OAI211_X1 U14352 ( .C1(n12588), .C2(n12006), .A(n11979), .B(n11978), .ZN(
        P3_U3173) );
  XNOR2_X1 U14353 ( .A(n11981), .B(n11980), .ZN(n11982) );
  XNOR2_X1 U14354 ( .A(n11983), .B(n11982), .ZN(n11989) );
  NOR2_X1 U14355 ( .A1(n12006), .A2(n12634), .ZN(n11988) );
  NAND2_X1 U14356 ( .A1(n12272), .A2(n14730), .ZN(n11984) );
  OAI21_X1 U14357 ( .B1(n11985), .B2(n14762), .A(n11984), .ZN(n12485) );
  AOI22_X1 U14358 ( .A1(n12019), .A2(n12485), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11986) );
  OAI21_X1 U14359 ( .B1(n14678), .B2(n12487), .A(n11986), .ZN(n11987) );
  AOI211_X1 U14360 ( .C1(n11989), .C2(n14668), .A(n11988), .B(n11987), .ZN(
        n11990) );
  INV_X1 U14361 ( .A(n11990), .ZN(P3_U3174) );
  XNOR2_X1 U14362 ( .A(n11991), .B(n12363), .ZN(n11996) );
  INV_X1 U14363 ( .A(n12375), .ZN(n11993) );
  OAI22_X1 U14364 ( .A1(n12178), .A2(n14760), .B1(n12396), .B2(n14762), .ZN(
        n12372) );
  AOI22_X1 U14365 ( .A1(n12372), .A2(n12019), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11992) );
  OAI21_X1 U14366 ( .B1(n11993), .B2(n14678), .A(n11992), .ZN(n11994) );
  AOI21_X1 U14367 ( .B1(n12578), .B2(n14675), .A(n11994), .ZN(n11995) );
  OAI21_X1 U14368 ( .B1(n11996), .B2(n12023), .A(n11995), .ZN(P3_U3175) );
  OAI211_X1 U14369 ( .C1(n11999), .C2(n11998), .A(n11997), .B(n14668), .ZN(
        n12005) );
  NOR2_X1 U14370 ( .A1(n14678), .A2(n12421), .ZN(n12002) );
  NAND2_X1 U14371 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n14045)
         );
  OAI21_X1 U14372 ( .B1(n12000), .B2(n12420), .A(n14045), .ZN(n12001) );
  AOI211_X1 U14373 ( .C1(n12003), .C2(n12271), .A(n12002), .B(n12001), .ZN(
        n12004) );
  OAI211_X1 U14374 ( .C1(n12600), .C2(n12006), .A(n12005), .B(n12004), .ZN(
        P3_U3178) );
  XOR2_X1 U14375 ( .A(n12008), .B(n12007), .Z(n12013) );
  OAI22_X1 U14376 ( .A1(n12189), .A2(n14762), .B1(n12009), .B2(n14760), .ZN(
        n12323) );
  AOI22_X1 U14377 ( .A1(n12323), .A2(n12019), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12010) );
  OAI21_X1 U14378 ( .B1(n12327), .B2(n14678), .A(n12010), .ZN(n12011) );
  AOI21_X1 U14379 ( .B1(n12500), .B2(n14675), .A(n12011), .ZN(n12012) );
  OAI21_X1 U14380 ( .B1(n12013), .B2(n12023), .A(n12012), .ZN(P3_U3180) );
  XNOR2_X1 U14381 ( .A(n12014), .B(n12468), .ZN(n12015) );
  XNOR2_X1 U14382 ( .A(n12016), .B(n12015), .ZN(n12024) );
  NAND2_X1 U14383 ( .A1(n12272), .A2(n14731), .ZN(n12017) );
  OAI21_X1 U14384 ( .B1(n12018), .B2(n14760), .A(n12017), .ZN(n12456) );
  AOI22_X1 U14385 ( .A1(n12019), .A2(n12456), .B1(P3_REG3_REG_15__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12020) );
  OAI21_X1 U14386 ( .B1(n14678), .B2(n12460), .A(n12020), .ZN(n12021) );
  AOI21_X1 U14387 ( .B1(n12616), .B2(n14675), .A(n12021), .ZN(n12022) );
  OAI21_X1 U14388 ( .B1(n12024), .B2(n12023), .A(n12022), .ZN(P3_U3181) );
  INV_X1 U14389 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13822) );
  NAND2_X1 U14390 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12038), .ZN(n12027) );
  AOI22_X1 U14391 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n13822), .B1(n12041), 
        .B2(n12027), .ZN(n12031) );
  INV_X1 U14392 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U14393 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(n12029), .B1(
        P1_DATAO_REG_31__SCAN_IN), .B2(n12028), .ZN(n12030) );
  XNOR2_X1 U14394 ( .A(n12031), .B(n12030), .ZN(n12638) );
  INV_X1 U14395 ( .A(SI_31_), .ZN(n12642) );
  NOR2_X1 U14396 ( .A1(n8601), .A2(n12642), .ZN(n12032) );
  AOI21_X1 U14397 ( .B1(n12638), .B2(n8611), .A(n12032), .ZN(n12051) );
  NAND2_X1 U14398 ( .A1(n6457), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12036) );
  NAND2_X1 U14399 ( .A1(n8719), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12035) );
  NAND2_X1 U14400 ( .A1(n12033), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n12034) );
  NAND4_X1 U14401 ( .A1(n12037), .A2(n12036), .A3(n12035), .A4(n12034), .ZN(
        n14049) );
  NAND2_X1 U14402 ( .A1(n12051), .A2(n14049), .ZN(n12047) );
  AOI22_X1 U14403 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n12038), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n13822), .ZN(n12039) );
  INV_X1 U14404 ( .A(n12039), .ZN(n12040) );
  XNOR2_X1 U14405 ( .A(n12041), .B(n12040), .ZN(n12643) );
  NAND2_X1 U14406 ( .A1(n12643), .A2(n12042), .ZN(n12045) );
  INV_X1 U14407 ( .A(SI_30_), .ZN(n12645) );
  OR2_X1 U14408 ( .A1(n12043), .A2(n12645), .ZN(n12044) );
  NAND2_X1 U14409 ( .A1(n12045), .A2(n12044), .ZN(n14057) );
  INV_X1 U14410 ( .A(n12261), .ZN(n12050) );
  NAND2_X1 U14411 ( .A1(n14057), .A2(n12050), .ZN(n12046) );
  INV_X1 U14412 ( .A(n14049), .ZN(n12049) );
  AOI21_X1 U14413 ( .B1(n14057), .B2(n12049), .A(n12206), .ZN(n12048) );
  NAND2_X1 U14414 ( .A1(n12052), .A2(n12049), .ZN(n12243) );
  OR2_X1 U14415 ( .A1(n14057), .A2(n12050), .ZN(n12214) );
  XNOR2_X1 U14416 ( .A(n12056), .B(n12055), .ZN(n12213) );
  NAND2_X1 U14417 ( .A1(n12266), .A2(n12183), .ZN(n12192) );
  INV_X1 U14418 ( .A(n12062), .ZN(n12057) );
  AOI21_X1 U14419 ( .B1(n12422), .B2(n12058), .A(n12057), .ZN(n12059) );
  AND2_X1 U14420 ( .A1(n12217), .A2(n12059), .ZN(n12067) );
  INV_X1 U14421 ( .A(n12060), .ZN(n12061) );
  NAND2_X1 U14422 ( .A1(n12062), .A2(n12061), .ZN(n12064) );
  NAND2_X1 U14423 ( .A1(n12064), .A2(n12063), .ZN(n12065) );
  NOR2_X1 U14424 ( .A1(n12216), .A2(n12065), .ZN(n12066) );
  MUX2_X1 U14425 ( .A(n12067), .B(n12066), .S(n12076), .Z(n12162) );
  NAND2_X1 U14426 ( .A1(n12072), .A2(n12068), .ZN(n12071) );
  MUX2_X1 U14427 ( .A(n12071), .B(n12070), .S(n12069), .Z(n12075) );
  NAND2_X1 U14428 ( .A1(n12073), .A2(n12076), .ZN(n12074) );
  NAND3_X1 U14429 ( .A1(n12075), .A2(n12077), .A3(n12074), .ZN(n12079) );
  NAND3_X1 U14430 ( .A1(n12079), .A2(n8968), .A3(n12078), .ZN(n12084) );
  NAND2_X1 U14431 ( .A1(n12087), .A2(n12080), .ZN(n12081) );
  NAND2_X1 U14432 ( .A1(n12081), .A2(n12183), .ZN(n12083) );
  INV_X1 U14433 ( .A(n12086), .ZN(n12082) );
  AOI21_X1 U14434 ( .B1(n12084), .B2(n12083), .A(n12082), .ZN(n12092) );
  AOI21_X1 U14435 ( .B1(n12086), .B2(n12085), .A(n12183), .ZN(n12091) );
  NOR2_X1 U14436 ( .A1(n12087), .A2(n12183), .ZN(n12089) );
  NOR2_X1 U14437 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  OAI21_X1 U14438 ( .B1(n12092), .B2(n12091), .A(n12090), .ZN(n12096) );
  MUX2_X1 U14439 ( .A(n12094), .B(n12093), .S(n12076), .Z(n12095) );
  NAND3_X1 U14440 ( .A1(n12096), .A2(n12218), .A3(n12095), .ZN(n12100) );
  NAND2_X1 U14441 ( .A1(n12106), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U14442 ( .A1(n12098), .A2(n12076), .ZN(n12099) );
  NAND2_X1 U14443 ( .A1(n12100), .A2(n12099), .ZN(n12104) );
  AOI21_X1 U14444 ( .B1(n12103), .B2(n12101), .A(n12076), .ZN(n12102) );
  AOI21_X1 U14445 ( .B1(n12104), .B2(n12103), .A(n12102), .ZN(n12112) );
  OAI21_X1 U14446 ( .B1(n12076), .B2(n12106), .A(n12105), .ZN(n12111) );
  NAND2_X1 U14447 ( .A1(n12107), .A2(n14826), .ZN(n12108) );
  MUX2_X1 U14448 ( .A(n12109), .B(n12108), .S(n12183), .Z(n12110) );
  OAI211_X1 U14449 ( .C1(n12112), .C2(n12111), .A(n12222), .B(n12110), .ZN(
        n12117) );
  INV_X1 U14450 ( .A(n12227), .ZN(n12116) );
  MUX2_X1 U14451 ( .A(n12114), .B(n12113), .S(n12076), .Z(n12115) );
  NAND3_X1 U14452 ( .A1(n12117), .A2(n12116), .A3(n12115), .ZN(n12122) );
  MUX2_X1 U14453 ( .A(n14732), .B(n12118), .S(n12076), .Z(n12120) );
  NAND2_X1 U14454 ( .A1(n12120), .A2(n12119), .ZN(n12121) );
  AOI21_X1 U14455 ( .B1(n12122), .B2(n12121), .A(n14735), .ZN(n12129) );
  MUX2_X1 U14456 ( .A(n12124), .B(n12123), .S(n12076), .Z(n12125) );
  NAND2_X1 U14457 ( .A1(n12125), .A2(n12229), .ZN(n12128) );
  AND2_X1 U14458 ( .A1(n12135), .A2(n12126), .ZN(n12127) );
  OAI22_X1 U14459 ( .A1(n12129), .A2(n12128), .B1(n12076), .B2(n12127), .ZN(
        n12133) );
  AOI21_X1 U14460 ( .B1(n12132), .B2(n12130), .A(n12183), .ZN(n12131) );
  AOI21_X1 U14461 ( .B1(n12133), .B2(n12132), .A(n12131), .ZN(n12142) );
  INV_X1 U14462 ( .A(n12138), .ZN(n12134) );
  AND2_X1 U14463 ( .A1(n12134), .A2(n12136), .ZN(n12484) );
  OAI21_X1 U14464 ( .B1(n12183), .B2(n12135), .A(n12484), .ZN(n12141) );
  INV_X1 U14465 ( .A(n12136), .ZN(n12137) );
  MUX2_X1 U14466 ( .A(n12138), .B(n12137), .S(n12183), .Z(n12139) );
  NOR2_X1 U14467 ( .A1(n12139), .A2(n12464), .ZN(n12140) );
  INV_X1 U14468 ( .A(n12454), .ZN(n12451) );
  OAI211_X1 U14469 ( .C1(n12142), .C2(n12141), .A(n12140), .B(n12451), .ZN(
        n12149) );
  NAND2_X1 U14470 ( .A1(n12154), .A2(n12433), .ZN(n12144) );
  OR2_X1 U14471 ( .A1(n12616), .A2(n12468), .ZN(n12143) );
  OAI211_X1 U14472 ( .C1(n12454), .C2(n12145), .A(n12144), .B(n12143), .ZN(
        n12146) );
  NAND2_X1 U14473 ( .A1(n12146), .A2(n12183), .ZN(n12148) );
  INV_X1 U14474 ( .A(n12151), .ZN(n12147) );
  AOI21_X1 U14475 ( .B1(n12149), .B2(n12148), .A(n12147), .ZN(n12157) );
  OAI211_X1 U14476 ( .C1(n12454), .C2(n12152), .A(n12151), .B(n12150), .ZN(
        n12153) );
  AND2_X1 U14477 ( .A1(n12153), .A2(n12076), .ZN(n12156) );
  NAND3_X1 U14478 ( .A1(n12154), .A2(n12076), .A3(n12433), .ZN(n12155) );
  OAI21_X1 U14479 ( .B1(n12157), .B2(n12156), .A(n12155), .ZN(n12158) );
  NAND3_X1 U14480 ( .A1(n12158), .A2(n12432), .A3(n12422), .ZN(n12161) );
  INV_X1 U14481 ( .A(n12217), .ZN(n12159) );
  MUX2_X1 U14482 ( .A(n12216), .B(n12159), .S(n12076), .Z(n12160) );
  AOI21_X1 U14483 ( .B1(n12162), .B2(n12161), .A(n12160), .ZN(n12163) );
  AND2_X1 U14484 ( .A1(n12393), .A2(n12163), .ZN(n12174) );
  INV_X1 U14485 ( .A(n12164), .ZN(n12169) );
  OR2_X1 U14486 ( .A1(n12170), .A2(n12169), .ZN(n12380) );
  NAND2_X1 U14487 ( .A1(n12400), .A2(n12383), .ZN(n12166) );
  MUX2_X1 U14488 ( .A(n12166), .B(n12165), .S(n12076), .Z(n12167) );
  NAND2_X1 U14489 ( .A1(n12378), .A2(n12167), .ZN(n12173) );
  INV_X1 U14490 ( .A(n12168), .ZN(n12175) );
  MUX2_X1 U14491 ( .A(n12170), .B(n12169), .S(n12076), .Z(n12171) );
  INV_X1 U14492 ( .A(n12171), .ZN(n12172) );
  OAI211_X1 U14493 ( .C1(n12174), .C2(n12173), .A(n12371), .B(n12172), .ZN(
        n12180) );
  NAND3_X1 U14494 ( .A1(n12180), .A2(n12360), .A3(n12175), .ZN(n12182) );
  INV_X1 U14495 ( .A(n12176), .ZN(n12177) );
  NOR2_X1 U14496 ( .A1(n12239), .A2(n12177), .ZN(n12179) );
  AOI22_X1 U14497 ( .A1(n12180), .A2(n12179), .B1(n12178), .B2(n12572), .ZN(
        n12181) );
  MUX2_X1 U14498 ( .A(n12182), .B(n12181), .S(n12076), .Z(n12188) );
  NAND2_X1 U14499 ( .A1(n12350), .A2(n6498), .ZN(n12186) );
  XNOR2_X1 U14500 ( .A(n12184), .B(n12183), .ZN(n12185) );
  NAND2_X1 U14501 ( .A1(n12186), .A2(n12185), .ZN(n12187) );
  NAND3_X1 U14502 ( .A1(n12343), .A2(n12189), .A3(n12076), .ZN(n12190) );
  OAI211_X1 U14503 ( .C1(n12343), .C2(n12192), .A(n12191), .B(n12190), .ZN(
        n12196) );
  MUX2_X1 U14504 ( .A(n12194), .B(n12193), .S(n12076), .Z(n12195) );
  NAND2_X1 U14505 ( .A1(n12201), .A2(n12197), .ZN(n12198) );
  NAND2_X1 U14506 ( .A1(n12300), .A2(n12198), .ZN(n12202) );
  INV_X1 U14507 ( .A(n12203), .ZN(n12204) );
  INV_X1 U14508 ( .A(n12206), .ZN(n12207) );
  NAND2_X1 U14509 ( .A1(n12208), .A2(n12207), .ZN(n12209) );
  NAND2_X1 U14510 ( .A1(n12209), .A2(n12214), .ZN(n12210) );
  NAND2_X1 U14511 ( .A1(n12210), .A2(n12215), .ZN(n12211) );
  OAI22_X1 U14512 ( .A1(n12213), .A2(n12212), .B1(n12254), .B2(n12247), .ZN(
        n12252) );
  INV_X1 U14513 ( .A(n12215), .ZN(n12244) );
  NAND2_X1 U14514 ( .A1(n7055), .A2(n12217), .ZN(n12404) );
  INV_X1 U14515 ( .A(n12464), .ZN(n12474) );
  NAND4_X1 U14516 ( .A1(n12220), .A2(n12219), .A3(n8968), .A4(n12218), .ZN(
        n12225) );
  INV_X1 U14517 ( .A(n9945), .ZN(n12223) );
  NAND4_X1 U14518 ( .A1(n14742), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12224) );
  NOR2_X1 U14519 ( .A1(n12225), .A2(n12224), .ZN(n12231) );
  INV_X1 U14520 ( .A(n14735), .ZN(n12230) );
  NOR2_X1 U14521 ( .A1(n12227), .A2(n12226), .ZN(n12228) );
  NAND4_X1 U14522 ( .A1(n12231), .A2(n12230), .A3(n12229), .A4(n12228), .ZN(
        n12233) );
  NOR2_X1 U14523 ( .A1(n12233), .A2(n12232), .ZN(n12234) );
  AND4_X1 U14524 ( .A1(n12432), .A2(n12474), .A3(n12484), .A4(n12234), .ZN(
        n12235) );
  NAND4_X1 U14525 ( .A1(n12235), .A2(n12422), .A3(n12443), .A4(n12451), .ZN(
        n12236) );
  NOR2_X1 U14526 ( .A1(n12404), .A2(n12236), .ZN(n12237) );
  NAND4_X1 U14527 ( .A1(n12371), .A2(n12378), .A3(n12237), .A4(n12393), .ZN(
        n12238) );
  NOR3_X1 U14528 ( .A1(n12239), .A2(n12325), .A3(n12238), .ZN(n12240) );
  XNOR2_X1 U14529 ( .A(n12246), .B(n12245), .ZN(n12250) );
  INV_X1 U14530 ( .A(n12247), .ZN(n12248) );
  INV_X1 U14531 ( .A(n14769), .ZN(n14780) );
  NOR2_X1 U14532 ( .A1(n12252), .A2(n12251), .ZN(n12260) );
  INV_X1 U14533 ( .A(n12253), .ZN(n12255) );
  NOR4_X1 U14534 ( .A1(n14762), .A2(n12255), .A3(n12654), .A4(n12254), .ZN(
        n12258) );
  OAI21_X1 U14535 ( .B1(n12259), .B2(n12256), .A(P3_B_REG_SCAN_IN), .ZN(n12257) );
  OAI22_X1 U14536 ( .A1(n12260), .A2(n12259), .B1(n12258), .B2(n12257), .ZN(
        P3_U3296) );
  MUX2_X1 U14537 ( .A(n14049), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12280), .Z(
        P3_U3522) );
  MUX2_X1 U14538 ( .A(n12261), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12280), .Z(
        P3_U3521) );
  MUX2_X1 U14539 ( .A(n12262), .B(P3_DATAO_REG_29__SCAN_IN), .S(n12280), .Z(
        P3_U3520) );
  MUX2_X1 U14540 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12263), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14541 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12264), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14542 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12265), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14543 ( .A(n12266), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12280), .Z(
        P3_U3516) );
  MUX2_X1 U14544 ( .A(n12362), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12280), .Z(
        P3_U3515) );
  MUX2_X1 U14545 ( .A(n12267), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12280), .Z(
        P3_U3514) );
  MUX2_X1 U14546 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12363), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14547 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12268), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14548 ( .A(n12269), .B(P3_DATAO_REG_20__SCAN_IN), .S(n12280), .Z(
        P3_U3511) );
  MUX2_X1 U14549 ( .A(n12270), .B(P3_DATAO_REG_19__SCAN_IN), .S(n12280), .Z(
        P3_U3510) );
  MUX2_X1 U14550 ( .A(n12434), .B(P3_DATAO_REG_18__SCAN_IN), .S(n12280), .Z(
        P3_U3509) );
  MUX2_X1 U14551 ( .A(n12271), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12280), .Z(
        P3_U3508) );
  MUX2_X1 U14552 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12433), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14553 ( .A(n12272), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12280), .Z(
        P3_U3505) );
  MUX2_X1 U14554 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12273), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14555 ( .A(n14729), .B(P3_DATAO_REG_11__SCAN_IN), .S(n12280), .Z(
        P3_U3502) );
  MUX2_X1 U14556 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12274), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14557 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n14732), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U14558 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12275), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14559 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12276), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U14560 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12277), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14561 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12278), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14562 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12279), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14563 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9045), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U14564 ( .A(n12281), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12280), .Z(
        P3_U3491) );
  AOI21_X1 U14565 ( .B1(n12459), .B2(n12283), .A(n12282), .ZN(n12298) );
  OAI21_X1 U14566 ( .B1(P3_REG1_REG_15__SCAN_IN), .B2(n12285), .A(n12284), 
        .ZN(n12296) );
  AOI21_X1 U14567 ( .B1(n12288), .B2(n12287), .A(n12286), .ZN(n12294) );
  INV_X1 U14568 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n12289) );
  NOR2_X1 U14569 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12289), .ZN(n12291) );
  INV_X1 U14570 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14930) );
  NOR2_X1 U14571 ( .A1(n14724), .A2(n14930), .ZN(n12290) );
  AOI211_X1 U14572 ( .C1(n14686), .C2(n12292), .A(n12291), .B(n12290), .ZN(
        n12293) );
  OAI21_X1 U14573 ( .B1(n12294), .B2(n14036), .A(n12293), .ZN(n12295) );
  AOI21_X1 U14574 ( .B1(n14703), .B2(n12296), .A(n12295), .ZN(n12297) );
  OAI21_X1 U14575 ( .B1(n12298), .B2(n14708), .A(n12297), .ZN(P3_U3197) );
  XNOR2_X1 U14576 ( .A(n12299), .B(n12300), .ZN(n12555) );
  INV_X1 U14577 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12305) );
  AOI21_X1 U14578 ( .B1(n12301), .B2(n12300), .A(n12418), .ZN(n12304) );
  AOI21_X1 U14579 ( .B1(n12304), .B2(n12303), .A(n12302), .ZN(n12550) );
  MUX2_X1 U14580 ( .A(n12305), .B(n12550), .S(n14791), .Z(n12309) );
  INV_X1 U14581 ( .A(n12306), .ZN(n12307) );
  AOI22_X1 U14582 ( .A1(n12552), .A2(n6433), .B1(n14772), .B2(n12307), .ZN(
        n12308) );
  OAI211_X1 U14583 ( .C1(n12493), .C2(n12555), .A(n12309), .B(n12308), .ZN(
        P3_U3205) );
  XNOR2_X1 U14584 ( .A(n12310), .B(n12311), .ZN(n12557) );
  XNOR2_X1 U14585 ( .A(n12313), .B(n12312), .ZN(n12315) );
  OAI222_X1 U14586 ( .A1(n14760), .A2(n12316), .B1(n12315), .B2(n12418), .C1(
        n14762), .C2(n12314), .ZN(n12556) );
  MUX2_X1 U14587 ( .A(P3_REG2_REG_27__SCAN_IN), .B(n12556), .S(n14791), .Z(
        n12317) );
  INV_X1 U14588 ( .A(n12317), .ZN(n12320) );
  AOI22_X1 U14589 ( .A1(n12497), .A2(n6433), .B1(n14772), .B2(n12318), .ZN(
        n12319) );
  OAI211_X1 U14590 ( .C1(n12493), .C2(n12557), .A(n12320), .B(n12319), .ZN(
        P3_U3206) );
  XNOR2_X1 U14591 ( .A(n12322), .B(n12321), .ZN(n12324) );
  AOI21_X1 U14592 ( .B1(n12324), .B2(n14778), .A(n12323), .ZN(n12503) );
  XNOR2_X1 U14593 ( .A(n12326), .B(n12325), .ZN(n12501) );
  INV_X1 U14594 ( .A(n12327), .ZN(n12328) );
  AOI22_X1 U14595 ( .A1(n14793), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n14772), 
        .B2(n12328), .ZN(n12329) );
  OAI21_X1 U14596 ( .B1(n12330), .B2(n12355), .A(n12329), .ZN(n12331) );
  AOI21_X1 U14597 ( .B1(n12501), .B2(n14737), .A(n12331), .ZN(n12332) );
  OAI21_X1 U14598 ( .B1(n12503), .B2(n14793), .A(n12332), .ZN(P3_U3207) );
  AOI21_X1 U14599 ( .B1(n12333), .B2(n12335), .A(n6536), .ZN(n12563) );
  INV_X1 U14600 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12340) );
  OAI211_X1 U14601 ( .C1(n12336), .C2(n12335), .A(n12334), .B(n14778), .ZN(
        n12338) );
  NAND2_X1 U14602 ( .A1(n12338), .A2(n12337), .ZN(n12561) );
  INV_X1 U14603 ( .A(n12561), .ZN(n12339) );
  MUX2_X1 U14604 ( .A(n12340), .B(n12339), .S(n14791), .Z(n12345) );
  INV_X1 U14605 ( .A(n12341), .ZN(n12342) );
  AOI22_X1 U14606 ( .A1(n12343), .A2(n6433), .B1(n14772), .B2(n12342), .ZN(
        n12344) );
  OAI211_X1 U14607 ( .C1(n12493), .C2(n12563), .A(n12345), .B(n12344), .ZN(
        P3_U3208) );
  XNOR2_X1 U14608 ( .A(n12346), .B(n12350), .ZN(n12349) );
  INV_X1 U14609 ( .A(n12347), .ZN(n12348) );
  OAI21_X1 U14610 ( .B1(n12349), .B2(n12418), .A(n12348), .ZN(n12506) );
  INV_X1 U14611 ( .A(n12506), .ZN(n12358) );
  XNOR2_X1 U14612 ( .A(n12351), .B(n12350), .ZN(n12507) );
  INV_X1 U14613 ( .A(n12352), .ZN(n12353) );
  AOI22_X1 U14614 ( .A1(n14793), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n14772), 
        .B2(n12353), .ZN(n12354) );
  OAI21_X1 U14615 ( .B1(n12569), .B2(n12355), .A(n12354), .ZN(n12356) );
  AOI21_X1 U14616 ( .B1(n12507), .B2(n14737), .A(n12356), .ZN(n12357) );
  OAI21_X1 U14617 ( .B1(n12358), .B2(n14793), .A(n12357), .ZN(P3_U3209) );
  XNOR2_X1 U14618 ( .A(n12359), .B(n12360), .ZN(n12575) );
  INV_X1 U14619 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12365) );
  XNOR2_X1 U14620 ( .A(n12361), .B(n12360), .ZN(n12364) );
  AOI222_X1 U14621 ( .A1(n14778), .A2(n12364), .B1(n12363), .B2(n14731), .C1(
        n12362), .C2(n14730), .ZN(n12570) );
  MUX2_X1 U14622 ( .A(n12365), .B(n12570), .S(n14791), .Z(n12368) );
  AOI22_X1 U14623 ( .A1(n12572), .A2(n6433), .B1(n14772), .B2(n12366), .ZN(
        n12367) );
  OAI211_X1 U14624 ( .C1(n12493), .C2(n12575), .A(n12368), .B(n12367), .ZN(
        P3_U3210) );
  XOR2_X1 U14625 ( .A(n12371), .B(n12369), .Z(n12581) );
  INV_X1 U14626 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12374) );
  XOR2_X1 U14627 ( .A(n12371), .B(n12370), .Z(n12373) );
  AOI21_X1 U14628 ( .B1(n12373), .B2(n14778), .A(n12372), .ZN(n12576) );
  MUX2_X1 U14629 ( .A(n12374), .B(n12576), .S(n14791), .Z(n12377) );
  AOI22_X1 U14630 ( .A1(n12578), .A2(n6433), .B1(n14772), .B2(n12375), .ZN(
        n12376) );
  OAI211_X1 U14631 ( .C1(n12493), .C2(n12581), .A(n12377), .B(n12376), .ZN(
        P3_U3211) );
  XNOR2_X1 U14632 ( .A(n12379), .B(n12378), .ZN(n12584) );
  INV_X1 U14633 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12386) );
  XNOR2_X1 U14634 ( .A(n12381), .B(n12380), .ZN(n12382) );
  OAI222_X1 U14635 ( .A1(n14760), .A2(n12384), .B1(n14762), .B2(n12383), .C1(
        n12382), .C2(n12418), .ZN(n12582) );
  INV_X1 U14636 ( .A(n12582), .ZN(n12385) );
  MUX2_X1 U14637 ( .A(n12386), .B(n12385), .S(n14791), .Z(n12390) );
  AOI22_X1 U14638 ( .A1(n12388), .A2(n6433), .B1(n14772), .B2(n12387), .ZN(
        n12389) );
  OAI211_X1 U14639 ( .C1(n12493), .C2(n12584), .A(n12390), .B(n12389), .ZN(
        P3_U3212) );
  XNOR2_X1 U14640 ( .A(n12392), .B(n12391), .ZN(n12589) );
  XNOR2_X1 U14641 ( .A(n12393), .B(n12394), .ZN(n12395) );
  OAI222_X1 U14642 ( .A1(n14760), .A2(n12396), .B1(n14762), .B2(n12420), .C1(
        n12418), .C2(n12395), .ZN(n12587) );
  INV_X1 U14643 ( .A(n12587), .ZN(n12397) );
  MUX2_X1 U14644 ( .A(n12398), .B(n12397), .S(n14791), .Z(n12402) );
  AOI22_X1 U14645 ( .A1(n12400), .A2(n6433), .B1(n14772), .B2(n12399), .ZN(
        n12401) );
  OAI211_X1 U14646 ( .C1(n12493), .C2(n12589), .A(n12402), .B(n12401), .ZN(
        P3_U3213) );
  XOR2_X1 U14647 ( .A(n12404), .B(n12403), .Z(n12594) );
  INV_X1 U14648 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12409) );
  XNOR2_X1 U14649 ( .A(n12405), .B(n12404), .ZN(n12407) );
  OAI21_X1 U14650 ( .B1(n12407), .B2(n12418), .A(n12406), .ZN(n12592) );
  INV_X1 U14651 ( .A(n12592), .ZN(n12408) );
  MUX2_X1 U14652 ( .A(n12409), .B(n12408), .S(n14791), .Z(n12413) );
  AOI22_X1 U14653 ( .A1(n12411), .A2(n6433), .B1(n14772), .B2(n12410), .ZN(
        n12412) );
  OAI211_X1 U14654 ( .C1(n12493), .C2(n12594), .A(n12413), .B(n12412), .ZN(
        P3_U3214) );
  AOI21_X1 U14655 ( .B1(n12422), .B2(n12416), .A(n12415), .ZN(n12417) );
  OAI222_X1 U14656 ( .A1(n14760), .A2(n12420), .B1(n14762), .B2(n12419), .C1(
        n12418), .C2(n12417), .ZN(n12524) );
  INV_X1 U14657 ( .A(n12524), .ZN(n12429) );
  OAI22_X1 U14658 ( .A1(n14791), .A2(n7723), .B1(n12421), .B2(n14785), .ZN(
        n12426) );
  NOR2_X1 U14659 ( .A1(n12423), .A2(n12422), .ZN(n12523) );
  INV_X1 U14660 ( .A(n12525), .ZN(n12424) );
  NOR3_X1 U14661 ( .A1(n12523), .A2(n12424), .A3(n12493), .ZN(n12425) );
  AOI211_X1 U14662 ( .C1(n6433), .C2(n12427), .A(n12426), .B(n12425), .ZN(
        n12428) );
  OAI21_X1 U14663 ( .B1(n12429), .B2(n14793), .A(n12428), .ZN(P3_U3215) );
  XOR2_X1 U14664 ( .A(n12432), .B(n12430), .Z(n12606) );
  XOR2_X1 U14665 ( .A(n12432), .B(n12431), .Z(n12435) );
  AOI222_X1 U14666 ( .A1(n14778), .A2(n12435), .B1(n12434), .B2(n14730), .C1(
        n12433), .C2(n14731), .ZN(n12601) );
  MUX2_X1 U14667 ( .A(n14931), .B(n12601), .S(n14791), .Z(n12439) );
  INV_X1 U14668 ( .A(n12436), .ZN(n12437) );
  AOI22_X1 U14669 ( .A1(n12603), .A2(n6433), .B1(n12437), .B2(n14772), .ZN(
        n12438) );
  OAI211_X1 U14670 ( .C1(n12493), .C2(n12606), .A(n12439), .B(n12438), .ZN(
        P3_U3216) );
  OAI21_X1 U14671 ( .B1(n12441), .B2(n12443), .A(n12440), .ZN(n12442) );
  INV_X1 U14672 ( .A(n12442), .ZN(n12612) );
  XNOR2_X1 U14673 ( .A(n12444), .B(n12443), .ZN(n12446) );
  AOI21_X1 U14674 ( .B1(n12446), .B2(n14778), .A(n12445), .ZN(n12607) );
  MUX2_X1 U14675 ( .A(n12447), .B(n12607), .S(n14791), .Z(n12450) );
  AOI22_X1 U14676 ( .A1(n12609), .A2(n6433), .B1(n14772), .B2(n12448), .ZN(
        n12449) );
  OAI211_X1 U14677 ( .C1(n12493), .C2(n12612), .A(n12450), .B(n12449), .ZN(
        P3_U3217) );
  XNOR2_X1 U14678 ( .A(n12452), .B(n12451), .ZN(n12619) );
  OAI211_X1 U14679 ( .C1(n12455), .C2(n12454), .A(n12453), .B(n14778), .ZN(
        n12458) );
  INV_X1 U14680 ( .A(n12456), .ZN(n12457) );
  AND2_X1 U14681 ( .A1(n12458), .A2(n12457), .ZN(n12613) );
  MUX2_X1 U14682 ( .A(n12459), .B(n12613), .S(n14791), .Z(n12463) );
  INV_X1 U14683 ( .A(n12460), .ZN(n12461) );
  AOI22_X1 U14684 ( .A1(n12616), .A2(n6433), .B1(n14772), .B2(n12461), .ZN(
        n12462) );
  OAI211_X1 U14685 ( .C1(n12493), .C2(n12619), .A(n12463), .B(n12462), .ZN(
        P3_U3218) );
  OR2_X1 U14686 ( .A1(n12465), .A2(n12464), .ZN(n12466) );
  NAND3_X1 U14687 ( .A1(n12467), .A2(n14778), .A3(n12466), .ZN(n12472) );
  OAI22_X1 U14688 ( .A1(n12469), .A2(n14762), .B1(n12468), .B2(n14760), .ZN(
        n12470) );
  INV_X1 U14689 ( .A(n12470), .ZN(n12471) );
  NAND2_X1 U14690 ( .A1(n12472), .A2(n12471), .ZN(n12620) );
  MUX2_X1 U14691 ( .A(n12620), .B(P3_REG2_REG_14__SCAN_IN), .S(n14793), .Z(
        n12473) );
  INV_X1 U14692 ( .A(n12473), .ZN(n12481) );
  XNOR2_X1 U14693 ( .A(n12475), .B(n12474), .ZN(n12625) );
  NAND2_X1 U14694 ( .A1(n6433), .A2(n12476), .ZN(n12477) );
  OAI21_X1 U14695 ( .B1(n12478), .B2(n14785), .A(n12477), .ZN(n12479) );
  AOI21_X1 U14696 ( .B1(n12625), .B2(n14737), .A(n12479), .ZN(n12480) );
  NAND2_X1 U14697 ( .A1(n12481), .A2(n12480), .ZN(P3_U3219) );
  XOR2_X1 U14698 ( .A(n12484), .B(n12482), .Z(n12631) );
  INV_X1 U14699 ( .A(n12631), .ZN(n12492) );
  XOR2_X1 U14700 ( .A(n12484), .B(n12483), .Z(n12486) );
  AOI21_X1 U14701 ( .B1(n12486), .B2(n14778), .A(n12485), .ZN(n12629) );
  MUX2_X1 U14702 ( .A(n12629), .B(n14910), .S(n14793), .Z(n12491) );
  INV_X1 U14703 ( .A(n12634), .ZN(n12489) );
  INV_X1 U14704 ( .A(n12487), .ZN(n12488) );
  AOI22_X1 U14705 ( .A1(n6433), .A2(n12489), .B1(n14772), .B2(n12488), .ZN(
        n12490) );
  OAI211_X1 U14706 ( .C1(n12493), .C2(n12492), .A(n12491), .B(n12490), .ZN(
        P3_U3220) );
  INV_X1 U14707 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12494) );
  MUX2_X1 U14708 ( .A(n12494), .B(n12550), .S(n14868), .Z(n12496) );
  NAND2_X1 U14709 ( .A1(n12552), .A2(n12536), .ZN(n12495) );
  OAI211_X1 U14710 ( .C1(n12540), .C2(n12555), .A(n12496), .B(n12495), .ZN(
        P3_U3487) );
  MUX2_X1 U14711 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n12556), .S(n14868), .Z(
        n12499) );
  OAI22_X1 U14712 ( .A1(n12557), .A2(n12540), .B1(n8902), .B2(n12548), .ZN(
        n12498) );
  OR2_X1 U14713 ( .A1(n12499), .A2(n12498), .ZN(P3_U3486) );
  AOI22_X1 U14714 ( .A1(n12501), .A2(n14848), .B1(n14821), .B2(n12500), .ZN(
        n12502) );
  NAND2_X1 U14715 ( .A1(n12503), .A2(n12502), .ZN(n12560) );
  MUX2_X1 U14716 ( .A(P3_REG1_REG_26__SCAN_IN), .B(n12560), .S(n14868), .Z(
        P3_U3485) );
  MUX2_X1 U14717 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12561), .S(n14868), .Z(
        n12505) );
  OAI22_X1 U14718 ( .A1(n12563), .A2(n12540), .B1(n12562), .B2(n12548), .ZN(
        n12504) );
  OR2_X1 U14719 ( .A1(n12505), .A2(n12504), .ZN(P3_U3484) );
  INV_X1 U14720 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n12508) );
  AOI21_X1 U14721 ( .B1(n14848), .B2(n12507), .A(n12506), .ZN(n12566) );
  MUX2_X1 U14722 ( .A(n12508), .B(n12566), .S(n14868), .Z(n12509) );
  OAI21_X1 U14723 ( .B1(n12569), .B2(n12548), .A(n12509), .ZN(P3_U3483) );
  INV_X1 U14724 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12510) );
  MUX2_X1 U14725 ( .A(n12510), .B(n12570), .S(n14868), .Z(n12512) );
  NAND2_X1 U14726 ( .A1(n12572), .A2(n12536), .ZN(n12511) );
  OAI211_X1 U14727 ( .C1(n12540), .C2(n12575), .A(n12512), .B(n12511), .ZN(
        P3_U3482) );
  INV_X1 U14728 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12513) );
  MUX2_X1 U14729 ( .A(n12513), .B(n12576), .S(n14868), .Z(n12515) );
  NAND2_X1 U14730 ( .A1(n12578), .A2(n12536), .ZN(n12514) );
  OAI211_X1 U14731 ( .C1(n12540), .C2(n12581), .A(n12515), .B(n12514), .ZN(
        P3_U3481) );
  MUX2_X1 U14732 ( .A(P3_REG1_REG_21__SCAN_IN), .B(n12582), .S(n14868), .Z(
        n12517) );
  OAI22_X1 U14733 ( .A1(n12584), .A2(n12540), .B1(n12583), .B2(n12548), .ZN(
        n12516) );
  OR2_X1 U14734 ( .A1(n12517), .A2(n12516), .ZN(P3_U3480) );
  MUX2_X1 U14735 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12587), .S(n14868), .Z(
        n12519) );
  OAI22_X1 U14736 ( .A1(n12589), .A2(n12540), .B1(n12588), .B2(n12548), .ZN(
        n12518) );
  OR2_X1 U14737 ( .A1(n12519), .A2(n12518), .ZN(P3_U3479) );
  MUX2_X1 U14738 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12592), .S(n14868), .Z(
        n12521) );
  OAI22_X1 U14739 ( .A1(n12594), .A2(n12540), .B1(n12593), .B2(n12548), .ZN(
        n12520) );
  OR2_X1 U14740 ( .A1(n12521), .A2(n12520), .ZN(P3_U3478) );
  INV_X1 U14741 ( .A(n14848), .ZN(n12522) );
  NOR2_X1 U14742 ( .A1(n12523), .A2(n12522), .ZN(n12526) );
  AOI21_X1 U14743 ( .B1(n12526), .B2(n12525), .A(n12524), .ZN(n12597) );
  MUX2_X1 U14744 ( .A(n12527), .B(n12597), .S(n14868), .Z(n12528) );
  OAI21_X1 U14745 ( .B1(n12600), .B2(n12548), .A(n12528), .ZN(P3_U3477) );
  INV_X1 U14746 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12529) );
  MUX2_X1 U14747 ( .A(n12529), .B(n12601), .S(n14868), .Z(n12531) );
  NAND2_X1 U14748 ( .A1(n12603), .A2(n12536), .ZN(n12530) );
  OAI211_X1 U14749 ( .C1(n12540), .C2(n12606), .A(n12531), .B(n12530), .ZN(
        P3_U3476) );
  MUX2_X1 U14750 ( .A(n12532), .B(n12607), .S(n14868), .Z(n12534) );
  NAND2_X1 U14751 ( .A1(n12609), .A2(n12536), .ZN(n12533) );
  OAI211_X1 U14752 ( .C1(n12612), .C2(n12540), .A(n12534), .B(n12533), .ZN(
        P3_U3475) );
  INV_X1 U14753 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12535) );
  MUX2_X1 U14754 ( .A(n12535), .B(n12613), .S(n14868), .Z(n12538) );
  NAND2_X1 U14755 ( .A1(n12616), .A2(n12536), .ZN(n12537) );
  OAI211_X1 U14756 ( .C1(n12619), .C2(n12540), .A(n12538), .B(n12537), .ZN(
        P3_U3474) );
  INV_X1 U14757 ( .A(n14868), .ZN(n14866) );
  MUX2_X1 U14758 ( .A(n12620), .B(P3_REG1_REG_14__SCAN_IN), .S(n14866), .Z(
        n12539) );
  INV_X1 U14759 ( .A(n12539), .ZN(n12543) );
  INV_X1 U14760 ( .A(n12540), .ZN(n12545) );
  NOR2_X1 U14761 ( .A1(n12623), .A2(n12548), .ZN(n12541) );
  AOI21_X1 U14762 ( .B1(n12625), .B2(n12545), .A(n12541), .ZN(n12542) );
  NAND2_X1 U14763 ( .A1(n12543), .A2(n12542), .ZN(P3_U3473) );
  INV_X1 U14764 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n12544) );
  MUX2_X1 U14765 ( .A(n12629), .B(n12544), .S(n14866), .Z(n12547) );
  NAND2_X1 U14766 ( .A1(n12631), .A2(n12545), .ZN(n12546) );
  OAI211_X1 U14767 ( .C1(n12548), .C2(n12634), .A(n12547), .B(n12546), .ZN(
        P3_U3472) );
  MUX2_X1 U14768 ( .A(P3_REG1_REG_0__SCAN_IN), .B(n12549), .S(n14868), .Z(
        P3_U3459) );
  INV_X1 U14769 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12551) );
  MUX2_X1 U14770 ( .A(n12551), .B(n12550), .S(n14851), .Z(n12554) );
  INV_X1 U14771 ( .A(n12635), .ZN(n12615) );
  NAND2_X1 U14772 ( .A1(n12552), .A2(n12615), .ZN(n12553) );
  OAI211_X1 U14773 ( .C1(n12555), .C2(n12622), .A(n12554), .B(n12553), .ZN(
        P3_U3455) );
  MUX2_X1 U14774 ( .A(P3_REG0_REG_27__SCAN_IN), .B(n12556), .S(n14851), .Z(
        n12559) );
  OAI22_X1 U14775 ( .A1(n12557), .A2(n12622), .B1(n8902), .B2(n12635), .ZN(
        n12558) );
  OR2_X1 U14776 ( .A1(n12559), .A2(n12558), .ZN(P3_U3454) );
  MUX2_X1 U14777 ( .A(P3_REG0_REG_26__SCAN_IN), .B(n12560), .S(n14851), .Z(
        P3_U3453) );
  MUX2_X1 U14778 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12561), .S(n14851), .Z(
        n12565) );
  OAI22_X1 U14779 ( .A1(n12563), .A2(n12622), .B1(n12562), .B2(n12635), .ZN(
        n12564) );
  OR2_X1 U14780 ( .A1(n12565), .A2(n12564), .ZN(P3_U3452) );
  INV_X1 U14781 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n12567) );
  MUX2_X1 U14782 ( .A(n12567), .B(n12566), .S(n14851), .Z(n12568) );
  OAI21_X1 U14783 ( .B1(n12569), .B2(n12635), .A(n12568), .ZN(P3_U3451) );
  INV_X1 U14784 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12571) );
  MUX2_X1 U14785 ( .A(n12571), .B(n12570), .S(n14851), .Z(n12574) );
  NAND2_X1 U14786 ( .A1(n12572), .A2(n12615), .ZN(n12573) );
  OAI211_X1 U14787 ( .C1(n12575), .C2(n12622), .A(n12574), .B(n12573), .ZN(
        P3_U3450) );
  INV_X1 U14788 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12577) );
  MUX2_X1 U14789 ( .A(n12577), .B(n12576), .S(n14851), .Z(n12580) );
  NAND2_X1 U14790 ( .A1(n12578), .A2(n12615), .ZN(n12579) );
  OAI211_X1 U14791 ( .C1(n12581), .C2(n12622), .A(n12580), .B(n12579), .ZN(
        P3_U3449) );
  MUX2_X1 U14792 ( .A(P3_REG0_REG_21__SCAN_IN), .B(n12582), .S(n14851), .Z(
        n12586) );
  OAI22_X1 U14793 ( .A1(n12584), .A2(n12622), .B1(n12583), .B2(n12635), .ZN(
        n12585) );
  OR2_X1 U14794 ( .A1(n12586), .A2(n12585), .ZN(P3_U3448) );
  MUX2_X1 U14795 ( .A(P3_REG0_REG_20__SCAN_IN), .B(n12587), .S(n14851), .Z(
        n12591) );
  OAI22_X1 U14796 ( .A1(n12589), .A2(n12622), .B1(n12588), .B2(n12635), .ZN(
        n12590) );
  OR2_X1 U14797 ( .A1(n12591), .A2(n12590), .ZN(P3_U3447) );
  MUX2_X1 U14798 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12592), .S(n14851), .Z(
        n12596) );
  OAI22_X1 U14799 ( .A1(n12594), .A2(n12622), .B1(n12593), .B2(n12635), .ZN(
        n12595) );
  OR2_X1 U14800 ( .A1(n12596), .A2(n12595), .ZN(P3_U3446) );
  INV_X1 U14801 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12598) );
  MUX2_X1 U14802 ( .A(n12598), .B(n12597), .S(n14851), .Z(n12599) );
  OAI21_X1 U14803 ( .B1(n12600), .B2(n12635), .A(n12599), .ZN(P3_U3444) );
  INV_X1 U14804 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12602) );
  MUX2_X1 U14805 ( .A(n12602), .B(n12601), .S(n14851), .Z(n12605) );
  NAND2_X1 U14806 ( .A1(n12603), .A2(n12615), .ZN(n12604) );
  OAI211_X1 U14807 ( .C1(n12606), .C2(n12622), .A(n12605), .B(n12604), .ZN(
        P3_U3441) );
  INV_X1 U14808 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12608) );
  MUX2_X1 U14809 ( .A(n12608), .B(n12607), .S(n14851), .Z(n12611) );
  NAND2_X1 U14810 ( .A1(n12609), .A2(n12615), .ZN(n12610) );
  OAI211_X1 U14811 ( .C1(n12612), .C2(n12622), .A(n12611), .B(n12610), .ZN(
        P3_U3438) );
  INV_X1 U14812 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12614) );
  MUX2_X1 U14813 ( .A(n12614), .B(n12613), .S(n14851), .Z(n12618) );
  NAND2_X1 U14814 ( .A1(n12616), .A2(n12615), .ZN(n12617) );
  OAI211_X1 U14815 ( .C1(n12619), .C2(n12622), .A(n12618), .B(n12617), .ZN(
        P3_U3435) );
  MUX2_X1 U14816 ( .A(n12620), .B(P3_REG0_REG_14__SCAN_IN), .S(n14849), .Z(
        n12621) );
  INV_X1 U14817 ( .A(n12621), .ZN(n12627) );
  INV_X1 U14818 ( .A(n12622), .ZN(n12630) );
  NOR2_X1 U14819 ( .A1(n12635), .A2(n12623), .ZN(n12624) );
  AOI21_X1 U14820 ( .B1(n12625), .B2(n12630), .A(n12624), .ZN(n12626) );
  NAND2_X1 U14821 ( .A1(n12627), .A2(n12626), .ZN(P3_U3432) );
  INV_X1 U14822 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n12628) );
  MUX2_X1 U14823 ( .A(n12629), .B(n12628), .S(n14849), .Z(n12633) );
  NAND2_X1 U14824 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  OAI211_X1 U14825 ( .C1(n12635), .C2(n12634), .A(n12633), .B(n12632), .ZN(
        P3_U3429) );
  MUX2_X1 U14826 ( .A(P3_D_REG_1__SCAN_IN), .B(n12637), .S(n12636), .Z(
        P3_U3377) );
  NAND2_X1 U14827 ( .A1(n12638), .A2(n13948), .ZN(n12641) );
  OR4_X1 U14828 ( .A1(n12639), .A2(P3_IR_REG_30__SCAN_IN), .A3(P3_U3151), .A4(
        n7646), .ZN(n12640) );
  OAI211_X1 U14829 ( .C1(n12661), .C2(n12642), .A(n12641), .B(n12640), .ZN(
        P3_U3264) );
  INV_X1 U14830 ( .A(n12643), .ZN(n12644) );
  OAI222_X1 U14831 ( .A1(P3_U3151), .A2(n12646), .B1(n12661), .B2(n12645), 
        .C1(n12657), .C2(n12644), .ZN(P3_U3265) );
  INV_X1 U14832 ( .A(n12647), .ZN(n12649) );
  OAI222_X1 U14833 ( .A1(n12661), .A2(n12650), .B1(n12664), .B2(n12649), .C1(
        P3_U3151), .C2(n12648), .ZN(P3_U3266) );
  INV_X1 U14834 ( .A(n12651), .ZN(n12652) );
  OAI222_X1 U14835 ( .A1(P3_U3151), .A2(n12654), .B1(n12661), .B2(n12653), 
        .C1(n12657), .C2(n12652), .ZN(P3_U3267) );
  INV_X1 U14836 ( .A(n12655), .ZN(n12656) );
  OAI222_X1 U14837 ( .A1(P3_U3151), .A2(n12659), .B1(n12661), .B2(n12658), 
        .C1(n12657), .C2(n12656), .ZN(P3_U3268) );
  INV_X1 U14838 ( .A(n12660), .ZN(n12663) );
  OAI222_X1 U14839 ( .A1(P3_U3151), .A2(n12665), .B1(n12664), .B2(n12663), 
        .C1(n12662), .C2(n12661), .ZN(P3_U3269) );
  MUX2_X1 U14840 ( .A(n12666), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AOI22_X1 U14841 ( .A1(n12882), .A2(n12754), .B1(n12824), .B2(n12884), .ZN(
        n12904) );
  OAI22_X1 U14842 ( .A1(n12744), .A2(n12904), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12670), .ZN(n12671) );
  AOI21_X1 U14843 ( .B1(n12909), .B2(n12758), .A(n12671), .ZN(n12672) );
  OAI211_X1 U14844 ( .C1(n12911), .C2(n12761), .A(n12673), .B(n12672), .ZN(
        P2_U3186) );
  INV_X1 U14845 ( .A(n13116), .ZN(n12970) );
  OAI211_X1 U14846 ( .C1(n12674), .C2(n12676), .A(n12675), .B(n12763), .ZN(
        n12681) );
  AOI22_X1 U14847 ( .A1(n12754), .A2(n12874), .B1(n12878), .B2(n12824), .ZN(
        n12963) );
  INV_X1 U14848 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n12677) );
  OAI22_X1 U14849 ( .A1(n12744), .A2(n12963), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12677), .ZN(n12678) );
  AOI21_X1 U14850 ( .B1(n12679), .B2(n12758), .A(n12678), .ZN(n12680) );
  OAI211_X1 U14851 ( .C1(n12970), .C2(n12761), .A(n12681), .B(n12680), .ZN(
        P2_U3188) );
  OAI21_X1 U14852 ( .B1(n12684), .B2(n12683), .A(n6952), .ZN(n12685) );
  NAND2_X1 U14853 ( .A1(n12685), .A2(n12763), .ZN(n12690) );
  NAND2_X1 U14854 ( .A1(n12869), .A2(n12824), .ZN(n12687) );
  NAND2_X1 U14855 ( .A1(n12864), .A2(n12754), .ZN(n12686) );
  NAND2_X1 U14856 ( .A1(n12687), .A2(n12686), .ZN(n13019) );
  AND2_X1 U14857 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12820) );
  NOR2_X1 U14858 ( .A1(n12742), .A2(n13023), .ZN(n12688) );
  AOI211_X1 U14859 ( .C1(n12757), .C2(n13019), .A(n12820), .B(n12688), .ZN(
        n12689) );
  OAI211_X1 U14860 ( .C1(n7072), .C2(n12761), .A(n12690), .B(n12689), .ZN(
        P2_U3191) );
  OAI211_X1 U14861 ( .C1(n12693), .C2(n12692), .A(n12691), .B(n12763), .ZN(
        n12697) );
  AOI22_X1 U14862 ( .A1(n12869), .A2(n12754), .B1(n12824), .B2(n12874), .ZN(
        n12990) );
  INV_X1 U14863 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n12694) );
  OAI22_X1 U14864 ( .A1(n12990), .A2(n12744), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12694), .ZN(n12695) );
  AOI21_X1 U14865 ( .B1(n12996), .B2(n12758), .A(n12695), .ZN(n12696) );
  OAI211_X1 U14866 ( .C1(n12998), .C2(n12761), .A(n12697), .B(n12696), .ZN(
        P2_U3195) );
  OAI21_X1 U14867 ( .B1(n12699), .B2(n12698), .A(n12763), .ZN(n12707) );
  INV_X1 U14868 ( .A(n12934), .ZN(n12703) );
  OR2_X1 U14869 ( .A1(n12881), .A2(n12756), .ZN(n12700) );
  OAI21_X1 U14870 ( .B1(n12701), .B2(n12848), .A(n12700), .ZN(n12932) );
  AOI22_X1 U14871 ( .A1(n12757), .A2(n12932), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12702) );
  OAI21_X1 U14872 ( .B1(n12703), .B2(n12742), .A(n12702), .ZN(n12704) );
  AOI21_X1 U14873 ( .B1(n13105), .B2(n12747), .A(n12704), .ZN(n12705) );
  OAI21_X1 U14874 ( .B1(n12707), .B2(n12706), .A(n12705), .ZN(P2_U3197) );
  AOI21_X1 U14875 ( .B1(n12710), .B2(n12709), .A(n12708), .ZN(n12714) );
  INV_X1 U14876 ( .A(n12860), .ZN(n12835) );
  OAI22_X1 U14877 ( .A1(n12837), .A2(n12756), .B1(n12835), .B2(n12848), .ZN(
        n13049) );
  NAND2_X1 U14878 ( .A1(n13049), .A2(n12757), .ZN(n12711) );
  NAND2_X1 U14879 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14538)
         );
  OAI211_X1 U14880 ( .C1(n12742), .C2(n13054), .A(n12711), .B(n14538), .ZN(
        n12712) );
  AOI21_X1 U14881 ( .B1(n13146), .B2(n12747), .A(n12712), .ZN(n12713) );
  OAI21_X1 U14882 ( .B1(n12714), .B2(n12749), .A(n12713), .ZN(P2_U3200) );
  OAI211_X1 U14883 ( .C1(n12717), .C2(n12716), .A(n12715), .B(n12763), .ZN(
        n12721) );
  AOI22_X1 U14884 ( .A1(n12754), .A2(n12877), .B1(n12880), .B2(n12824), .ZN(
        n12945) );
  OAI22_X1 U14885 ( .A1(n12744), .A2(n12945), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12718), .ZN(n12719) );
  AOI21_X1 U14886 ( .B1(n12954), .B2(n12758), .A(n12719), .ZN(n12720) );
  OAI211_X1 U14887 ( .C1(n13110), .C2(n12761), .A(n12721), .B(n12720), .ZN(
        P2_U3201) );
  INV_X1 U14888 ( .A(n12722), .ZN(n12724) );
  NAND2_X1 U14889 ( .A1(n12724), .A2(n12723), .ZN(n12725) );
  XNOR2_X1 U14890 ( .A(n12726), .B(n12725), .ZN(n12731) );
  INV_X1 U14891 ( .A(n12867), .ZN(n12727) );
  OAI22_X1 U14892 ( .A1(n12840), .A2(n12756), .B1(n12727), .B2(n12848), .ZN(
        n13005) );
  AOI22_X1 U14893 ( .A1(n13005), .A2(n12757), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12728) );
  OAI21_X1 U14894 ( .B1(n13008), .B2(n12742), .A(n12728), .ZN(n12729) );
  AOI21_X1 U14895 ( .B1(n13131), .B2(n12747), .A(n12729), .ZN(n12730) );
  OAI21_X1 U14896 ( .B1(n12731), .B2(n12749), .A(n12730), .ZN(P2_U3205) );
  AOI211_X1 U14897 ( .C1(n12734), .C2(n12733), .A(n12749), .B(n12732), .ZN(
        n12735) );
  INV_X1 U14898 ( .A(n12735), .ZN(n12739) );
  AOI22_X1 U14899 ( .A1(n12872), .A2(n12754), .B1(n12824), .B2(n12877), .ZN(
        n12975) );
  OAI22_X1 U14900 ( .A1(n12975), .A2(n12744), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12736), .ZN(n12737) );
  AOI21_X1 U14901 ( .B1(n12979), .B2(n12758), .A(n12737), .ZN(n12738) );
  OAI211_X1 U14902 ( .C1(n12981), .C2(n12761), .A(n12739), .B(n12738), .ZN(
        P2_U3207) );
  XNOR2_X1 U14903 ( .A(n12741), .B(n12740), .ZN(n12750) );
  NOR2_X1 U14904 ( .A1(n12742), .A2(n13037), .ZN(n12746) );
  AOI22_X1 U14905 ( .A1(n12867), .A2(n12824), .B1(n12754), .B2(n12863), .ZN(
        n13033) );
  NAND2_X1 U14906 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n12794)
         );
  OAI21_X1 U14907 ( .B1(n13033), .B2(n12744), .A(n12794), .ZN(n12745) );
  AOI211_X1 U14908 ( .C1(n13141), .C2(n12747), .A(n12746), .B(n12745), .ZN(
        n12748) );
  OAI21_X1 U14909 ( .B1(n12750), .B2(n12749), .A(n12748), .ZN(P2_U3210) );
  OAI21_X1 U14910 ( .B1(n12753), .B2(n12752), .A(n12751), .ZN(n12764) );
  NAND2_X1 U14911 ( .A1(n12880), .A2(n12754), .ZN(n12755) );
  OAI21_X1 U14912 ( .B1(n12883), .B2(n12756), .A(n12755), .ZN(n12918) );
  AOI22_X1 U14913 ( .A1(n12757), .A2(n12918), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12760) );
  NAND2_X1 U14914 ( .A1(n12758), .A2(n12922), .ZN(n12759) );
  OAI211_X1 U14915 ( .C1(n12924), .C2(n12761), .A(n12760), .B(n12759), .ZN(
        n12762) );
  AOI21_X1 U14916 ( .B1(n12764), .B2(n12763), .A(n12762), .ZN(n12765) );
  INV_X1 U14917 ( .A(n12765), .ZN(P2_U3212) );
  MUX2_X1 U14918 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n12766), .S(n12783), .Z(
        P2_U3562) );
  MUX2_X1 U14919 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n12767), .S(n12783), .Z(
        P2_U3561) );
  MUX2_X1 U14920 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12768), .S(n12783), .Z(
        P2_U3560) );
  MUX2_X1 U14921 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n12884), .S(n12783), .Z(
        P2_U3559) );
  MUX2_X1 U14922 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n12769), .S(n12783), .Z(
        P2_U3558) );
  MUX2_X1 U14923 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n12882), .S(n12783), .Z(
        P2_U3557) );
  MUX2_X1 U14924 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n12880), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U14925 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n12878), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U14926 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n12877), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U14927 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n12874), .S(P2_U3947), .Z(
        P2_U3553) );
  MUX2_X1 U14928 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n12872), .S(P2_U3947), .Z(
        P2_U3552) );
  MUX2_X1 U14929 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n12869), .S(P2_U3947), .Z(
        P2_U3551) );
  MUX2_X1 U14930 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n12867), .S(P2_U3947), .Z(
        P2_U3550) );
  MUX2_X1 U14931 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n12864), .S(n12783), .Z(
        P2_U3549) );
  MUX2_X1 U14932 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n12863), .S(n12783), .Z(
        P2_U3548) );
  MUX2_X1 U14933 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n12860), .S(n12783), .Z(
        P2_U3547) );
  MUX2_X1 U14934 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n12856), .S(n12783), .Z(
        P2_U3546) );
  MUX2_X1 U14935 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n12770), .S(n12783), .Z(
        P2_U3545) );
  MUX2_X1 U14936 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n12771), .S(n12783), .Z(
        P2_U3544) );
  MUX2_X1 U14937 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n12772), .S(n12783), .Z(
        P2_U3543) );
  MUX2_X1 U14938 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n12773), .S(n12783), .Z(
        P2_U3542) );
  MUX2_X1 U14939 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n12774), .S(n12783), .Z(
        P2_U3541) );
  MUX2_X1 U14940 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n12775), .S(n12783), .Z(
        P2_U3540) );
  MUX2_X1 U14941 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n12776), .S(n12783), .Z(
        P2_U3539) );
  MUX2_X1 U14942 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n12777), .S(n12783), .Z(
        P2_U3538) );
  MUX2_X1 U14943 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n12778), .S(n12783), .Z(
        P2_U3537) );
  MUX2_X1 U14944 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n12779), .S(n12783), .Z(
        P2_U3536) );
  MUX2_X1 U14945 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n12780), .S(n12783), .Z(
        P2_U3535) );
  MUX2_X1 U14946 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n12781), .S(n12783), .Z(
        P2_U3534) );
  MUX2_X1 U14947 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n12782), .S(n12783), .Z(
        P2_U3533) );
  MUX2_X1 U14948 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n11293), .S(n12783), .Z(
        P2_U3532) );
  MUX2_X1 U14949 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n11289), .S(n12783), .Z(
        P2_U3531) );
  NOR2_X1 U14950 ( .A1(n12785), .A2(n12786), .ZN(n12787) );
  NOR2_X1 U14951 ( .A1(n12788), .A2(n14501), .ZN(n12789) );
  INV_X1 U14952 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n14506) );
  XNOR2_X1 U14953 ( .A(n12788), .B(n14501), .ZN(n14507) );
  NOR2_X1 U14954 ( .A1(n14506), .A2(n14507), .ZN(n14505) );
  XNOR2_X1 U14955 ( .A(n14522), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n14518) );
  XNOR2_X1 U14956 ( .A(n14536), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n14528) );
  INV_X1 U14957 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n12791) );
  NAND2_X1 U14958 ( .A1(n12792), .A2(n12791), .ZN(n12807) );
  OAI21_X1 U14959 ( .B1(n12792), .B2(n12791), .A(n12807), .ZN(n12793) );
  INV_X1 U14960 ( .A(n12793), .ZN(n12804) );
  OAI21_X1 U14961 ( .B1(n12815), .B2(n12809), .A(n12794), .ZN(n12802) );
  XNOR2_X1 U14962 ( .A(n14497), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n14493) );
  NOR2_X1 U14963 ( .A1(n12797), .A2(n14501), .ZN(n12798) );
  INV_X1 U14964 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14503) );
  XNOR2_X1 U14965 ( .A(n14522), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n14515) );
  XNOR2_X1 U14966 ( .A(n14536), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14532) );
  AOI211_X1 U14967 ( .C1(n12800), .C2(n12799), .A(n12811), .B(n14531), .ZN(
        n12801) );
  AOI211_X1 U14968 ( .C1(n14442), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n12802), 
        .B(n12801), .ZN(n12803) );
  OAI21_X1 U14969 ( .B1(n12804), .B2(n14527), .A(n12803), .ZN(P2_U3232) );
  NAND2_X1 U14970 ( .A1(n12805), .A2(n12809), .ZN(n12806) );
  NAND2_X1 U14971 ( .A1(n12807), .A2(n12806), .ZN(n12808) );
  XOR2_X1 U14972 ( .A(n12808), .B(P2_REG2_REG_19__SCAN_IN), .Z(n12818) );
  INV_X1 U14973 ( .A(n12818), .ZN(n12816) );
  NOR2_X1 U14974 ( .A1(n12810), .A2(n12809), .ZN(n12812) );
  XOR2_X1 U14975 ( .A(n12813), .B(P2_REG1_REG_19__SCAN_IN), .Z(n12817) );
  INV_X1 U14976 ( .A(n13146), .ZN(n13057) );
  NAND2_X1 U14977 ( .A1(n13074), .A2(n13057), .ZN(n13051) );
  XNOR2_X1 U14978 ( .A(n13083), .B(n12828), .ZN(n12821) );
  NAND2_X1 U14979 ( .A1(n12821), .A2(n12952), .ZN(n13082) );
  NAND2_X1 U14980 ( .A1(n12822), .A2(P2_B_REG_SCAN_IN), .ZN(n12823) );
  NAND2_X1 U14981 ( .A1(n12824), .A2(n12823), .ZN(n12846) );
  OR2_X1 U14982 ( .A1(n12825), .A2(n12846), .ZN(n13084) );
  NOR2_X1 U14983 ( .A1(n14557), .A2(n13084), .ZN(n12830) );
  NOR2_X1 U14984 ( .A1(n13083), .A2(n13076), .ZN(n12826) );
  AOI211_X1 U14985 ( .C1(n14557), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12830), 
        .B(n12826), .ZN(n12827) );
  OAI21_X1 U14986 ( .B1(n13082), .B2(n12953), .A(n12827), .ZN(P2_U3234) );
  OAI211_X1 U14987 ( .C1(n13086), .C2(n12852), .A(n12828), .B(n12952), .ZN(
        n13085) );
  NOR2_X1 U14988 ( .A1(n13086), .A2(n13076), .ZN(n12829) );
  AOI211_X1 U14989 ( .C1(n14557), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12830), 
        .B(n12829), .ZN(n12831) );
  OAI21_X1 U14990 ( .B1(n12953), .B2(n13085), .A(n12831), .ZN(P2_U3235) );
  INV_X1 U14991 ( .A(n12832), .ZN(n12858) );
  INV_X1 U14992 ( .A(n13066), .ZN(n12836) );
  INV_X1 U14993 ( .A(n13141), .ZN(n13040) );
  NAND2_X1 U14994 ( .A1(n13040), .A2(n12864), .ZN(n12838) );
  INV_X1 U14995 ( .A(n13026), .ZN(n13017) );
  NAND2_X1 U14996 ( .A1(n12970), .A2(n12877), .ZN(n12841) );
  INV_X1 U14997 ( .A(n12950), .ZN(n12842) );
  INV_X1 U14998 ( .A(n12938), .ZN(n12930) );
  XNOR2_X1 U14999 ( .A(n12845), .B(n12886), .ZN(n12851) );
  OAI22_X1 U15000 ( .A1(n12849), .A2(n12848), .B1(n12847), .B2(n12846), .ZN(
        n12850) );
  AOI21_X2 U15001 ( .B1(n12851), .B2(n14548), .A(n12850), .ZN(n13090) );
  INV_X1 U15002 ( .A(n13088), .ZN(n12855) );
  AOI22_X1 U15003 ( .A1(n14557), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n12853), 
        .B2(n14553), .ZN(n12854) );
  OAI21_X1 U15004 ( .B1(n12855), .B2(n13076), .A(n12854), .ZN(n12887) );
  NAND2_X1 U15005 ( .A1(n13151), .A2(n12860), .ZN(n12861) );
  INV_X1 U15006 ( .A(n13031), .ZN(n13042) );
  OR2_X1 U15007 ( .A1(n13141), .A2(n12864), .ZN(n12865) );
  NAND2_X1 U15008 ( .A1(n13136), .A2(n12867), .ZN(n12866) );
  OR2_X1 U15009 ( .A1(n13136), .A2(n12867), .ZN(n12868) );
  NOR2_X1 U15010 ( .A1(n13131), .A2(n12869), .ZN(n12870) );
  INV_X1 U15011 ( .A(n12999), .ZN(n12871) );
  OR2_X1 U15012 ( .A1(n13126), .A2(n12872), .ZN(n12873) );
  XNOR2_X1 U15013 ( .A(n12888), .B(n12889), .ZN(n13095) );
  AOI21_X1 U15014 ( .B1(n6530), .B2(n12889), .A(n12946), .ZN(n12892) );
  AOI21_X1 U15015 ( .B1(n12892), .B2(n12891), .A(n12890), .ZN(n13094) );
  OAI21_X1 U15016 ( .B1(n12893), .B2(n13071), .A(n13094), .ZN(n12894) );
  NAND2_X1 U15017 ( .A1(n12894), .A2(n14554), .ZN(n12902) );
  INV_X1 U15018 ( .A(n12908), .ZN(n12897) );
  INV_X1 U15019 ( .A(n12895), .ZN(n12896) );
  AOI211_X1 U15020 ( .C1(n7078), .C2(n12897), .A(n9339), .B(n12896), .ZN(
        n13092) );
  INV_X1 U15021 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n12898) );
  OAI22_X1 U15022 ( .A1(n12899), .A2(n13076), .B1(n14554), .B2(n12898), .ZN(
        n12900) );
  AOI21_X1 U15023 ( .B1(n13092), .B2(n13078), .A(n12900), .ZN(n12901) );
  OAI211_X1 U15024 ( .C1(n13081), .C2(n13095), .A(n12902), .B(n12901), .ZN(
        P2_U3237) );
  XNOR2_X1 U15025 ( .A(n12903), .B(n12912), .ZN(n12906) );
  INV_X1 U15026 ( .A(n12904), .ZN(n12905) );
  AOI21_X1 U15027 ( .B1(n12906), .B2(n14548), .A(n12905), .ZN(n13098) );
  NOR2_X1 U15028 ( .A1(n12911), .A2(n12921), .ZN(n12907) );
  AOI22_X1 U15029 ( .A1(n14557), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n12909), 
        .B2(n14553), .ZN(n12910) );
  OAI21_X1 U15030 ( .B1(n12911), .B2(n13076), .A(n12910), .ZN(n12915) );
  XNOR2_X1 U15031 ( .A(n12913), .B(n12912), .ZN(n13099) );
  NOR2_X1 U15032 ( .A1(n13099), .A2(n13081), .ZN(n12914) );
  AOI211_X1 U15033 ( .C1(n13078), .C2(n7590), .A(n12915), .B(n12914), .ZN(
        n12916) );
  OAI21_X1 U15034 ( .B1(n13098), .B2(n14557), .A(n12916), .ZN(P2_U3238) );
  XNOR2_X1 U15035 ( .A(n12917), .B(n12926), .ZN(n12919) );
  AOI21_X1 U15036 ( .B1(n12919), .B2(n14548), .A(n12918), .ZN(n13102) );
  NOR2_X1 U15037 ( .A1(n12924), .A2(n7602), .ZN(n12920) );
  AOI22_X1 U15038 ( .A1(n14557), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n12922), 
        .B2(n14553), .ZN(n12923) );
  OAI21_X1 U15039 ( .B1(n12924), .B2(n13076), .A(n12923), .ZN(n12928) );
  XOR2_X1 U15040 ( .A(n12926), .B(n12925), .Z(n13103) );
  NOR2_X1 U15041 ( .A1(n13103), .A2(n13081), .ZN(n12927) );
  AOI211_X1 U15042 ( .C1(n7604), .C2(n13078), .A(n12928), .B(n12927), .ZN(
        n12929) );
  OAI21_X1 U15043 ( .B1(n13102), .B2(n14557), .A(n12929), .ZN(P2_U3239) );
  XNOR2_X1 U15044 ( .A(n12931), .B(n12930), .ZN(n12933) );
  AOI21_X1 U15045 ( .B1(n12933), .B2(n14548), .A(n12932), .ZN(n13107) );
  AOI211_X1 U15046 ( .C1(n13105), .C2(n12951), .A(n9339), .B(n7602), .ZN(
        n13104) );
  AOI22_X1 U15047 ( .A1(n14557), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n12934), 
        .B2(n14553), .ZN(n12935) );
  OAI21_X1 U15048 ( .B1(n12936), .B2(n13076), .A(n12935), .ZN(n12942) );
  OAI21_X1 U15049 ( .B1(n12939), .B2(n12938), .A(n12937), .ZN(n12940) );
  INV_X1 U15050 ( .A(n12940), .ZN(n13108) );
  NOR2_X1 U15051 ( .A1(n13108), .A2(n13081), .ZN(n12941) );
  AOI211_X1 U15052 ( .C1(n13104), .C2(n13078), .A(n12942), .B(n12941), .ZN(
        n12943) );
  OAI21_X1 U15053 ( .B1(n13107), .B2(n14557), .A(n12943), .ZN(P2_U3240) );
  XNOR2_X1 U15054 ( .A(n12944), .B(n12950), .ZN(n12947) );
  OAI21_X1 U15055 ( .B1(n12947), .B2(n12946), .A(n12945), .ZN(n13111) );
  INV_X1 U15056 ( .A(n13111), .ZN(n12959) );
  AOI21_X1 U15057 ( .B1(n12950), .B2(n12949), .A(n12948), .ZN(n13113) );
  OAI211_X1 U15058 ( .C1(n13110), .C2(n12968), .A(n12952), .B(n12951), .ZN(
        n13109) );
  NOR2_X1 U15059 ( .A1(n13109), .A2(n12953), .ZN(n12957) );
  AOI22_X1 U15060 ( .A1(n14557), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n12954), 
        .B2(n14553), .ZN(n12955) );
  OAI21_X1 U15061 ( .B1(n13110), .B2(n13076), .A(n12955), .ZN(n12956) );
  AOI211_X1 U15062 ( .C1(n13113), .C2(n10296), .A(n12957), .B(n12956), .ZN(
        n12958) );
  OAI21_X1 U15063 ( .B1(n12959), .B2(n14557), .A(n12958), .ZN(P2_U3241) );
  XNOR2_X1 U15064 ( .A(n12960), .B(n12961), .ZN(n13119) );
  XNOR2_X1 U15065 ( .A(n12962), .B(n12961), .ZN(n12965) );
  INV_X1 U15066 ( .A(n12963), .ZN(n12964) );
  AOI21_X1 U15067 ( .B1(n12965), .B2(n14548), .A(n12964), .ZN(n13118) );
  OAI21_X1 U15068 ( .B1(n12966), .B2(n13071), .A(n13118), .ZN(n12967) );
  NAND2_X1 U15069 ( .A1(n12967), .A2(n14554), .ZN(n12973) );
  AOI211_X1 U15070 ( .C1(n13116), .C2(n12978), .A(n9339), .B(n12968), .ZN(
        n13115) );
  INV_X1 U15071 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n12969) );
  OAI22_X1 U15072 ( .A1(n12970), .A2(n13076), .B1(n12969), .B2(n14554), .ZN(
        n12971) );
  AOI21_X1 U15073 ( .B1(n13115), .B2(n13078), .A(n12971), .ZN(n12972) );
  OAI211_X1 U15074 ( .C1(n13119), .C2(n13081), .A(n12973), .B(n12972), .ZN(
        P2_U3242) );
  XOR2_X1 U15075 ( .A(n12974), .B(n12982), .Z(n12977) );
  INV_X1 U15076 ( .A(n12975), .ZN(n12976) );
  AOI21_X1 U15077 ( .B1(n12977), .B2(n14548), .A(n12976), .ZN(n13123) );
  AOI211_X1 U15078 ( .C1(n13121), .C2(n12993), .A(n9339), .B(n6751), .ZN(
        n13120) );
  AOI22_X1 U15079 ( .A1(n14557), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n12979), 
        .B2(n14553), .ZN(n12980) );
  OAI21_X1 U15080 ( .B1(n12981), .B2(n13076), .A(n12980), .ZN(n12987) );
  AND2_X1 U15081 ( .A1(n12983), .A2(n12982), .ZN(n12985) );
  OR2_X1 U15082 ( .A1(n12985), .A2(n12984), .ZN(n13124) );
  NOR2_X1 U15083 ( .A1(n13124), .A2(n13081), .ZN(n12986) );
  AOI211_X1 U15084 ( .C1(n13120), .C2(n13078), .A(n12987), .B(n12986), .ZN(
        n12988) );
  OAI21_X1 U15085 ( .B1(n13123), .B2(n14557), .A(n12988), .ZN(P2_U3243) );
  XNOR2_X1 U15086 ( .A(n12989), .B(n12999), .ZN(n12992) );
  INV_X1 U15087 ( .A(n12990), .ZN(n12991) );
  AOI21_X1 U15088 ( .B1(n12992), .B2(n14548), .A(n12991), .ZN(n13128) );
  INV_X1 U15089 ( .A(n13007), .ZN(n12995) );
  INV_X1 U15090 ( .A(n12993), .ZN(n12994) );
  AOI211_X1 U15091 ( .C1(n13126), .C2(n12995), .A(n9339), .B(n12994), .ZN(
        n13125) );
  AOI22_X1 U15092 ( .A1(P2_REG2_REG_21__SCAN_IN), .A2(n14557), .B1(n12996), 
        .B2(n14553), .ZN(n12997) );
  OAI21_X1 U15093 ( .B1(n12998), .B2(n13076), .A(n12997), .ZN(n13002) );
  XNOR2_X1 U15094 ( .A(n13000), .B(n12999), .ZN(n13129) );
  NOR2_X1 U15095 ( .A1(n13129), .A2(n13081), .ZN(n13001) );
  AOI211_X1 U15096 ( .C1(n13125), .C2(n13078), .A(n13002), .B(n13001), .ZN(
        n13003) );
  OAI21_X1 U15097 ( .B1(n13128), .B2(n14557), .A(n13003), .ZN(P2_U3244) );
  XNOR2_X1 U15098 ( .A(n13004), .B(n13012), .ZN(n13006) );
  AOI21_X1 U15099 ( .B1(n13006), .B2(n14548), .A(n13005), .ZN(n13133) );
  AOI211_X1 U15100 ( .C1(n13131), .C2(n13021), .A(n9339), .B(n13007), .ZN(
        n13130) );
  INV_X1 U15101 ( .A(n13131), .ZN(n13011) );
  INV_X1 U15102 ( .A(n13008), .ZN(n13009) );
  AOI22_X1 U15103 ( .A1(n14557), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n13009), 
        .B2(n14553), .ZN(n13010) );
  OAI21_X1 U15104 ( .B1(n13011), .B2(n13076), .A(n13010), .ZN(n13015) );
  XNOR2_X1 U15105 ( .A(n13013), .B(n13012), .ZN(n13134) );
  NOR2_X1 U15106 ( .A1(n13134), .A2(n13081), .ZN(n13014) );
  AOI211_X1 U15107 ( .C1(n13130), .C2(n13078), .A(n13015), .B(n13014), .ZN(
        n13016) );
  OAI21_X1 U15108 ( .B1(n13133), .B2(n14557), .A(n13016), .ZN(P2_U3245) );
  XNOR2_X1 U15109 ( .A(n13018), .B(n13017), .ZN(n13020) );
  AOI21_X1 U15110 ( .B1(n13020), .B2(n14548), .A(n13019), .ZN(n13138) );
  INV_X1 U15111 ( .A(n13021), .ZN(n13022) );
  AOI211_X1 U15112 ( .C1(n13136), .C2(n13036), .A(n9339), .B(n13022), .ZN(
        n13135) );
  INV_X1 U15113 ( .A(n13023), .ZN(n13024) );
  AOI22_X1 U15114 ( .A1(n14557), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13024), 
        .B2(n14553), .ZN(n13025) );
  OAI21_X1 U15115 ( .B1(n7072), .B2(n13076), .A(n13025), .ZN(n13029) );
  XNOR2_X1 U15116 ( .A(n13027), .B(n13026), .ZN(n13139) );
  NOR2_X1 U15117 ( .A1(n13139), .A2(n13081), .ZN(n13028) );
  AOI211_X1 U15118 ( .C1(n13135), .C2(n13078), .A(n13029), .B(n13028), .ZN(
        n13030) );
  OAI21_X1 U15119 ( .B1(n13138), .B2(n14557), .A(n13030), .ZN(P2_U3246) );
  XNOR2_X1 U15120 ( .A(n13032), .B(n13031), .ZN(n13035) );
  INV_X1 U15121 ( .A(n13033), .ZN(n13034) );
  AOI21_X1 U15122 ( .B1(n13035), .B2(n14548), .A(n13034), .ZN(n13143) );
  AOI211_X1 U15123 ( .C1(n13141), .C2(n13051), .A(n9339), .B(n7073), .ZN(
        n13140) );
  INV_X1 U15124 ( .A(n13037), .ZN(n13038) );
  AOI22_X1 U15125 ( .A1(n14557), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13038), 
        .B2(n14553), .ZN(n13039) );
  OAI21_X1 U15126 ( .B1(n13040), .B2(n13076), .A(n13039), .ZN(n13046) );
  OAI21_X1 U15127 ( .B1(n13043), .B2(n13042), .A(n13041), .ZN(n13044) );
  INV_X1 U15128 ( .A(n13044), .ZN(n13144) );
  NOR2_X1 U15129 ( .A1(n13144), .A2(n13081), .ZN(n13045) );
  AOI211_X1 U15130 ( .C1(n13140), .C2(n13078), .A(n13046), .B(n13045), .ZN(
        n13047) );
  OAI21_X1 U15131 ( .B1(n13143), .B2(n14557), .A(n13047), .ZN(P2_U3247) );
  XNOR2_X1 U15132 ( .A(n13048), .B(n13058), .ZN(n13050) );
  AOI21_X1 U15133 ( .B1(n13050), .B2(n14548), .A(n13049), .ZN(n13148) );
  INV_X1 U15134 ( .A(n13074), .ZN(n13053) );
  INV_X1 U15135 ( .A(n13051), .ZN(n13052) );
  AOI211_X1 U15136 ( .C1(n13146), .C2(n13053), .A(n9339), .B(n13052), .ZN(
        n13145) );
  INV_X1 U15137 ( .A(n13054), .ZN(n13055) );
  AOI22_X1 U15138 ( .A1(n14557), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13055), 
        .B2(n14553), .ZN(n13056) );
  OAI21_X1 U15139 ( .B1(n13057), .B2(n13076), .A(n13056), .ZN(n13061) );
  XNOR2_X1 U15140 ( .A(n13059), .B(n13058), .ZN(n13149) );
  NOR2_X1 U15141 ( .A1(n13149), .A2(n13081), .ZN(n13060) );
  AOI211_X1 U15142 ( .C1(n13145), .C2(n13078), .A(n13061), .B(n13060), .ZN(
        n13062) );
  OAI21_X1 U15143 ( .B1(n13148), .B2(n14557), .A(n13062), .ZN(P2_U3248) );
  NAND2_X1 U15144 ( .A1(n13063), .A2(n13066), .ZN(n13064) );
  NAND2_X1 U15145 ( .A1(n13065), .A2(n13064), .ZN(n13154) );
  XNOR2_X1 U15146 ( .A(n13066), .B(n13067), .ZN(n13070) );
  INV_X1 U15147 ( .A(n13068), .ZN(n13069) );
  AOI21_X1 U15148 ( .B1(n13070), .B2(n14548), .A(n13069), .ZN(n13153) );
  OAI21_X1 U15149 ( .B1(n13072), .B2(n13071), .A(n13153), .ZN(n13073) );
  NAND2_X1 U15150 ( .A1(n13073), .A2(n14554), .ZN(n13080) );
  AOI211_X1 U15151 ( .C1(n13151), .C2(n13075), .A(n9339), .B(n13074), .ZN(
        n13150) );
  INV_X1 U15152 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n14956) );
  OAI22_X1 U15153 ( .A1(n7458), .A2(n13076), .B1(n14554), .B2(n14956), .ZN(
        n13077) );
  AOI21_X1 U15154 ( .B1(n13150), .B2(n13078), .A(n13077), .ZN(n13079) );
  OAI211_X1 U15155 ( .C1(n13154), .C2(n13081), .A(n13080), .B(n13079), .ZN(
        P2_U3249) );
  OAI211_X1 U15156 ( .C1(n13083), .C2(n14627), .A(n13082), .B(n13084), .ZN(
        n13176) );
  MUX2_X1 U15157 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13176), .S(n14663), .Z(
        P2_U3530) );
  OAI211_X1 U15158 ( .C1(n13086), .C2(n14627), .A(n13085), .B(n13084), .ZN(
        n13177) );
  MUX2_X1 U15159 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13177), .S(n14663), .Z(
        P2_U3529) );
  AOI21_X1 U15160 ( .B1(n14637), .B2(n13088), .A(n13087), .ZN(n13089) );
  MUX2_X1 U15161 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13178), .S(n14663), .Z(
        P2_U3528) );
  OAI211_X1 U15162 ( .C1(n14583), .C2(n13095), .A(n13094), .B(n13093), .ZN(
        n13179) );
  MUX2_X1 U15163 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13179), .S(n14663), .Z(
        P2_U3527) );
  AOI21_X1 U15164 ( .B1(n14637), .B2(n13096), .A(n7590), .ZN(n13097) );
  OAI211_X1 U15165 ( .C1(n14583), .C2(n13099), .A(n13098), .B(n13097), .ZN(
        n13180) );
  MUX2_X1 U15166 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13180), .S(n14663), .Z(
        P2_U3526) );
  AOI21_X1 U15167 ( .B1(n14637), .B2(n13100), .A(n7604), .ZN(n13101) );
  OAI211_X1 U15168 ( .C1(n14583), .C2(n13103), .A(n13102), .B(n13101), .ZN(
        n13181) );
  MUX2_X1 U15169 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13181), .S(n14663), .Z(
        P2_U3525) );
  AOI21_X1 U15170 ( .B1(n14637), .B2(n13105), .A(n13104), .ZN(n13106) );
  OAI211_X1 U15171 ( .C1(n14583), .C2(n13108), .A(n13107), .B(n13106), .ZN(
        n13182) );
  MUX2_X1 U15172 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13182), .S(n14663), .Z(
        P2_U3524) );
  OAI21_X1 U15173 ( .B1(n13110), .B2(n14627), .A(n13109), .ZN(n13112) );
  AOI211_X1 U15174 ( .C1(n13113), .C2(n14614), .A(n13112), .B(n13111), .ZN(
        n13114) );
  INV_X1 U15175 ( .A(n13114), .ZN(n13183) );
  MUX2_X1 U15176 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13183), .S(n14663), .Z(
        P2_U3523) );
  AOI21_X1 U15177 ( .B1(n14637), .B2(n13116), .A(n13115), .ZN(n13117) );
  OAI211_X1 U15178 ( .C1(n14583), .C2(n13119), .A(n13118), .B(n13117), .ZN(
        n13184) );
  MUX2_X1 U15179 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13184), .S(n14663), .Z(
        P2_U3522) );
  AOI21_X1 U15180 ( .B1(n14637), .B2(n13121), .A(n13120), .ZN(n13122) );
  OAI211_X1 U15181 ( .C1(n14583), .C2(n13124), .A(n13123), .B(n13122), .ZN(
        n13185) );
  MUX2_X1 U15182 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13185), .S(n14663), .Z(
        P2_U3521) );
  AOI21_X1 U15183 ( .B1(n14637), .B2(n13126), .A(n13125), .ZN(n13127) );
  OAI211_X1 U15184 ( .C1(n14583), .C2(n13129), .A(n13128), .B(n13127), .ZN(
        n13186) );
  MUX2_X1 U15185 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13186), .S(n14663), .Z(
        P2_U3520) );
  AOI21_X1 U15186 ( .B1(n14637), .B2(n13131), .A(n13130), .ZN(n13132) );
  OAI211_X1 U15187 ( .C1(n14583), .C2(n13134), .A(n13133), .B(n13132), .ZN(
        n13187) );
  MUX2_X1 U15188 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13187), .S(n14663), .Z(
        P2_U3519) );
  AOI21_X1 U15189 ( .B1(n14637), .B2(n13136), .A(n13135), .ZN(n13137) );
  OAI211_X1 U15190 ( .C1(n14583), .C2(n13139), .A(n13138), .B(n13137), .ZN(
        n13188) );
  MUX2_X1 U15191 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13188), .S(n14663), .Z(
        P2_U3518) );
  AOI21_X1 U15192 ( .B1(n14637), .B2(n13141), .A(n13140), .ZN(n13142) );
  OAI211_X1 U15193 ( .C1(n14583), .C2(n13144), .A(n13143), .B(n13142), .ZN(
        n13189) );
  MUX2_X1 U15194 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13189), .S(n14663), .Z(
        P2_U3517) );
  AOI21_X1 U15195 ( .B1(n14637), .B2(n13146), .A(n13145), .ZN(n13147) );
  OAI211_X1 U15196 ( .C1(n14583), .C2(n13149), .A(n13148), .B(n13147), .ZN(
        n13190) );
  MUX2_X1 U15197 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13190), .S(n14663), .Z(
        P2_U3516) );
  AOI21_X1 U15198 ( .B1(n14637), .B2(n13151), .A(n13150), .ZN(n13152) );
  OAI211_X1 U15199 ( .C1(n14583), .C2(n13154), .A(n13153), .B(n13152), .ZN(
        n13191) );
  MUX2_X1 U15200 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13191), .S(n14663), .Z(
        P2_U3515) );
  AOI21_X1 U15201 ( .B1(n14637), .B2(n13156), .A(n13155), .ZN(n13157) );
  OAI211_X1 U15202 ( .C1(n14583), .C2(n13159), .A(n13158), .B(n13157), .ZN(
        n13192) );
  MUX2_X1 U15203 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n13192), .S(n14663), .Z(
        P2_U3514) );
  OAI21_X1 U15204 ( .B1(n13161), .B2(n14627), .A(n13160), .ZN(n13163) );
  AOI211_X1 U15205 ( .C1(n13164), .C2(n14614), .A(n13163), .B(n13162), .ZN(
        n13194) );
  NAND2_X1 U15206 ( .A1(n14661), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n13165) );
  OAI21_X1 U15207 ( .B1(n13194), .B2(n14661), .A(n13165), .ZN(P2_U3513) );
  AOI21_X1 U15208 ( .B1(n14637), .B2(n13167), .A(n13166), .ZN(n13168) );
  OAI211_X1 U15209 ( .C1(n14583), .C2(n13170), .A(n13169), .B(n13168), .ZN(
        n13195) );
  MUX2_X1 U15210 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n13195), .S(n14663), .Z(
        P2_U3512) );
  AOI21_X1 U15211 ( .B1(n14637), .B2(n13172), .A(n13171), .ZN(n13173) );
  OAI211_X1 U15212 ( .C1(n14583), .C2(n13175), .A(n13174), .B(n13173), .ZN(
        n13196) );
  MUX2_X1 U15213 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n13196), .S(n14663), .Z(
        P2_U3511) );
  MUX2_X1 U15214 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13176), .S(n14648), .Z(
        P2_U3498) );
  MUX2_X1 U15215 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13177), .S(n14648), .Z(
        P2_U3497) );
  MUX2_X1 U15216 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13178), .S(n14648), .Z(
        P2_U3496) );
  MUX2_X1 U15217 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13179), .S(n14648), .Z(
        P2_U3495) );
  MUX2_X1 U15218 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13180), .S(n14648), .Z(
        P2_U3494) );
  MUX2_X1 U15219 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13181), .S(n14648), .Z(
        P2_U3493) );
  MUX2_X1 U15220 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13182), .S(n14648), .Z(
        P2_U3492) );
  MUX2_X1 U15221 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13183), .S(n14648), .Z(
        P2_U3491) );
  MUX2_X1 U15222 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13184), .S(n14648), .Z(
        P2_U3490) );
  MUX2_X1 U15223 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13185), .S(n14648), .Z(
        P2_U3489) );
  MUX2_X1 U15224 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13186), .S(n14648), .Z(
        P2_U3488) );
  MUX2_X1 U15225 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13187), .S(n14648), .Z(
        P2_U3487) );
  MUX2_X1 U15226 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13188), .S(n14648), .Z(
        P2_U3486) );
  MUX2_X1 U15227 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13189), .S(n14648), .Z(
        P2_U3484) );
  MUX2_X1 U15228 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13190), .S(n14648), .Z(
        P2_U3481) );
  MUX2_X1 U15229 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13191), .S(n14648), .Z(
        P2_U3478) );
  MUX2_X1 U15230 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n13192), .S(n14648), .Z(
        P2_U3475) );
  NAND2_X1 U15231 ( .A1(n14646), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n13193) );
  OAI21_X1 U15232 ( .B1(n13194), .B2(n14646), .A(n13193), .ZN(P2_U3472) );
  MUX2_X1 U15233 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n13195), .S(n14648), .Z(
        P2_U3469) );
  MUX2_X1 U15234 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n13196), .S(n14648), .Z(
        P2_U3466) );
  INV_X1 U15235 ( .A(n11567), .ZN(n13821) );
  NOR4_X1 U15236 ( .A1(n7216), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13197), .A4(
        P2_U3088), .ZN(n13198) );
  AOI21_X1 U15237 ( .B1(P1_DATAO_REG_31__SCAN_IN), .B2(n6626), .A(n13198), 
        .ZN(n13199) );
  OAI21_X1 U15238 ( .B1(n13821), .B2(n13213), .A(n13199), .ZN(P2_U3296) );
  INV_X1 U15239 ( .A(n13200), .ZN(n13827) );
  OAI222_X1 U15240 ( .A1(P2_U3088), .A2(n13201), .B1(n13213), .B2(n13827), 
        .C1(n14963), .C2(n13210), .ZN(P2_U3298) );
  INV_X1 U15241 ( .A(n11551), .ZN(n13829) );
  AOI21_X1 U15242 ( .B1(n6626), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13202), 
        .ZN(n13203) );
  OAI21_X1 U15243 ( .B1(n13829), .B2(n13213), .A(n13203), .ZN(P2_U3299) );
  INV_X1 U15244 ( .A(n13204), .ZN(n13832) );
  OAI222_X1 U15245 ( .A1(P2_U3088), .A2(n13206), .B1(n13213), .B2(n13832), 
        .C1(n13205), .C2(n13210), .ZN(P2_U3300) );
  INV_X1 U15246 ( .A(n13207), .ZN(n13209) );
  INV_X1 U15247 ( .A(n13208), .ZN(n13836) );
  OAI222_X1 U15248 ( .A1(P2_U3088), .A2(n13209), .B1(n13213), .B2(n13836), 
        .C1(n6922), .C2(n13210), .ZN(P2_U3301) );
  OAI222_X1 U15249 ( .A1(n13214), .A2(P2_U3088), .B1(n13213), .B2(n13212), 
        .C1(n13211), .C2(n13210), .ZN(P2_U3302) );
  INV_X1 U15250 ( .A(n13215), .ZN(n13216) );
  MUX2_X1 U15251 ( .A(n13216), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  AOI22_X1 U15252 ( .A1(n14087), .A2(n13608), .B1(n13547), .B2(n6454), .ZN(
        n13571) );
  OAI22_X1 U15253 ( .A1(n13334), .A2(n13571), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13220), .ZN(n13221) );
  AOI21_X1 U15254 ( .B1(n13326), .B2(n13579), .A(n13221), .ZN(n13222) );
  INV_X1 U15255 ( .A(n13223), .ZN(n13224) );
  AOI21_X1 U15256 ( .B1(n13226), .B2(n13225), .A(n13224), .ZN(n13233) );
  NAND2_X1 U15257 ( .A1(n14073), .A2(n13342), .ZN(n13227) );
  NAND2_X1 U15258 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14218)
         );
  OAI211_X1 U15259 ( .C1(n13228), .C2(n13313), .A(n13227), .B(n14218), .ZN(
        n13229) );
  AOI21_X1 U15260 ( .B1(n13230), .B2(n13326), .A(n13229), .ZN(n13232) );
  NAND2_X1 U15261 ( .A1(n14136), .A2(n14075), .ZN(n13231) );
  OAI211_X1 U15262 ( .C1(n13233), .C2(n14078), .A(n13232), .B(n13231), .ZN(
        P1_U3215) );
  INV_X1 U15263 ( .A(n13778), .ZN(n13646) );
  NOR3_X1 U15264 ( .A1(n6491), .A2(n6720), .A3(n13235), .ZN(n13238) );
  INV_X1 U15265 ( .A(n13236), .ZN(n13237) );
  OAI21_X1 U15266 ( .B1(n13238), .B2(n13237), .A(n13320), .ZN(n13242) );
  AOI22_X1 U15267 ( .A1(n13513), .A2(n14087), .B1(n6454), .B2(n6879), .ZN(
        n13642) );
  OAI22_X1 U15268 ( .A1(n13642), .A2(n13334), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13239), .ZN(n13240) );
  AOI21_X1 U15269 ( .B1(n13643), .B2(n13326), .A(n13240), .ZN(n13241) );
  OAI211_X1 U15270 ( .C1(n13646), .C2(n13329), .A(n13242), .B(n13241), .ZN(
        P1_U3216) );
  INV_X1 U15271 ( .A(n13700), .ZN(n14104) );
  INV_X1 U15272 ( .A(n13243), .ZN(n13246) );
  OAI21_X1 U15273 ( .B1(n13246), .B2(n13245), .A(n13244), .ZN(n13248) );
  NAND3_X1 U15274 ( .A1(n13248), .A2(n13320), .A3(n13247), .ZN(n13252) );
  INV_X1 U15275 ( .A(n13695), .ZN(n13250) );
  AOI22_X1 U15276 ( .A1(n13256), .A2(n6454), .B1(n14087), .B2(n13507), .ZN(
        n14102) );
  NAND2_X1 U15277 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13489)
         );
  OAI21_X1 U15278 ( .B1(n14102), .B2(n13334), .A(n13489), .ZN(n13249) );
  AOI21_X1 U15279 ( .B1(n13250), .B2(n13326), .A(n13249), .ZN(n13251) );
  OAI211_X1 U15280 ( .C1(n14104), .C2(n13329), .A(n13252), .B(n13251), .ZN(
        P1_U3219) );
  INV_X1 U15281 ( .A(n13253), .ZN(n13302) );
  AOI21_X1 U15282 ( .B1(n13255), .B2(n13254), .A(n13302), .ZN(n13261) );
  NOR2_X1 U15283 ( .A1(n14083), .A2(n13669), .ZN(n13259) );
  AOI22_X1 U15284 ( .A1(n13513), .A2(n6454), .B1(n14087), .B2(n13256), .ZN(
        n13791) );
  OAI22_X1 U15285 ( .A1(n13791), .A2(n13334), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13257), .ZN(n13258) );
  AOI211_X1 U15286 ( .C1(n13529), .C2(n14075), .A(n13259), .B(n13258), .ZN(
        n13260) );
  OAI21_X1 U15287 ( .B1(n13261), .B2(n14078), .A(n13260), .ZN(P1_U3223) );
  OAI21_X1 U15288 ( .B1(n13264), .B2(n13263), .A(n13262), .ZN(n13265) );
  NAND2_X1 U15289 ( .A1(n13265), .A2(n13320), .ZN(n13271) );
  OAI22_X1 U15290 ( .A1(n13313), .A2(n15021), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13266), .ZN(n13269) );
  NOR2_X1 U15291 ( .A1(n13267), .A2(n13607), .ZN(n13268) );
  AOI211_X1 U15292 ( .C1(n13611), .C2(n13326), .A(n13269), .B(n13268), .ZN(
        n13270) );
  OAI211_X1 U15293 ( .C1(n13534), .C2(n13329), .A(n13271), .B(n13270), .ZN(
        P1_U3225) );
  INV_X1 U15294 ( .A(n13272), .ZN(n14071) );
  INV_X1 U15295 ( .A(n13273), .ZN(n13275) );
  NOR3_X1 U15296 ( .A1(n14071), .A2(n13275), .A3(n13274), .ZN(n13278) );
  INV_X1 U15297 ( .A(n13276), .ZN(n13277) );
  OAI21_X1 U15298 ( .B1(n13278), .B2(n13277), .A(n13320), .ZN(n13283) );
  NAND2_X1 U15299 ( .A1(n14073), .A2(n13340), .ZN(n13279) );
  NAND2_X1 U15300 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14267)
         );
  OAI211_X1 U15301 ( .C1(n13525), .C2(n13313), .A(n13279), .B(n14267), .ZN(
        n13280) );
  AOI21_X1 U15302 ( .B1(n13281), .B2(n13326), .A(n13280), .ZN(n13282) );
  OAI211_X1 U15303 ( .C1(n13522), .C2(n13329), .A(n13283), .B(n13282), .ZN(
        P1_U3228) );
  OAI21_X1 U15304 ( .B1(n13286), .B2(n13285), .A(n13284), .ZN(n13287) );
  NAND2_X1 U15305 ( .A1(n13287), .A2(n13320), .ZN(n13291) );
  AOI22_X1 U15306 ( .A1(n14087), .A2(n13516), .B1(n13533), .B2(n6454), .ZN(
        n13625) );
  OAI22_X1 U15307 ( .A1(n13334), .A2(n13625), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13288), .ZN(n13289) );
  AOI21_X1 U15308 ( .B1(n13326), .B2(n13630), .A(n13289), .ZN(n13290) );
  OAI211_X1 U15309 ( .C1(n13772), .C2(n13329), .A(n13291), .B(n13290), .ZN(
        P1_U3229) );
  XNOR2_X1 U15310 ( .A(n13293), .B(n13292), .ZN(n13299) );
  AOI22_X1 U15311 ( .A1(n14074), .A2(n13678), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13295) );
  NAND2_X1 U15312 ( .A1(n14073), .A2(n13709), .ZN(n13294) );
  OAI211_X1 U15313 ( .C1(n14083), .C2(n13296), .A(n13295), .B(n13294), .ZN(
        n13297) );
  AOI21_X1 U15314 ( .B1(n7031), .B2(n14075), .A(n13297), .ZN(n13298) );
  OAI21_X1 U15315 ( .B1(n13299), .B2(n14078), .A(n13298), .ZN(P1_U3233) );
  NOR3_X1 U15316 ( .A1(n13302), .A2(n6721), .A3(n13301), .ZN(n13303) );
  OAI21_X1 U15317 ( .B1(n13303), .B2(n6491), .A(n13320), .ZN(n13308) );
  AND2_X1 U15318 ( .A1(n13516), .A2(n6454), .ZN(n13304) );
  AOI21_X1 U15319 ( .B1(n13678), .B2(n14087), .A(n13304), .ZN(n13784) );
  INV_X1 U15320 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13305) );
  OAI22_X1 U15321 ( .A1(n13784), .A2(n13334), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13305), .ZN(n13306) );
  AOI21_X1 U15322 ( .B1(n13657), .B2(n13326), .A(n13306), .ZN(n13307) );
  OAI211_X1 U15323 ( .C1(n13329), .C2(n13786), .A(n13308), .B(n13307), .ZN(
        P1_U3235) );
  INV_X1 U15324 ( .A(n13717), .ZN(n14111) );
  OAI21_X1 U15325 ( .B1(n13310), .B2(n13309), .A(n13243), .ZN(n13311) );
  NAND2_X1 U15326 ( .A1(n13311), .A2(n13320), .ZN(n13316) );
  INV_X1 U15327 ( .A(n13709), .ZN(n13527) );
  NAND2_X1 U15328 ( .A1(n14073), .A2(n14086), .ZN(n13312) );
  NAND2_X1 U15329 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14286)
         );
  OAI211_X1 U15330 ( .C1(n13527), .C2(n13313), .A(n13312), .B(n14286), .ZN(
        n13314) );
  AOI21_X1 U15331 ( .B1(n13716), .B2(n13326), .A(n13314), .ZN(n13315) );
  OAI211_X1 U15332 ( .C1(n14111), .C2(n13329), .A(n13316), .B(n13315), .ZN(
        P1_U3238) );
  OAI21_X1 U15333 ( .B1(n13319), .B2(n13318), .A(n13317), .ZN(n13321) );
  NAND2_X1 U15334 ( .A1(n13321), .A2(n13320), .ZN(n13328) );
  NAND2_X1 U15335 ( .A1(n13556), .A2(n6454), .ZN(n13323) );
  NAND2_X1 U15336 ( .A1(n13533), .A2(n14087), .ZN(n13322) );
  AND2_X1 U15337 ( .A1(n13323), .A2(n13322), .ZN(n13754) );
  OAI22_X1 U15338 ( .A1(n13334), .A2(n13754), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13324), .ZN(n13325) );
  AOI21_X1 U15339 ( .B1(n13326), .B2(n13594), .A(n13325), .ZN(n13327) );
  OAI211_X1 U15340 ( .C1(n13756), .C2(n13329), .A(n13328), .B(n13327), .ZN(
        P1_U3240) );
  XNOR2_X1 U15341 ( .A(n13331), .B(n13330), .ZN(n13339) );
  NOR2_X1 U15342 ( .A1(n14083), .A2(n13332), .ZN(n13336) );
  NAND2_X1 U15343 ( .A1(P1_REG3_REG_15__SCAN_IN), .A2(P1_U3086), .ZN(n14233)
         );
  OAI21_X1 U15344 ( .B1(n13334), .B2(n13333), .A(n14233), .ZN(n13335) );
  AOI211_X1 U15345 ( .C1(n13337), .C2(n14075), .A(n13336), .B(n13335), .ZN(
        n13338) );
  OAI21_X1 U15346 ( .B1(n13339), .B2(n14078), .A(n13338), .ZN(P1_U3241) );
  MUX2_X1 U15347 ( .A(n13494), .B(P1_DATAO_REG_31__SCAN_IN), .S(n15020), .Z(
        P1_U3591) );
  MUX2_X1 U15348 ( .A(n13543), .B(P1_DATAO_REG_30__SCAN_IN), .S(n15020), .Z(
        P1_U3590) );
  MUX2_X1 U15349 ( .A(n13557), .B(P1_DATAO_REG_29__SCAN_IN), .S(n15020), .Z(
        P1_U3589) );
  MUX2_X1 U15350 ( .A(n13547), .B(P1_DATAO_REG_28__SCAN_IN), .S(n15020), .Z(
        P1_U3588) );
  MUX2_X1 U15351 ( .A(n13556), .B(P1_DATAO_REG_27__SCAN_IN), .S(n15020), .Z(
        P1_U3587) );
  MUX2_X1 U15352 ( .A(n13533), .B(P1_DATAO_REG_25__SCAN_IN), .S(n15020), .Z(
        P1_U3585) );
  MUX2_X1 U15353 ( .A(n6879), .B(P1_DATAO_REG_24__SCAN_IN), .S(n15020), .Z(
        P1_U3584) );
  MUX2_X1 U15354 ( .A(n13516), .B(P1_DATAO_REG_23__SCAN_IN), .S(n15020), .Z(
        P1_U3583) );
  MUX2_X1 U15355 ( .A(n13513), .B(P1_DATAO_REG_22__SCAN_IN), .S(n15020), .Z(
        P1_U3582) );
  MUX2_X1 U15356 ( .A(n13678), .B(P1_DATAO_REG_21__SCAN_IN), .S(n15020), .Z(
        P1_U3581) );
  MUX2_X1 U15357 ( .A(n13709), .B(P1_DATAO_REG_19__SCAN_IN), .S(n15020), .Z(
        P1_U3579) );
  MUX2_X1 U15358 ( .A(n13507), .B(P1_DATAO_REG_18__SCAN_IN), .S(n15020), .Z(
        P1_U3578) );
  MUX2_X1 U15359 ( .A(n14086), .B(P1_DATAO_REG_17__SCAN_IN), .S(n15020), .Z(
        P1_U3577) );
  MUX2_X1 U15360 ( .A(n13340), .B(P1_DATAO_REG_16__SCAN_IN), .S(n15020), .Z(
        P1_U3576) );
  MUX2_X1 U15361 ( .A(n14088), .B(P1_DATAO_REG_15__SCAN_IN), .S(n15020), .Z(
        P1_U3575) );
  MUX2_X1 U15362 ( .A(n13341), .B(P1_DATAO_REG_14__SCAN_IN), .S(n15020), .Z(
        P1_U3574) );
  MUX2_X1 U15363 ( .A(n13342), .B(P1_DATAO_REG_13__SCAN_IN), .S(n15020), .Z(
        P1_U3573) );
  MUX2_X1 U15364 ( .A(n13343), .B(P1_DATAO_REG_12__SCAN_IN), .S(n15020), .Z(
        P1_U3572) );
  MUX2_X1 U15365 ( .A(n13344), .B(P1_DATAO_REG_11__SCAN_IN), .S(n15020), .Z(
        P1_U3571) );
  MUX2_X1 U15366 ( .A(n13345), .B(P1_DATAO_REG_10__SCAN_IN), .S(n15020), .Z(
        P1_U3570) );
  MUX2_X1 U15367 ( .A(n13346), .B(P1_DATAO_REG_9__SCAN_IN), .S(n15020), .Z(
        P1_U3569) );
  MUX2_X1 U15368 ( .A(n13347), .B(P1_DATAO_REG_8__SCAN_IN), .S(n15020), .Z(
        P1_U3568) );
  MUX2_X1 U15369 ( .A(n13348), .B(P1_DATAO_REG_7__SCAN_IN), .S(n15020), .Z(
        P1_U3567) );
  MUX2_X1 U15370 ( .A(n13349), .B(P1_DATAO_REG_6__SCAN_IN), .S(n15020), .Z(
        P1_U3566) );
  MUX2_X1 U15371 ( .A(n13350), .B(P1_DATAO_REG_5__SCAN_IN), .S(n15020), .Z(
        P1_U3565) );
  MUX2_X1 U15372 ( .A(n13351), .B(P1_DATAO_REG_4__SCAN_IN), .S(n15020), .Z(
        P1_U3564) );
  MUX2_X1 U15373 ( .A(n13352), .B(P1_DATAO_REG_3__SCAN_IN), .S(n15020), .Z(
        P1_U3563) );
  MUX2_X1 U15374 ( .A(n13353), .B(P1_DATAO_REG_2__SCAN_IN), .S(n15020), .Z(
        P1_U3562) );
  MUX2_X1 U15375 ( .A(n13354), .B(P1_DATAO_REG_1__SCAN_IN), .S(n15020), .Z(
        P1_U3561) );
  MUX2_X1 U15376 ( .A(n13355), .B(P1_DATAO_REG_0__SCAN_IN), .S(n15020), .Z(
        P1_U3560) );
  INV_X1 U15377 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n13357) );
  INV_X1 U15378 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n13356) );
  OAI22_X1 U15379 ( .A1(n14288), .A2(n13357), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13356), .ZN(n13358) );
  AOI21_X1 U15380 ( .B1(n13359), .B2(n14276), .A(n13358), .ZN(n13367) );
  OAI211_X1 U15381 ( .C1(n13362), .C2(n13361), .A(n14226), .B(n13360), .ZN(
        n13366) );
  OAI211_X1 U15382 ( .C1(n13364), .C2(n13368), .A(n14280), .B(n13363), .ZN(
        n13365) );
  NAND3_X1 U15383 ( .A1(n13367), .A2(n13366), .A3(n13365), .ZN(P1_U3244) );
  INV_X1 U15384 ( .A(n13368), .ZN(n13369) );
  MUX2_X1 U15385 ( .A(n13370), .B(n13369), .S(n13492), .Z(n13373) );
  AOI21_X1 U15386 ( .B1(n7373), .B2(n13371), .A(n15020), .ZN(n13372) );
  OAI21_X1 U15387 ( .B1(n13373), .B2(n13828), .A(n13372), .ZN(n13410) );
  INV_X1 U15388 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n13374) );
  OAI22_X1 U15389 ( .A1(n14288), .A2(n14986), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13374), .ZN(n13375) );
  AOI21_X1 U15390 ( .B1(n13376), .B2(n14276), .A(n13375), .ZN(n13385) );
  OAI211_X1 U15391 ( .C1(n13379), .C2(n13378), .A(n14280), .B(n13377), .ZN(
        n13384) );
  OAI211_X1 U15392 ( .C1(n13382), .C2(n13381), .A(n14226), .B(n13380), .ZN(
        n13383) );
  NAND4_X1 U15393 ( .A1(n13410), .A2(n13385), .A3(n13384), .A4(n13383), .ZN(
        P1_U3245) );
  NAND2_X1 U15394 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n13386) );
  OAI21_X1 U15395 ( .B1(n14288), .B2(n6843), .A(n13386), .ZN(n13387) );
  AOI21_X1 U15396 ( .B1(n14276), .B2(n13388), .A(n13387), .ZN(n13397) );
  OAI211_X1 U15397 ( .C1(n13391), .C2(n13390), .A(n14226), .B(n13389), .ZN(
        n13396) );
  OAI211_X1 U15398 ( .C1(n13394), .C2(n13393), .A(n14280), .B(n13392), .ZN(
        n13395) );
  NAND3_X1 U15399 ( .A1(n13397), .A2(n13396), .A3(n13395), .ZN(P1_U3246) );
  OAI21_X1 U15400 ( .B1(n14288), .B2(n6932), .A(n13398), .ZN(n13399) );
  AOI21_X1 U15401 ( .B1(n14276), .B2(n13400), .A(n13399), .ZN(n13409) );
  OAI211_X1 U15402 ( .C1(n13403), .C2(n13402), .A(n14226), .B(n13401), .ZN(
        n13408) );
  OAI211_X1 U15403 ( .C1(n13406), .C2(n13405), .A(n14280), .B(n13404), .ZN(
        n13407) );
  NAND4_X1 U15404 ( .A1(n13410), .A2(n13409), .A3(n13408), .A4(n13407), .ZN(
        P1_U3247) );
  NAND2_X1 U15405 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n13411) );
  OAI21_X1 U15406 ( .B1(n14288), .B2(n13903), .A(n13411), .ZN(n13412) );
  AOI21_X1 U15407 ( .B1(n14276), .B2(n13413), .A(n13412), .ZN(n13422) );
  OAI211_X1 U15408 ( .C1(n13416), .C2(n13415), .A(n14226), .B(n13414), .ZN(
        n13421) );
  OAI211_X1 U15409 ( .C1(n13419), .C2(n13418), .A(n14280), .B(n13417), .ZN(
        n13420) );
  NAND3_X1 U15410 ( .A1(n13422), .A2(n13421), .A3(n13420), .ZN(P1_U3249) );
  OAI21_X1 U15411 ( .B1(n14288), .B2(n14911), .A(n13423), .ZN(n13424) );
  AOI21_X1 U15412 ( .B1(n14276), .B2(n13425), .A(n13424), .ZN(n13434) );
  OAI211_X1 U15413 ( .C1(n13428), .C2(n13427), .A(n14226), .B(n13426), .ZN(
        n13433) );
  OAI211_X1 U15414 ( .C1(n13431), .C2(n13430), .A(n14280), .B(n13429), .ZN(
        n13432) );
  NAND3_X1 U15415 ( .A1(n13434), .A2(n13433), .A3(n13432), .ZN(P1_U3250) );
  OAI211_X1 U15416 ( .C1(n13437), .C2(n13436), .A(n13435), .B(n14226), .ZN(
        n13446) );
  NAND2_X1 U15417 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n13438)
         );
  OAI21_X1 U15418 ( .B1(n14288), .B2(n13877), .A(n13438), .ZN(n13439) );
  AOI21_X1 U15419 ( .B1(n14276), .B2(n13440), .A(n13439), .ZN(n13445) );
  OAI211_X1 U15420 ( .C1(n13443), .C2(n13442), .A(n14280), .B(n13441), .ZN(
        n13444) );
  NAND3_X1 U15421 ( .A1(n13446), .A2(n13445), .A3(n13444), .ZN(P1_U3253) );
  INV_X1 U15422 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14270) );
  INV_X1 U15423 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n13447) );
  OR2_X1 U15424 ( .A1(n14239), .A2(n13447), .ZN(n13449) );
  NAND2_X1 U15425 ( .A1(n14239), .A2(n13447), .ZN(n13448) );
  AND2_X1 U15426 ( .A1(n13449), .A2(n13448), .ZN(n14236) );
  INV_X1 U15427 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n13450) );
  MUX2_X1 U15428 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n13450), .S(n14211), .Z(
        n14208) );
  OR2_X1 U15429 ( .A1(n13451), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n13452) );
  NAND2_X1 U15430 ( .A1(n13453), .A2(n13452), .ZN(n14192) );
  INV_X1 U15431 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n13454) );
  MUX2_X1 U15432 ( .A(n13454), .B(P1_REG1_REG_13__SCAN_IN), .S(n14190), .Z(
        n14191) );
  NOR2_X1 U15433 ( .A1(n14192), .A2(n14191), .ZN(n14193) );
  AOI21_X1 U15434 ( .B1(n14190), .B2(P1_REG1_REG_13__SCAN_IN), .A(n14193), 
        .ZN(n14209) );
  NAND2_X1 U15435 ( .A1(n14208), .A2(n14209), .ZN(n14207) );
  OR2_X1 U15436 ( .A1(n14211), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n13455) );
  NAND2_X1 U15437 ( .A1(n14207), .A2(n13455), .ZN(n13456) );
  NAND2_X1 U15438 ( .A1(n14230), .A2(n13456), .ZN(n13457) );
  XNOR2_X1 U15439 ( .A(n13456), .B(n13473), .ZN(n14225) );
  INV_X1 U15440 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14224) );
  NAND2_X1 U15441 ( .A1(n14225), .A2(n14224), .ZN(n14223) );
  NAND2_X1 U15442 ( .A1(n13457), .A2(n14223), .ZN(n14237) );
  NOR2_X1 U15443 ( .A1(n14236), .A2(n14237), .ZN(n14238) );
  AOI21_X1 U15444 ( .B1(n14239), .B2(P1_REG1_REG_16__SCAN_IN), .A(n14238), 
        .ZN(n14253) );
  INV_X1 U15445 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n13458) );
  OR2_X1 U15446 ( .A1(n14258), .A2(n13458), .ZN(n13460) );
  NAND2_X1 U15447 ( .A1(n14258), .A2(n13458), .ZN(n13459) );
  NAND2_X1 U15448 ( .A1(n13460), .A2(n13459), .ZN(n14256) );
  INV_X1 U15449 ( .A(n14256), .ZN(n13461) );
  NOR2_X1 U15450 ( .A1(n14253), .A2(n13461), .ZN(n14254) );
  AOI21_X1 U15451 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n14258), .A(n14254), 
        .ZN(n13462) );
  XNOR2_X1 U15452 ( .A(n13479), .B(n13462), .ZN(n14271) );
  NOR2_X1 U15453 ( .A1(n14270), .A2(n14271), .ZN(n14272) );
  NOR2_X1 U15454 ( .A1(n13462), .A2(n13479), .ZN(n13463) );
  NOR2_X1 U15455 ( .A1(n14272), .A2(n13463), .ZN(n13464) );
  INV_X1 U15456 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14109) );
  XOR2_X1 U15457 ( .A(n13464), .B(n14109), .Z(n13483) );
  OR2_X1 U15458 ( .A1(n14239), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13466) );
  NAND2_X1 U15459 ( .A1(n14239), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n13465) );
  NAND2_X1 U15460 ( .A1(n13466), .A2(n13465), .ZN(n14243) );
  INV_X1 U15461 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n13467) );
  MUX2_X1 U15462 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n13467), .S(n14211), .Z(
        n14214) );
  NAND2_X1 U15463 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n14190), .ZN(n13471) );
  OR2_X1 U15464 ( .A1(n14190), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n13468) );
  NAND2_X1 U15465 ( .A1(n13468), .A2(n13471), .ZN(n14196) );
  NAND2_X1 U15466 ( .A1(n13470), .A2(n13469), .ZN(n14197) );
  OR2_X1 U15467 ( .A1(n14196), .A2(n14197), .ZN(n14198) );
  NAND2_X1 U15468 ( .A1(n13471), .A2(n14198), .ZN(n14213) );
  NAND2_X1 U15469 ( .A1(n14214), .A2(n14213), .ZN(n14212) );
  NAND2_X1 U15470 ( .A1(n14211), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n13472) );
  AND2_X1 U15471 ( .A1(n14212), .A2(n13472), .ZN(n13474) );
  NAND2_X1 U15472 ( .A1(n13474), .A2(n14230), .ZN(n13475) );
  XNOR2_X1 U15473 ( .A(n13474), .B(n13473), .ZN(n14221) );
  NAND2_X1 U15474 ( .A1(n14221), .A2(n11002), .ZN(n14220) );
  NAND2_X1 U15475 ( .A1(n13475), .A2(n14220), .ZN(n14244) );
  NOR2_X1 U15476 ( .A1(n14243), .A2(n14244), .ZN(n14245) );
  AOI21_X1 U15477 ( .B1(n14239), .B2(P1_REG2_REG_16__SCAN_IN), .A(n14245), 
        .ZN(n14260) );
  OR2_X1 U15478 ( .A1(n14258), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13477) );
  NAND2_X1 U15479 ( .A1(n14258), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n13476) );
  NAND2_X1 U15480 ( .A1(n13477), .A2(n13476), .ZN(n14261) );
  NOR2_X1 U15481 ( .A1(n14260), .A2(n14261), .ZN(n14259) );
  AOI21_X1 U15482 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n14258), .A(n14259), 
        .ZN(n13478) );
  NOR2_X1 U15483 ( .A1(n13478), .A2(n13479), .ZN(n13480) );
  XNOR2_X1 U15484 ( .A(n13479), .B(n13478), .ZN(n14278) );
  NOR2_X1 U15485 ( .A1(n8316), .A2(n14278), .ZN(n14277) );
  NOR2_X1 U15486 ( .A1(n13480), .A2(n14277), .ZN(n13481) );
  XNOR2_X1 U15487 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n13481), .ZN(n13482) );
  AOI22_X1 U15488 ( .A1(n13483), .A2(n14226), .B1(n13482), .B2(n14280), .ZN(
        n13488) );
  INV_X1 U15489 ( .A(n13482), .ZN(n13485) );
  NOR2_X1 U15490 ( .A1(n13483), .A2(n14284), .ZN(n13484) );
  AOI211_X1 U15491 ( .C1(n14280), .C2(n13485), .A(n14276), .B(n13484), .ZN(
        n13487) );
  MUX2_X1 U15492 ( .A(n13488), .B(n13487), .S(n13486), .Z(n13490) );
  OAI211_X1 U15493 ( .C1(n7275), .C2(n14288), .A(n13490), .B(n13489), .ZN(
        P1_U3262) );
  NOR2_X2 U15494 ( .A1(n13778), .A2(n13655), .ZN(n13641) );
  NAND2_X1 U15495 ( .A1(n13772), .A2(n13641), .ZN(n13629) );
  OR2_X2 U15496 ( .A1(n13491), .A2(n13606), .ZN(n13592) );
  NAND2_X1 U15497 ( .A1(n13541), .A2(n13736), .ZN(n13497) );
  XNOR2_X1 U15498 ( .A(n13733), .B(n13497), .ZN(n13731) );
  NAND2_X1 U15499 ( .A1(n13731), .A2(n13725), .ZN(n13496) );
  NAND2_X1 U15500 ( .A1(n13492), .A2(P1_B_REG_SCAN_IN), .ZN(n13493) );
  AND2_X1 U15501 ( .A1(n6454), .A2(n13493), .ZN(n13542) );
  NAND2_X1 U15502 ( .A1(n13542), .A2(n13494), .ZN(n13734) );
  NOR2_X1 U15503 ( .A1(n14315), .A2(n13734), .ZN(n13498) );
  AOI21_X1 U15504 ( .B1(n14315), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13498), 
        .ZN(n13495) );
  OAI211_X1 U15505 ( .C1(n13733), .C2(n14298), .A(n13496), .B(n13495), .ZN(
        P1_U3263) );
  OAI211_X1 U15506 ( .C1(n13541), .C2(n13736), .A(n9843), .B(n13497), .ZN(
        n13735) );
  NAND2_X1 U15507 ( .A1(n14315), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13500) );
  INV_X1 U15508 ( .A(n13498), .ZN(n13499) );
  OAI211_X1 U15509 ( .C1(n13736), .C2(n14298), .A(n13500), .B(n13499), .ZN(
        n13501) );
  INV_X1 U15510 ( .A(n13501), .ZN(n13502) );
  OAI21_X1 U15511 ( .B1(n13735), .B2(n13720), .A(n13502), .ZN(P1_U3264) );
  INV_X1 U15512 ( .A(n13533), .ZN(n13519) );
  INV_X1 U15513 ( .A(n13503), .ZN(n13504) );
  AND2_X1 U15514 ( .A1(n13717), .A2(n13507), .ZN(n13509) );
  OR2_X1 U15515 ( .A1(n13717), .A2(n13507), .ZN(n13508) );
  OR2_X1 U15516 ( .A1(n13700), .A2(n13709), .ZN(n13510) );
  NAND2_X1 U15517 ( .A1(n13511), .A2(n13510), .ZN(n13683) );
  OR2_X1 U15518 ( .A1(n13799), .A2(n13528), .ZN(n13512) );
  INV_X1 U15519 ( .A(n13531), .ZN(n13654) );
  OR2_X1 U15520 ( .A1(n13661), .A2(n13513), .ZN(n13514) );
  NAND2_X1 U15521 ( .A1(n13515), .A2(n13514), .ZN(n13649) );
  INV_X1 U15522 ( .A(n13638), .ZN(n13648) );
  NAND2_X1 U15523 ( .A1(n13778), .A2(n13516), .ZN(n13517) );
  NAND2_X1 U15524 ( .A1(n13772), .A2(n13607), .ZN(n13518) );
  NAND2_X1 U15525 ( .A1(n13522), .A2(n14086), .ZN(n13523) );
  INV_X1 U15526 ( .A(n13529), .ZN(n13793) );
  INV_X1 U15527 ( .A(n13587), .ZN(n13590) );
  NAND2_X1 U15528 ( .A1(n13554), .A2(n13537), .ZN(n13540) );
  NAND2_X1 U15529 ( .A1(n13741), .A2(n14313), .ZN(n13551) );
  NAND2_X1 U15530 ( .A1(n13543), .A2(n13542), .ZN(n13738) );
  INV_X1 U15531 ( .A(n13544), .ZN(n13545) );
  OAI22_X1 U15532 ( .A1(n13546), .A2(n13738), .B1(n13545), .B2(n14093), .ZN(
        n13549) );
  NAND2_X1 U15533 ( .A1(n13547), .A2(n14087), .ZN(n13737) );
  NOR2_X1 U15534 ( .A1(n14315), .A2(n13737), .ZN(n13548) );
  AOI211_X1 U15535 ( .C1(n14322), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13549), 
        .B(n13548), .ZN(n13550) );
  OAI211_X1 U15536 ( .C1(n13739), .C2(n14298), .A(n13551), .B(n13550), .ZN(
        n13552) );
  AOI21_X1 U15537 ( .B1(n13742), .B2(n13977), .A(n13552), .ZN(n13553) );
  OAI21_X1 U15538 ( .B1(n13743), .B2(n13675), .A(n13553), .ZN(P1_U3356) );
  OAI21_X1 U15539 ( .B1(n13560), .B2(n13559), .A(n13558), .ZN(n13748) );
  INV_X1 U15540 ( .A(n13748), .ZN(n13567) );
  AOI21_X1 U15541 ( .B1(n13745), .B2(n13577), .A(n14352), .ZN(n13562) );
  NAND2_X1 U15542 ( .A1(n13744), .A2(n14313), .ZN(n13565) );
  AOI22_X1 U15543 ( .A1(n14322), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n13563), 
        .B2(n14311), .ZN(n13564) );
  OAI211_X1 U15544 ( .C1(n6825), .C2(n14298), .A(n13565), .B(n13564), .ZN(
        n13566) );
  AOI21_X1 U15545 ( .B1(n13567), .B2(n14308), .A(n13566), .ZN(n13568) );
  OAI21_X1 U15546 ( .B1(n13747), .B2(n14322), .A(n13568), .ZN(P1_U3265) );
  OAI21_X1 U15547 ( .B1(n13576), .B2(n13570), .A(n13569), .ZN(n13573) );
  INV_X1 U15548 ( .A(n13571), .ZN(n13572) );
  AOI21_X1 U15549 ( .B1(n13573), .B2(n14373), .A(n13572), .ZN(n13752) );
  INV_X1 U15550 ( .A(n13753), .ZN(n13584) );
  AOI21_X1 U15551 ( .B1(n13750), .B2(n13592), .A(n14352), .ZN(n13578) );
  AND2_X1 U15552 ( .A1(n13578), .A2(n13577), .ZN(n13749) );
  NAND2_X1 U15553 ( .A1(n13749), .A2(n14313), .ZN(n13581) );
  AOI22_X1 U15554 ( .A1(n14322), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n13579), 
        .B2(n14311), .ZN(n13580) );
  OAI211_X1 U15555 ( .C1(n13582), .C2(n14298), .A(n13581), .B(n13580), .ZN(
        n13583) );
  AOI21_X1 U15556 ( .B1(n13584), .B2(n14308), .A(n13583), .ZN(n13585) );
  OAI21_X1 U15557 ( .B1(n13752), .B2(n14322), .A(n13585), .ZN(P1_U3266) );
  OAI21_X1 U15558 ( .B1(n13588), .B2(n13587), .A(n13586), .ZN(n13760) );
  OAI21_X1 U15559 ( .B1(n13591), .B2(n13590), .A(n13589), .ZN(n13758) );
  INV_X1 U15560 ( .A(n13606), .ZN(n13593) );
  OAI211_X1 U15561 ( .C1(n13756), .C2(n13593), .A(n9843), .B(n13592), .ZN(
        n13755) );
  INV_X1 U15562 ( .A(n13594), .ZN(n13595) );
  OAI22_X1 U15563 ( .A1(n14315), .A2(n13754), .B1(n13595), .B2(n14093), .ZN(
        n13597) );
  NOR2_X1 U15564 ( .A1(n13756), .A2(n14298), .ZN(n13596) );
  AOI211_X1 U15565 ( .C1(n14322), .C2(P1_REG2_REG_26__SCAN_IN), .A(n13597), 
        .B(n13596), .ZN(n13598) );
  OAI21_X1 U15566 ( .B1(n13720), .B2(n13755), .A(n13598), .ZN(n13599) );
  AOI21_X1 U15567 ( .B1(n13758), .B2(n13977), .A(n13599), .ZN(n13600) );
  OAI21_X1 U15568 ( .B1(n13675), .B2(n13760), .A(n13600), .ZN(P1_U3267) );
  XNOR2_X1 U15569 ( .A(n13602), .B(n13601), .ZN(n13770) );
  NOR2_X1 U15570 ( .A1(n13604), .A2(n13603), .ZN(n13761) );
  NOR2_X1 U15571 ( .A1(n13761), .A2(n13675), .ZN(n13620) );
  NAND2_X1 U15572 ( .A1(n13763), .A2(n13629), .ZN(n13605) );
  NAND2_X1 U15573 ( .A1(n13606), .A2(n13605), .ZN(n13765) );
  OR2_X1 U15574 ( .A1(n13607), .A2(n13963), .ZN(n13610) );
  NAND2_X1 U15575 ( .A1(n13608), .A2(n6454), .ZN(n13609) );
  NAND2_X1 U15576 ( .A1(n13610), .A2(n13609), .ZN(n13762) );
  INV_X1 U15577 ( .A(n13762), .ZN(n13615) );
  NAND2_X1 U15578 ( .A1(n14315), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13614) );
  INV_X1 U15579 ( .A(n13611), .ZN(n13612) );
  OR2_X1 U15580 ( .A1(n14093), .A2(n13612), .ZN(n13613) );
  OAI211_X1 U15581 ( .C1(n14322), .C2(n13615), .A(n13614), .B(n13613), .ZN(
        n13616) );
  AOI21_X1 U15582 ( .B1(n13763), .B2(n14310), .A(n13616), .ZN(n13617) );
  OAI21_X1 U15583 ( .B1(n13765), .B2(n13618), .A(n13617), .ZN(n13619) );
  AOI21_X1 U15584 ( .B1(n13620), .B2(n13767), .A(n13619), .ZN(n13621) );
  OAI21_X1 U15585 ( .B1(n13770), .B2(n13705), .A(n13621), .ZN(P1_U3268) );
  OAI211_X1 U15586 ( .C1(n13624), .C2(n13623), .A(n13622), .B(n14373), .ZN(
        n13626) );
  NAND2_X1 U15587 ( .A1(n13626), .A2(n13625), .ZN(n13773) );
  INV_X1 U15588 ( .A(n13773), .ZN(n13636) );
  OAI21_X1 U15589 ( .B1(n6518), .B2(n13628), .A(n13627), .ZN(n13775) );
  OAI211_X1 U15590 ( .C1(n13772), .C2(n13641), .A(n9843), .B(n13629), .ZN(
        n13771) );
  AOI22_X1 U15591 ( .A1(n14315), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n13630), 
        .B2(n14311), .ZN(n13633) );
  NAND2_X1 U15592 ( .A1(n13631), .A2(n14310), .ZN(n13632) );
  OAI211_X1 U15593 ( .C1(n13771), .C2(n13720), .A(n13633), .B(n13632), .ZN(
        n13634) );
  AOI21_X1 U15594 ( .B1(n13775), .B2(n14308), .A(n13634), .ZN(n13635) );
  OAI21_X1 U15595 ( .B1(n13636), .B2(n14322), .A(n13635), .ZN(P1_U3269) );
  AOI21_X1 U15596 ( .B1(n13639), .B2(n13638), .A(n13637), .ZN(n13783) );
  AND2_X1 U15597 ( .A1(n13778), .A2(n13655), .ZN(n13640) );
  INV_X1 U15598 ( .A(n13642), .ZN(n13777) );
  AOI22_X1 U15599 ( .A1(n13777), .A2(n13970), .B1(n13643), .B2(n14311), .ZN(
        n13645) );
  NAND2_X1 U15600 ( .A1(n14315), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n13644) );
  OAI211_X1 U15601 ( .C1(n13646), .C2(n14298), .A(n13645), .B(n13644), .ZN(
        n13647) );
  AOI21_X1 U15602 ( .B1(n7607), .B2(n14313), .A(n13647), .ZN(n13651) );
  NAND2_X1 U15603 ( .A1(n13649), .A2(n13648), .ZN(n13779) );
  NAND3_X1 U15604 ( .A1(n13780), .A2(n13779), .A3(n14308), .ZN(n13650) );
  OAI211_X1 U15605 ( .C1(n13783), .C2(n13705), .A(n13651), .B(n13650), .ZN(
        P1_U3270) );
  XNOR2_X1 U15606 ( .A(n13652), .B(n13654), .ZN(n13790) );
  XNOR2_X1 U15607 ( .A(n13653), .B(n13654), .ZN(n13788) );
  AOI21_X1 U15608 ( .B1(n13668), .B2(n13661), .A(n14352), .ZN(n13656) );
  NAND2_X1 U15609 ( .A1(n13656), .A2(n13655), .ZN(n13785) );
  NAND2_X1 U15610 ( .A1(n13657), .A2(n14311), .ZN(n13659) );
  NAND2_X1 U15611 ( .A1(n14315), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n13658) );
  OAI211_X1 U15612 ( .C1(n13784), .C2(n14315), .A(n13659), .B(n13658), .ZN(
        n13660) );
  AOI21_X1 U15613 ( .B1(n13661), .B2(n14310), .A(n13660), .ZN(n13662) );
  OAI21_X1 U15614 ( .B1(n13785), .B2(n13720), .A(n13662), .ZN(n13663) );
  AOI21_X1 U15615 ( .B1(n13788), .B2(n14308), .A(n13663), .ZN(n13664) );
  OAI21_X1 U15616 ( .B1(n13790), .B2(n13705), .A(n13664), .ZN(P1_U3271) );
  XOR2_X1 U15617 ( .A(n13667), .B(n13665), .Z(n13797) );
  XOR2_X1 U15618 ( .A(n13667), .B(n13666), .Z(n13795) );
  OAI211_X1 U15619 ( .C1(n7028), .C2(n13793), .A(n9843), .B(n13668), .ZN(
        n13792) );
  OAI22_X1 U15620 ( .A1(n13791), .A2(n14322), .B1(n13669), .B2(n14093), .ZN(
        n13671) );
  NOR2_X1 U15621 ( .A1(n13793), .A2(n14298), .ZN(n13670) );
  AOI211_X1 U15622 ( .C1(n14322), .C2(P1_REG2_REG_21__SCAN_IN), .A(n13671), 
        .B(n13670), .ZN(n13672) );
  OAI21_X1 U15623 ( .B1(n13720), .B2(n13792), .A(n13672), .ZN(n13673) );
  AOI21_X1 U15624 ( .B1(n13795), .B2(n13977), .A(n13673), .ZN(n13674) );
  OAI21_X1 U15625 ( .B1(n13675), .B2(n13797), .A(n13674), .ZN(P1_U3272) );
  OAI211_X1 U15626 ( .C1(n13677), .C2(n13684), .A(n13676), .B(n14373), .ZN(
        n13680) );
  AOI22_X1 U15627 ( .A1(n13678), .A2(n6454), .B1(n14087), .B2(n13709), .ZN(
        n13679) );
  NAND2_X1 U15628 ( .A1(n13680), .A2(n13679), .ZN(n13800) );
  INV_X1 U15629 ( .A(n13800), .ZN(n13692) );
  INV_X1 U15630 ( .A(n13681), .ZN(n13682) );
  AOI21_X1 U15631 ( .B1(n13684), .B2(n13683), .A(n13682), .ZN(n13802) );
  OAI211_X1 U15632 ( .C1(n13799), .C2(n13686), .A(n9843), .B(n13685), .ZN(
        n13798) );
  NOR2_X1 U15633 ( .A1(n13798), .A2(n13720), .ZN(n13690) );
  AOI22_X1 U15634 ( .A1(n14315), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n13687), 
        .B2(n14311), .ZN(n13688) );
  OAI21_X1 U15635 ( .B1(n13799), .B2(n14298), .A(n13688), .ZN(n13689) );
  AOI211_X1 U15636 ( .C1(n13802), .C2(n14308), .A(n13690), .B(n13689), .ZN(
        n13691) );
  OAI21_X1 U15637 ( .B1(n14322), .B2(n13692), .A(n13691), .ZN(P1_U3273) );
  AOI21_X1 U15638 ( .B1(n13701), .B2(n13694), .A(n13693), .ZN(n14105) );
  OAI21_X1 U15639 ( .B1(n13695), .B2(n14093), .A(n14102), .ZN(n13696) );
  MUX2_X1 U15640 ( .A(n13696), .B(P1_REG2_REG_19__SCAN_IN), .S(n14322), .Z(
        n13699) );
  XNOR2_X1 U15641 ( .A(n13715), .B(n13700), .ZN(n13697) );
  NAND2_X1 U15642 ( .A1(n13697), .A2(n9843), .ZN(n14103) );
  NOR2_X1 U15643 ( .A1(n14103), .A2(n13720), .ZN(n13698) );
  AOI211_X1 U15644 ( .C1(n14310), .C2(n13700), .A(n13699), .B(n13698), .ZN(
        n13704) );
  XNOR2_X1 U15645 ( .A(n13702), .B(n13701), .ZN(n14108) );
  NAND2_X1 U15646 ( .A1(n14108), .A2(n14308), .ZN(n13703) );
  OAI211_X1 U15647 ( .C1(n14105), .C2(n13705), .A(n13704), .B(n13703), .ZN(
        P1_U3274) );
  XNOR2_X1 U15648 ( .A(n13706), .B(n13707), .ZN(n14113) );
  XNOR2_X1 U15649 ( .A(n6489), .B(n13707), .ZN(n13708) );
  NAND2_X1 U15650 ( .A1(n13708), .A2(n14373), .ZN(n13711) );
  AOI22_X1 U15651 ( .A1(n13709), .A2(n6454), .B1(n14087), .B2(n14086), .ZN(
        n13710) );
  NAND2_X1 U15652 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  AOI21_X1 U15653 ( .B1(n14113), .B2(n14403), .A(n13712), .ZN(n14115) );
  NAND2_X1 U15654 ( .A1(n6482), .A2(n13717), .ZN(n13713) );
  NAND2_X1 U15655 ( .A1(n13713), .A2(n9843), .ZN(n13714) );
  OR2_X1 U15656 ( .A1(n13715), .A2(n13714), .ZN(n14110) );
  AOI22_X1 U15657 ( .A1(n14315), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n13716), 
        .B2(n14311), .ZN(n13719) );
  NAND2_X1 U15658 ( .A1(n13717), .A2(n14310), .ZN(n13718) );
  OAI211_X1 U15659 ( .C1(n14110), .C2(n13720), .A(n13719), .B(n13718), .ZN(
        n13721) );
  AOI21_X1 U15660 ( .B1(n14113), .B2(n14304), .A(n13721), .ZN(n13722) );
  OAI21_X1 U15661 ( .B1(n14115), .B2(n14322), .A(n13722), .ZN(P1_U3275) );
  OAI21_X1 U15662 ( .B1(n14308), .B2(n13977), .A(n13723), .ZN(n13730) );
  OAI21_X1 U15663 ( .B1(n14310), .B2(n13725), .A(n13724), .ZN(n13729) );
  AOI22_X1 U15664 ( .A1(n13970), .A2(n13726), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n14311), .ZN(n13728) );
  NAND2_X1 U15665 ( .A1(n14315), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n13727) );
  NAND4_X1 U15666 ( .A1(n13730), .A2(n13729), .A3(n13728), .A4(n13727), .ZN(
        P1_U3293) );
  NAND2_X1 U15667 ( .A1(n13731), .A2(n9843), .ZN(n13732) );
  OAI211_X1 U15668 ( .C1(n13733), .C2(n14417), .A(n13732), .B(n13734), .ZN(
        n13804) );
  MUX2_X1 U15669 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n13804), .S(n14441), .Z(
        P1_U3559) );
  OAI211_X1 U15670 ( .C1(n13736), .C2(n14417), .A(n13735), .B(n13734), .ZN(
        n13805) );
  MUX2_X1 U15671 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n13805), .S(n14441), .Z(
        P1_U3558) );
  OAI211_X1 U15672 ( .C1(n13739), .C2(n14417), .A(n13738), .B(n13737), .ZN(
        n13740) );
  MUX2_X1 U15673 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n13806), .S(n14441), .Z(
        P1_U3557) );
  OAI211_X1 U15674 ( .C1(n14368), .C2(n13748), .A(n13747), .B(n13746), .ZN(
        n13807) );
  MUX2_X1 U15675 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n13807), .S(n14441), .Z(
        P1_U3556) );
  AOI21_X1 U15676 ( .B1(n14397), .B2(n13750), .A(n13749), .ZN(n13751) );
  OAI211_X1 U15677 ( .C1(n14368), .C2(n13753), .A(n13752), .B(n13751), .ZN(
        n13808) );
  MUX2_X1 U15678 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n13808), .S(n14441), .Z(
        P1_U3555) );
  OAI211_X1 U15679 ( .C1(n13756), .C2(n14417), .A(n13755), .B(n13754), .ZN(
        n13757) );
  AOI21_X1 U15680 ( .B1(n13758), .B2(n14373), .A(n13757), .ZN(n13759) );
  OAI21_X1 U15681 ( .B1(n14368), .B2(n13760), .A(n13759), .ZN(n13809) );
  MUX2_X1 U15682 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n13809), .S(n14441), .Z(
        P1_U3554) );
  NOR2_X1 U15683 ( .A1(n13761), .A2(n14368), .ZN(n13768) );
  AOI21_X1 U15684 ( .B1(n13763), .B2(n14397), .A(n13762), .ZN(n13764) );
  OAI21_X1 U15685 ( .B1(n13765), .B2(n14352), .A(n13764), .ZN(n13766) );
  AOI21_X1 U15686 ( .B1(n13768), .B2(n13767), .A(n13766), .ZN(n13769) );
  OAI21_X1 U15687 ( .B1(n13770), .B2(n14379), .A(n13769), .ZN(n13810) );
  MUX2_X1 U15688 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n13810), .S(n14441), .Z(
        P1_U3553) );
  OAI21_X1 U15689 ( .B1(n13772), .B2(n14417), .A(n13771), .ZN(n13774) );
  AOI211_X1 U15690 ( .C1(n14421), .C2(n13775), .A(n13774), .B(n13773), .ZN(
        n13776) );
  INV_X1 U15691 ( .A(n13776), .ZN(n13811) );
  MUX2_X1 U15692 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n13811), .S(n14441), .Z(
        P1_U3552) );
  AOI211_X1 U15693 ( .C1(n14397), .C2(n13778), .A(n13777), .B(n7607), .ZN(
        n13782) );
  NAND3_X1 U15694 ( .A1(n13780), .A2(n13779), .A3(n14421), .ZN(n13781) );
  OAI211_X1 U15695 ( .C1(n13783), .C2(n14379), .A(n13782), .B(n13781), .ZN(
        n13812) );
  MUX2_X1 U15696 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n13812), .S(n14441), .Z(
        P1_U3551) );
  OAI211_X1 U15697 ( .C1(n14417), .C2(n13786), .A(n13785), .B(n13784), .ZN(
        n13787) );
  AOI21_X1 U15698 ( .B1(n13788), .B2(n14421), .A(n13787), .ZN(n13789) );
  OAI21_X1 U15699 ( .B1(n13790), .B2(n14379), .A(n13789), .ZN(n13813) );
  MUX2_X1 U15700 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n13813), .S(n14441), .Z(
        P1_U3550) );
  OAI211_X1 U15701 ( .C1(n13793), .C2(n14417), .A(n13792), .B(n13791), .ZN(
        n13794) );
  AOI21_X1 U15702 ( .B1(n13795), .B2(n14373), .A(n13794), .ZN(n13796) );
  OAI21_X1 U15703 ( .B1(n14368), .B2(n13797), .A(n13796), .ZN(n13814) );
  MUX2_X1 U15704 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n13814), .S(n14441), .Z(
        P1_U3549) );
  OAI21_X1 U15705 ( .B1(n13799), .B2(n14417), .A(n13798), .ZN(n13801) );
  AOI211_X1 U15706 ( .C1(n13802), .C2(n14421), .A(n13801), .B(n13800), .ZN(
        n13803) );
  INV_X1 U15707 ( .A(n13803), .ZN(n13815) );
  MUX2_X1 U15708 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n13815), .S(n14441), .Z(
        P1_U3548) );
  MUX2_X1 U15709 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n13804), .S(n14425), .Z(
        P1_U3527) );
  MUX2_X1 U15710 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n13805), .S(n14425), .Z(
        P1_U3526) );
  MUX2_X1 U15711 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n13806), .S(n14425), .Z(
        P1_U3525) );
  MUX2_X1 U15712 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n13807), .S(n14425), .Z(
        P1_U3524) );
  MUX2_X1 U15713 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n13808), .S(n14425), .Z(
        P1_U3523) );
  MUX2_X1 U15714 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n13809), .S(n14425), .Z(
        P1_U3522) );
  MUX2_X1 U15715 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n13810), .S(n14425), .Z(
        P1_U3521) );
  MUX2_X1 U15716 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n13811), .S(n14425), .Z(
        P1_U3520) );
  MUX2_X1 U15717 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n13812), .S(n14425), .Z(
        P1_U3519) );
  MUX2_X1 U15718 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n13813), .S(n14425), .Z(
        P1_U3518) );
  MUX2_X1 U15719 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n13814), .S(n14425), .Z(
        P1_U3517) );
  MUX2_X1 U15720 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n13815), .S(n14425), .Z(
        P1_U3516) );
  NOR4_X1 U15721 ( .A1(n13817), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), 
        .A4(n13816), .ZN(n13818) );
  AOI21_X1 U15722 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(n13819), .A(n13818), 
        .ZN(n13820) );
  OAI21_X1 U15723 ( .B1(n13821), .B2(n13837), .A(n13820), .ZN(P1_U3324) );
  OAI222_X1 U15724 ( .A1(n13837), .A2(n13824), .B1(n13823), .B2(P1_U3086), 
        .C1(n13822), .C2(n13833), .ZN(P1_U3325) );
  OAI222_X1 U15725 ( .A1(n13837), .A2(n13827), .B1(n13826), .B2(P1_U3086), 
        .C1(n13825), .C2(n13833), .ZN(P1_U3326) );
  OAI222_X1 U15726 ( .A1(n13833), .A2(n13830), .B1(n13837), .B2(n13829), .C1(
        P1_U3086), .C2(n13828), .ZN(P1_U3327) );
  OAI222_X1 U15727 ( .A1(n13837), .A2(n13832), .B1(n8530), .B2(P1_U3086), .C1(
        n13831), .C2(n13833), .ZN(P1_U3328) );
  OAI222_X1 U15728 ( .A1(n13837), .A2(n13836), .B1(P1_U3086), .B2(n13835), 
        .C1(n13834), .C2(n13833), .ZN(P1_U3329) );
  MUX2_X1 U15729 ( .A(n13839), .B(n13838), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  MUX2_X1 U15730 ( .A(n13840), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15731 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14252) );
  AND2_X1 U15732 ( .A1(n14252), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n13865) );
  INV_X1 U15733 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14235) );
  NOR2_X1 U15734 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14235), .ZN(n13864) );
  INV_X1 U15735 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14206) );
  XOR2_X1 U15736 ( .A(n14913), .B(P1_ADDR_REG_12__SCAN_IN), .Z(n13922) );
  XOR2_X1 U15737 ( .A(n14698), .B(P1_ADDR_REG_9__SCAN_IN), .Z(n13915) );
  INV_X1 U15738 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n13855) );
  INV_X1 U15739 ( .A(n13889), .ZN(n13888) );
  XNOR2_X1 U15740 ( .A(n14986), .B(P3_ADDR_REG_2__SCAN_IN), .ZN(n13885) );
  NOR2_X1 U15741 ( .A1(n13845), .A2(n6941), .ZN(n13847) );
  NOR2_X1 U15742 ( .A1(P3_ADDR_REG_6__SCAN_IN), .A2(n13903), .ZN(n13849) );
  INV_X1 U15743 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n13848) );
  NOR2_X1 U15744 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n13850), .ZN(n13852) );
  XNOR2_X1 U15745 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n13850), .ZN(n13907) );
  XNOR2_X1 U15746 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(n13853), .ZN(n13880) );
  NAND2_X1 U15747 ( .A1(n13915), .A2(n13914), .ZN(n13856) );
  NOR2_X1 U15748 ( .A1(n13877), .A2(n13878), .ZN(n13858) );
  INV_X1 U15749 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n14723) );
  NAND2_X1 U15750 ( .A1(n13877), .A2(n13878), .ZN(n13857) );
  XNOR2_X1 U15751 ( .A(n13860), .B(P1_ADDR_REG_11__SCAN_IN), .ZN(n13875) );
  NAND2_X1 U15752 ( .A1(n13922), .A2(n13921), .ZN(n13861) );
  INV_X1 U15753 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n14960) );
  NAND2_X1 U15754 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n14960), .ZN(n13862) );
  XOR2_X1 U15755 ( .A(n14916), .B(P3_ADDR_REG_14__SCAN_IN), .Z(n13872) );
  NAND2_X1 U15756 ( .A1(n13871), .A2(n13872), .ZN(n13863) );
  OAI22_X1 U15757 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(n14930), .B1(n13864), 
        .B2(n13870), .ZN(n13931) );
  OAI22_X1 U15758 ( .A1(n13865), .A2(n13931), .B1(P3_ADDR_REG_16__SCAN_IN), 
        .B2(n14252), .ZN(n13866) );
  NOR2_X1 U15759 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n13866), .ZN(n13868) );
  INV_X1 U15760 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14269) );
  XNOR2_X1 U15761 ( .A(n14269), .B(n13866), .ZN(n13935) );
  AND2_X1 U15762 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n13935), .ZN(n13867) );
  NOR2_X1 U15763 ( .A1(n13868), .A2(n13867), .ZN(n13990) );
  INV_X1 U15764 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14289) );
  XNOR2_X1 U15765 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n14289), .ZN(n13989) );
  XNOR2_X1 U15766 ( .A(n13990), .B(n13989), .ZN(n13937) );
  XNOR2_X1 U15767 ( .A(n14930), .B(P1_ADDR_REG_15__SCAN_IN), .ZN(n13869) );
  XOR2_X1 U15768 ( .A(n13870), .B(n13869), .Z(n13927) );
  INV_X1 U15769 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14500) );
  XOR2_X1 U15770 ( .A(n13872), .B(n13871), .Z(n14181) );
  INV_X1 U15771 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n13926) );
  XOR2_X1 U15772 ( .A(n14960), .B(P1_ADDR_REG_13__SCAN_IN), .Z(n13874) );
  XNOR2_X1 U15773 ( .A(n13874), .B(n13873), .ZN(n14178) );
  INV_X1 U15774 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n13920) );
  XOR2_X1 U15775 ( .A(n13876), .B(n13875), .Z(n14173) );
  INV_X1 U15776 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14489) );
  XOR2_X1 U15777 ( .A(n13877), .B(P3_ADDR_REG_10__SCAN_IN), .Z(n13879) );
  XNOR2_X1 U15778 ( .A(n13879), .B(n13878), .ZN(n13953) );
  XOR2_X1 U15779 ( .A(n13881), .B(n13880), .Z(n13913) );
  OR2_X1 U15780 ( .A1(n13883), .A2(n13884), .ZN(n13897) );
  INV_X1 U15781 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14454) );
  INV_X1 U15782 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14965) );
  XNOR2_X1 U15783 ( .A(n13885), .B(n13886), .ZN(n13941) );
  XNOR2_X1 U15784 ( .A(n13888), .B(n13887), .ZN(n13890) );
  NAND2_X1 U15785 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n13890), .ZN(n13892) );
  AOI21_X1 U15786 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n9671), .A(n13889), .ZN(
        n15029) );
  INV_X1 U15787 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15028) );
  NOR2_X1 U15788 ( .A1(n15029), .A2(n15028), .ZN(n15037) );
  NAND2_X1 U15789 ( .A1(n13892), .A2(n13891), .ZN(n13942) );
  NAND2_X1 U15790 ( .A1(n13941), .A2(n13942), .ZN(n13893) );
  NOR2_X1 U15791 ( .A1(n13941), .A2(n13942), .ZN(n13940) );
  XOR2_X1 U15792 ( .A(n6843), .B(n13894), .Z(n15033) );
  NAND2_X1 U15793 ( .A1(n15034), .A2(n15033), .ZN(n13895) );
  NOR2_X1 U15794 ( .A1(n15034), .A2(n15033), .ZN(n15032) );
  AOI21_X1 U15795 ( .B1(n14454), .B2(n13895), .A(n15032), .ZN(n15024) );
  NAND2_X1 U15796 ( .A1(n13902), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n13906) );
  XNOR2_X1 U15797 ( .A(n13903), .B(P3_ADDR_REG_6__SCAN_IN), .ZN(n13904) );
  XNOR2_X1 U15798 ( .A(n13905), .B(n13904), .ZN(n13944) );
  NAND2_X1 U15799 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n13908), .ZN(n13911) );
  XOR2_X1 U15800 ( .A(n14911), .B(n13907), .Z(n15031) );
  XNOR2_X1 U15801 ( .A(n13915), .B(n13914), .ZN(n13917) );
  NAND2_X1 U15802 ( .A1(n13916), .A2(n13917), .ZN(n13918) );
  NAND2_X1 U15803 ( .A1(n14173), .A2(n14174), .ZN(n13919) );
  NOR2_X1 U15804 ( .A1(n14173), .A2(n14174), .ZN(n14172) );
  XNOR2_X1 U15805 ( .A(n13922), .B(n13921), .ZN(n13924) );
  NAND2_X1 U15806 ( .A1(n14178), .A2(n14179), .ZN(n13925) );
  XOR2_X1 U15807 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n14252), .Z(n13932) );
  XOR2_X1 U15808 ( .A(n13932), .B(n13931), .Z(n13933) );
  XNOR2_X1 U15809 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n13935), .ZN(n13984) );
  INV_X1 U15810 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14541) );
  AOI21_X1 U15811 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n13938) );
  OAI21_X1 U15812 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n13938), 
        .ZN(U28) );
  AOI21_X1 U15813 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n13939) );
  OAI21_X1 U15814 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n13939), 
        .ZN(U29) );
  AOI21_X1 U15815 ( .B1(n13942), .B2(n13941), .A(n13940), .ZN(n13943) );
  XOR2_X1 U15816 ( .A(n13943), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U15817 ( .A(n13945), .B(n13944), .Z(SUB_1596_U57) );
  INV_X1 U15818 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n14477) );
  XOR2_X1 U15819 ( .A(n14477), .B(n13946), .Z(SUB_1596_U55) );
  AOI22_X1 U15820 ( .A1(n13949), .A2(n13948), .B1(SI_18_), .B2(n13947), .ZN(
        n13950) );
  OAI21_X1 U15821 ( .B1(P3_U3151), .B2(n13951), .A(n13950), .ZN(P3_U3277) );
  XOR2_X1 U15822 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n13952), .Z(SUB_1596_U54) );
  AOI21_X1 U15823 ( .B1(n13954), .B2(n13953), .A(n6622), .ZN(n13955) );
  XOR2_X1 U15824 ( .A(n13955), .B(P2_ADDR_REG_10__SCAN_IN), .Z(SUB_1596_U70)
         );
  INV_X1 U15825 ( .A(n14400), .ZN(n14392) );
  OAI21_X1 U15826 ( .B1(n13957), .B2(n14417), .A(n13956), .ZN(n13959) );
  AOI211_X1 U15827 ( .C1(n14392), .C2(n13960), .A(n13959), .B(n13958), .ZN(
        n13962) );
  INV_X1 U15828 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U15829 ( .A1(n14425), .A2(n13962), .B1(n13961), .B2(n14423), .ZN(
        P1_U3495) );
  AOI22_X1 U15830 ( .A1(n14441), .A2(n13962), .B1(n9600), .B2(n14438), .ZN(
        P1_U3540) );
  INV_X1 U15831 ( .A(n14145), .ZN(n13968) );
  OAI22_X1 U15832 ( .A1(n13966), .A2(n13965), .B1(n13964), .B2(n13963), .ZN(
        n14144) );
  INV_X1 U15833 ( .A(n14144), .ZN(n13967) );
  OAI211_X1 U15834 ( .C1(n13968), .C2(n14094), .A(n13967), .B(n13970), .ZN(
        n13969) );
  OAI21_X1 U15835 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n13970), .A(n13969), 
        .ZN(n13980) );
  XNOR2_X1 U15836 ( .A(n13972), .B(n13971), .ZN(n14149) );
  XNOR2_X1 U15837 ( .A(n13973), .B(n14145), .ZN(n13974) );
  NOR2_X1 U15838 ( .A1(n13974), .A2(n14352), .ZN(n14143) );
  XNOR2_X1 U15839 ( .A(n13976), .B(n13975), .ZN(n14147) );
  INV_X1 U15840 ( .A(n14147), .ZN(n13978) );
  AOI222_X1 U15841 ( .A1(n14308), .A2(n14149), .B1(n14313), .B2(n14143), .C1(
        n13978), .C2(n13977), .ZN(n13979) );
  OAI211_X1 U15842 ( .C1(n13981), .C2(n14093), .A(n13980), .B(n13979), .ZN(
        P1_U3280) );
  OAI21_X1 U15843 ( .B1(n13984), .B2(n13983), .A(n13982), .ZN(n13985) );
  XOR2_X1 U15844 ( .A(n13985), .B(n14541), .Z(SUB_1596_U63) );
  NOR2_X1 U15845 ( .A1(n13990), .A2(n13989), .ZN(n13991) );
  AOI21_X1 U15846 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n14289), .A(n13991), 
        .ZN(n13995) );
  XNOR2_X1 U15847 ( .A(n13992), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n13993) );
  XNOR2_X1 U15848 ( .A(n13993), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n13994) );
  XNOR2_X1 U15849 ( .A(n13995), .B(n13994), .ZN(n13996) );
  XNOR2_X1 U15850 ( .A(n13997), .B(n13996), .ZN(SUB_1596_U4) );
  AOI22_X1 U15851 ( .A1(n14686), .A2(n13998), .B1(n14664), .B2(
        P3_ADDR_REG_16__SCAN_IN), .ZN(n14014) );
  INV_X1 U15852 ( .A(n13999), .ZN(n14001) );
  NAND2_X1 U15853 ( .A1(n14001), .A2(n14000), .ZN(n14002) );
  XNOR2_X1 U15854 ( .A(n14003), .B(n14002), .ZN(n14008) );
  OAI21_X1 U15855 ( .B1(n14006), .B2(n14005), .A(n14004), .ZN(n14007) );
  AOI22_X1 U15856 ( .A1(n14008), .A2(n14713), .B1(n14703), .B2(n14007), .ZN(
        n14013) );
  OAI221_X1 U15857 ( .B1(n14010), .B2(n6526), .C1(n14010), .C2(n14009), .A(
        n14040), .ZN(n14011) );
  NAND4_X1 U15858 ( .A1(n14014), .A2(n14013), .A3(n14012), .A4(n14011), .ZN(
        P3_U3198) );
  AOI22_X1 U15859 ( .A1(n14686), .A2(n14015), .B1(n14664), .B2(
        P3_ADDR_REG_17__SCAN_IN), .ZN(n14028) );
  OAI21_X1 U15860 ( .B1(P3_REG1_REG_17__SCAN_IN), .B2(n14017), .A(n14016), 
        .ZN(n14022) );
  AOI211_X1 U15861 ( .C1(n14020), .C2(n14019), .A(n14036), .B(n14018), .ZN(
        n14021) );
  AOI21_X1 U15862 ( .B1(n14703), .B2(n14022), .A(n14021), .ZN(n14027) );
  NAND2_X1 U15863 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(P3_U3151), .ZN(n14026)
         );
  OAI221_X1 U15864 ( .B1(n14024), .B2(n14931), .C1(n14024), .C2(n14023), .A(
        n14040), .ZN(n14025) );
  NAND4_X1 U15865 ( .A1(n14028), .A2(n14027), .A3(n14026), .A4(n14025), .ZN(
        P3_U3199) );
  AOI22_X1 U15866 ( .A1(n14686), .A2(n14029), .B1(n14664), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14047) );
  OAI21_X1 U15867 ( .B1(n14032), .B2(n14031), .A(n14030), .ZN(n14039) );
  AOI21_X1 U15868 ( .B1(n14035), .B2(n14034), .A(n14033), .ZN(n14037) );
  NOR2_X1 U15869 ( .A1(n14037), .A2(n14036), .ZN(n14038) );
  AOI21_X1 U15870 ( .B1(n14703), .B2(n14039), .A(n14038), .ZN(n14046) );
  OAI221_X1 U15871 ( .B1(n14043), .B2(n14042), .C1(n14043), .C2(n14041), .A(
        n14040), .ZN(n14044) );
  NAND4_X1 U15872 ( .A1(n14047), .A2(n14046), .A3(n14045), .A4(n14044), .ZN(
        P3_U3200) );
  AOI22_X1 U15873 ( .A1(n14050), .A2(n14772), .B1(n14056), .B2(n14791), .ZN(
        n14054) );
  AOI22_X1 U15874 ( .A1(n12052), .A2(n6433), .B1(n14793), .B2(
        P3_REG2_REG_31__SCAN_IN), .ZN(n14051) );
  NAND2_X1 U15875 ( .A1(n14054), .A2(n14051), .ZN(P3_U3202) );
  AOI22_X1 U15876 ( .A1(n14057), .A2(n6433), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14793), .ZN(n14053) );
  NAND2_X1 U15877 ( .A1(n14054), .A2(n14053), .ZN(P3_U3203) );
  AOI21_X1 U15878 ( .B1(n12052), .B2(n14821), .A(n14056), .ZN(n14065) );
  INV_X1 U15879 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U15880 ( .A1(n14868), .A2(n14065), .B1(n14055), .B2(n14866), .ZN(
        P3_U3490) );
  AOI21_X1 U15881 ( .B1(n14057), .B2(n14821), .A(n14056), .ZN(n14067) );
  INV_X1 U15882 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14058) );
  AOI22_X1 U15883 ( .A1(n14868), .A2(n14067), .B1(n14058), .B2(n14866), .ZN(
        P3_U3489) );
  AOI21_X1 U15884 ( .B1(n14060), .B2(n14848), .A(n14059), .ZN(n14061) );
  AND2_X1 U15885 ( .A1(n14062), .A2(n14061), .ZN(n14069) );
  INV_X1 U15886 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U15887 ( .A1(n14868), .A2(n14069), .B1(n14063), .B2(n14866), .ZN(
        P3_U3470) );
  INV_X1 U15888 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U15889 ( .A1(n14851), .A2(n14065), .B1(n14064), .B2(n14849), .ZN(
        P3_U3458) );
  INV_X1 U15890 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n14066) );
  AOI22_X1 U15891 ( .A1(n14851), .A2(n14067), .B1(n14066), .B2(n14849), .ZN(
        P3_U3457) );
  INV_X1 U15892 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14068) );
  AOI22_X1 U15893 ( .A1(n14851), .A2(n14069), .B1(n14068), .B2(n14849), .ZN(
        P3_U3423) );
  AOI21_X1 U15894 ( .B1(n14072), .B2(n14070), .A(n14071), .ZN(n14079) );
  AOI22_X1 U15895 ( .A1(n14074), .A2(n14086), .B1(n14073), .B2(n14088), .ZN(
        n14077) );
  NAND2_X1 U15896 ( .A1(n14089), .A2(n14075), .ZN(n14076) );
  OAI211_X1 U15897 ( .C1(n14079), .C2(n14078), .A(n14077), .B(n14076), .ZN(
        n14080) );
  INV_X1 U15898 ( .A(n14080), .ZN(n14082) );
  NAND2_X1 U15899 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(P1_U3086), .ZN(n14250)
         );
  OAI211_X1 U15900 ( .C1(n14083), .C2(n14092), .A(n14082), .B(n14250), .ZN(
        P1_U3226) );
  XNOR2_X1 U15901 ( .A(n14084), .B(n14099), .ZN(n14085) );
  AOI222_X1 U15902 ( .A1(n14088), .A2(n14087), .B1(n14086), .B2(n6454), .C1(
        n14373), .C2(n14085), .ZN(n14127) );
  INV_X1 U15903 ( .A(n14127), .ZN(n14097) );
  NAND2_X1 U15904 ( .A1(n14090), .A2(n14089), .ZN(n14125) );
  AND3_X1 U15905 ( .A1(n14125), .A2(n14091), .A3(n14124), .ZN(n14096) );
  OAI22_X1 U15906 ( .A1(n14128), .A2(n14094), .B1(n14093), .B2(n14092), .ZN(
        n14095) );
  NOR3_X1 U15907 ( .A1(n14097), .A2(n14096), .A3(n14095), .ZN(n14101) );
  XNOR2_X1 U15908 ( .A(n14098), .B(n14099), .ZN(n14130) );
  AOI22_X1 U15909 ( .A1(n14130), .A2(n14308), .B1(P1_REG2_REG_16__SCAN_IN), 
        .B2(n14322), .ZN(n14100) );
  OAI21_X1 U15910 ( .B1(n14322), .B2(n14101), .A(n14100), .ZN(P1_U3277) );
  OAI211_X1 U15911 ( .C1(n14104), .C2(n14417), .A(n14103), .B(n14102), .ZN(
        n14107) );
  NOR2_X1 U15912 ( .A1(n14105), .A2(n14379), .ZN(n14106) );
  AOI211_X1 U15913 ( .C1(n14108), .C2(n14421), .A(n14107), .B(n14106), .ZN(
        n14157) );
  AOI22_X1 U15914 ( .A1(n14441), .A2(n14157), .B1(n14109), .B2(n14438), .ZN(
        P1_U3547) );
  OAI21_X1 U15915 ( .B1(n14111), .B2(n14417), .A(n14110), .ZN(n14112) );
  AOI21_X1 U15916 ( .B1(n14113), .B2(n14392), .A(n14112), .ZN(n14114) );
  AND2_X1 U15917 ( .A1(n14115), .A2(n14114), .ZN(n14159) );
  AOI22_X1 U15918 ( .A1(n14441), .A2(n14159), .B1(n14270), .B2(n14438), .ZN(
        P1_U3546) );
  NAND2_X1 U15919 ( .A1(n14116), .A2(n14397), .ZN(n14117) );
  OAI211_X1 U15920 ( .C1(n14119), .C2(n14352), .A(n14118), .B(n14117), .ZN(
        n14122) );
  NOR2_X1 U15921 ( .A1(n14120), .A2(n14379), .ZN(n14121) );
  AOI211_X1 U15922 ( .C1(n14123), .C2(n14421), .A(n14122), .B(n14121), .ZN(
        n14161) );
  AOI22_X1 U15923 ( .A1(n14441), .A2(n14161), .B1(n13458), .B2(n14438), .ZN(
        P1_U3545) );
  NAND3_X1 U15924 ( .A1(n14125), .A2(n9843), .A3(n14124), .ZN(n14126) );
  OAI211_X1 U15925 ( .C1(n14128), .C2(n14417), .A(n14127), .B(n14126), .ZN(
        n14129) );
  AOI21_X1 U15926 ( .B1(n14130), .B2(n14421), .A(n14129), .ZN(n14163) );
  AOI22_X1 U15927 ( .A1(n14441), .A2(n14163), .B1(n13447), .B2(n14438), .ZN(
        P1_U3544) );
  OAI21_X1 U15928 ( .B1(n14132), .B2(n14417), .A(n14131), .ZN(n14134) );
  AOI211_X1 U15929 ( .C1(n14135), .C2(n14421), .A(n14134), .B(n14133), .ZN(
        n14165) );
  AOI22_X1 U15930 ( .A1(n14441), .A2(n14165), .B1(n14224), .B2(n14438), .ZN(
        P1_U3543) );
  AOI22_X1 U15931 ( .A1(n14137), .A2(n9843), .B1(n14397), .B2(n14136), .ZN(
        n14141) );
  NAND3_X1 U15932 ( .A1(n14139), .A2(n14138), .A3(n14421), .ZN(n14140) );
  AOI22_X1 U15933 ( .A1(n14441), .A2(n14167), .B1(n13450), .B2(n14438), .ZN(
        P1_U3542) );
  AOI211_X1 U15934 ( .C1(n14397), .C2(n14145), .A(n14144), .B(n14143), .ZN(
        n14146) );
  OAI21_X1 U15935 ( .B1(n14147), .B2(n14379), .A(n14146), .ZN(n14148) );
  AOI21_X1 U15936 ( .B1(n14149), .B2(n14421), .A(n14148), .ZN(n14169) );
  AOI22_X1 U15937 ( .A1(n14441), .A2(n14169), .B1(n13454), .B2(n14438), .ZN(
        P1_U3541) );
  OAI211_X1 U15938 ( .C1(n14152), .C2(n14417), .A(n14151), .B(n14150), .ZN(
        n14153) );
  AOI21_X1 U15939 ( .B1(n14154), .B2(n14421), .A(n14153), .ZN(n14171) );
  AOI22_X1 U15940 ( .A1(n14441), .A2(n14171), .B1(n14155), .B2(n14438), .ZN(
        P1_U3539) );
  INV_X1 U15941 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14156) );
  AOI22_X1 U15942 ( .A1(n14425), .A2(n14157), .B1(n14156), .B2(n14423), .ZN(
        P1_U3515) );
  INV_X1 U15943 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U15944 ( .A1(n14425), .A2(n14159), .B1(n14158), .B2(n14423), .ZN(
        P1_U3513) );
  INV_X1 U15945 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14160) );
  AOI22_X1 U15946 ( .A1(n14425), .A2(n14161), .B1(n14160), .B2(n14423), .ZN(
        P1_U3510) );
  INV_X1 U15947 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14162) );
  AOI22_X1 U15948 ( .A1(n14425), .A2(n14163), .B1(n14162), .B2(n14423), .ZN(
        P1_U3507) );
  INV_X1 U15949 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14164) );
  AOI22_X1 U15950 ( .A1(n14425), .A2(n14165), .B1(n14164), .B2(n14423), .ZN(
        P1_U3504) );
  INV_X1 U15951 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n14166) );
  AOI22_X1 U15952 ( .A1(n14425), .A2(n14167), .B1(n14166), .B2(n14423), .ZN(
        P1_U3501) );
  INV_X1 U15953 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14168) );
  AOI22_X1 U15954 ( .A1(n14425), .A2(n14169), .B1(n14168), .B2(n14423), .ZN(
        P1_U3498) );
  INV_X1 U15955 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U15956 ( .A1(n14425), .A2(n14171), .B1(n14170), .B2(n14423), .ZN(
        P1_U3492) );
  AOI21_X1 U15957 ( .B1(n14174), .B2(n14173), .A(n14172), .ZN(n14175) );
  XOR2_X1 U15958 ( .A(n14175), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U15959 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14176), .ZN(SUB_1596_U68)
         );
  AOI21_X1 U15960 ( .B1(n14179), .B2(n14178), .A(n14177), .ZN(n14180) );
  XOR2_X1 U15961 ( .A(n14180), .B(P2_ADDR_REG_13__SCAN_IN), .Z(SUB_1596_U67)
         );
  AOI21_X1 U15962 ( .B1(n14182), .B2(n14181), .A(n6589), .ZN(n14183) );
  XOR2_X1 U15963 ( .A(n14183), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  INV_X1 U15964 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14513) );
  NOR2_X1 U15965 ( .A1(n14185), .A2(n14184), .ZN(n14186) );
  XNOR2_X1 U15966 ( .A(n14513), .B(n14186), .ZN(SUB_1596_U65) );
  INV_X1 U15967 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U15968 ( .A1(n14188), .A2(n14187), .ZN(n14189) );
  XNOR2_X1 U15969 ( .A(n14525), .B(n14189), .ZN(SUB_1596_U64) );
  INV_X1 U15970 ( .A(n14190), .ZN(n14202) );
  NAND2_X1 U15971 ( .A1(n14192), .A2(n14191), .ZN(n14195) );
  NOR2_X1 U15972 ( .A1(n14284), .A2(n14193), .ZN(n14194) );
  NAND2_X1 U15973 ( .A1(n14195), .A2(n14194), .ZN(n14201) );
  NAND2_X1 U15974 ( .A1(n14197), .A2(n14196), .ZN(n14199) );
  NAND3_X1 U15975 ( .A1(n14199), .A2(n14280), .A3(n14198), .ZN(n14200) );
  OAI211_X1 U15976 ( .C1(n14231), .C2(n14202), .A(n14201), .B(n14200), .ZN(
        n14203) );
  INV_X1 U15977 ( .A(n14203), .ZN(n14205) );
  OAI211_X1 U15978 ( .C1(n14206), .C2(n14288), .A(n14205), .B(n14204), .ZN(
        P1_U3256) );
  OAI21_X1 U15979 ( .B1(n14209), .B2(n14208), .A(n14207), .ZN(n14210) );
  NAND2_X1 U15980 ( .A1(n14226), .A2(n14210), .ZN(n14217) );
  NAND2_X1 U15981 ( .A1(n14276), .A2(n14211), .ZN(n14216) );
  OAI211_X1 U15982 ( .C1(n14214), .C2(n14213), .A(n14280), .B(n14212), .ZN(
        n14215) );
  AND3_X1 U15983 ( .A1(n14217), .A2(n14216), .A3(n14215), .ZN(n14219) );
  OAI211_X1 U15984 ( .C1(n14916), .C2(n14288), .A(n14219), .B(n14218), .ZN(
        P1_U3257) );
  OAI21_X1 U15985 ( .B1(n14221), .B2(n11002), .A(n14220), .ZN(n14222) );
  NAND2_X1 U15986 ( .A1(n14222), .A2(n14280), .ZN(n14229) );
  OAI21_X1 U15987 ( .B1(n14225), .B2(n14224), .A(n14223), .ZN(n14227) );
  NAND2_X1 U15988 ( .A1(n14227), .A2(n14226), .ZN(n14228) );
  OAI211_X1 U15989 ( .C1(n14231), .C2(n14230), .A(n14229), .B(n14228), .ZN(
        n14232) );
  INV_X1 U15990 ( .A(n14232), .ZN(n14234) );
  OAI211_X1 U15991 ( .C1(n14235), .C2(n14288), .A(n14234), .B(n14233), .ZN(
        P1_U3258) );
  NAND2_X1 U15992 ( .A1(n14237), .A2(n14236), .ZN(n14242) );
  NOR2_X1 U15993 ( .A1(n14284), .A2(n14238), .ZN(n14241) );
  AND2_X1 U15994 ( .A1(n14276), .A2(n14239), .ZN(n14240) );
  AOI21_X1 U15995 ( .B1(n14242), .B2(n14241), .A(n14240), .ZN(n14249) );
  NAND2_X1 U15996 ( .A1(n14244), .A2(n14243), .ZN(n14247) );
  INV_X1 U15997 ( .A(n14245), .ZN(n14246) );
  NAND3_X1 U15998 ( .A1(n14247), .A2(n14280), .A3(n14246), .ZN(n14248) );
  AND2_X1 U15999 ( .A1(n14249), .A2(n14248), .ZN(n14251) );
  OAI211_X1 U16000 ( .C1(n14252), .C2(n14288), .A(n14251), .B(n14250), .ZN(
        P1_U3259) );
  INV_X1 U16001 ( .A(n14253), .ZN(n14257) );
  INV_X1 U16002 ( .A(n14254), .ZN(n14255) );
  OAI21_X1 U16003 ( .B1(n14257), .B2(n14256), .A(n14255), .ZN(n14265) );
  NAND2_X1 U16004 ( .A1(n14276), .A2(n14258), .ZN(n14264) );
  AOI21_X1 U16005 ( .B1(n14261), .B2(n14260), .A(n14259), .ZN(n14262) );
  NAND2_X1 U16006 ( .A1(n14280), .A2(n14262), .ZN(n14263) );
  OAI211_X1 U16007 ( .C1(n14284), .C2(n14265), .A(n14264), .B(n14263), .ZN(
        n14266) );
  INV_X1 U16008 ( .A(n14266), .ZN(n14268) );
  OAI211_X1 U16009 ( .C1(n14269), .C2(n14288), .A(n14268), .B(n14267), .ZN(
        P1_U3260) );
  NAND2_X1 U16010 ( .A1(n14271), .A2(n14270), .ZN(n14274) );
  INV_X1 U16011 ( .A(n14272), .ZN(n14273) );
  NAND2_X1 U16012 ( .A1(n14274), .A2(n14273), .ZN(n14283) );
  NAND2_X1 U16013 ( .A1(n14276), .A2(n14275), .ZN(n14282) );
  AOI21_X1 U16014 ( .B1(n14278), .B2(n8316), .A(n14277), .ZN(n14279) );
  NAND2_X1 U16015 ( .A1(n14280), .A2(n14279), .ZN(n14281) );
  OAI211_X1 U16016 ( .C1(n14284), .C2(n14283), .A(n14282), .B(n14281), .ZN(
        n14285) );
  INV_X1 U16017 ( .A(n14285), .ZN(n14287) );
  OAI211_X1 U16018 ( .C1(n14289), .C2(n14288), .A(n14287), .B(n14286), .ZN(
        P1_U3261) );
  XNOR2_X1 U16019 ( .A(n14290), .B(n14291), .ZN(n14391) );
  XNOR2_X1 U16020 ( .A(n14292), .B(n14291), .ZN(n14294) );
  OAI21_X1 U16021 ( .B1(n14294), .B2(n14379), .A(n14293), .ZN(n14295) );
  AOI21_X1 U16022 ( .B1(n14391), .B2(n14403), .A(n14295), .ZN(n14388) );
  AOI22_X1 U16023 ( .A1(n14315), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n14296), 
        .B2(n14311), .ZN(n14297) );
  OAI21_X1 U16024 ( .B1(n14298), .B2(n14387), .A(n14297), .ZN(n14299) );
  INV_X1 U16025 ( .A(n14299), .ZN(n14306) );
  INV_X1 U16026 ( .A(n14300), .ZN(n14302) );
  OAI211_X1 U16027 ( .C1(n14387), .C2(n14302), .A(n14301), .B(n9843), .ZN(
        n14386) );
  INV_X1 U16028 ( .A(n14386), .ZN(n14303) );
  AOI22_X1 U16029 ( .A1(n14391), .A2(n14304), .B1(n14313), .B2(n14303), .ZN(
        n14305) );
  OAI211_X1 U16030 ( .C1(n14315), .C2(n14388), .A(n14306), .B(n14305), .ZN(
        P1_U3287) );
  NAND2_X1 U16031 ( .A1(n14308), .A2(n14307), .ZN(n14319) );
  NAND2_X1 U16032 ( .A1(n14310), .A2(n14309), .ZN(n14318) );
  AOI22_X1 U16033 ( .A1(n14313), .A2(n14312), .B1(n14311), .B2(n8025), .ZN(
        n14317) );
  NAND2_X1 U16034 ( .A1(n14315), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n14316) );
  AND4_X1 U16035 ( .A1(n14319), .A2(n14318), .A3(n14317), .A4(n14316), .ZN(
        n14320) );
  OAI21_X1 U16036 ( .B1(n14322), .B2(n14321), .A(n14320), .ZN(P1_U3290) );
  INV_X1 U16037 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14323) );
  NOR2_X1 U16038 ( .A1(n14350), .A2(n14323), .ZN(P1_U3294) );
  INV_X1 U16039 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14903) );
  NOR2_X1 U16040 ( .A1(n14350), .A2(n14903), .ZN(P1_U3295) );
  INV_X1 U16041 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14324) );
  NOR2_X1 U16042 ( .A1(n14350), .A2(n14324), .ZN(P1_U3296) );
  INV_X1 U16043 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14325) );
  NOR2_X1 U16044 ( .A1(n14350), .A2(n14325), .ZN(P1_U3297) );
  INV_X1 U16045 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14326) );
  NOR2_X1 U16046 ( .A1(n14350), .A2(n14326), .ZN(P1_U3298) );
  INV_X1 U16047 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14327) );
  NOR2_X1 U16048 ( .A1(n14350), .A2(n14327), .ZN(P1_U3299) );
  INV_X1 U16049 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14328) );
  NOR2_X1 U16050 ( .A1(n14350), .A2(n14328), .ZN(P1_U3300) );
  INV_X1 U16051 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14329) );
  NOR2_X1 U16052 ( .A1(n14350), .A2(n14329), .ZN(P1_U3301) );
  INV_X1 U16053 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14330) );
  NOR2_X1 U16054 ( .A1(n14350), .A2(n14330), .ZN(P1_U3302) );
  INV_X1 U16055 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14991) );
  NOR2_X1 U16056 ( .A1(n14350), .A2(n14991), .ZN(P1_U3303) );
  INV_X1 U16057 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14331) );
  NOR2_X1 U16058 ( .A1(n14350), .A2(n14331), .ZN(P1_U3304) );
  INV_X1 U16059 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14332) );
  NOR2_X1 U16060 ( .A1(n14350), .A2(n14332), .ZN(P1_U3305) );
  INV_X1 U16061 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14333) );
  NOR2_X1 U16062 ( .A1(n14350), .A2(n14333), .ZN(P1_U3306) );
  INV_X1 U16063 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14334) );
  NOR2_X1 U16064 ( .A1(n14350), .A2(n14334), .ZN(P1_U3307) );
  INV_X1 U16065 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14335) );
  NOR2_X1 U16066 ( .A1(n14350), .A2(n14335), .ZN(P1_U3308) );
  INV_X1 U16067 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14336) );
  NOR2_X1 U16068 ( .A1(n14350), .A2(n14336), .ZN(P1_U3309) );
  INV_X1 U16069 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14337) );
  NOR2_X1 U16070 ( .A1(n14350), .A2(n14337), .ZN(P1_U3310) );
  INV_X1 U16071 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14338) );
  NOR2_X1 U16072 ( .A1(n14350), .A2(n14338), .ZN(P1_U3311) );
  INV_X1 U16073 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14339) );
  NOR2_X1 U16074 ( .A1(n14350), .A2(n14339), .ZN(P1_U3312) );
  INV_X1 U16075 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14340) );
  NOR2_X1 U16076 ( .A1(n14350), .A2(n14340), .ZN(P1_U3313) );
  INV_X1 U16077 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14341) );
  NOR2_X1 U16078 ( .A1(n14350), .A2(n14341), .ZN(P1_U3314) );
  INV_X1 U16079 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14941) );
  NOR2_X1 U16080 ( .A1(n14350), .A2(n14941), .ZN(P1_U3315) );
  INV_X1 U16081 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14342) );
  NOR2_X1 U16082 ( .A1(n14350), .A2(n14342), .ZN(P1_U3316) );
  INV_X1 U16083 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14343) );
  NOR2_X1 U16084 ( .A1(n14350), .A2(n14343), .ZN(P1_U3317) );
  INV_X1 U16085 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14344) );
  NOR2_X1 U16086 ( .A1(n14350), .A2(n14344), .ZN(P1_U3318) );
  INV_X1 U16087 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14345) );
  NOR2_X1 U16088 ( .A1(n14350), .A2(n14345), .ZN(P1_U3319) );
  INV_X1 U16089 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14346) );
  NOR2_X1 U16090 ( .A1(n14350), .A2(n14346), .ZN(P1_U3320) );
  INV_X1 U16091 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14347) );
  NOR2_X1 U16092 ( .A1(n14350), .A2(n14347), .ZN(P1_U3321) );
  INV_X1 U16093 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14348) );
  NOR2_X1 U16094 ( .A1(n14350), .A2(n14348), .ZN(P1_U3322) );
  INV_X1 U16095 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14349) );
  NOR2_X1 U16096 ( .A1(n14350), .A2(n14349), .ZN(P1_U3323) );
  OAI22_X1 U16097 ( .A1(n14353), .A2(n14352), .B1(n14351), .B2(n14417), .ZN(
        n14355) );
  AOI211_X1 U16098 ( .C1(n14392), .C2(n14356), .A(n14355), .B(n14354), .ZN(
        n14426) );
  INV_X1 U16099 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n14357) );
  AOI22_X1 U16100 ( .A1(n14425), .A2(n14426), .B1(n14357), .B2(n14423), .ZN(
        P1_U3462) );
  INV_X1 U16101 ( .A(n14358), .ZN(n14359) );
  OAI21_X1 U16102 ( .B1(n6815), .B2(n14417), .A(n14359), .ZN(n14361) );
  AOI211_X1 U16103 ( .C1(n14392), .C2(n14362), .A(n14361), .B(n14360), .ZN(
        n14428) );
  INV_X1 U16104 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n14363) );
  AOI22_X1 U16105 ( .A1(n14425), .A2(n14428), .B1(n14363), .B2(n14423), .ZN(
        P1_U3465) );
  INV_X1 U16106 ( .A(n14364), .ZN(n14366) );
  OAI211_X1 U16107 ( .C1(n14367), .C2(n14417), .A(n14366), .B(n14365), .ZN(
        n14371) );
  NOR2_X1 U16108 ( .A1(n14369), .A2(n14368), .ZN(n14370) );
  AOI211_X1 U16109 ( .C1(n14373), .C2(n14372), .A(n14371), .B(n14370), .ZN(
        n14430) );
  INV_X1 U16110 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14374) );
  AOI22_X1 U16111 ( .A1(n14425), .A2(n14430), .B1(n14374), .B2(n14423), .ZN(
        P1_U3471) );
  AOI21_X1 U16112 ( .B1(n14397), .B2(n14376), .A(n14375), .ZN(n14378) );
  OAI211_X1 U16113 ( .C1(n14380), .C2(n14379), .A(n14378), .B(n14377), .ZN(
        n14383) );
  NOR2_X1 U16114 ( .A1(n14381), .A2(n14400), .ZN(n14382) );
  AOI211_X1 U16115 ( .C1(n14384), .C2(n14403), .A(n14383), .B(n14382), .ZN(
        n14432) );
  INV_X1 U16116 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14385) );
  AOI22_X1 U16117 ( .A1(n14425), .A2(n14432), .B1(n14385), .B2(n14423), .ZN(
        P1_U3474) );
  OAI21_X1 U16118 ( .B1(n14387), .B2(n14417), .A(n14386), .ZN(n14390) );
  INV_X1 U16119 ( .A(n14388), .ZN(n14389) );
  AOI211_X1 U16120 ( .C1(n14392), .C2(n14391), .A(n14390), .B(n14389), .ZN(
        n14433) );
  INV_X1 U16121 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n14393) );
  AOI22_X1 U16122 ( .A1(n14425), .A2(n14433), .B1(n14393), .B2(n14423), .ZN(
        P1_U3477) );
  INV_X1 U16123 ( .A(n14399), .ZN(n14402) );
  AOI211_X1 U16124 ( .C1(n14397), .C2(n14396), .A(n14395), .B(n14394), .ZN(
        n14398) );
  OAI21_X1 U16125 ( .B1(n14400), .B2(n14399), .A(n14398), .ZN(n14401) );
  AOI21_X1 U16126 ( .B1(n14403), .B2(n14402), .A(n14401), .ZN(n14434) );
  INV_X1 U16127 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14404) );
  AOI22_X1 U16128 ( .A1(n14425), .A2(n14434), .B1(n14404), .B2(n14423), .ZN(
        P1_U3480) );
  OAI211_X1 U16129 ( .C1(n6822), .C2(n14417), .A(n14406), .B(n14405), .ZN(
        n14407) );
  AOI21_X1 U16130 ( .B1(n14408), .B2(n14421), .A(n14407), .ZN(n14436) );
  INV_X1 U16131 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14409) );
  AOI22_X1 U16132 ( .A1(n14425), .A2(n14436), .B1(n14409), .B2(n14423), .ZN(
        P1_U3483) );
  OAI211_X1 U16133 ( .C1(n14412), .C2(n14417), .A(n14411), .B(n14410), .ZN(
        n14413) );
  AOI21_X1 U16134 ( .B1(n14414), .B2(n14421), .A(n14413), .ZN(n14437) );
  INV_X1 U16135 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14966) );
  AOI22_X1 U16136 ( .A1(n14425), .A2(n14437), .B1(n14966), .B2(n14423), .ZN(
        P1_U3486) );
  OAI211_X1 U16137 ( .C1(n14418), .C2(n14417), .A(n14416), .B(n14415), .ZN(
        n14420) );
  AOI211_X1 U16138 ( .C1(n14422), .C2(n14421), .A(n14420), .B(n14419), .ZN(
        n14440) );
  INV_X1 U16139 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14424) );
  AOI22_X1 U16140 ( .A1(n14425), .A2(n14440), .B1(n14424), .B2(n14423), .ZN(
        P1_U3489) );
  AOI22_X1 U16141 ( .A1(n14441), .A2(n14426), .B1(n9410), .B2(n14438), .ZN(
        P1_U3529) );
  AOI22_X1 U16142 ( .A1(n14441), .A2(n14428), .B1(n14427), .B2(n14438), .ZN(
        P1_U3530) );
  AOI22_X1 U16143 ( .A1(n14441), .A2(n14430), .B1(n14429), .B2(n14438), .ZN(
        P1_U3532) );
  INV_X1 U16144 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14431) );
  AOI22_X1 U16145 ( .A1(n14441), .A2(n14432), .B1(n14431), .B2(n14438), .ZN(
        P1_U3533) );
  AOI22_X1 U16146 ( .A1(n14441), .A2(n14433), .B1(n9416), .B2(n14438), .ZN(
        P1_U3534) );
  AOI22_X1 U16147 ( .A1(n14441), .A2(n14434), .B1(n9418), .B2(n14438), .ZN(
        P1_U3535) );
  AOI22_X1 U16148 ( .A1(n14441), .A2(n14436), .B1(n14435), .B2(n14438), .ZN(
        P1_U3536) );
  AOI22_X1 U16149 ( .A1(n14441), .A2(n14437), .B1(n9459), .B2(n14438), .ZN(
        P1_U3537) );
  AOI22_X1 U16150 ( .A1(n14441), .A2(n14440), .B1(n14439), .B2(n14438), .ZN(
        P1_U3538) );
  NOR2_X1 U16151 ( .A1(n14442), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI211_X1 U16152 ( .C1(n14445), .C2(n14444), .A(n14443), .B(n14527), .ZN(
        n14450) );
  AOI211_X1 U16153 ( .C1(n14448), .C2(n14447), .A(n14446), .B(n14531), .ZN(
        n14449) );
  AOI211_X1 U16154 ( .C1(n14537), .C2(n14451), .A(n14450), .B(n14449), .ZN(
        n14453) );
  NAND2_X1 U16155 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n14452) );
  OAI211_X1 U16156 ( .C1(n14540), .C2(n14454), .A(n14453), .B(n14452), .ZN(
        P2_U3217) );
  INV_X1 U16157 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15027) );
  AOI211_X1 U16158 ( .C1(n14457), .C2(n14456), .A(n14527), .B(n14455), .ZN(
        n14462) );
  AOI211_X1 U16159 ( .C1(n14460), .C2(n14459), .A(n14531), .B(n14458), .ZN(
        n14461) );
  AOI211_X1 U16160 ( .C1(n14537), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n14465) );
  OAI211_X1 U16161 ( .C1(n14540), .C2(n15027), .A(n14465), .B(n14464), .ZN(
        P2_U3219) );
  AOI211_X1 U16162 ( .C1(n14468), .C2(n14467), .A(n14527), .B(n14466), .ZN(
        n14473) );
  AOI211_X1 U16163 ( .C1(n14471), .C2(n14470), .A(n14531), .B(n14469), .ZN(
        n14472) );
  AOI211_X1 U16164 ( .C1(n14537), .C2(n14474), .A(n14473), .B(n14472), .ZN(
        n14476) );
  OAI211_X1 U16165 ( .C1(n14477), .C2(n14540), .A(n14476), .B(n14475), .ZN(
        P2_U3222) );
  AOI211_X1 U16166 ( .C1(n14480), .C2(n14479), .A(n14527), .B(n14478), .ZN(
        n14485) );
  AOI211_X1 U16167 ( .C1(n14483), .C2(n14482), .A(n14531), .B(n14481), .ZN(
        n14484) );
  AOI211_X1 U16168 ( .C1(n14537), .C2(n14486), .A(n14485), .B(n14484), .ZN(
        n14488) );
  OAI211_X1 U16169 ( .C1(n14489), .C2(n14540), .A(n14488), .B(n14487), .ZN(
        P2_U3224) );
  AOI211_X1 U16170 ( .C1(n14491), .C2(n11014), .A(n14490), .B(n14527), .ZN(
        n14496) );
  AOI211_X1 U16171 ( .C1(n14494), .C2(n14493), .A(n14492), .B(n14531), .ZN(
        n14495) );
  AOI211_X1 U16172 ( .C1(n14537), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14499) );
  OAI211_X1 U16173 ( .C1(n14500), .C2(n14540), .A(n14499), .B(n14498), .ZN(
        P2_U3228) );
  INV_X1 U16174 ( .A(n14501), .ZN(n14510) );
  AOI211_X1 U16175 ( .C1(n14504), .C2(n14503), .A(n14502), .B(n14531), .ZN(
        n14509) );
  AOI211_X1 U16176 ( .C1(n14507), .C2(n14506), .A(n14505), .B(n14527), .ZN(
        n14508) );
  AOI211_X1 U16177 ( .C1(n14537), .C2(n14510), .A(n14509), .B(n14508), .ZN(
        n14512) );
  NAND2_X1 U16178 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n14511)
         );
  OAI211_X1 U16179 ( .C1(n14513), .C2(n14540), .A(n14512), .B(n14511), .ZN(
        P2_U3229) );
  AOI211_X1 U16180 ( .C1(n14516), .C2(n14515), .A(n14514), .B(n14531), .ZN(
        n14521) );
  AOI211_X1 U16181 ( .C1(n14519), .C2(n14518), .A(n14517), .B(n14527), .ZN(
        n14520) );
  AOI211_X1 U16182 ( .C1(n14537), .C2(n14522), .A(n14521), .B(n14520), .ZN(
        n14524) );
  OAI211_X1 U16183 ( .C1(n14525), .C2(n14540), .A(n14524), .B(n14523), .ZN(
        P2_U3230) );
  AOI211_X1 U16184 ( .C1(n14529), .C2(n14528), .A(n14527), .B(n14526), .ZN(
        n14535) );
  AOI211_X1 U16185 ( .C1(n14533), .C2(n14532), .A(n14531), .B(n14530), .ZN(
        n14534) );
  AOI211_X1 U16186 ( .C1(n14537), .C2(n14536), .A(n14535), .B(n14534), .ZN(
        n14539) );
  OAI211_X1 U16187 ( .C1(n14541), .C2(n14540), .A(n14539), .B(n14538), .ZN(
        P2_U3231) );
  INV_X1 U16188 ( .A(n14542), .ZN(n14547) );
  INV_X1 U16189 ( .A(n14543), .ZN(n14544) );
  NAND2_X1 U16190 ( .A1(n14545), .A2(n14544), .ZN(n14568) );
  OAI22_X1 U16191 ( .A1(n14567), .A2(n14547), .B1(n14546), .B2(n14568), .ZN(
        n14552) );
  NOR2_X1 U16192 ( .A1(n14549), .A2(n14548), .ZN(n14551) );
  OAI21_X1 U16193 ( .B1(n14551), .B2(n14567), .A(n14550), .ZN(n14569) );
  AOI211_X1 U16194 ( .C1(n14553), .C2(P2_REG3_REG_0__SCAN_IN), .A(n14552), .B(
        n14569), .ZN(n14555) );
  AOI22_X1 U16195 ( .A1(n14557), .A2(n14556), .B1(n14555), .B2(n14554), .ZN(
        P2_U3265) );
  INV_X1 U16196 ( .A(n14566), .ZN(n14563) );
  AND2_X1 U16197 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14560), .ZN(P2_U3266) );
  AND2_X1 U16198 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14560), .ZN(P2_U3267) );
  AND2_X1 U16199 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14560), .ZN(P2_U3268) );
  AND2_X1 U16200 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14560), .ZN(P2_U3269) );
  AND2_X1 U16201 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14560), .ZN(P2_U3270) );
  AND2_X1 U16202 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14560), .ZN(P2_U3271) );
  AND2_X1 U16203 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14560), .ZN(P2_U3272) );
  AND2_X1 U16204 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14560), .ZN(P2_U3273) );
  AND2_X1 U16205 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14560), .ZN(P2_U3274) );
  AND2_X1 U16206 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14560), .ZN(P2_U3275) );
  AND2_X1 U16207 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14560), .ZN(P2_U3276) );
  AND2_X1 U16208 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14560), .ZN(P2_U3277) );
  AND2_X1 U16209 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14560), .ZN(P2_U3278) );
  AND2_X1 U16210 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14560), .ZN(P2_U3279) );
  AND2_X1 U16211 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14560), .ZN(P2_U3280) );
  INV_X1 U16212 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n14977) );
  NOR2_X1 U16213 ( .A1(n14559), .A2(n14977), .ZN(P2_U3281) );
  AND2_X1 U16214 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14560), .ZN(P2_U3282) );
  AND2_X1 U16215 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14560), .ZN(P2_U3283) );
  AND2_X1 U16216 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14560), .ZN(P2_U3284) );
  AND2_X1 U16217 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14560), .ZN(P2_U3285) );
  INV_X1 U16218 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n14972) );
  NOR2_X1 U16219 ( .A1(n14559), .A2(n14972), .ZN(P2_U3286) );
  INV_X1 U16220 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n14933) );
  NOR2_X1 U16221 ( .A1(n14559), .A2(n14933), .ZN(P2_U3287) );
  AND2_X1 U16222 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14560), .ZN(P2_U3288) );
  AND2_X1 U16223 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14560), .ZN(P2_U3289) );
  AND2_X1 U16224 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14560), .ZN(P2_U3290) );
  AND2_X1 U16225 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14560), .ZN(P2_U3291) );
  AND2_X1 U16226 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14560), .ZN(P2_U3292) );
  AND2_X1 U16227 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14560), .ZN(P2_U3293) );
  AND2_X1 U16228 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14560), .ZN(P2_U3294) );
  AND2_X1 U16229 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14560), .ZN(P2_U3295) );
  AOI22_X1 U16230 ( .A1(n14566), .A2(n14562), .B1(n14561), .B2(n14563), .ZN(
        P2_U3416) );
  AOI22_X1 U16231 ( .A1(n14566), .A2(n14565), .B1(n14564), .B2(n14563), .ZN(
        P2_U3417) );
  INV_X1 U16232 ( .A(n14567), .ZN(n14571) );
  INV_X1 U16233 ( .A(n14568), .ZN(n14570) );
  AOI211_X1 U16234 ( .C1(n14571), .C2(n14630), .A(n14570), .B(n14569), .ZN(
        n14650) );
  INV_X1 U16235 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14962) );
  AOI22_X1 U16236 ( .A1(n14648), .A2(n14650), .B1(n14962), .B2(n14646), .ZN(
        P2_U3430) );
  OAI21_X1 U16237 ( .B1(n10046), .B2(n14627), .A(n14572), .ZN(n14574) );
  AOI211_X1 U16238 ( .C1(n14614), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14652) );
  INV_X1 U16239 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14576) );
  AOI22_X1 U16240 ( .A1(n14648), .A2(n14652), .B1(n14576), .B2(n14646), .ZN(
        P2_U3436) );
  AOI211_X1 U16241 ( .C1(n14637), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        n14581) );
  OAI211_X1 U16242 ( .C1(n14583), .C2(n14582), .A(n14581), .B(n14580), .ZN(
        n14584) );
  INV_X1 U16243 ( .A(n14584), .ZN(n14653) );
  INV_X1 U16244 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U16245 ( .A1(n14648), .A2(n14653), .B1(n14585), .B2(n14646), .ZN(
        P2_U3439) );
  INV_X1 U16246 ( .A(n14586), .ZN(n14591) );
  OAI21_X1 U16247 ( .B1(n14588), .B2(n14627), .A(n14587), .ZN(n14590) );
  AOI211_X1 U16248 ( .C1(n14630), .C2(n14591), .A(n14590), .B(n14589), .ZN(
        n14655) );
  INV_X1 U16249 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16250 ( .A1(n14648), .A2(n14655), .B1(n14592), .B2(n14646), .ZN(
        P2_U3442) );
  INV_X1 U16251 ( .A(n14593), .ZN(n14598) );
  OAI21_X1 U16252 ( .B1(n14595), .B2(n14627), .A(n14594), .ZN(n14597) );
  AOI211_X1 U16253 ( .C1(n14630), .C2(n14598), .A(n14597), .B(n14596), .ZN(
        n14656) );
  INV_X1 U16254 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14599) );
  AOI22_X1 U16255 ( .A1(n14648), .A2(n14656), .B1(n14599), .B2(n14646), .ZN(
        P2_U3445) );
  NOR2_X1 U16256 ( .A1(n14600), .A2(n9575), .ZN(n14606) );
  INV_X1 U16257 ( .A(n14601), .ZN(n14604) );
  OAI211_X1 U16258 ( .C1(n14604), .C2(n14627), .A(n14603), .B(n14602), .ZN(
        n14605) );
  AOI211_X1 U16259 ( .C1(n14607), .C2(n14630), .A(n14606), .B(n14605), .ZN(
        n14657) );
  INV_X1 U16260 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14608) );
  AOI22_X1 U16261 ( .A1(n14648), .A2(n14657), .B1(n14608), .B2(n14646), .ZN(
        P2_U3448) );
  OAI21_X1 U16262 ( .B1(n14610), .B2(n14627), .A(n14609), .ZN(n14613) );
  INV_X1 U16263 ( .A(n14611), .ZN(n14612) );
  AOI211_X1 U16264 ( .C1(n14615), .C2(n14614), .A(n14613), .B(n14612), .ZN(
        n14658) );
  INV_X1 U16265 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14616) );
  AOI22_X1 U16266 ( .A1(n14648), .A2(n14658), .B1(n14616), .B2(n14646), .ZN(
        P2_U3451) );
  NOR2_X1 U16267 ( .A1(n14620), .A2(n9575), .ZN(n14622) );
  NAND2_X1 U16268 ( .A1(n14617), .A2(n14637), .ZN(n14619) );
  OAI211_X1 U16269 ( .C1(n14620), .C2(n14641), .A(n14619), .B(n14618), .ZN(
        n14621) );
  NOR3_X1 U16270 ( .A1(n14623), .A2(n14622), .A3(n14621), .ZN(n14659) );
  INV_X1 U16271 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14624) );
  AOI22_X1 U16272 ( .A1(n14648), .A2(n14659), .B1(n14624), .B2(n14646), .ZN(
        P2_U3454) );
  INV_X1 U16273 ( .A(n14632), .ZN(n14631) );
  INV_X1 U16274 ( .A(n14625), .ZN(n14626) );
  OAI21_X1 U16275 ( .B1(n14628), .B2(n14627), .A(n14626), .ZN(n14629) );
  AOI21_X1 U16276 ( .B1(n14631), .B2(n14630), .A(n14629), .ZN(n14634) );
  OR2_X1 U16277 ( .A1(n14632), .A2(n9575), .ZN(n14633) );
  INV_X1 U16278 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14636) );
  AOI22_X1 U16279 ( .A1(n14648), .A2(n14660), .B1(n14636), .B2(n14646), .ZN(
        P2_U3457) );
  NOR2_X1 U16280 ( .A1(n14642), .A2(n9575), .ZN(n14644) );
  NAND2_X1 U16281 ( .A1(n14638), .A2(n14637), .ZN(n14640) );
  OAI211_X1 U16282 ( .C1(n14642), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14643) );
  NOR3_X1 U16283 ( .A1(n14645), .A2(n14644), .A3(n14643), .ZN(n14662) );
  INV_X1 U16284 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14647) );
  AOI22_X1 U16285 ( .A1(n14648), .A2(n14662), .B1(n14647), .B2(n14646), .ZN(
        P2_U3460) );
  AOI22_X1 U16286 ( .A1(n14663), .A2(n14650), .B1(n14649), .B2(n14661), .ZN(
        P2_U3499) );
  INV_X1 U16287 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n14651) );
  AOI22_X1 U16288 ( .A1(n14663), .A2(n14652), .B1(n14651), .B2(n14661), .ZN(
        P2_U3501) );
  INV_X1 U16289 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n14973) );
  AOI22_X1 U16290 ( .A1(n14663), .A2(n14653), .B1(n14973), .B2(n14661), .ZN(
        P2_U3502) );
  INV_X1 U16291 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14654) );
  AOI22_X1 U16292 ( .A1(n14663), .A2(n14655), .B1(n14654), .B2(n14661), .ZN(
        P2_U3503) );
  INV_X1 U16293 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14990) );
  AOI22_X1 U16294 ( .A1(n14663), .A2(n14656), .B1(n14990), .B2(n14661), .ZN(
        P2_U3504) );
  AOI22_X1 U16295 ( .A1(n14663), .A2(n14657), .B1(n9489), .B2(n14661), .ZN(
        P2_U3505) );
  AOI22_X1 U16296 ( .A1(n14663), .A2(n14658), .B1(n9682), .B2(n14661), .ZN(
        P2_U3506) );
  AOI22_X1 U16297 ( .A1(n14663), .A2(n14659), .B1(n10003), .B2(n14661), .ZN(
        P2_U3507) );
  AOI22_X1 U16298 ( .A1(n14663), .A2(n14660), .B1(n10004), .B2(n14661), .ZN(
        P2_U3508) );
  AOI22_X1 U16299 ( .A1(n14663), .A2(n14662), .B1(n10529), .B2(n14661), .ZN(
        P2_U3509) );
  NOR2_X1 U16300 ( .A1(P3_U3897), .A2(n14664), .ZN(P3_U3150) );
  OAI21_X1 U16301 ( .B1(n14667), .B2(n14666), .A(n14665), .ZN(n14674) );
  OAI211_X1 U16302 ( .C1(n14671), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14672) );
  INV_X1 U16303 ( .A(n14672), .ZN(n14673) );
  AOI211_X1 U16304 ( .C1(n14676), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14677) );
  OAI21_X1 U16305 ( .B1(n14679), .B2(n14678), .A(n14677), .ZN(P3_U3153) );
  AOI21_X1 U16306 ( .B1(n14681), .B2(n14976), .A(n14680), .ZN(n14694) );
  OAI21_X1 U16307 ( .B1(n14683), .B2(P3_REG1_REG_9__SCAN_IN), .A(n14682), .ZN(
        n14684) );
  AOI22_X1 U16308 ( .A1(n14686), .A2(n14685), .B1(n14703), .B2(n14684), .ZN(
        n14693) );
  INV_X1 U16309 ( .A(n14711), .ZN(n14690) );
  AND2_X1 U16310 ( .A1(n14711), .A2(n14687), .ZN(n14689) );
  OAI22_X1 U16311 ( .A1(n14712), .A2(n14690), .B1(n14689), .B2(n14688), .ZN(
        n14691) );
  NAND2_X1 U16312 ( .A1(n14691), .A2(n14713), .ZN(n14692) );
  OAI211_X1 U16313 ( .C1(n14694), .C2(n14708), .A(n14693), .B(n14692), .ZN(
        n14695) );
  INV_X1 U16314 ( .A(n14695), .ZN(n14697) );
  NAND2_X1 U16315 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(P3_U3151), .ZN(n14696) );
  OAI211_X1 U16316 ( .C1(n14698), .C2(n14724), .A(n14697), .B(n14696), .ZN(
        P3_U3191) );
  OAI21_X1 U16317 ( .B1(n14701), .B2(n14700), .A(n14699), .ZN(n14704) );
  AOI21_X1 U16318 ( .B1(n14704), .B2(n14703), .A(n14702), .ZN(n14722) );
  AOI21_X1 U16319 ( .B1(n14707), .B2(n14706), .A(n14705), .ZN(n14709) );
  OR2_X1 U16320 ( .A1(n14709), .A2(n14708), .ZN(n14717) );
  AND3_X1 U16321 ( .A1(n14712), .A2(n14711), .A3(n14710), .ZN(n14714) );
  OAI21_X1 U16322 ( .B1(n14715), .B2(n14714), .A(n14713), .ZN(n14716) );
  OAI211_X1 U16323 ( .C1(n14719), .C2(n14718), .A(n14717), .B(n14716), .ZN(
        n14720) );
  INV_X1 U16324 ( .A(n14720), .ZN(n14721) );
  OAI211_X1 U16325 ( .C1(n14724), .C2(n14723), .A(n14722), .B(n14721), .ZN(
        P3_U3192) );
  AND2_X1 U16326 ( .A1(n14725), .A2(n14821), .ZN(n14846) );
  AOI22_X1 U16327 ( .A1(n14726), .A2(n14846), .B1(n14793), .B2(
        P3_REG2_REG_10__SCAN_IN), .ZN(n14740) );
  OAI211_X1 U16328 ( .C1(n14728), .C2(n14735), .A(n14727), .B(n14778), .ZN(
        n14734) );
  AOI22_X1 U16329 ( .A1(n14732), .A2(n14731), .B1(n14730), .B2(n14729), .ZN(
        n14733) );
  NAND2_X1 U16330 ( .A1(n14734), .A2(n14733), .ZN(n14845) );
  XNOR2_X1 U16331 ( .A(n14736), .B(n14735), .ZN(n14847) );
  AND2_X1 U16332 ( .A1(n14847), .A2(n14737), .ZN(n14738) );
  AOI21_X1 U16333 ( .B1(n14791), .B2(n14845), .A(n14738), .ZN(n14739) );
  OAI211_X1 U16334 ( .C1(n14741), .C2(n14785), .A(n14740), .B(n14739), .ZN(
        P3_U3223) );
  OR2_X1 U16335 ( .A1(n14743), .A2(n14742), .ZN(n14744) );
  NAND2_X1 U16336 ( .A1(n14745), .A2(n14744), .ZN(n14822) );
  INV_X1 U16337 ( .A(n14822), .ZN(n14752) );
  OAI211_X1 U16338 ( .C1(n14746), .C2(n14748), .A(n14747), .B(n14778), .ZN(
        n14749) );
  INV_X1 U16339 ( .A(n14749), .ZN(n14750) );
  AOI211_X1 U16340 ( .C1(n14843), .C2(n14822), .A(n14751), .B(n14750), .ZN(
        n14824) );
  OAI21_X1 U16341 ( .B1(n14752), .B2(n14770), .A(n14824), .ZN(n14753) );
  MUX2_X1 U16342 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n14753), .S(n14791), .Z(
        n14754) );
  AOI21_X1 U16343 ( .B1(n6433), .B2(n14820), .A(n14754), .ZN(n14755) );
  OAI21_X1 U16344 ( .B1(n14756), .B2(n14785), .A(n14755), .ZN(P3_U3227) );
  XNOR2_X1 U16345 ( .A(n14757), .B(n14759), .ZN(n14800) );
  XNOR2_X1 U16346 ( .A(n14758), .B(n14759), .ZN(n14765) );
  OAI22_X1 U16347 ( .A1(n14763), .A2(n14762), .B1(n14761), .B2(n14760), .ZN(
        n14764) );
  AOI21_X1 U16348 ( .B1(n14765), .B2(n14778), .A(n14764), .ZN(n14766) );
  OAI21_X1 U16349 ( .B1(n14800), .B2(n14783), .A(n14766), .ZN(n14801) );
  NOR2_X1 U16350 ( .A1(n14767), .A2(n14837), .ZN(n14802) );
  INV_X1 U16351 ( .A(n14802), .ZN(n14768) );
  OAI22_X1 U16352 ( .A1(n14800), .A2(n14770), .B1(n14769), .B2(n14768), .ZN(
        n14771) );
  AOI211_X1 U16353 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n14772), .A(n14801), .B(
        n14771), .ZN(n14773) );
  AOI22_X1 U16354 ( .A1(n14793), .A2(n14774), .B1(n14773), .B2(n14791), .ZN(
        P3_U3231) );
  XNOR2_X1 U16355 ( .A(n9945), .B(n14775), .ZN(n14794) );
  XNOR2_X1 U16356 ( .A(n14776), .B(n9945), .ZN(n14779) );
  AOI21_X1 U16357 ( .B1(n14779), .B2(n14778), .A(n14777), .ZN(n14795) );
  NAND3_X1 U16358 ( .A1(n14781), .A2(n14821), .A3(n14780), .ZN(n14782) );
  OAI211_X1 U16359 ( .C1(n14783), .C2(n14794), .A(n14795), .B(n14782), .ZN(
        n14784) );
  INV_X1 U16360 ( .A(n14784), .ZN(n14792) );
  OAI22_X1 U16361 ( .A1(n14787), .A2(n14794), .B1(n14786), .B2(n14785), .ZN(
        n14788) );
  INV_X1 U16362 ( .A(n14788), .ZN(n14789) );
  OAI221_X1 U16363 ( .B1(n14793), .B2(n14792), .C1(n14791), .C2(n14790), .A(
        n14789), .ZN(P3_U3232) );
  INV_X1 U16364 ( .A(n14794), .ZN(n14798) );
  OAI21_X1 U16365 ( .B1(n14796), .B2(n14837), .A(n14795), .ZN(n14797) );
  AOI21_X1 U16366 ( .B1(n14848), .B2(n14798), .A(n14797), .ZN(n14852) );
  INV_X1 U16367 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U16368 ( .A1(n14851), .A2(n14852), .B1(n14799), .B2(n14849), .ZN(
        P3_U3393) );
  INV_X1 U16369 ( .A(n14800), .ZN(n14803) );
  AOI211_X1 U16370 ( .C1(n14803), .C2(n14833), .A(n14802), .B(n14801), .ZN(
        n14853) );
  INV_X1 U16371 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n14804) );
  AOI22_X1 U16372 ( .A1(n14851), .A2(n14853), .B1(n14804), .B2(n14849), .ZN(
        P3_U3396) );
  INV_X1 U16373 ( .A(n14805), .ZN(n14806) );
  AOI211_X1 U16374 ( .C1(n14833), .C2(n14808), .A(n14807), .B(n14806), .ZN(
        n14855) );
  INV_X1 U16375 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14809) );
  AOI22_X1 U16376 ( .A1(n14851), .A2(n14855), .B1(n14809), .B2(n14849), .ZN(
        P3_U3399) );
  INV_X1 U16377 ( .A(n14810), .ZN(n14812) );
  AOI211_X1 U16378 ( .C1(n14813), .C2(n14833), .A(n14812), .B(n14811), .ZN(
        n14857) );
  INV_X1 U16379 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n14814) );
  AOI22_X1 U16380 ( .A1(n14851), .A2(n14857), .B1(n14814), .B2(n14849), .ZN(
        P3_U3402) );
  INV_X1 U16381 ( .A(n14815), .ZN(n14817) );
  AOI211_X1 U16382 ( .C1(n14818), .C2(n14833), .A(n14817), .B(n14816), .ZN(
        n14858) );
  INV_X1 U16383 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n14819) );
  AOI22_X1 U16384 ( .A1(n14851), .A2(n14858), .B1(n14819), .B2(n14849), .ZN(
        P3_U3405) );
  AOI22_X1 U16385 ( .A1(n14822), .A2(n14833), .B1(n14821), .B2(n14820), .ZN(
        n14823) );
  AND2_X1 U16386 ( .A1(n14824), .A2(n14823), .ZN(n14860) );
  INV_X1 U16387 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n14825) );
  AOI22_X1 U16388 ( .A1(n14851), .A2(n14860), .B1(n14825), .B2(n14849), .ZN(
        P3_U3408) );
  INV_X1 U16389 ( .A(n14833), .ZN(n14838) );
  OAI22_X1 U16390 ( .A1(n14827), .A2(n14838), .B1(n14837), .B2(n14826), .ZN(
        n14828) );
  NOR2_X1 U16391 ( .A1(n14829), .A2(n14828), .ZN(n14861) );
  INV_X1 U16392 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n14830) );
  AOI22_X1 U16393 ( .A1(n14851), .A2(n14861), .B1(n14830), .B2(n14849), .ZN(
        P3_U3411) );
  AOI211_X1 U16394 ( .C1(n14834), .C2(n14833), .A(n14832), .B(n14831), .ZN(
        n14863) );
  INV_X1 U16395 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n14835) );
  AOI22_X1 U16396 ( .A1(n14851), .A2(n14863), .B1(n14835), .B2(n14849), .ZN(
        P3_U3414) );
  INV_X1 U16397 ( .A(n14839), .ZN(n14842) );
  OAI22_X1 U16398 ( .A1(n14839), .A2(n14838), .B1(n14837), .B2(n14836), .ZN(
        n14841) );
  AOI211_X1 U16399 ( .C1(n14843), .C2(n14842), .A(n14841), .B(n14840), .ZN(
        n14865) );
  INV_X1 U16400 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n14844) );
  AOI22_X1 U16401 ( .A1(n14851), .A2(n14865), .B1(n14844), .B2(n14849), .ZN(
        P3_U3417) );
  AOI211_X1 U16402 ( .C1(n14848), .C2(n14847), .A(n14846), .B(n14845), .ZN(
        n14867) );
  INV_X1 U16403 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n14850) );
  AOI22_X1 U16404 ( .A1(n14851), .A2(n14867), .B1(n14850), .B2(n14849), .ZN(
        P3_U3420) );
  AOI22_X1 U16405 ( .A1(n14868), .A2(n14852), .B1(n9745), .B2(n14866), .ZN(
        P3_U3460) );
  AOI22_X1 U16406 ( .A1(n14868), .A2(n14853), .B1(n7740), .B2(n14866), .ZN(
        P3_U3461) );
  INV_X1 U16407 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n14854) );
  AOI22_X1 U16408 ( .A1(n14868), .A2(n14855), .B1(n14854), .B2(n14866), .ZN(
        P3_U3462) );
  AOI22_X1 U16409 ( .A1(n14868), .A2(n14857), .B1(n14856), .B2(n14866), .ZN(
        P3_U3463) );
  AOI22_X1 U16410 ( .A1(n14868), .A2(n14858), .B1(n7747), .B2(n14866), .ZN(
        P3_U3464) );
  AOI22_X1 U16411 ( .A1(n14868), .A2(n14860), .B1(n14859), .B2(n14866), .ZN(
        P3_U3465) );
  AOI22_X1 U16412 ( .A1(n14868), .A2(n14861), .B1(n7750), .B2(n14866), .ZN(
        P3_U3466) );
  AOI22_X1 U16413 ( .A1(n14868), .A2(n14863), .B1(n14862), .B2(n14866), .ZN(
        P3_U3467) );
  INV_X1 U16414 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n14864) );
  AOI22_X1 U16415 ( .A1(n14868), .A2(n14865), .B1(n14864), .B2(n14866), .ZN(
        P3_U3468) );
  AOI22_X1 U16416 ( .A1(n14868), .A2(n14867), .B1(n14944), .B2(n14866), .ZN(
        P3_U3469) );
  NOR2_X1 U16417 ( .A1(keyinput16), .A2(keyinput24), .ZN(n14869) );
  NAND3_X1 U16418 ( .A1(keyinput58), .A2(keyinput59), .A3(n14869), .ZN(n14873)
         );
  NAND4_X1 U16419 ( .A1(keyinput47), .A2(keyinput38), .A3(keyinput42), .A4(
        keyinput26), .ZN(n14872) );
  NAND4_X1 U16420 ( .A1(keyinput19), .A2(keyinput22), .A3(keyinput14), .A4(
        keyinput33), .ZN(n14871) );
  NAND4_X1 U16421 ( .A1(keyinput32), .A2(keyinput44), .A3(keyinput8), .A4(
        keyinput36), .ZN(n14870) );
  NOR4_X1 U16422 ( .A1(n14873), .A2(n14872), .A3(n14871), .A4(n14870), .ZN(
        n15019) );
  NAND2_X1 U16423 ( .A1(keyinput45), .A2(keyinput13), .ZN(n14874) );
  NOR3_X1 U16424 ( .A1(keyinput54), .A2(keyinput11), .A3(n14874), .ZN(n14880)
         );
  NOR3_X1 U16425 ( .A1(keyinput34), .A2(keyinput57), .A3(keyinput20), .ZN(
        n14879) );
  NAND3_X1 U16426 ( .A1(keyinput43), .A2(keyinput6), .A3(keyinput35), .ZN(
        n14877) );
  INV_X1 U16427 ( .A(keyinput18), .ZN(n14875) );
  NAND3_X1 U16428 ( .A1(keyinput5), .A2(keyinput30), .A3(n14875), .ZN(n14876)
         );
  NOR4_X1 U16429 ( .A1(keyinput56), .A2(keyinput31), .A3(n14877), .A4(n14876), 
        .ZN(n14878) );
  NAND4_X1 U16430 ( .A1(n14880), .A2(keyinput17), .A3(n14879), .A4(n14878), 
        .ZN(n14893) );
  NAND4_X1 U16431 ( .A1(keyinput10), .A2(keyinput0), .A3(keyinput23), .A4(
        keyinput21), .ZN(n14892) );
  NOR2_X1 U16432 ( .A1(keyinput1), .A2(keyinput40), .ZN(n14885) );
  NAND3_X1 U16433 ( .A1(keyinput15), .A2(keyinput12), .A3(keyinput50), .ZN(
        n14883) );
  INV_X1 U16434 ( .A(keyinput62), .ZN(n14881) );
  NAND3_X1 U16435 ( .A1(keyinput53), .A2(keyinput9), .A3(n14881), .ZN(n14882)
         );
  NOR4_X1 U16436 ( .A1(keyinput4), .A2(keyinput52), .A3(n14883), .A4(n14882), 
        .ZN(n14884) );
  NAND4_X1 U16437 ( .A1(keyinput28), .A2(keyinput46), .A3(n14885), .A4(n14884), 
        .ZN(n14891) );
  NOR4_X1 U16438 ( .A1(keyinput63), .A2(keyinput55), .A3(keyinput51), .A4(
        keyinput39), .ZN(n14889) );
  NOR4_X1 U16439 ( .A1(keyinput27), .A2(keyinput7), .A3(keyinput3), .A4(
        keyinput2), .ZN(n14888) );
  NOR4_X1 U16440 ( .A1(keyinput41), .A2(keyinput37), .A3(keyinput61), .A4(
        keyinput49), .ZN(n14887) );
  NOR4_X1 U16441 ( .A1(keyinput25), .A2(keyinput29), .A3(keyinput60), .A4(
        keyinput48), .ZN(n14886) );
  NAND4_X1 U16442 ( .A1(n14889), .A2(n14888), .A3(n14887), .A4(n14886), .ZN(
        n14890) );
  NOR4_X1 U16443 ( .A1(n14893), .A2(n14892), .A3(n14891), .A4(n14890), .ZN(
        n15018) );
  INV_X1 U16444 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14895) );
  AOI22_X1 U16445 ( .A1(n14896), .A2(keyinput45), .B1(keyinput13), .B2(n14895), 
        .ZN(n14894) );
  OAI221_X1 U16446 ( .B1(n14896), .B2(keyinput45), .C1(n14895), .C2(keyinput13), .A(n14894), .ZN(n14908) );
  AOI22_X1 U16447 ( .A1(n14899), .A2(keyinput54), .B1(keyinput11), .B2(n14898), 
        .ZN(n14897) );
  OAI221_X1 U16448 ( .B1(n14899), .B2(keyinput54), .C1(n14898), .C2(keyinput11), .A(n14897), .ZN(n14907) );
  AOI22_X1 U16449 ( .A1(n14901), .A2(keyinput17), .B1(n11572), .B2(keyinput34), 
        .ZN(n14900) );
  OAI221_X1 U16450 ( .B1(n14901), .B2(keyinput17), .C1(n11572), .C2(keyinput34), .A(n14900), .ZN(n14906) );
  AOI22_X1 U16451 ( .A1(n14904), .A2(keyinput57), .B1(keyinput20), .B2(n14903), 
        .ZN(n14902) );
  OAI221_X1 U16452 ( .B1(n14904), .B2(keyinput57), .C1(n14903), .C2(keyinput20), .A(n14902), .ZN(n14905) );
  NOR4_X1 U16453 ( .A1(n14908), .A2(n14907), .A3(n14906), .A4(n14905), .ZN(
        n14954) );
  AOI22_X1 U16454 ( .A1(n14911), .A2(keyinput18), .B1(n14910), .B2(keyinput30), 
        .ZN(n14909) );
  OAI221_X1 U16455 ( .B1(n14911), .B2(keyinput18), .C1(n14910), .C2(keyinput30), .A(n14909), .ZN(n14922) );
  AOI22_X1 U16456 ( .A1(n14913), .A2(keyinput43), .B1(n10645), .B2(keyinput56), 
        .ZN(n14912) );
  OAI221_X1 U16457 ( .B1(n14913), .B2(keyinput43), .C1(n10645), .C2(keyinput56), .A(n14912), .ZN(n14921) );
  INV_X1 U16458 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14915) );
  AOI22_X1 U16459 ( .A1(n14916), .A2(keyinput5), .B1(n14915), .B2(keyinput31), 
        .ZN(n14914) );
  OAI221_X1 U16460 ( .B1(n14916), .B2(keyinput5), .C1(n14915), .C2(keyinput31), 
        .A(n14914), .ZN(n14920) );
  XOR2_X1 U16461 ( .A(n10211), .B(keyinput35), .Z(n14918) );
  XNOR2_X1 U16462 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput6), .ZN(n14917) );
  NAND2_X1 U16463 ( .A1(n14918), .A2(n14917), .ZN(n14919) );
  NOR4_X1 U16464 ( .A1(n14922), .A2(n14921), .A3(n14920), .A4(n14919), .ZN(
        n14953) );
  INV_X1 U16465 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n14925) );
  AOI22_X1 U16466 ( .A1(n14925), .A2(keyinput10), .B1(n14924), .B2(keyinput0), 
        .ZN(n14923) );
  OAI221_X1 U16467 ( .B1(n14925), .B2(keyinput10), .C1(n14924), .C2(keyinput0), 
        .A(n14923), .ZN(n14937) );
  INV_X1 U16468 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n14927) );
  AOI22_X1 U16469 ( .A1(n14928), .A2(keyinput23), .B1(keyinput21), .B2(n14927), 
        .ZN(n14926) );
  OAI221_X1 U16470 ( .B1(n14928), .B2(keyinput23), .C1(n14927), .C2(keyinput21), .A(n14926), .ZN(n14936) );
  AOI22_X1 U16471 ( .A1(n14931), .A2(keyinput28), .B1(keyinput1), .B2(n14930), 
        .ZN(n14929) );
  OAI221_X1 U16472 ( .B1(n14931), .B2(keyinput28), .C1(n14930), .C2(keyinput1), 
        .A(n14929), .ZN(n14935) );
  AOI22_X1 U16473 ( .A1(n9416), .A2(keyinput40), .B1(n14933), .B2(keyinput46), 
        .ZN(n14932) );
  OAI221_X1 U16474 ( .B1(n9416), .B2(keyinput40), .C1(n14933), .C2(keyinput46), 
        .A(n14932), .ZN(n14934) );
  NOR4_X1 U16475 ( .A1(n14937), .A2(n14936), .A3(n14935), .A4(n14934), .ZN(
        n14952) );
  AOI22_X1 U16476 ( .A1(n14939), .A2(keyinput9), .B1(n13458), .B2(keyinput53), 
        .ZN(n14938) );
  OAI221_X1 U16477 ( .B1(n14939), .B2(keyinput9), .C1(n13458), .C2(keyinput53), 
        .A(n14938), .ZN(n14950) );
  AOI22_X1 U16478 ( .A1(n12374), .A2(keyinput12), .B1(keyinput50), .B2(n14941), 
        .ZN(n14940) );
  OAI221_X1 U16479 ( .B1(n12374), .B2(keyinput12), .C1(n14941), .C2(keyinput50), .A(n14940), .ZN(n14949) );
  INV_X1 U16480 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14943) );
  AOI22_X1 U16481 ( .A1(n14944), .A2(keyinput4), .B1(keyinput15), .B2(n14943), 
        .ZN(n14942) );
  OAI221_X1 U16482 ( .B1(n14944), .B2(keyinput4), .C1(n14943), .C2(keyinput15), 
        .A(n14942), .ZN(n14948) );
  XNOR2_X1 U16483 ( .A(P3_IR_REG_0__SCAN_IN), .B(keyinput62), .ZN(n14946) );
  XNOR2_X1 U16484 ( .A(P2_REG2_REG_2__SCAN_IN), .B(keyinput52), .ZN(n14945) );
  NAND2_X1 U16485 ( .A1(n14946), .A2(n14945), .ZN(n14947) );
  NOR4_X1 U16486 ( .A1(n14950), .A2(n14949), .A3(n14948), .A4(n14947), .ZN(
        n14951) );
  NAND4_X1 U16487 ( .A1(n14954), .A2(n14953), .A3(n14952), .A4(n14951), .ZN(
        n15017) );
  AOI22_X1 U16488 ( .A1(n14957), .A2(keyinput60), .B1(n14956), .B2(keyinput22), 
        .ZN(n14955) );
  OAI221_X1 U16489 ( .B1(n14957), .B2(keyinput60), .C1(n14956), .C2(keyinput22), .A(n14955), .ZN(n14970) );
  AOI22_X1 U16490 ( .A1(n14960), .A2(keyinput63), .B1(n14959), .B2(keyinput39), 
        .ZN(n14958) );
  OAI221_X1 U16491 ( .B1(n14960), .B2(keyinput63), .C1(n14959), .C2(keyinput39), .A(n14958), .ZN(n14969) );
  AOI22_X1 U16492 ( .A1(n14963), .A2(keyinput25), .B1(keyinput48), .B2(n14962), 
        .ZN(n14961) );
  OAI221_X1 U16493 ( .B1(n14963), .B2(keyinput25), .C1(n14962), .C2(keyinput48), .A(n14961), .ZN(n14968) );
  AOI22_X1 U16494 ( .A1(n14966), .A2(keyinput51), .B1(keyinput36), .B2(n14965), 
        .ZN(n14964) );
  OAI221_X1 U16495 ( .B1(n14966), .B2(keyinput51), .C1(n14965), .C2(keyinput36), .A(n14964), .ZN(n14967) );
  NOR4_X1 U16496 ( .A1(n14970), .A2(n14969), .A3(n14968), .A4(n14967), .ZN(
        n15015) );
  AOI22_X1 U16497 ( .A1(n14973), .A2(keyinput55), .B1(n14972), .B2(keyinput7), 
        .ZN(n14971) );
  OAI221_X1 U16498 ( .B1(n14973), .B2(keyinput55), .C1(n14972), .C2(keyinput7), 
        .A(n14971), .ZN(n14984) );
  AOI22_X1 U16499 ( .A1(n14976), .A2(keyinput29), .B1(P3_U3151), .B2(
        keyinput16), .ZN(n14974) );
  OAI221_X1 U16500 ( .B1(n14976), .B2(keyinput29), .C1(P3_U3151), .C2(
        keyinput16), .A(n14974), .ZN(n14983) );
  XNOR2_X1 U16501 ( .A(n14977), .B(keyinput32), .ZN(n14982) );
  XNOR2_X1 U16502 ( .A(P2_IR_REG_20__SCAN_IN), .B(keyinput47), .ZN(n14980) );
  XNOR2_X1 U16503 ( .A(P3_REG3_REG_18__SCAN_IN), .B(keyinput38), .ZN(n14979)
         );
  XNOR2_X1 U16504 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput8), .ZN(n14978) );
  NAND3_X1 U16505 ( .A1(n14980), .A2(n14979), .A3(n14978), .ZN(n14981) );
  NOR4_X1 U16506 ( .A1(n14984), .A2(n14983), .A3(n14982), .A4(n14981), .ZN(
        n15014) );
  INV_X1 U16507 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n14987) );
  AOI22_X1 U16508 ( .A1(n14987), .A2(keyinput49), .B1(keyinput42), .B2(n14986), 
        .ZN(n14985) );
  OAI221_X1 U16509 ( .B1(n14987), .B2(keyinput49), .C1(n14986), .C2(keyinput42), .A(n14985), .ZN(n14998) );
  AOI22_X1 U16510 ( .A1(n14990), .A2(keyinput2), .B1(keyinput41), .B2(n14989), 
        .ZN(n14988) );
  OAI221_X1 U16511 ( .B1(n14990), .B2(keyinput2), .C1(n14989), .C2(keyinput41), 
        .A(n14988), .ZN(n14997) );
  XNOR2_X1 U16512 ( .A(n14991), .B(keyinput26), .ZN(n14996) );
  XNOR2_X1 U16513 ( .A(P3_IR_REG_14__SCAN_IN), .B(keyinput3), .ZN(n14994) );
  XNOR2_X1 U16514 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput24), .ZN(n14993) );
  XNOR2_X1 U16515 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput27), .ZN(n14992)
         );
  NAND3_X1 U16516 ( .A1(n14994), .A2(n14993), .A3(n14992), .ZN(n14995) );
  NOR4_X1 U16517 ( .A1(n14998), .A2(n14997), .A3(n14996), .A4(n14995), .ZN(
        n15013) );
  AOI22_X1 U16518 ( .A1(n15000), .A2(keyinput58), .B1(keyinput14), .B2(n9434), 
        .ZN(n14999) );
  OAI221_X1 U16519 ( .B1(n15000), .B2(keyinput58), .C1(n9434), .C2(keyinput14), 
        .A(n14999), .ZN(n15011) );
  INV_X1 U16520 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n15003) );
  INV_X1 U16521 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n15002) );
  AOI22_X1 U16522 ( .A1(n15003), .A2(keyinput61), .B1(keyinput19), .B2(n15002), 
        .ZN(n15001) );
  OAI221_X1 U16523 ( .B1(n15003), .B2(keyinput61), .C1(n15002), .C2(keyinput19), .A(n15001), .ZN(n15010) );
  XNOR2_X1 U16524 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput33), .ZN(n15006)
         );
  XNOR2_X1 U16525 ( .A(P3_IR_REG_9__SCAN_IN), .B(keyinput44), .ZN(n15005) );
  XNOR2_X1 U16526 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput59), .ZN(n15004) );
  NAND3_X1 U16527 ( .A1(n15006), .A2(n15005), .A3(n15004), .ZN(n15009) );
  XNOR2_X1 U16528 ( .A(n15007), .B(keyinput37), .ZN(n15008) );
  NOR4_X1 U16529 ( .A1(n15011), .A2(n15010), .A3(n15009), .A4(n15008), .ZN(
        n15012) );
  NAND4_X1 U16530 ( .A1(n15015), .A2(n15014), .A3(n15013), .A4(n15012), .ZN(
        n15016) );
  AOI211_X1 U16531 ( .C1(n15019), .C2(n15018), .A(n15017), .B(n15016), .ZN(
        n15023) );
  MUX2_X1 U16532 ( .A(n15021), .B(n6922), .S(n15020), .Z(n15022) );
  XNOR2_X1 U16533 ( .A(n15023), .B(n15022), .ZN(P1_U3586) );
  XOR2_X1 U16534 ( .A(n15025), .B(n15024), .Z(SUB_1596_U59) );
  XOR2_X1 U16535 ( .A(n15027), .B(n15026), .Z(SUB_1596_U58) );
  AOI21_X1 U16536 ( .B1(n15029), .B2(n15028), .A(n15037), .ZN(SUB_1596_U53) );
  XOR2_X1 U16537 ( .A(n15030), .B(n15031), .Z(SUB_1596_U56) );
  AOI21_X1 U16538 ( .B1(n15034), .B2(n15033), .A(n15032), .ZN(n15035) );
  XOR2_X1 U16539 ( .A(n15035), .B(P2_ADDR_REG_3__SCAN_IN), .Z(SUB_1596_U60) );
  XOR2_X1 U16540 ( .A(n15037), .B(n15036), .Z(SUB_1596_U5) );
  AND4_X1 U9730 ( .A1(n9020), .A2(n9019), .A3(n9018), .A4(n9936), .ZN(n9825)
         );
  NAND2_X1 U7213 ( .A1(n11026), .A2(n9299), .ZN(n10758) );
  CLKBUF_X1 U7249 ( .A(n9354), .Z(n9864) );
  INV_X2 U7310 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7373) );
endmodule

