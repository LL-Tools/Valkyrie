

module b22_C_2inp_gates_syn ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, SUB_1596_U4, 
        SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, 
        SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, 
        SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, 
        SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53, U29, U28, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, 
        P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, 
        P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556, P1_U3557, 
        P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588, P1_U3589, 
        P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U4016, 
        P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, 
        P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, 
        P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, 
        P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, 
        P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442, P2_U3445, 
        P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463, P2_U3466, 
        P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484, P2_U3486, 
        P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492, P2_U3493, 
        P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, 
        P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, 
        P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, 
        P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, 
        P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527, P2_U3528, 
        P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, 
        P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552, P2_U3553, 
        P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559, P2_U3560, 
        P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211, P2_U3210, 
        P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, 
        P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, 
        P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, 
        P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087, P2_U3947, 
        P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290, P3_U3289, 
        P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283, P3_U3282, 
        P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276, P3_U3275, 
        P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269, P3_U3268, 
        P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377, P3_U3263, 
        P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257, P3_U3256, 
        P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250, P3_U3249, 
        P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243, P3_U3242, 
        P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236, P3_U3235, 
        P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402, P3_U3405, 
        P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423, P3_U3426, 
        P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444, P3_U3446, 
        P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452, P3_U3453, 
        P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459, P3_U3460, 
        P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466, P3_U3467, 
        P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473, P3_U3474, 
        P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480, P3_U3481, 
        P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487, P3_U3488, 
        P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230, P3_U3229, 
        P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223, P3_U3222, 
        P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216, P3_U3215, 
        P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209, P3_U3208, 
        P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202, P3_U3201, 
        P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195, P3_U3194, 
        P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188, P3_U3187, 
        P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491, P3_U3492, 
        P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498, P3_U3499, 
        P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505, P3_U3506, 
        P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512, P3_U3513, 
        P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519, P3_U3520, 
        P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179, P3_U3178, 
        P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172, P3_U3171, 
        P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165, P3_U3164, 
        P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158, P3_U3157, 
        P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150, P3_U3897, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6399, n6400, n6401, n6402, n6403, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837;

  NAND2_X1 U7147 ( .A1(n7479), .A2(n6503), .ZN(n13179) );
  INV_X4 U7148 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  CLKBUF_X2 U7149 ( .A(n12225), .Z(n6446) );
  NAND2_X1 U7150 ( .A1(n6685), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8431) );
  INV_X2 U7151 ( .A(n10936), .ZN(n13139) );
  INV_X1 U7152 ( .A(n6403), .ZN(n6406) );
  BUF_X2 U7153 ( .A(n6402), .Z(n13492) );
  INV_X2 U7154 ( .A(n10554), .ZN(n6409) );
  INV_X2 U7155 ( .A(n10810), .ZN(n9380) );
  NAND2_X1 U7156 ( .A1(n12418), .A2(n12422), .ZN(n12414) );
  NAND2_X2 U7158 ( .A1(n7992), .A2(n7994), .ZN(n8595) );
  AND2_X1 U7159 ( .A1(n10296), .A2(n8209), .ZN(n8055) );
  OAI21_X1 U7160 ( .B1(n8209), .B2(n10161), .A(n6425), .ZN(n8087) );
  NOR2_X1 U7162 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8006) );
  NAND2_X1 U7163 ( .A1(n8209), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n6425) );
  INV_X4 U7164 ( .A(n6402), .ZN(n6440) );
  NOR2_X1 U7165 ( .A1(n15335), .A2(n14107), .ZN(n14326) );
  NOR2_X1 U7166 ( .A1(n15263), .A2(n15261), .ZN(n11029) );
  NOR2_X1 U7167 ( .A1(n9817), .A2(n10025), .ZN(n6965) );
  INV_X2 U7168 ( .A(n10717), .ZN(n10936) );
  NAND2_X1 U7169 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n8095) );
  AND2_X1 U7170 ( .A1(n10884), .A2(n13578), .ZN(n10554) );
  INV_X1 U7171 ( .A(n9418), .ZN(n9395) );
  AND2_X1 U7172 ( .A1(n14759), .A2(n14760), .ZN(n15041) );
  XNOR2_X1 U7173 ( .A(n11571), .B(n6410), .ZN(n14510) );
  INV_X1 U7174 ( .A(n9591), .ZN(n9991) );
  INV_X1 U7175 ( .A(n6443), .ZN(n12360) );
  INV_X1 U7177 ( .A(n9291), .ZN(n10243) );
  INV_X1 U7178 ( .A(n14482), .ZN(n10825) );
  NAND2_X1 U7179 ( .A1(n11054), .A2(n14148), .ZN(n14303) );
  INV_X1 U7180 ( .A(n14325), .ZN(n6410) );
  XNOR2_X1 U7181 ( .A(n8208), .B(SI_10_), .ZN(n8205) );
  OAI21_X1 U7182 ( .B1(n8209), .B2(n10157), .A(n7340), .ZN(n8068) );
  NAND2_X1 U7183 ( .A1(n13075), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9500) );
  NAND2_X2 U7184 ( .A1(n8281), .A2(n8280), .ZN(n14009) );
  OR2_X1 U7185 ( .A1(n13218), .A2(n13110), .ZN(n13219) );
  INV_X1 U7186 ( .A(n13294), .ZN(n13579) );
  INV_X1 U7187 ( .A(n6403), .ZN(n6405) );
  NAND2_X1 U7188 ( .A1(n7363), .A2(n8393), .ZN(n14065) );
  NAND2_X1 U7189 ( .A1(n6579), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8851) );
  XNOR2_X1 U7190 ( .A(n8068), .B(SI_3_), .ZN(n8067) );
  XNOR2_X1 U7191 ( .A(n8392), .B(P2_IR_REG_19__SCAN_IN), .ZN(n13672) );
  AOI21_X1 U7192 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n8748), .A(n15830), .ZN(
        n15822) );
  NAND2_X1 U7193 ( .A1(n15228), .A2(n15445), .ZN(n15227) );
  OR2_X1 U7194 ( .A1(n7393), .A2(n6943), .ZN(n6399) );
  OR2_X1 U7195 ( .A1(n8052), .A2(n10150), .ZN(n6400) );
  AND2_X1 U7196 ( .A1(n7631), .A2(n6538), .ZN(n6401) );
  AND3_X1 U7197 ( .A1(n7901), .A2(n13294), .A3(n13672), .ZN(n6402) );
  OR2_X2 U7198 ( .A1(n8469), .A2(n11335), .ZN(n8416) );
  NAND2_X2 U7199 ( .A1(n8415), .A2(n8414), .ZN(n8469) );
  NAND2_X1 U7200 ( .A1(n6714), .A2(n8908), .ZN(n9453) );
  INV_X1 U7201 ( .A(n8039), .ZN(n8017) );
  NAND2_X2 U7202 ( .A1(n9733), .A2(n9732), .ZN(n9752) );
  INV_X2 U7203 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n15703) );
  OAI21_X2 U7204 ( .B1(n11842), .B2(n11841), .A(n11843), .ZN(n11928) );
  NAND2_X2 U7205 ( .A1(n11802), .A2(n11801), .ZN(n11842) );
  XNOR2_X2 U7206 ( .A(n12638), .B(n12646), .ZN(n12636) );
  NAND2_X2 U7207 ( .A1(n7037), .A2(n12611), .ZN(n12638) );
  AOI21_X2 U7208 ( .B1(n6998), .B2(n6996), .A(n6585), .ZN(n6995) );
  XNOR2_X2 U7209 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n6829) );
  AND2_X2 U7210 ( .A1(n12424), .A2(n12419), .ZN(n12526) );
  NOR4_X2 U7211 ( .A1(n14927), .A2(n14950), .A3(n14998), .A4(n14518), .ZN(
        n14519) );
  XNOR2_X2 U7212 ( .A(n8851), .B(n8850), .ZN(n14482) );
  XNOR2_X2 U7213 ( .A(n14009), .B(n13386), .ZN(n13889) );
  INV_X1 U7214 ( .A(n15261), .ZN(n15286) );
  OAI211_X2 U7215 ( .C1(n6434), .C2(n10267), .A(n8935), .B(n8934), .ZN(n15261)
         );
  NAND2_X2 U7216 ( .A1(n9489), .A2(n9490), .ZN(n13081) );
  NAND2_X4 U7217 ( .A1(n9022), .A2(n9021), .ZN(n14325) );
  AOI21_X2 U7218 ( .B1(n12910), .B2(n12914), .A(n12470), .ZN(n12900) );
  XNOR2_X2 U7219 ( .A(n12593), .B(n12600), .ZN(n12594) );
  NAND2_X2 U7220 ( .A1(n7202), .A2(n11690), .ZN(n12593) );
  XNOR2_X2 U7221 ( .A(n8868), .B(n8867), .ZN(n8871) );
  AOI21_X2 U7222 ( .B1(n7650), .B2(n7652), .A(n6569), .ZN(n7649) );
  INV_X1 U7223 ( .A(n10554), .ZN(n6403) );
  NAND2_X1 U7225 ( .A1(n6513), .A2(n12778), .ZN(n12934) );
  AOI21_X1 U7226 ( .B1(n12511), .B2(n12510), .A(n7317), .ZN(n7316) );
  NAND2_X1 U7227 ( .A1(n7348), .A2(n7357), .ZN(n13155) );
  NAND2_X1 U7228 ( .A1(n6704), .A2(n6708), .ZN(n12791) );
  NAND2_X1 U7229 ( .A1(n14945), .A2(n14943), .ZN(n14926) );
  NAND2_X1 U7230 ( .A1(n9331), .A2(n9330), .ZN(n14840) );
  NAND2_X1 U7231 ( .A1(n6653), .A2(n9121), .ZN(n15149) );
  INV_X1 U7232 ( .A(n11729), .ZN(n6407) );
  AND2_X1 U7233 ( .A1(n10077), .A2(n12436), .ZN(n11265) );
  INV_X2 U7234 ( .A(n6445), .ZN(n12220) );
  INV_X1 U7235 ( .A(n12414), .ZN(n7416) );
  INV_X1 U7236 ( .A(n14319), .ZN(n11406) );
  INV_X2 U7237 ( .A(n14993), .ZN(n6408) );
  NAND2_X1 U7238 ( .A1(n14302), .A2(n14303), .ZN(n11052) );
  NAND2_X2 U7239 ( .A1(n7169), .A2(n10643), .ZN(n12407) );
  NAND2_X1 U7240 ( .A1(n8988), .A2(n8987), .ZN(n14313) );
  NAND2_X1 U7241 ( .A1(n9645), .A2(n9644), .ZN(n12435) );
  NAND3_X2 U7242 ( .A1(n9541), .A2(n7138), .A3(n7643), .ZN(n12580) );
  INV_X1 U7243 ( .A(n14551), .ZN(n14107) );
  INV_X1 U7244 ( .A(n14554), .ZN(n11402) );
  BUF_X2 U7245 ( .A(n9533), .Z(n12583) );
  INV_X1 U7246 ( .A(n9514), .ZN(n7152) );
  NAND2_X1 U7247 ( .A1(n12584), .A2(n7809), .ZN(n10737) );
  AND3_X1 U7248 ( .A1(n8929), .A2(n8927), .A3(n8928), .ZN(n7797) );
  CLKBUF_X2 U7249 ( .A(n14312), .Z(n14441) );
  AND2_X1 U7250 ( .A1(n9540), .A2(n9539), .ZN(n7138) );
  NAND4_X1 U7251 ( .A1(n8083), .A2(n8082), .A3(n8081), .A4(n8080), .ZN(n13608)
         );
  INV_X1 U7252 ( .A(n13609), .ZN(n7395) );
  NOR2_X2 U7253 ( .A1(n10824), .A2(n10825), .ZN(n15264) );
  INV_X2 U7254 ( .A(n11937), .ZN(n9504) );
  AND2_X1 U7255 ( .A1(n14483), .A2(n14482), .ZN(n14292) );
  INV_X2 U7257 ( .A(n12201), .ZN(n7069) );
  INV_X4 U7258 ( .A(n8398), .ZN(n8596) );
  INV_X1 U7260 ( .A(n13578), .ZN(n7902) );
  INV_X2 U7261 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n10140) );
  NAND2_X1 U7262 ( .A1(n7506), .A2(n7505), .ZN(n14487) );
  OAI211_X1 U7263 ( .C1(n8700), .C2(n14040), .A(n8698), .B(n8699), .ZN(n13931)
         );
  XNOR2_X1 U7264 ( .A(n6432), .B(n13565), .ZN(n8700) );
  AOI21_X1 U7265 ( .B1(n12118), .B2(n15311), .A(n12117), .ZN(n15063) );
  OAI21_X1 U7266 ( .B1(n7706), .B2(n10085), .A(n7705), .ZN(n6673) );
  NAND2_X1 U7267 ( .A1(n8804), .A2(n8683), .ZN(n6432) );
  AND3_X1 U7268 ( .A1(n6431), .A2(n7034), .A3(n8612), .ZN(n8699) );
  NOR2_X1 U7269 ( .A1(n14813), .A2(n14812), .ZN(n14814) );
  NAND2_X1 U7270 ( .A1(n8807), .A2(n8604), .ZN(n6431) );
  NAND2_X1 U7271 ( .A1(n13699), .A2(n8682), .ZN(n8801) );
  NAND2_X1 U7272 ( .A1(n7006), .A2(n6534), .ZN(n13148) );
  NAND2_X1 U7273 ( .A1(n14829), .A2(n12104), .ZN(n14813) );
  NAND2_X1 U7274 ( .A1(n7874), .A2(n6550), .ZN(n13524) );
  NOR3_X1 U7275 ( .A1(n15075), .A2(n15074), .A3(n15073), .ZN(n7213) );
  OR2_X1 U7276 ( .A1(n12753), .A2(n15570), .ZN(n6962) );
  INV_X1 U7277 ( .A(n13488), .ZN(n7874) );
  NAND2_X1 U7278 ( .A1(n14849), .A2(n6423), .ZN(n14829) );
  AND2_X1 U7279 ( .A1(n14849), .A2(n12107), .ZN(n14831) );
  NAND2_X1 U7280 ( .A1(n13698), .A2(n13697), .ZN(n13699) );
  AOI21_X1 U7281 ( .B1(n7223), .B2(n7222), .A(n12774), .ZN(n12999) );
  OR2_X1 U7282 ( .A1(n13179), .A2(n12010), .ZN(n7010) );
  OR3_X1 U7283 ( .A1(n13963), .A2(n13962), .A3(n13961), .ZN(n14056) );
  NAND2_X1 U7284 ( .A1(n6429), .A2(n6399), .ZN(n13698) );
  NAND2_X1 U7285 ( .A1(n6762), .A2(n6500), .ZN(n14749) );
  AND2_X1 U7286 ( .A1(n6711), .A2(n7227), .ZN(n6486) );
  OR2_X1 U7287 ( .A1(n7708), .A2(n6915), .ZN(n6914) );
  AND2_X1 U7288 ( .A1(n10105), .A2(n7665), .ZN(n7664) );
  AOI21_X1 U7289 ( .B1(n10092), .B2(n10091), .A(n10090), .ZN(n10093) );
  NAND2_X1 U7290 ( .A1(n6944), .A2(n6460), .ZN(n6429) );
  NOR3_X1 U7291 ( .A1(n13683), .A2(n6409), .A3(n6882), .ZN(n8697) );
  NAND2_X1 U7292 ( .A1(n14847), .A2(n14848), .ZN(n6670) );
  NAND2_X1 U7293 ( .A1(n6830), .A2(n8787), .ZN(n15242) );
  NAND2_X1 U7294 ( .A1(n15243), .A2(n15485), .ZN(n15240) );
  OR2_X1 U7295 ( .A1(n12767), .A2(n13065), .ZN(n10105) );
  NAND2_X1 U7296 ( .A1(n12100), .A2(n6422), .ZN(n14847) );
  XNOR2_X1 U7297 ( .A(n12298), .B(n12235), .ZN(n12299) );
  NAND2_X1 U7298 ( .A1(n12100), .A2(n12099), .ZN(n14866) );
  OR2_X1 U7299 ( .A1(n12352), .A2(n12351), .ZN(n12384) );
  INV_X1 U7300 ( .A(n6831), .ZN(n6830) );
  XNOR2_X1 U7301 ( .A(n12352), .B(n9999), .ZN(n12767) );
  NAND2_X1 U7302 ( .A1(n12135), .A2(n12134), .ZN(n14861) );
  NOR2_X1 U7303 ( .A1(n7316), .A2(n12781), .ZN(n7183) );
  NAND2_X1 U7304 ( .A1(n12038), .A2(n12037), .ZN(n14499) );
  NAND2_X1 U7305 ( .A1(n6831), .A2(n7639), .ZN(n15243) );
  OAI21_X1 U7306 ( .B1(n12219), .B2(n7862), .A(n7860), .ZN(n12338) );
  OAI21_X1 U7307 ( .B1(n12809), .B2(n7661), .A(n7659), .ZN(n12782) );
  NAND2_X1 U7308 ( .A1(n7829), .A2(n7827), .ZN(n12352) );
  AND2_X1 U7309 ( .A1(n7087), .A2(n6455), .ZN(n12298) );
  NAND2_X1 U7310 ( .A1(n13446), .A2(n12035), .ZN(n14095) );
  NAND2_X1 U7311 ( .A1(n13450), .A2(n13449), .ZN(n13676) );
  OAI21_X1 U7312 ( .B1(n7687), .B2(n7392), .A(n8681), .ZN(n7391) );
  NAND2_X1 U7313 ( .A1(n7253), .A2(n7257), .ZN(n7551) );
  INV_X1 U7314 ( .A(n7348), .ZN(n13154) );
  AOI21_X1 U7315 ( .B1(n7690), .B2(n7688), .A(n6572), .ZN(n7687) );
  NAND2_X1 U7316 ( .A1(n8594), .A2(n8593), .ZN(n13460) );
  AND2_X1 U7317 ( .A1(n14867), .A2(n14869), .ZN(n12133) );
  OAI21_X1 U7318 ( .B1(n7574), .B2(n7573), .A(n14243), .ZN(n7572) );
  NAND2_X1 U7319 ( .A1(n8784), .A2(n8783), .ZN(n15239) );
  NAND2_X1 U7320 ( .A1(n12027), .A2(n12026), .ZN(n14758) );
  XNOR2_X1 U7321 ( .A(n6418), .B(n13448), .ZN(n14474) );
  NAND2_X1 U7322 ( .A1(n14252), .A2(n6995), .ZN(n6994) );
  NAND2_X1 U7323 ( .A1(n9400), .A2(n9399), .ZN(n14787) );
  AND2_X1 U7324 ( .A1(n12102), .A2(n12099), .ZN(n6422) );
  NAND2_X1 U7325 ( .A1(n6659), .A2(n6658), .ZN(n14867) );
  NOR2_X1 U7326 ( .A1(n7689), .A2(n8462), .ZN(n7394) );
  INV_X1 U7327 ( .A(n7689), .ZN(n7690) );
  INV_X1 U7328 ( .A(n14885), .ZN(n6659) );
  OAI21_X1 U7329 ( .B1(n12029), .B2(n7896), .A(n7893), .ZN(n6418) );
  XNOR2_X1 U7330 ( .A(n12029), .B(n12028), .ZN(n14098) );
  AOI21_X1 U7331 ( .B1(n7491), .B2(n6453), .A(n6582), .ZN(n7490) );
  NAND2_X1 U7332 ( .A1(n13736), .A2(n13535), .ZN(n7689) );
  AND3_X1 U7333 ( .A1(n6876), .A2(n6878), .A3(n6875), .ZN(n13753) );
  AND2_X1 U7334 ( .A1(n7339), .A2(n13202), .ZN(n7491) );
  INV_X1 U7335 ( .A(n14222), .ZN(n6993) );
  OAI21_X1 U7336 ( .B1(n7283), .B2(n13382), .A(n7281), .ZN(n7909) );
  AND2_X1 U7337 ( .A1(n14830), .A2(n12107), .ZN(n6423) );
  AND2_X1 U7338 ( .A1(n14887), .A2(n14884), .ZN(n14885) );
  NAND2_X1 U7339 ( .A1(n14947), .A2(n14390), .ZN(n14945) );
  NAND2_X1 U7340 ( .A1(n8592), .A2(n8591), .ZN(n12029) );
  NOR2_X1 U7341 ( .A1(n15479), .A2(n15478), .ZN(n15477) );
  NAND2_X1 U7342 ( .A1(n9368), .A2(n9367), .ZN(n15060) );
  XNOR2_X1 U7343 ( .A(n14840), .B(n14542), .ZN(n14830) );
  NAND2_X1 U7344 ( .A1(n8531), .A2(n8530), .ZN(n13940) );
  XNOR2_X1 U7345 ( .A(n13948), .B(n13475), .ZN(n13736) );
  OR2_X1 U7346 ( .A1(n11987), .A2(n6453), .ZN(n7339) );
  NAND2_X1 U7347 ( .A1(n6700), .A2(n6561), .ZN(n7419) );
  NAND2_X1 U7348 ( .A1(n7128), .A2(n7127), .ZN(n8592) );
  XNOR2_X1 U7349 ( .A(n8560), .B(n8545), .ZN(n11806) );
  NAND2_X1 U7350 ( .A1(n14967), .A2(n12096), .ZN(n14947) );
  NAND2_X1 U7351 ( .A1(n7782), .A2(n6610), .ZN(n14967) );
  NAND3_X1 U7352 ( .A1(n6511), .A2(n7583), .A3(n9175), .ZN(n14122) );
  AND2_X1 U7353 ( .A1(n13133), .A2(n11986), .ZN(n11987) );
  OR2_X1 U7354 ( .A1(n13791), .A2(n13421), .ZN(n7387) );
  NAND2_X1 U7355 ( .A1(n8452), .A2(n8451), .ZN(n14058) );
  NAND2_X1 U7356 ( .A1(n6583), .A2(n14402), .ZN(n7801) );
  AND2_X1 U7357 ( .A1(n8502), .A2(n8501), .ZN(n13475) );
  AOI21_X1 U7358 ( .B1(n13652), .B2(n13651), .A(n15459), .ZN(n15479) );
  AND2_X1 U7359 ( .A1(n7580), .A2(n9221), .ZN(n7579) );
  NAND2_X1 U7360 ( .A1(n9350), .A2(n9349), .ZN(n15065) );
  XNOR2_X1 U7361 ( .A(n9290), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n15197) );
  OAI21_X1 U7362 ( .B1(n8544), .B2(n7886), .A(n7884), .ZN(n8566) );
  NAND2_X1 U7363 ( .A1(n11864), .A2(n7582), .ZN(n7583) );
  NAND2_X1 U7364 ( .A1(n9309), .A2(n9308), .ZN(n15078) );
  AND2_X1 U7365 ( .A1(n8487), .A2(n8486), .ZN(n13437) );
  NAND2_X1 U7366 ( .A1(n8524), .A2(n8523), .ZN(n13592) );
  NAND2_X1 U7367 ( .A1(n8479), .A2(n8478), .ZN(n13956) );
  NAND2_X1 U7368 ( .A1(n6696), .A2(n6694), .ZN(n12862) );
  NAND2_X1 U7369 ( .A1(n8429), .A2(n8428), .ZN(n13432) );
  NAND2_X1 U7370 ( .A1(n8518), .A2(n8517), .ZN(n13722) );
  XNOR2_X1 U7371 ( .A(n15096), .B(n14545), .ZN(n14907) );
  NAND2_X1 U7372 ( .A1(n6417), .A2(n8528), .ZN(n8544) );
  OR2_X1 U7373 ( .A1(n13906), .A2(n6951), .ZN(n6955) );
  NOR2_X1 U7374 ( .A1(n9150), .A2(n7584), .ZN(n7582) );
  XNOR2_X1 U7375 ( .A(n6433), .B(n8492), .ZN(n11562) );
  NAND2_X1 U7376 ( .A1(n8418), .A2(n8417), .ZN(n13972) );
  XNOR2_X1 U7377 ( .A(n8427), .B(n8440), .ZN(n11493) );
  OAI21_X1 U7378 ( .B1(n8490), .B2(n11745), .A(n8491), .ZN(n6433) );
  OR2_X1 U7379 ( .A1(n8527), .A2(n8526), .ZN(n6417) );
  NAND2_X1 U7380 ( .A1(n11958), .A2(n12084), .ZN(n12090) );
  OAI211_X1 U7381 ( .C1(n7363), .C2(n13139), .A(n7360), .B(n7359), .ZN(n13204)
         );
  OR2_X1 U7382 ( .A1(n15230), .A2(n7313), .ZN(n7311) );
  NAND2_X1 U7383 ( .A1(n6414), .A2(n8513), .ZN(n8527) );
  NAND2_X1 U7384 ( .A1(n11775), .A2(n7323), .ZN(n11778) );
  AND2_X1 U7385 ( .A1(n6952), .A2(n6615), .ZN(n6956) );
  XNOR2_X1 U7386 ( .A(n8426), .B(n8441), .ZN(n11454) );
  NAND2_X1 U7387 ( .A1(n8348), .A2(n8347), .ZN(n13821) );
  NAND2_X1 U7388 ( .A1(n8477), .A2(n6415), .ZN(n6414) );
  NAND2_X1 U7389 ( .A1(n11214), .A2(n8146), .ZN(n7363) );
  NAND2_X1 U7390 ( .A1(n9230), .A2(n9229), .ZN(n15109) );
  NAND2_X1 U7391 ( .A1(n8425), .A2(n8416), .ZN(n8426) );
  INV_X1 U7392 ( .A(n14361), .ZN(n15006) );
  AND2_X1 U7393 ( .A1(n14386), .A2(n14368), .ZN(n14987) );
  NAND2_X1 U7394 ( .A1(n8477), .A2(n8476), .ZN(n8506) );
  XNOR2_X1 U7395 ( .A(n8386), .B(n8385), .ZN(n11214) );
  OR2_X1 U7396 ( .A1(n15130), .A2(n14370), .ZN(n14386) );
  NAND2_X1 U7397 ( .A1(n6960), .A2(n8668), .ZN(n6958) );
  NAND2_X1 U7398 ( .A1(n8364), .A2(n8363), .ZN(n14073) );
  NAND2_X1 U7399 ( .A1(n8469), .A2(n8468), .ZN(n8477) );
  NAND2_X1 U7400 ( .A1(n8839), .A2(n8838), .ZN(n14960) );
  NAND2_X1 U7401 ( .A1(n11794), .A2(n11793), .ZN(n11849) );
  OAI22_X1 U7402 ( .A1(n8382), .A2(n8405), .B1(n8408), .B2(n11103), .ZN(n8386)
         );
  OR2_X1 U7403 ( .A1(n13357), .A2(n13356), .ZN(n13362) );
  NAND2_X1 U7404 ( .A1(n8300), .A2(n8299), .ZN(n13866) );
  NAND2_X1 U7405 ( .A1(n9202), .A2(n9201), .ZN(n15130) );
  XNOR2_X1 U7406 ( .A(n13365), .B(n13601), .ZN(n11729) );
  NAND2_X1 U7407 ( .A1(n9181), .A2(n9180), .ZN(n15122) );
  NAND2_X1 U7408 ( .A1(n9856), .A2(n9855), .ZN(n13038) );
  NAND2_X1 U7409 ( .A1(n8238), .A2(n8237), .ZN(n14085) );
  NAND2_X1 U7410 ( .A1(n8408), .A2(n8407), .ZN(n8415) );
  AOI21_X1 U7411 ( .B1(n7020), .B2(n11359), .A(n7019), .ZN(n7018) );
  NAND2_X1 U7412 ( .A1(n8324), .A2(n8323), .ZN(n13996) );
  NAND2_X1 U7413 ( .A1(n6419), .A2(n7880), .ZN(n8408) );
  NAND2_X1 U7414 ( .A1(n10498), .A2(n8962), .ZN(n6653) );
  XNOR2_X1 U7415 ( .A(n8295), .B(n8294), .ZN(n10829) );
  AOI21_X1 U7416 ( .B1(n8359), .B2(n6472), .A(n8344), .ZN(n7358) );
  NAND2_X2 U7417 ( .A1(n8215), .A2(n8214), .ZN(n13365) );
  NAND2_X1 U7418 ( .A1(n7002), .A2(n9141), .ZN(n15144) );
  XNOR2_X1 U7419 ( .A(n14350), .B(n14549), .ZN(n11799) );
  NAND2_X1 U7420 ( .A1(n8337), .A2(n7881), .ZN(n6419) );
  XNOR2_X1 U7421 ( .A(n8290), .B(n8308), .ZN(n10763) );
  XNOR2_X1 U7422 ( .A(n6669), .B(n8258), .ZN(n10498) );
  NOR2_X1 U7423 ( .A1(n14026), .A2(n13352), .ZN(n7767) );
  OAI21_X1 U7424 ( .B1(n8290), .B2(n8308), .A(n8289), .ZN(n8295) );
  OAI21_X1 U7425 ( .B1(n8227), .B2(n8226), .A(n8254), .ZN(n6669) );
  NAND2_X1 U7426 ( .A1(n8277), .A2(n8289), .ZN(n8290) );
  AND2_X1 U7427 ( .A1(n7844), .A2(n7842), .ZN(n7841) );
  AND2_X1 U7428 ( .A1(n7612), .A2(n7613), .ZN(n15588) );
  NAND2_X1 U7429 ( .A1(n8314), .A2(n8313), .ZN(n8337) );
  NAND2_X1 U7430 ( .A1(n8196), .A2(n8195), .ZN(n14026) );
  NAND2_X1 U7431 ( .A1(n6426), .A2(n9075), .ZN(n14350) );
  XNOR2_X1 U7432 ( .A(n8227), .B(n8226), .ZN(n10457) );
  INV_X1 U7433 ( .A(n12286), .ZN(n13062) );
  NAND2_X1 U7434 ( .A1(n8349), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8368) );
  NAND2_X1 U7435 ( .A1(n10284), .A2(n8962), .ZN(n6426) );
  NAND2_X1 U7436 ( .A1(n8253), .A2(n8249), .ZN(n8227) );
  AOI21_X1 U7437 ( .B1(n7083), .B2(n7081), .A(n6524), .ZN(n7080) );
  OR2_X1 U7438 ( .A1(n8312), .A2(n10497), .ZN(n8277) );
  NAND2_X1 U7439 ( .A1(n7411), .A2(n7412), .ZN(n10961) );
  NAND2_X1 U7440 ( .A1(n9059), .A2(n9058), .ZN(n14344) );
  INV_X1 U7441 ( .A(n12534), .ZN(n7081) );
  NAND2_X1 U7442 ( .A1(n8193), .A2(n7878), .ZN(n7877) );
  XNOR2_X1 U7443 ( .A(n11220), .B(n11228), .ZN(n11218) );
  NAND2_X1 U7444 ( .A1(n12443), .A2(n12442), .ZN(n12534) );
  NOR2_X1 U7445 ( .A1(n6408), .A2(n10903), .ZN(n15024) );
  XNOR2_X1 U7446 ( .A(n8190), .B(n8188), .ZN(n10239) );
  NAND2_X1 U7447 ( .A1(n15540), .A2(n10687), .ZN(n11220) );
  OR2_X1 U7448 ( .A1(n9766), .A2(n9765), .ZN(n7736) );
  NAND2_X1 U7449 ( .A1(n8190), .A2(n8189), .ZN(n8193) );
  NAND2_X1 U7450 ( .A1(n9037), .A2(n9036), .ZN(n15335) );
  INV_X1 U7451 ( .A(n12532), .ZN(n11267) );
  NAND2_X1 U7452 ( .A1(n9754), .A2(n9753), .ZN(n9766) );
  NAND2_X1 U7453 ( .A1(n6421), .A2(n8168), .ZN(n8190) );
  NAND2_X1 U7454 ( .A1(n8111), .A2(n8110), .ZN(n14036) );
  INV_X1 U7455 ( .A(n11052), .ZN(n14503) );
  NAND2_X1 U7456 ( .A1(n8129), .A2(n8128), .ZN(n15525) );
  CLKBUF_X3 U7457 ( .A(n12225), .Z(n6445) );
  OR2_X1 U7458 ( .A1(n11520), .A2(n12574), .ZN(n12454) );
  AND2_X1 U7459 ( .A1(n12439), .A2(n6461), .ZN(n12532) );
  OAI21_X1 U7460 ( .B1(n7617), .B2(n10447), .A(n7616), .ZN(n15545) );
  NAND2_X1 U7461 ( .A1(n10581), .A2(n10580), .ZN(n12225) );
  XNOR2_X1 U7462 ( .A(n11096), .B(n12579), .ZN(n12524) );
  XNOR2_X1 U7463 ( .A(n10683), .B(n10431), .ZN(n10681) );
  AND2_X1 U7464 ( .A1(n9603), .A2(n7134), .ZN(n9604) );
  NAND2_X1 U7465 ( .A1(n9622), .A2(n9621), .ZN(n11096) );
  AND2_X1 U7466 ( .A1(n7807), .A2(n7809), .ZN(n7808) );
  OAI21_X1 U7467 ( .B1(n6495), .B2(n7346), .A(n8276), .ZN(n7345) );
  INV_X1 U7468 ( .A(n14148), .ZN(n15293) );
  NAND2_X1 U7469 ( .A1(n10430), .A2(n10429), .ZN(n10683) );
  NAND2_X1 U7470 ( .A1(n8125), .A2(n8124), .ZN(n8143) );
  INV_X1 U7471 ( .A(n14556), .ZN(n11054) );
  NAND2_X2 U7472 ( .A1(n8930), .A2(n7797), .ZN(n14557) );
  INV_X2 U7473 ( .A(n6494), .ZN(n9397) );
  OAI211_X1 U7474 ( .C1(n9291), .C2(n14589), .A(n8948), .B(n8947), .ZN(n14148)
         );
  AND2_X2 U7475 ( .A1(n10107), .A2(n10244), .ZN(P1_U4016) );
  AND2_X1 U7476 ( .A1(n6760), .A2(n9028), .ZN(n11571) );
  OAI211_X1 U7477 ( .C1(SI_5_), .C2(n9989), .A(n9574), .B(n9573), .ZN(n10985)
         );
  INV_X1 U7478 ( .A(n12980), .ZN(n6411) );
  INV_X1 U7479 ( .A(n15512), .ZN(n6751) );
  NAND4_X2 U7480 ( .A1(n9632), .A2(n9631), .A3(n9630), .A4(n9629), .ZN(n12579)
         );
  NAND4_X1 U7481 ( .A1(n9508), .A2(n9506), .A3(n9505), .A4(n9507), .ZN(n12584)
         );
  AND3_X1 U7482 ( .A1(n8882), .A2(n8881), .A3(n8880), .ZN(n8883) );
  NAND4_X2 U7483 ( .A1(n8961), .A2(n8960), .A3(n8959), .A4(n8958), .ZN(n14555)
         );
  AOI21_X1 U7484 ( .B1(n7881), .B2(n7883), .A(n8340), .ZN(n7880) );
  NAND4_X2 U7485 ( .A1(n8983), .A2(n8982), .A3(n8981), .A4(n8980), .ZN(n14554)
         );
  AND2_X1 U7486 ( .A1(n8476), .A2(n6416), .ZN(n6415) );
  INV_X1 U7487 ( .A(n7167), .ZN(n12368) );
  OR2_X1 U7488 ( .A1(n6437), .A2(n8924), .ZN(n8929) );
  AND2_X1 U7489 ( .A1(n7879), .A2(n8252), .ZN(n7878) );
  INV_X2 U7490 ( .A(n8174), .ZN(n13496) );
  INV_X2 U7491 ( .A(n9846), .ZN(n6442) );
  INV_X1 U7492 ( .A(n9522), .ZN(n9617) );
  CLKBUF_X3 U7493 ( .A(n14312), .Z(n6412) );
  AND2_X2 U7494 ( .A1(n8876), .A2(n10808), .ZN(n10810) );
  OAI21_X1 U7495 ( .B1(n8077), .B2(n7292), .A(n6477), .ZN(n13606) );
  AOI21_X1 U7496 ( .B1(n8475), .B2(n8474), .A(n8473), .ZN(n8476) );
  INV_X1 U7497 ( .A(n7882), .ZN(n7881) );
  NAND2_X1 U7498 ( .A1(n8848), .A2(n10182), .ZN(n10106) );
  XNOR2_X1 U7499 ( .A(n8066), .B(n8067), .ZN(n10167) );
  AND2_X1 U7500 ( .A1(n7542), .A2(n6400), .ZN(n8066) );
  INV_X2 U7501 ( .A(n9207), .ZN(n14427) );
  CLKBUF_X2 U7502 ( .A(n10015), .Z(n6443) );
  AND2_X1 U7503 ( .A1(n9425), .A2(n9430), .ZN(n8848) );
  CLKBUF_X3 U7504 ( .A(n9453), .Z(n6439) );
  AND2_X1 U7505 ( .A1(n8911), .A2(n8910), .ZN(n10904) );
  INV_X2 U7506 ( .A(n8077), .ZN(n8597) );
  AND4_X1 U7507 ( .A1(n8027), .A2(n8026), .A3(n8025), .A4(n8024), .ZN(n13293)
         );
  CLKBUF_X1 U7508 ( .A(n9453), .Z(n6437) );
  OAI21_X1 U7509 ( .B1(n9568), .B2(n7720), .A(n7717), .ZN(n9656) );
  INV_X1 U7510 ( .A(n8505), .ZN(n6416) );
  NAND2_X2 U7511 ( .A1(n7069), .A2(n11937), .ZN(n10015) );
  NAND2_X1 U7512 ( .A1(n13580), .A2(n13578), .ZN(n13571) );
  AND2_X1 U7513 ( .A1(n11461), .A2(n10097), .ZN(n12549) );
  INV_X1 U7514 ( .A(n8925), .ZN(n9207) );
  XNOR2_X1 U7515 ( .A(n9840), .B(P3_IR_REG_19__SCAN_IN), .ZN(n12548) );
  AND2_X1 U7516 ( .A1(n10010), .A2(n10009), .ZN(n10097) );
  INV_X1 U7517 ( .A(n8871), .ZN(n8908) );
  NAND2_X1 U7518 ( .A1(n8844), .A2(n8846), .ZN(n11564) );
  OR2_X1 U7519 ( .A1(n8205), .A2(n8192), .ZN(n7879) );
  NOR2_X1 U7520 ( .A1(n13284), .A2(n7902), .ZN(n7901) );
  INV_X1 U7521 ( .A(n8085), .ZN(n8084) );
  XNOR2_X1 U7522 ( .A(n9556), .B(n9555), .ZN(n15550) );
  XNOR2_X1 U7523 ( .A(n8087), .B(n6424), .ZN(n8085) );
  NAND2_X1 U7524 ( .A1(n6712), .A2(n7136), .ZN(n9489) );
  XNOR2_X1 U7525 ( .A(n8849), .B(P1_IR_REG_21__SCAN_IN), .ZN(n14483) );
  NAND2_X1 U7526 ( .A1(n7675), .A2(n7672), .ZN(n12205) );
  INV_X1 U7527 ( .A(n12202), .ZN(n6714) );
  XNOR2_X1 U7528 ( .A(n7004), .B(n15784), .ZN(n13294) );
  NAND2_X1 U7529 ( .A1(n8583), .A2(n8613), .ZN(n13284) );
  INV_X1 U7530 ( .A(n7992), .ZN(n14096) );
  XNOR2_X1 U7531 ( .A(n10006), .B(P3_IR_REG_22__SCAN_IN), .ZN(n12560) );
  NAND2_X1 U7532 ( .A1(n8866), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8868) );
  OR2_X1 U7533 ( .A1(n9588), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U7534 ( .A1(n8613), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7004) );
  XNOR2_X1 U7535 ( .A(n8106), .B(SI_5_), .ZN(n8103) );
  NAND2_X2 U7536 ( .A1(n7875), .A2(P1_U3086), .ZN(n15189) );
  NAND2_X2 U7537 ( .A1(n7875), .A2(P2_U3088), .ZN(n14099) );
  MUX2_X1 U7538 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9492), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n7172) );
  XNOR2_X1 U7539 ( .A(n10036), .B(P3_IR_REG_26__SCAN_IN), .ZN(n10048) );
  OR2_X1 U7540 ( .A1(n9501), .A2(n13074), .ZN(n7338) );
  NAND2_X1 U7541 ( .A1(n8825), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U7542 ( .A1(n9602), .A2(n9601), .ZN(n10680) );
  OAI21_X1 U7543 ( .B1(n10042), .B2(P3_IR_REG_25__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n10036) );
  XNOR2_X1 U7544 ( .A(n8052), .B(SI_2_), .ZN(n8053) );
  OR2_X1 U7545 ( .A1(n8588), .A2(n6543), .ZN(n7675) );
  NOR2_X1 U7546 ( .A1(n10000), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n9818) );
  AND2_X1 U7547 ( .A1(n6740), .A2(n7954), .ZN(n7586) );
  NAND3_X1 U7548 ( .A1(n7086), .A2(n9640), .A3(n7851), .ZN(n10042) );
  NAND2_X1 U7549 ( .A1(n9637), .A2(n7615), .ZN(n10634) );
  AND2_X1 U7550 ( .A1(n7086), .A2(n9640), .ZN(n10004) );
  AND2_X1 U7551 ( .A1(n8580), .A2(n8584), .ZN(n8588) );
  INV_X1 U7552 ( .A(n8017), .ZN(n6413) );
  NAND3_X1 U7553 ( .A1(n6966), .A2(n6964), .A3(n6965), .ZN(n9491) );
  AND2_X1 U7554 ( .A1(n7850), .A2(n10002), .ZN(n7086) );
  AND4_X1 U7555 ( .A1(n7960), .A2(n8818), .A3(n8827), .A4(n7464), .ZN(n6738)
         );
  NOR2_X1 U7556 ( .A1(n7587), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6740) );
  NOR2_X1 U7557 ( .A1(n8071), .A2(n8001), .ZN(n8580) );
  NOR2_X1 U7558 ( .A1(n7980), .A2(n7979), .ZN(n7981) );
  NOR2_X1 U7559 ( .A1(n7978), .A2(n8108), .ZN(n7982) );
  INV_X1 U7560 ( .A(n8944), .ZN(n8827) );
  NAND2_X1 U7561 ( .A1(n7210), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n6428) );
  NAND2_X1 U7562 ( .A1(n7234), .A2(n7553), .ZN(n7552) );
  NAND2_X1 U7563 ( .A1(n7409), .A2(n9480), .ZN(n9637) );
  NAND4_X1 U7564 ( .A1(n9770), .A2(n9789), .A3(n9485), .A4(n9484), .ZN(n9816)
         );
  AND4_X1 U7565 ( .A1(n8819), .A2(n8853), .A3(n8859), .A4(n8856), .ZN(n7954)
         );
  AND2_X2 U7566 ( .A1(n10140), .A2(n6890), .ZN(n7409) );
  NAND4_X1 U7567 ( .A1(n7983), .A2(n8579), .A3(n15784), .A4(n8634), .ZN(n8622)
         );
  AND4_X1 U7568 ( .A1(n8832), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(n7960)
         );
  NAND3_X1 U7569 ( .A1(n15703), .A2(n9819), .A3(n9481), .ZN(n10001) );
  AND4_X1 U7570 ( .A1(n8834), .A2(n8816), .A3(n8815), .A4(n8828), .ZN(n8818)
         );
  NAND4_X1 U7571 ( .A1(n9478), .A2(n9555), .A3(n9477), .A4(n9476), .ZN(n9638)
         );
  INV_X1 U7572 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n7237) );
  NOR2_X1 U7573 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n8834) );
  NOR2_X1 U7574 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n8819) );
  INV_X1 U7575 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7236) );
  INV_X1 U7576 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n8828) );
  INV_X1 U7577 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7235) );
  NOR2_X1 U7578 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n8815) );
  NOR2_X1 U7579 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8816) );
  NOR2_X1 U7580 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n8812) );
  NOR2_X1 U7581 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n8813) );
  INV_X4 U7582 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7583 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n8859) );
  INV_X1 U7584 ( .A(SI_4_), .ZN(n6424) );
  NOR2_X1 U7585 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8005) );
  NOR2_X1 U7586 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8004) );
  INV_X1 U7587 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8002) );
  INV_X1 U7588 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8003) );
  INV_X4 U7589 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  NOR2_X1 U7590 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n7476) );
  NOR2_X1 U7591 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7477) );
  NOR2_X1 U7592 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n7478) );
  INV_X1 U7593 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7998) );
  INV_X1 U7594 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7977) );
  INV_X1 U7595 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n8072) );
  INV_X1 U7596 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8000) );
  INV_X1 U7597 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n9699) );
  INV_X1 U7598 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8634) );
  NOR2_X1 U7600 ( .A1(P3_IR_REG_7__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n9478) );
  INV_X1 U7601 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n9485) );
  INV_X1 U7602 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n9484) );
  INV_X1 U7603 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n9476) );
  INV_X1 U7604 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n9819) );
  NOR2_X1 U7605 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .ZN(
        n7983) );
  INV_X1 U7606 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n9789) );
  INV_X1 U7607 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n9555) );
  INV_X1 U7608 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n9770) );
  NOR2_X1 U7609 ( .A1(P3_IR_REG_11__SCAN_IN), .A2(P3_IR_REG_9__SCAN_IN), .ZN(
        n9483) );
  NOR2_X1 U7610 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n9482) );
  INV_X1 U7611 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n8579) );
  NAND3_X1 U7612 ( .A1(n6420), .A2(n6552), .A3(n7161), .ZN(n13488) );
  NAND2_X1 U7613 ( .A1(n6420), .A2(n7161), .ZN(n13491) );
  AND2_X1 U7614 ( .A1(n7162), .A2(n13511), .ZN(n6420) );
  MUX2_X1 U7615 ( .A(n10166), .B(n10152), .S(n8039), .Z(n8052) );
  NAND2_X2 U7616 ( .A1(n6428), .A2(n7552), .ZN(n8039) );
  NAND2_X1 U7617 ( .A1(n8166), .A2(n8165), .ZN(n6421) );
  XNOR2_X1 U7618 ( .A(n8207), .B(n8205), .ZN(n10284) );
  NAND3_X1 U7619 ( .A1(n7774), .A2(n6427), .A3(n14362), .ZN(n6654) );
  NAND2_X1 U7620 ( .A1(n6736), .A2(n6734), .ZN(n6427) );
  NAND2_X1 U7621 ( .A1(n7774), .A2(n6427), .ZN(n12092) );
  NAND2_X1 U7622 ( .A1(n6430), .A2(n8145), .ZN(n8166) );
  NAND3_X1 U7623 ( .A1(n7552), .A2(P2_DATAO_REG_3__SCAN_IN), .A3(n6428), .ZN(
        n7340) );
  NAND2_X1 U7624 ( .A1(n8017), .A2(n8013), .ZN(n8913) );
  NAND2_X2 U7625 ( .A1(n6657), .A2(n8493), .ZN(n13948) );
  NAND2_X1 U7626 ( .A1(n8143), .A2(n8142), .ZN(n6430) );
  OR2_X1 U7627 ( .A1(n9637), .A2(P3_IR_REG_3__SCAN_IN), .ZN(n9601) );
  INV_X1 U7628 ( .A(n9637), .ZN(n9640) );
  OAI222_X1 U7629 ( .A1(P3_U3151), .A2(n12201), .B1(n13090), .B2(n12200), .C1(
        n12199), .C2(n13095), .ZN(P3_U3266) );
  AOI21_X1 U7630 ( .B1(n12773), .B2(n6818), .A(n12834), .ZN(n7222) );
  NAND2_X1 U7631 ( .A1(n7653), .A2(n7654), .ZN(n12773) );
  MUX2_X2 U7632 ( .A(P3_REG1_REG_27__SCAN_IN), .B(n13005), .S(n15665), .Z(
        P3_U3486) );
  NOR2_X2 U7633 ( .A1(n13742), .A2(n13722), .ZN(n13725) );
  OR2_X1 U7634 ( .A1(n10015), .A2(n10686), .ZN(n9540) );
  AOI22_X2 U7635 ( .A1(n12693), .A2(n12692), .B1(P3_REG1_REG_16__SCAN_IN), 
        .B2(n12701), .ZN(n12712) );
  NAND3_X2 U7636 ( .A1(n8826), .A2(n7265), .A3(n7263), .ZN(n6434) );
  NAND3_X1 U7637 ( .A1(n8826), .A2(n7265), .A3(n7263), .ZN(n6435) );
  NAND3_X1 U7638 ( .A1(n8826), .A2(n7265), .A3(n7263), .ZN(n9291) );
  OAI21_X1 U7639 ( .B1(n7776), .B2(n14516), .A(n11852), .ZN(n7775) );
  NAND2_X1 U7640 ( .A1(n15293), .A2(n14556), .ZN(n14302) );
  NAND4_X2 U7641 ( .A1(n8943), .A2(n8942), .A3(n8941), .A4(n8940), .ZN(n14556)
         );
  NOR2_X2 U7642 ( .A1(n9491), .A2(n7205), .ZN(n9501) );
  NAND2_X2 U7643 ( .A1(n12402), .A2(n12401), .ZN(n10589) );
  AOI21_X1 U7644 ( .B1(n10962), .B2(n9608), .A(n9607), .ZN(n9610) );
  NOR2_X2 U7645 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8886) );
  INV_X1 U7646 ( .A(n6494), .ZN(n6436) );
  NAND2_X1 U7647 ( .A1(n10106), .A2(n14292), .ZN(n6494) );
  NOR2_X2 U7648 ( .A1(n11556), .A2(n14344), .ZN(n11530) );
  INV_X1 U7649 ( .A(n7554), .ZN(n7455) );
  NAND2_X2 U7650 ( .A1(n11778), .A2(n9764), .ZN(n11765) );
  INV_X1 U7651 ( .A(n9846), .ZN(n6441) );
  INV_X2 U7652 ( .A(n9846), .ZN(n10012) );
  AOI21_X2 U7653 ( .B1(n11134), .B2(n6722), .A(n6593), .ZN(n11480) );
  CLKBUF_X1 U7654 ( .A(n12225), .Z(n6444) );
  NAND2_X1 U7655 ( .A1(n13081), .A2(n13085), .ZN(n6447) );
  NAND2_X1 U7656 ( .A1(n13081), .A2(n13085), .ZN(n6448) );
  OAI21_X2 U7657 ( .B1(n11249), .B2(n7082), .A(n7080), .ZN(n11430) );
  NAND2_X2 U7658 ( .A1(n9677), .A2(n9676), .ZN(n11249) );
  AOI21_X2 U7659 ( .B1(n7055), .B2(n12979), .A(n9534), .ZN(n10964) );
  NOR2_X1 U7660 ( .A1(n9878), .A2(n7079), .ZN(n7078) );
  INV_X1 U7661 ( .A(n9864), .ZN(n7079) );
  INV_X1 U7662 ( .A(n9780), .ZN(n7652) );
  AND2_X1 U7663 ( .A1(n9877), .A2(n9876), .ZN(n12320) );
  NOR2_X1 U7664 ( .A1(n9638), .A2(n10001), .ZN(n7850) );
  INV_X1 U7665 ( .A(n12223), .ZN(n7867) );
  NAND2_X1 U7666 ( .A1(n12372), .A2(n12371), .ZN(n12517) );
  NAND2_X1 U7667 ( .A1(n15545), .A2(n6911), .ZN(n10694) );
  NAND2_X1 U7668 ( .A1(n6905), .A2(n11219), .ZN(n15567) );
  NAND2_X1 U7669 ( .A1(n15545), .A2(n10693), .ZN(n6905) );
  OR2_X1 U7670 ( .A1(n12932), .A2(n12345), .ZN(n12514) );
  NAND2_X1 U7671 ( .A1(n12414), .A2(n10768), .ZN(n9606) );
  NAND2_X1 U7672 ( .A1(n10736), .A2(n7152), .ZN(n10582) );
  NAND2_X1 U7673 ( .A1(n9514), .A2(n10736), .ZN(n12402) );
  OR2_X1 U7674 ( .A1(n12944), .A2(n12821), .ZN(n12497) );
  NOR2_X1 U7675 ( .A1(n13869), .A2(n6954), .ZN(n6953) );
  NAND2_X1 U7676 ( .A1(n10296), .A2(n7875), .ZN(n13495) );
  NOR2_X1 U7677 ( .A1(n14286), .A2(n11494), .ZN(n10245) );
  NAND2_X1 U7678 ( .A1(n8722), .A2(n7164), .ZN(n8733) );
  NAND2_X1 U7679 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n7165), .ZN(n7164) );
  INV_X1 U7680 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n7165) );
  NAND2_X2 U7681 ( .A1(n9504), .A2(n12201), .ZN(n9846) );
  AOI21_X1 U7682 ( .B1(n7831), .B2(n7833), .A(n7828), .ZN(n7827) );
  INV_X1 U7683 ( .A(n12515), .ZN(n7828) );
  INV_X1 U7684 ( .A(n12862), .ZN(n6700) );
  NAND2_X1 U7685 ( .A1(n7075), .A2(n7074), .ZN(n7663) );
  AOI21_X1 U7686 ( .B1(n7076), .B2(n7077), .A(n6560), .ZN(n7074) );
  AND2_X1 U7687 ( .A1(n12893), .A2(n7059), .ZN(n7058) );
  OAI21_X1 U7688 ( .B1(n11765), .B2(n7060), .A(n7061), .ZN(n7056) );
  NAND2_X1 U7689 ( .A1(n7992), .A2(n7993), .ZN(n8398) );
  INV_X1 U7690 ( .A(n8055), .ZN(n8174) );
  NAND2_X1 U7691 ( .A1(n14529), .A2(n14492), .ZN(n14530) );
  OAI21_X1 U7692 ( .B1(n6556), .B2(n7252), .A(n14756), .ZN(n7245) );
  NOR2_X1 U7693 ( .A1(n14861), .A2(n7246), .ZN(n7243) );
  OAI21_X1 U7694 ( .B1(n14866), .B2(n6476), .A(n6589), .ZN(n6762) );
  AND2_X1 U7695 ( .A1(n13303), .A2(n13302), .ZN(n13313) );
  INV_X1 U7696 ( .A(n6851), .ZN(n6850) );
  OAI21_X1 U7697 ( .B1(n6412), .B2(n6853), .A(n6852), .ZN(n6851) );
  NAND2_X1 U7698 ( .A1(n6412), .A2(n14295), .ZN(n6852) );
  AOI22_X1 U7699 ( .A1(n14036), .A2(n13492), .B1(n6440), .B2(n13606), .ZN(
        n13336) );
  AOI21_X1 U7700 ( .B1(n7331), .B2(n7330), .A(n7329), .ZN(n7328) );
  NAND2_X1 U7701 ( .A1(n12429), .A2(n12512), .ZN(n7336) );
  NAND2_X1 U7702 ( .A1(n14351), .A2(n6874), .ZN(n6871) );
  NAND2_X1 U7703 ( .A1(n7531), .A2(n14353), .ZN(n7530) );
  INV_X1 U7704 ( .A(n14354), .ZN(n7531) );
  NAND2_X1 U7705 ( .A1(n6462), .A2(n6554), .ZN(n6872) );
  INV_X1 U7706 ( .A(n13387), .ZN(n7285) );
  INV_X1 U7707 ( .A(n13374), .ZN(n6750) );
  NOR2_X1 U7708 ( .A1(n14407), .A2(n14406), .ZN(n7535) );
  AND2_X1 U7709 ( .A1(n7916), .A2(n7297), .ZN(n7296) );
  INV_X1 U7710 ( .A(n13423), .ZN(n7297) );
  INV_X1 U7711 ( .A(n8288), .ZN(n7941) );
  INV_X1 U7712 ( .A(n14411), .ZN(n7524) );
  INV_X1 U7713 ( .A(n14410), .ZN(n7525) );
  NOR2_X1 U7714 ( .A1(n6912), .A2(n11219), .ZN(n6911) );
  NAND2_X1 U7715 ( .A1(n12612), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7608) );
  INV_X1 U7716 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n9624) );
  OR2_X1 U7717 ( .A1(n13512), .A2(n13510), .ZN(n7162) );
  NOR2_X1 U7718 ( .A1(n7524), .A2(n7525), .ZN(n7523) );
  AND2_X1 U7719 ( .A1(n8107), .A2(n8088), .ZN(n6989) );
  NAND2_X1 U7720 ( .A1(n8707), .A2(n8706), .ZN(n8708) );
  INV_X1 U7721 ( .A(n12268), .ZN(n7863) );
  INV_X1 U7722 ( .A(n12517), .ZN(n12547) );
  NAND2_X1 U7723 ( .A1(n7603), .A2(n6628), .ZN(n7602) );
  AOI21_X1 U7724 ( .B1(n9950), .B2(n7660), .A(n6576), .ZN(n7659) );
  INV_X1 U7725 ( .A(n7956), .ZN(n7660) );
  NAND2_X1 U7726 ( .A1(n7826), .A2(n12457), .ZN(n7823) );
  NAND2_X1 U7727 ( .A1(n7130), .A2(n7144), .ZN(n12418) );
  INV_X1 U7728 ( .A(n12582), .ZN(n7144) );
  NOR2_X1 U7729 ( .A1(n9989), .A2(SI_3_), .ZN(n7135) );
  OR2_X1 U7730 ( .A1(n12249), .A2(n12333), .ZN(n12541) );
  NAND2_X1 U7731 ( .A1(n11826), .A2(n11677), .ZN(n12471) );
  INV_X1 U7732 ( .A(n10025), .ZN(n7851) );
  AOI21_X1 U7733 ( .B1(n7716), .B2(n9852), .A(n7715), .ZN(n7714) );
  INV_X1 U7734 ( .A(n9865), .ZN(n7715) );
  NAND2_X1 U7735 ( .A1(n9658), .A2(n9657), .ZN(n9680) );
  NOR2_X1 U7736 ( .A1(n6782), .A2(n9548), .ZN(n7744) );
  AND2_X1 U7737 ( .A1(n10168), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n9548) );
  INV_X1 U7738 ( .A(n9545), .ZN(n6782) );
  NAND2_X1 U7739 ( .A1(n10170), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n9550) );
  NAND2_X1 U7740 ( .A1(n7354), .A2(n11996), .ZN(n7353) );
  INV_X1 U7741 ( .A(n11995), .ZN(n7354) );
  NAND2_X1 U7742 ( .A1(n7436), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U7743 ( .A1(n15497), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7435) );
  AND2_X1 U7744 ( .A1(n8578), .A2(n8556), .ZN(n6774) );
  NAND2_X1 U7745 ( .A1(n6778), .A2(n8504), .ZN(n13717) );
  NOR2_X1 U7746 ( .A1(n13534), .A2(n7693), .ZN(n7692) );
  INV_X1 U7747 ( .A(n8679), .ZN(n7693) );
  NAND2_X1 U7748 ( .A1(n6686), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8394) );
  INV_X1 U7749 ( .A(n8368), .ZN(n6686) );
  AND2_X1 U7750 ( .A1(n8247), .A2(n6771), .ZN(n6770) );
  NAND2_X1 U7751 ( .A1(n8225), .A2(n6407), .ZN(n6771) );
  OR2_X1 U7752 ( .A1(n8667), .A2(n7683), .ZN(n7685) );
  INV_X1 U7753 ( .A(n8665), .ZN(n7683) );
  NAND2_X1 U7754 ( .A1(n11358), .A2(n8658), .ZN(n8662) );
  AOI21_X1 U7755 ( .B1(n6940), .B2(n7381), .A(n13546), .ZN(n6939) );
  OR2_X1 U7756 ( .A1(n11003), .A2(n6941), .ZN(n6937) );
  INV_X1 U7757 ( .A(n7381), .ZN(n6941) );
  NOR2_X1 U7758 ( .A1(n12144), .A2(n13540), .ZN(n7678) );
  XNOR2_X1 U7759 ( .A(n7395), .B(n13286), .ZN(n10113) );
  OR2_X1 U7760 ( .A1(n9370), .A2(n9369), .ZN(n9404) );
  NAND2_X1 U7761 ( .A1(n9310), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n9333) );
  NAND2_X1 U7762 ( .A1(n9310), .A2(n7278), .ZN(n9352) );
  AND2_X1 U7763 ( .A1(n6735), .A2(n11851), .ZN(n6734) );
  NAND2_X1 U7764 ( .A1(n6508), .A2(n11848), .ZN(n6735) );
  INV_X1 U7765 ( .A(n11409), .ZN(n11481) );
  INV_X1 U7766 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U7767 ( .A1(n8315), .A2(n10780), .ZN(n8358) );
  NAND2_X1 U7768 ( .A1(n8337), .A2(n8336), .ZN(n8359) );
  AND2_X1 U7769 ( .A1(n15782), .A2(P3_ADDR_REG_6__SCAN_IN), .ZN(n6660) );
  AOI21_X1 U7770 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(n8728), .A(n8727), .ZN(
        n8782) );
  NOR2_X1 U7771 ( .A1(n8779), .A2(n8778), .ZN(n8727) );
  NAND2_X1 U7772 ( .A1(n10578), .A2(n12549), .ZN(n10581) );
  XNOR2_X1 U7773 ( .A(n9604), .B(n6444), .ZN(n10649) );
  NAND2_X1 U7774 ( .A1(n6514), .A2(n7870), .ZN(n7869) );
  NOR2_X1 U7775 ( .A1(n11638), .A2(n7872), .ZN(n7871) );
  OR2_X1 U7776 ( .A1(n7116), .A2(n7177), .ZN(n7113) );
  AND2_X1 U7777 ( .A1(n11824), .A2(n7117), .ZN(n7116) );
  NAND2_X1 U7778 ( .A1(n6449), .A2(n7118), .ZN(n7117) );
  NAND2_X1 U7779 ( .A1(n7178), .A2(n6449), .ZN(n7114) );
  NAND2_X1 U7780 ( .A1(n10531), .A2(n10163), .ZN(n10548) );
  NAND2_X1 U7781 ( .A1(n6913), .A2(n6571), .ZN(n7706) );
  AOI21_X1 U7782 ( .B1(n12518), .B2(n12546), .A(n12517), .ZN(n6916) );
  NAND2_X1 U7783 ( .A1(n10624), .A2(n10401), .ZN(n10402) );
  NAND2_X1 U7784 ( .A1(n10402), .A2(n10680), .ZN(n10406) );
  AOI21_X1 U7785 ( .B1(n15543), .B2(n7619), .A(n7618), .ZN(n7616) );
  INV_X1 U7786 ( .A(n15544), .ZN(n7618) );
  NAND2_X1 U7787 ( .A1(n6977), .A2(n6458), .ZN(n6971) );
  OAI21_X1 U7788 ( .B1(n15565), .B2(n6978), .A(n11696), .ZN(n6977) );
  NAND2_X1 U7789 ( .A1(n11693), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n12588) );
  NAND2_X1 U7790 ( .A1(n7605), .A2(n7601), .ZN(n7600) );
  AND2_X1 U7791 ( .A1(n12587), .A2(n12646), .ZN(n7601) );
  INV_X1 U7792 ( .A(n12377), .ZN(n9998) );
  AND2_X1 U7793 ( .A1(n9891), .A2(n9890), .ZN(n12837) );
  AND2_X1 U7794 ( .A1(n12843), .A2(n9892), .ZN(n7662) );
  NOR2_X1 U7795 ( .A1(n10078), .A2(n7825), .ZN(n7824) );
  INV_X1 U7796 ( .A(n12457), .ZN(n7825) );
  AND2_X1 U7797 ( .A1(n12466), .A2(n12471), .ZN(n12538) );
  NOR2_X1 U7798 ( .A1(n9989), .A2(n10143), .ZN(n9497) );
  AOI21_X1 U7799 ( .B1(n12771), .B2(n9991), .A(n9980), .ZN(n12230) );
  NAND2_X1 U7800 ( .A1(n7830), .A2(n7832), .ZN(n12778) );
  AOI21_X1 U7801 ( .B1(n6708), .B2(n6706), .A(n7835), .ZN(n6705) );
  INV_X1 U7802 ( .A(n12982), .ZN(n12836) );
  AOI21_X1 U7803 ( .B1(n7078), .B2(n12872), .A(n6568), .ZN(n7076) );
  AOI21_X1 U7804 ( .B1(n7649), .B2(n7651), .A(n7062), .ZN(n7061) );
  INV_X1 U7805 ( .A(n7430), .ZN(n7429) );
  NAND2_X1 U7806 ( .A1(n11265), .A2(n7838), .ZN(n7428) );
  NAND2_X1 U7807 ( .A1(n10876), .A2(n12512), .ZN(n12838) );
  OR2_X1 U7808 ( .A1(n12560), .A2(n12400), .ZN(n15626) );
  INV_X1 U7809 ( .A(n10548), .ZN(n10543) );
  OAI21_X1 U7810 ( .B1(n11934), .B2(n11933), .A(n11935), .ZN(n12354) );
  AOI21_X1 U7811 ( .B1(n7758), .B2(n7747), .A(n7745), .ZN(n9940) );
  NOR2_X1 U7812 ( .A1(n7752), .A2(n7748), .ZN(n7747) );
  NOR2_X1 U7813 ( .A1(n7749), .A2(n7746), .ZN(n7745) );
  OR2_X1 U7814 ( .A1(n9895), .A2(n9894), .ZN(n7756) );
  NAND2_X1 U7815 ( .A1(n9837), .A2(n9836), .ZN(n9853) );
  AOI21_X1 U7816 ( .B1(n7729), .B2(n7730), .A(n6797), .ZN(n6796) );
  INV_X1 U7817 ( .A(n9800), .ZN(n6797) );
  INV_X1 U7818 ( .A(n7731), .ZN(n7730) );
  NAND2_X1 U7819 ( .A1(n10179), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U7820 ( .A1(n11997), .A2(n11996), .ZN(n13111) );
  INV_X1 U7821 ( .A(n7011), .ZN(n7009) );
  AOI21_X1 U7822 ( .B1(n7011), .B2(n7008), .A(n6575), .ZN(n7007) );
  INV_X1 U7823 ( .A(n13162), .ZN(n7008) );
  NAND2_X1 U7824 ( .A1(n7497), .A2(n13099), .ZN(n7014) );
  AND2_X1 U7825 ( .A1(n7495), .A2(n6616), .ZN(n7494) );
  AND3_X1 U7826 ( .A1(n10562), .A2(n10561), .A3(n10560), .ZN(n10567) );
  INV_X1 U7827 ( .A(n13284), .ZN(n13580) );
  AND2_X1 U7828 ( .A1(n8437), .A2(n8436), .ZN(n13430) );
  AND2_X1 U7829 ( .A1(n8401), .A2(n8400), .ZN(n13203) );
  AND4_X1 U7830 ( .A1(n8100), .A2(n8099), .A3(n8098), .A4(n8097), .ZN(n13330)
         );
  INV_X1 U7831 ( .A(n7993), .ZN(n7994) );
  AOI21_X1 U7832 ( .B1(n15409), .B2(n7450), .A(n6578), .ZN(n7449) );
  INV_X1 U7833 ( .A(n10367), .ZN(n7450) );
  OR2_X1 U7834 ( .A1(n15494), .A2(n15493), .ZN(n7436) );
  INV_X1 U7835 ( .A(n7391), .ZN(n7390) );
  NAND2_X1 U7836 ( .A1(n6958), .A2(n13889), .ZN(n6951) );
  AND2_X1 U7837 ( .A1(n10563), .A2(n10307), .ZN(n13880) );
  NAND2_X1 U7838 ( .A1(n8152), .A2(n8151), .ZN(n14031) );
  AOI21_X1 U7839 ( .B1(n8628), .B2(n11490), .A(n11624), .ZN(n15502) );
  XNOR2_X1 U7840 ( .A(n8635), .B(n8634), .ZN(n11449) );
  XNOR2_X1 U7841 ( .A(n7036), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U7842 ( .A1(n14091), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7036) );
  INV_X1 U7843 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U7844 ( .A1(n8618), .A2(n8617), .ZN(n8620) );
  INV_X1 U7845 ( .A(n8616), .ZN(n8618) );
  AND2_X1 U7846 ( .A1(n7998), .A2(n7977), .ZN(n7698) );
  NOR2_X1 U7847 ( .A1(n14160), .A2(n7575), .ZN(n7574) );
  INV_X1 U7848 ( .A(n9270), .ZN(n7575) );
  AND2_X1 U7849 ( .A1(n14446), .A2(n14443), .ZN(n14444) );
  NAND2_X1 U7851 ( .A1(n14478), .A2(n14477), .ZN(n14743) );
  OR2_X1 U7852 ( .A1(n14095), .A2(n12036), .ZN(n12038) );
  NOR2_X1 U7853 ( .A1(n14780), .A2(n7549), .ZN(n7548) );
  INV_X1 U7854 ( .A(n7550), .ZN(n7549) );
  NOR2_X1 U7855 ( .A1(n7794), .A2(n7792), .ZN(n7791) );
  NAND2_X1 U7856 ( .A1(n7790), .A2(n14797), .ZN(n7788) );
  XNOR2_X1 U7857 ( .A(n14750), .B(n14806), .ZN(n14797) );
  NAND2_X1 U7858 ( .A1(n14796), .A2(n12106), .ZN(n14755) );
  NAND2_X1 U7859 ( .A1(n11562), .A2(n8962), .ZN(n9331) );
  INV_X1 U7860 ( .A(n12097), .ZN(n7804) );
  NAND2_X1 U7861 ( .A1(n7803), .A2(n14402), .ZN(n7802) );
  NAND2_X1 U7862 ( .A1(n15042), .A2(n15327), .ZN(n7271) );
  NAND2_X1 U7863 ( .A1(n8858), .A2(n9443), .ZN(n14286) );
  MUX2_X1 U7864 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8854), .S(
        P1_IR_REG_22__SCAN_IN), .Z(n8858) );
  AND2_X1 U7865 ( .A1(n8724), .A2(P3_ADDR_REG_12__SCAN_IN), .ZN(n6661) );
  NOR2_X1 U7866 ( .A1(n8733), .A2(n8734), .ZN(n8723) );
  NAND3_X1 U7867 ( .A1(n6819), .A2(n6820), .A3(n6532), .ZN(n8774) );
  AND2_X1 U7868 ( .A1(n15230), .A2(n7313), .ZN(n7312) );
  NAND2_X1 U7869 ( .A1(n9958), .A2(n9957), .ZN(n12932) );
  AOI21_X1 U7870 ( .B1(n7099), .B2(n7097), .A(n6637), .ZN(n7096) );
  AND2_X1 U7871 ( .A1(n10878), .A2(n12512), .ZN(n12982) );
  NAND2_X1 U7872 ( .A1(n9863), .A2(n9862), .ZN(n12887) );
  NAND2_X1 U7873 ( .A1(n10625), .A2(n10626), .ZN(n10624) );
  NAND2_X1 U7874 ( .A1(n13123), .A2(n11987), .ZN(n13206) );
  NAND2_X1 U7875 ( .A1(n13230), .A2(n7217), .ZN(n6934) );
  AOI21_X1 U7876 ( .B1(n8697), .B2(n13919), .A(n8693), .ZN(n8694) );
  AOI21_X1 U7877 ( .B1(n7568), .B2(n7570), .A(n6564), .ZN(n7566) );
  AOI21_X1 U7878 ( .B1(n14736), .B2(n14737), .A(n6490), .ZN(n6692) );
  NAND2_X1 U7879 ( .A1(n15239), .A2(n15472), .ZN(n15236) );
  NAND2_X1 U7880 ( .A1(n6656), .A2(n6655), .ZN(n15238) );
  INV_X1 U7881 ( .A(n8783), .ZN(n6655) );
  INV_X1 U7882 ( .A(n8784), .ZN(n6656) );
  NAND2_X1 U7883 ( .A1(n12398), .A2(n12397), .ZN(n7330) );
  NAND2_X1 U7884 ( .A1(n12396), .A2(n12400), .ZN(n12395) );
  AOI21_X1 U7885 ( .B1(n13321), .B2(n13322), .A(n6529), .ZN(n6718) );
  OR2_X1 U7886 ( .A1(n13316), .A2(n13317), .ZN(n6720) );
  NAND2_X1 U7887 ( .A1(n13314), .A2(n13315), .ZN(n6715) );
  INV_X1 U7888 ( .A(n6590), .ZN(n7908) );
  INV_X1 U7889 ( .A(n13331), .ZN(n7907) );
  NAND2_X1 U7890 ( .A1(n6849), .A2(n14297), .ZN(n14305) );
  OAI21_X1 U7891 ( .B1(n15251), .B2(n14296), .A(n6850), .ZN(n6849) );
  NAND2_X1 U7892 ( .A1(n13344), .A2(n6475), .ZN(n6732) );
  NAND2_X1 U7893 ( .A1(n6847), .A2(n6547), .ZN(n6846) );
  INV_X1 U7894 ( .A(n14308), .ZN(n6847) );
  INV_X1 U7895 ( .A(n14311), .ZN(n7538) );
  INV_X1 U7896 ( .A(n6732), .ZN(n6727) );
  NAND2_X1 U7897 ( .A1(n13339), .A2(n6733), .ZN(n6729) );
  NOR2_X1 U7898 ( .A1(n13344), .A2(n6475), .ZN(n7903) );
  AOI21_X1 U7899 ( .B1(n12430), .B2(n12513), .A(n7209), .ZN(n7337) );
  NAND2_X1 U7900 ( .A1(n12433), .A2(n12530), .ZN(n7335) );
  OR2_X1 U7901 ( .A1(n6522), .A2(n7291), .ZN(n7289) );
  NAND2_X1 U7902 ( .A1(n6522), .A2(n7291), .ZN(n7290) );
  NAND2_X1 U7903 ( .A1(n6872), .A2(n6871), .ZN(n14355) );
  AND2_X1 U7904 ( .A1(n7533), .A2(n14354), .ZN(n7532) );
  INV_X1 U7905 ( .A(n14353), .ZN(n7533) );
  AOI21_X1 U7906 ( .B1(n12472), .B2(n12471), .A(n12513), .ZN(n12474) );
  AOI21_X1 U7907 ( .B1(n7321), .B2(n7322), .A(n7320), .ZN(n7319) );
  AND2_X1 U7908 ( .A1(n12469), .A2(n7325), .ZN(n7322) );
  INV_X1 U7909 ( .A(n12474), .ZN(n7321) );
  OAI22_X1 U7910 ( .A1(n12474), .A2(n12472), .B1(n12473), .B2(n13062), .ZN(
        n7320) );
  OAI21_X1 U7911 ( .B1(n14358), .B2(n14359), .A(n14360), .ZN(n14366) );
  NAND2_X1 U7912 ( .A1(n7526), .A2(n7530), .ZN(n14359) );
  NAND2_X1 U7913 ( .A1(n6872), .A2(n6870), .ZN(n7526) );
  NAND2_X1 U7914 ( .A1(n14366), .A2(n14367), .ZN(n14365) );
  NAND2_X1 U7915 ( .A1(n6577), .A2(n13393), .ZN(n7910) );
  NOR2_X1 U7916 ( .A1(n6567), .A2(n7282), .ZN(n7281) );
  NAND2_X1 U7917 ( .A1(n6818), .A2(n12544), .ZN(n6817) );
  NOR3_X1 U7918 ( .A1(n6786), .A2(n12893), .A3(n12909), .ZN(n6785) );
  OR2_X1 U7919 ( .A1(n12506), .A2(n12512), .ZN(n7315) );
  NAND2_X1 U7920 ( .A1(n12509), .A2(n12512), .ZN(n7317) );
  OR2_X1 U7921 ( .A1(n13008), .A2(n12566), .ZN(n9950) );
  AOI21_X1 U7922 ( .B1(n13456), .B2(n6440), .A(n13455), .ZN(n13512) );
  NAND2_X1 U7923 ( .A1(n7915), .A2(n13423), .ZN(n7914) );
  INV_X1 U7924 ( .A(n7919), .ZN(n7915) );
  NOR2_X1 U7925 ( .A1(n7293), .A2(n6452), .ZN(n6758) );
  NAND2_X1 U7926 ( .A1(n6595), .A2(n6480), .ZN(n7293) );
  AND2_X1 U7927 ( .A1(n7912), .A2(n13422), .ZN(n7911) );
  NAND2_X1 U7928 ( .A1(n7913), .A2(n13423), .ZN(n7912) );
  AND2_X1 U7929 ( .A1(n7296), .A2(n6617), .ZN(n7295) );
  NAND2_X1 U7930 ( .A1(n13781), .A2(n13817), .ZN(n6678) );
  OR4_X1 U7931 ( .A1(n13554), .A2(n6407), .A3(n13553), .A4(n13907), .ZN(n13555) );
  INV_X1 U7932 ( .A(n8504), .ZN(n6781) );
  OAI21_X1 U7933 ( .B1(n11808), .B2(n7927), .A(n8272), .ZN(n7926) );
  AOI21_X1 U7934 ( .B1(n7939), .B2(n13889), .A(n8335), .ZN(n7938) );
  NAND2_X1 U7935 ( .A1(n8376), .A2(n8377), .ZN(n7937) );
  NOR2_X1 U7936 ( .A1(n7937), .A2(n7940), .ZN(n7936) );
  NOR4_X1 U7937 ( .A1(n14755), .A2(n14520), .A3(n14887), .A4(n14869), .ZN(
        n14521) );
  NOR2_X1 U7938 ( .A1(n7519), .A2(n14412), .ZN(n7518) );
  INV_X1 U7939 ( .A(n7522), .ZN(n7519) );
  NAND2_X1 U7940 ( .A1(n6597), .A2(n14408), .ZN(n6867) );
  NAND2_X1 U7941 ( .A1(n7514), .A2(n7513), .ZN(n7512) );
  NAND2_X1 U7942 ( .A1(n7522), .A2(n14413), .ZN(n7513) );
  INV_X1 U7943 ( .A(n7518), .ZN(n7514) );
  OR2_X1 U7944 ( .A1(n7520), .A2(n7517), .ZN(n7516) );
  AOI21_X1 U7945 ( .B1(n7523), .B2(n7522), .A(n7521), .ZN(n7520) );
  NOR2_X1 U7946 ( .A1(n7259), .A2(n7255), .ZN(n7254) );
  INV_X1 U7947 ( .A(n7261), .ZN(n7255) );
  NOR2_X1 U7948 ( .A1(n7888), .A2(n8559), .ZN(n7887) );
  INV_X1 U7949 ( .A(n7890), .ZN(n7888) );
  INV_X1 U7950 ( .A(n7891), .ZN(n7885) );
  AOI21_X1 U7951 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8414) );
  NAND2_X1 U7952 ( .A1(n8067), .A2(n8069), .ZN(n7541) );
  INV_X1 U7953 ( .A(n9626), .ZN(n9625) );
  INV_X1 U7954 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n6929) );
  NOR2_X1 U7955 ( .A1(n12213), .A2(n7103), .ZN(n7102) );
  INV_X1 U7956 ( .A(n7109), .ZN(n7103) );
  INV_X1 U7957 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n10023) );
  INV_X1 U7958 ( .A(n10528), .ZN(n10410) );
  NAND2_X1 U7959 ( .A1(n10627), .A2(n10413), .ZN(n10415) );
  NAND2_X1 U7960 ( .A1(n6650), .A2(n15567), .ZN(n15569) );
  NOR2_X1 U7961 ( .A1(n15588), .A2(n6904), .ZN(n11692) );
  NOR2_X1 U7962 ( .A1(n15597), .A2(n11691), .ZN(n6904) );
  OAI21_X1 U7963 ( .B1(n6896), .B2(n6900), .A(n6902), .ZN(n7592) );
  INV_X1 U7964 ( .A(n6897), .ZN(n6902) );
  NAND2_X1 U7965 ( .A1(n7599), .A2(n6623), .ZN(n6900) );
  NAND2_X1 U7966 ( .A1(n12660), .A2(n12659), .ZN(n12684) );
  INV_X1 U7967 ( .A(n12351), .ZN(n12519) );
  INV_X1 U7968 ( .A(n6919), .ZN(n6917) );
  NOR2_X1 U7969 ( .A1(n9857), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n7225) );
  NOR2_X1 U7970 ( .A1(n9793), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n7226) );
  INV_X1 U7971 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n9741) );
  INV_X1 U7972 ( .A(n9743), .ZN(n9742) );
  AND2_X1 U7973 ( .A1(n9741), .A2(n6927), .ZN(n6926) );
  INV_X1 U7974 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n6927) );
  NAND2_X1 U7975 ( .A1(n9625), .A2(n9624), .ZN(n9646) );
  NAND2_X1 U7976 ( .A1(n12583), .A2(n12990), .ZN(n12404) );
  INV_X1 U7977 ( .A(n12820), .ZN(n12544) );
  INV_X1 U7978 ( .A(n9693), .ZN(n7084) );
  NOR2_X1 U7979 ( .A1(n10961), .A2(n12529), .ZN(n11090) );
  INV_X1 U7980 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n9487) );
  INV_X1 U7981 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n9486) );
  INV_X1 U7982 ( .A(n7703), .ZN(n7702) );
  OAI21_X1 U7983 ( .B1(n9953), .B2(n7704), .A(n9971), .ZN(n7703) );
  INV_X1 U7984 ( .A(n9955), .ZN(n7704) );
  INV_X1 U7985 ( .A(n7724), .ZN(n7719) );
  NOR2_X1 U7986 ( .A1(n9611), .A2(n7725), .ZN(n7724) );
  INV_X1 U7987 ( .A(n9552), .ZN(n7725) );
  NAND2_X1 U7988 ( .A1(n10196), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n9634) );
  INV_X1 U7989 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6890) );
  NAND2_X1 U7990 ( .A1(n10709), .A2(n13238), .ZN(n7487) );
  NAND2_X1 U7991 ( .A1(n10555), .A2(n6409), .ZN(n10710) );
  NAND2_X1 U7992 ( .A1(n13231), .A2(n13232), .ZN(n7486) );
  NAND2_X1 U7993 ( .A1(n10710), .A2(n10711), .ZN(n10709) );
  XNOR2_X1 U7994 ( .A(n10717), .B(n6751), .ZN(n13231) );
  NAND2_X1 U7995 ( .A1(n6460), .A2(n8680), .ZN(n6943) );
  AND2_X1 U7996 ( .A1(n13538), .A2(n7934), .ZN(n7933) );
  OR2_X1 U7997 ( .A1(n13718), .A2(n7935), .ZN(n7934) );
  INV_X1 U7998 ( .A(n8525), .ZN(n7935) );
  INV_X1 U7999 ( .A(n13537), .ZN(n7932) );
  INV_X1 U8000 ( .A(n6780), .ZN(n6779) );
  OAI21_X1 U8001 ( .B1(n7922), .B2(n6781), .A(n7933), .ZN(n6780) );
  NAND2_X1 U8002 ( .A1(n6779), .A2(n6781), .ZN(n6777) );
  OR2_X1 U8003 ( .A1(n14058), .A2(n13426), .ZN(n8463) );
  NAND2_X1 U8004 ( .A1(n13791), .A2(n6879), .ZN(n7769) );
  INV_X1 U8005 ( .A(n8366), .ZN(n8349) );
  NOR2_X1 U8006 ( .A1(n13866), .A2(n14009), .ZN(n7759) );
  AND2_X1 U8007 ( .A1(n6518), .A2(n8162), .ZN(n7024) );
  NAND2_X1 U8008 ( .A1(n6888), .A2(n7013), .ZN(n6886) );
  NAND2_X1 U8009 ( .A1(n8651), .A2(n13916), .ZN(n8032) );
  NAND2_X1 U8010 ( .A1(n13304), .A2(n6751), .ZN(n8051) );
  OR2_X1 U8011 ( .A1(n13460), .A2(n13456), .ZN(n7773) );
  AND2_X1 U8012 ( .A1(n13725), .A2(n13712), .ZN(n13707) );
  OR2_X1 U8013 ( .A1(n13754), .A2(n13948), .ZN(n13742) );
  NOR2_X1 U8014 ( .A1(n13820), .A2(n7769), .ZN(n13787) );
  AND2_X1 U8015 ( .A1(n10106), .A2(n10808), .ZN(n8888) );
  INV_X1 U8016 ( .A(n8888), .ZN(n9301) );
  OAI21_X1 U8017 ( .B1(n11148), .B2(n11077), .A(n11076), .ZN(n8975) );
  INV_X1 U8018 ( .A(n9125), .ZN(n8863) );
  INV_X1 U8019 ( .A(n9301), .ZN(n9401) );
  NOR2_X1 U8020 ( .A1(n7796), .A2(n7795), .ZN(n7794) );
  OAI22_X1 U8021 ( .A1(n14830), .A2(n7249), .B1(n14542), .B2(n14840), .ZN(
        n7248) );
  NAND2_X1 U8022 ( .A1(n12137), .A2(n12136), .ZN(n7249) );
  NOR2_X1 U8023 ( .A1(n7277), .A2(n7276), .ZN(n7275) );
  INV_X1 U8024 ( .A(n9232), .ZN(n9231) );
  NOR2_X1 U8025 ( .A1(n14382), .A2(n7262), .ZN(n7261) );
  INV_X1 U8026 ( .A(n12127), .ZN(n7262) );
  INV_X1 U8027 ( .A(n9024), .ZN(n7272) );
  INV_X1 U8028 ( .A(n11133), .ZN(n6723) );
  INV_X1 U8029 ( .A(n14292), .ZN(n10808) );
  NAND2_X1 U8030 ( .A1(n14362), .A2(n7242), .ZN(n7241) );
  INV_X1 U8031 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15756) );
  INV_X1 U8032 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n8856) );
  INV_X1 U8033 ( .A(n7897), .ZN(n7896) );
  AOI21_X1 U8034 ( .B1(n7897), .B2(n7895), .A(n7894), .ZN(n7893) );
  INV_X1 U8035 ( .A(n13445), .ZN(n7894) );
  INV_X1 U8036 ( .A(n12028), .ZN(n7895) );
  INV_X1 U8037 ( .A(n8565), .ZN(n7127) );
  NAND2_X1 U8038 ( .A1(n8543), .A2(n13091), .ZN(n7890) );
  NAND2_X1 U8039 ( .A1(n7892), .A2(SI_26_), .ZN(n7891) );
  INV_X1 U8040 ( .A(n8543), .ZN(n7892) );
  NOR2_X1 U8041 ( .A1(n8443), .A2(n8442), .ZN(n8470) );
  INV_X1 U8042 ( .A(n7509), .ZN(n7508) );
  AND2_X1 U8043 ( .A1(n8358), .A2(n8317), .ZN(n8336) );
  NAND2_X1 U8044 ( .A1(n7635), .A2(n7633), .ZN(n8705) );
  NAND2_X1 U8045 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n7634), .ZN(n7633) );
  INV_X1 U8046 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n7634) );
  XNOR2_X1 U8047 ( .A(n8708), .B(n15756), .ZN(n8749) );
  NAND2_X1 U8048 ( .A1(n15215), .A2(n7632), .ZN(n6834) );
  AND2_X1 U8049 ( .A1(n7107), .A2(n7106), .ZN(n7105) );
  NAND2_X1 U8050 ( .A1(n12212), .A2(n12328), .ZN(n7106) );
  OR2_X1 U8051 ( .A1(n12213), .A2(n7108), .ZN(n7107) );
  NAND2_X1 U8052 ( .A1(n12287), .A2(n7109), .ZN(n7108) );
  NAND2_X1 U8053 ( .A1(n12288), .A2(n7102), .ZN(n7101) );
  AND2_X1 U8054 ( .A1(n7867), .A2(n7966), .ZN(n7866) );
  NAND2_X1 U8055 ( .A1(n6596), .A2(n7867), .ZN(n7865) );
  AND2_X1 U8056 ( .A1(n10653), .A2(n10980), .ZN(n10857) );
  INV_X1 U8057 ( .A(n12584), .ZN(n7807) );
  INV_X1 U8058 ( .A(n12261), .ZN(n7856) );
  AOI21_X1 U8059 ( .B1(n7113), .B2(n7114), .A(n7111), .ZN(n7110) );
  INV_X1 U8060 ( .A(n11827), .ZN(n7111) );
  XNOR2_X1 U8061 ( .A(n6811), .B(n12548), .ZN(n12550) );
  NAND2_X1 U8062 ( .A1(n6812), .A2(n12547), .ZN(n6811) );
  NOR2_X1 U8063 ( .A1(n6814), .A2(n6813), .ZN(n6812) );
  NAND2_X1 U8064 ( .A1(n7706), .A2(n12521), .ZN(n7705) );
  AND2_X1 U8065 ( .A1(n12366), .A2(n12365), .ZN(n12755) );
  NAND2_X1 U8066 ( .A1(n13097), .A2(n10049), .ZN(n10531) );
  AND3_X1 U8067 ( .A1(n9779), .A2(n9778), .A3(n9777), .ZN(n11677) );
  OR2_X1 U8068 ( .A1(n10015), .A2(n15657), .ZN(n9581) );
  OR2_X1 U8069 ( .A1(n10015), .A2(n10390), .ZN(n9594) );
  AOI21_X1 U8070 ( .B1(n10410), .B2(n10409), .A(n10411), .ZN(n10522) );
  AND2_X1 U8071 ( .A1(n10617), .A2(n7373), .ZN(n10516) );
  NAND2_X1 U8072 ( .A1(n10528), .A2(n7374), .ZN(n7373) );
  INV_X1 U8073 ( .A(n10383), .ZN(n7374) );
  INV_X1 U8074 ( .A(n10406), .ZN(n7598) );
  NAND2_X1 U8075 ( .A1(n10406), .A2(n7597), .ZN(n7593) );
  NAND2_X1 U8076 ( .A1(n7614), .A2(n15566), .ZN(n15572) );
  NOR2_X1 U8077 ( .A1(n11219), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6910) );
  INV_X1 U8078 ( .A(n6907), .ZN(n6906) );
  NAND2_X1 U8079 ( .A1(n11241), .A2(n11694), .ZN(n15583) );
  INV_X1 U8080 ( .A(n15564), .ZN(n6974) );
  NOR2_X1 U8081 ( .A1(n7143), .A2(n12585), .ZN(n11693) );
  AND2_X1 U8082 ( .A1(n11692), .A2(n12600), .ZN(n7143) );
  INV_X1 U8083 ( .A(n12586), .ZN(n12585) );
  OR2_X1 U8084 ( .A1(n11692), .A2(n12600), .ZN(n12586) );
  NAND2_X1 U8085 ( .A1(n6967), .A2(n6968), .ZN(n12602) );
  AOI21_X1 U8086 ( .B1(n6969), .B2(n6975), .A(n6591), .ZN(n6968) );
  NAND2_X1 U8087 ( .A1(n7602), .A2(n6903), .ZN(n12630) );
  NAND2_X1 U8088 ( .A1(n6468), .A2(n6625), .ZN(n12632) );
  NOR2_X1 U8089 ( .A1(n6983), .A2(n12619), .ZN(n6982) );
  INV_X1 U8090 ( .A(n6985), .ZN(n6983) );
  INV_X1 U8091 ( .A(n12603), .ZN(n6980) );
  OAI21_X1 U8092 ( .B1(n12640), .B2(n7041), .A(n7039), .ZN(n12673) );
  INV_X1 U8093 ( .A(n7040), .ZN(n7039) );
  OAI21_X1 U8094 ( .B1(n12639), .B2(n7041), .A(n12658), .ZN(n7040) );
  INV_X1 U8095 ( .A(n12653), .ZN(n7041) );
  AND2_X1 U8096 ( .A1(n7592), .A2(n12683), .ZN(n12677) );
  OR2_X1 U8097 ( .A1(n12685), .A2(n12686), .ZN(n7367) );
  OR2_X1 U8098 ( .A1(n12713), .A2(n15723), .ZN(n7050) );
  XNOR2_X1 U8099 ( .A(n12736), .B(n6986), .ZN(n12726) );
  NOR2_X1 U8100 ( .A1(n7049), .A2(n7047), .ZN(n7046) );
  INV_X1 U8101 ( .A(n12747), .ZN(n7047) );
  OR2_X1 U8102 ( .A1(n9976), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n12756) );
  OR2_X1 U8103 ( .A1(n9945), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9961) );
  NAND2_X1 U8104 ( .A1(n6592), .A2(n6467), .ZN(n7420) );
  NAND2_X1 U8105 ( .A1(n12490), .A2(n7423), .ZN(n7422) );
  INV_X1 U8106 ( .A(n12491), .ZN(n7423) );
  NAND2_X1 U8107 ( .A1(n6710), .A2(n7818), .ZN(n11767) );
  AND2_X1 U8108 ( .A1(n12538), .A2(n7819), .ZN(n7818) );
  NAND2_X1 U8109 ( .A1(n7821), .A2(n7820), .ZN(n7819) );
  OAI21_X1 U8110 ( .B1(n12414), .B2(n12408), .A(n12418), .ZN(n7415) );
  NAND2_X1 U8111 ( .A1(n12977), .A2(n10074), .ZN(n10075) );
  INV_X1 U8112 ( .A(n12979), .ZN(n10074) );
  NAND2_X1 U8113 ( .A1(n9515), .A2(n10582), .ZN(n7055) );
  AOI21_X1 U8114 ( .B1(n12198), .B2(n9956), .A(n9990), .ZN(n12387) );
  INV_X1 U8115 ( .A(n7655), .ZN(n7654) );
  OAI21_X1 U8116 ( .B1(n12779), .B2(n7656), .A(n9969), .ZN(n7655) );
  NAND2_X1 U8117 ( .A1(n12809), .A2(n7956), .ZN(n12794) );
  OR2_X1 U8118 ( .A1(n12817), .A2(n12820), .ZN(n12815) );
  AND2_X1 U8119 ( .A1(n9910), .A2(n9909), .ZN(n12821) );
  INV_X1 U8120 ( .A(n7078), .ZN(n7077) );
  AND2_X1 U8121 ( .A1(n6467), .A2(n12389), .ZN(n12852) );
  AOI21_X1 U8122 ( .B1(n6697), .B2(n12539), .A(n6695), .ZN(n6694) );
  NAND2_X1 U8123 ( .A1(n12900), .A2(n6697), .ZN(n6696) );
  INV_X1 U8124 ( .A(n7810), .ZN(n6695) );
  AND2_X1 U8125 ( .A1(n12540), .A2(n9831), .ZN(n7670) );
  NAND2_X1 U8126 ( .A1(n12877), .A2(n12876), .ZN(n12875) );
  AND2_X1 U8127 ( .A1(n12482), .A2(n12390), .ZN(n7816) );
  AND2_X1 U8128 ( .A1(n6528), .A2(n12872), .ZN(n7814) );
  INV_X1 U8129 ( .A(n6584), .ZN(n7059) );
  OR2_X1 U8130 ( .A1(n12900), .A2(n12539), .ZN(n6702) );
  INV_X1 U8131 ( .A(n7651), .ZN(n7650) );
  OAI21_X1 U8132 ( .B1(n11764), .B2(n7652), .A(n9797), .ZN(n7651) );
  NOR2_X1 U8133 ( .A1(n12465), .A2(n12470), .ZN(n12914) );
  NAND2_X1 U8134 ( .A1(n11764), .A2(n11765), .ZN(n11763) );
  NAND2_X1 U8135 ( .A1(n9774), .A2(n9773), .ZN(n11826) );
  INV_X1 U8136 ( .A(n6509), .ZN(n7826) );
  NAND2_X1 U8137 ( .A1(n11435), .A2(n12454), .ZN(n11591) );
  INV_X1 U8138 ( .A(n7846), .ZN(n7840) );
  INV_X1 U8139 ( .A(n12448), .ZN(n7839) );
  INV_X1 U8140 ( .A(n12533), .ZN(n7842) );
  NOR2_X1 U8141 ( .A1(n12534), .A2(n7847), .ZN(n7846) );
  INV_X1 U8142 ( .A(n12439), .ZN(n7847) );
  INV_X1 U8143 ( .A(n7845), .ZN(n7844) );
  OAI21_X1 U8144 ( .B1(n12534), .B2(n6461), .A(n12442), .ZN(n7845) );
  INV_X1 U8145 ( .A(n15626), .ZN(n12933) );
  OR2_X1 U8146 ( .A1(n12513), .A2(n12522), .ZN(n10535) );
  AND2_X1 U8147 ( .A1(n13096), .A2(n10035), .ZN(n7090) );
  NAND2_X1 U8148 ( .A1(n10052), .A2(n7958), .ZN(n7091) );
  NAND2_X1 U8149 ( .A1(n9987), .A2(n9986), .ZN(n11934) );
  INV_X1 U8150 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n9502) );
  NAND2_X1 U8151 ( .A1(n9942), .A2(n9941), .ZN(n9954) );
  NAND2_X1 U8152 ( .A1(n9940), .A2(n9939), .ZN(n9942) );
  NOR2_X1 U8153 ( .A1(n7125), .A2(n7124), .ZN(n7123) );
  NOR2_X1 U8154 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7124) );
  AOI21_X1 U8155 ( .B1(n9899), .B2(n7751), .A(n7755), .ZN(n7753) );
  AOI21_X1 U8156 ( .B1(n6487), .B2(n7713), .A(n6649), .ZN(n6784) );
  AOI21_X1 U8157 ( .B1(n7714), .B2(n7712), .A(n7711), .ZN(n7710) );
  INV_X1 U8158 ( .A(n9867), .ZN(n7711) );
  INV_X1 U8159 ( .A(n9852), .ZN(n7712) );
  AND2_X1 U8160 ( .A1(n9867), .A2(n9854), .ZN(n9865) );
  INV_X1 U8161 ( .A(n9851), .ZN(n7716) );
  NAND2_X1 U8162 ( .A1(n6791), .A2(n6790), .ZN(n9834) );
  AOI21_X1 U8163 ( .B1(n6793), .B2(n6795), .A(n6635), .ZN(n6790) );
  NAND2_X1 U8164 ( .A1(n9766), .A2(n6793), .ZN(n6791) );
  AOI21_X1 U8165 ( .B1(n7731), .B2(n7733), .A(n9798), .ZN(n7729) );
  AOI21_X1 U8166 ( .B1(n7734), .B2(n9765), .A(n7732), .ZN(n7731) );
  INV_X1 U8167 ( .A(n9782), .ZN(n7732) );
  AND2_X1 U8168 ( .A1(n9782), .A2(n9768), .ZN(n9781) );
  XNOR2_X1 U8169 ( .A(n9752), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n9750) );
  NAND2_X1 U8170 ( .A1(n6799), .A2(n6798), .ZN(n9731) );
  AOI21_X1 U8171 ( .B1(n6801), .B2(n6802), .A(n6586), .ZN(n6798) );
  NAND2_X1 U8172 ( .A1(n9680), .A2(n6801), .ZN(n6799) );
  INV_X1 U8173 ( .A(n9678), .ZN(n6807) );
  AOI21_X1 U8174 ( .B1(n9679), .B2(n6806), .A(n6804), .ZN(n6803) );
  INV_X1 U8175 ( .A(n9694), .ZN(n6804) );
  INV_X1 U8176 ( .A(n9680), .ZN(n6809) );
  AND2_X1 U8177 ( .A1(n7722), .A2(n7726), .ZN(n7721) );
  INV_X1 U8178 ( .A(n9614), .ZN(n7722) );
  NAND2_X1 U8179 ( .A1(n9568), .A2(n7724), .ZN(n7723) );
  NAND2_X1 U8180 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n7727), .ZN(n7726) );
  INV_X1 U8181 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n7727) );
  OAI21_X1 U8182 ( .B1(n9546), .B2(n7741), .A(n7738), .ZN(n9570) );
  AOI21_X1 U8183 ( .B1(n7740), .B2(n7742), .A(n7739), .ZN(n7738) );
  INV_X1 U8184 ( .A(n9550), .ZN(n7739) );
  AND2_X1 U8185 ( .A1(n9552), .A2(n9551), .ZN(n9569) );
  NAND2_X1 U8186 ( .A1(n9546), .A2(n7744), .ZN(n7743) );
  NAND2_X1 U8187 ( .A1(n10166), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n9545) );
  NAND2_X1 U8188 ( .A1(n13099), .A2(n11968), .ZN(n13104) );
  NAND2_X1 U8189 ( .A1(n11044), .A2(n6838), .ZN(n6837) );
  NAND2_X1 U8190 ( .A1(n6838), .A2(n11043), .ZN(n6836) );
  NOR2_X1 U8191 ( .A1(n11977), .A2(n7496), .ZN(n7501) );
  INV_X1 U8192 ( .A(n13180), .ZN(n7482) );
  NAND2_X1 U8193 ( .A1(n7017), .A2(n6549), .ZN(n7016) );
  OAI22_X1 U8194 ( .A1(n13154), .A2(n6456), .B1(n6450), .B2(n7348), .ZN(n7017)
         );
  NAND2_X1 U8195 ( .A1(n13153), .A2(n6450), .ZN(n7347) );
  NAND2_X1 U8196 ( .A1(n11999), .A2(n11998), .ZN(n12002) );
  AND2_X1 U8197 ( .A1(n12000), .A2(n13115), .ZN(n7184) );
  XNOR2_X1 U8198 ( .A(n10720), .B(n10719), .ZN(n13190) );
  NAND2_X1 U8199 ( .A1(n10936), .A2(n7362), .ZN(n7359) );
  NAND2_X1 U8200 ( .A1(n7363), .A2(n7361), .ZN(n7360) );
  NOR2_X1 U8201 ( .A1(n10936), .A2(n7362), .ZN(n7361) );
  NAND2_X1 U8202 ( .A1(n7159), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n8267) );
  INV_X1 U8203 ( .A(n8242), .ZN(n7159) );
  NAND2_X1 U8204 ( .A1(n7158), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8283) );
  INV_X1 U8205 ( .A(n8267), .ZN(n7158) );
  NAND2_X1 U8206 ( .A1(n7348), .A2(n6456), .ZN(n7349) );
  NAND2_X1 U8207 ( .A1(n13155), .A2(n6450), .ZN(n7352) );
  AND2_X1 U8208 ( .A1(n13579), .A2(n13580), .ZN(n10563) );
  INV_X1 U8209 ( .A(n8595), .ZN(n8519) );
  AND3_X1 U8210 ( .A1(n8287), .A2(n8286), .A3(n8285), .ZN(n13386) );
  AND4_X1 U8211 ( .A1(n8161), .A2(n8160), .A3(n8159), .A4(n8158), .ZN(n13345)
         );
  NAND2_X1 U8212 ( .A1(n6665), .A2(n6664), .ZN(n15372) );
  OR2_X1 U8213 ( .A1(n15379), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U8214 ( .A1(n15379), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6664) );
  NAND2_X1 U8215 ( .A1(n6668), .A2(n15409), .ZN(n7448) );
  INV_X1 U8216 ( .A(n13629), .ZN(n6668) );
  OR2_X1 U8217 ( .A1(n10359), .A2(n10360), .ZN(n10946) );
  AND2_X1 U8218 ( .A1(n15428), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7445) );
  AND2_X1 U8219 ( .A1(n15456), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7443) );
  AOI21_X1 U8220 ( .B1(P2_REG1_REG_16__SCAN_IN), .B2(n15482), .A(n15477), .ZN(
        n15494) );
  NAND2_X1 U8221 ( .A1(n7432), .A2(n7431), .ZN(n13654) );
  INV_X1 U8222 ( .A(n7434), .ZN(n7433) );
  NAND2_X1 U8223 ( .A1(n7434), .A2(n13663), .ZN(n7431) );
  NOR2_X1 U8224 ( .A1(n13654), .A2(n13987), .ZN(n13659) );
  NOR2_X1 U8225 ( .A1(n13693), .A2(n7773), .ZN(n13683) );
  AND2_X1 U8226 ( .A1(n8683), .A2(n8577), .ZN(n13561) );
  NAND2_X1 U8227 ( .A1(n13725), .A2(n6881), .ZN(n13693) );
  INV_X1 U8228 ( .A(n7692), .ZN(n7688) );
  NAND2_X1 U8229 ( .A1(n12048), .A2(n7692), .ZN(n7691) );
  NAND2_X1 U8230 ( .A1(n12049), .A2(n13558), .ZN(n12048) );
  AND2_X1 U8231 ( .A1(n8462), .A2(n8439), .ZN(n7929) );
  NOR3_X1 U8232 ( .A1(n13820), .A2(n13432), .A3(n7769), .ZN(n13770) );
  NAND2_X1 U8233 ( .A1(n13800), .A2(n8404), .ZN(n7030) );
  NAND2_X1 U8234 ( .A1(n7032), .A2(n8403), .ZN(n13803) );
  INV_X1 U8235 ( .A(n13800), .ZN(n7032) );
  AND2_X1 U8236 ( .A1(n7695), .A2(n8676), .ZN(n7694) );
  NAND2_X1 U8237 ( .A1(n8675), .A2(n7696), .ZN(n7695) );
  INV_X1 U8238 ( .A(n8674), .ZN(n7696) );
  NAND2_X1 U8239 ( .A1(n7122), .A2(n6479), .ZN(n7389) );
  INV_X1 U8240 ( .A(n13829), .ZN(n7122) );
  INV_X1 U8241 ( .A(n8675), .ZN(n7697) );
  NAND2_X1 U8242 ( .A1(n7389), .A2(n8673), .ZN(n13816) );
  NAND2_X1 U8243 ( .A1(n8274), .A2(n8273), .ZN(n13877) );
  NAND2_X1 U8244 ( .A1(n8664), .A2(n7682), .ZN(n7681) );
  NAND2_X1 U8245 ( .A1(n11730), .A2(n11729), .ZN(n6769) );
  NAND2_X1 U8246 ( .A1(n7026), .A2(n6518), .ZN(n7025) );
  NAND2_X1 U8247 ( .A1(n13549), .A2(n7027), .ZN(n7026) );
  NAND2_X1 U8248 ( .A1(n8163), .A2(n8162), .ZN(n7027) );
  NAND2_X1 U8249 ( .A1(n11359), .A2(n7024), .ZN(n7023) );
  NOR2_X1 U8250 ( .A1(n6501), .A2(n11171), .ZN(n7401) );
  NOR2_X1 U8251 ( .A1(n6501), .A2(n7403), .ZN(n7402) );
  INV_X1 U8252 ( .A(n8656), .ZN(n7403) );
  NAND2_X1 U8253 ( .A1(n6942), .A2(n7399), .ZN(n11358) );
  INV_X1 U8254 ( .A(n7400), .ZN(n7399) );
  NAND2_X1 U8255 ( .A1(n6937), .A2(n6533), .ZN(n6942) );
  OAI21_X1 U8256 ( .B1(n7401), .B2(n7402), .A(n8657), .ZN(n7400) );
  NOR2_X1 U8257 ( .A1(n11319), .A2(n15525), .ZN(n11364) );
  NAND2_X1 U8258 ( .A1(n6937), .A2(n6939), .ZN(n7671) );
  NOR2_X1 U8259 ( .A1(n13543), .A2(n7384), .ZN(n7380) );
  INV_X1 U8260 ( .A(n8655), .ZN(n7384) );
  NOR2_X1 U8261 ( .A1(n7382), .A2(n6544), .ZN(n7381) );
  AND2_X1 U8262 ( .A1(n8655), .A2(n7383), .ZN(n7382) );
  INV_X1 U8263 ( .A(n8654), .ZN(n7383) );
  NAND2_X1 U8264 ( .A1(n7678), .A2(n10113), .ZN(n7677) );
  NAND2_X1 U8265 ( .A1(n8652), .A2(n10113), .ZN(n7676) );
  AND2_X1 U8266 ( .A1(n7943), .A2(n13545), .ZN(n7942) );
  INV_X1 U8267 ( .A(n10113), .ZN(n13542) );
  NAND2_X1 U8268 ( .A1(n8651), .A2(n7216), .ZN(n7962) );
  AND2_X1 U8269 ( .A1(n8050), .A2(n8051), .ZN(n13540) );
  OR2_X1 U8270 ( .A1(n13304), .A2(n6751), .ZN(n8050) );
  XNOR2_X1 U8271 ( .A(n13571), .B(n13579), .ZN(n8686) );
  OR2_X1 U8272 ( .A1(n14095), .A2(n13495), .ZN(n13498) );
  NOR2_X1 U8273 ( .A1(n6752), .A2(n6542), .ZN(n15512) );
  NAND2_X1 U8274 ( .A1(n8049), .A2(n6753), .ZN(n6752) );
  AND2_X1 U8275 ( .A1(n8638), .A2(n8637), .ZN(n10559) );
  AND3_X1 U8276 ( .A1(n7987), .A2(n6539), .A3(n7986), .ZN(n7988) );
  AND2_X1 U8277 ( .A1(n7985), .A2(n7984), .ZN(n7986) );
  XNOR2_X1 U8278 ( .A(n8012), .B(n8011), .ZN(n10307) );
  NAND2_X1 U8279 ( .A1(n8010), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8012) );
  INV_X1 U8280 ( .A(n8010), .ZN(n7674) );
  OR2_X1 U8281 ( .A1(n8623), .A2(n8622), .ZN(n8625) );
  OR2_X1 U8282 ( .A1(n8633), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n8616) );
  INV_X1 U8283 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7999) );
  AND2_X1 U8284 ( .A1(n8150), .A2(n8170), .ZN(n10369) );
  AND2_X1 U8285 ( .A1(n8057), .A2(n8071), .ZN(n10317) );
  NAND2_X1 U8286 ( .A1(n14252), .A2(n14251), .ZN(n6999) );
  OR2_X1 U8287 ( .A1(n9187), .A2(n14207), .ZN(n9232) );
  NAND2_X1 U8288 ( .A1(n9292), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n9312) );
  INV_X1 U8289 ( .A(n9293), .ZN(n9292) );
  INV_X1 U8290 ( .A(n7572), .ZN(n7571) );
  INV_X1 U8291 ( .A(n9288), .ZN(n7573) );
  AOI21_X1 U8292 ( .B1(n7579), .B2(n9222), .A(n7577), .ZN(n7576) );
  INV_X1 U8293 ( .A(n14201), .ZN(n7577) );
  INV_X1 U8294 ( .A(n6438), .ZN(n9388) );
  OR2_X1 U8295 ( .A1(n10260), .A2(n10261), .ZN(n10466) );
  XNOR2_X1 U8296 ( .A(n14727), .B(n14726), .ZN(n14734) );
  NAND2_X1 U8297 ( .A1(n7795), .A2(n14750), .ZN(n7550) );
  AND2_X1 U8298 ( .A1(n9404), .A2(n9371), .ZN(n14263) );
  NAND2_X1 U8299 ( .A1(n14836), .A2(n6464), .ZN(n14819) );
  AND2_X1 U8300 ( .A1(n9352), .A2(n9334), .ZN(n14841) );
  INV_X1 U8301 ( .A(n7974), .ZN(n6658) );
  NAND2_X1 U8302 ( .A1(n7551), .A2(n6474), .ZN(n14868) );
  OR2_X1 U8303 ( .A1(n9274), .A2(n9273), .ZN(n9293) );
  AOI21_X1 U8304 ( .B1(n7801), .B2(n7802), .A(n7800), .ZN(n7799) );
  INV_X1 U8305 ( .A(n14907), .ZN(n7800) );
  INV_X1 U8306 ( .A(n12129), .ZN(n7259) );
  NAND2_X1 U8307 ( .A1(n14974), .A2(n15124), .ZN(n14975) );
  OR2_X1 U8308 ( .A1(n11928), .A2(n14516), .ZN(n11926) );
  OR2_X1 U8309 ( .A1(n6724), .A2(n7963), .ZN(n6721) );
  NAND2_X1 U8310 ( .A1(n11485), .A2(n11799), .ZN(n11794) );
  NAND2_X1 U8311 ( .A1(n7240), .A2(n11471), .ZN(n11551) );
  NAND2_X1 U8312 ( .A1(n7239), .A2(n6681), .ZN(n6680) );
  NAND3_X1 U8313 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n9001) );
  OAI21_X1 U8314 ( .B1(n15279), .B2(n8892), .A(n11021), .ZN(n15255) );
  NAND2_X1 U8315 ( .A1(n8866), .A2(n8824), .ZN(n8826) );
  OR2_X1 U8316 ( .A1(n10257), .A2(P1_IR_REG_27__SCAN_IN), .ZN(n7265) );
  NAND2_X1 U8317 ( .A1(n14286), .A2(n11494), .ZN(n10824) );
  INV_X1 U8318 ( .A(n15041), .ZN(n7475) );
  INV_X1 U8319 ( .A(n15040), .ZN(n7474) );
  INV_X1 U8320 ( .A(n15336), .ZN(n15344) );
  NAND2_X1 U8321 ( .A1(n15294), .A2(n15320), .ZN(n15327) );
  NAND2_X1 U8322 ( .A1(n15264), .A2(n14738), .ZN(n15030) );
  INV_X1 U8323 ( .A(n15327), .ZN(n15340) );
  AND3_X1 U8324 ( .A1(n10244), .A2(P1_STATE_REG_SCAN_IN), .A3(n10106), .ZN(
        n10813) );
  INV_X1 U8325 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n8820) );
  NOR2_X1 U8326 ( .A1(n12033), .A2(n7898), .ZN(n7897) );
  INV_X1 U8327 ( .A(n12031), .ZN(n7898) );
  XNOR2_X1 U8328 ( .A(n8847), .B(P1_IR_REG_26__SCAN_IN), .ZN(n10182) );
  XNOR2_X1 U8329 ( .A(n8845), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9430) );
  NAND2_X1 U8330 ( .A1(n7510), .A2(n8859), .ZN(n7509) );
  INV_X1 U8331 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n8850) );
  NAND2_X1 U8332 ( .A1(n8886), .A2(n8817), .ZN(n8944) );
  INV_X1 U8333 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8817) );
  NAND2_X1 U8334 ( .A1(n8743), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n8742) );
  XNOR2_X1 U8335 ( .A(n8705), .B(n15781), .ZN(n8738) );
  NAND2_X1 U8336 ( .A1(n6682), .A2(n8712), .ZN(n8757) );
  NAND2_X1 U8337 ( .A1(n8752), .A2(n14620), .ZN(n6682) );
  OAI21_X1 U8338 ( .B1(P3_ADDR_REG_8__SCAN_IN), .B2(n8719), .A(n8718), .ZN(
        n8735) );
  NAND2_X1 U8339 ( .A1(n8721), .A2(n6683), .ZN(n8770) );
  NAND2_X1 U8340 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(n6684), .ZN(n6683) );
  OAI22_X1 U8341 ( .A1(n8776), .A2(n8725), .B1(P1_ADDR_REG_13__SCAN_IN), .B2(
        n8726), .ZN(n8779) );
  AOI21_X2 U8342 ( .B1(n15231), .B2(n6504), .A(n7303), .ZN(n8784) );
  NAND2_X1 U8343 ( .A1(n7305), .A2(n7304), .ZN(n7303) );
  NAND2_X1 U8344 ( .A1(n6454), .A2(n7312), .ZN(n7304) );
  NAND2_X1 U8345 ( .A1(n15221), .A2(n8790), .ZN(n15201) );
  NAND2_X1 U8346 ( .A1(n7859), .A2(n7857), .ZN(n12228) );
  AOI21_X1 U8347 ( .B1(n7860), .B2(n7862), .A(n7858), .ZN(n7857) );
  NAND2_X1 U8348 ( .A1(n10642), .A2(n10641), .ZN(n10652) );
  INV_X1 U8349 ( .A(n13044), .ZN(n12249) );
  NAND2_X1 U8350 ( .A1(n7864), .A2(n7865), .ZN(n12267) );
  NAND2_X1 U8351 ( .A1(n12219), .A2(n7866), .ZN(n7864) );
  AND2_X1 U8352 ( .A1(n9814), .A2(n9813), .ZN(n12281) );
  INV_X1 U8353 ( .A(n12320), .ZN(n12570) );
  INV_X1 U8354 ( .A(n12281), .ZN(n12916) );
  OAI211_X1 U8355 ( .C1(n12363), .C2(n15696), .A(n9796), .B(n9795), .ZN(n12905) );
  NOR2_X1 U8356 ( .A1(n6889), .A2(n10398), .ZN(n10515) );
  NOR2_X1 U8357 ( .A1(n10528), .A2(n6566), .ZN(n6889) );
  AND2_X1 U8358 ( .A1(n10406), .A2(n10403), .ZN(n10664) );
  NAND2_X1 U8359 ( .A1(n10664), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10663) );
  NAND2_X1 U8360 ( .A1(n10439), .A2(n10440), .ZN(n10689) );
  NAND2_X1 U8361 ( .A1(n12604), .A2(n12603), .ZN(n12615) );
  AND2_X1 U8362 ( .A1(n7048), .A2(n7045), .ZN(n12748) );
  INV_X1 U8363 ( .A(n7049), .ZN(n7045) );
  NAND2_X1 U8364 ( .A1(n12712), .A2(n7050), .ZN(n7048) );
  NAND2_X1 U8365 ( .A1(n15598), .A2(n6986), .ZN(n7378) );
  INV_X1 U8366 ( .A(n12728), .ZN(n7379) );
  AND2_X1 U8367 ( .A1(n12726), .A2(n12727), .ZN(n7377) );
  AND2_X1 U8368 ( .A1(n10126), .A2(n7168), .ZN(n15591) );
  NAND2_X1 U8369 ( .A1(n12934), .A2(n12978), .ZN(n6667) );
  OR2_X1 U8370 ( .A1(n12783), .A2(n12834), .ZN(n6711) );
  NAND2_X1 U8371 ( .A1(n9902), .A2(n9901), .ZN(n12944) );
  NAND2_X1 U8372 ( .A1(n7663), .A2(n9892), .ZN(n12833) );
  NOR2_X1 U8373 ( .A1(n9989), .A2(SI_4_), .ZN(n7132) );
  NOR2_X1 U8374 ( .A1(n10509), .A2(n15608), .ZN(n12762) );
  NAND2_X1 U8375 ( .A1(n10543), .A2(n10508), .ZN(n15610) );
  NAND2_X1 U8376 ( .A1(n12762), .A2(n12933), .ZN(n12828) );
  NAND2_X2 U8377 ( .A1(n10509), .A2(n15610), .ZN(n15616) );
  INV_X1 U8378 ( .A(n12375), .ZN(n12924) );
  NAND2_X1 U8379 ( .A1(n12370), .A2(n12369), .ZN(n12925) );
  NAND2_X1 U8380 ( .A1(n13098), .A2(n6448), .ZN(n12941) );
  NAND2_X1 U8381 ( .A1(n7070), .A2(n10021), .ZN(n12764) );
  NOR2_X1 U8382 ( .A1(n10020), .A2(n10019), .ZN(n10021) );
  NAND2_X1 U8383 ( .A1(n9975), .A2(n9974), .ZN(n13001) );
  XNOR2_X1 U8384 ( .A(n12770), .B(n12769), .ZN(n13004) );
  NAND2_X1 U8385 ( .A1(n9869), .A2(n9868), .ZN(n13032) );
  NAND2_X1 U8386 ( .A1(n7952), .A2(n9831), .ZN(n12886) );
  NAND2_X1 U8387 ( .A1(n9806), .A2(n9805), .ZN(n13056) );
  NAND2_X1 U8388 ( .A1(n7137), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7136) );
  NAND2_X1 U8389 ( .A1(n7006), .A2(n7007), .ZN(n12017) );
  NAND2_X1 U8390 ( .A1(n13933), .A2(n13280), .ZN(n12022) );
  INV_X1 U8391 ( .A(n12016), .ZN(n7005) );
  NAND2_X1 U8392 ( .A1(n12187), .A2(n7003), .ZN(n12197) );
  AND2_X1 U8393 ( .A1(n12188), .A2(n11657), .ZN(n7003) );
  NAND2_X1 U8394 ( .A1(n11953), .A2(n11667), .ZN(n7502) );
  INV_X1 U8395 ( .A(n13251), .ZN(n7015) );
  NAND2_X1 U8396 ( .A1(n13229), .A2(n13609), .ZN(n6935) );
  NAND2_X1 U8397 ( .A1(n10727), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13277) );
  INV_X1 U8398 ( .A(n13227), .ZN(n13280) );
  INV_X1 U8399 ( .A(n13437), .ZN(n13593) );
  INV_X1 U8400 ( .A(n13203), .ZN(n13782) );
  INV_X1 U8401 ( .A(n13126), .ZN(n13596) );
  INV_X1 U8402 ( .A(n13392), .ZN(n13881) );
  INV_X1 U8403 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n7292) );
  OR2_X1 U8404 ( .A1(n8077), .A2(n7991), .ZN(n7996) );
  AND3_X1 U8405 ( .A1(n6947), .A2(n6949), .A3(n6950), .ZN(n6946) );
  INV_X1 U8406 ( .A(n13293), .ZN(n13612) );
  AND2_X1 U8407 ( .A1(n15419), .A2(n10948), .ZN(n10950) );
  AOI21_X1 U8408 ( .B1(n13671), .B2(n15486), .A(n7441), .ZN(n7440) );
  NAND2_X1 U8409 ( .A1(n8557), .A2(n6773), .ZN(n7034) );
  AOI21_X1 U8410 ( .B1(n7199), .B2(n13897), .A(n7196), .ZN(n13721) );
  NAND2_X1 U8411 ( .A1(n7198), .A2(n7197), .ZN(n7196) );
  NAND2_X1 U8412 ( .A1(n13716), .A2(n7200), .ZN(n7199) );
  NAND2_X1 U8413 ( .A1(n15507), .A2(n8649), .ZN(n13843) );
  AND2_X1 U8414 ( .A1(n15538), .A2(n15524), .ZN(n14023) );
  NAND2_X1 U8415 ( .A1(n7142), .A2(n15522), .ZN(n7141) );
  INV_X1 U8416 ( .A(n11948), .ZN(n7142) );
  NOR2_X1 U8417 ( .A1(n13942), .A2(n7193), .ZN(n14050) );
  NAND2_X1 U8418 ( .A1(n7195), .A2(n7194), .ZN(n7193) );
  INV_X1 U8419 ( .A(n13943), .ZN(n7194) );
  NAND2_X1 U8420 ( .A1(n13944), .A2(n15522), .ZN(n7195) );
  AND2_X1 U8421 ( .A1(n15533), .A2(n15524), .ZN(n14086) );
  NAND2_X1 U8422 ( .A1(n8630), .A2(n8629), .ZN(n15506) );
  INV_X1 U8423 ( .A(n15507), .ZN(n15509) );
  NAND2_X1 U8424 ( .A1(n14221), .A2(n7574), .ZN(n14159) );
  NAND2_X1 U8425 ( .A1(n9348), .A2(n9347), .ZN(n14178) );
  AND2_X1 U8426 ( .A1(n14840), .A2(n15336), .ZN(n15073) );
  OAI21_X1 U8427 ( .B1(n14252), .B2(n6997), .A(n6995), .ZN(n14223) );
  NAND2_X1 U8428 ( .A1(n14532), .A2(n6861), .ZN(n6860) );
  INV_X1 U8429 ( .A(n14533), .ZN(n6861) );
  INV_X1 U8430 ( .A(n14532), .ZN(n6854) );
  AOI21_X1 U8431 ( .B1(n14421), .B2(n7507), .A(n14473), .ZN(n7505) );
  NOR2_X1 U8432 ( .A1(n14423), .A2(n14422), .ZN(n14445) );
  AND2_X1 U8433 ( .A1(n14486), .A2(n11451), .ZN(n6855) );
  INV_X1 U8434 ( .A(n14538), .ZN(n6857) );
  OR2_X1 U8435 ( .A1(n9190), .A2(n9189), .ZN(n14954) );
  AND2_X1 U8436 ( .A1(n11372), .A2(n11371), .ZN(n11373) );
  XNOR2_X1 U8437 ( .A(n7544), .B(n14757), .ZN(n15042) );
  AOI21_X1 U8438 ( .B1(n7548), .B2(n7546), .A(n7972), .ZN(n7545) );
  INV_X1 U8439 ( .A(n7548), .ZN(n7547) );
  XNOR2_X1 U8440 ( .A(n14752), .B(n14757), .ZN(n15043) );
  OAI21_X1 U8441 ( .B1(n14749), .B2(n7787), .A(n7783), .ZN(n7793) );
  AOI21_X1 U8442 ( .B1(n7786), .B2(n7785), .A(n7784), .ZN(n7783) );
  NAND2_X1 U8443 ( .A1(n14833), .A2(n15008), .ZN(n12115) );
  NAND2_X1 U8444 ( .A1(n6496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U8445 ( .A1(n7630), .A2(n8759), .ZN(n7629) );
  INV_X1 U8446 ( .A(n15823), .ZN(n6828) );
  INV_X1 U8447 ( .A(n8768), .ZN(n7301) );
  NAND2_X1 U8448 ( .A1(n15220), .A2(n15431), .ZN(n15218) );
  OR2_X1 U8449 ( .A1(n15231), .A2(n7312), .ZN(n7310) );
  INV_X1 U8450 ( .A(n8787), .ZN(n7639) );
  INV_X1 U8451 ( .A(n12401), .ZN(n7332) );
  NOR2_X1 U8452 ( .A1(n12401), .A2(n12513), .ZN(n7329) );
  NAND2_X1 U8453 ( .A1(n7908), .A2(n7907), .ZN(n7905) );
  NAND2_X1 U8454 ( .A1(n6590), .A2(n13331), .ZN(n7906) );
  NAND2_X1 U8455 ( .A1(n14307), .A2(n6846), .ZN(n6845) );
  NAND2_X1 U8456 ( .A1(n6731), .A2(n6730), .ZN(n13355) );
  OAI21_X1 U8457 ( .B1(n6729), .B2(n6728), .A(n6726), .ZN(n6731) );
  AOI21_X1 U8458 ( .B1(n6727), .B2(n13349), .A(n13348), .ZN(n6726) );
  NAND2_X1 U8459 ( .A1(n12438), .A2(n12532), .ZN(n7333) );
  AOI21_X1 U8460 ( .B1(n7337), .B2(n7336), .A(n7335), .ZN(n7334) );
  NOR2_X1 U8461 ( .A1(n7287), .A2(n6546), .ZN(n7286) );
  INV_X1 U8462 ( .A(n7289), .ZN(n7287) );
  AND2_X1 U8463 ( .A1(n6873), .A2(n6871), .ZN(n6870) );
  INV_X1 U8464 ( .A(n7532), .ZN(n6873) );
  NAND2_X1 U8465 ( .A1(n7529), .A2(n7527), .ZN(n14357) );
  AOI21_X1 U8466 ( .B1(n7532), .B2(n7530), .A(n7528), .ZN(n7527) );
  INV_X1 U8467 ( .A(n14358), .ZN(n7528) );
  NAND2_X1 U8468 ( .A1(n7900), .A2(n6747), .ZN(n6746) );
  NOR2_X1 U8469 ( .A1(n6749), .A2(n6748), .ZN(n6747) );
  INV_X1 U8470 ( .A(n6546), .ZN(n6749) );
  OAI21_X1 U8471 ( .B1(n7318), .B2(n6481), .A(n7319), .ZN(n12475) );
  INV_X1 U8472 ( .A(n12488), .ZN(n7180) );
  NOR2_X1 U8473 ( .A1(n7285), .A2(n13388), .ZN(n7282) );
  AND2_X1 U8474 ( .A1(n7285), .A2(n13388), .ZN(n7284) );
  AND2_X1 U8475 ( .A1(n14376), .A2(n14377), .ZN(n14378) );
  NAND2_X1 U8476 ( .A1(n14365), .A2(n6517), .ZN(n14377) );
  AOI22_X1 U8477 ( .A1(n14375), .A2(n14374), .B1(n14373), .B2(n14372), .ZN(
        n14376) );
  NAND2_X1 U8478 ( .A1(n7918), .A2(n7917), .ZN(n7916) );
  INV_X1 U8479 ( .A(n13416), .ZN(n7917) );
  INV_X1 U8480 ( .A(n13417), .ZN(n7918) );
  NOR4_X1 U8481 ( .A1(n14507), .A2(n14506), .A3(n14505), .A4(n14504), .ZN(
        n14512) );
  INV_X1 U8482 ( .A(n14403), .ZN(n7537) );
  NOR2_X1 U8483 ( .A1(n12539), .A2(n6788), .ZN(n6787) );
  NAND2_X1 U8484 ( .A1(n12537), .A2(n6469), .ZN(n6788) );
  NOR2_X1 U8485 ( .A1(n12533), .A2(n12534), .ZN(n6789) );
  NAND2_X1 U8486 ( .A1(n12494), .A2(n6555), .ZN(n7327) );
  INV_X1 U8487 ( .A(n7916), .ZN(n7913) );
  AND2_X1 U8488 ( .A1(n13416), .A2(n13417), .ZN(n7919) );
  OR2_X1 U8489 ( .A1(n6868), .A2(n6865), .ZN(n6864) );
  AND2_X1 U8490 ( .A1(n7536), .A2(n14408), .ZN(n6868) );
  AND2_X1 U8491 ( .A1(n7536), .A2(n6866), .ZN(n6865) );
  AOI21_X1 U8492 ( .B1(n14407), .B2(n14406), .A(n7537), .ZN(n7536) );
  INV_X1 U8493 ( .A(n7535), .ZN(n7534) );
  NAND2_X1 U8494 ( .A1(n7344), .A2(n6537), .ZN(n7343) );
  NAND2_X1 U8495 ( .A1(n7596), .A2(n7598), .ZN(n7594) );
  OAI211_X1 U8496 ( .C1(n7602), .C2(n7590), .A(n12657), .B(n6898), .ZN(n6897)
         );
  NAND2_X1 U8497 ( .A1(n7606), .A2(n6899), .ZN(n6898) );
  NOR2_X1 U8498 ( .A1(n12646), .A2(n7590), .ZN(n6899) );
  NAND2_X1 U8499 ( .A1(n6921), .A2(n6920), .ZN(n6919) );
  INV_X1 U8500 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U8501 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_22__SCAN_IN), .ZN(
        n7140) );
  NOR2_X1 U8502 ( .A1(n13736), .A2(n7923), .ZN(n7922) );
  INV_X1 U8503 ( .A(n8489), .ZN(n7923) );
  INV_X1 U8504 ( .A(n9312), .ZN(n9310) );
  NOR2_X1 U8505 ( .A1(n9332), .A2(n9311), .ZN(n7278) );
  NAND2_X1 U8506 ( .A1(n14557), .A2(n15286), .ZN(n14287) );
  INV_X1 U8507 ( .A(n12091), .ZN(n7242) );
  INV_X1 U8508 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9896) );
  INV_X1 U8509 ( .A(n8358), .ZN(n7883) );
  OAI21_X1 U8510 ( .B1(n8336), .B2(n7883), .A(n8379), .ZN(n7882) );
  INV_X1 U8511 ( .A(n7343), .ZN(n7342) );
  NAND2_X1 U8512 ( .A1(n8260), .A2(n10283), .ZN(n8276) );
  NAND2_X1 U8513 ( .A1(n8209), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n6674) );
  AOI21_X1 U8514 ( .B1(n7312), .B2(n7311), .A(n15234), .ZN(n7309) );
  XNOR2_X1 U8515 ( .A(n6446), .B(n7130), .ZN(n10653) );
  AND2_X1 U8516 ( .A1(n11639), .A2(n12575), .ZN(n7872) );
  NAND2_X1 U8517 ( .A1(n11640), .A2(n11641), .ZN(n7870) );
  INV_X1 U8518 ( .A(n7868), .ZN(n7118) );
  NOR2_X1 U8519 ( .A1(n12781), .A2(n12523), .ZN(n6815) );
  NOR2_X1 U8520 ( .A1(n12545), .A2(n6817), .ZN(n6816) );
  INV_X1 U8521 ( .A(n6571), .ZN(n6813) );
  NAND2_X1 U8522 ( .A1(n7183), .A2(n7182), .ZN(n7708) );
  AOI21_X1 U8523 ( .B1(n12511), .B2(n12507), .A(n7315), .ZN(n7314) );
  OAI21_X1 U8524 ( .B1(n13085), .B2(P3_REG2_REG_1__SCAN_IN), .A(n7375), .ZN(
        n10383) );
  NAND2_X1 U8525 ( .A1(n13085), .A2(n10382), .ZN(n7375) );
  OR2_X1 U8526 ( .A1(n10446), .A2(n10682), .ZN(n10447) );
  OAI21_X1 U8527 ( .B1(n6911), .B2(n6909), .A(n6908), .ZN(n6907) );
  NAND2_X1 U8528 ( .A1(n11219), .A2(n6912), .ZN(n6908) );
  AND2_X1 U8529 ( .A1(n6971), .A2(n6970), .ZN(n6969) );
  INV_X1 U8530 ( .A(n15593), .ZN(n6970) );
  NAND2_X1 U8531 ( .A1(n12694), .A2(n6895), .ZN(n12696) );
  NAND2_X1 U8532 ( .A1(n12701), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n6895) );
  AOI21_X1 U8533 ( .B1(n7832), .B2(n7835), .A(n6502), .ZN(n7831) );
  NAND2_X1 U8534 ( .A1(n12506), .A2(n12509), .ZN(n7834) );
  AND2_X1 U8535 ( .A1(n9997), .A2(n12385), .ZN(n12377) );
  INV_X1 U8536 ( .A(n9950), .ZN(n7661) );
  INV_X1 U8537 ( .A(n12779), .ZN(n12781) );
  INV_X1 U8538 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n6924) );
  INV_X1 U8539 ( .A(n7824), .ZN(n7820) );
  NOR2_X1 U8540 ( .A1(n7822), .A2(n7427), .ZN(n7426) );
  INV_X1 U8541 ( .A(n12454), .ZN(n7427) );
  NOR2_X1 U8542 ( .A1(n9705), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U8543 ( .A1(n9633), .A2(n7647), .ZN(n7646) );
  INV_X1 U8544 ( .A(n9633), .ZN(n7648) );
  NAND2_X1 U8545 ( .A1(n9625), .A2(n6519), .ZN(n9669) );
  NAND2_X1 U8546 ( .A1(n12580), .A2(n10971), .ZN(n12427) );
  INV_X1 U8547 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n9536) );
  NAND2_X1 U8548 ( .A1(n6447), .A2(n8017), .ZN(n9522) );
  NAND2_X1 U8549 ( .A1(n7659), .A2(n7661), .ZN(n7656) );
  NOR2_X1 U8550 ( .A1(n12779), .A2(n7658), .ZN(n7657) );
  INV_X1 U8551 ( .A(n7659), .ZN(n7658) );
  AND2_X1 U8552 ( .A1(n13001), .A2(n12230), .ZN(n10081) );
  OR2_X1 U8553 ( .A1(n13001), .A2(n12230), .ZN(n12515) );
  INV_X1 U8554 ( .A(n6708), .ZN(n6707) );
  INV_X1 U8555 ( .A(n7424), .ZN(n6706) );
  NOR2_X1 U8556 ( .A1(n12505), .A2(n7425), .ZN(n7424) );
  INV_X1 U8557 ( .A(n12501), .ZN(n7425) );
  AOI21_X1 U8558 ( .B1(n7424), .B2(n12820), .A(n6709), .ZN(n6708) );
  AOI21_X1 U8559 ( .B1(n7814), .B2(n7812), .A(n7811), .ZN(n7810) );
  INV_X1 U8560 ( .A(n12487), .ZN(n7811) );
  INV_X1 U8561 ( .A(n7816), .ZN(n7812) );
  NOR2_X1 U8562 ( .A1(n7813), .A2(n6699), .ZN(n6697) );
  INV_X1 U8563 ( .A(n7814), .ZN(n7813) );
  NOR2_X1 U8564 ( .A1(n7840), .A2(n7839), .ZN(n7838) );
  INV_X1 U8565 ( .A(n12580), .ZN(n7154) );
  NAND2_X1 U8566 ( .A1(n7156), .A2(n9479), .ZN(n10052) );
  AND2_X1 U8567 ( .A1(n7750), .A2(n7754), .ZN(n7749) );
  NOR2_X1 U8568 ( .A1(n9924), .A2(n7755), .ZN(n7754) );
  NAND2_X1 U8569 ( .A1(n9899), .A2(n7751), .ZN(n7750) );
  INV_X1 U8570 ( .A(n9923), .ZN(n7746) );
  NAND2_X1 U8571 ( .A1(n7757), .A2(n9923), .ZN(n7748) );
  INV_X1 U8572 ( .A(n9894), .ZN(n7757) );
  INV_X1 U8573 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n10003) );
  NAND2_X1 U8574 ( .A1(n10004), .A2(n10003), .ZN(n10009) );
  NOR2_X1 U8575 ( .A1(n9817), .A2(n9816), .ZN(n10002) );
  INV_X1 U8576 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9835) );
  AOI21_X1 U8577 ( .B1(n6796), .B2(n6794), .A(n6633), .ZN(n6793) );
  INV_X1 U8578 ( .A(n7729), .ZN(n6794) );
  INV_X1 U8579 ( .A(n6796), .ZN(n6795) );
  INV_X1 U8580 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9751) );
  AOI21_X1 U8581 ( .B1(n6803), .B2(n6805), .A(n6587), .ZN(n6801) );
  INV_X1 U8582 ( .A(n6803), .ZN(n6802) );
  INV_X1 U8583 ( .A(n7744), .ZN(n7740) );
  NOR2_X1 U8584 ( .A1(n8302), .A2(n8301), .ZN(n8325) );
  NOR2_X1 U8585 ( .A1(n7481), .A2(n7351), .ZN(n7350) );
  INV_X1 U8586 ( .A(n7353), .ZN(n7351) );
  OR2_X1 U8587 ( .A1(n13180), .A2(n12002), .ZN(n7481) );
  INV_X1 U8588 ( .A(n8393), .ZN(n7362) );
  OR3_X1 U8589 ( .A1(n13488), .A2(n13487), .A3(n13486), .ZN(n13516) );
  NAND2_X1 U8590 ( .A1(n6757), .A2(n7294), .ZN(n13435) );
  AOI21_X1 U8591 ( .B1(n7911), .B2(n6557), .A(n7295), .ZN(n7294) );
  NAND2_X1 U8592 ( .A1(n6759), .A2(n6758), .ZN(n6757) );
  NOR2_X1 U8593 ( .A1(n13524), .A2(n13473), .ZN(n13521) );
  AND2_X1 U8594 ( .A1(n7149), .A2(n13556), .ZN(n13557) );
  NOR2_X1 U8595 ( .A1(n8677), .A2(n6678), .ZN(n6677) );
  NOR2_X1 U8596 ( .A1(n13801), .A2(n7150), .ZN(n7149) );
  INV_X1 U8597 ( .A(n13704), .ZN(n6675) );
  INV_X1 U8598 ( .A(n13760), .ZN(n6676) );
  NOR2_X1 U8599 ( .A1(n13940), .A2(n13933), .ZN(n6881) );
  NOR2_X1 U8600 ( .A1(n8535), .A2(n8534), .ZN(n7160) );
  NOR2_X1 U8601 ( .A1(n8480), .A2(n13117), .ZN(n6687) );
  INV_X1 U8602 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8282) );
  NAND2_X1 U8603 ( .A1(n6770), .A2(n6772), .ZN(n6768) );
  INV_X1 U8604 ( .A(n7926), .ZN(n7925) );
  INV_X1 U8605 ( .A(n8225), .ZN(n6772) );
  INV_X1 U8606 ( .A(n8663), .ZN(n7684) );
  AND2_X1 U8607 ( .A1(n11710), .A2(n7024), .ZN(n7020) );
  INV_X1 U8608 ( .A(n11709), .ZN(n7019) );
  NOR2_X1 U8609 ( .A1(n13365), .A2(n7766), .ZN(n7765) );
  INV_X1 U8610 ( .A(n7401), .ZN(n6936) );
  INV_X1 U8611 ( .A(n8102), .ZN(n6765) );
  INV_X1 U8612 ( .A(n11185), .ZN(n7946) );
  NOR2_X1 U8613 ( .A1(n7946), .A2(n7947), .ZN(n7945) );
  INV_X1 U8614 ( .A(n8065), .ZN(n7947) );
  AND2_X1 U8615 ( .A1(n8102), .A2(n8101), .ZN(n13545) );
  AND2_X1 U8616 ( .A1(n7215), .A2(n8032), .ZN(n13541) );
  INV_X1 U8617 ( .A(n13916), .ZN(n7216) );
  INV_X1 U8618 ( .A(n7220), .ZN(n7219) );
  OAI21_X1 U8619 ( .B1(n7938), .B2(n7937), .A(n8378), .ZN(n7220) );
  OAI21_X1 U8620 ( .B1(n13877), .B2(n13889), .A(n8288), .ZN(n13870) );
  OR2_X1 U8621 ( .A1(n13495), .A2(n10165), .ZN(n6753) );
  OR2_X1 U8622 ( .A1(n8147), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8149) );
  OR2_X1 U8623 ( .A1(n14105), .A2(n9055), .ZN(n7558) );
  OR2_X1 U8624 ( .A1(n9222), .A2(n9178), .ZN(n7580) );
  NOR2_X1 U8625 ( .A1(n11311), .A2(n9124), .ZN(n7273) );
  AND2_X1 U8626 ( .A1(n8864), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9184) );
  XNOR2_X1 U8627 ( .A(n14527), .B(n14738), .ZN(n14529) );
  NAND2_X1 U8628 ( .A1(n6869), .A2(n7512), .ZN(n7511) );
  NAND2_X1 U8629 ( .A1(n7518), .A2(n7523), .ZN(n7515) );
  NAND2_X1 U8630 ( .A1(n7971), .A2(n7247), .ZN(n7246) );
  INV_X1 U8631 ( .A(n7248), .ZN(n7247) );
  AND2_X1 U8632 ( .A1(n6464), .A2(n7470), .ZN(n7469) );
  NAND2_X1 U8633 ( .A1(n14860), .A2(n7779), .ZN(n7778) );
  NOR2_X1 U8634 ( .A1(n14830), .A2(n7251), .ZN(n7250) );
  INV_X1 U8635 ( .A(n12136), .ZN(n7251) );
  INV_X1 U8636 ( .A(n7258), .ZN(n7257) );
  NAND2_X1 U8637 ( .A1(n7543), .A2(n7254), .ZN(n7253) );
  OAI21_X1 U8638 ( .B1(n6459), .B2(n7259), .A(n14912), .ZN(n7258) );
  NOR2_X1 U8639 ( .A1(n15096), .A2(n15104), .ZN(n7467) );
  NOR2_X1 U8640 ( .A1(n14975), .A2(n14960), .ZN(n14933) );
  NAND2_X1 U8641 ( .A1(n14344), .A2(n14343), .ZN(n6725) );
  INV_X1 U8642 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n9060) );
  NOR2_X1 U8643 ( .A1(n11470), .A2(n14501), .ZN(n6681) );
  AND4_X1 U8644 ( .A1(n7456), .A2(n11406), .A3(n11051), .A4(n6410), .ZN(n11476) );
  INV_X1 U8645 ( .A(n14553), .ZN(n11405) );
  NAND2_X1 U8646 ( .A1(n11405), .A2(n14319), .ZN(n11409) );
  NAND2_X1 U8647 ( .A1(n11479), .A2(n11409), .ZN(n14504) );
  NOR2_X1 U8648 ( .A1(n14309), .A2(n14313), .ZN(n7456) );
  NAND2_X1 U8649 ( .A1(n14287), .A2(n14289), .ZN(n14502) );
  NAND2_X1 U8650 ( .A1(n7464), .A2(n8823), .ZN(n7264) );
  AOI21_X1 U8651 ( .B1(n7887), .B2(n7885), .A(n6634), .ZN(n7884) );
  INV_X1 U8652 ( .A(n7887), .ZN(n7886) );
  XNOR2_X1 U8653 ( .A(n8506), .B(n8508), .ZN(n8490) );
  AND2_X1 U8654 ( .A1(n6466), .A2(n8853), .ZN(n6862) );
  OAI211_X1 U8655 ( .C1(n8104), .C2(n6990), .A(n6988), .B(n8121), .ZN(n8125)
         );
  NAND2_X1 U8656 ( .A1(n7642), .A2(n8710), .ZN(n8711) );
  XNOR2_X1 U8657 ( .A(n8711), .B(n7641), .ZN(n8752) );
  INV_X1 U8658 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7641) );
  NAND2_X1 U8659 ( .A1(n8716), .A2(n8717), .ZN(n8761) );
  NOR2_X1 U8660 ( .A1(n8720), .A2(n7166), .ZN(n8766) );
  AND2_X1 U8661 ( .A1(n14664), .A2(P3_ADDR_REG_9__SCAN_IN), .ZN(n7166) );
  INV_X1 U8662 ( .A(n7622), .ZN(n7620) );
  NOR2_X1 U8663 ( .A1(n7622), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7621) );
  NOR2_X1 U8664 ( .A1(n15224), .A2(n7625), .ZN(n7622) );
  NAND2_X1 U8665 ( .A1(n15224), .A2(n7625), .ZN(n7623) );
  AOI21_X1 U8666 ( .B1(n7309), .B2(n7307), .A(P2_ADDR_REG_14__SCAN_IN), .ZN(
        n7306) );
  INV_X1 U8667 ( .A(n7311), .ZN(n7307) );
  NAND2_X1 U8668 ( .A1(n7306), .A2(n7308), .ZN(n7305) );
  INV_X1 U8669 ( .A(n7309), .ZN(n7308) );
  AOI22_X1 U8670 ( .A1(n8782), .A2(n8729), .B1(P3_ADDR_REG_15__SCAN_IN), .B2(
        n11631), .ZN(n8785) );
  INV_X1 U8671 ( .A(n12339), .ZN(n7858) );
  OR2_X1 U8672 ( .A1(n11672), .A2(n12573), .ZN(n7868) );
  AND2_X1 U8673 ( .A1(n6519), .A2(n9668), .ZN(n6928) );
  INV_X1 U8674 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n9668) );
  INV_X1 U8675 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10657) );
  NAND2_X1 U8676 ( .A1(n7094), .A2(n7208), .ZN(n10916) );
  INV_X1 U8677 ( .A(n10873), .ZN(n7094) );
  INV_X1 U8678 ( .A(n12214), .ZN(n7207) );
  INV_X1 U8679 ( .A(n7099), .ZN(n7098) );
  INV_X1 U8680 ( .A(n7102), .ZN(n7097) );
  AND2_X1 U8681 ( .A1(n7105), .A2(n7100), .ZN(n7099) );
  INV_X1 U8682 ( .A(n12241), .ZN(n7100) );
  NAND2_X1 U8683 ( .A1(n7093), .A2(n7092), .ZN(n11637) );
  AOI21_X1 U8684 ( .B1(n10915), .B2(n10874), .A(n6540), .ZN(n7092) );
  OR2_X1 U8685 ( .A1(n12211), .A2(n12281), .ZN(n7109) );
  NAND4_X1 U8686 ( .A1(n9535), .A2(n9536), .A3(n10657), .A4(n6930), .ZN(n9626)
         );
  INV_X1 U8687 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n6930) );
  AOI21_X1 U8688 ( .B1(n6506), .B2(n7861), .A(n6451), .ZN(n7860) );
  INV_X1 U8689 ( .A(n7866), .ZN(n7861) );
  INV_X1 U8690 ( .A(n6506), .ZN(n7862) );
  NAND2_X1 U8691 ( .A1(n9992), .A2(n9991), .ZN(n12366) );
  AOI21_X1 U8692 ( .B1(n12792), .B2(n9991), .A(n9949), .ZN(n12269) );
  NOR2_X1 U8693 ( .A1(n9530), .A2(n7410), .ZN(n10398) );
  NAND2_X1 U8694 ( .A1(n6644), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n15547) );
  AND2_X1 U8695 ( .A1(n15553), .A2(n7370), .ZN(n6963) );
  NAND2_X1 U8696 ( .A1(n7371), .A2(n10688), .ZN(n7370) );
  INV_X1 U8697 ( .A(n10440), .ZN(n7371) );
  AND2_X1 U8698 ( .A1(n15567), .A2(n10694), .ZN(n10695) );
  NAND2_X1 U8699 ( .A1(n15561), .A2(n11224), .ZN(n11686) );
  NAND2_X1 U8700 ( .A1(n7613), .A2(n6489), .ZN(n15585) );
  NAND2_X1 U8701 ( .A1(n7038), .A2(n6516), .ZN(n12610) );
  XNOR2_X1 U8702 ( .A(n12684), .B(n12661), .ZN(n12664) );
  AND2_X1 U8703 ( .A1(n7367), .A2(n7366), .ZN(n12704) );
  NAND2_X1 U8704 ( .A1(n12701), .A2(n12702), .ZN(n7366) );
  NOR2_X1 U8705 ( .A1(n12704), .A2(n12703), .ZN(n12723) );
  AND2_X1 U8706 ( .A1(n12713), .A2(n15723), .ZN(n7049) );
  AOI21_X1 U8707 ( .B1(n7043), .B2(n7046), .A(n6652), .ZN(n7042) );
  INV_X1 U8708 ( .A(n7050), .ZN(n7043) );
  NOR2_X1 U8709 ( .A1(n12723), .A2(n7364), .ZN(n12736) );
  NOR2_X1 U8710 ( .A1(n12713), .A2(n7365), .ZN(n7364) );
  INV_X1 U8711 ( .A(n12725), .ZN(n7365) );
  AND2_X1 U8712 ( .A1(n12514), .A2(n12768), .ZN(n12779) );
  NAND2_X1 U8713 ( .A1(n6918), .A2(n9928), .ZN(n9945) );
  OR2_X1 U8714 ( .A1(n9885), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9903) );
  NAND2_X1 U8715 ( .A1(n7225), .A2(n9870), .ZN(n9885) );
  INV_X1 U8716 ( .A(n7225), .ZN(n9871) );
  NAND2_X1 U8717 ( .A1(n7226), .A2(n6922), .ZN(n9857) );
  AND2_X1 U8718 ( .A1(n6488), .A2(n6923), .ZN(n6922) );
  INV_X1 U8719 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U8720 ( .A1(n7226), .A2(n6488), .ZN(n9842) );
  NAND2_X1 U8721 ( .A1(n7226), .A2(n9807), .ZN(n9824) );
  INV_X1 U8722 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n6925) );
  INV_X1 U8723 ( .A(n7226), .ZN(n9808) );
  NAND2_X1 U8724 ( .A1(n9742), .A2(n9741), .ZN(n9758) );
  NAND2_X1 U8725 ( .A1(n9742), .A2(n6926), .ZN(n9775) );
  NAND2_X1 U8726 ( .A1(n7224), .A2(n11514), .ZN(n9743) );
  OR2_X1 U8727 ( .A1(n9686), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9705) );
  INV_X1 U8728 ( .A(n7224), .ZN(n9722) );
  NAND2_X1 U8729 ( .A1(n11092), .A2(n7209), .ZN(n11091) );
  CLKBUF_X1 U8730 ( .A(n12524), .Z(n7209) );
  NAND2_X1 U8731 ( .A1(n7413), .A2(n12424), .ZN(n7412) );
  NAND2_X1 U8732 ( .A1(n9535), .A2(n10657), .ZN(n9576) );
  NOR2_X1 U8733 ( .A1(n12755), .A2(n12754), .ZN(n12993) );
  NOR2_X1 U8734 ( .A1(n12772), .A2(n9982), .ZN(n7072) );
  AND2_X1 U8735 ( .A1(n13001), .A2(n12565), .ZN(n9982) );
  NOR2_X1 U8736 ( .A1(n12374), .A2(n12754), .ZN(n10020) );
  NAND2_X1 U8737 ( .A1(n12795), .A2(n12981), .ZN(n7230) );
  NAND2_X1 U8738 ( .A1(n7203), .A2(n12801), .ZN(n12809) );
  AND2_X1 U8739 ( .A1(n9922), .A2(n12806), .ZN(n7204) );
  NAND2_X1 U8740 ( .A1(n11767), .A2(n12471), .ZN(n12910) );
  AND2_X1 U8741 ( .A1(n6509), .A2(n12457), .ZN(n12536) );
  INV_X1 U8742 ( .A(n7083), .ZN(n7082) );
  NOR2_X1 U8743 ( .A1(n9712), .A2(n7084), .ZN(n7083) );
  INV_X1 U8744 ( .A(n10121), .ZN(n10530) );
  AOI21_X1 U8745 ( .B1(n7702), .B2(n7704), .A(n6648), .ZN(n7700) );
  NAND2_X1 U8746 ( .A1(n7137), .A2(n7206), .ZN(n7205) );
  OAI21_X1 U8747 ( .B1(n6713), .B2(n13074), .A(P3_IR_REG_28__SCAN_IN), .ZN(
        n6712) );
  INV_X1 U8748 ( .A(n9493), .ZN(n6713) );
  NAND2_X1 U8749 ( .A1(n10042), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7119) );
  NAND2_X1 U8750 ( .A1(n10004), .A2(n7849), .ZN(n10022) );
  NOR2_X1 U8751 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n7849) );
  OR2_X1 U8752 ( .A1(n9786), .A2(P3_IR_REG_15__SCAN_IN), .ZN(n9788) );
  INV_X1 U8753 ( .A(n9767), .ZN(n7735) );
  OR2_X1 U8754 ( .A1(n9714), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U8755 ( .A1(n9639), .A2(n9640), .ZN(n10000) );
  INV_X1 U8756 ( .A(n9818), .ZN(n9661) );
  INV_X1 U8757 ( .A(n7721), .ZN(n7720) );
  AOI21_X1 U8758 ( .B1(n7719), .B2(n7721), .A(n7718), .ZN(n7717) );
  INV_X1 U8759 ( .A(n9634), .ZN(n7718) );
  XNOR2_X1 U8760 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n9525) );
  NAND2_X1 U8761 ( .A1(n9494), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n9523) );
  INV_X1 U8762 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8198) );
  OR2_X1 U8763 ( .A1(n13231), .A2(n13232), .ZN(n7483) );
  INV_X1 U8764 ( .A(n8394), .ZN(n6685) );
  INV_X1 U8765 ( .A(n7163), .ZN(n8453) );
  AND2_X1 U8766 ( .A1(n13190), .A2(n10718), .ZN(n6838) );
  INV_X1 U8767 ( .A(n11968), .ZN(n7499) );
  OR2_X1 U8768 ( .A1(n11043), .A2(n11044), .ZN(n13188) );
  NAND2_X1 U8769 ( .A1(n8178), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8199) );
  INV_X1 U8770 ( .A(n8180), .ZN(n8178) );
  NAND2_X1 U8771 ( .A1(n8216), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8242) );
  INV_X1 U8772 ( .A(n8218), .ZN(n8216) );
  AND2_X1 U8773 ( .A1(n12179), .A2(n11952), .ZN(n11953) );
  NAND2_X1 U8774 ( .A1(n7504), .A2(n11665), .ZN(n11954) );
  NAND2_X1 U8775 ( .A1(n8112), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n8131) );
  INV_X1 U8776 ( .A(n8114), .ZN(n8112) );
  AND2_X1 U8777 ( .A1(n7488), .A2(n7012), .ZN(n7011) );
  NAND2_X1 U8778 ( .A1(n12010), .A2(n13162), .ZN(n7012) );
  AND2_X1 U8779 ( .A1(n13267), .A2(n12012), .ZN(n7488) );
  XNOR2_X1 U8780 ( .A(n13866), .B(n13139), .ZN(n12062) );
  NAND2_X1 U8781 ( .A1(n13104), .A2(n11972), .ZN(n12064) );
  AND2_X1 U8782 ( .A1(n8542), .A2(n8541), .ZN(n13466) );
  OR2_X1 U8783 ( .A1(n13741), .A2(n8595), .ZN(n8502) );
  AND2_X1 U8784 ( .A1(n8460), .A2(n8459), .ZN(n13426) );
  AND2_X1 U8785 ( .A1(n8374), .A2(n8373), .ZN(n13409) );
  AND2_X1 U8786 ( .A1(n8334), .A2(n8333), .ZN(n13397) );
  AND3_X1 U8787 ( .A1(n8307), .A2(n8306), .A3(n8305), .ZN(n13392) );
  AND3_X1 U8788 ( .A1(n8246), .A2(n8245), .A3(n8244), .ZN(n13372) );
  AND4_X1 U8789 ( .A1(n8204), .A2(n8203), .A3(n8202), .A4(n8201), .ZN(n13358)
         );
  AND4_X1 U8790 ( .A1(n8137), .A2(n8136), .A3(n8135), .A4(n8134), .ZN(n13343)
         );
  OR2_X1 U8791 ( .A1(n8077), .A2(n8033), .ZN(n8038) );
  NAND2_X1 U8792 ( .A1(n7994), .A2(n6478), .ZN(n6947) );
  NAND2_X1 U8793 ( .A1(n15372), .A2(n10302), .ZN(n15376) );
  NAND2_X1 U8794 ( .A1(n10344), .A2(n10345), .ZN(n10343) );
  AND2_X1 U8795 ( .A1(n10946), .A2(n10945), .ZN(n15421) );
  NOR2_X1 U8796 ( .A1(n7451), .A2(n7447), .ZN(n7446) );
  INV_X1 U8797 ( .A(n10370), .ZN(n7451) );
  INV_X1 U8798 ( .A(n7449), .ZN(n7447) );
  AND2_X1 U8799 ( .A1(n11751), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7444) );
  OR2_X1 U8800 ( .A1(n15449), .A2(n15450), .ZN(n15446) );
  AND2_X1 U8801 ( .A1(n13649), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7442) );
  AND2_X1 U8802 ( .A1(n15462), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n15459) );
  NOR2_X1 U8803 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n8389) );
  AND2_X1 U8804 ( .A1(n6774), .A2(n6603), .ZN(n6773) );
  INV_X1 U8805 ( .A(n7160), .ZN(n8548) );
  NAND2_X1 U8806 ( .A1(n7390), .A2(n6551), .ZN(n6944) );
  AND2_X1 U8807 ( .A1(n6777), .A2(n7931), .ZN(n6776) );
  AOI21_X1 U8808 ( .B1(n7933), .B2(n7935), .A(n7932), .ZN(n7931) );
  INV_X1 U8809 ( .A(n13562), .ZN(n13697) );
  NAND2_X1 U8810 ( .A1(n7201), .A2(n13559), .ZN(n7200) );
  INV_X1 U8811 ( .A(n13717), .ZN(n7201) );
  NAND2_X1 U8812 ( .A1(n13720), .A2(n13880), .ZN(n7198) );
  NAND2_X1 U8813 ( .A1(n13719), .A2(n13878), .ZN(n7197) );
  NAND2_X1 U8814 ( .A1(n6687), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8535) );
  NAND2_X1 U8815 ( .A1(n7163), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n8480) );
  INV_X1 U8816 ( .A(n6687), .ZN(n8495) );
  NOR2_X1 U8817 ( .A1(n14058), .A2(n7769), .ZN(n6878) );
  NAND2_X1 U8818 ( .A1(n7386), .A2(n7387), .ZN(n7385) );
  AND3_X1 U8819 ( .A1(n14070), .A2(n13842), .A3(n13883), .ZN(n6877) );
  OR2_X1 U8820 ( .A1(n13829), .A2(n13858), .ZN(n13860) );
  NAND2_X1 U8821 ( .A1(n13883), .A2(n8688), .ZN(n13884) );
  OR2_X1 U8822 ( .A1(n14085), .A2(n7768), .ZN(n13900) );
  NAND2_X1 U8823 ( .A1(n7928), .A2(n11808), .ZN(n11812) );
  NAND2_X1 U8824 ( .A1(n11583), .A2(n7767), .ZN(n11733) );
  NAND2_X1 U8825 ( .A1(n11583), .A2(n11614), .ZN(n11719) );
  NAND2_X1 U8826 ( .A1(n8130), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8156) );
  INV_X1 U8827 ( .A(n8131), .ZN(n8130) );
  NAND2_X1 U8828 ( .A1(n8154), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n8180) );
  INV_X1 U8829 ( .A(n8156), .ZN(n8154) );
  AND2_X1 U8830 ( .A1(n11366), .A2(n11364), .ZN(n11583) );
  NOR2_X1 U8831 ( .A1(n11207), .A2(n14036), .ZN(n6883) );
  INV_X1 U8832 ( .A(n6886), .ZN(n6884) );
  NAND2_X1 U8833 ( .A1(n11003), .A2(n11002), .ZN(n11005) );
  NAND2_X1 U8834 ( .A1(n11192), .A2(n11191), .ZN(n11321) );
  NAND2_X1 U8835 ( .A1(n10108), .A2(n8065), .ZN(n11006) );
  NAND2_X1 U8836 ( .A1(n6887), .A2(n6888), .ZN(n11010) );
  INV_X1 U8837 ( .A(n11207), .ZN(n6887) );
  INV_X1 U8838 ( .A(n13878), .ZN(n13273) );
  NAND2_X1 U8839 ( .A1(n13612), .A2(n13296), .ZN(n12142) );
  INV_X1 U8840 ( .A(n13541), .ZN(n12151) );
  NOR2_X1 U8841 ( .A1(n13916), .A2(n13296), .ZN(n12147) );
  NOR2_X1 U8842 ( .A1(n13675), .A2(n7771), .ZN(n7770) );
  NAND2_X1 U8843 ( .A1(n7772), .A2(n13694), .ZN(n7771) );
  INV_X1 U8844 ( .A(n7773), .ZN(n7772) );
  AND2_X1 U8845 ( .A1(n8808), .A2(n13460), .ZN(n6882) );
  NOR2_X1 U8846 ( .A1(n13939), .A2(n7189), .ZN(n7188) );
  AND2_X1 U8847 ( .A1(n13940), .A2(n15524), .ZN(n7189) );
  NAND2_X1 U8848 ( .A1(n10113), .A2(n10114), .ZN(n10112) );
  OR2_X1 U8849 ( .A1(n7678), .A2(n8652), .ZN(n10114) );
  AND3_X1 U8850 ( .A1(n15508), .A2(n10562), .A3(n8701), .ZN(n8810) );
  AND2_X1 U8851 ( .A1(n13294), .A2(n13284), .ZN(n10884) );
  OR2_X1 U8852 ( .A1(n8149), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U8853 ( .A1(n7218), .A2(n7998), .ZN(n8048) );
  INV_X1 U8854 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9494) );
  NAND2_X1 U8855 ( .A1(n8857), .A2(n8856), .ZN(n9443) );
  INV_X1 U8856 ( .A(n8855), .ZN(n8857) );
  AND2_X1 U8857 ( .A1(n14261), .A2(n7569), .ZN(n7568) );
  OR2_X1 U8858 ( .A1(n14179), .A2(n7570), .ZN(n7569) );
  INV_X1 U8859 ( .A(n9366), .ZN(n7570) );
  NAND2_X1 U8860 ( .A1(n9231), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9246) );
  NAND2_X1 U8861 ( .A1(n15018), .A2(n8888), .ZN(n9418) );
  NOR2_X1 U8862 ( .A1(n11568), .A2(n7560), .ZN(n7559) );
  INV_X1 U8863 ( .A(n7563), .ZN(n7560) );
  OR2_X1 U8864 ( .A1(n9033), .A2(n9034), .ZN(n7563) );
  NAND2_X1 U8865 ( .A1(n7562), .A2(n7564), .ZN(n7561) );
  INV_X1 U8866 ( .A(n14104), .ZN(n7562) );
  NAND2_X1 U8867 ( .A1(n11864), .A2(n9119), .ZN(n14168) );
  NAND2_X1 U8868 ( .A1(n9184), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9187) );
  NAND2_X1 U8869 ( .A1(n9231), .A2(n7275), .ZN(n9257) );
  INV_X1 U8870 ( .A(n14251), .ZN(n6996) );
  INV_X1 U8871 ( .A(n6998), .ZN(n6997) );
  NAND2_X1 U8872 ( .A1(n8863), .A2(n7273), .ZN(n9165) );
  NAND2_X1 U8873 ( .A1(n8863), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9142) );
  INV_X1 U8874 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n11311) );
  NOR2_X1 U8875 ( .A1(n9301), .A2(n12036), .ZN(n7001) );
  OR2_X1 U8876 ( .A1(n9155), .A2(n14229), .ZN(n7585) );
  INV_X1 U8877 ( .A(n9119), .ZN(n7584) );
  NAND2_X1 U8878 ( .A1(n8862), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n9125) );
  INV_X1 U8879 ( .A(n9106), .ZN(n8862) );
  XNOR2_X1 U8880 ( .A(n8938), .B(n9380), .ZN(n8953) );
  NOR2_X1 U8881 ( .A1(n6523), .A2(n7556), .ZN(n7555) );
  INV_X1 U8882 ( .A(n11079), .ZN(n7556) );
  INV_X1 U8883 ( .A(n9418), .ZN(n9324) );
  AND2_X1 U8884 ( .A1(n14122), .A2(n9178), .ZN(n14189) );
  OR2_X1 U8885 ( .A1(n6437), .A2(n10611), .ZN(n8882) );
  INV_X1 U8886 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14591) );
  INV_X1 U8887 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14664) );
  NAND2_X1 U8888 ( .A1(n6689), .A2(n6688), .ZN(n11372) );
  INV_X1 U8889 ( .A(n11304), .ZN(n6688) );
  INV_X1 U8890 ( .A(n11303), .ZN(n6689) );
  XNOR2_X1 U8891 ( .A(n11901), .B(n11908), .ZN(n11899) );
  OR2_X1 U8892 ( .A1(n11905), .A2(n11906), .ZN(n14687) );
  OR2_X1 U8893 ( .A1(n11913), .A2(n11914), .ZN(n14696) );
  OR2_X1 U8894 ( .A1(n14711), .A2(n14712), .ZN(n14729) );
  OR2_X1 U8895 ( .A1(n14783), .A2(n14758), .ZN(n14759) );
  NOR2_X1 U8896 ( .A1(n14759), .A2(n14499), .ZN(n14744) );
  INV_X1 U8897 ( .A(n14797), .ZN(n7546) );
  INV_X1 U8898 ( .A(n7791), .ZN(n7785) );
  INV_X1 U8899 ( .A(n14751), .ZN(n7784) );
  NAND2_X1 U8900 ( .A1(n14803), .A2(n15046), .ZN(n14783) );
  AND2_X1 U8901 ( .A1(n14836), .A2(n7468), .ZN(n14803) );
  AND2_X1 U8902 ( .A1(n7469), .A2(n7795), .ZN(n7468) );
  NAND2_X1 U8903 ( .A1(n7796), .A2(n15010), .ZN(n12116) );
  AND2_X1 U8904 ( .A1(n14871), .A2(n14859), .ZN(n14836) );
  NAND2_X1 U8905 ( .A1(n14836), .A2(n14843), .ZN(n14837) );
  AND2_X1 U8906 ( .A1(n9300), .A2(n9299), .ZN(n14852) );
  AND2_X1 U8907 ( .A1(n14934), .A2(n7465), .ZN(n14871) );
  AND2_X1 U8908 ( .A1(n6465), .A2(n14877), .ZN(n7465) );
  AND2_X1 U8909 ( .A1(n7275), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n7274) );
  NAND2_X1 U8910 ( .A1(n14934), .A2(n6465), .ZN(n14889) );
  NAND2_X1 U8911 ( .A1(n7551), .A2(n12131), .ZN(n14883) );
  AND2_X1 U8912 ( .A1(n14934), .A2(n14921), .ZN(n14915) );
  NAND2_X1 U8913 ( .A1(n7782), .A2(n14386), .ZN(n14965) );
  INV_X1 U8914 ( .A(n14987), .ZN(n14998) );
  NAND2_X1 U8915 ( .A1(n15014), .A2(n7458), .ZN(n7461) );
  NOR2_X1 U8916 ( .A1(n7462), .A2(n15130), .ZN(n7458) );
  NAND2_X1 U8917 ( .A1(n7460), .A2(n7459), .ZN(n15017) );
  NOR2_X1 U8918 ( .A1(n15136), .A2(n7462), .ZN(n7460) );
  NOR2_X1 U8919 ( .A1(n7953), .A2(n7462), .ZN(n15015) );
  NOR2_X1 U8920 ( .A1(n7953), .A2(n15149), .ZN(n11923) );
  OAI21_X1 U8921 ( .B1(n11849), .B2(n6508), .A(n11848), .ZN(n11850) );
  OR2_X1 U8922 ( .A1(n11850), .A2(n11844), .ZN(n11921) );
  OR2_X1 U8923 ( .A1(n9061), .A2(n9060), .ZN(n9077) );
  OR2_X1 U8924 ( .A1(n9077), .A2(n9076), .ZN(n9106) );
  NAND2_X1 U8925 ( .A1(n7272), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9039) );
  NAND2_X1 U8926 ( .A1(n8861), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9024) );
  NOR2_X1 U8927 ( .A1(n6553), .A2(n6723), .ZN(n6722) );
  INV_X1 U8928 ( .A(n14313), .ZN(n11345) );
  NAND2_X1 U8929 ( .A1(n11051), .A2(n11058), .ZN(n11139) );
  AND2_X1 U8930 ( .A1(n11029), .A2(n15293), .ZN(n11051) );
  CLKBUF_X1 U8931 ( .A(n14502), .Z(n15256) );
  INV_X1 U8932 ( .A(n14557), .ZN(n14298) );
  AND2_X1 U8933 ( .A1(n10245), .A2(n14571), .ZN(n15008) );
  INV_X1 U8934 ( .A(n15010), .ZN(n14855) );
  NAND2_X1 U8935 ( .A1(n15264), .A2(n14526), .ZN(n15018) );
  INV_X1 U8936 ( .A(n15296), .ZN(n15311) );
  INV_X1 U8937 ( .A(n15264), .ZN(n15280) );
  INV_X1 U8938 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n15781) );
  NOR2_X1 U8939 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), .ZN(
        n7463) );
  NAND2_X1 U8940 ( .A1(n7889), .A2(n7890), .ZN(n8560) );
  NAND2_X1 U8941 ( .A1(n8544), .A2(n7891), .ZN(n7889) );
  NAND2_X1 U8942 ( .A1(n7954), .A2(n7510), .ZN(n7781) );
  XNOR2_X1 U8943 ( .A(n8449), .B(n8448), .ZN(n9289) );
  NAND2_X1 U8944 ( .A1(n7588), .A2(n6466), .ZN(n8852) );
  NAND2_X1 U8945 ( .A1(n8359), .A2(n8358), .ZN(n8380) );
  NAND2_X1 U8946 ( .A1(n9057), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9101) );
  OR2_X1 U8947 ( .A1(n9056), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n9057) );
  OR2_X1 U8948 ( .A1(n9019), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n9056) );
  OR2_X1 U8949 ( .A1(n8984), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U8950 ( .A1(n8104), .A2(n8105), .ZN(n6991) );
  OR2_X1 U8951 ( .A1(n8944), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8963) );
  NAND2_X1 U8952 ( .A1(n8829), .A2(n8828), .ZN(n8984) );
  INV_X1 U8953 ( .A(n8963), .ZN(n8829) );
  INV_X1 U8954 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n8743) );
  NAND2_X1 U8955 ( .A1(n7638), .A2(n7636), .ZN(n8740) );
  NAND2_X1 U8956 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n7637), .ZN(n7636) );
  INV_X1 U8957 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n7637) );
  XNOR2_X1 U8958 ( .A(n8749), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n8750) );
  AND2_X1 U8959 ( .A1(n8765), .A2(n6834), .ZN(n6833) );
  NAND2_X1 U8960 ( .A1(n7115), .A2(n6449), .ZN(n11825) );
  NAND2_X1 U8961 ( .A1(n11671), .A2(n7868), .ZN(n7115) );
  AND2_X1 U8962 ( .A1(n9921), .A2(n9920), .ZN(n12839) );
  NAND2_X1 U8963 ( .A1(n10916), .A2(n10915), .ZN(n11424) );
  NAND2_X1 U8964 ( .A1(n7101), .A2(n7105), .ZN(n12242) );
  NAND2_X1 U8965 ( .A1(n7101), .A2(n7099), .ZN(n12243) );
  XNOR2_X1 U8966 ( .A(n10869), .B(n12578), .ZN(n11290) );
  INV_X1 U8967 ( .A(n7808), .ZN(n12399) );
  NAND2_X1 U8968 ( .A1(n12309), .A2(n12216), .ZN(n12260) );
  INV_X1 U8969 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11514) );
  AOI21_X1 U8970 ( .B1(n10779), .B2(n9956), .A(n9792), .ZN(n12286) );
  AOI21_X1 U8971 ( .B1(n12299), .B2(n12821), .A(n7157), .ZN(n12302) );
  NAND2_X1 U8972 ( .A1(n10652), .A2(n10651), .ZN(n10863) );
  NAND2_X1 U8973 ( .A1(n12311), .A2(n12310), .ZN(n12309) );
  AOI21_X1 U8974 ( .B1(n7854), .B2(n7853), .A(n6636), .ZN(n7852) );
  INV_X1 U8975 ( .A(n12310), .ZN(n7853) );
  NAND2_X1 U8976 ( .A1(n7104), .A2(n7109), .ZN(n12331) );
  OR2_X1 U8977 ( .A1(n12288), .A2(n12287), .ZN(n7104) );
  AND2_X1 U8978 ( .A1(n9968), .A2(n9967), .ZN(n12345) );
  INV_X1 U8979 ( .A(n12347), .ZN(n12285) );
  OAI21_X1 U8980 ( .B1(n11671), .B2(n7114), .A(n7113), .ZN(n11828) );
  INV_X1 U8981 ( .A(n12349), .ZN(n12308) );
  NAND2_X1 U8982 ( .A1(n10538), .A2(n10537), .ZN(n12340) );
  NAND2_X1 U8983 ( .A1(n6673), .A2(n6671), .ZN(n12555) );
  INV_X1 U8984 ( .A(n6672), .ZN(n6671) );
  OAI21_X1 U8985 ( .B1(n12553), .B2(n12552), .A(n12551), .ZN(n6672) );
  INV_X1 U8986 ( .A(n12345), .ZN(n12795) );
  INV_X1 U8987 ( .A(n12839), .ZN(n12567) );
  INV_X1 U8988 ( .A(n12821), .ZN(n12568) );
  OR2_X1 U8989 ( .A1(n10531), .A2(n13072), .ZN(n12571) );
  OR2_X1 U8990 ( .A1(n9596), .A2(n9623), .ZN(n9631) );
  OR2_X1 U8991 ( .A1(n10015), .A2(n9560), .ZN(n9566) );
  OR2_X1 U8992 ( .A1(n9596), .A2(n9578), .ZN(n9579) );
  OR2_X1 U8993 ( .A1(n10015), .A2(n9516), .ZN(n9521) );
  NAND2_X1 U8994 ( .A1(n10515), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n10514) );
  OAI21_X1 U8995 ( .B1(n10664), .B2(n7598), .A(n7596), .ZN(n10445) );
  NAND2_X1 U8996 ( .A1(n10689), .A2(n10688), .ZN(n15552) );
  NAND2_X1 U8997 ( .A1(n6976), .A2(n11234), .ZN(n11697) );
  NAND2_X1 U8998 ( .A1(n15564), .A2(n15565), .ZN(n6976) );
  NAND2_X1 U8999 ( .A1(n7611), .A2(n7610), .ZN(n7612) );
  OR2_X1 U9000 ( .A1(n15584), .A2(n11271), .ZN(n7610) );
  NAND2_X1 U9001 ( .A1(n6972), .A2(n6971), .ZN(n15594) );
  NAND2_X1 U9002 ( .A1(n6974), .A2(n6973), .ZN(n6972) );
  NAND2_X1 U9003 ( .A1(n12588), .A2(n12586), .ZN(n7604) );
  NOR2_X1 U9004 ( .A1(n12630), .A2(n6901), .ZN(n12613) );
  NAND2_X1 U9005 ( .A1(n7599), .A2(n7600), .ZN(n6901) );
  NAND2_X1 U9006 ( .A1(n12615), .A2(n6985), .ZN(n12618) );
  NAND2_X1 U9007 ( .A1(n12632), .A2(n12631), .ZN(n7589) );
  AOI21_X1 U9008 ( .B1(n6982), .B2(n6980), .A(n6594), .ZN(n6979) );
  INV_X1 U9009 ( .A(n6982), .ZN(n6981) );
  NAND2_X1 U9010 ( .A1(n12648), .A2(n12647), .ZN(n12660) );
  NAND2_X1 U9011 ( .A1(n12640), .A2(n12639), .ZN(n12654) );
  NOR2_X1 U9012 ( .A1(n6893), .A2(n12677), .ZN(n12678) );
  NAND2_X1 U9013 ( .A1(n6894), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n6893) );
  NOR2_X1 U9014 ( .A1(n7591), .A2(n12677), .ZN(n12655) );
  NAND2_X1 U9015 ( .A1(n12675), .A2(n12674), .ZN(n12693) );
  INV_X1 U9016 ( .A(n7367), .ZN(n12700) );
  XNOR2_X1 U9017 ( .A(n12712), .B(n12713), .ZN(n12714) );
  OR2_X1 U9018 ( .A1(n10125), .A2(n10123), .ZN(n15570) );
  XNOR2_X1 U9019 ( .A(n7052), .B(n7051), .ZN(n12750) );
  INV_X1 U9020 ( .A(n12749), .ZN(n7051) );
  OAI21_X1 U9021 ( .B1(n12712), .B2(n7044), .A(n7042), .ZN(n7052) );
  INV_X1 U9022 ( .A(n7046), .ZN(n7044) );
  NAND2_X1 U9023 ( .A1(n9927), .A2(n9926), .ZN(n12803) );
  NOR2_X1 U9024 ( .A1(n12843), .A2(n7418), .ZN(n7417) );
  INV_X1 U9025 ( .A(n7420), .ZN(n7418) );
  NAND2_X1 U9026 ( .A1(n7419), .A2(n7420), .ZN(n12844) );
  NAND2_X1 U9027 ( .A1(n7817), .A2(n7821), .ZN(n11768) );
  NAND2_X1 U9028 ( .A1(n11591), .A2(n7824), .ZN(n7817) );
  NAND2_X1 U9029 ( .A1(n7414), .A2(n6693), .ZN(n10976) );
  AOI21_X1 U9030 ( .B1(n10782), .B2(n10783), .A(n12411), .ZN(n10772) );
  INV_X1 U9031 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n9535) );
  XNOR2_X1 U9032 ( .A(n7055), .B(n12979), .ZN(n12987) );
  INV_X1 U9033 ( .A(n15616), .ZN(n15618) );
  INV_X1 U9034 ( .A(n12968), .ZN(n12976) );
  NAND2_X1 U9035 ( .A1(n12359), .A2(n12358), .ZN(n12375) );
  NAND2_X1 U9036 ( .A1(n12935), .A2(n7407), .ZN(n13005) );
  AND2_X1 U9037 ( .A1(n12932), .A2(n12933), .ZN(n7408) );
  NAND2_X1 U9038 ( .A1(n9944), .A2(n9943), .ZN(n13008) );
  AOI21_X1 U9039 ( .B1(n7231), .B2(n12986), .A(n7228), .ZN(n13006) );
  NAND2_X1 U9040 ( .A1(n7230), .A2(n7229), .ZN(n7228) );
  XNOR2_X1 U9041 ( .A(n12794), .B(n12793), .ZN(n7231) );
  NAND2_X1 U9042 ( .A1(n12796), .A2(n12982), .ZN(n7229) );
  INV_X1 U9043 ( .A(n12803), .ZN(n13012) );
  INV_X1 U9044 ( .A(n12941), .ZN(n13020) );
  NAND2_X1 U9045 ( .A1(n9884), .A2(n9883), .ZN(n13027) );
  NAND2_X1 U9046 ( .A1(n7073), .A2(n7076), .ZN(n12856) );
  OR2_X1 U9047 ( .A1(n12877), .A2(n7077), .ZN(n7073) );
  NAND2_X1 U9048 ( .A1(n7421), .A2(n12490), .ZN(n12853) );
  NAND2_X1 U9049 ( .A1(n12862), .A2(n12491), .ZN(n7421) );
  NAND2_X1 U9050 ( .A1(n12875), .A2(n9864), .ZN(n12865) );
  AND2_X1 U9051 ( .A1(n12879), .A2(n12878), .ZN(n13037) );
  NAND2_X1 U9052 ( .A1(n7815), .A2(n7814), .ZN(n12871) );
  AND2_X1 U9053 ( .A1(n7815), .A2(n6528), .ZN(n12873) );
  NAND2_X1 U9054 ( .A1(n12891), .A2(n7816), .ZN(n7815) );
  AOI21_X1 U9055 ( .B1(n11165), .B2(n9956), .A(n9841), .ZN(n13044) );
  NOR2_X1 U9056 ( .A1(n6520), .A2(n10079), .ZN(n12883) );
  NAND2_X1 U9057 ( .A1(n9823), .A2(n9822), .ZN(n13050) );
  NAND2_X1 U9058 ( .A1(n7649), .A2(n7059), .ZN(n7057) );
  NAND2_X1 U9059 ( .A1(n7649), .A2(n7063), .ZN(n12902) );
  NAND2_X1 U9060 ( .A1(n11765), .A2(n7650), .ZN(n7063) );
  NAND2_X1 U9061 ( .A1(n11763), .A2(n9780), .ZN(n12915) );
  OAI21_X1 U9062 ( .B1(n11591), .B2(n7826), .A(n12457), .ZN(n11774) );
  NAND2_X1 U9063 ( .A1(n9740), .A2(n9739), .ZN(n11644) );
  NAND2_X1 U9064 ( .A1(n9721), .A2(n9720), .ZN(n11520) );
  OAI21_X1 U9065 ( .B1(n7837), .B2(n11265), .A(n7836), .ZN(n11437) );
  INV_X1 U9066 ( .A(n7841), .ZN(n7837) );
  AOI21_X1 U9067 ( .B1(n7841), .B2(n7840), .A(n7839), .ZN(n7836) );
  NAND2_X1 U9068 ( .A1(n7085), .A2(n9693), .ZN(n11337) );
  NAND2_X1 U9069 ( .A1(n11249), .A2(n12534), .ZN(n7085) );
  NAND2_X1 U9070 ( .A1(n7843), .A2(n7844), .ZN(n11339) );
  NAND2_X1 U9071 ( .A1(n11265), .A2(n7846), .ZN(n7843) );
  AOI21_X1 U9072 ( .B1(n11265), .B2(n12439), .A(n7848), .ZN(n11251) );
  AND2_X1 U9073 ( .A1(n15654), .A2(n12933), .ZN(n13061) );
  NAND2_X1 U9074 ( .A1(n9529), .A2(n10142), .ZN(n9513) );
  AND2_X1 U9075 ( .A1(n10530), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10163) );
  NAND2_X1 U9076 ( .A1(n7089), .A2(n6525), .ZN(n10044) );
  INV_X1 U9077 ( .A(n10163), .ZN(n13072) );
  NOR2_X1 U9078 ( .A1(P3_IR_REG_28__SCAN_IN), .A2(n7669), .ZN(n7668) );
  NAND2_X1 U9079 ( .A1(n9502), .A2(n7206), .ZN(n7669) );
  XNOR2_X1 U9080 ( .A(n12354), .B(n11936), .ZN(n12367) );
  XNOR2_X1 U9081 ( .A(n11934), .B(n9988), .ZN(n12198) );
  NAND2_X1 U9082 ( .A1(n7701), .A2(n9955), .ZN(n9972) );
  NAND2_X1 U9083 ( .A1(n9954), .A2(n9953), .ZN(n7701) );
  INV_X1 U9084 ( .A(n10048), .ZN(n10037) );
  OAI21_X1 U9085 ( .B1(n7756), .B2(n7752), .A(n7753), .ZN(n9925) );
  NAND2_X1 U9086 ( .A1(n9900), .A2(n9899), .ZN(n9913) );
  NAND2_X1 U9087 ( .A1(n7756), .A2(n9893), .ZN(n9900) );
  NAND2_X1 U9088 ( .A1(n7709), .A2(n7710), .ZN(n9880) );
  OR2_X1 U9089 ( .A1(n9853), .A2(n7713), .ZN(n7709) );
  INV_X1 U9090 ( .A(n10097), .ZN(n11334) );
  OAI21_X1 U9091 ( .B1(n9853), .B2(n7716), .A(n9852), .ZN(n9866) );
  INV_X1 U9092 ( .A(SI_18_), .ZN(n11103) );
  INV_X1 U9093 ( .A(SI_17_), .ZN(n10928) );
  NAND2_X1 U9094 ( .A1(n6792), .A2(n6796), .ZN(n9815) );
  NAND2_X1 U9095 ( .A1(n9766), .A2(n7729), .ZN(n6792) );
  INV_X1 U9096 ( .A(SI_16_), .ZN(n10780) );
  XNOR2_X1 U9097 ( .A(n9799), .B(n9798), .ZN(n10779) );
  NAND2_X1 U9098 ( .A1(n7728), .A2(n7731), .ZN(n9799) );
  NAND2_X1 U9099 ( .A1(n9766), .A2(n7734), .ZN(n7728) );
  NAND2_X1 U9100 ( .A1(n7736), .A2(n9767), .ZN(n9784) );
  INV_X1 U9101 ( .A(SI_15_), .ZN(n10637) );
  INV_X1 U9102 ( .A(SI_13_), .ZN(n10283) );
  INV_X1 U9103 ( .A(SI_12_), .ZN(n10233) );
  INV_X1 U9104 ( .A(SI_11_), .ZN(n10201) );
  NAND2_X1 U9105 ( .A1(n6800), .A2(n6803), .ZN(n9713) );
  NAND2_X1 U9106 ( .A1(n9680), .A2(n6806), .ZN(n6800) );
  NAND2_X1 U9107 ( .A1(n6808), .A2(n9678), .ZN(n9696) );
  NAND2_X1 U9108 ( .A1(n6809), .A2(n6810), .ZN(n6808) );
  NAND2_X1 U9109 ( .A1(n7723), .A2(n7721), .ZN(n9635) );
  NAND2_X1 U9110 ( .A1(n7723), .A2(n7726), .ZN(n9615) );
  NAND2_X1 U9111 ( .A1(n9568), .A2(n9552), .ZN(n9612) );
  NAND2_X1 U9112 ( .A1(n7743), .A2(n7742), .ZN(n9586) );
  NAND2_X1 U9113 ( .A1(n7743), .A2(n9547), .ZN(n9584) );
  NAND2_X1 U9114 ( .A1(n9546), .A2(n9545), .ZN(n9599) );
  NOR2_X1 U9115 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_2__SCAN_IN), .ZN(
        n7053) );
  NOR2_X1 U9116 ( .A1(n13074), .A2(n9480), .ZN(n7054) );
  MUX2_X1 U9117 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9495), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n9496) );
  OR2_X1 U9118 ( .A1(n10723), .A2(n10724), .ZN(n10299) );
  AND3_X1 U9119 ( .A1(n8271), .A2(n8270), .A3(n8269), .ZN(n13552) );
  INV_X1 U9120 ( .A(n13204), .ZN(n11988) );
  AND2_X1 U9121 ( .A1(n8357), .A2(n8356), .ZN(n13126) );
  NAND2_X1 U9122 ( .A1(n13188), .A2(n6838), .ZN(n13187) );
  AND2_X1 U9123 ( .A1(n11962), .A2(n6840), .ZN(n6839) );
  INV_X1 U9124 ( .A(n13214), .ZN(n6840) );
  INV_X1 U9125 ( .A(n7501), .ZN(n7500) );
  OR2_X1 U9126 ( .A1(n13180), .A2(n6521), .ZN(n7356) );
  OAI21_X1 U9127 ( .B1(n13218), .B2(n12002), .A(n6521), .ZN(n7480) );
  NAND2_X1 U9128 ( .A1(n6835), .A2(n12166), .ZN(n12171) );
  NAND2_X1 U9129 ( .A1(n12197), .A2(n11660), .ZN(n6835) );
  NAND2_X1 U9130 ( .A1(n12090), .A2(n11962), .ZN(n13213) );
  INV_X1 U9131 ( .A(n13277), .ZN(n13261) );
  NAND2_X1 U9132 ( .A1(n11954), .A2(n11953), .ZN(n12184) );
  NAND2_X1 U9133 ( .A1(n7014), .A2(n7494), .ZN(n13252) );
  AOI21_X1 U9134 ( .B1(n13179), .B2(n13162), .A(n6841), .ZN(n13264) );
  NAND2_X1 U9135 ( .A1(n7011), .A2(n13270), .ZN(n6841) );
  NOR2_X1 U9136 ( .A1(n13577), .A2(n13580), .ZN(n7148) );
  OR2_X1 U9137 ( .A1(n13143), .A2(n8595), .ZN(n8576) );
  NAND2_X1 U9138 ( .A1(n8555), .A2(n8554), .ZN(n13591) );
  INV_X1 U9139 ( .A(n13466), .ZN(n13720) );
  INV_X1 U9140 ( .A(n13475), .ZN(n13719) );
  INV_X1 U9141 ( .A(n13426), .ZN(n13594) );
  INV_X1 U9142 ( .A(n13397), .ZN(n13598) );
  OR2_X1 U9143 ( .A1(n8077), .A2(n8078), .ZN(n8082) );
  NAND2_X1 U9144 ( .A1(n13629), .A2(n10367), .ZN(n15408) );
  INV_X1 U9145 ( .A(n7436), .ZN(n15491) );
  INV_X1 U9146 ( .A(n7431), .ZN(n13660) );
  NAND2_X1 U9147 ( .A1(n8802), .A2(n8578), .ZN(n8803) );
  OR2_X1 U9148 ( .A1(n13698), .A2(n13697), .ZN(n13932) );
  OR2_X1 U9149 ( .A1(n7393), .A2(n7392), .ZN(n6945) );
  NAND2_X1 U9150 ( .A1(n7687), .A2(n7393), .ZN(n13715) );
  NAND2_X1 U9151 ( .A1(n7690), .A2(n7691), .ZN(n13734) );
  NAND2_X1 U9152 ( .A1(n7691), .A2(n13535), .ZN(n13732) );
  NAND2_X1 U9153 ( .A1(n11562), .A2(n8146), .ZN(n6657) );
  NAND2_X1 U9154 ( .A1(n7930), .A2(n8439), .ZN(n12050) );
  NAND2_X1 U9155 ( .A1(n13803), .A2(n8404), .ZN(n13780) );
  NAND2_X1 U9156 ( .A1(n7388), .A2(n7694), .ZN(n13778) );
  NAND2_X1 U9157 ( .A1(n6510), .A2(n8674), .ZN(n13795) );
  NAND2_X1 U9158 ( .A1(n6955), .A2(n6956), .ZN(n13864) );
  NAND2_X1 U9159 ( .A1(n6957), .A2(n6960), .ZN(n13890) );
  OR2_X1 U9160 ( .A1(n13906), .A2(n8668), .ZN(n6957) );
  NAND2_X1 U9161 ( .A1(n7686), .A2(n8665), .ZN(n11809) );
  NAND2_X1 U9162 ( .A1(n11728), .A2(n6407), .ZN(n7686) );
  NAND2_X1 U9163 ( .A1(n7023), .A2(n7025), .ZN(n11711) );
  INV_X1 U9164 ( .A(n7398), .ZN(n7964) );
  AOI21_X1 U9165 ( .B1(n7671), .B2(n7402), .A(n7401), .ZN(n7398) );
  NAND2_X1 U9166 ( .A1(n11188), .A2(n8102), .ZN(n11327) );
  NAND2_X1 U9167 ( .A1(n11003), .A2(n7380), .ZN(n6938) );
  INV_X1 U9168 ( .A(n13904), .ZN(n13917) );
  AND2_X1 U9169 ( .A1(n13913), .A2(n13568), .ZN(n13919) );
  INV_X1 U9170 ( .A(n13919), .ZN(n13744) );
  AND2_X1 U9171 ( .A1(n15538), .A2(n13927), .ZN(n7764) );
  INV_X1 U9172 ( .A(n15538), .ZN(n15536) );
  AND2_X1 U9173 ( .A1(n15533), .A2(n13927), .ZN(n7763) );
  NAND2_X1 U9174 ( .A1(n7190), .A2(n7186), .ZN(n14049) );
  INV_X1 U9175 ( .A(n7187), .ZN(n7186) );
  INV_X1 U9176 ( .A(n13938), .ZN(n7190) );
  OAI21_X1 U9177 ( .B1(n13941), .B2(n14040), .A(n7188), .ZN(n7187) );
  OR3_X1 U9178 ( .A1(n13992), .A2(n13991), .A3(n13990), .ZN(n14071) );
  NAND2_X1 U9179 ( .A1(n7397), .A2(n8146), .ZN(n7396) );
  INV_X1 U9180 ( .A(n10167), .ZN(n7397) );
  AND2_X1 U9181 ( .A1(n10723), .A2(n8636), .ZN(n15507) );
  AND2_X1 U9182 ( .A1(n8011), .A2(n7990), .ZN(n7948) );
  NAND2_X1 U9183 ( .A1(n7404), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7035) );
  NOR2_X1 U9184 ( .A1(n7674), .A2(n7673), .ZN(n7672) );
  NOR2_X1 U9185 ( .A1(n8009), .A2(n8008), .ZN(n7673) );
  INV_X1 U9186 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n15780) );
  XNOR2_X1 U9187 ( .A(n8627), .B(n8626), .ZN(n11624) );
  INV_X1 U9188 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U9189 ( .A1(n8624), .A2(n8625), .ZN(n11490) );
  NAND2_X1 U9190 ( .A1(n8619), .A2(n8620), .ZN(n11563) );
  INV_X1 U9191 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11509) );
  INV_X1 U9192 ( .A(n13672), .ZN(n13568) );
  INV_X1 U9193 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10900) );
  INV_X1 U9194 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10751) );
  INV_X1 U9195 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10830) );
  INV_X1 U9196 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10494) );
  INV_X1 U9197 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10500) );
  INV_X1 U9198 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10458) );
  XNOR2_X1 U9199 ( .A(n8194), .B(P2_IR_REG_10__SCAN_IN), .ZN(n15428) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10240) );
  INV_X1 U9201 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10235) );
  INV_X1 U9202 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10199) );
  INV_X1 U9203 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10177) );
  INV_X1 U9204 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10152) );
  OAI211_X1 U9205 ( .C1(P2_IR_REG_2__SCAN_IN), .C2(P2_IR_REG_31__SCAN_IN), .A(
        n7452), .B(n8048), .ZN(n10350) );
  NAND2_X1 U9206 ( .A1(n8047), .A2(n7453), .ZN(n7452) );
  NOR2_X1 U9207 ( .A1(n7989), .A2(n7998), .ZN(n7453) );
  INV_X1 U9208 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10153) );
  MUX2_X1 U9209 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8018), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8019) );
  AND2_X1 U9210 ( .A1(n9414), .A2(n9413), .ZN(n14794) );
  OR2_X1 U9211 ( .A1(n9465), .A2(n6439), .ZN(n9414) );
  NAND2_X1 U9212 ( .A1(n6511), .A2(n7583), .ZN(n14124) );
  AND2_X1 U9213 ( .A1(n14282), .A2(n15008), .ZN(n14264) );
  AND2_X1 U9214 ( .A1(n6999), .A2(n6526), .ZN(n14154) );
  NAND2_X1 U9215 ( .A1(n6999), .A2(n6998), .ZN(n14152) );
  NAND2_X1 U9216 ( .A1(n7561), .A2(n7563), .ZN(n11569) );
  NAND2_X1 U9217 ( .A1(n10290), .A2(n8921), .ZN(n10605) );
  NAND2_X1 U9218 ( .A1(n8896), .A2(n8922), .ZN(n10608) );
  NAND2_X1 U9219 ( .A1(n14221), .A2(n9270), .ZN(n14161) );
  INV_X1 U9220 ( .A(n14954), .ZN(n14384) );
  AND2_X1 U9221 ( .A1(n7583), .A2(n7585), .ZN(n14231) );
  NAND2_X1 U9222 ( .A1(n14159), .A2(n9288), .ZN(n14242) );
  OR2_X1 U9223 ( .A1(n9224), .A2(n9225), .ZN(n7581) );
  NAND2_X1 U9224 ( .A1(n7557), .A2(n11080), .ZN(n11159) );
  OR2_X1 U9225 ( .A1(n9451), .A2(n9447), .ZN(n14271) );
  AND2_X1 U9226 ( .A1(n14218), .A2(n15336), .ZN(n14269) );
  INV_X1 U9227 ( .A(n14271), .ZN(n14273) );
  INV_X1 U9228 ( .A(n14794), .ZN(n14761) );
  NAND2_X1 U9229 ( .A1(n9377), .A2(n9376), .ZN(n14753) );
  NAND2_X1 U9230 ( .A1(n9359), .A2(n9358), .ZN(n14833) );
  OR2_X1 U9231 ( .A1(n14181), .A2(n6439), .ZN(n9359) );
  NAND2_X1 U9232 ( .A1(n9340), .A2(n9339), .ZN(n14542) );
  NAND2_X1 U9233 ( .A1(n9320), .A2(n9319), .ZN(n14832) );
  OR2_X1 U9234 ( .A1(n14134), .A2(n6438), .ZN(n9320) );
  INV_X1 U9235 ( .A(n14852), .ZN(n14543) );
  NAND2_X1 U9236 ( .A1(n9281), .A2(n9280), .ZN(n14544) );
  INV_X1 U9237 ( .A(n11571), .ZN(n14552) );
  NAND2_X1 U9238 ( .A1(n10466), .A2(n10465), .ZN(n14641) );
  OR2_X1 U9239 ( .A1(n10476), .A2(n10475), .ZN(n10843) );
  INV_X1 U9240 ( .A(n14499), .ZN(n15036) );
  NAND2_X1 U9241 ( .A1(n14791), .A2(n7550), .ZN(n14779) );
  AND2_X1 U9242 ( .A1(n14791), .A2(n7548), .ZN(n14778) );
  NAND2_X1 U9243 ( .A1(n7789), .A2(n7788), .ZN(n14777) );
  AND2_X1 U9244 ( .A1(n7789), .A2(n7786), .ZN(n14775) );
  NAND2_X1 U9245 ( .A1(n7798), .A2(n7801), .ZN(n14897) );
  OR2_X1 U9246 ( .A1(n14926), .A2(n7802), .ZN(n7798) );
  NAND2_X1 U9247 ( .A1(n7805), .A2(n12097), .ZN(n14913) );
  OR2_X1 U9248 ( .A1(n14926), .A2(n14927), .ZN(n7805) );
  INV_X1 U9249 ( .A(n7256), .ZN(n14911) );
  AOI21_X1 U9250 ( .B1(n7260), .B2(n6459), .A(n7259), .ZN(n7256) );
  NAND2_X1 U9251 ( .A1(n7260), .A2(n14380), .ZN(n14928) );
  NAND2_X1 U9252 ( .A1(n7543), .A2(n12127), .ZN(n14951) );
  NAND2_X1 U9253 ( .A1(n12092), .A2(n12091), .ZN(n15003) );
  NAND2_X1 U9254 ( .A1(n11926), .A2(n11845), .ZN(n11846) );
  NAND2_X1 U9255 ( .A1(n7239), .A2(n14507), .ZN(n15303) );
  INV_X1 U9256 ( .A(n15268), .ZN(n14982) );
  OR2_X1 U9257 ( .A1(n14476), .A2(n10188), .ZN(n7454) );
  OAI22_X1 U9258 ( .A1(n12036), .A2(n10189), .B1(n10264), .B2(n9291), .ZN(
        n7554) );
  OR2_X1 U9259 ( .A1(n10814), .A2(n15030), .ZN(n14977) );
  INV_X1 U9260 ( .A(n14994), .ZN(n15260) );
  NAND2_X1 U9261 ( .A1(n6756), .A2(n6559), .ZN(n15161) );
  OR2_X1 U9262 ( .A1(n15043), .A2(n15296), .ZN(n6756) );
  AND2_X1 U9263 ( .A1(n7475), .A2(n7474), .ZN(n7270) );
  INV_X1 U9264 ( .A(n6679), .ZN(n15062) );
  NAND2_X1 U9265 ( .A1(n7214), .A2(n7213), .ZN(n15168) );
  INV_X1 U9266 ( .A(n15076), .ZN(n7214) );
  OR3_X1 U9267 ( .A1(n15127), .A2(n15126), .A3(n15125), .ZN(n15176) );
  AND3_X1 U9268 ( .A1(n8822), .A2(n7954), .A3(n6737), .ZN(n6739) );
  AND2_X1 U9269 ( .A1(n8823), .A2(n8867), .ZN(n7806) );
  NAND2_X1 U9270 ( .A1(n7899), .A2(n7897), .ZN(n13446) );
  INV_X1 U9271 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n15767) );
  INV_X1 U9272 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n11495) );
  OR2_X1 U9273 ( .A1(n9226), .A2(n7509), .ZN(n6579) );
  INV_X1 U9274 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10896) );
  INV_X1 U9275 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10831) );
  INV_X1 U9276 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10764) );
  XNOR2_X1 U9277 ( .A(n9161), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11627) );
  AND2_X1 U9278 ( .A1(n9160), .A2(n9140), .ZN(n11377) );
  INV_X1 U9279 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n15769) );
  INV_X1 U9280 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10464) );
  INV_X1 U9281 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10286) );
  INV_X1 U9282 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10242) );
  INV_X1 U9283 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10238) );
  INV_X1 U9284 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10196) );
  INV_X1 U9285 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n10179) );
  INV_X1 U9286 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n10170) );
  INV_X1 U9287 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10168) );
  XNOR2_X1 U9288 ( .A(n8946), .B(n8945), .ZN(n14589) );
  INV_X1 U9289 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10166) );
  NOR2_X1 U9290 ( .A1(n8746), .A2(n15835), .ZN(n15206) );
  INV_X1 U9291 ( .A(n15210), .ZN(n7626) );
  XNOR2_X1 U9292 ( .A(n8774), .B(n8773), .ZN(n15228) );
  NAND3_X1 U9293 ( .A1(n15240), .A2(n15242), .A3(n7640), .ZN(n15222) );
  INV_X1 U9294 ( .A(n6530), .ZN(n7640) );
  NAND2_X1 U9295 ( .A1(n15240), .A2(n15242), .ZN(n8791) );
  OAI21_X1 U9296 ( .B1(n15201), .B2(n15202), .A(n13647), .ZN(n7300) );
  NAND2_X1 U9297 ( .A1(n15201), .A2(n15202), .ZN(n15200) );
  OAI21_X1 U9298 ( .B1(n12735), .B2(n7377), .A(n15595), .ZN(n7376) );
  INV_X1 U9299 ( .A(n7171), .ZN(n7170) );
  OAI21_X1 U9300 ( .B1(n12767), .B2(n12922), .A(n12766), .ZN(n7171) );
  MUX2_X1 U9301 ( .A(n12775), .B(n12999), .S(n15616), .Z(n12776) );
  NOR2_X1 U9302 ( .A1(n15665), .A2(n10089), .ZN(n10090) );
  NAND2_X1 U9303 ( .A1(n6632), .A2(n10104), .ZN(n7665) );
  AOI21_X1 U9304 ( .B1(n12024), .B2(n13148), .A(n12023), .ZN(n12025) );
  NAND2_X1 U9305 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  AOI21_X1 U9306 ( .B1(n12017), .B2(n12016), .A(n13250), .ZN(n12024) );
  NAND2_X1 U9307 ( .A1(n13229), .A2(n7217), .ZN(n10707) );
  OAI21_X1 U9308 ( .B1(n13123), .B2(n6453), .A(n7491), .ZN(n13210) );
  AND2_X1 U9309 ( .A1(n6935), .A2(n6934), .ZN(n13247) );
  NAND2_X1 U9310 ( .A1(n6933), .A2(n6932), .ZN(P2_U3532) );
  NAND2_X1 U9311 ( .A1(n13611), .A2(n7217), .ZN(n6932) );
  OR2_X1 U9312 ( .A1(n13611), .A2(n10188), .ZN(n6933) );
  NAND2_X1 U9313 ( .A1(n7033), .A2(n13913), .ZN(n7965) );
  INV_X1 U9314 ( .A(n8695), .ZN(n8696) );
  INV_X1 U9315 ( .A(n8699), .ZN(n7033) );
  OR2_X1 U9316 ( .A1(n15538), .A2(n8600), .ZN(n7145) );
  NOR2_X1 U9317 ( .A1(n6624), .A2(n7950), .ZN(n7949) );
  NAND2_X1 U9318 ( .A1(n8811), .A2(n15538), .ZN(n7951) );
  NOR2_X1 U9319 ( .A1(n15538), .A2(n15711), .ZN(n7950) );
  NAND2_X1 U9320 ( .A1(n7192), .A2(n7191), .ZN(n13946) );
  OR2_X1 U9321 ( .A1(n15538), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n7191) );
  NAND2_X1 U9322 ( .A1(n14050), .A2(n15538), .ZN(n7192) );
  AOI21_X1 U9323 ( .B1(P2_REG0_REG_28__SCAN_IN), .B2(n15531), .A(n6626), .ZN(
        n7232) );
  NAND2_X1 U9324 ( .A1(n8811), .A2(n15533), .ZN(n7233) );
  AOI21_X1 U9325 ( .B1(n14487), .B2(n6855), .A(n6857), .ZN(n6856) );
  NAND2_X1 U9326 ( .A1(n6854), .A2(n11451), .ZN(n6858) );
  NAND2_X1 U9327 ( .A1(n6691), .A2(n6690), .ZN(n14741) );
  NAND2_X1 U9328 ( .A1(n6558), .A2(n6692), .ZN(n6691) );
  NAND2_X1 U9329 ( .A1(n14739), .A2(n14526), .ZN(n6690) );
  NAND2_X1 U9330 ( .A1(n7473), .A2(n7472), .ZN(P1_U3557) );
  NAND2_X1 U9331 ( .A1(n15365), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n7472) );
  NAND2_X1 U9332 ( .A1(n15161), .A2(n15367), .ZN(n7473) );
  NAND2_X1 U9333 ( .A1(n6755), .A2(n6754), .ZN(P1_U3525) );
  NAND2_X1 U9334 ( .A1(n15353), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6754) );
  NAND2_X1 U9335 ( .A1(n15161), .A2(n15354), .ZN(n6755) );
  NAND2_X1 U9336 ( .A1(n7212), .A2(n7211), .ZN(P1_U3520) );
  NAND2_X1 U9337 ( .A1(n15353), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U9338 ( .A1(n15168), .A2(n15354), .ZN(n7212) );
  INV_X1 U9339 ( .A(n6662), .ZN(n15827) );
  NAND2_X1 U9340 ( .A1(n15216), .A2(n15215), .ZN(n15214) );
  NAND2_X1 U9341 ( .A1(n15212), .A2(n8765), .ZN(n15216) );
  NAND2_X1 U9342 ( .A1(n15225), .A2(n15224), .ZN(n15223) );
  NAND2_X1 U9343 ( .A1(n7624), .A2(n15218), .ZN(n15225) );
  NOR2_X1 U9344 ( .A1(n15231), .A2(n15230), .ZN(n15229) );
  NAND2_X1 U9345 ( .A1(n7310), .A2(n6454), .ZN(n15233) );
  INV_X1 U9346 ( .A(n15238), .ZN(n15237) );
  OR2_X1 U9347 ( .A1(n11673), .A2(n11674), .ZN(n6449) );
  NAND2_X1 U9348 ( .A1(n7543), .A2(n7261), .ZN(n7260) );
  AND2_X1 U9349 ( .A1(n11995), .A2(n7355), .ZN(n6450) );
  INV_X1 U9350 ( .A(n7606), .ZN(n7605) );
  OAI21_X1 U9351 ( .B1(n12586), .B2(n12587), .A(n7608), .ZN(n7606) );
  AND2_X1 U9352 ( .A1(n12226), .A2(n12822), .ZN(n6451) );
  AND2_X1 U9353 ( .A1(n6484), .A2(n13410), .ZN(n6452) );
  AND2_X1 U9354 ( .A1(n13204), .A2(n11989), .ZN(n6453) );
  AND2_X1 U9355 ( .A1(n15234), .A2(n7311), .ZN(n6454) );
  INV_X1 U9356 ( .A(n14806), .ZN(n7795) );
  NAND2_X1 U9357 ( .A1(n12317), .A2(n12569), .ZN(n6455) );
  AND2_X1 U9358 ( .A1(n7357), .A2(n11996), .ZN(n6456) );
  AND2_X1 U9359 ( .A1(n7759), .A2(n13857), .ZN(n6457) );
  OR2_X1 U9360 ( .A1(n11695), .A2(n11694), .ZN(n6458) );
  NOR2_X1 U9361 ( .A1(n12130), .A2(n14381), .ZN(n6459) );
  OR2_X1 U9362 ( .A1(n13940), .A2(n13720), .ZN(n6460) );
  NAND2_X1 U9363 ( .A1(n11272), .A2(n12577), .ZN(n6461) );
  AND2_X1 U9364 ( .A1(n14349), .A2(n14348), .ZN(n6462) );
  AND2_X1 U9365 ( .A1(n13883), .A2(n6457), .ZN(n6463) );
  AND2_X1 U9366 ( .A1(n14843), .A2(n7471), .ZN(n6464) );
  AND2_X1 U9367 ( .A1(n7467), .A2(n7466), .ZN(n6465) );
  AND2_X1 U9368 ( .A1(n7508), .A2(n8850), .ZN(n6466) );
  NAND2_X1 U9369 ( .A1(n7924), .A2(n8489), .ZN(n13735) );
  OR2_X1 U9370 ( .A1(n13027), .A2(n12837), .ZN(n6467) );
  AND2_X1 U9371 ( .A1(n7600), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6468) );
  INV_X1 U9372 ( .A(n11852), .ZN(n7777) );
  AND3_X1 U9373 ( .A1(n11436), .A2(n12536), .A3(n6789), .ZN(n6469) );
  AND4_X1 U9374 ( .A1(n12532), .A2(n7647), .A3(n12531), .A4(n12530), .ZN(n6470) );
  AND4_X1 U9375 ( .A1(n12519), .A2(n12515), .A3(n12514), .A4(n12513), .ZN(
        n6471) );
  AND3_X1 U9376 ( .A1(n8381), .A2(n8358), .A3(SI_18_), .ZN(n6472) );
  INV_X1 U9377 ( .A(n10874), .ZN(n7208) );
  NOR2_X1 U9378 ( .A1(n7697), .A2(n13817), .ZN(n6473) );
  AND2_X1 U9379 ( .A1(n6573), .A2(n12131), .ZN(n6474) );
  AND2_X1 U9380 ( .A1(n13341), .A2(n13340), .ZN(n6475) );
  OR2_X1 U9381 ( .A1(n7780), .A2(n14869), .ZN(n6476) );
  AND3_X1 U9382 ( .A1(n8117), .A2(n8116), .A3(n8118), .ZN(n6477) );
  AND2_X1 U9383 ( .A1(n14096), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6478) );
  AND2_X1 U9384 ( .A1(n8672), .A2(n7969), .ZN(n6479) );
  INV_X1 U9385 ( .A(n6975), .ZN(n6973) );
  NAND2_X1 U9386 ( .A1(n11234), .A2(n6458), .ZN(n6975) );
  OR2_X1 U9387 ( .A1(n6507), .A2(n7298), .ZN(n6480) );
  OR2_X1 U9388 ( .A1(n15144), .A2(n15149), .ZN(n7462) );
  OR2_X1 U9389 ( .A1(n12474), .A2(n6581), .ZN(n6481) );
  INV_X1 U9390 ( .A(n14352), .ZN(n6874) );
  NOR2_X1 U9391 ( .A1(n15584), .A2(n11235), .ZN(n6482) );
  AND2_X1 U9392 ( .A1(n8756), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n6483) );
  AND2_X1 U9393 ( .A1(n13407), .A2(n13406), .ZN(n6484) );
  AND2_X1 U9394 ( .A1(n10692), .A2(n10691), .ZN(n6485) );
  INV_X1 U9395 ( .A(n7959), .ZN(n7346) );
  INV_X1 U9396 ( .A(n7493), .ZN(n12152) );
  AND2_X1 U9397 ( .A1(n7710), .A2(n9879), .ZN(n6487) );
  NAND2_X1 U9398 ( .A1(n7606), .A2(n12637), .ZN(n6903) );
  INV_X1 U9399 ( .A(n9679), .ZN(n6810) );
  INV_X1 U9400 ( .A(n7714), .ZN(n7713) );
  INV_X1 U9401 ( .A(n12893), .ZN(n6701) );
  AND2_X1 U9402 ( .A1(n7089), .A2(n10048), .ZN(n10202) );
  AND2_X1 U9403 ( .A1(n9807), .A2(n6924), .ZN(n6488) );
  AND2_X1 U9404 ( .A1(n15583), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n6489) );
  INV_X1 U9405 ( .A(n6623), .ZN(n7590) );
  NAND2_X1 U9406 ( .A1(n8076), .A2(n8075), .ZN(n13320) );
  INV_X1 U9407 ( .A(n13320), .ZN(n7013) );
  NOR2_X2 U9408 ( .A1(n12152), .A2(n7492), .ZN(n14040) );
  INV_X1 U9409 ( .A(n14040), .ZN(n15522) );
  OR2_X1 U9410 ( .A1(n14735), .A2(n14526), .ZN(n6490) );
  INV_X1 U9411 ( .A(n9893), .ZN(n7751) );
  OR2_X1 U9412 ( .A1(n15538), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6491) );
  OR2_X1 U9413 ( .A1(n15533), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6492) );
  AND3_X1 U9414 ( .A1(n15691), .A2(n9870), .A3(n6917), .ZN(n6493) );
  INV_X1 U9415 ( .A(n8239), .ZN(n8304) );
  INV_X1 U9416 ( .A(n10736), .ZN(n7151) );
  NAND2_X2 U9417 ( .A1(n8884), .A2(n8883), .ZN(n8892) );
  AND2_X1 U9418 ( .A1(n7876), .A2(n8259), .ZN(n6495) );
  INV_X1 U9419 ( .A(n12864), .ZN(n7181) );
  NAND2_X1 U9420 ( .A1(n9570), .A2(n9569), .ZN(n9568) );
  OR2_X1 U9421 ( .A1(n9226), .A2(P1_IR_REG_18__SCAN_IN), .ZN(n6496) );
  INV_X1 U9422 ( .A(n12539), .ZN(n7062) );
  NAND2_X1 U9423 ( .A1(n6769), .A2(n8225), .ZN(n11810) );
  XNOR2_X1 U9424 ( .A(n10007), .B(P3_IR_REG_21__SCAN_IN), .ZN(n12400) );
  INV_X1 U9425 ( .A(n12400), .ZN(n11461) );
  AND2_X1 U9426 ( .A1(n14836), .A2(n7469), .ZN(n6497) );
  INV_X1 U9427 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n13074) );
  AND2_X1 U9428 ( .A1(n7010), .A2(n13162), .ZN(n6498) );
  AND2_X1 U9429 ( .A1(n14934), .A2(n7467), .ZN(n6499) );
  NOR3_X1 U9430 ( .A1(n14755), .A2(n12113), .A3(n12112), .ZN(n6500) );
  NOR2_X1 U9431 ( .A1(n15525), .A2(n13605), .ZN(n6501) );
  OR2_X1 U9432 ( .A1(n10081), .A2(n10080), .ZN(n6502) );
  AND2_X1 U9433 ( .A1(n7016), .A2(n7356), .ZN(n6503) );
  OR2_X1 U9434 ( .A1(n7306), .A2(n6454), .ZN(n6504) );
  AND2_X1 U9435 ( .A1(n13338), .A2(n13337), .ZN(n6505) );
  NAND2_X1 U9436 ( .A1(n8177), .A2(n8176), .ZN(n13352) );
  AND2_X1 U9437 ( .A1(n7865), .A2(n7863), .ZN(n6506) );
  AND2_X1 U9438 ( .A1(n13412), .A2(n13411), .ZN(n6507) );
  NOR2_X1 U9439 ( .A1(n9583), .A2(n7737), .ZN(n7742) );
  NOR2_X1 U9440 ( .A1(n15154), .A2(n11920), .ZN(n6508) );
  OR2_X1 U9441 ( .A1(n11644), .A2(n12573), .ZN(n6509) );
  INV_X1 U9442 ( .A(n10693), .ZN(n6912) );
  NAND4_X1 U9443 ( .A1(n8063), .A2(n8064), .A3(n8062), .A4(n8061), .ZN(n13609)
         );
  OAI21_X1 U9444 ( .B1(n9529), .B2(P3_IR_REG_0__SCAN_IN), .A(n9513), .ZN(
        n10756) );
  INV_X1 U9445 ( .A(n10756), .ZN(n7809) );
  OR2_X1 U9446 ( .A1(n13816), .A2(n13817), .ZN(n6510) );
  AND2_X1 U9447 ( .A1(n7585), .A2(n9159), .ZN(n6511) );
  AND3_X1 U9448 ( .A1(n9581), .A2(n9579), .A3(n9580), .ZN(n6512) );
  OR2_X1 U9449 ( .A1(n12780), .A2(n12779), .ZN(n6513) );
  OR3_X1 U9450 ( .A1(n11639), .A2(n12574), .A3(n12575), .ZN(n6514) );
  XOR2_X1 U9451 ( .A(n13567), .B(n13672), .Z(n6515) );
  OR2_X1 U9452 ( .A1(n12595), .A2(n12600), .ZN(n6516) );
  AND4_X1 U9453 ( .A1(n15006), .A2(n14368), .A3(n15009), .A4(n6412), .ZN(n6517) );
  NAND2_X1 U9454 ( .A1(n12202), .A2(n8871), .ZN(n9079) );
  OR2_X1 U9455 ( .A1(n13352), .A2(n8187), .ZN(n6518) );
  AND2_X1 U9456 ( .A1(n9624), .A2(n6929), .ZN(n6519) );
  AND2_X1 U9457 ( .A1(n6702), .A2(n6698), .ZN(n6520) );
  INV_X1 U9458 ( .A(n13546), .ZN(n6766) );
  NAND2_X1 U9459 ( .A1(n12048), .A2(n8679), .ZN(n13759) );
  NAND2_X1 U9460 ( .A1(n11812), .A2(n8247), .ZN(n13895) );
  NAND2_X1 U9461 ( .A1(n12815), .A2(n12501), .ZN(n12800) );
  INV_X1 U9462 ( .A(n8678), .ZN(n13765) );
  NAND2_X1 U9463 ( .A1(n13112), .A2(n12001), .ZN(n6521) );
  AND2_X1 U9464 ( .A1(n13360), .A2(n13359), .ZN(n6522) );
  AND2_X1 U9465 ( .A1(n11148), .A2(n11077), .ZN(n6523) );
  NAND2_X1 U9466 ( .A1(n8569), .A2(n8568), .ZN(n13456) );
  INV_X1 U9467 ( .A(n13456), .ZN(n6880) );
  INV_X1 U9468 ( .A(n11996), .ZN(n7355) );
  INV_X1 U9469 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7990) );
  AOI21_X1 U9470 ( .B1(n14805), .B2(n9388), .A(n9391), .ZN(n14750) );
  NAND4_X1 U9471 ( .A1(n9521), .A2(n9520), .A3(n9519), .A4(n9518), .ZN(n9533)
         );
  AND2_X1 U9472 ( .A1(n11499), .A2(n10919), .ZN(n6524) );
  INV_X1 U9473 ( .A(n13349), .ZN(n6728) );
  AND2_X1 U9474 ( .A1(n10048), .A2(n10040), .ZN(n6525) );
  NAND2_X1 U9475 ( .A1(n9242), .A2(n9241), .ZN(n6526) );
  INV_X1 U9476 ( .A(n14860), .ZN(n7780) );
  OR2_X1 U9477 ( .A1(n13820), .A2(n14065), .ZN(n6527) );
  NAND2_X1 U9478 ( .A1(n13044), .A2(n12333), .ZN(n6528) );
  AND2_X1 U9479 ( .A1(n13317), .A2(n13316), .ZN(n6529) );
  XOR2_X1 U9480 ( .A(n8789), .B(n8788), .Z(n6530) );
  AND2_X1 U9481 ( .A1(n13529), .A2(n13528), .ZN(n6531) );
  OR2_X1 U9482 ( .A1(n7622), .A2(n7623), .ZN(n6532) );
  AND2_X1 U9483 ( .A1(n6939), .A2(n6936), .ZN(n6533) );
  AND2_X1 U9484 ( .A1(n7007), .A2(n7005), .ZN(n6534) );
  AND3_X1 U9485 ( .A1(n12885), .A2(n12872), .A3(n6785), .ZN(n6535) );
  INV_X1 U9486 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8011) );
  AND2_X1 U9487 ( .A1(n7387), .A2(n8673), .ZN(n6536) );
  NAND2_X1 U9488 ( .A1(n8547), .A2(n8546), .ZN(n13933) );
  OR2_X1 U9489 ( .A1(n8308), .A2(SI_14_), .ZN(n6537) );
  OR2_X1 U9490 ( .A1(n8760), .A2(n8759), .ZN(n6538) );
  AND3_X1 U9491 ( .A1(n7478), .A2(n7477), .A3(n7476), .ZN(n6539) );
  AND2_X1 U9492 ( .A1(n11423), .A2(n12576), .ZN(n6540) );
  AND2_X1 U9493 ( .A1(n9617), .A2(n10146), .ZN(n6541) );
  NAND2_X1 U9494 ( .A1(n9000), .A2(n8999), .ZN(n14319) );
  AND2_X1 U9495 ( .A1(n8046), .A2(n10314), .ZN(n6542) );
  NAND2_X1 U9496 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), 
        .ZN(n6543) );
  NOR2_X1 U9497 ( .A1(n13328), .A2(n13607), .ZN(n6544) );
  OR2_X1 U9498 ( .A1(n14409), .A2(n7534), .ZN(n6545) );
  INV_X1 U9499 ( .A(n8404), .ZN(n7031) );
  AND2_X1 U9500 ( .A1(n9558), .A2(n9559), .ZN(n10971) );
  INV_X1 U9501 ( .A(n10971), .ZN(n7155) );
  NAND4_X1 U9502 ( .A1(n7140), .A2(n10005), .A3(n10031), .A4(n9479), .ZN(
        n10025) );
  AND2_X1 U9503 ( .A1(n13364), .A2(n13363), .ZN(n6546) );
  INV_X1 U9504 ( .A(n15202), .ZN(n6827) );
  INV_X1 U9505 ( .A(n7833), .ZN(n7832) );
  NAND2_X1 U9506 ( .A1(n12779), .A2(n7834), .ZN(n7833) );
  NAND2_X1 U9507 ( .A1(n8791), .A2(n6530), .ZN(n8790) );
  NAND3_X1 U9508 ( .A1(n14290), .A2(n14303), .A3(n14289), .ZN(n6547) );
  INV_X1 U9509 ( .A(n7822), .ZN(n7821) );
  OAI21_X1 U9510 ( .B1(n10078), .B2(n7823), .A(n12463), .ZN(n7822) );
  OR2_X1 U9511 ( .A1(n15215), .A2(n7632), .ZN(n6548) );
  AND2_X1 U9512 ( .A1(n7350), .A2(n7347), .ZN(n6549) );
  NAND2_X1 U9513 ( .A1(n13487), .A2(n13486), .ZN(n6550) );
  NAND2_X1 U9514 ( .A1(n13940), .A2(n13720), .ZN(n6551) );
  NAND2_X1 U9515 ( .A1(n13490), .A2(n13489), .ZN(n6552) );
  NOR2_X1 U9516 ( .A1(n14554), .A2(n11345), .ZN(n6553) );
  INV_X1 U9517 ( .A(n13675), .ZN(n14047) );
  NAND2_X1 U9518 ( .A1(n13498), .A2(n13497), .ZN(n13675) );
  OR2_X1 U9519 ( .A1(n6874), .A2(n14351), .ZN(n6554) );
  INV_X1 U9520 ( .A(n12508), .ZN(n6709) );
  AND2_X1 U9521 ( .A1(n12835), .A2(n12495), .ZN(n6555) );
  OR2_X1 U9522 ( .A1(n7248), .A2(n7250), .ZN(n6556) );
  AND2_X1 U9523 ( .A1(n12462), .A2(n12463), .ZN(n12537) );
  INV_X1 U9524 ( .A(n12537), .ZN(n7323) );
  OR2_X1 U9525 ( .A1(n7914), .A2(n6562), .ZN(n6557) );
  NAND2_X1 U9526 ( .A1(n12515), .A2(n9981), .ZN(n12769) );
  INV_X1 U9527 ( .A(n12769), .ZN(n6818) );
  OR2_X1 U9528 ( .A1(n14734), .A2(n14733), .ZN(n6558) );
  AND2_X1 U9529 ( .A1(n7271), .A2(n7270), .ZN(n6559) );
  AND2_X1 U9530 ( .A1(n13027), .A2(n12569), .ZN(n6560) );
  AND2_X1 U9531 ( .A1(n6467), .A2(n12490), .ZN(n6561) );
  AND2_X1 U9532 ( .A1(n6507), .A2(n7298), .ZN(n6562) );
  AND2_X1 U9533 ( .A1(n14327), .A2(n11521), .ZN(n6563) );
  AND2_X1 U9534 ( .A1(n9384), .A2(n9383), .ZN(n6564) );
  NAND2_X1 U9535 ( .A1(n14848), .A2(n12101), .ZN(n14869) );
  INV_X1 U9536 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n9479) );
  INV_X1 U9537 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7206) );
  INV_X1 U9538 ( .A(n13153), .ZN(n7357) );
  INV_X1 U9539 ( .A(n8680), .ZN(n7392) );
  AND2_X1 U9540 ( .A1(n12309), .A2(n7854), .ZN(n6565) );
  INV_X1 U9541 ( .A(n14413), .ZN(n7517) );
  AND2_X1 U9542 ( .A1(n10140), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6566) );
  AND2_X1 U9543 ( .A1(n13062), .A2(n12293), .ZN(n12470) );
  NOR2_X1 U9544 ( .A1(n6577), .A2(n13393), .ZN(n6567) );
  NOR2_X1 U9545 ( .A1(n13032), .A2(n12570), .ZN(n6568) );
  NOR2_X1 U9546 ( .A1(n12286), .A2(n12293), .ZN(n6569) );
  AND2_X1 U9547 ( .A1(n12803), .A2(n12822), .ZN(n12505) );
  OR2_X1 U9548 ( .A1(n6401), .A2(n13626), .ZN(n6570) );
  INV_X1 U9549 ( .A(n14412), .ZN(n7521) );
  NAND2_X1 U9550 ( .A1(n12375), .A2(n12755), .ZN(n6571) );
  NAND2_X1 U9551 ( .A1(n8339), .A2(n10928), .ZN(n8381) );
  AND2_X1 U9552 ( .A1(n13948), .A2(n13719), .ZN(n6572) );
  INV_X1 U9553 ( .A(n15060), .ZN(n7470) );
  NOR2_X1 U9554 ( .A1(n14907), .A2(n7974), .ZN(n6573) );
  INV_X1 U9555 ( .A(n8892), .ZN(n6853) );
  AND2_X1 U9556 ( .A1(n15009), .A2(n6436), .ZN(n6574) );
  NOR2_X1 U9557 ( .A1(n12013), .A2(n12014), .ZN(n6575) );
  NOR2_X1 U9558 ( .A1(n9951), .A2(n12269), .ZN(n6576) );
  INV_X1 U9559 ( .A(n6699), .ZN(n6698) );
  NAND2_X1 U9560 ( .A1(n6701), .A2(n12394), .ZN(n6699) );
  INV_X1 U9561 ( .A(n7409), .ZN(n9530) );
  AND2_X1 U9562 ( .A1(n13390), .A2(n13389), .ZN(n6577) );
  AND2_X1 U9563 ( .A1(n10369), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6578) );
  AND2_X1 U9564 ( .A1(n7310), .A2(n7311), .ZN(n6580) );
  NAND2_X1 U9565 ( .A1(n9590), .A2(n7131), .ZN(n15627) );
  INV_X1 U9566 ( .A(n15627), .ZN(n7130) );
  OR2_X1 U9567 ( .A1(n7324), .A2(n7323), .ZN(n6581) );
  INV_X1 U9568 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8823) );
  XNOR2_X1 U9569 ( .A(n13676), .B(n13530), .ZN(n13566) );
  INV_X1 U9570 ( .A(n13566), .ZN(n7161) );
  INV_X1 U9571 ( .A(n7940), .ZN(n7939) );
  OR2_X1 U9572 ( .A1(n13809), .A2(n7941), .ZN(n7940) );
  AND2_X1 U9573 ( .A1(n11992), .A2(n11991), .ZN(n6582) );
  INV_X1 U9574 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n10005) );
  OR2_X1 U9575 ( .A1(n14912), .A2(n7804), .ZN(n6583) );
  INV_X1 U9576 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10161) );
  INV_X1 U9577 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10157) );
  AND2_X1 U9578 ( .A1(n13056), .A2(n12916), .ZN(n6584) );
  AND2_X1 U9579 ( .A1(n8671), .A2(n8670), .ZN(n13833) );
  AND2_X1 U9580 ( .A1(n9254), .A2(n9253), .ZN(n6585) );
  INV_X1 U9581 ( .A(n7787), .ZN(n7786) );
  NAND2_X1 U9582 ( .A1(n7788), .A2(n14780), .ZN(n7787) );
  AND2_X1 U9583 ( .A1(n10464), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6586) );
  AND2_X1 U9584 ( .A1(n10458), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n6587) );
  AND2_X1 U9585 ( .A1(n12129), .A2(n12128), .ZN(n14927) );
  INV_X1 U9586 ( .A(n14927), .ZN(n7803) );
  INV_X1 U9587 ( .A(n14409), .ZN(n6866) );
  AND2_X1 U9588 ( .A1(n7993), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6588) );
  INV_X1 U9589 ( .A(n13375), .ZN(n6748) );
  INV_X1 U9590 ( .A(n11234), .ZN(n6978) );
  AND2_X1 U9591 ( .A1(n12109), .A2(n7778), .ZN(n6589) );
  INV_X1 U9592 ( .A(n6461), .ZN(n7848) );
  AND2_X1 U9593 ( .A1(n13327), .A2(n13326), .ZN(n6590) );
  NOR2_X1 U9594 ( .A1(n11699), .A2(n11698), .ZN(n6591) );
  INV_X1 U9595 ( .A(n12509), .ZN(n7835) );
  NAND2_X1 U9596 ( .A1(n12389), .A2(n7422), .ZN(n6592) );
  AND2_X1 U9597 ( .A1(n14554), .A2(n11345), .ZN(n6593) );
  AND2_X1 U9598 ( .A1(n12646), .A2(n12645), .ZN(n6594) );
  OR2_X1 U9599 ( .A1(n15136), .A2(n12093), .ZN(n14371) );
  INV_X1 U9600 ( .A(n7971), .ZN(n7252) );
  INV_X1 U9601 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7464) );
  OR2_X1 U9602 ( .A1(n7911), .A2(n7296), .ZN(n6595) );
  INV_X1 U9603 ( .A(n6918), .ZN(n9929) );
  AND2_X1 U9604 ( .A1(n7225), .A2(n6493), .ZN(n6918) );
  INV_X1 U9605 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n15751) );
  INV_X1 U9606 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U9607 ( .A1(n12224), .A2(n6455), .ZN(n6596) );
  OR2_X1 U9608 ( .A1(n7535), .A2(n6866), .ZN(n6597) );
  NAND2_X1 U9609 ( .A1(n6945), .A2(n7390), .ZN(n13702) );
  NAND2_X1 U9610 ( .A1(n6877), .A2(n6457), .ZN(n13820) );
  INV_X1 U9611 ( .A(n13820), .ZN(n6875) );
  OR2_X1 U9612 ( .A1(n13972), .A2(n13595), .ZN(n6598) );
  AND3_X1 U9613 ( .A1(n12729), .A2(n7379), .A3(n7378), .ZN(n6599) );
  AND2_X1 U9614 ( .A1(n13368), .A2(n13375), .ZN(n6600) );
  INV_X1 U9615 ( .A(n12545), .ZN(n9999) );
  NAND2_X1 U9616 ( .A1(n12519), .A2(n9998), .ZN(n12545) );
  OR2_X1 U9617 ( .A1(n13410), .A2(n6484), .ZN(n6601) );
  AND2_X1 U9618 ( .A1(n12547), .A2(n12373), .ZN(n6602) );
  INV_X1 U9619 ( .A(n14877), .ZN(n15084) );
  NAND2_X1 U9620 ( .A1(n15197), .A2(n6434), .ZN(n14877) );
  NOR2_X1 U9621 ( .A1(n8684), .A2(n13836), .ZN(n6603) );
  AND2_X1 U9622 ( .A1(n6881), .A2(n6880), .ZN(n6604) );
  NOR2_X1 U9623 ( .A1(n12003), .A2(n7480), .ZN(n6605) );
  INV_X1 U9624 ( .A(n6961), .ZN(n6960) );
  INV_X1 U9625 ( .A(n8247), .ZN(n7927) );
  AND2_X1 U9626 ( .A1(n9013), .A2(n11080), .ZN(n6606) );
  AND2_X1 U9627 ( .A1(n7906), .A2(n13334), .ZN(n6607) );
  OR2_X1 U9628 ( .A1(n13050), .A2(n12328), .ZN(n12390) );
  NAND2_X1 U9629 ( .A1(n14813), .A2(n14812), .ZN(n6608) );
  AND2_X1 U9630 ( .A1(n12508), .A2(n9937), .ZN(n12807) );
  INV_X1 U9631 ( .A(n12807), .ZN(n12801) );
  NAND2_X1 U9632 ( .A1(n14456), .A2(n14455), .ZN(n6609) );
  INV_X1 U9633 ( .A(n12843), .ZN(n12835) );
  NAND2_X1 U9634 ( .A1(n12497), .A2(n9911), .ZN(n12843) );
  AND2_X1 U9635 ( .A1(n12095), .A2(n14386), .ZN(n6610) );
  AND2_X1 U9636 ( .A1(n6732), .A2(n6728), .ZN(n6611) );
  AND2_X1 U9637 ( .A1(n12454), .A2(n12455), .ZN(n11436) );
  INV_X1 U9638 ( .A(n12469), .ZN(n7324) );
  INV_X1 U9639 ( .A(n7178), .ZN(n7177) );
  AND2_X1 U9640 ( .A1(n7629), .A2(n7626), .ZN(n6612) );
  NOR2_X1 U9641 ( .A1(n8311), .A2(n8310), .ZN(n6613) );
  NAND2_X1 U9642 ( .A1(n9386), .A2(n9385), .ZN(n14806) );
  AND2_X1 U9643 ( .A1(n6867), .A2(n6545), .ZN(n6614) );
  NAND2_X1 U9644 ( .A1(n14009), .A2(n13599), .ZN(n6615) );
  NAND2_X1 U9645 ( .A1(n11981), .A2(n11980), .ZN(n6616) );
  OR2_X1 U9646 ( .A1(n7919), .A2(n6562), .ZN(n6617) );
  INV_X1 U9647 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7510) );
  AND2_X1 U9648 ( .A1(n7516), .A2(n7515), .ZN(n6618) );
  AND2_X1 U9649 ( .A1(n7925), .A2(n6768), .ZN(n6619) );
  AND2_X1 U9650 ( .A1(n14371), .A2(n7241), .ZN(n6620) );
  AND2_X1 U9651 ( .A1(n13557), .A2(n6677), .ZN(n6621) );
  INV_X1 U9652 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8867) );
  AND2_X1 U9653 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n6622) );
  INV_X1 U9654 ( .A(n8822), .ZN(n7587) );
  INV_X1 U9655 ( .A(n7855), .ZN(n7854) );
  NAND2_X1 U9656 ( .A1(n7856), .A2(n12216), .ZN(n7855) );
  INV_X1 U9657 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n7989) );
  INV_X1 U9658 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U9659 ( .A1(n8686), .A2(n13568), .ZN(n7493) );
  NAND2_X1 U9660 ( .A1(n8589), .A2(n8623), .ZN(n13578) );
  AND2_X1 U9661 ( .A1(n10044), .A2(n10043), .ZN(n10578) );
  INV_X1 U9662 ( .A(n12526), .ZN(n7413) );
  INV_X1 U9663 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n7410) );
  AND2_X1 U9664 ( .A1(n10567), .A2(n10564), .ZN(n13270) );
  NAND2_X1 U9665 ( .A1(n7428), .A2(n7429), .ZN(n11435) );
  INV_X1 U9666 ( .A(n14065), .ZN(n6879) );
  XNOR2_X1 U9667 ( .A(n14555), .B(n14309), .ZN(n14501) );
  INV_X2 U9668 ( .A(n12512), .ZN(n12513) );
  INV_X1 U9669 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7174) );
  INV_X1 U9670 ( .A(n12587), .ZN(n7607) );
  INV_X1 U9671 ( .A(n12784), .ZN(n7227) );
  AND2_X1 U9672 ( .A1(n12657), .A2(n12628), .ZN(n6623) );
  NAND2_X1 U9673 ( .A1(n11091), .A2(n9633), .ZN(n11256) );
  OAI21_X1 U9674 ( .B1(n11188), .B2(n6766), .A(n6763), .ZN(n11166) );
  NAND2_X1 U9675 ( .A1(n7021), .A2(n7018), .ZN(n11730) );
  NAND2_X1 U9676 ( .A1(n8664), .A2(n8663), .ZN(n11728) );
  NAND2_X1 U9677 ( .A1(n11134), .A2(n11133), .ZN(n11344) );
  NAND2_X1 U9678 ( .A1(n7671), .A2(n8656), .ZN(n11170) );
  NAND2_X1 U9679 ( .A1(n11005), .A2(n8654), .ZN(n11181) );
  NAND2_X1 U9680 ( .A1(n6938), .A2(n7381), .ZN(n11318) );
  INV_X1 U9681 ( .A(n15065), .ZN(n7471) );
  OAI211_X1 U9682 ( .C1(n11480), .C2(n6724), .A(n11484), .B(n6721), .ZN(n11485) );
  AND2_X1 U9683 ( .A1(n7498), .A2(n11976), .ZN(n7497) );
  AND2_X1 U9684 ( .A1(n13456), .A2(n14023), .ZN(n6624) );
  OR2_X1 U9685 ( .A1(n11796), .A2(n15154), .ZN(n7953) );
  INV_X1 U9686 ( .A(n7953), .ZN(n7459) );
  AND3_X1 U9687 ( .A1(n7602), .A2(n7599), .A3(n6903), .ZN(n6625) );
  OR2_X1 U9688 ( .A1(n14877), .A2(n14543), .ZN(n14848) );
  INV_X1 U9689 ( .A(n14848), .ZN(n7779) );
  AND2_X1 U9690 ( .A1(n13456), .A2(n14086), .ZN(n6626) );
  AND2_X1 U9691 ( .A1(n7561), .A2(n7559), .ZN(n11567) );
  AND2_X1 U9692 ( .A1(n9849), .A2(n9848), .ZN(n12333) );
  INV_X1 U9693 ( .A(n12333), .ZN(n12895) );
  AND2_X1 U9694 ( .A1(n6702), .A2(n12394), .ZN(n6627) );
  NOR2_X1 U9695 ( .A1(n12587), .A2(n12646), .ZN(n6628) );
  INV_X1 U9696 ( .A(n6806), .ZN(n6805) );
  NOR2_X1 U9697 ( .A1(n9695), .A2(n6807), .ZN(n6806) );
  INV_X1 U9698 ( .A(n7734), .ZN(n7733) );
  NOR2_X1 U9699 ( .A1(n9783), .A2(n7735), .ZN(n7734) );
  INV_X1 U9700 ( .A(n12822), .ZN(n12796) );
  AND2_X1 U9701 ( .A1(n9936), .A2(n9935), .ZN(n12822) );
  INV_X1 U9702 ( .A(n12328), .ZN(n12903) );
  AND2_X1 U9703 ( .A1(n9830), .A2(n9829), .ZN(n12328) );
  NAND2_X1 U9704 ( .A1(n13883), .A2(n7759), .ZN(n7760) );
  AND2_X1 U9705 ( .A1(n12615), .A2(n6982), .ZN(n6629) );
  OR2_X1 U9706 ( .A1(n9885), .A2(n6919), .ZN(n6630) );
  AND2_X1 U9707 ( .A1(n11851), .A2(n11921), .ZN(n6631) );
  NAND2_X2 U9708 ( .A1(n9272), .A2(n9271), .ZN(n14891) );
  INV_X1 U9709 ( .A(n14891), .ZN(n7466) );
  INV_X1 U9710 ( .A(n12524), .ZN(n7647) );
  OR2_X1 U9711 ( .A1(n12763), .A2(n15653), .ZN(n6632) );
  INV_X1 U9712 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n12078) );
  AND2_X1 U9713 ( .A1(n10900), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n6633) );
  AND2_X1 U9714 ( .A1(n8561), .A2(SI_27_), .ZN(n6634) );
  AND2_X1 U9715 ( .A1(n10896), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6635) );
  NOR2_X1 U9716 ( .A1(n12218), .A2(n12570), .ZN(n6636) );
  AND2_X1 U9717 ( .A1(n7207), .A2(n12895), .ZN(n6637) );
  OR2_X1 U9718 ( .A1(n14053), .A2(n14079), .ZN(n6638) );
  AND2_X1 U9719 ( .A1(n7273), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n6639) );
  INV_X1 U9720 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7597) );
  AND2_X1 U9721 ( .A1(n6926), .A2(n6925), .ZN(n6640) );
  AND2_X1 U9722 ( .A1(n7604), .A2(n7607), .ZN(n6641) );
  AND2_X1 U9723 ( .A1(n7302), .A2(n7301), .ZN(n15219) );
  INV_X1 U9724 ( .A(n15219), .ZN(n7624) );
  AND2_X1 U9725 ( .A1(n7589), .A2(n6623), .ZN(n6642) );
  INV_X1 U9726 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n10031) );
  NOR2_X1 U9727 ( .A1(n12521), .A2(n12560), .ZN(n6643) );
  AND2_X1 U9728 ( .A1(n10447), .A2(n15543), .ZN(n6644) );
  NAND2_X1 U9729 ( .A1(n8058), .A2(n7396), .ZN(n13286) );
  INV_X1 U9730 ( .A(n13286), .ZN(n6888) );
  INV_X1 U9731 ( .A(n15468), .ZN(n7441) );
  INV_X2 U9732 ( .A(n15353), .ZN(n15354) );
  INV_X2 U9733 ( .A(n15365), .ZN(n15367) );
  INV_X1 U9734 ( .A(n9899), .ZN(n7752) );
  AND2_X1 U9735 ( .A1(P3_U3897), .A2(n13081), .ZN(n15595) );
  NAND2_X1 U9736 ( .A1(n13630), .A2(n13631), .ZN(n13629) );
  OAI211_X1 U9737 ( .C1(SI_2_), .C2(n9989), .A(n9532), .B(n9531), .ZN(n12990)
         );
  INV_X1 U9738 ( .A(n12990), .ZN(n7169) );
  AND2_X1 U9739 ( .A1(n13499), .A2(n8590), .ZN(n13836) );
  INV_X1 U9740 ( .A(n13836), .ZN(n13897) );
  NAND2_X1 U9741 ( .A1(n6738), .A2(n7586), .ZN(n6645) );
  NAND2_X1 U9742 ( .A1(n7456), .A2(n11051), .ZN(n7457) );
  INV_X1 U9743 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n7276) );
  INV_X1 U9744 ( .A(n9912), .ZN(n7755) );
  NAND2_X1 U9745 ( .A1(n15408), .A2(n15409), .ZN(n6646) );
  AND2_X1 U9746 ( .A1(n7448), .A2(n7449), .ZN(n6647) );
  AND2_X1 U9747 ( .A1(n11807), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6648) );
  INV_X1 U9748 ( .A(n6885), .ZN(n11192) );
  OR2_X1 U9749 ( .A1(n6886), .A2(n11207), .ZN(n6885) );
  AND2_X1 U9750 ( .A1(n11495), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6649) );
  AND2_X1 U9751 ( .A1(n10694), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n6650) );
  AND2_X1 U9752 ( .A1(n7278), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6651) );
  INV_X1 U9753 ( .A(n12746), .ZN(n6986) );
  INV_X1 U9754 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n6920) );
  INV_X1 U9755 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n8821) );
  AND2_X1 U9756 ( .A1(n7593), .A2(n10405), .ZN(n7596) );
  AND2_X1 U9757 ( .A1(n12746), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n6652) );
  INV_X1 U9758 ( .A(n10688), .ZN(n7372) );
  AND2_X1 U9759 ( .A1(n10098), .A2(n10011), .ZN(n12834) );
  INV_X1 U9760 ( .A(n12834), .ZN(n12986) );
  XNOR2_X1 U9761 ( .A(n7035), .B(n7990), .ZN(n7993) );
  INV_X1 U9762 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6948) );
  INV_X1 U9763 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7553) );
  INV_X1 U9764 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7313) );
  INV_X1 U9765 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n6684) );
  INV_X1 U9766 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7632) );
  INV_X1 U9767 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n7619) );
  INV_X1 U9768 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n6909) );
  NAND2_X1 U9769 ( .A1(n7878), .A2(n8205), .ZN(n7876) );
  NAND2_X1 U9770 ( .A1(n6654), .A2(n6620), .ZN(n14988) );
  NAND2_X1 U9771 ( .A1(n14896), .A2(n12098), .ZN(n14880) );
  NAND2_X1 U9772 ( .A1(n8041), .A2(n8042), .ZN(n8045) );
  NAND2_X1 U9773 ( .A1(n8029), .A2(n8913), .ZN(n8042) );
  NAND2_X1 U9774 ( .A1(n7238), .A2(n7799), .ZN(n14896) );
  OR2_X1 U9775 ( .A1(n15149), .A2(n11853), .ZN(n11851) );
  XNOR2_X2 U9776 ( .A(n7299), .B(n8763), .ZN(n15213) );
  NAND2_X2 U9777 ( .A1(n6662), .A2(n6570), .ZN(n7299) );
  NAND3_X1 U9778 ( .A1(n7628), .A2(n7627), .A3(n6612), .ZN(n7631) );
  XNOR2_X2 U9779 ( .A(n8755), .B(n8754), .ZN(n15825) );
  NAND2_X1 U9780 ( .A1(n6739), .A2(n6738), .ZN(n15182) );
  AND2_X2 U9781 ( .A1(n14530), .A2(n14531), .ZN(n14532) );
  NAND2_X1 U9782 ( .A1(n7056), .A2(n7058), .ZN(n7952) );
  OAI21_X1 U9783 ( .B1(n12764), .B2(n12763), .A(n15665), .ZN(n7153) );
  XNOR2_X1 U9784 ( .A(n7072), .B(n12545), .ZN(n7071) );
  NAND2_X1 U9785 ( .A1(n7071), .A2(n12986), .ZN(n7070) );
  NOR2_X1 U9786 ( .A1(n12773), .A2(n6818), .ZN(n12772) );
  XNOR2_X1 U9787 ( .A(n10415), .B(n10414), .ZN(n10665) );
  NAND2_X1 U9788 ( .A1(n8761), .A2(n8762), .ZN(n8718) );
  NAND2_X1 U9789 ( .A1(n8770), .A2(n8771), .ZN(n8722) );
  AOI21_X2 U9790 ( .B1(n8757), .B2(n8713), .A(n6660), .ZN(n8715) );
  NAND2_X1 U9791 ( .A1(n8766), .A2(n8767), .ZN(n8721) );
  NAND2_X1 U9792 ( .A1(n6670), .A2(n14860), .ZN(n14849) );
  INV_X1 U9793 ( .A(n11851), .ZN(n7776) );
  NOR2_X2 U9794 ( .A1(n8723), .A2(n6661), .ZN(n8776) );
  NAND2_X1 U9795 ( .A1(n6931), .A2(n7385), .ZN(n8678) );
  NAND2_X1 U9796 ( .A1(n6959), .A2(n8669), .ZN(n13829) );
  NAND2_X1 U9797 ( .A1(n6828), .A2(n8759), .ZN(n7628) );
  OR2_X2 U9798 ( .A1(n15828), .A2(n15829), .ZN(n6662) );
  OAI21_X2 U9799 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(n8747), .A(n15205), .ZN(
        n15831) );
  XNOR2_X1 U9800 ( .A(n8744), .B(n8745), .ZN(n15836) );
  NOR2_X1 U9801 ( .A1(n15836), .A2(n15837), .ZN(n15835) );
  NAND3_X1 U9802 ( .A1(n6663), .A2(n9475), .A3(n9474), .ZN(P1_U3220) );
  NAND2_X1 U9803 ( .A1(n9450), .A2(n7957), .ZN(n6663) );
  NAND2_X1 U9804 ( .A1(n14988), .A2(n14987), .ZN(n7782) );
  NAND2_X1 U9805 ( .A1(n7578), .A2(n7576), .ZN(n14204) );
  OAI22_X1 U9806 ( .A1(n14104), .A2(n7558), .B1(n7559), .B2(n9055), .ZN(n11875) );
  NAND2_X1 U9807 ( .A1(n10757), .A2(n10758), .ZN(n14141) );
  NAND2_X1 U9808 ( .A1(n7173), .A2(n6608), .ZN(n15064) );
  NAND2_X1 U9809 ( .A1(n15064), .A2(n15311), .ZN(n15071) );
  NAND2_X1 U9810 ( .A1(n14868), .A2(n12133), .ZN(n12135) );
  NAND2_X1 U9811 ( .A1(n14972), .A2(n12126), .ZN(n7543) );
  NOR2_X1 U9812 ( .A1(n14816), .A2(n14815), .ZN(n14818) );
  OAI21_X1 U9813 ( .B1(n15058), .B2(n15340), .A(n15061), .ZN(n6679) );
  INV_X1 U9814 ( .A(n11057), .ZN(n7239) );
  NAND2_X1 U9815 ( .A1(n15437), .A2(n15438), .ZN(n15436) );
  OAI21_X1 U9816 ( .B1(n13670), .B2(n15492), .A(n7440), .ZN(n7439) );
  AOI21_X1 U9817 ( .B1(n7439), .B2(n13672), .A(n7438), .ZN(n7437) );
  NOR2_X1 U9818 ( .A1(n11748), .A2(n11747), .ZN(n13648) );
  NOR2_X1 U9819 ( .A1(n10956), .A2(n10955), .ZN(n11746) );
  NAND3_X1 U9820 ( .A1(n6666), .A2(n9654), .A3(n7644), .ZN(n11266) );
  NAND2_X1 U9821 ( .A1(n11092), .A2(n7645), .ZN(n6666) );
  AND2_X2 U9822 ( .A1(n6486), .A2(n6667), .ZN(n12935) );
  NAND2_X1 U9823 ( .A1(n7433), .A2(n13653), .ZN(n7432) );
  NAND2_X2 U9824 ( .A1(n9850), .A2(n12541), .ZN(n12877) );
  NOR2_X1 U9825 ( .A1(n15423), .A2(n7445), .ZN(n10956) );
  NOR2_X1 U9826 ( .A1(n15451), .A2(n7443), .ZN(n11748) );
  NOR2_X1 U9827 ( .A1(n11746), .A2(n7444), .ZN(n15437) );
  NAND2_X2 U9828 ( .A1(n12404), .A2(n12407), .ZN(n12979) );
  NOR2_X1 U9829 ( .A1(n13648), .A2(n7442), .ZN(n13650) );
  XNOR2_X1 U9830 ( .A(n13650), .B(n13652), .ZN(n15462) );
  OAI21_X1 U9831 ( .B1(n13673), .B2(n13672), .A(n7437), .ZN(P2_U3233) );
  INV_X1 U9832 ( .A(n7314), .ZN(n7182) );
  NAND3_X1 U9833 ( .A1(n6914), .A2(n7707), .A3(n6916), .ZN(n6913) );
  NAND2_X1 U9834 ( .A1(n7327), .A2(n12496), .ZN(n7326) );
  NAND2_X1 U9835 ( .A1(n12489), .A2(n7179), .ZN(n12493) );
  OAI21_X1 U9836 ( .B1(n7334), .B2(n7333), .A(n12440), .ZN(n12441) );
  NAND2_X1 U9837 ( .A1(n12503), .A2(n12502), .ZN(n12511) );
  AOI21_X1 U9838 ( .B1(n12406), .B2(n7328), .A(n12405), .ZN(n12412) );
  NAND2_X1 U9839 ( .A1(n8402), .A2(n8404), .ZN(n13801) );
  OAI21_X1 U9840 ( .B1(n8209), .B2(n10289), .A(n6674), .ZN(n8208) );
  NAND3_X1 U9841 ( .A1(n6621), .A2(n6676), .A3(n6675), .ZN(n13560) );
  NAND3_X2 U9842 ( .A1(n7960), .A2(n8818), .A3(n8827), .ZN(n9226) );
  INV_X4 U9843 ( .A(n12036), .ZN(n8962) );
  NAND3_X1 U9844 ( .A1(n6680), .A2(n11468), .A3(n11469), .ZN(n7240) );
  XNOR2_X2 U9845 ( .A(n8715), .B(P3_ADDR_REG_7__SCAN_IN), .ZN(n8737) );
  NAND2_X1 U9846 ( .A1(n7160), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n8570) );
  OAI211_X1 U9847 ( .C1(n13583), .C2(n7902), .A(n6515), .B(n7148), .ZN(n13587)
         );
  INV_X1 U9848 ( .A(n8566), .ZN(n7128) );
  NAND3_X1 U9849 ( .A1(n7414), .A2(n12424), .A3(n6693), .ZN(n7411) );
  NAND3_X1 U9850 ( .A1(n10782), .A2(n10783), .A3(n7416), .ZN(n6693) );
  OR2_X1 U9851 ( .A1(n12817), .A2(n6707), .ZN(n6703) );
  NAND2_X1 U9852 ( .A1(n12817), .A2(n7424), .ZN(n6704) );
  NAND2_X1 U9853 ( .A1(n6703), .A2(n6705), .ZN(n7830) );
  NAND2_X1 U9854 ( .A1(n11435), .A2(n7426), .ZN(n6710) );
  AND2_X2 U9855 ( .A1(n6714), .A2(n8871), .ZN(n8925) );
  NAND3_X1 U9856 ( .A1(n13310), .A2(n13309), .A3(n13311), .ZN(n6716) );
  NAND3_X1 U9857 ( .A1(n6716), .A2(n6720), .A3(n6715), .ZN(n6719) );
  NAND3_X1 U9858 ( .A1(n7905), .A2(n13325), .A3(n6717), .ZN(n7904) );
  NAND2_X1 U9859 ( .A1(n6719), .A2(n6718), .ZN(n6717) );
  NAND3_X1 U9860 ( .A1(n11482), .A2(n6563), .A3(n6725), .ZN(n6724) );
  NAND2_X1 U9861 ( .A1(n6729), .A2(n6611), .ZN(n6730) );
  NOR2_X1 U9862 ( .A1(n7903), .A2(n6505), .ZN(n6733) );
  NAND2_X1 U9863 ( .A1(n11849), .A2(n11848), .ZN(n6736) );
  AND2_X1 U9864 ( .A1(n7510), .A2(n7806), .ZN(n6737) );
  INV_X2 U9865 ( .A(n9226), .ZN(n7588) );
  NAND3_X1 U9866 ( .A1(n6742), .A2(n6741), .A3(n6748), .ZN(n6743) );
  NAND2_X1 U9867 ( .A1(n13369), .A2(n13368), .ZN(n6741) );
  NAND2_X1 U9868 ( .A1(n7900), .A2(n6546), .ZN(n6742) );
  NAND2_X1 U9869 ( .A1(n13369), .A2(n6600), .ZN(n6745) );
  NAND2_X1 U9870 ( .A1(n6744), .A2(n6743), .ZN(n13380) );
  NAND3_X1 U9871 ( .A1(n6746), .A2(n6745), .A3(n6750), .ZN(n6744) );
  NAND3_X1 U9872 ( .A1(n13405), .A2(n13404), .A3(n6601), .ZN(n6759) );
  NAND2_X1 U9873 ( .A1(n11571), .A2(n14325), .ZN(n11521) );
  OAI211_X1 U9874 ( .C1(n6438), .C2(n14109), .A(n9026), .B(n9027), .ZN(n6761)
         );
  INV_X1 U9875 ( .A(n6761), .ZN(n6760) );
  NAND2_X1 U9876 ( .A1(n6765), .A2(n13546), .ZN(n6764) );
  AND2_X1 U9877 ( .A1(n6764), .A2(n8119), .ZN(n6763) );
  NAND2_X1 U9878 ( .A1(n11327), .A2(n13546), .ZN(n11326) );
  NAND2_X1 U9879 ( .A1(n11166), .A2(n8138), .ZN(n8140) );
  NAND2_X1 U9880 ( .A1(n11730), .A2(n6770), .ZN(n6767) );
  NAND2_X1 U9881 ( .A1(n6767), .A2(n6619), .ZN(n8274) );
  NAND2_X1 U9882 ( .A1(n8557), .A2(n6774), .ZN(n8807) );
  NAND2_X1 U9883 ( .A1(n8557), .A2(n8556), .ZN(n7921) );
  NAND2_X1 U9884 ( .A1(n7924), .A2(n6779), .ZN(n6775) );
  NAND2_X1 U9885 ( .A1(n6775), .A2(n6776), .ZN(n13687) );
  NAND2_X1 U9886 ( .A1(n7924), .A2(n7922), .ZN(n6778) );
  NAND2_X1 U9887 ( .A1(n9853), .A2(n6487), .ZN(n6783) );
  NAND2_X1 U9888 ( .A1(n6783), .A2(n6784), .ZN(n9895) );
  NAND3_X1 U9889 ( .A1(n12497), .A2(n9911), .A3(n6535), .ZN(n12542) );
  NAND3_X1 U9890 ( .A1(n6787), .A2(n12538), .A3(n6470), .ZN(n6786) );
  NAND4_X1 U9891 ( .A1(n12543), .A2(n6816), .A3(n12546), .A4(n6815), .ZN(n6814) );
  NAND2_X1 U9892 ( .A1(n15219), .A2(n7620), .ZN(n6819) );
  NAND2_X1 U9893 ( .A1(n15220), .A2(n7621), .ZN(n6820) );
  XNOR2_X1 U9894 ( .A(n6821), .B(P2_ADDR_REG_18__SCAN_IN), .ZN(SUB_1596_U62)
         );
  NAND3_X1 U9895 ( .A1(n6824), .A2(n6823), .A3(n6822), .ZN(n6821) );
  NAND3_X1 U9896 ( .A1(n15221), .A2(n6827), .A3(n8790), .ZN(n6822) );
  NAND2_X1 U9897 ( .A1(n6826), .A2(n15202), .ZN(n6823) );
  NAND2_X1 U9898 ( .A1(n6825), .A2(n15202), .ZN(n6824) );
  INV_X1 U9899 ( .A(n8790), .ZN(n6826) );
  INV_X1 U9900 ( .A(n15221), .ZN(n6825) );
  NAND2_X2 U9901 ( .A1(n15825), .A2(n15824), .ZN(n15823) );
  NAND2_X1 U9902 ( .A1(n8741), .A2(n6829), .ZN(n7638) );
  XNOR2_X1 U9903 ( .A(n8742), .B(n6829), .ZN(n8744) );
  AND2_X2 U9904 ( .A1(n15238), .A2(n15236), .ZN(n6831) );
  NAND2_X1 U9905 ( .A1(n6833), .A2(n15212), .ZN(n6832) );
  NAND2_X1 U9906 ( .A1(n6832), .A2(n6548), .ZN(n8769) );
  INV_X1 U9907 ( .A(n8769), .ZN(n7302) );
  NAND2_X1 U9908 ( .A1(n11120), .A2(n11119), .ZN(n12187) );
  NAND3_X1 U9909 ( .A1(n6837), .A2(n10721), .A3(n6836), .ZN(n11118) );
  NAND2_X2 U9910 ( .A1(n12090), .A2(n6839), .ZN(n13099) );
  NAND2_X1 U9911 ( .A1(n7698), .A2(n7218), .ZN(n8071) );
  NAND3_X1 U9913 ( .A1(n6842), .A2(n14324), .A3(n14338), .ZN(n14342) );
  NAND2_X1 U9914 ( .A1(n6843), .A2(n14315), .ZN(n6842) );
  OAI21_X1 U9915 ( .B1(n6848), .B2(n6845), .A(n6844), .ZN(n6843) );
  NAND2_X1 U9916 ( .A1(n14310), .A2(n7538), .ZN(n6844) );
  OAI21_X1 U9917 ( .B1(n14310), .B2(n7538), .A(n14306), .ZN(n6848) );
  NAND3_X1 U9918 ( .A1(n6859), .A2(n6858), .A3(n6856), .ZN(P1_U3242) );
  NAND3_X1 U9919 ( .A1(n6860), .A2(n11451), .A3(n14534), .ZN(n6859) );
  NAND2_X1 U9920 ( .A1(n7588), .A2(n6862), .ZN(n8855) );
  NAND2_X1 U9921 ( .A1(n8855), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8854) );
  NAND2_X1 U9922 ( .A1(n14404), .A2(n6864), .ZN(n6863) );
  NAND2_X1 U9923 ( .A1(n6863), .A2(n6614), .ZN(n6869) );
  INV_X1 U9924 ( .A(n13432), .ZN(n6876) );
  NOR2_X4 U9925 ( .A1(n13900), .A2(n14014), .ZN(n13883) );
  NAND3_X1 U9926 ( .A1(n13883), .A2(n6457), .A3(n13842), .ZN(n13841) );
  INV_X1 U9927 ( .A(n14058), .ZN(n13228) );
  NAND2_X1 U9928 ( .A1(n13725), .A2(n6604), .ZN(n8808) );
  NAND3_X1 U9929 ( .A1(n11191), .A2(n6884), .A3(n6883), .ZN(n11319) );
  NAND2_X1 U9930 ( .A1(n9530), .A2(n9496), .ZN(n10528) );
  INV_X1 U9931 ( .A(n7591), .ZN(n6894) );
  NAND2_X1 U9932 ( .A1(n6891), .A2(n12676), .ZN(n12694) );
  OAI21_X1 U9933 ( .B1(n7591), .B2(n12662), .A(n6892), .ZN(n6891) );
  INV_X1 U9934 ( .A(n12677), .ZN(n6892) );
  NAND3_X1 U9935 ( .A1(n6468), .A2(n7602), .A3(n6903), .ZN(n6896) );
  OAI21_X1 U9936 ( .B1(n15545), .B2(n6910), .A(n6906), .ZN(n7614) );
  NAND3_X1 U9937 ( .A1(n12520), .A2(n12546), .A3(n12519), .ZN(n6915) );
  NAND2_X1 U9938 ( .A1(n9742), .A2(n6640), .ZN(n9793) );
  NAND2_X1 U9939 ( .A1(n9625), .A2(n6928), .ZN(n9686) );
  NAND3_X1 U9940 ( .A1(n9535), .A2(n10657), .A3(n9536), .ZN(n9562) );
  AOI21_X2 U9941 ( .B1(n8678), .B2(n8677), .A(n7975), .ZN(n12049) );
  NAND3_X1 U9942 ( .A1(n7389), .A2(n6536), .A3(n6473), .ZN(n6931) );
  INV_X1 U9943 ( .A(n7380), .ZN(n6940) );
  NAND2_X1 U9944 ( .A1(n6946), .A2(n7996), .ZN(n7217) );
  NAND2_X2 U9945 ( .A1(n7994), .A2(n14096), .ZN(n8239) );
  NAND3_X1 U9946 ( .A1(n7992), .A2(n7994), .A3(P2_REG3_REG_1__SCAN_IN), .ZN(
        n6949) );
  NAND2_X1 U9947 ( .A1(n7992), .A2(n6588), .ZN(n6950) );
  NAND2_X1 U9948 ( .A1(n6953), .A2(n6955), .ZN(n6959) );
  NAND3_X1 U9949 ( .A1(n6958), .A2(n6961), .A3(n13889), .ZN(n6952) );
  INV_X1 U9950 ( .A(n6956), .ZN(n6954) );
  NOR2_X1 U9951 ( .A1(n13905), .A2(n13552), .ZN(n6961) );
  NAND3_X1 U9952 ( .A1(n12752), .A2(n6962), .A3(n12751), .ZN(P3_U3201) );
  AOI21_X1 U9953 ( .B1(n6963), .B2(n7372), .A(n6485), .ZN(n7369) );
  NAND2_X1 U9954 ( .A1(n10439), .A2(n6963), .ZN(n7368) );
  NOR3_X2 U9955 ( .A1(n9816), .A2(n9488), .A3(n10001), .ZN(n6966) );
  NAND4_X1 U9956 ( .A1(n6966), .A2(n6964), .A3(n6965), .A4(n7206), .ZN(n9493)
         );
  INV_X1 U9957 ( .A(n9817), .ZN(n9736) );
  NOR2_X2 U9958 ( .A1(n9637), .A2(n9638), .ZN(n6964) );
  NAND2_X1 U9959 ( .A1(n15564), .A2(n6969), .ZN(n6967) );
  OAI21_X1 U9960 ( .B1(n12604), .B2(n6981), .A(n6979), .ZN(n6984) );
  INV_X1 U9961 ( .A(n6984), .ZN(n12648) );
  OR2_X1 U9962 ( .A1(n12616), .A2(n12617), .ZN(n6985) );
  NAND3_X1 U9963 ( .A1(n6987), .A2(n7235), .A3(P3_ADDR_REG_19__SCAN_IN), .ZN(
        n7234) );
  INV_X2 U9964 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n6987) );
  OAI21_X1 U9965 ( .B1(n15500), .B2(n6987), .A(n13674), .ZN(n7438) );
  NAND2_X1 U9966 ( .A1(n7877), .A2(n6495), .ZN(n8275) );
  NAND2_X1 U9967 ( .A1(n7147), .A2(n8088), .ZN(n8105) );
  NAND2_X1 U9968 ( .A1(n7147), .A2(n6989), .ZN(n6988) );
  INV_X1 U9969 ( .A(n8107), .ZN(n6990) );
  NAND2_X1 U9970 ( .A1(n6991), .A2(n8107), .ZN(n8122) );
  NAND2_X2 U9971 ( .A1(n6994), .A2(n6992), .ZN(n14221) );
  AOI21_X2 U9972 ( .B1(n6995), .B2(n6997), .A(n6993), .ZN(n6992) );
  AND2_X2 U9973 ( .A1(n14153), .A2(n6526), .ZN(n6998) );
  OAI21_X1 U9974 ( .B1(n9141), .B2(n9301), .A(n7000), .ZN(n9148) );
  AOI21_X1 U9975 ( .B1(n10455), .B2(n7001), .A(n6574), .ZN(n7000) );
  NAND2_X1 U9976 ( .A1(n10455), .A2(n8962), .ZN(n7002) );
  NAND2_X1 U9977 ( .A1(n7579), .A2(n14122), .ZN(n7578) );
  OR2_X2 U9978 ( .A1(n13179), .A2(n7009), .ZN(n7006) );
  XNOR2_X1 U9979 ( .A(n10936), .B(n7013), .ZN(n10719) );
  NAND3_X1 U9980 ( .A1(n7485), .A2(n7483), .A3(n7484), .ZN(n11044) );
  NAND3_X2 U9981 ( .A1(n7494), .A2(n7014), .A3(n7015), .ZN(n13123) );
  NAND2_X1 U9982 ( .A1(n7022), .A2(n11710), .ZN(n7021) );
  INV_X1 U9983 ( .A(n7025), .ZN(n7022) );
  OAI21_X1 U9984 ( .B1(n11359), .B2(n8163), .A(n8162), .ZN(n11578) );
  INV_X1 U9985 ( .A(n7028), .ZN(n7029) );
  OAI21_X1 U9986 ( .B1(n8403), .B2(n7031), .A(n13781), .ZN(n7028) );
  NAND2_X1 U9987 ( .A1(n7030), .A2(n7029), .ZN(n13779) );
  NAND2_X1 U9988 ( .A1(n14096), .A2(n7993), .ZN(n8077) );
  NAND2_X1 U9989 ( .A1(n12610), .A2(n12609), .ZN(n7037) );
  NAND2_X1 U9990 ( .A1(n12594), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7038) );
  NAND2_X1 U9991 ( .A1(n11218), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n11222) );
  NAND2_X1 U9992 ( .A1(n15541), .A2(n15542), .ZN(n15540) );
  NAND2_X1 U9993 ( .A1(n10681), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n10685) );
  NAND2_X1 U9994 ( .A1(n10418), .A2(n10419), .ZN(n10430) );
  XNOR2_X1 U9995 ( .A(n12673), .B(n12661), .ZN(n12672) );
  AOI21_X1 U9996 ( .B1(n9530), .B2(n7054), .A(n7053), .ZN(n7615) );
  OAI22_X1 U9997 ( .A1(n7061), .A2(n6584), .B1(n11765), .B2(n7057), .ZN(n12894) );
  INV_X1 U9998 ( .A(n7649), .ZN(n7060) );
  NAND2_X2 U9999 ( .A1(n7069), .A2(n9504), .ZN(n9591) );
  OAI211_X2 U10000 ( .C1(n9846), .C2(n10742), .A(n7067), .B(n7064), .ZN(n9514)
         );
  AND2_X1 U10001 ( .A1(n7066), .A2(n7065), .ZN(n7064) );
  NAND3_X1 U10002 ( .A1(n7069), .A2(n9504), .A3(P3_REG3_REG_1__SCAN_IN), .ZN(
        n7065) );
  NAND2_X1 U10003 ( .A1(n12201), .A2(n11937), .ZN(n9596) );
  NAND3_X1 U10004 ( .A1(n12201), .A2(n11937), .A3(P3_REG0_REG_1__SCAN_IN), 
        .ZN(n7066) );
  NAND2_X1 U10005 ( .A1(n7069), .A2(n7068), .ZN(n7067) );
  AND2_X1 U10006 ( .A1(n11937), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7068) );
  XNOR2_X2 U10007 ( .A(n9500), .B(n9499), .ZN(n11937) );
  XNOR2_X2 U10008 ( .A(n7338), .B(n9502), .ZN(n12201) );
  NAND2_X1 U10009 ( .A1(n12877), .A2(n7076), .ZN(n7075) );
  OAI21_X2 U10010 ( .B1(n11430), .B2(n11436), .A(n9729), .ZN(n11596) );
  INV_X1 U10011 ( .A(n12319), .ZN(n12219) );
  OR2_X1 U10012 ( .A1(n12319), .A2(n7088), .ZN(n7087) );
  INV_X1 U10013 ( .A(n7966), .ZN(n7088) );
  NAND3_X1 U10014 ( .A1(n10038), .A2(n7091), .A3(n7090), .ZN(n7089) );
  NAND2_X1 U10015 ( .A1(n10873), .A2(n10915), .ZN(n7093) );
  OR2_X1 U10016 ( .A1(n12288), .A2(n7098), .ZN(n7095) );
  NAND2_X1 U10017 ( .A1(n7095), .A2(n7096), .ZN(n12311) );
  NAND2_X1 U10018 ( .A1(n11671), .A2(n7113), .ZN(n7112) );
  NAND2_X1 U10019 ( .A1(n7112), .A2(n7110), .ZN(n12208) );
  NAND3_X1 U10020 ( .A1(n7139), .A2(n9609), .A3(n9610), .ZN(n11092) );
  OAI21_X1 U10021 ( .B1(n12311), .B2(n7855), .A(n7852), .ZN(n12319) );
  AOI21_X2 U10022 ( .B1(n7873), .B2(n7871), .A(n7869), .ZN(n11671) );
  AOI21_X1 U10023 ( .B1(n12210), .B2(n12905), .A(n12276), .ZN(n12288) );
  NOR2_X1 U10024 ( .A1(n12277), .A2(n12278), .ZN(n12276) );
  XNOR2_X1 U10025 ( .A(n7119), .B(P3_IR_REG_25__SCAN_IN), .ZN(n10047) );
  NAND2_X1 U10026 ( .A1(n6411), .A2(n9604), .ZN(n12408) );
  NAND4_X2 U10027 ( .A1(n9593), .A2(n9592), .A3(n9597), .A4(n9594), .ZN(n12980) );
  OAI211_X1 U10028 ( .C1(n10863), .C2(n10862), .A(n7961), .B(n11290), .ZN(
        n7120) );
  NAND3_X1 U10029 ( .A1(n7120), .A2(n7121), .A3(n10871), .ZN(n10873) );
  NAND2_X1 U10030 ( .A1(n10867), .A2(n10868), .ZN(n7121) );
  NAND2_X1 U10031 ( .A1(n10598), .A2(n10599), .ZN(n10642) );
  NAND2_X1 U10032 ( .A1(n11594), .A2(n9749), .ZN(n11775) );
  NAND2_X1 U10033 ( .A1(n7645), .A2(n7648), .ZN(n7644) );
  OAI21_X1 U10034 ( .B1(n12209), .B2(n12918), .A(n12208), .ZN(n12277) );
  NOR2_X2 U10035 ( .A1(n15820), .A2(n8751), .ZN(n8754) );
  NAND2_X2 U10036 ( .A1(n15213), .A2(n15801), .ZN(n15212) );
  NAND2_X1 U10037 ( .A1(n8801), .A2(n13561), .ZN(n8804) );
  NAND2_X1 U10038 ( .A1(n13931), .A2(n15538), .ZN(n7146) );
  NAND2_X1 U10039 ( .A1(n14926), .A2(n7801), .ZN(n7238) );
  NAND2_X1 U10040 ( .A1(n7126), .A2(n7123), .ZN(n10046) );
  INV_X1 U10041 ( .A(n10042), .ZN(n7125) );
  OR2_X1 U10042 ( .A1(n10041), .A2(n10031), .ZN(n7126) );
  NAND2_X1 U10043 ( .A1(n7899), .A2(n12031), .ZN(n12034) );
  NAND2_X1 U10044 ( .A1(n8045), .A2(n8044), .ZN(n8054) );
  NAND2_X1 U10045 ( .A1(n7129), .A2(n6609), .ZN(n14468) );
  INV_X1 U10046 ( .A(n14457), .ZN(n7129) );
  AND2_X1 U10047 ( .A1(n9617), .A2(n10145), .ZN(n7133) );
  NAND3_X1 U10048 ( .A1(n10963), .A2(n10964), .A3(n9608), .ZN(n7139) );
  NOR2_X2 U10049 ( .A1(n7416), .A2(n10783), .ZN(n10963) );
  NOR2_X1 U10050 ( .A1(n7133), .A2(n7132), .ZN(n7131) );
  INV_X1 U10051 ( .A(n7244), .ZN(n14816) );
  INV_X1 U10052 ( .A(n10047), .ZN(n13096) );
  INV_X1 U10053 ( .A(n10004), .ZN(n10026) );
  INV_X1 U10054 ( .A(n9604), .ZN(n10789) );
  NOR2_X1 U10055 ( .A1(n6541), .A2(n7135), .ZN(n7134) );
  OAI21_X1 U10056 ( .B1(n10584), .B2(n6444), .A(n10583), .ZN(n10596) );
  NAND3_X1 U10057 ( .A1(n9483), .A2(n9482), .A3(n9699), .ZN(n9817) );
  NAND2_X1 U10058 ( .A1(n9818), .A2(n10002), .ZN(n9839) );
  OAI21_X1 U10059 ( .B1(n12841), .B2(n12544), .A(n7204), .ZN(n7203) );
  NAND3_X1 U10060 ( .A1(n7988), .A2(n8297), .A3(n7948), .ZN(n14091) );
  NAND2_X1 U10061 ( .A1(n13749), .A2(n8488), .ZN(n7924) );
  NAND2_X1 U10062 ( .A1(n13779), .A2(n8424), .ZN(n13767) );
  NAND3_X1 U10063 ( .A1(n11940), .A2(n11944), .A3(n7141), .ZN(n8811) );
  NAND2_X1 U10064 ( .A1(n8803), .A2(n8804), .ZN(n11948) );
  AND2_X2 U10065 ( .A1(n7982), .A2(n7981), .ZN(n8297) );
  NAND2_X1 U10066 ( .A1(n10109), .A2(n13542), .ZN(n10108) );
  INV_X1 U10067 ( .A(n7217), .ZN(n8651) );
  NAND2_X1 U10068 ( .A1(n7146), .A2(n7145), .ZN(P2_U3528) );
  AOI21_X1 U10069 ( .B1(n8807), .B2(n7920), .A(n13146), .ZN(n11940) );
  NAND2_X1 U10070 ( .A1(n7233), .A2(n7232), .ZN(P2_U3495) );
  NAND2_X1 U10071 ( .A1(n7951), .A2(n7949), .ZN(P2_U3527) );
  NAND2_X1 U10072 ( .A1(n7609), .A2(n11235), .ZN(n7613) );
  OAI211_X1 U10073 ( .C1(n12731), .C2(n12730), .A(n6599), .B(n7376), .ZN(
        P3_U3200) );
  NAND2_X2 U10074 ( .A1(n6512), .A2(n9582), .ZN(n12582) );
  NAND2_X2 U10075 ( .A1(n7151), .A2(n7152), .ZN(n12401) );
  INV_X1 U10076 ( .A(n13148), .ZN(n13138) );
  NAND2_X1 U10077 ( .A1(n8140), .A2(n8139), .ZN(n11359) );
  NAND2_X1 U10078 ( .A1(n13541), .A2(n8031), .ZN(n12148) );
  NAND3_X1 U10079 ( .A1(n7539), .A2(n8085), .A3(n7541), .ZN(n7147) );
  NAND2_X4 U10080 ( .A1(n12202), .A2(n8908), .ZN(n14432) );
  NAND2_X2 U10081 ( .A1(n11865), .A2(n11866), .ZN(n11864) );
  NAND2_X1 U10082 ( .A1(n8992), .A2(n7555), .ZN(n7557) );
  NAND2_X1 U10083 ( .A1(n11875), .A2(n9071), .ZN(n9094) );
  NAND2_X1 U10084 ( .A1(n7567), .A2(n9366), .ZN(n14260) );
  NAND3_X1 U10085 ( .A1(n13833), .A2(n13858), .A3(n13869), .ZN(n7150) );
  NAND2_X1 U10086 ( .A1(n9577), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U10087 ( .A1(n11199), .A2(n8051), .ZN(n10109) );
  NAND2_X1 U10088 ( .A1(n7153), .A2(n10093), .ZN(P3_U3488) );
  INV_X1 U10089 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n9481) );
  NAND2_X1 U10090 ( .A1(n9608), .A2(n12526), .ZN(n9609) );
  NAND2_X2 U10091 ( .A1(n7154), .A2(n7155), .ZN(n12425) );
  NAND2_X1 U10092 ( .A1(n10052), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10041) );
  INV_X1 U10093 ( .A(n10050), .ZN(n7156) );
  AND2_X1 U10094 ( .A1(n12298), .A2(n12297), .ZN(n7157) );
  NAND2_X4 U10095 ( .A1(n13081), .A2(n13085), .ZN(n9529) );
  AND2_X1 U10096 ( .A1(n10965), .A2(n12529), .ZN(n9608) );
  NOR2_X2 U10097 ( .A1(n9497), .A2(n9498), .ZN(n10736) );
  NAND2_X1 U10098 ( .A1(n8093), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n8114) );
  NAND2_X2 U10099 ( .A1(n8689), .A2(n8571), .ZN(n13143) );
  NAND2_X1 U10100 ( .A1(n8325), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8366) );
  AOI21_X1 U10101 ( .B1(n13485), .B2(n13484), .A(n7280), .ZN(n7279) );
  NOR2_X2 U10102 ( .A1(n8431), .A2(n8430), .ZN(n7163) );
  OAI21_X1 U10103 ( .B1(n8066), .B2(n8067), .A(n8069), .ZN(n8086) );
  NAND2_X2 U10104 ( .A1(n15222), .A2(n15501), .ZN(n15221) );
  INV_X1 U10105 ( .A(n8742), .ZN(n8741) );
  NAND2_X1 U10106 ( .A1(n7300), .A2(n15200), .ZN(n8800) );
  BUF_X1 U10108 ( .A(n13085), .Z(n7168) );
  NAND2_X1 U10109 ( .A1(n12765), .A2(n7170), .ZN(P3_U3204) );
  OR2_X1 U10110 ( .A1(n12581), .A2(n10805), .ZN(n10965) );
  INV_X2 U10111 ( .A(n9529), .ZN(n9804) );
  NAND2_X1 U10112 ( .A1(n7663), .A2(n7662), .ZN(n12841) );
  NAND2_X4 U10113 ( .A1(n7172), .A2(n9493), .ZN(n13085) );
  INV_X1 U10114 ( .A(n13801), .ZN(n8403) );
  OAI21_X1 U10115 ( .B1(n8345), .B2(n8359), .A(n7358), .ZN(n8382) );
  INV_X1 U10116 ( .A(n14814), .ZN(n7173) );
  XNOR2_X2 U10117 ( .A(n8897), .B(n7174), .ZN(n12202) );
  INV_X1 U10118 ( .A(n7345), .ZN(n7344) );
  NAND2_X1 U10119 ( .A1(n7341), .A2(n7175), .ZN(n8314) );
  INV_X1 U10120 ( .A(n7176), .ZN(n7175) );
  OAI21_X1 U10121 ( .B1(n7343), .B2(n7959), .A(n6613), .ZN(n7176) );
  INV_X4 U10122 ( .A(n8209), .ZN(n7875) );
  NAND2_X1 U10123 ( .A1(n11823), .A2(n12572), .ZN(n7178) );
  NOR2_X1 U10124 ( .A1(n7181), .A2(n7180), .ZN(n7179) );
  AOI21_X1 U10125 ( .B1(n7326), .B2(n12544), .A(n12801), .ZN(n12503) );
  INV_X1 U10126 ( .A(n7742), .ZN(n7741) );
  NOR2_X2 U10127 ( .A1(n13111), .A2(n7184), .ZN(n12003) );
  AND2_X2 U10128 ( .A1(n7489), .A2(n7490), .ZN(n7348) );
  INV_X1 U10129 ( .A(n11972), .ZN(n7496) );
  OAI21_X1 U10130 ( .B1(n7877), .B2(n7346), .A(n7344), .ZN(n8312) );
  NAND2_X1 U10131 ( .A1(n8054), .A2(n8053), .ZN(n7542) );
  NAND2_X1 U10132 ( .A1(n7542), .A2(n7540), .ZN(n7539) );
  MUX2_X1 U10133 ( .A(n14294), .B(n14293), .S(n14436), .Z(n14296) );
  INV_X2 U10134 ( .A(n14312), .ZN(n14436) );
  OAI21_X1 U10135 ( .B1(n14424), .B2(n10825), .A(n7185), .ZN(n14312) );
  NAND2_X1 U10136 ( .A1(n14424), .A2(n14483), .ZN(n7185) );
  NAND2_X1 U10137 ( .A1(n13716), .A2(n8525), .ZN(n13703) );
  NAND2_X1 U10138 ( .A1(n13767), .A2(n8438), .ZN(n7930) );
  INV_X1 U10139 ( .A(n8297), .ZN(n8278) );
  NAND3_X1 U10140 ( .A1(n7988), .A2(n8297), .A3(n8011), .ZN(n7404) );
  NAND2_X1 U10141 ( .A1(n15590), .A2(n15589), .ZN(n7202) );
  INV_X1 U10142 ( .A(n10582), .ZN(n10584) );
  NAND2_X1 U10143 ( .A1(n7217), .A2(n7216), .ZN(n7215) );
  NAND2_X1 U10144 ( .A1(n7221), .A2(n7219), .ZN(n13800) );
  NAND3_X1 U10145 ( .A1(n8004), .A2(n8006), .A3(n8005), .ZN(n8231) );
  NAND3_X1 U10146 ( .A1(n7237), .A2(n7236), .A3(P2_ADDR_REG_19__SCAN_IN), .ZN(
        n7210) );
  NAND2_X1 U10147 ( .A1(n8207), .A2(n8206), .ZN(n8253) );
  NAND2_X1 U10148 ( .A1(n14052), .A2(n6638), .ZN(P2_U3492) );
  NAND2_X1 U10149 ( .A1(n7930), .A2(n7929), .ZN(n12052) );
  NAND2_X1 U10150 ( .A1(n13877), .A2(n7936), .ZN(n7221) );
  CLKBUF_X3 U10151 ( .A(n9617), .Z(n9956) );
  XNOR2_X1 U10152 ( .A(n12524), .B(n12220), .ZN(n11288) );
  INV_X1 U10153 ( .A(n12772), .ZN(n7223) );
  NAND2_X1 U10154 ( .A1(n9960), .A2(n9959), .ZN(n9976) );
  INV_X4 U10155 ( .A(n8039), .ZN(n8209) );
  NAND2_X1 U10156 ( .A1(n12003), .A2(n7482), .ZN(n7479) );
  AND4_X1 U10157 ( .A1(n10861), .A2(n10860), .A3(n10990), .A4(n11288), .ZN(
        n7961) );
  INV_X1 U10158 ( .A(n11637), .ZN(n7873) );
  NAND2_X1 U10159 ( .A1(n13717), .A2(n13718), .ZN(n13716) );
  NAND2_X1 U10160 ( .A1(n11551), .A2(n14318), .ZN(n11472) );
  AOI21_X1 U10161 ( .B1(n14861), .B2(n7250), .A(n7248), .ZN(n7244) );
  OAI21_X1 U10162 ( .B1(n14861), .B2(n12137), .A(n12136), .ZN(n14828) );
  NOR2_X1 U10163 ( .A1(n7243), .A2(n7245), .ZN(n14792) );
  NAND2_X4 U10164 ( .A1(n6434), .A2(n7875), .ZN(n14476) );
  NAND2_X1 U10165 ( .A1(n10257), .A2(n7264), .ZN(n7263) );
  NAND2_X1 U10166 ( .A1(n7268), .A2(n7266), .ZN(n12121) );
  INV_X1 U10167 ( .A(n7267), .ZN(n7266) );
  OAI21_X1 U10168 ( .B1(n11844), .B2(n7269), .A(n7777), .ZN(n7267) );
  NAND2_X1 U10169 ( .A1(n11928), .A2(n11845), .ZN(n7268) );
  INV_X1 U10170 ( .A(n11845), .ZN(n7269) );
  NAND2_X1 U10171 ( .A1(n7272), .A2(n6622), .ZN(n9061) );
  NAND2_X1 U10172 ( .A1(n8863), .A2(n6639), .ZN(n9204) );
  NAND2_X1 U10173 ( .A1(n9231), .A2(n7274), .ZN(n9274) );
  INV_X1 U10174 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n7277) );
  NAND2_X1 U10175 ( .A1(n9310), .A2(n6651), .ZN(n9370) );
  OAI21_X2 U10176 ( .B1(n7279), .B2(n6531), .A(n13533), .ZN(n13583) );
  NAND3_X1 U10177 ( .A1(n13527), .A2(n13525), .A3(n13526), .ZN(n7280) );
  OR2_X1 U10178 ( .A1(n13381), .A2(n7284), .ZN(n7283) );
  NAND2_X1 U10179 ( .A1(n13362), .A2(n7290), .ZN(n7288) );
  NAND2_X1 U10180 ( .A1(n7288), .A2(n7289), .ZN(n7900) );
  NAND2_X1 U10181 ( .A1(n7288), .A2(n7286), .ZN(n13369) );
  INV_X1 U10182 ( .A(n13361), .ZN(n7291) );
  INV_X1 U10183 ( .A(n13413), .ZN(n7298) );
  INV_X1 U10184 ( .A(n7299), .ZN(n8764) );
  NAND2_X1 U10185 ( .A1(n12584), .A2(n10756), .ZN(n12396) );
  INV_X1 U10186 ( .A(n12461), .ZN(n7318) );
  NAND2_X1 U10187 ( .A1(n12464), .A2(n12538), .ZN(n7325) );
  AOI21_X1 U10188 ( .B1(n7808), .B2(n11461), .A(n7332), .ZN(n7331) );
  NAND2_X1 U10189 ( .A1(n7877), .A2(n7342), .ZN(n7341) );
  NAND2_X1 U10190 ( .A1(n13155), .A2(n11995), .ZN(n11997) );
  NAND3_X1 U10191 ( .A1(n7352), .A2(n7353), .A3(n7349), .ZN(n13218) );
  NAND2_X1 U10192 ( .A1(n7368), .A2(n7369), .ZN(n11226) );
  NAND2_X1 U10193 ( .A1(n7694), .A2(n6598), .ZN(n7386) );
  NAND3_X1 U10194 ( .A1(n6473), .A2(n7389), .A3(n8673), .ZN(n7388) );
  NAND2_X1 U10195 ( .A1(n7394), .A2(n12049), .ZN(n7393) );
  NAND2_X1 U10196 ( .A1(n7406), .A2(n7405), .ZN(P3_U3454) );
  OR2_X1 U10197 ( .A1(n15654), .A2(n9965), .ZN(n7405) );
  NAND2_X1 U10198 ( .A1(n13005), .A2(n15654), .ZN(n7406) );
  AOI21_X1 U10199 ( .B1(n12934), .B2(n6643), .A(n7408), .ZN(n7407) );
  INV_X1 U10200 ( .A(n7415), .ZN(n7414) );
  NAND2_X1 U10201 ( .A1(n7419), .A2(n7417), .ZN(n12946) );
  OAI21_X1 U10202 ( .B1(n7841), .B2(n7839), .A(n11436), .ZN(n7430) );
  NAND2_X1 U10203 ( .A1(n7448), .A2(n7446), .ZN(n10953) );
  NAND2_X2 U10204 ( .A1(n7455), .A2(n7454), .ZN(n14295) );
  NAND3_X1 U10205 ( .A1(n7456), .A2(n11406), .A3(n11051), .ZN(n11415) );
  INV_X1 U10206 ( .A(n7457), .ZN(n11350) );
  NOR2_X2 U10207 ( .A1(n7461), .A2(n7953), .ZN(n14974) );
  NAND3_X1 U10208 ( .A1(n7588), .A2(n7463), .A3(n7586), .ZN(n8866) );
  NAND2_X1 U10209 ( .A1(n7588), .A2(n7586), .ZN(n8825) );
  NAND4_X1 U10210 ( .A1(n7486), .A2(n10712), .A3(n10710), .A4(n10711), .ZN(
        n7484) );
  NAND3_X1 U10211 ( .A1(n7487), .A2(n13237), .A3(n7486), .ZN(n7485) );
  NAND2_X1 U10212 ( .A1(n13123), .A2(n7491), .ZN(n7489) );
  NOR2_X1 U10213 ( .A1(n12152), .A2(n13897), .ZN(n10377) );
  NAND2_X2 U10214 ( .A1(n7493), .A2(n13571), .ZN(n10717) );
  INV_X1 U10215 ( .A(n13285), .ZN(n7492) );
  NOR2_X1 U10216 ( .A1(n11203), .A2(n7493), .ZN(n11204) );
  OAI211_X1 U10217 ( .C1(n11012), .C2(n7493), .A(n11009), .B(n11008), .ZN(
        n15519) );
  NOR2_X1 U10218 ( .A1(n14029), .A2(n7493), .ZN(n11715) );
  NAND3_X1 U10219 ( .A1(n7498), .A2(n11976), .A3(n7500), .ZN(n7495) );
  NAND2_X1 U10220 ( .A1(n7499), .A2(n7501), .ZN(n7498) );
  OAI21_X1 U10221 ( .B1(n13099), .B2(n7500), .A(n7497), .ZN(n12077) );
  INV_X1 U10222 ( .A(n11666), .ZN(n7504) );
  NAND3_X1 U10223 ( .A1(n7503), .A2(n11957), .A3(n7502), .ZN(n11958) );
  NAND2_X1 U10224 ( .A1(n11666), .A2(n11953), .ZN(n7503) );
  NAND2_X1 U10225 ( .A1(n14445), .A2(n14444), .ZN(n7506) );
  AND2_X1 U10226 ( .A1(n14444), .A2(n14420), .ZN(n7507) );
  NAND2_X1 U10227 ( .A1(n7511), .A2(n6618), .ZN(n14417) );
  NAND2_X1 U10228 ( .A1(n7524), .A2(n7525), .ZN(n7522) );
  NAND2_X1 U10229 ( .A1(n14355), .A2(n7530), .ZN(n7529) );
  AND2_X1 U10230 ( .A1(n8069), .A2(n6400), .ZN(n7540) );
  OAI21_X1 U10231 ( .B1(n14792), .B2(n7547), .A(n7545), .ZN(n7544) );
  NAND2_X1 U10232 ( .A1(n14792), .A2(n14797), .ZN(n14791) );
  NAND2_X2 U10233 ( .A1(n6435), .A2(n8209), .ZN(n12036) );
  NAND2_X1 U10234 ( .A1(n7557), .A2(n6606), .ZN(n9018) );
  INV_X1 U10235 ( .A(n14105), .ZN(n7564) );
  NAND2_X1 U10236 ( .A1(n14178), .A2(n7568), .ZN(n7565) );
  NAND2_X1 U10237 ( .A1(n7565), .A2(n7566), .ZN(n14116) );
  NAND2_X1 U10238 ( .A1(n14178), .A2(n14179), .ZN(n7567) );
  OAI21_X2 U10239 ( .B1(n14221), .B2(n7573), .A(n7571), .ZN(n14241) );
  NAND2_X2 U10240 ( .A1(n14204), .A2(n7581), .ZN(n14252) );
  NAND3_X1 U10241 ( .A1(n8896), .A2(n8922), .A3(n10605), .ZN(n10606) );
  NAND2_X1 U10242 ( .A1(n10606), .A2(n8922), .ZN(n10757) );
  NOR2_X1 U10243 ( .A1(n9226), .A2(n7781), .ZN(n8840) );
  NAND2_X1 U10244 ( .A1(n12121), .A2(n12120), .ZN(n15005) );
  XNOR2_X1 U10245 ( .A(n8120), .B(n8122), .ZN(n10180) );
  NAND2_X1 U10246 ( .A1(n11476), .A2(n11475), .ZN(n11556) );
  OR2_X2 U10247 ( .A1(n14295), .A2(n15276), .ZN(n15263) );
  NOR2_X1 U10248 ( .A1(n7592), .A2(n12683), .ZN(n7591) );
  NAND2_X1 U10249 ( .A1(n10664), .A2(n7596), .ZN(n7595) );
  NAND3_X1 U10250 ( .A1(n7595), .A2(n10444), .A3(n7594), .ZN(n10446) );
  INV_X1 U10251 ( .A(n12588), .ZN(n7603) );
  NAND3_X1 U10252 ( .A1(n12588), .A2(n7605), .A3(n12646), .ZN(n7599) );
  INV_X1 U10253 ( .A(n11241), .ZN(n7609) );
  NAND2_X1 U10254 ( .A1(n11241), .A2(n6482), .ZN(n7611) );
  NAND2_X1 U10255 ( .A1(n7613), .A2(n15583), .ZN(n11242) );
  INV_X1 U10256 ( .A(n15543), .ZN(n7617) );
  INV_X1 U10257 ( .A(P2_ADDR_REG_11__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U10258 ( .A1(n15823), .A2(n6483), .ZN(n7627) );
  NAND3_X1 U10259 ( .A1(n7628), .A2(n7629), .A3(n7627), .ZN(n15211) );
  NAND2_X1 U10260 ( .A1(n15823), .A2(n8756), .ZN(n8760) );
  INV_X1 U10261 ( .A(n8756), .ZN(n7630) );
  INV_X1 U10262 ( .A(n7631), .ZN(n15209) );
  NAND2_X1 U10263 ( .A1(n8740), .A2(n8739), .ZN(n7635) );
  NAND2_X2 U10264 ( .A1(n15227), .A2(n8775), .ZN(n15231) );
  NAND2_X1 U10265 ( .A1(n8749), .A2(n8709), .ZN(n7642) );
  AND2_X1 U10266 ( .A1(n7646), .A2(n9653), .ZN(n7645) );
  NAND2_X1 U10267 ( .A1(n12809), .A2(n7657), .ZN(n7653) );
  NAND2_X1 U10268 ( .A1(n12764), .A2(n10104), .ZN(n7666) );
  NAND2_X1 U10269 ( .A1(n7666), .A2(n7664), .ZN(P3_U3456) );
  NAND2_X1 U10270 ( .A1(n7667), .A2(n7668), .ZN(n13075) );
  INV_X1 U10271 ( .A(n9491), .ZN(n7667) );
  NAND2_X1 U10272 ( .A1(n7952), .A2(n7670), .ZN(n9850) );
  NAND3_X1 U10273 ( .A1(n7677), .A2(n7676), .A3(n8653), .ZN(n11003) );
  NAND2_X1 U10274 ( .A1(n7681), .A2(n7679), .ZN(n13906) );
  INV_X1 U10275 ( .A(n7680), .ZN(n7679) );
  OAI21_X1 U10276 ( .B1(n7685), .B2(n6407), .A(n8666), .ZN(n7680) );
  NOR2_X1 U10277 ( .A1(n7685), .A2(n7684), .ZN(n7682) );
  NAND2_X1 U10278 ( .A1(n9954), .A2(n7702), .ZN(n7699) );
  NAND2_X1 U10279 ( .A1(n7699), .A2(n7700), .ZN(n9985) );
  NAND3_X1 U10280 ( .A1(n7708), .A2(n12546), .A3(n6471), .ZN(n7707) );
  INV_X1 U10281 ( .A(n9547), .ZN(n7737) );
  INV_X1 U10282 ( .A(n9895), .ZN(n7758) );
  INV_X1 U10283 ( .A(n7760), .ZN(n13865) );
  NAND2_X1 U10284 ( .A1(n7761), .A2(n6492), .ZN(n14042) );
  NAND2_X1 U10285 ( .A1(n13925), .A2(n7763), .ZN(n7761) );
  NAND2_X1 U10286 ( .A1(n7762), .A2(n6491), .ZN(n13926) );
  NAND2_X1 U10287 ( .A1(n13925), .A2(n7764), .ZN(n7762) );
  NAND2_X1 U10288 ( .A1(n11583), .A2(n7765), .ZN(n7768) );
  INV_X1 U10289 ( .A(n7767), .ZN(n7766) );
  INV_X1 U10290 ( .A(n7768), .ZN(n11816) );
  NAND2_X1 U10291 ( .A1(n13707), .A2(n7770), .ZN(n13682) );
  INV_X1 U10292 ( .A(n7775), .ZN(n7774) );
  NAND2_X1 U10293 ( .A1(n14749), .A2(n7791), .ZN(n7789) );
  AOI21_X1 U10294 ( .B1(n14749), .B2(n14796), .A(n14797), .ZN(n14799) );
  INV_X1 U10295 ( .A(n7794), .ZN(n7790) );
  INV_X1 U10296 ( .A(n14796), .ZN(n7792) );
  INV_X1 U10297 ( .A(n7793), .ZN(n14752) );
  INV_X1 U10298 ( .A(n14750), .ZN(n7796) );
  NAND3_X1 U10299 ( .A1(n8930), .A2(n15261), .A3(n7797), .ZN(n14289) );
  NAND2_X2 U10300 ( .A1(n15182), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U10301 ( .A1(n7808), .A2(n12402), .ZN(n10586) );
  NOR2_X1 U10302 ( .A1(n10459), .A2(n7808), .ZN(n12525) );
  XNOR2_X1 U10303 ( .A(n10589), .B(n7808), .ZN(n10744) );
  NAND2_X1 U10304 ( .A1(n12791), .A2(n7831), .ZN(n7829) );
  OAI21_X1 U10305 ( .B1(n12791), .B2(n12506), .A(n12509), .ZN(n12780) );
  INV_X1 U10306 ( .A(n10022), .ZN(n10024) );
  NAND2_X1 U10307 ( .A1(n12219), .A2(n7860), .ZN(n7859) );
  MUX2_X1 U10308 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n8209), .Z(n8015) );
  MUX2_X1 U10309 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8209), .Z(n8106) );
  MUX2_X1 U10310 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8209), .Z(n8123) );
  MUX2_X1 U10311 ( .A(n9511), .B(n9512), .S(n8209), .Z(n10142) );
  MUX2_X1 U10312 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8209), .Z(n8144) );
  MUX2_X1 U10313 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n8017), .Z(n8167) );
  MUX2_X1 U10314 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n8209), .Z(n8191) );
  MUX2_X1 U10315 ( .A(n9915), .B(SI_24_), .S(n7875), .Z(n13098) );
  NAND2_X1 U10316 ( .A1(n8193), .A2(n8192), .ZN(n8207) );
  NAND2_X1 U10317 ( .A1(n12029), .A2(n12028), .ZN(n7899) );
  NAND3_X1 U10318 ( .A1(n13294), .A2(n13672), .A3(n13578), .ZN(n13285) );
  NAND2_X1 U10319 ( .A1(n7904), .A2(n6607), .ZN(n13339) );
  NAND2_X1 U10320 ( .A1(n7909), .A2(n7910), .ZN(n13400) );
  AOI21_X1 U10321 ( .B1(n7921), .B2(n13561), .A(n13836), .ZN(n7920) );
  INV_X1 U10322 ( .A(n11810), .ZN(n7928) );
  NAND2_X1 U10323 ( .A1(n10108), .A2(n7945), .ZN(n7944) );
  NAND2_X1 U10324 ( .A1(n7944), .A2(n7942), .ZN(n11188) );
  OR2_X1 U10325 ( .A1(n7946), .A2(n13543), .ZN(n7943) );
  NAND2_X1 U10326 ( .A1(n11006), .A2(n13543), .ZN(n11186) );
  NAND2_X1 U10327 ( .A1(n8297), .A2(n7988), .ZN(n8010) );
  NAND2_X1 U10328 ( .A1(n13753), .A2(n13758), .ZN(n13754) );
  XNOR2_X1 U10329 ( .A(n6401), .B(n13626), .ZN(n15828) );
  NAND4_X4 U10330 ( .A1(n9567), .A2(n9566), .A3(n9565), .A4(n9564), .ZN(n12581) );
  OR2_X2 U10331 ( .A1(n12363), .A2(n9563), .ZN(n9564) );
  INV_X1 U10332 ( .A(n8753), .ZN(n8755) );
  CLKBUF_X1 U10333 ( .A(n11075), .Z(n14142) );
  OR2_X1 U10334 ( .A1(n9596), .A2(n9595), .ZN(n9597) );
  AND2_X1 U10335 ( .A1(n12580), .A2(n7155), .ZN(n9607) );
  INV_X2 U10336 ( .A(n10296), .ZN(n8046) );
  XOR2_X1 U10337 ( .A(n14830), .B(n14828), .Z(n15072) );
  AND2_X1 U10338 ( .A1(n10053), .A2(n10052), .ZN(n10121) );
  NAND2_X1 U10339 ( .A1(n13931), .A2(n15533), .ZN(n8704) );
  NAND2_X1 U10340 ( .A1(n12384), .A2(n6602), .ZN(n12381) );
  INV_X1 U10341 ( .A(n13883), .ZN(n13899) );
  AND2_X1 U10342 ( .A1(n13521), .A2(n13483), .ZN(n13484) );
  AND2_X1 U10343 ( .A1(n13290), .A2(n13289), .ZN(n13308) );
  OR3_X1 U10344 ( .A1(n13524), .A2(n13523), .A3(n13522), .ZN(n13525) );
  INV_X1 U10345 ( .A(n6520), .ZN(n12891) );
  OAI22_X1 U10346 ( .A1(n13435), .A2(n13434), .B1(n13441), .B2(n13440), .ZN(
        n13444) );
  INV_X1 U10347 ( .A(n13676), .ZN(n14043) );
  OAI21_X1 U10348 ( .B1(n8700), .B2(n13908), .A(n8694), .ZN(n8695) );
  INV_X1 U10349 ( .A(n14516), .ZN(n11844) );
  NAND2_X1 U10350 ( .A1(n8588), .A2(n8579), .ZN(n8613) );
  AND2_X1 U10351 ( .A1(n8003), .A2(n8002), .ZN(n7955) );
  OR2_X1 U10352 ( .A1(n13012), .A2(n12822), .ZN(n7956) );
  AND2_X1 U10353 ( .A1(n9449), .A2(n14273), .ZN(n7957) );
  AND3_X1 U10354 ( .A1(n10030), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_IR_REG_24__SCAN_IN), .ZN(n7958) );
  AND2_X1 U10355 ( .A1(n8276), .A2(n8262), .ZN(n7959) );
  INV_X1 U10356 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n15184) );
  INV_X1 U10357 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n8780) );
  AND2_X1 U10358 ( .A1(n14510), .A2(n11479), .ZN(n7963) );
  OR2_X1 U10359 ( .A1(n12317), .A2(n12569), .ZN(n7966) );
  AND3_X1 U10360 ( .A1(n12380), .A2(n12379), .A3(n12378), .ZN(n7967) );
  OR2_X1 U10361 ( .A1(n14188), .A2(n14187), .ZN(n7968) );
  INV_X1 U10362 ( .A(n14973), .ZN(n12095) );
  OR2_X1 U10363 ( .A1(n13996), .A2(n13598), .ZN(n7969) );
  AND2_X1 U10364 ( .A1(n13996), .A2(n13397), .ZN(n7970) );
  AND2_X1 U10365 ( .A1(n14755), .A2(n14812), .ZN(n7971) );
  AND2_X1 U10366 ( .A1(n14787), .A2(n14761), .ZN(n7972) );
  NOR4_X1 U10367 ( .A1(n13561), .A2(n13560), .A3(n13559), .A4(n13558), .ZN(
        n7973) );
  INV_X1 U10368 ( .A(n12971), .ZN(n10091) );
  AND3_X2 U10369 ( .A1(n10073), .A2(n10507), .A3(n10072), .ZN(n15665) );
  NOR2_X1 U10370 ( .A1(n14891), .A2(n14544), .ZN(n7974) );
  NOR2_X1 U10371 ( .A1(n13432), .A2(n13783), .ZN(n7975) );
  OR2_X1 U10372 ( .A1(n13610), .A2(n6751), .ZN(n7976) );
  INV_X1 U10373 ( .A(n15335), .ZN(n11475) );
  NOR2_X1 U10374 ( .A1(n8375), .A2(n7970), .ZN(n8376) );
  INV_X1 U10375 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n9477) );
  INV_X1 U10376 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8301) );
  INV_X1 U10377 ( .A(n8613), .ZN(n8614) );
  NAND2_X1 U10378 ( .A1(n14190), .A2(n14275), .ZN(n9217) );
  INV_X1 U10379 ( .A(n9204), .ZN(n8864) );
  AND3_X1 U10380 ( .A1(n8821), .A2(n8820), .A3(n8843), .ZN(n8822) );
  NAND2_X1 U10381 ( .A1(n12401), .A2(n6444), .ZN(n10583) );
  OR2_X1 U10382 ( .A1(n12932), .A2(n12795), .ZN(n9969) );
  AND2_X1 U10383 ( .A1(n10764), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n9765) );
  INV_X1 U10384 ( .A(n12150), .ZN(n8031) );
  OAI21_X1 U10385 ( .B1(n13540), .B2(n7962), .A(n7976), .ZN(n8652) );
  INV_X1 U10386 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n7984) );
  NAND2_X1 U10387 ( .A1(n9306), .A2(n9305), .ZN(n9307) );
  INV_X1 U10388 ( .A(n9267), .ZN(n9268) );
  INV_X1 U10389 ( .A(n9266), .ZN(n9269) );
  INV_X1 U10390 ( .A(n9220), .ZN(n9221) );
  INV_X1 U10391 ( .A(n8975), .ZN(n8976) );
  INV_X1 U10392 ( .A(n14753), .ZN(n14793) );
  INV_X1 U10393 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n9076) );
  INV_X1 U10394 ( .A(n8205), .ZN(n8206) );
  NOR2_X1 U10395 ( .A1(n12230), .A2(n12836), .ZN(n10019) );
  INV_X1 U10396 ( .A(n12564), .ZN(n12385) );
  AND2_X1 U10397 ( .A1(n10123), .A2(n9529), .ZN(n10878) );
  INV_X1 U10398 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n9499) );
  INV_X1 U10399 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n9480) );
  INV_X1 U10400 ( .A(n14009), .ZN(n8688) );
  INV_X1 U10401 ( .A(n8611), .ZN(n8612) );
  NAND2_X1 U10402 ( .A1(n6405), .A2(n13672), .ZN(n10568) );
  INV_X1 U10403 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n9897) );
  OR2_X1 U10404 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  INV_X1 U10405 ( .A(n9252), .ZN(n9253) );
  INV_X1 U10406 ( .A(n14974), .ZN(n14991) );
  INV_X1 U10407 ( .A(n14787), .ZN(n15046) );
  NAND2_X1 U10408 ( .A1(n8338), .A2(SI_17_), .ZN(n8360) );
  NOR2_X1 U10409 ( .A1(n8735), .A2(n8736), .ZN(n8720) );
  INV_X1 U10410 ( .A(n12887), .ZN(n12485) );
  OR2_X1 U10411 ( .A1(n12215), .A2(n12485), .ZN(n12216) );
  OR2_X1 U10412 ( .A1(n10099), .A2(n10098), .ZN(n10541) );
  INV_X1 U10413 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n10621) );
  INV_X1 U10414 ( .A(n15595), .ZN(n15576) );
  OR2_X1 U10415 ( .A1(n10085), .A2(n12513), .ZN(n10529) );
  NOR2_X1 U10416 ( .A1(n10064), .A2(n10063), .ZN(n10100) );
  INV_X1 U10417 ( .A(n10081), .ZN(n9981) );
  OR2_X1 U10418 ( .A1(n10505), .A2(n10100), .ZN(n10540) );
  AND2_X1 U10419 ( .A1(n10242), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n9679) );
  INV_X1 U10420 ( .A(n12020), .ZN(n12021) );
  INV_X1 U10421 ( .A(n11667), .ZN(n11665) );
  INV_X1 U10422 ( .A(n13275), .ZN(n13263) );
  OR2_X1 U10423 ( .A1(n13260), .A2(n8595), .ZN(n8542) );
  INV_X1 U10424 ( .A(n10300), .ZN(n10323) );
  INV_X1 U10425 ( .A(n13766), .ZN(n8677) );
  AND2_X1 U10426 ( .A1(n13536), .A2(n13535), .ZN(n13760) );
  OR3_X1 U10427 ( .A1(n14021), .A2(n14020), .A3(n14019), .ZN(n14083) );
  AND2_X1 U10428 ( .A1(n10884), .A2(n13570), .ZN(n15524) );
  OR2_X1 U10429 ( .A1(n8235), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n8263) );
  INV_X1 U10430 ( .A(n14550), .ZN(n14343) );
  INV_X1 U10431 ( .A(n15011), .ZN(n14370) );
  INV_X1 U10432 ( .A(n14833), .ZN(n14216) );
  INV_X1 U10433 ( .A(n14262), .ZN(n14279) );
  OR2_X1 U10434 ( .A1(n14873), .A2(n6439), .ZN(n9300) );
  INV_X1 U10435 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n15782) );
  INV_X1 U10436 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n14207) );
  INV_X1 U10437 ( .A(n11476), .ZN(n11558) );
  INV_X1 U10438 ( .A(n15008), .ZN(n14853) );
  OR2_X1 U10439 ( .A1(n6408), .A2(n10826), .ZN(n14994) );
  NOR2_X2 U10440 ( .A1(n10824), .A2(n9446), .ZN(n15336) );
  NAND2_X1 U10441 ( .A1(n9429), .A2(n9428), .ZN(n11462) );
  AND3_X1 U10442 ( .A1(n10182), .A2(n9427), .A3(n9426), .ZN(n9439) );
  AND2_X1 U10443 ( .A1(n8381), .A2(n8360), .ZN(n8379) );
  AND2_X1 U10444 ( .A1(n10547), .A2(n10546), .ZN(n12347) );
  INV_X1 U10445 ( .A(n15570), .ZN(n15586) );
  NAND2_X1 U10446 ( .A1(n10088), .A2(n10087), .ZN(n12978) );
  INV_X1 U10447 ( .A(n12828), .ZN(n12913) );
  INV_X1 U10448 ( .A(n15610), .ZN(n12912) );
  INV_X1 U10449 ( .A(n12767), .ZN(n10092) );
  AND2_X1 U10450 ( .A1(n15665), .A2(n12933), .ZN(n12968) );
  INV_X1 U10451 ( .A(n12838), .ZN(n12981) );
  OR2_X1 U10452 ( .A1(n12978), .A2(n6643), .ZN(n15630) );
  AOI21_X1 U10453 ( .B1(n10202), .B2(n10164), .A(n10039), .ZN(n10502) );
  AND2_X1 U10454 ( .A1(n9852), .A2(n9838), .ZN(n9851) );
  AND2_X1 U10455 ( .A1(n10567), .A2(n13574), .ZN(n13275) );
  INV_X1 U10456 ( .A(n15492), .ZN(n15460) );
  INV_X1 U10457 ( .A(n13643), .ZN(n15482) );
  AND2_X1 U10458 ( .A1(n10323), .A2(n10322), .ZN(n15486) );
  AND2_X1 U10459 ( .A1(n10563), .A2(n8605), .ZN(n13878) );
  NAND2_X2 U10460 ( .A1(n8650), .A2(n13843), .ZN(n13913) );
  INV_X1 U10461 ( .A(n15506), .ZN(n10561) );
  AND2_X1 U10462 ( .A1(n8236), .A2(n8263), .ZN(n11754) );
  AND2_X1 U10463 ( .A1(n10293), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14262) );
  INV_X1 U10464 ( .A(n10605), .ZN(n10609) );
  NAND2_X1 U10465 ( .A1(n12116), .A2(n12115), .ZN(n12117) );
  AND2_X1 U10466 ( .A1(n10245), .A2(n15193), .ZN(n15010) );
  INV_X1 U10467 ( .A(n14504), .ZN(n11346) );
  NAND2_X2 U10468 ( .A1(n14762), .A2(n14977), .ZN(n14993) );
  INV_X1 U10469 ( .A(n14743), .ZN(n15028) );
  AND2_X1 U10470 ( .A1(n10816), .A2(n10815), .ZN(n15296) );
  INV_X1 U10471 ( .A(n9439), .ZN(n10184) );
  INV_X1 U10472 ( .A(n8772), .ZN(n8773) );
  AND2_X1 U10473 ( .A1(n10133), .A2(n10132), .ZN(n15539) );
  NAND2_X1 U10474 ( .A1(n10544), .A2(n10543), .ZN(n12349) );
  AND2_X1 U10475 ( .A1(n12366), .A2(n10017), .ZN(n12374) );
  INV_X1 U10476 ( .A(n12837), .ZN(n12569) );
  INV_X1 U10477 ( .A(n11677), .ZN(n12918) );
  INV_X1 U10478 ( .A(n15539), .ZN(n15605) );
  INV_X1 U10479 ( .A(n15591), .ZN(n12730) );
  NAND2_X1 U10480 ( .A1(n15616), .A2(n10773), .ZN(n12922) );
  INV_X1 U10481 ( .A(n12789), .ZN(n11276) );
  INV_X1 U10482 ( .A(n15665), .ZN(n15663) );
  NAND2_X1 U10483 ( .A1(n15654), .A2(n15630), .ZN(n13065) );
  INV_X1 U10484 ( .A(n15654), .ZN(n15653) );
  AND2_X2 U10485 ( .A1(n10103), .A2(n10543), .ZN(n15654) );
  INV_X1 U10486 ( .A(n12548), .ZN(n12743) );
  INV_X1 U10487 ( .A(SI_14_), .ZN(n10497) );
  INV_X1 U10488 ( .A(n13956), .ZN(n13758) );
  AND2_X1 U10489 ( .A1(n10566), .A2(n13843), .ZN(n13227) );
  INV_X1 U10490 ( .A(n13530), .ZN(n13679) );
  INV_X1 U10491 ( .A(n13430), .ZN(n13783) );
  INV_X1 U10492 ( .A(n13345), .ZN(n13604) );
  NAND2_X1 U10493 ( .A1(n15432), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15468) );
  INV_X1 U10494 ( .A(n15368), .ZN(n15500) );
  INV_X1 U10495 ( .A(n13913), .ZN(n13894) );
  AND2_X1 U10496 ( .A1(n11724), .A2(n8687), .ZN(n13908) );
  AND2_X2 U10497 ( .A1(n8810), .A2(n10561), .ZN(n15538) );
  AND2_X2 U10498 ( .A1(n8810), .A2(n15506), .ZN(n15533) );
  INV_X1 U10499 ( .A(n15533), .ZN(n15531) );
  NOR2_X1 U10500 ( .A1(n15509), .A2(n15502), .ZN(n15503) );
  INV_X1 U10501 ( .A(n15503), .ZN(n15504) );
  INV_X1 U10502 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10767) );
  XNOR2_X1 U10503 ( .A(n9445), .B(n9444), .ZN(n10244) );
  INV_X1 U10504 ( .A(n14269), .ZN(n14285) );
  INV_X1 U10505 ( .A(n15247), .ZN(n14742) );
  INV_X1 U10506 ( .A(n15024), .ZN(n14925) );
  OR2_X1 U10507 ( .A1(n6408), .A2(n15296), .ZN(n15026) );
  OR2_X1 U10508 ( .A1(n15033), .A2(n15032), .ZN(n15365) );
  NAND2_X1 U10509 ( .A1(n15063), .A2(n15062), .ZN(n15166) );
  AND3_X1 U10510 ( .A1(n15352), .A2(n15351), .A3(n15350), .ZN(n15366) );
  OR2_X1 U10511 ( .A1(n15033), .A2(n11463), .ZN(n15353) );
  NAND2_X1 U10512 ( .A1(n10813), .A2(n10184), .ZN(n15666) );
  INV_X1 U10513 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n11807) );
  INV_X1 U10514 ( .A(n14483), .ZN(n11494) );
  INV_X1 U10515 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10748) );
  INV_X2 U10516 ( .A(n12571), .ZN(P3_U3897) );
  NOR2_X1 U10517 ( .A1(P2_U3088), .A2(n10299), .ZN(P2_U3947) );
  NAND2_X1 U10518 ( .A1(n7965), .A2(n8696), .ZN(P2_U3236) );
  NAND2_X1 U10519 ( .A1(n7218), .A2(n8006), .ZN(n7978) );
  NAND3_X1 U10520 ( .A1(n8072), .A2(n8000), .A3(n7977), .ZN(n8108) );
  NAND2_X1 U10521 ( .A1(n8005), .A2(n8004), .ZN(n7980) );
  NAND3_X1 U10522 ( .A1(n8003), .A2(n7998), .A3(n8002), .ZN(n7979) );
  INV_X1 U10523 ( .A(n8622), .ZN(n7987) );
  NOR2_X1 U10524 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n7985) );
  INV_X1 U10525 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n7991) );
  INV_X1 U10526 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U10527 ( .A1(n8626), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n7997) );
  NOR2_X1 U10528 ( .A1(n8622), .A2(n7997), .ZN(n8009) );
  XNOR2_X1 U10529 ( .A(n7989), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8008) );
  NAND3_X1 U10530 ( .A1(n8072), .A2(n8000), .A3(n7999), .ZN(n8001) );
  NAND2_X1 U10531 ( .A1(n6539), .A2(n7955), .ZN(n8007) );
  NOR2_X2 U10532 ( .A1(n8007), .A2(n8231), .ZN(n8584) );
  AND2_X1 U10533 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n8013) );
  AND2_X1 U10534 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U10535 ( .A1(n8039), .A2(n8014), .ZN(n8029) );
  INV_X1 U10536 ( .A(SI_1_), .ZN(n10143) );
  XNOR2_X1 U10537 ( .A(n8042), .B(n10143), .ZN(n8016) );
  XNOR2_X1 U10538 ( .A(n8016), .B(n8015), .ZN(n10189) );
  NAND2_X1 U10539 ( .A1(n8055), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8021) );
  NAND2_X1 U10540 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8018) );
  INV_X1 U10541 ( .A(n7218), .ZN(n8047) );
  NAND2_X1 U10542 ( .A1(n8019), .A2(n8047), .ZN(n15379) );
  INV_X1 U10543 ( .A(n15379), .ZN(n10312) );
  NAND2_X1 U10544 ( .A1(n8046), .A2(n10312), .ZN(n8020) );
  OAI211_X2 U10545 ( .C1(n13495), .C2(n10189), .A(n8021), .B(n8020), .ZN(
        n13916) );
  NAND2_X1 U10546 ( .A1(n8596), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8027) );
  INV_X1 U10547 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n8022) );
  OR2_X1 U10548 ( .A1(n8077), .A2(n8022), .ZN(n8026) );
  INV_X1 U10549 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10887) );
  OR2_X1 U10550 ( .A1(n8595), .A2(n10887), .ZN(n8025) );
  INV_X1 U10551 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n8023) );
  OR2_X1 U10552 ( .A1(n8239), .A2(n8023), .ZN(n8024) );
  NAND2_X1 U10553 ( .A1(n7875), .A2(SI_0_), .ZN(n8028) );
  NAND2_X1 U10554 ( .A1(n8028), .A2(n9494), .ZN(n8030) );
  AND2_X1 U10555 ( .A1(n8029), .A2(n8030), .ZN(n14103) );
  MUX2_X1 U10556 ( .A(P2_IR_REG_0__SCAN_IN), .B(n14103), .S(n10296), .Z(n13296) );
  NAND2_X1 U10557 ( .A1(n13293), .A2(n13296), .ZN(n12150) );
  NAND2_X1 U10558 ( .A1(n12148), .A2(n8032), .ZN(n11200) );
  INV_X1 U10559 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10560 ( .A1(n8596), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8037) );
  INV_X1 U10561 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n11208) );
  OR2_X1 U10562 ( .A1(n8595), .A2(n11208), .ZN(n8036) );
  INV_X1 U10563 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n8034) );
  OR2_X1 U10564 ( .A1(n8239), .A2(n8034), .ZN(n8035) );
  INV_X1 U10566 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n10188) );
  AOI21_X1 U10567 ( .B1(n8039), .B2(P1_DATAO_REG_1__SCAN_IN), .A(SI_1_), .ZN(
        n8040) );
  OAI21_X1 U10568 ( .B1(n8039), .B2(n10188), .A(n8040), .ZN(n8041) );
  NAND2_X1 U10569 ( .A1(n8039), .A2(n10153), .ZN(n8043) );
  OAI211_X1 U10570 ( .C1(P2_DATAO_REG_1__SCAN_IN), .C2(n6413), .A(n8043), .B(
        SI_1_), .ZN(n8044) );
  XNOR2_X1 U10571 ( .A(n8054), .B(n8053), .ZN(n10165) );
  INV_X1 U10572 ( .A(n10350), .ZN(n10314) );
  NAND2_X1 U10573 ( .A1(n8055), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U10574 ( .A1(n11200), .A2(n13540), .ZN(n11199) );
  INV_X1 U10575 ( .A(SI_2_), .ZN(n10150) );
  NAND2_X1 U10576 ( .A1(n8048), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8056) );
  MUX2_X1 U10577 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8056), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8057) );
  AOI22_X1 U10578 ( .A1(n8055), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n8046), .B2(
        n10317), .ZN(n8058) );
  NAND2_X1 U10579 ( .A1(n8596), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8064) );
  INV_X1 U10580 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n8059) );
  OR2_X1 U10581 ( .A1(n8077), .A2(n8059), .ZN(n8063) );
  OR2_X1 U10582 ( .A1(n8595), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8062) );
  INV_X1 U10583 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n8060) );
  OR2_X1 U10584 ( .A1(n8239), .A2(n8060), .ZN(n8061) );
  NAND2_X1 U10585 ( .A1(n7395), .A2(n13286), .ZN(n8065) );
  NAND2_X1 U10586 ( .A1(n8068), .A2(SI_3_), .ZN(n8069) );
  XNOR2_X1 U10587 ( .A(n8086), .B(n8084), .ZN(n10160) );
  INV_X2 U10588 ( .A(n13495), .ZN(n8146) );
  NAND2_X1 U10589 ( .A1(n10160), .A2(n8146), .ZN(n8076) );
  NAND2_X1 U10590 ( .A1(n8071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8070) );
  MUX2_X1 U10591 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8070), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n8074) );
  INV_X1 U10592 ( .A(n8071), .ZN(n8073) );
  NAND2_X1 U10593 ( .A1(n8073), .A2(n8072), .ZN(n8089) );
  NAND2_X1 U10594 ( .A1(n8074), .A2(n8089), .ZN(n15403) );
  INV_X1 U10595 ( .A(n15403), .ZN(n10320) );
  AOI22_X1 U10596 ( .A1(n8055), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n8046), .B2(
        n10320), .ZN(n8075) );
  NAND2_X1 U10597 ( .A1(n8596), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n8083) );
  INV_X1 U10598 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n8078) );
  OAI21_X1 U10599 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n8095), .ZN(n13184) );
  OR2_X1 U10600 ( .A1(n8595), .A2(n13184), .ZN(n8081) );
  INV_X1 U10601 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n8079) );
  OR2_X1 U10602 ( .A1(n8239), .A2(n8079), .ZN(n8080) );
  XNOR2_X1 U10603 ( .A(n13320), .B(n13608), .ZN(n13543) );
  INV_X1 U10604 ( .A(n13608), .ZN(n11183) );
  NAND2_X1 U10605 ( .A1(n13320), .A2(n11183), .ZN(n11185) );
  NAND2_X1 U10606 ( .A1(n8087), .A2(SI_4_), .ZN(n8088) );
  XNOR2_X1 U10607 ( .A(n8103), .B(n8105), .ZN(n10176) );
  NAND2_X1 U10608 ( .A1(n10176), .A2(n8146), .ZN(n8092) );
  NAND2_X1 U10609 ( .A1(n8089), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8090) );
  XNOR2_X1 U10610 ( .A(n8090), .B(P2_IR_REG_5__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U10611 ( .A1(n8055), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n8046), .B2(
        n10362), .ZN(n8091) );
  NAND2_X1 U10612 ( .A1(n8092), .A2(n8091), .ZN(n13328) );
  NAND2_X1 U10613 ( .A1(n8597), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n8100) );
  INV_X1 U10614 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n10311) );
  OR2_X1 U10615 ( .A1(n8398), .A2(n10311), .ZN(n8099) );
  INV_X1 U10616 ( .A(n8095), .ZN(n8093) );
  INV_X1 U10617 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10618 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  NAND2_X1 U10619 ( .A1(n8114), .A2(n8096), .ZN(n11194) );
  OR2_X1 U10620 ( .A1(n8595), .A2(n11194), .ZN(n8098) );
  INV_X1 U10621 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10301) );
  OR2_X1 U10622 ( .A1(n8239), .A2(n10301), .ZN(n8097) );
  NAND2_X1 U10623 ( .A1(n13328), .A2(n13330), .ZN(n8102) );
  OR2_X1 U10624 ( .A1(n13328), .A2(n13330), .ZN(n8101) );
  INV_X1 U10625 ( .A(n8103), .ZN(n8104) );
  NAND2_X1 U10626 ( .A1(n8106), .A2(SI_5_), .ZN(n8107) );
  XNOR2_X1 U10627 ( .A(n8123), .B(SI_6_), .ZN(n8120) );
  NAND2_X1 U10628 ( .A1(n10180), .A2(n8146), .ZN(n8111) );
  NOR2_X1 U10629 ( .A1(n8048), .A2(n8108), .ZN(n8233) );
  INV_X1 U10630 ( .A(n8233), .ZN(n8587) );
  NAND2_X1 U10631 ( .A1(n8587), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8109) );
  XNOR2_X1 U10632 ( .A(n8109), .B(P2_IR_REG_6__SCAN_IN), .ZN(n13615) );
  AOI22_X1 U10633 ( .A1(n13496), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n8046), 
        .B2(n13615), .ZN(n8110) );
  INV_X1 U10634 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10353) );
  OR2_X1 U10635 ( .A1(n8398), .A2(n10353), .ZN(n8118) );
  INV_X1 U10636 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10637 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  NAND2_X1 U10638 ( .A1(n8131), .A2(n8115), .ZN(n11322) );
  OR2_X1 U10639 ( .A1(n8595), .A2(n11322), .ZN(n8117) );
  INV_X1 U10640 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10365) );
  OR2_X1 U10641 ( .A1(n8239), .A2(n10365), .ZN(n8116) );
  XNOR2_X1 U10642 ( .A(n14036), .B(n13606), .ZN(n13546) );
  INV_X1 U10643 ( .A(n13606), .ZN(n11182) );
  NAND2_X1 U10644 ( .A1(n14036), .A2(n11182), .ZN(n8119) );
  INV_X1 U10645 ( .A(n8120), .ZN(n8121) );
  NAND2_X1 U10646 ( .A1(n8123), .A2(SI_6_), .ZN(n8124) );
  XNOR2_X1 U10647 ( .A(n8144), .B(SI_7_), .ZN(n8141) );
  XNOR2_X1 U10648 ( .A(n8143), .B(n8141), .ZN(n10194) );
  NAND2_X1 U10649 ( .A1(n10194), .A2(n8146), .ZN(n8129) );
  INV_X1 U10650 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8126) );
  NAND2_X1 U10651 ( .A1(n8233), .A2(n8126), .ZN(n8147) );
  NAND2_X1 U10652 ( .A1(n8147), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8127) );
  XNOR2_X1 U10653 ( .A(n8127), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13628) );
  AOI22_X1 U10654 ( .A1(n8046), .A2(n13628), .B1(n13496), .B2(
        P1_DATAO_REG_7__SCAN_IN), .ZN(n8128) );
  NAND2_X1 U10655 ( .A1(n8597), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n8137) );
  INV_X1 U10656 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n11175) );
  OR2_X1 U10657 ( .A1(n8398), .A2(n11175), .ZN(n8136) );
  INV_X1 U10658 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U10659 ( .A1(n8131), .A2(n11125), .ZN(n8132) );
  NAND2_X1 U10660 ( .A1(n8156), .A2(n8132), .ZN(n11174) );
  OR2_X1 U10661 ( .A1(n8595), .A2(n11174), .ZN(n8135) );
  INV_X1 U10662 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8133) );
  OR2_X1 U10663 ( .A1(n8239), .A2(n8133), .ZN(n8134) );
  OR2_X1 U10664 ( .A1(n15525), .A2(n13343), .ZN(n8138) );
  NAND2_X1 U10665 ( .A1(n15525), .A2(n13343), .ZN(n8139) );
  INV_X1 U10666 ( .A(n8141), .ZN(n8142) );
  NAND2_X1 U10667 ( .A1(n8144), .A2(SI_7_), .ZN(n8145) );
  XNOR2_X1 U10668 ( .A(n8167), .B(SI_8_), .ZN(n8164) );
  XNOR2_X1 U10669 ( .A(n8166), .B(n8164), .ZN(n10234) );
  NAND2_X1 U10670 ( .A1(n10234), .A2(n8146), .ZN(n8152) );
  NAND2_X1 U10671 ( .A1(n8149), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8148) );
  MUX2_X1 U10672 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8148), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n8150) );
  AOI22_X1 U10673 ( .A1(n10369), .A2(n8046), .B1(n13496), .B2(
        P1_DATAO_REG_8__SCAN_IN), .ZN(n8151) );
  NAND2_X1 U10674 ( .A1(n8596), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n8161) );
  INV_X1 U10675 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n8153) );
  OR2_X1 U10676 ( .A1(n8077), .A2(n8153), .ZN(n8160) );
  INV_X1 U10677 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n8155) );
  NAND2_X1 U10678 ( .A1(n8156), .A2(n8155), .ZN(n8157) );
  NAND2_X1 U10679 ( .A1(n8180), .A2(n8157), .ZN(n12192) );
  OR2_X1 U10680 ( .A1(n8595), .A2(n12192), .ZN(n8159) );
  INV_X1 U10681 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10368) );
  OR2_X1 U10682 ( .A1(n8239), .A2(n10368), .ZN(n8158) );
  AND2_X1 U10683 ( .A1(n14031), .A2(n13345), .ZN(n8163) );
  OR2_X1 U10684 ( .A1(n14031), .A2(n13345), .ZN(n8162) );
  INV_X1 U10685 ( .A(n8164), .ZN(n8165) );
  NAND2_X1 U10686 ( .A1(n8167), .A2(SI_8_), .ZN(n8168) );
  XNOR2_X1 U10687 ( .A(n8191), .B(SI_9_), .ZN(n8188) );
  NAND2_X1 U10688 ( .A1(n10239), .A2(n8146), .ZN(n8177) );
  NAND2_X1 U10689 ( .A1(n8170), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8169) );
  MUX2_X1 U10690 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8169), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n8173) );
  INV_X1 U10691 ( .A(n8170), .ZN(n8172) );
  INV_X1 U10692 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8171) );
  NAND2_X1 U10693 ( .A1(n8172), .A2(n8171), .ZN(n8212) );
  NAND2_X1 U10694 ( .A1(n8173), .A2(n8212), .ZN(n10944) );
  OAI22_X1 U10695 ( .A1(n10944), .A2(n10296), .B1(n8174), .B2(n10240), .ZN(
        n8175) );
  INV_X1 U10696 ( .A(n8175), .ZN(n8176) );
  INV_X1 U10697 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n11612) );
  OR2_X1 U10698 ( .A1(n8398), .A2(n11612), .ZN(n8186) );
  INV_X1 U10699 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n15718) );
  OR2_X1 U10700 ( .A1(n8077), .A2(n15718), .ZN(n8185) );
  INV_X1 U10701 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n8179) );
  NAND2_X1 U10702 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  NAND2_X1 U10703 ( .A1(n8199), .A2(n8181), .ZN(n12162) );
  OR2_X1 U10704 ( .A1(n8595), .A2(n12162), .ZN(n8184) );
  INV_X1 U10705 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n8182) );
  OR2_X1 U10706 ( .A1(n8239), .A2(n8182), .ZN(n8183) );
  NAND4_X1 U10707 ( .A1(n8186), .A2(n8185), .A3(n8184), .A4(n8183), .ZN(n13603) );
  OR2_X1 U10708 ( .A1(n13352), .A2(n13603), .ZN(n8659) );
  NAND2_X1 U10709 ( .A1(n13352), .A2(n13603), .ZN(n11712) );
  NAND2_X1 U10710 ( .A1(n8659), .A2(n11712), .ZN(n13549) );
  INV_X1 U10711 ( .A(n13603), .ZN(n8187) );
  INV_X1 U10712 ( .A(n8188), .ZN(n8189) );
  NAND2_X1 U10713 ( .A1(n8191), .A2(SI_9_), .ZN(n8192) );
  NAND2_X1 U10714 ( .A1(n10284), .A2(n8146), .ZN(n8196) );
  NAND2_X1 U10715 ( .A1(n8212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8194) );
  AOI22_X1 U10716 ( .A1(n15428), .A2(n8046), .B1(n13496), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n8195) );
  NAND2_X1 U10717 ( .A1(n8597), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n8204) );
  INV_X1 U10718 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8197) );
  OR2_X1 U10719 ( .A1(n8239), .A2(n8197), .ZN(n8203) );
  OR2_X2 U10720 ( .A1(n8199), .A2(n8198), .ZN(n8218) );
  NAND2_X1 U10721 ( .A1(n8199), .A2(n8198), .ZN(n8200) );
  NAND2_X1 U10722 ( .A1(n8218), .A2(n8200), .ZN(n11720) );
  OR2_X1 U10723 ( .A1(n8595), .A2(n11720), .ZN(n8202) );
  INV_X1 U10724 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10947) );
  OR2_X1 U10725 ( .A1(n8398), .A2(n10947), .ZN(n8201) );
  OR2_X1 U10726 ( .A1(n14026), .A2(n13358), .ZN(n11710) );
  NAND2_X1 U10727 ( .A1(n14026), .A2(n13358), .ZN(n11709) );
  NAND2_X1 U10728 ( .A1(n8208), .A2(SI_10_), .ZN(n8249) );
  MUX2_X1 U10729 ( .A(n10464), .B(n10458), .S(n6413), .Z(n8210) );
  NAND2_X1 U10730 ( .A1(n8210), .A2(n10201), .ZN(n8254) );
  INV_X1 U10731 ( .A(n8210), .ZN(n8211) );
  NAND2_X1 U10732 ( .A1(n8211), .A2(SI_11_), .ZN(n8248) );
  NAND2_X1 U10733 ( .A1(n8254), .A2(n8248), .ZN(n8226) );
  NAND2_X1 U10734 ( .A1(n10457), .A2(n8146), .ZN(n8215) );
  OAI21_X1 U10735 ( .B1(n8212), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8213) );
  XNOR2_X1 U10736 ( .A(n8213), .B(P2_IR_REG_11__SCAN_IN), .ZN(n11751) );
  AOI22_X1 U10737 ( .A1(n11751), .A2(n8046), .B1(n13496), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U10738 ( .A1(n8597), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n8224) );
  INV_X1 U10739 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11735) );
  OR2_X1 U10740 ( .A1(n8398), .A2(n11735), .ZN(n8223) );
  INV_X1 U10741 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n8217) );
  NAND2_X1 U10742 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  NAND2_X1 U10743 ( .A1(n8242), .A2(n8219), .ZN(n12175) );
  OR2_X1 U10744 ( .A1(n8595), .A2(n12175), .ZN(n8222) );
  INV_X1 U10745 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8220) );
  OR2_X1 U10746 ( .A1(n8239), .A2(n8220), .ZN(n8221) );
  NAND4_X1 U10747 ( .A1(n8224), .A2(n8223), .A3(n8222), .A4(n8221), .ZN(n13601) );
  INV_X1 U10748 ( .A(n13601), .ZN(n13367) );
  NAND2_X1 U10749 ( .A1(n13365), .A2(n13367), .ZN(n8225) );
  MUX2_X1 U10750 ( .A(n15769), .B(n10500), .S(n6413), .Z(n8228) );
  NAND2_X1 U10751 ( .A1(n8228), .A2(n10233), .ZN(n8255) );
  INV_X1 U10752 ( .A(n8228), .ZN(n8229) );
  NAND2_X1 U10753 ( .A1(n8229), .A2(SI_12_), .ZN(n8230) );
  NAND2_X1 U10754 ( .A1(n8255), .A2(n8230), .ZN(n8251) );
  INV_X1 U10755 ( .A(n8251), .ZN(n8258) );
  NAND2_X1 U10756 ( .A1(n10498), .A2(n8146), .ZN(n8238) );
  INV_X1 U10757 ( .A(n8231), .ZN(n8232) );
  NAND2_X1 U10758 ( .A1(n8233), .A2(n8232), .ZN(n8235) );
  NAND2_X1 U10759 ( .A1(n8235), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8234) );
  MUX2_X1 U10760 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8234), .S(
        P2_IR_REG_12__SCAN_IN), .Z(n8236) );
  AOI22_X1 U10761 ( .A1(n13496), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n8046), 
        .B2(n11754), .ZN(n8237) );
  INV_X1 U10762 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15765) );
  OR2_X1 U10763 ( .A1(n8077), .A2(n15765), .ZN(n8241) );
  INV_X1 U10764 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n15667) );
  OR2_X1 U10765 ( .A1(n8239), .A2(n15667), .ZN(n8240) );
  AND2_X1 U10766 ( .A1(n8241), .A2(n8240), .ZN(n8246) );
  NAND2_X1 U10767 ( .A1(n8242), .A2(n12078), .ZN(n8243) );
  AND2_X1 U10768 ( .A1(n8267), .A2(n8243), .ZN(n12083) );
  NAND2_X1 U10769 ( .A1(n12083), .A2(n8519), .ZN(n8245) );
  INV_X1 U10770 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11755) );
  OR2_X1 U10771 ( .A1(n8398), .A2(n11755), .ZN(n8244) );
  XNOR2_X1 U10772 ( .A(n14085), .B(n13372), .ZN(n13553) );
  OR2_X1 U10773 ( .A1(n14085), .A2(n13372), .ZN(n8247) );
  NAND2_X1 U10774 ( .A1(n8249), .A2(n8248), .ZN(n8250) );
  NOR2_X1 U10775 ( .A1(n8251), .A2(n8250), .ZN(n8252) );
  INV_X1 U10776 ( .A(n8254), .ZN(n8257) );
  INV_X1 U10777 ( .A(n8255), .ZN(n8256) );
  AOI21_X1 U10778 ( .B1(n8258), .B2(n8257), .A(n8256), .ZN(n8259) );
  MUX2_X1 U10779 ( .A(n9751), .B(n10494), .S(n7875), .Z(n8260) );
  INV_X1 U10780 ( .A(n8260), .ZN(n8261) );
  NAND2_X1 U10781 ( .A1(n8261), .A2(SI_13_), .ZN(n8262) );
  XNOR2_X1 U10782 ( .A(n8275), .B(n7959), .ZN(n10455) );
  NAND2_X1 U10783 ( .A1(n10455), .A2(n8146), .ZN(n8266) );
  NAND2_X1 U10784 ( .A1(n8263), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8264) );
  XNOR2_X1 U10785 ( .A(n8264), .B(P2_IR_REG_13__SCAN_IN), .ZN(n15456) );
  AOI22_X1 U10786 ( .A1(n13496), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n8046), 
        .B2(n15456), .ZN(n8265) );
  NAND2_X2 U10787 ( .A1(n8266), .A2(n8265), .ZN(n14014) );
  INV_X1 U10788 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n15668) );
  NAND2_X1 U10789 ( .A1(n8267), .A2(n15668), .ZN(n8268) );
  NAND2_X1 U10790 ( .A1(n8283), .A2(n8268), .ZN(n13901) );
  OR2_X1 U10791 ( .A1(n13901), .A2(n8595), .ZN(n8271) );
  AOI22_X1 U10792 ( .A1(n8304), .A2(P2_REG1_REG_13__SCAN_IN), .B1(n8597), .B2(
        P2_REG0_REG_13__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10793 ( .A1(n8596), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n8269) );
  NAND2_X1 U10794 ( .A1(n14014), .A2(n13552), .ZN(n8272) );
  OR2_X1 U10795 ( .A1(n14014), .A2(n13552), .ZN(n8273) );
  NAND2_X1 U10796 ( .A1(n8312), .A2(n10497), .ZN(n8289) );
  MUX2_X1 U10797 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n7875), .Z(n8308) );
  NAND2_X1 U10798 ( .A1(n10763), .A2(n8146), .ZN(n8281) );
  NAND2_X1 U10799 ( .A1(n8278), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8279) );
  XNOR2_X1 U10800 ( .A(n8279), .B(P2_IR_REG_14__SCAN_IN), .ZN(n13649) );
  AOI22_X1 U10801 ( .A1(n13496), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n8046), 
        .B2(n13649), .ZN(n8280) );
  OR2_X2 U10802 ( .A1(n8283), .A2(n8282), .ZN(n8302) );
  NAND2_X1 U10803 ( .A1(n8283), .A2(n8282), .ZN(n8284) );
  NAND2_X1 U10804 ( .A1(n8302), .A2(n8284), .ZN(n13886) );
  OR2_X1 U10805 ( .A1(n13886), .A2(n8595), .ZN(n8287) );
  AOI22_X1 U10806 ( .A1(n8596), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8597), .B2(
        P2_REG0_REG_14__SCAN_IN), .ZN(n8286) );
  NAND2_X1 U10807 ( .A1(n8304), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n8285) );
  NAND2_X1 U10808 ( .A1(n14009), .A2(n13386), .ZN(n8288) );
  MUX2_X1 U10809 ( .A(n10831), .B(n10830), .S(n7875), .Z(n8291) );
  NAND2_X1 U10810 ( .A1(n8291), .A2(n10637), .ZN(n8313) );
  INV_X1 U10811 ( .A(n8291), .ZN(n8292) );
  NAND2_X1 U10812 ( .A1(n8292), .A2(SI_15_), .ZN(n8293) );
  NAND2_X1 U10813 ( .A1(n8313), .A2(n8293), .ZN(n8311) );
  INV_X1 U10814 ( .A(n8311), .ZN(n8294) );
  NAND2_X1 U10815 ( .A1(n10829), .A2(n8146), .ZN(n8300) );
  INV_X1 U10816 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8296) );
  NAND2_X1 U10817 ( .A1(n8297), .A2(n8296), .ZN(n8391) );
  NAND2_X1 U10818 ( .A1(n8391), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8298) );
  XNOR2_X1 U10819 ( .A(n8298), .B(P2_IR_REG_15__SCAN_IN), .ZN(n13652) );
  AOI22_X1 U10820 ( .A1(n13496), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n8046), 
        .B2(n13652), .ZN(n8299) );
  INV_X1 U10821 ( .A(n8325), .ZN(n8327) );
  NAND2_X1 U10822 ( .A1(n8302), .A2(n8301), .ZN(n8303) );
  AND2_X1 U10823 ( .A1(n8327), .A2(n8303), .ZN(n13872) );
  NAND2_X1 U10824 ( .A1(n13872), .A2(n8519), .ZN(n8307) );
  AOI22_X1 U10825 ( .A1(n8596), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8597), .B2(
        P2_REG0_REG_15__SCAN_IN), .ZN(n8306) );
  NAND2_X1 U10826 ( .A1(n8304), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8305) );
  AND2_X1 U10827 ( .A1(n13866), .A2(n13392), .ZN(n13809) );
  INV_X1 U10828 ( .A(n8308), .ZN(n8309) );
  NOR2_X1 U10829 ( .A1(n8309), .A2(n10497), .ZN(n8310) );
  MUX2_X1 U10830 ( .A(n10748), .B(n10751), .S(n7875), .Z(n8315) );
  INV_X1 U10831 ( .A(n8315), .ZN(n8316) );
  NAND2_X1 U10832 ( .A1(n8316), .A2(SI_16_), .ZN(n8317) );
  XNOR2_X1 U10833 ( .A(n8337), .B(n8336), .ZN(n10747) );
  NAND2_X1 U10834 ( .A1(n10747), .A2(n8146), .ZN(n8324) );
  OR2_X1 U10835 ( .A1(n8391), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U10836 ( .A1(n8319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8318) );
  MUX2_X1 U10837 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8318), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n8322) );
  INV_X1 U10838 ( .A(n8319), .ZN(n8321) );
  INV_X1 U10839 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10840 ( .A1(n8321), .A2(n8320), .ZN(n8361) );
  NAND2_X1 U10841 ( .A1(n8322), .A2(n8361), .ZN(n13643) );
  AOI22_X1 U10842 ( .A1(n8046), .A2(n15482), .B1(n13496), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n8323) );
  INV_X1 U10843 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8326) );
  NAND2_X1 U10844 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  NAND2_X1 U10845 ( .A1(n8366), .A2(n8328), .ZN(n13854) );
  OR2_X1 U10846 ( .A1(n13854), .A2(n8595), .ZN(n8334) );
  INV_X1 U10847 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U10848 ( .A1(n8597), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10849 ( .A1(n8596), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8329) );
  OAI211_X1 U10850 ( .C1(n8331), .C2(n8239), .A(n8330), .B(n8329), .ZN(n8332)
         );
  INV_X1 U10851 ( .A(n8332), .ZN(n8333) );
  OR2_X1 U10852 ( .A1(n13996), .A2(n13397), .ZN(n13811) );
  OAI21_X1 U10853 ( .B1(n13866), .B2(n13392), .A(n13811), .ZN(n8335) );
  MUX2_X1 U10854 ( .A(n10896), .B(n10900), .S(n7875), .Z(n8339) );
  INV_X1 U10855 ( .A(n8339), .ZN(n8338) );
  NAND2_X1 U10856 ( .A1(n8360), .A2(n11103), .ZN(n8345) );
  INV_X1 U10857 ( .A(n8381), .ZN(n8340) );
  NAND2_X1 U10858 ( .A1(n8340), .A2(n11103), .ZN(n8343) );
  INV_X1 U10859 ( .A(n8360), .ZN(n8341) );
  NAND2_X1 U10860 ( .A1(n8341), .A2(SI_18_), .ZN(n8342) );
  OAI211_X1 U10861 ( .C1(n8345), .C2(n8358), .A(n8343), .B(n8342), .ZN(n8344)
         );
  MUX2_X1 U10862 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n7875), .Z(n8409) );
  XNOR2_X1 U10863 ( .A(n8382), .B(n8409), .ZN(n10924) );
  NAND2_X1 U10864 ( .A1(n10924), .A2(n8146), .ZN(n8348) );
  OAI21_X1 U10865 ( .B1(n8361), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8346) );
  XNOR2_X1 U10866 ( .A(n8346), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13663) );
  AOI22_X1 U10867 ( .A1(n13663), .A2(n8046), .B1(n13496), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n8347) );
  INV_X1 U10868 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10869 ( .A1(n8368), .A2(n8350), .ZN(n8351) );
  AND2_X1 U10870 ( .A1(n8394), .A2(n8351), .ZN(n13822) );
  NAND2_X1 U10871 ( .A1(n13822), .A2(n8519), .ZN(n8357) );
  INV_X1 U10872 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8354) );
  NAND2_X1 U10873 ( .A1(n8304), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8353) );
  NAND2_X1 U10874 ( .A1(n8597), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n8352) );
  OAI211_X1 U10875 ( .C1(n8398), .C2(n8354), .A(n8353), .B(n8352), .ZN(n8355)
         );
  INV_X1 U10876 ( .A(n8355), .ZN(n8356) );
  NAND2_X1 U10877 ( .A1(n13821), .A2(n13126), .ZN(n8377) );
  XNOR2_X1 U10878 ( .A(n8380), .B(n8379), .ZN(n10895) );
  NAND2_X1 U10879 ( .A1(n10895), .A2(n8146), .ZN(n8364) );
  NAND2_X1 U10880 ( .A1(n8361), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8362) );
  XNOR2_X1 U10881 ( .A(n8362), .B(P2_IR_REG_17__SCAN_IN), .ZN(n15497) );
  AOI22_X1 U10882 ( .A1(n15497), .A2(n8046), .B1(n13496), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n8363) );
  INV_X1 U10883 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8365) );
  NAND2_X1 U10884 ( .A1(n8366), .A2(n8365), .ZN(n8367) );
  NAND2_X1 U10885 ( .A1(n8368), .A2(n8367), .ZN(n13844) );
  OR2_X1 U10886 ( .A1(n13844), .A2(n8595), .ZN(n8374) );
  INV_X1 U10887 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8371) );
  NAND2_X1 U10888 ( .A1(n8597), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n8370) );
  NAND2_X1 U10889 ( .A1(n8596), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8369) );
  OAI211_X1 U10890 ( .C1(n8239), .C2(n8371), .A(n8370), .B(n8369), .ZN(n8372)
         );
  INV_X1 U10891 ( .A(n8372), .ZN(n8373) );
  NAND2_X1 U10892 ( .A1(n14073), .A2(n13409), .ZN(n8670) );
  INV_X1 U10893 ( .A(n8670), .ZN(n8375) );
  NOR2_X1 U10894 ( .A1(n14073), .A2(n13409), .ZN(n13812) );
  INV_X1 U10895 ( .A(n13821), .ZN(n14070) );
  AOI22_X1 U10896 ( .A1(n8377), .A2(n13812), .B1(n14070), .B2(n13596), .ZN(
        n8378) );
  INV_X1 U10897 ( .A(n8409), .ZN(n8405) );
  MUX2_X1 U10898 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n7875), .Z(n8383) );
  NAND2_X1 U10899 ( .A1(n8383), .A2(SI_19_), .ZN(n8412) );
  INV_X1 U10900 ( .A(n8383), .ZN(n8384) );
  INV_X1 U10901 ( .A(SI_19_), .ZN(n11164) );
  NAND2_X1 U10902 ( .A1(n8384), .A2(n11164), .ZN(n8410) );
  NAND2_X1 U10903 ( .A1(n8412), .A2(n8410), .ZN(n8385) );
  INV_X1 U10904 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8388) );
  INV_X1 U10905 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n8387) );
  NAND3_X1 U10906 ( .A1(n8389), .A2(n8388), .A3(n8387), .ZN(n8390) );
  OAI21_X1 U10907 ( .B1(n8391), .B2(n8390), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8392) );
  AOI22_X1 U10908 ( .A1(n13496), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n13672), 
        .B2(n8046), .ZN(n8393) );
  INV_X1 U10909 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n15722) );
  NAND2_X1 U10910 ( .A1(n8394), .A2(n15722), .ZN(n8395) );
  NAND2_X1 U10911 ( .A1(n8431), .A2(n8395), .ZN(n13128) );
  OR2_X1 U10912 ( .A1(n13128), .A2(n8595), .ZN(n8401) );
  INV_X1 U10913 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n13667) );
  NAND2_X1 U10914 ( .A1(n8304), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10915 ( .A1(n8597), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n8396) );
  OAI211_X1 U10916 ( .C1(n8398), .C2(n13667), .A(n8397), .B(n8396), .ZN(n8399)
         );
  INV_X1 U10917 ( .A(n8399), .ZN(n8400) );
  NAND2_X1 U10918 ( .A1(n14065), .A2(n13203), .ZN(n8404) );
  OR2_X1 U10919 ( .A1(n14065), .A2(n13203), .ZN(n8402) );
  OAI21_X1 U10920 ( .B1(n11103), .B2(n8405), .A(n8412), .ZN(n8406) );
  INV_X1 U10921 ( .A(n8406), .ZN(n8407) );
  NOR2_X1 U10922 ( .A1(n8409), .A2(SI_18_), .ZN(n8413) );
  INV_X1 U10923 ( .A(n8410), .ZN(n8411) );
  INV_X1 U10924 ( .A(SI_20_), .ZN(n11335) );
  NAND2_X1 U10925 ( .A1(n8469), .A2(n11335), .ZN(n8425) );
  MUX2_X1 U10926 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(P1_DATAO_REG_20__SCAN_IN), 
        .S(n7875), .Z(n8441) );
  NAND2_X1 U10927 ( .A1(n11454), .A2(n8146), .ZN(n8418) );
  NAND2_X1 U10928 ( .A1(n13496), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8417) );
  XNOR2_X1 U10929 ( .A(n8431), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n13788) );
  NAND2_X1 U10930 ( .A1(n13788), .A2(n8519), .ZN(n8423) );
  INV_X1 U10931 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n15804) );
  NAND2_X1 U10932 ( .A1(n8596), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n8420) );
  NAND2_X1 U10933 ( .A1(n8304), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n8419) );
  OAI211_X1 U10934 ( .C1(n8077), .C2(n15804), .A(n8420), .B(n8419), .ZN(n8421)
         );
  INV_X1 U10935 ( .A(n8421), .ZN(n8422) );
  NAND2_X1 U10936 ( .A1(n8423), .A2(n8422), .ZN(n13595) );
  XNOR2_X1 U10937 ( .A(n13972), .B(n13595), .ZN(n13781) );
  INV_X1 U10938 ( .A(n13595), .ZN(n13421) );
  NAND2_X1 U10939 ( .A1(n13972), .A2(n13421), .ZN(n8424) );
  OAI21_X1 U10940 ( .B1(n8426), .B2(n8441), .A(n8425), .ZN(n8427) );
  MUX2_X1 U10941 ( .A(n11495), .B(n11509), .S(n7875), .Z(n8445) );
  XNOR2_X1 U10942 ( .A(n8445), .B(SI_21_), .ZN(n8440) );
  NAND2_X1 U10943 ( .A1(n11493), .A2(n8146), .ZN(n8429) );
  NAND2_X1 U10944 ( .A1(n13496), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8428) );
  INV_X1 U10945 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n13196) );
  INV_X1 U10946 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13157) );
  OAI21_X1 U10947 ( .B1(n8431), .B2(n13196), .A(n13157), .ZN(n8432) );
  NAND2_X1 U10948 ( .A1(P2_REG3_REG_20__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n8430) );
  AND2_X1 U10949 ( .A1(n8432), .A2(n8453), .ZN(n13772) );
  NAND2_X1 U10950 ( .A1(n13772), .A2(n8519), .ZN(n8437) );
  INV_X1 U10951 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n15733) );
  NAND2_X1 U10952 ( .A1(n8596), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n8434) );
  NAND2_X1 U10953 ( .A1(n8304), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n8433) );
  OAI211_X1 U10954 ( .C1(n8077), .C2(n15733), .A(n8434), .B(n8433), .ZN(n8435)
         );
  INV_X1 U10955 ( .A(n8435), .ZN(n8436) );
  OR2_X1 U10956 ( .A1(n13432), .A2(n13430), .ZN(n8438) );
  NAND2_X1 U10957 ( .A1(n13432), .A2(n13430), .ZN(n8439) );
  NAND2_X1 U10958 ( .A1(n8441), .A2(SI_20_), .ZN(n8464) );
  NAND2_X1 U10959 ( .A1(n8469), .A2(n8464), .ZN(n8444) );
  INV_X1 U10960 ( .A(n8440), .ZN(n8443) );
  NOR2_X1 U10961 ( .A1(n8441), .A2(SI_20_), .ZN(n8442) );
  NAND2_X1 U10962 ( .A1(n8444), .A2(n8470), .ZN(n8447) );
  INV_X1 U10963 ( .A(n8445), .ZN(n8446) );
  NAND2_X1 U10964 ( .A1(n8446), .A2(SI_21_), .ZN(n8466) );
  NAND2_X1 U10965 ( .A1(n8447), .A2(n8466), .ZN(n8449) );
  INV_X1 U10966 ( .A(SI_22_), .ZN(n8448) );
  MUX2_X1 U10967 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n7875), .Z(n8472) );
  INV_X1 U10968 ( .A(n8472), .ZN(n8450) );
  XNOR2_X1 U10969 ( .A(n9289), .B(n8450), .ZN(n11949) );
  NAND2_X1 U10970 ( .A1(n11949), .A2(n8146), .ZN(n8452) );
  NAND2_X1 U10971 ( .A1(n13496), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n8451) );
  INV_X1 U10972 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n13221) );
  NAND2_X1 U10973 ( .A1(n8453), .A2(n13221), .ZN(n8454) );
  NAND2_X1 U10974 ( .A1(n8480), .A2(n8454), .ZN(n12057) );
  OR2_X1 U10975 ( .A1(n12057), .A2(n8595), .ZN(n8460) );
  INV_X1 U10976 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8457) );
  NAND2_X1 U10977 ( .A1(n8597), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n8456) );
  NAND2_X1 U10978 ( .A1(n8596), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n8455) );
  OAI211_X1 U10979 ( .C1(n8239), .C2(n8457), .A(n8456), .B(n8455), .ZN(n8458)
         );
  INV_X1 U10980 ( .A(n8458), .ZN(n8459) );
  NAND2_X1 U10981 ( .A1(n14058), .A2(n13426), .ZN(n8461) );
  NAND2_X1 U10982 ( .A1(n8463), .A2(n8461), .ZN(n13558) );
  INV_X1 U10983 ( .A(n13558), .ZN(n8462) );
  NAND2_X1 U10984 ( .A1(n12052), .A2(n8463), .ZN(n13749) );
  INV_X1 U10985 ( .A(n8464), .ZN(n8467) );
  NAND2_X1 U10986 ( .A1(n8472), .A2(SI_22_), .ZN(n8465) );
  NAND2_X1 U10987 ( .A1(n8466), .A2(n8465), .ZN(n8471) );
  NOR2_X1 U10988 ( .A1(n8467), .A2(n8471), .ZN(n8468) );
  INV_X1 U10989 ( .A(n8470), .ZN(n8475) );
  INV_X1 U10990 ( .A(n8471), .ZN(n8474) );
  NOR2_X1 U10991 ( .A1(n8472), .A2(SI_22_), .ZN(n8473) );
  MUX2_X1 U10992 ( .A(n9897), .B(n9896), .S(n7875), .Z(n8508) );
  XNOR2_X1 U10993 ( .A(n8490), .B(SI_23_), .ZN(n11448) );
  NAND2_X1 U10994 ( .A1(n11448), .A2(n8146), .ZN(n8479) );
  NAND2_X1 U10995 ( .A1(n13496), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n8478) );
  INV_X1 U10996 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n13117) );
  NAND2_X1 U10997 ( .A1(n8480), .A2(n13117), .ZN(n8481) );
  AND2_X1 U10998 ( .A1(n8495), .A2(n8481), .ZN(n13752) );
  NAND2_X1 U10999 ( .A1(n13752), .A2(n8519), .ZN(n8487) );
  INV_X1 U11000 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n8484) );
  NAND2_X1 U11001 ( .A1(n8597), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8483) );
  NAND2_X1 U11002 ( .A1(n8596), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n8482) );
  OAI211_X1 U11003 ( .C1(n8239), .C2(n8484), .A(n8483), .B(n8482), .ZN(n8485)
         );
  INV_X1 U11004 ( .A(n8485), .ZN(n8486) );
  NAND2_X1 U11005 ( .A1(n13956), .A2(n13437), .ZN(n8488) );
  OR2_X1 U11006 ( .A1(n13956), .A2(n13437), .ZN(n8489) );
  OR2_X1 U11007 ( .A1(n8506), .A2(n8508), .ZN(n8491) );
  MUX2_X1 U11008 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n7875), .Z(n8511) );
  XNOR2_X1 U11009 ( .A(n8511), .B(SI_24_), .ZN(n8492) );
  NAND2_X1 U11010 ( .A1(n13496), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8493) );
  INV_X1 U11011 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8494) );
  NAND2_X1 U11012 ( .A1(n8495), .A2(n8494), .ZN(n8496) );
  NAND2_X1 U11013 ( .A1(n8535), .A2(n8496), .ZN(n13741) );
  INV_X1 U11014 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n8499) );
  NAND2_X1 U11015 ( .A1(n8597), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8498) );
  NAND2_X1 U11016 ( .A1(n8596), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n8497) );
  OAI211_X1 U11017 ( .C1(n8499), .C2(n8239), .A(n8498), .B(n8497), .ZN(n8500)
         );
  INV_X1 U11018 ( .A(n8500), .ZN(n8501) );
  INV_X1 U11019 ( .A(n13736), .ZN(n8503) );
  NAND2_X1 U11020 ( .A1(n13948), .A2(n13475), .ZN(n8504) );
  INV_X1 U11021 ( .A(n8508), .ZN(n8510) );
  OAI22_X1 U11022 ( .A1(n8510), .A2(SI_23_), .B1(n8511), .B2(SI_24_), .ZN(
        n8505) );
  INV_X1 U11023 ( .A(SI_23_), .ZN(n11745) );
  INV_X1 U11024 ( .A(SI_24_), .ZN(n8507) );
  OAI21_X1 U11025 ( .B1(n8508), .B2(n11745), .A(n8507), .ZN(n8512) );
  AND2_X1 U11026 ( .A1(SI_24_), .A2(SI_23_), .ZN(n8509) );
  AOI22_X1 U11027 ( .A1(n8512), .A2(n8511), .B1(n8510), .B2(n8509), .ZN(n8513)
         );
  MUX2_X1 U11028 ( .A(n15767), .B(n11492), .S(n7875), .Z(n8514) );
  INV_X1 U11029 ( .A(SI_25_), .ZN(n13094) );
  NAND2_X1 U11030 ( .A1(n8514), .A2(n13094), .ZN(n8528) );
  INV_X1 U11031 ( .A(n8514), .ZN(n8515) );
  NAND2_X1 U11032 ( .A1(n8515), .A2(SI_25_), .ZN(n8516) );
  NAND2_X1 U11033 ( .A1(n8528), .A2(n8516), .ZN(n8526) );
  XNOR2_X1 U11034 ( .A(n8527), .B(n8526), .ZN(n11488) );
  NAND2_X1 U11035 ( .A1(n11488), .A2(n8146), .ZN(n8518) );
  NAND2_X1 U11036 ( .A1(n13496), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8517) );
  XNOR2_X1 U11037 ( .A(n8535), .B(P2_REG3_REG_25__SCAN_IN), .ZN(n13726) );
  NAND2_X1 U11038 ( .A1(n13726), .A2(n8519), .ZN(n8524) );
  INV_X1 U11039 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n13945) );
  NAND2_X1 U11040 ( .A1(n8596), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8521) );
  NAND2_X1 U11041 ( .A1(n8597), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n8520) );
  OAI211_X1 U11042 ( .C1(n13945), .C2(n8239), .A(n8521), .B(n8520), .ZN(n8522)
         );
  INV_X1 U11043 ( .A(n8522), .ZN(n8523) );
  XNOR2_X1 U11044 ( .A(n13722), .B(n13592), .ZN(n13718) );
  INV_X1 U11045 ( .A(n13592), .ZN(n13257) );
  NAND2_X1 U11046 ( .A1(n13722), .A2(n13257), .ZN(n8525) );
  INV_X1 U11047 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n11621) );
  MUX2_X1 U11048 ( .A(n11621), .B(n15780), .S(n7875), .Z(n8543) );
  XNOR2_X1 U11049 ( .A(n8543), .B(SI_26_), .ZN(n8529) );
  XNOR2_X1 U11050 ( .A(n8544), .B(n8529), .ZN(n11620) );
  NAND2_X1 U11051 ( .A1(n11620), .A2(n8146), .ZN(n8531) );
  NAND2_X1 U11052 ( .A1(n13496), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n8530) );
  INV_X1 U11053 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8533) );
  INV_X1 U11054 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8532) );
  OAI21_X1 U11055 ( .B1(n8535), .B2(n8533), .A(n8532), .ZN(n8536) );
  NAND2_X1 U11056 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(P2_REG3_REG_25__SCAN_IN), 
        .ZN(n8534) );
  NAND2_X1 U11057 ( .A1(n8536), .A2(n8548), .ZN(n13260) );
  INV_X1 U11058 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8539) );
  NAND2_X1 U11059 ( .A1(n8596), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U11060 ( .A1(n8597), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8537) );
  OAI211_X1 U11061 ( .C1(n8539), .C2(n8239), .A(n8538), .B(n8537), .ZN(n8540)
         );
  INV_X1 U11062 ( .A(n8540), .ZN(n8541) );
  OR2_X1 U11063 ( .A1(n13940), .A2(n13466), .ZN(n13538) );
  NAND2_X1 U11064 ( .A1(n13940), .A2(n13466), .ZN(n13537) );
  INV_X1 U11065 ( .A(SI_26_), .ZN(n13091) );
  INV_X1 U11066 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12206) );
  MUX2_X1 U11067 ( .A(n11807), .B(n12206), .S(n7875), .Z(n8558) );
  XNOR2_X1 U11068 ( .A(n8558), .B(SI_27_), .ZN(n8545) );
  NAND2_X1 U11069 ( .A1(n11806), .A2(n8146), .ZN(n8547) );
  NAND2_X1 U11070 ( .A1(n13496), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8546) );
  INV_X1 U11071 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n15791) );
  NAND2_X1 U11072 ( .A1(n8548), .A2(n15791), .ZN(n8549) );
  NAND2_X1 U11073 ( .A1(n8570), .A2(n8549), .ZN(n13692) );
  OR2_X1 U11074 ( .A1(n13692), .A2(n8595), .ZN(n8555) );
  INV_X1 U11075 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n8552) );
  NAND2_X1 U11076 ( .A1(n8596), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U11077 ( .A1(n8597), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8550) );
  OAI211_X1 U11078 ( .C1(n8552), .C2(n8239), .A(n8551), .B(n8550), .ZN(n8553)
         );
  INV_X1 U11079 ( .A(n8553), .ZN(n8554) );
  XNOR2_X1 U11080 ( .A(n13933), .B(n13591), .ZN(n13562) );
  NAND2_X1 U11081 ( .A1(n13687), .A2(n13562), .ZN(n8557) );
  INV_X1 U11082 ( .A(n13591), .ZN(n13135) );
  NAND2_X1 U11083 ( .A1(n13933), .A2(n13135), .ZN(n8556) );
  INV_X1 U11084 ( .A(n8558), .ZN(n8561) );
  NOR2_X1 U11085 ( .A1(n8561), .A2(SI_27_), .ZN(n8559) );
  INV_X1 U11086 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n15196) );
  INV_X1 U11087 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9973) );
  MUX2_X1 U11088 ( .A(n15196), .B(n9973), .S(n7875), .Z(n8562) );
  INV_X1 U11089 ( .A(SI_28_), .ZN(n13082) );
  NAND2_X1 U11090 ( .A1(n8562), .A2(n13082), .ZN(n8591) );
  INV_X1 U11091 ( .A(n8562), .ZN(n8563) );
  NAND2_X1 U11092 ( .A1(n8563), .A2(SI_28_), .ZN(n8564) );
  NAND2_X1 U11093 ( .A1(n8591), .A2(n8564), .ZN(n8565) );
  NAND2_X1 U11094 ( .A1(n8566), .A2(n8565), .ZN(n8567) );
  NAND2_X1 U11095 ( .A1(n8592), .A2(n8567), .ZN(n11861) );
  NAND2_X1 U11096 ( .A1(n11861), .A2(n8146), .ZN(n8569) );
  NAND2_X1 U11097 ( .A1(n13496), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8568) );
  INV_X1 U11098 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n13142) );
  OR2_X2 U11099 ( .A1(n8570), .A2(n13142), .ZN(n8689) );
  NAND2_X1 U11100 ( .A1(n8570), .A2(n13142), .ZN(n8571) );
  INV_X1 U11101 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n15711) );
  NAND2_X1 U11102 ( .A1(n8596), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11103 ( .A1(n8597), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n8572) );
  OAI211_X1 U11104 ( .C1(n15711), .C2(n8239), .A(n8573), .B(n8572), .ZN(n8574)
         );
  INV_X1 U11105 ( .A(n8574), .ZN(n8575) );
  NAND2_X2 U11106 ( .A1(n8576), .A2(n8575), .ZN(n13590) );
  NAND2_X1 U11107 ( .A1(n13456), .A2(n13590), .ZN(n8683) );
  OR2_X1 U11108 ( .A1(n13456), .A2(n13590), .ZN(n8577) );
  INV_X1 U11109 ( .A(n13561), .ZN(n8578) );
  NAND2_X1 U11110 ( .A1(n13579), .A2(n13672), .ZN(n13499) );
  NAND2_X1 U11111 ( .A1(n8584), .A2(n8580), .ZN(n8581) );
  NAND2_X1 U11112 ( .A1(n8581), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8582) );
  MUX2_X1 U11113 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8582), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n8583) );
  INV_X1 U11114 ( .A(n8584), .ZN(n8586) );
  XNOR2_X1 U11115 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_20__SCAN_IN), .ZN(
        n8585) );
  OAI21_X1 U11116 ( .B1(n8587), .B2(n8586), .A(n8585), .ZN(n8589) );
  INV_X1 U11117 ( .A(n8588), .ZN(n8623) );
  NAND2_X1 U11118 ( .A1(n13580), .A2(n7902), .ZN(n8590) );
  INV_X1 U11119 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n15190) );
  INV_X1 U11120 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14101) );
  MUX2_X1 U11121 ( .A(n15190), .B(n14101), .S(n7875), .Z(n12030) );
  XNOR2_X1 U11122 ( .A(n12030), .B(SI_29_), .ZN(n12028) );
  NAND2_X1 U11123 ( .A1(n14098), .A2(n8146), .ZN(n8594) );
  NAND2_X1 U11124 ( .A1(n13496), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8593) );
  OR2_X1 U11125 ( .A1(n8689), .A2(n8595), .ZN(n8603) );
  INV_X1 U11126 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n8600) );
  NAND2_X1 U11127 ( .A1(n8596), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n8599) );
  NAND2_X1 U11128 ( .A1(n8597), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8598) );
  OAI211_X1 U11129 ( .C1(n8239), .C2(n8600), .A(n8599), .B(n8598), .ZN(n8601)
         );
  INV_X1 U11130 ( .A(n8601), .ZN(n8602) );
  NAND2_X1 U11131 ( .A1(n8603), .A2(n8602), .ZN(n13589) );
  XNOR2_X1 U11132 ( .A(n13460), .B(n13589), .ZN(n8684) );
  INV_X1 U11133 ( .A(n8684), .ZN(n13565) );
  AOI211_X1 U11134 ( .C1(n6880), .C2(n13590), .A(n13836), .B(n13565), .ZN(
        n8604) );
  NAND3_X1 U11135 ( .A1(n6880), .A2(n13590), .A3(n13897), .ZN(n8610) );
  INV_X1 U11136 ( .A(n10307), .ZN(n8605) );
  INV_X1 U11137 ( .A(n12205), .ZN(n13575) );
  NAND2_X1 U11138 ( .A1(n13575), .A2(P2_B_REG_SCAN_IN), .ZN(n8606) );
  AND2_X1 U11139 ( .A1(n13880), .A2(n8606), .ZN(n13678) );
  INV_X1 U11140 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n13929) );
  NAND2_X1 U11141 ( .A1(n8596), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8608) );
  INV_X1 U11142 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n14045) );
  OR2_X1 U11143 ( .A1(n8077), .A2(n14045), .ZN(n8607) );
  OAI211_X1 U11144 ( .C1(n8239), .C2(n13929), .A(n8608), .B(n8607), .ZN(n13588) );
  AOI22_X1 U11145 ( .A1(n13590), .A2(n13878), .B1(n13678), .B2(n13588), .ZN(
        n8609) );
  OAI21_X1 U11146 ( .B1(n8684), .B2(n8610), .A(n8609), .ZN(n8611) );
  NAND2_X1 U11147 ( .A1(n8614), .A2(n15784), .ZN(n8633) );
  NAND2_X1 U11148 ( .A1(n8616), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8615) );
  MUX2_X1 U11149 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8615), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8619) );
  INV_X1 U11150 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8617) );
  XNOR2_X1 U11151 ( .A(n11563), .B(P2_B_REG_SCAN_IN), .ZN(n8628) );
  NAND2_X1 U11152 ( .A1(n8620), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8621) );
  MUX2_X1 U11153 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8621), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8624) );
  NAND2_X1 U11154 ( .A1(n8625), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8627) );
  INV_X1 U11155 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15505) );
  NAND2_X1 U11156 ( .A1(n15502), .A2(n15505), .ZN(n8630) );
  NAND2_X1 U11157 ( .A1(n11563), .A2(n11624), .ZN(n8629) );
  INV_X1 U11158 ( .A(n11490), .ZN(n8632) );
  NOR2_X1 U11159 ( .A1(n11563), .A2(n11624), .ZN(n8631) );
  NAND2_X1 U11160 ( .A1(n8632), .A2(n8631), .ZN(n10723) );
  NAND2_X1 U11161 ( .A1(n8633), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8635) );
  AND2_X1 U11162 ( .A1(n11449), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8636) );
  NAND2_X1 U11163 ( .A1(n13568), .A2(n13578), .ZN(n13570) );
  NAND2_X1 U11164 ( .A1(n10563), .A2(n13570), .ZN(n10570) );
  INV_X1 U11165 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15510) );
  NAND2_X1 U11166 ( .A1(n15502), .A2(n15510), .ZN(n8638) );
  NAND2_X1 U11167 ( .A1(n11490), .A2(n11624), .ZN(n8637) );
  NOR4_X1 U11168 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n8642) );
  NOR4_X1 U11169 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n8641) );
  NOR4_X1 U11170 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n8640) );
  NOR4_X1 U11171 ( .A1(P2_D_REG_21__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n8639) );
  NAND4_X1 U11172 ( .A1(n8642), .A2(n8641), .A3(n8640), .A4(n8639), .ZN(n8647)
         );
  NOR2_X1 U11173 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n15674) );
  NOR4_X1 U11174 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_3__SCAN_IN), .ZN(n8645) );
  NOR4_X1 U11175 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n8644) );
  NOR4_X1 U11176 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_7__SCAN_IN), .ZN(n8643) );
  NAND4_X1 U11177 ( .A1(n15674), .A2(n8645), .A3(n8644), .A4(n8643), .ZN(n8646) );
  OAI21_X1 U11178 ( .B1(n8647), .B2(n8646), .A(n15502), .ZN(n10562) );
  NAND2_X1 U11179 ( .A1(n10559), .A2(n10562), .ZN(n10569) );
  INV_X1 U11180 ( .A(n10569), .ZN(n8648) );
  NAND4_X1 U11181 ( .A1(n15506), .A2(n15507), .A3(n10570), .A4(n8648), .ZN(
        n8650) );
  INV_X1 U11182 ( .A(n10568), .ZN(n8649) );
  NAND2_X1 U11183 ( .A1(n12151), .A2(n12142), .ZN(n12144) );
  INV_X1 U11184 ( .A(n13304), .ZN(n13610) );
  OR2_X1 U11185 ( .A1(n13609), .A2(n13286), .ZN(n8653) );
  INV_X1 U11186 ( .A(n13543), .ZN(n11002) );
  OR2_X1 U11187 ( .A1(n13320), .A2(n13608), .ZN(n8654) );
  INV_X1 U11188 ( .A(n13330), .ZN(n13607) );
  NAND2_X1 U11189 ( .A1(n13328), .A2(n13607), .ZN(n8655) );
  OR2_X1 U11190 ( .A1(n14036), .A2(n13606), .ZN(n8656) );
  XNOR2_X1 U11191 ( .A(n15525), .B(n13343), .ZN(n11171) );
  INV_X1 U11192 ( .A(n13343), .ZN(n13605) );
  XNOR2_X1 U11193 ( .A(n14031), .B(n13604), .ZN(n11360) );
  INV_X1 U11194 ( .A(n11360), .ZN(n8657) );
  NAND2_X1 U11195 ( .A1(n14031), .A2(n13604), .ZN(n11576) );
  AND2_X1 U11196 ( .A1(n11712), .A2(n11576), .ZN(n8658) );
  INV_X1 U11197 ( .A(n13358), .ZN(n13602) );
  OAI21_X1 U11198 ( .B1(n14026), .B2(n13602), .A(n8659), .ZN(n8660) );
  INV_X1 U11199 ( .A(n8660), .ZN(n8661) );
  NAND2_X1 U11200 ( .A1(n8662), .A2(n8661), .ZN(n8664) );
  NAND2_X1 U11201 ( .A1(n14026), .A2(n13602), .ZN(n8663) );
  NAND2_X1 U11202 ( .A1(n13365), .A2(n13601), .ZN(n8665) );
  INV_X1 U11203 ( .A(n13372), .ZN(n13600) );
  AND2_X1 U11204 ( .A1(n14085), .A2(n13600), .ZN(n8667) );
  OR2_X1 U11205 ( .A1(n14085), .A2(n13600), .ZN(n8666) );
  INV_X1 U11206 ( .A(n13552), .ZN(n13879) );
  NOR2_X1 U11207 ( .A1(n14014), .A2(n13879), .ZN(n8668) );
  INV_X1 U11208 ( .A(n14014), .ZN(n13905) );
  INV_X1 U11209 ( .A(n13386), .ZN(n13599) );
  XNOR2_X1 U11210 ( .A(n13866), .B(n13881), .ZN(n13869) );
  OR2_X1 U11211 ( .A1(n13866), .A2(n13881), .ZN(n8669) );
  INV_X1 U11212 ( .A(n13812), .ZN(n8671) );
  INV_X1 U11213 ( .A(n13833), .ZN(n8672) );
  AND2_X1 U11214 ( .A1(n13996), .A2(n13598), .ZN(n13830) );
  INV_X1 U11215 ( .A(n13409), .ZN(n13597) );
  AOI22_X1 U11216 ( .A1(n8672), .A2(n13830), .B1(n14073), .B2(n13597), .ZN(
        n8673) );
  XNOR2_X1 U11217 ( .A(n13821), .B(n13596), .ZN(n13817) );
  OR2_X1 U11218 ( .A1(n13821), .A2(n13596), .ZN(n8674) );
  NAND2_X1 U11219 ( .A1(n14065), .A2(n13782), .ZN(n8675) );
  OR2_X1 U11220 ( .A1(n14065), .A2(n13782), .ZN(n8676) );
  INV_X1 U11221 ( .A(n13972), .ZN(n13791) );
  XNOR2_X1 U11222 ( .A(n13432), .B(n13783), .ZN(n13766) );
  NAND2_X1 U11223 ( .A1(n14058), .A2(n13594), .ZN(n8679) );
  AND2_X1 U11224 ( .A1(n13956), .A2(n13593), .ZN(n13534) );
  OR2_X1 U11225 ( .A1(n13956), .A2(n13593), .ZN(n13535) );
  OR2_X1 U11226 ( .A1(n13722), .A2(n13592), .ZN(n8680) );
  NAND2_X1 U11227 ( .A1(n13722), .A2(n13592), .ZN(n8681) );
  NAND2_X1 U11228 ( .A1(n13933), .A2(n13591), .ZN(n8682) );
  NOR2_X1 U11229 ( .A1(n13571), .A2(n13568), .ZN(n8685) );
  NAND2_X1 U11230 ( .A1(n13913), .A2(n8685), .ZN(n11724) );
  NAND2_X1 U11231 ( .A1(n13913), .A2(n12152), .ZN(n8687) );
  INV_X1 U11232 ( .A(n14085), .ZN(n12080) );
  INV_X1 U11233 ( .A(n13352), .ZN(n11614) );
  INV_X1 U11234 ( .A(n14031), .ZN(n11366) );
  NAND2_X1 U11235 ( .A1(n12147), .A2(n15512), .ZN(n11207) );
  INV_X1 U11236 ( .A(n13328), .ZN(n11191) );
  INV_X1 U11237 ( .A(n13996), .ZN(n13857) );
  INV_X1 U11238 ( .A(n14073), .ZN(n13842) );
  INV_X1 U11239 ( .A(n13940), .ZN(n13712) );
  INV_X1 U11240 ( .A(n13933), .ZN(n13694) );
  INV_X1 U11241 ( .A(n13460), .ZN(n8692) );
  AND2_X1 U11242 ( .A1(n10884), .A2(n7902), .ZN(n10565) );
  NAND2_X2 U11243 ( .A1(n13913), .A2(n10565), .ZN(n13904) );
  INV_X1 U11244 ( .A(n8689), .ZN(n8690) );
  INV_X1 U11245 ( .A(n13843), .ZN(n13915) );
  INV_X1 U11246 ( .A(n13913), .ZN(n13797) );
  AOI22_X1 U11247 ( .A1(n8690), .A2(n13915), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n13797), .ZN(n8691) );
  OAI21_X1 U11248 ( .B1(n8692), .B2(n13904), .A(n8691), .ZN(n8693) );
  AOI21_X1 U11249 ( .B1(n15524), .B2(n13460), .A(n8697), .ZN(n8698) );
  NOR2_X1 U11250 ( .A1(n10559), .A2(n15509), .ZN(n15508) );
  AND2_X1 U11251 ( .A1(n10568), .A2(n10570), .ZN(n8701) );
  INV_X1 U11252 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n8702) );
  OR2_X1 U11253 ( .A1(n15533), .A2(n8702), .ZN(n8703) );
  NAND2_X1 U11254 ( .A1(n8704), .A2(n8703), .ZN(P2_U3496) );
  INV_X1 U11255 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n8732) );
  INV_X1 U11256 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n8728) );
  INV_X1 U11257 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n8726) );
  INV_X1 U11258 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n8724) );
  INV_X1 U11259 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n15749) );
  XNOR2_X1 U11260 ( .A(P1_ADDR_REG_11__SCAN_IN), .B(P3_ADDR_REG_11__SCAN_IN), 
        .ZN(n8771) );
  INV_X1 U11261 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n15774) );
  XNOR2_X1 U11262 ( .A(P1_ADDR_REG_10__SCAN_IN), .B(P3_ADDR_REG_10__SCAN_IN), 
        .ZN(n8767) );
  INV_X1 U11263 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n8719) );
  XNOR2_X1 U11264 ( .A(P3_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n8762) );
  XNOR2_X1 U11265 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), 
        .ZN(n8739) );
  NAND2_X1 U11266 ( .A1(n8738), .A2(n14591), .ZN(n8707) );
  NAND2_X1 U11267 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n8705), .ZN(n8706) );
  NAND2_X1 U11268 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n8708), .ZN(n8710) );
  INV_X1 U11269 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8709) );
  NAND2_X1 U11270 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n8711), .ZN(n8712) );
  INV_X1 U11271 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14620) );
  INV_X1 U11272 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15560) );
  NAND2_X1 U11273 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n15560), .ZN(n8713) );
  INV_X1 U11274 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11275 ( .A1(n8715), .A2(n8714), .ZN(n8717) );
  NAND2_X1 U11276 ( .A1(n8737), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n8716) );
  XNOR2_X1 U11277 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(n14664), .ZN(n8736) );
  XNOR2_X1 U11278 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(n8724), .ZN(n8734) );
  INV_X1 U11279 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n11314) );
  NOR2_X1 U11280 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n11314), .ZN(n8725) );
  XOR2_X1 U11281 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .Z(n8778) );
  INV_X1 U11282 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n11631) );
  OR2_X1 U11283 ( .A1(n11631), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n8729) );
  INV_X1 U11284 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U11285 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n11916), .ZN(n8730) );
  INV_X1 U11286 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n15734) );
  AOI22_X1 U11287 ( .A1(n8785), .A2(n8730), .B1(P1_ADDR_REG_16__SCAN_IN), .B2(
        n15734), .ZN(n8789) );
  INV_X1 U11288 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14691) );
  XOR2_X1 U11289 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14691), .Z(n8788) );
  NAND2_X1 U11290 ( .A1(n8789), .A2(n8788), .ZN(n8731) );
  OAI21_X1 U11291 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(n8732), .A(n8731), .ZN(
        n8793) );
  XOR2_X1 U11292 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n8792) );
  XNOR2_X1 U11293 ( .A(n8793), .B(n8792), .ZN(n15202) );
  XOR2_X1 U11294 ( .A(n8734), .B(n8733), .Z(n8772) );
  XOR2_X1 U11295 ( .A(n8736), .B(n8735), .Z(n15215) );
  XNOR2_X1 U11296 ( .A(n8737), .B(P1_ADDR_REG_7__SCAN_IN), .ZN(n15829) );
  XNOR2_X1 U11297 ( .A(n8738), .B(P1_ADDR_REG_3__SCAN_IN), .ZN(n15832) );
  XOR2_X1 U11298 ( .A(n8740), .B(n8739), .Z(n15207) );
  INV_X1 U11299 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n8745) );
  NOR2_X1 U11300 ( .A1(n8744), .A2(n8745), .ZN(n8746) );
  OAI21_X1 U11301 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(n8743), .A(n8742), .ZN(
        n15826) );
  NAND2_X1 U11302 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15826), .ZN(n15837) );
  NOR2_X1 U11303 ( .A1(n15207), .A2(n15206), .ZN(n8747) );
  NAND2_X1 U11304 ( .A1(n15207), .A2(n15206), .ZN(n15205) );
  NAND2_X1 U11305 ( .A1(n15832), .A2(n15831), .ZN(n8748) );
  NOR2_X1 U11306 ( .A1(n15832), .A2(n15831), .ZN(n15830) );
  INV_X1 U11307 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n15407) );
  XNOR2_X1 U11308 ( .A(n15407), .B(n8750), .ZN(n15821) );
  NOR2_X1 U11309 ( .A1(n15822), .A2(n15821), .ZN(n15820) );
  NOR2_X1 U11310 ( .A1(n8750), .A2(n15407), .ZN(n8751) );
  XNOR2_X1 U11311 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n8752), .ZN(n8753) );
  NAND2_X1 U11312 ( .A1(n8754), .A2(n8753), .ZN(n8756) );
  INV_X1 U11313 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15824) );
  INV_X1 U11314 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n8759) );
  XNOR2_X1 U11315 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n8758) );
  XOR2_X1 U11316 ( .A(n8758), .B(n8757), .Z(n15210) );
  INV_X1 U11317 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n13626) );
  XNOR2_X1 U11318 ( .A(n8762), .B(n8761), .ZN(n8763) );
  NAND2_X1 U11319 ( .A1(n8764), .A2(n8763), .ZN(n8765) );
  INV_X1 U11320 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n15801) );
  XOR2_X1 U11321 ( .A(n8767), .B(n8766), .Z(n8768) );
  INV_X1 U11322 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n15431) );
  NAND2_X1 U11323 ( .A1(n8769), .A2(n8768), .ZN(n15220) );
  XNOR2_X1 U11324 ( .A(n8771), .B(n8770), .ZN(n15224) );
  NAND2_X1 U11325 ( .A1(n8772), .A2(n8774), .ZN(n8775) );
  INV_X1 U11326 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15445) );
  XNOR2_X1 U11327 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n8777) );
  XNOR2_X1 U11328 ( .A(n8777), .B(n8776), .ZN(n15230) );
  XNOR2_X1 U11329 ( .A(n8779), .B(n8778), .ZN(n15234) );
  XOR2_X1 U11330 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .Z(n8781) );
  XOR2_X1 U11331 ( .A(n8782), .B(n8781), .Z(n8783) );
  INV_X1 U11332 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n15472) );
  XNOR2_X1 U11333 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n8786) );
  XNOR2_X1 U11334 ( .A(n8786), .B(n8785), .ZN(n8787) );
  INV_X1 U11335 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15485) );
  INV_X1 U11336 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n15501) );
  INV_X1 U11337 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n8795) );
  NOR2_X1 U11338 ( .A1(n8793), .A2(n8792), .ZN(n8794) );
  AOI21_X1 U11339 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n8795), .A(n8794), .ZN(
        n8798) );
  XNOR2_X1 U11340 ( .A(P3_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n8796) );
  XOR2_X1 U11341 ( .A(n8796), .B(P1_ADDR_REG_19__SCAN_IN), .Z(n8797) );
  XNOR2_X1 U11342 ( .A(n8798), .B(n8797), .ZN(n8799) );
  XNOR2_X1 U11343 ( .A(n8800), .B(n8799), .ZN(SUB_1596_U4) );
  INV_X1 U11344 ( .A(n8801), .ZN(n8802) );
  NAND2_X1 U11345 ( .A1(n13589), .A2(n13880), .ZN(n8806) );
  NAND2_X1 U11346 ( .A1(n13591), .A2(n13878), .ZN(n8805) );
  NAND2_X1 U11347 ( .A1(n8806), .A2(n8805), .ZN(n13146) );
  AOI21_X1 U11348 ( .B1(n13693), .B2(n13456), .A(n6409), .ZN(n8809) );
  NAND2_X1 U11349 ( .A1(n8809), .A2(n8808), .ZN(n11944) );
  NOR2_X2 U11350 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8832) );
  NOR2_X1 U11351 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n8814) );
  NOR2_X1 U11352 ( .A1(n15184), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n8824) );
  NAND2_X1 U11353 ( .A1(n10895), .A2(n8962), .ZN(n8839) );
  INV_X1 U11354 ( .A(n8997), .ZN(n8831) );
  INV_X1 U11355 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8830) );
  NAND2_X1 U11356 ( .A1(n8831), .A2(n8830), .ZN(n9019) );
  NOR2_X1 U11357 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n8833) );
  INV_X1 U11358 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9135) );
  NAND4_X1 U11359 ( .A1(n8834), .A2(n8832), .A3(n8833), .A4(n9135), .ZN(n8835)
         );
  NOR2_X1 U11360 ( .A1(n9056), .A2(n8835), .ZN(n9195) );
  INV_X1 U11361 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U11362 ( .A1(n9195), .A2(n8836), .ZN(n9198) );
  OAI21_X1 U11363 ( .B1(n9198), .B2(P1_IR_REG_16__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8837) );
  XNOR2_X1 U11364 ( .A(n8837), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14715) );
  INV_X2 U11365 ( .A(n14476), .ZN(n9243) );
  AOI22_X1 U11366 ( .A1(n14715), .A2(n10243), .B1(P2_DATAO_REG_17__SCAN_IN), 
        .B2(n9243), .ZN(n8838) );
  INV_X1 U11367 ( .A(n8840), .ZN(n8841) );
  NAND2_X1 U11368 ( .A1(n8841), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8842) );
  MUX2_X1 U11369 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8842), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n8844) );
  NAND2_X1 U11370 ( .A1(n8840), .A2(n8843), .ZN(n8846) );
  INV_X1 U11371 ( .A(n11564), .ZN(n9425) );
  NAND2_X1 U11372 ( .A1(n8846), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8845) );
  OAI21_X1 U11373 ( .B1(n8846), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n8847) );
  NAND2_X1 U11374 ( .A1(n8852), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8849) );
  INV_X1 U11375 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8853) );
  XNOR2_X2 U11376 ( .A(n8860), .B(n8859), .ZN(n14526) );
  INV_X1 U11377 ( .A(n9001), .ZN(n8861) );
  NAND2_X1 U11378 ( .A1(n9187), .A2(n14207), .ZN(n8865) );
  NAND2_X1 U11379 ( .A1(n9232), .A2(n8865), .ZN(n14957) );
  NAND2_X1 U11380 ( .A1(n14427), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8870) );
  INV_X1 U11381 ( .A(n14432), .ZN(n9122) );
  NAND2_X1 U11382 ( .A1(n9122), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n8869) );
  AND2_X1 U11383 ( .A1(n8870), .A2(n8869), .ZN(n8873) );
  INV_X2 U11384 ( .A(n9079), .ZN(n9314) );
  NAND2_X1 U11385 ( .A1(n9408), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8872) );
  OAI211_X1 U11386 ( .C1(n14957), .C2(n6439), .A(n8873), .B(n8872), .ZN(n14969) );
  AOI22_X1 U11387 ( .A1(n14960), .A2(n9397), .B1(n9395), .B2(n14969), .ZN(
        n9223) );
  INV_X1 U11388 ( .A(n9223), .ZN(n9225) );
  NAND2_X1 U11389 ( .A1(n14960), .A2(n9401), .ZN(n8875) );
  NAND2_X1 U11390 ( .A1(n14969), .A2(n9397), .ZN(n8874) );
  NAND2_X1 U11391 ( .A1(n8875), .A2(n8874), .ZN(n8877) );
  INV_X1 U11392 ( .A(n14286), .ZN(n15198) );
  NAND2_X1 U11393 ( .A1(n15198), .A2(n14526), .ZN(n8876) );
  XNOR2_X1 U11394 ( .A(n8877), .B(n9380), .ZN(n9224) );
  INV_X1 U11395 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n8878) );
  OR2_X1 U11396 ( .A1(n14432), .A2(n8878), .ZN(n8884) );
  INV_X1 U11397 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n10611) );
  INV_X1 U11398 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n8879) );
  OR2_X1 U11399 ( .A1(n9079), .A2(n8879), .ZN(n8881) );
  NAND2_X1 U11400 ( .A1(n8925), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n8880) );
  NAND2_X1 U11401 ( .A1(n8892), .A2(n6436), .ZN(n8890) );
  NAND2_X1 U11402 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8885) );
  MUX2_X1 U11403 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8885), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8887) );
  INV_X1 U11404 ( .A(n8886), .ZN(n8931) );
  NAND2_X1 U11405 ( .A1(n8887), .A2(n8931), .ZN(n10264) );
  NAND2_X1 U11406 ( .A1(n14295), .A2(n8888), .ZN(n8889) );
  NAND2_X1 U11407 ( .A1(n8890), .A2(n8889), .ZN(n8891) );
  XNOR2_X1 U11408 ( .A(n8891), .B(n10810), .ZN(n8895) );
  AND2_X1 U11409 ( .A1(n14295), .A2(n6436), .ZN(n8893) );
  AOI21_X1 U11410 ( .B1(n8892), .B2(n9324), .A(n8893), .ZN(n8894) );
  OR2_X1 U11411 ( .A1(n8895), .A2(n8894), .ZN(n8896) );
  NAND2_X1 U11412 ( .A1(n8895), .A2(n8894), .ZN(n8922) );
  AOI22_X1 U11413 ( .A1(n7174), .A2(P1_REG2_REG_0__SCAN_IN), .B1(
        P1_IR_REG_30__SCAN_IN), .B2(P1_REG0_REG_0__SCAN_IN), .ZN(n8902) );
  INV_X1 U11414 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n8899) );
  NAND2_X1 U11415 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n8898) );
  OAI21_X1 U11416 ( .B1(n8899), .B2(P1_IR_REG_30__SCAN_IN), .A(n8898), .ZN(
        n8900) );
  NAND2_X1 U11417 ( .A1(n8897), .A2(n8900), .ZN(n8901) );
  OAI21_X1 U11418 ( .B1(n8897), .B2(n8902), .A(n8901), .ZN(n8903) );
  NAND2_X1 U11419 ( .A1(n8903), .A2(n8871), .ZN(n8911) );
  AOI22_X1 U11420 ( .A1(n7174), .A2(P1_REG3_REG_0__SCAN_IN), .B1(
        P1_REG1_REG_0__SCAN_IN), .B2(P1_IR_REG_30__SCAN_IN), .ZN(n8907) );
  INV_X1 U11421 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U11422 ( .A1(P1_IR_REG_30__SCAN_IN), .A2(P1_REG3_REG_0__SCAN_IN), 
        .ZN(n8904) );
  OAI21_X1 U11423 ( .B1(n8917), .B2(P1_IR_REG_30__SCAN_IN), .A(n8904), .ZN(
        n8905) );
  NAND2_X1 U11424 ( .A1(n8897), .A2(n8905), .ZN(n8906) );
  OAI21_X1 U11425 ( .B1(n8897), .B2(n8907), .A(n8906), .ZN(n8909) );
  NAND2_X1 U11426 ( .A1(n8909), .A2(n8908), .ZN(n8910) );
  OR2_X1 U11427 ( .A1(n9418), .A2(n10904), .ZN(n8916) );
  INV_X1 U11428 ( .A(SI_0_), .ZN(n9511) );
  INV_X1 U11429 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n9509) );
  OAI21_X1 U11430 ( .B1(n7875), .B2(n9511), .A(n9509), .ZN(n8912) );
  AND2_X1 U11431 ( .A1(n8913), .A2(n8912), .ZN(n15199) );
  MUX2_X1 U11432 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15199), .S(n6435), .Z(n15276)
         );
  INV_X1 U11433 ( .A(n10106), .ZN(n8914) );
  AOI22_X1 U11434 ( .A1(n15276), .A2(n6436), .B1(P1_IR_REG_0__SCAN_IN), .B2(
        n8914), .ZN(n8915) );
  AND2_X1 U11435 ( .A1(n8916), .A2(n8915), .ZN(n10292) );
  NOR2_X1 U11436 ( .A1(n10106), .A2(n8917), .ZN(n8918) );
  AOI21_X1 U11437 ( .B1(n15276), .B2(n9401), .A(n8918), .ZN(n8920) );
  INV_X1 U11438 ( .A(n10904), .ZN(n14558) );
  NAND2_X1 U11439 ( .A1(n14558), .A2(n6436), .ZN(n8919) );
  NAND2_X1 U11440 ( .A1(n8920), .A2(n8919), .ZN(n10291) );
  NAND2_X1 U11441 ( .A1(n10292), .A2(n10291), .ZN(n10290) );
  OR2_X1 U11442 ( .A1(n10291), .A2(n10810), .ZN(n8921) );
  INV_X1 U11443 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8923) );
  OR2_X1 U11444 ( .A1(n14432), .A2(n8923), .ZN(n8930) );
  INV_X1 U11445 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n8924) );
  NAND2_X1 U11446 ( .A1(n8925), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n8928) );
  INV_X1 U11447 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n8926) );
  OR2_X1 U11448 ( .A1(n9079), .A2(n8926), .ZN(n8927) );
  NAND2_X1 U11449 ( .A1(n14557), .A2(n6436), .ZN(n8937) );
  NAND2_X1 U11450 ( .A1(n8931), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8932) );
  MUX2_X1 U11451 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8932), .S(
        P1_IR_REG_2__SCAN_IN), .Z(n8933) );
  NAND2_X1 U11452 ( .A1(n8933), .A2(n8944), .ZN(n10267) );
  OR2_X1 U11453 ( .A1(n14476), .A2(n10166), .ZN(n8935) );
  OR2_X1 U11454 ( .A1(n12036), .A2(n10165), .ZN(n8934) );
  INV_X2 U11455 ( .A(n9301), .ZN(n9387) );
  NAND2_X1 U11456 ( .A1(n15261), .A2(n9401), .ZN(n8936) );
  NAND2_X1 U11457 ( .A1(n8937), .A2(n8936), .ZN(n8938) );
  AND2_X1 U11458 ( .A1(n15261), .A2(n6436), .ZN(n8939) );
  AOI21_X1 U11459 ( .B1(n14557), .B2(n9395), .A(n8939), .ZN(n8954) );
  XNOR2_X1 U11460 ( .A(n8953), .B(n8954), .ZN(n10758) );
  INV_X1 U11461 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10252) );
  OR2_X1 U11462 ( .A1(n14432), .A2(n10252), .ZN(n8943) );
  NAND2_X1 U11463 ( .A1(n9314), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n8942) );
  OR2_X1 U11464 ( .A1(n6439), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8941) );
  NAND2_X1 U11465 ( .A1(n8925), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n8940) );
  NAND2_X1 U11466 ( .A1(n14556), .A2(n6436), .ZN(n8950) );
  NAND2_X1 U11467 ( .A1(n8944), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8946) );
  INV_X1 U11468 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n8945) );
  OR2_X1 U11469 ( .A1(n10167), .A2(n12036), .ZN(n8948) );
  OR2_X1 U11470 ( .A1(n14476), .A2(n10168), .ZN(n8947) );
  NAND2_X1 U11471 ( .A1(n14148), .A2(n9387), .ZN(n8949) );
  NAND2_X1 U11472 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  XNOR2_X1 U11473 ( .A(n8951), .B(n9380), .ZN(n8974) );
  AND2_X1 U11474 ( .A1(n14148), .A2(n6436), .ZN(n8952) );
  AOI21_X1 U11475 ( .B1(n14556), .B2(n9395), .A(n8952), .ZN(n8972) );
  XNOR2_X1 U11476 ( .A(n8974), .B(n8972), .ZN(n14144) );
  INV_X1 U11477 ( .A(n8953), .ZN(n8955) );
  NAND2_X1 U11478 ( .A1(n8955), .A2(n8954), .ZN(n14140) );
  AND2_X1 U11479 ( .A1(n14144), .A2(n14140), .ZN(n8956) );
  NAND2_X1 U11480 ( .A1(n14141), .A2(n8956), .ZN(n11075) );
  NAND2_X1 U11481 ( .A1(n9314), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n8961) );
  NAND2_X1 U11482 ( .A1(n14427), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n8960) );
  XNOR2_X1 U11483 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11151) );
  OR2_X1 U11484 ( .A1(n6439), .A2(n11151), .ZN(n8959) );
  INV_X1 U11485 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n8957) );
  OR2_X1 U11486 ( .A1(n14432), .A2(n8957), .ZN(n8958) );
  NAND2_X1 U11487 ( .A1(n14555), .A2(n9397), .ZN(n8969) );
  NAND2_X1 U11488 ( .A1(n10160), .A2(n8962), .ZN(n8967) );
  NAND2_X1 U11489 ( .A1(n8963), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8964) );
  MUX2_X1 U11490 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8964), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n8965) );
  NAND2_X1 U11491 ( .A1(n8965), .A2(n8984), .ZN(n10272) );
  OR2_X1 U11492 ( .A1(n6435), .A2(n10272), .ZN(n8966) );
  OAI211_X1 U11493 ( .C1(n14476), .C2(n10170), .A(n8967), .B(n8966), .ZN(
        n14309) );
  NAND2_X1 U11494 ( .A1(n14309), .A2(n9387), .ZN(n8968) );
  NAND2_X1 U11495 ( .A1(n8969), .A2(n8968), .ZN(n8970) );
  XNOR2_X1 U11496 ( .A(n8970), .B(n10810), .ZN(n11148) );
  AND2_X1 U11497 ( .A1(n14309), .A2(n9397), .ZN(n8971) );
  AOI21_X1 U11498 ( .B1(n14555), .B2(n9395), .A(n8971), .ZN(n11077) );
  INV_X1 U11499 ( .A(n8972), .ZN(n8973) );
  NAND2_X1 U11500 ( .A1(n8974), .A2(n8973), .ZN(n11076) );
  NAND2_X1 U11501 ( .A1(n11075), .A2(n8976), .ZN(n8992) );
  NAND2_X1 U11502 ( .A1(n9314), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n8983) );
  NAND2_X1 U11503 ( .A1(n14427), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8982) );
  INV_X1 U11504 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n8978) );
  NAND2_X1 U11505 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8977) );
  NAND2_X1 U11506 ( .A1(n8978), .A2(n8977), .ZN(n8979) );
  NAND2_X1 U11507 ( .A1(n9001), .A2(n8979), .ZN(n11140) );
  OR2_X1 U11508 ( .A1(n6439), .A2(n11140), .ZN(n8981) );
  OR2_X1 U11509 ( .A1(n14432), .A2(n15360), .ZN(n8980) );
  NAND2_X1 U11510 ( .A1(n14554), .A2(n9397), .ZN(n8990) );
  NAND2_X1 U11511 ( .A1(n10176), .A2(n8962), .ZN(n8988) );
  NAND2_X1 U11512 ( .A1(n8984), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8985) );
  MUX2_X1 U11513 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8985), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n8986) );
  AND2_X1 U11514 ( .A1(n8986), .A2(n8997), .ZN(n14622) );
  AOI22_X1 U11515 ( .A1(n9243), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n10243), 
        .B2(n14622), .ZN(n8987) );
  NAND2_X1 U11516 ( .A1(n14313), .A2(n9387), .ZN(n8989) );
  NAND2_X1 U11517 ( .A1(n8990), .A2(n8989), .ZN(n8991) );
  XNOR2_X1 U11518 ( .A(n8991), .B(n10810), .ZN(n8993) );
  AOI22_X1 U11519 ( .A1(n14554), .A2(n9395), .B1(n6436), .B2(n14313), .ZN(
        n8994) );
  NAND2_X1 U11520 ( .A1(n8993), .A2(n8994), .ZN(n11079) );
  INV_X1 U11521 ( .A(n8993), .ZN(n8996) );
  INV_X1 U11522 ( .A(n8994), .ZN(n8995) );
  NAND2_X1 U11523 ( .A1(n8996), .A2(n8995), .ZN(n11080) );
  NAND2_X1 U11524 ( .A1(n10180), .A2(n8962), .ZN(n9000) );
  NAND2_X1 U11525 ( .A1(n8997), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8998) );
  XNOR2_X1 U11526 ( .A(n8998), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10481) );
  AOI22_X1 U11527 ( .A1(n9243), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n10243), 
        .B2(n10481), .ZN(n8999) );
  NAND2_X1 U11528 ( .A1(n14319), .A2(n9387), .ZN(n9009) );
  NAND2_X1 U11529 ( .A1(n9314), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11530 ( .A1(n14427), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9006) );
  INV_X1 U11531 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n15783) );
  NAND2_X1 U11532 ( .A1(n9001), .A2(n15783), .ZN(n9002) );
  NAND2_X1 U11533 ( .A1(n9024), .A2(n9002), .ZN(n11352) );
  OR2_X1 U11534 ( .A1(n6439), .A2(n11352), .ZN(n9005) );
  INV_X1 U11535 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n9003) );
  OR2_X1 U11536 ( .A1(n14432), .A2(n9003), .ZN(n9004) );
  NAND4_X2 U11537 ( .A1(n9007), .A2(n9006), .A3(n9005), .A4(n9004), .ZN(n14553) );
  NAND2_X1 U11538 ( .A1(n14553), .A2(n9397), .ZN(n9008) );
  NAND2_X1 U11539 ( .A1(n9009), .A2(n9008), .ZN(n9010) );
  XNOR2_X1 U11540 ( .A(n9010), .B(n9380), .ZN(n9014) );
  NAND2_X1 U11541 ( .A1(n14319), .A2(n9397), .ZN(n9012) );
  NAND2_X1 U11542 ( .A1(n14553), .A2(n9395), .ZN(n9011) );
  NAND2_X1 U11543 ( .A1(n9012), .A2(n9011), .ZN(n9015) );
  AND2_X1 U11544 ( .A1(n9014), .A2(n9015), .ZN(n11156) );
  INV_X1 U11545 ( .A(n11156), .ZN(n9013) );
  INV_X1 U11546 ( .A(n9014), .ZN(n9017) );
  INV_X1 U11547 ( .A(n9015), .ZN(n9016) );
  NAND2_X1 U11548 ( .A1(n9017), .A2(n9016), .ZN(n11155) );
  NAND2_X1 U11549 ( .A1(n9018), .A2(n11155), .ZN(n14104) );
  NAND2_X1 U11550 ( .A1(n10194), .A2(n8962), .ZN(n9022) );
  NAND2_X1 U11551 ( .A1(n9019), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9020) );
  XNOR2_X1 U11552 ( .A(n9020), .B(P1_IR_REG_7__SCAN_IN), .ZN(n14636) );
  AOI22_X1 U11553 ( .A1(n9243), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n10243), 
        .B2(n14636), .ZN(n9021) );
  NAND2_X1 U11554 ( .A1(n14325), .A2(n9387), .ZN(n9030) );
  NAND2_X1 U11555 ( .A1(n14427), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n9028) );
  NAND2_X1 U11556 ( .A1(n9314), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9027) );
  INV_X1 U11557 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n9023) );
  NAND2_X1 U11558 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  NAND2_X1 U11559 ( .A1(n9039), .A2(n9025), .ZN(n14109) );
  INV_X1 U11560 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10467) );
  OR2_X1 U11561 ( .A1(n14432), .A2(n10467), .ZN(n9026) );
  NAND2_X1 U11562 ( .A1(n14552), .A2(n9397), .ZN(n9029) );
  NAND2_X1 U11563 ( .A1(n9030), .A2(n9029), .ZN(n9031) );
  XNOR2_X1 U11564 ( .A(n9031), .B(n10810), .ZN(n9033) );
  AND2_X1 U11565 ( .A1(n14552), .A2(n9395), .ZN(n9032) );
  AOI21_X1 U11566 ( .B1(n14325), .B2(n6436), .A(n9032), .ZN(n9034) );
  XNOR2_X1 U11567 ( .A(n9033), .B(n9034), .ZN(n14105) );
  NAND2_X1 U11568 ( .A1(n10234), .A2(n8962), .ZN(n9037) );
  NAND2_X1 U11569 ( .A1(n9056), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9035) );
  XNOR2_X1 U11570 ( .A(n9035), .B(P1_IR_REG_8__SCAN_IN), .ZN(n14648) );
  AOI22_X1 U11571 ( .A1(n9243), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n10243), 
        .B2(n14648), .ZN(n9036) );
  NAND2_X1 U11572 ( .A1(n15335), .A2(n9401), .ZN(n9046) );
  NAND2_X1 U11573 ( .A1(n9314), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n9044) );
  NAND2_X1 U11574 ( .A1(n14427), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9043) );
  INV_X1 U11575 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U11576 ( .A1(n9039), .A2(n9038), .ZN(n9040) );
  NAND2_X1 U11577 ( .A1(n9061), .A2(n9040), .ZN(n11570) );
  OR2_X1 U11578 ( .A1(n6438), .A2(n11570), .ZN(n9042) );
  INV_X1 U11579 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10469) );
  OR2_X1 U11580 ( .A1(n14432), .A2(n10469), .ZN(n9041) );
  NAND4_X1 U11581 ( .A1(n9044), .A2(n9043), .A3(n9042), .A4(n9041), .ZN(n14551) );
  NAND2_X1 U11582 ( .A1(n14551), .A2(n6436), .ZN(n9045) );
  NAND2_X1 U11583 ( .A1(n9046), .A2(n9045), .ZN(n9047) );
  XNOR2_X1 U11584 ( .A(n9047), .B(n10810), .ZN(n9049) );
  AND2_X1 U11585 ( .A1(n14551), .A2(n9395), .ZN(n9048) );
  AOI21_X1 U11586 ( .B1(n15335), .B2(n9397), .A(n9048), .ZN(n9050) );
  NAND2_X1 U11587 ( .A1(n9049), .A2(n9050), .ZN(n9054) );
  INV_X1 U11588 ( .A(n9049), .ZN(n9052) );
  INV_X1 U11589 ( .A(n9050), .ZN(n9051) );
  NAND2_X1 U11590 ( .A1(n9052), .A2(n9051), .ZN(n9053) );
  NAND2_X1 U11591 ( .A1(n9054), .A2(n9053), .ZN(n11568) );
  INV_X1 U11592 ( .A(n9054), .ZN(n9055) );
  NAND2_X1 U11593 ( .A1(n10239), .A2(n8962), .ZN(n9059) );
  XNOR2_X1 U11594 ( .A(n9101), .B(P1_IR_REG_9__SCAN_IN), .ZN(n14666) );
  AOI22_X1 U11595 ( .A1(n9243), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n10243), 
        .B2(n14666), .ZN(n9058) );
  NAND2_X1 U11596 ( .A1(n14344), .A2(n9401), .ZN(n9068) );
  NAND2_X1 U11597 ( .A1(n14427), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9066) );
  NAND2_X1 U11598 ( .A1(n9314), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n9065) );
  NAND2_X1 U11599 ( .A1(n9061), .A2(n9060), .ZN(n9062) );
  NAND2_X1 U11600 ( .A1(n9077), .A2(n9062), .ZN(n11892) );
  OR2_X1 U11601 ( .A1(n6438), .A2(n11892), .ZN(n9064) );
  INV_X1 U11602 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10471) );
  OR2_X1 U11603 ( .A1(n14432), .A2(n10471), .ZN(n9063) );
  NAND4_X1 U11604 ( .A1(n9066), .A2(n9065), .A3(n9064), .A4(n9063), .ZN(n14550) );
  NAND2_X1 U11605 ( .A1(n14550), .A2(n9397), .ZN(n9067) );
  NAND2_X1 U11606 ( .A1(n9068), .A2(n9067), .ZN(n9069) );
  XNOR2_X1 U11607 ( .A(n9069), .B(n10810), .ZN(n11890) );
  AND2_X1 U11608 ( .A1(n14550), .A2(n9324), .ZN(n9070) );
  AOI21_X1 U11609 ( .B1(n14344), .B2(n9397), .A(n9070), .ZN(n9090) );
  NAND2_X1 U11610 ( .A1(n11890), .A2(n9090), .ZN(n9071) );
  INV_X1 U11611 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n9072) );
  NAND2_X1 U11612 ( .A1(n9101), .A2(n9072), .ZN(n9073) );
  NAND2_X1 U11613 ( .A1(n9073), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9074) );
  XNOR2_X1 U11614 ( .A(n9074), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U11615 ( .A1(n10243), .A2(n10841), .B1(n9243), .B2(
        P2_DATAO_REG_10__SCAN_IN), .ZN(n9075) );
  NAND2_X1 U11616 ( .A1(n14350), .A2(n9401), .ZN(n9086) );
  NAND2_X1 U11617 ( .A1(n14427), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9084) );
  NAND2_X1 U11618 ( .A1(n9122), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U11619 ( .A1(n9077), .A2(n9076), .ZN(n9078) );
  NAND2_X1 U11620 ( .A1(n9106), .A2(n9078), .ZN(n11884) );
  OR2_X1 U11621 ( .A1(n6438), .A2(n11884), .ZN(n9082) );
  INV_X1 U11622 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9080) );
  OR2_X1 U11623 ( .A1(n9079), .A2(n9080), .ZN(n9081) );
  NAND4_X1 U11624 ( .A1(n9084), .A2(n9083), .A3(n9082), .A4(n9081), .ZN(n14549) );
  NAND2_X1 U11625 ( .A1(n14549), .A2(n9397), .ZN(n9085) );
  NAND2_X1 U11626 ( .A1(n9086), .A2(n9085), .ZN(n9087) );
  XNOR2_X1 U11627 ( .A(n9087), .B(n9380), .ZN(n9095) );
  NAND2_X1 U11628 ( .A1(n14350), .A2(n9397), .ZN(n9089) );
  NAND2_X1 U11629 ( .A1(n14549), .A2(n9395), .ZN(n9088) );
  NAND2_X1 U11630 ( .A1(n9089), .A2(n9088), .ZN(n9096) );
  NAND2_X1 U11631 ( .A1(n9095), .A2(n9096), .ZN(n11877) );
  INV_X1 U11632 ( .A(n11890), .ZN(n9091) );
  INV_X1 U11633 ( .A(n9090), .ZN(n11874) );
  NAND2_X1 U11634 ( .A1(n9091), .A2(n11874), .ZN(n9092) );
  AND2_X1 U11635 ( .A1(n11877), .A2(n9092), .ZN(n9093) );
  NAND2_X1 U11636 ( .A1(n9094), .A2(n9093), .ZN(n11878) );
  INV_X1 U11637 ( .A(n9095), .ZN(n9098) );
  INV_X1 U11638 ( .A(n9096), .ZN(n9097) );
  NAND2_X1 U11639 ( .A1(n9098), .A2(n9097), .ZN(n11879) );
  NAND2_X1 U11640 ( .A1(n11878), .A2(n11879), .ZN(n11865) );
  NAND2_X1 U11641 ( .A1(n10457), .A2(n8962), .ZN(n9104) );
  INV_X1 U11642 ( .A(n8832), .ZN(n9099) );
  NAND2_X1 U11643 ( .A1(n9099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9100) );
  NAND2_X1 U11644 ( .A1(n9101), .A2(n9100), .ZN(n9120) );
  INV_X1 U11645 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U11646 ( .A(n9120), .B(n9102), .ZN(n14679) );
  AOI22_X1 U11647 ( .A1(P2_DATAO_REG_11__SCAN_IN), .A2(n9243), .B1(n14679), 
        .B2(n10243), .ZN(n9103) );
  NAND2_X2 U11648 ( .A1(n9104), .A2(n9103), .ZN(n15154) );
  NAND2_X1 U11649 ( .A1(n15154), .A2(n9401), .ZN(n9113) );
  NAND2_X1 U11650 ( .A1(n9408), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n9111) );
  NAND2_X1 U11651 ( .A1(n14427), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9110) );
  INV_X1 U11652 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U11653 ( .A1(n9106), .A2(n9105), .ZN(n9107) );
  NAND2_X1 U11654 ( .A1(n9125), .A2(n9107), .ZN(n11868) );
  OR2_X1 U11655 ( .A1(n6438), .A2(n11868), .ZN(n9109) );
  INV_X1 U11656 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10844) );
  OR2_X1 U11657 ( .A1(n14432), .A2(n10844), .ZN(n9108) );
  NAND4_X1 U11658 ( .A1(n9111), .A2(n9110), .A3(n9109), .A4(n9108), .ZN(n14548) );
  NAND2_X1 U11659 ( .A1(n14548), .A2(n9397), .ZN(n9112) );
  NAND2_X1 U11660 ( .A1(n9113), .A2(n9112), .ZN(n9114) );
  XNOR2_X1 U11661 ( .A(n9114), .B(n9380), .ZN(n9116) );
  AND2_X1 U11662 ( .A1(n14548), .A2(n9395), .ZN(n9115) );
  AOI21_X1 U11663 ( .B1(n15154), .B2(n9397), .A(n9115), .ZN(n9117) );
  XNOR2_X1 U11664 ( .A(n9116), .B(n9117), .ZN(n11866) );
  INV_X1 U11665 ( .A(n9116), .ZN(n9118) );
  NAND2_X1 U11666 ( .A1(n9118), .A2(n9117), .ZN(n9119) );
  OAI21_X1 U11667 ( .B1(n9120), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9136) );
  XNOR2_X1 U11668 ( .A(n9136), .B(P1_IR_REG_12__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U11669 ( .A1(n11305), .A2(n10243), .B1(n9243), .B2(
        P2_DATAO_REG_12__SCAN_IN), .ZN(n9121) );
  NAND2_X1 U11670 ( .A1(n15149), .A2(n9387), .ZN(n9132) );
  NAND2_X1 U11671 ( .A1(n9408), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n9130) );
  NAND2_X1 U11672 ( .A1(n9122), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9129) );
  INV_X1 U11673 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9123) );
  OR2_X1 U11674 ( .A1(n9207), .A2(n9123), .ZN(n9128) );
  INV_X1 U11675 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n9124) );
  NAND2_X1 U11676 ( .A1(n9125), .A2(n9124), .ZN(n9126) );
  NAND2_X1 U11677 ( .A1(n9142), .A2(n9126), .ZN(n14171) );
  OR2_X1 U11678 ( .A1(n6438), .A2(n14171), .ZN(n9127) );
  NAND4_X1 U11679 ( .A1(n9130), .A2(n9129), .A3(n9128), .A4(n9127), .ZN(n14547) );
  NAND2_X1 U11680 ( .A1(n14547), .A2(n9397), .ZN(n9131) );
  NAND2_X1 U11681 ( .A1(n9132), .A2(n9131), .ZN(n9133) );
  XNOR2_X1 U11682 ( .A(n9133), .B(n10810), .ZN(n9151) );
  AND2_X1 U11683 ( .A1(n14547), .A2(n9324), .ZN(n9134) );
  AOI21_X1 U11684 ( .B1(n15149), .B2(n9397), .A(n9134), .ZN(n9152) );
  XNOR2_X1 U11685 ( .A(n9151), .B(n9152), .ZN(n14169) );
  NAND2_X1 U11686 ( .A1(n9136), .A2(n9135), .ZN(n9137) );
  NAND2_X1 U11687 ( .A1(n9137), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9139) );
  INV_X1 U11688 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9138) );
  NAND2_X1 U11689 ( .A1(n9139), .A2(n9138), .ZN(n9160) );
  OR2_X1 U11690 ( .A1(n9139), .A2(n9138), .ZN(n9140) );
  AOI22_X1 U11691 ( .A1(n11377), .A2(n10243), .B1(n9243), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n9141) );
  NAND2_X1 U11692 ( .A1(n9408), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n9147) );
  NAND2_X1 U11693 ( .A1(n14427), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9146) );
  NAND2_X1 U11694 ( .A1(n9142), .A2(n11311), .ZN(n9143) );
  NAND2_X1 U11695 ( .A1(n9165), .A2(n9143), .ZN(n14234) );
  OR2_X1 U11696 ( .A1(n6439), .A2(n14234), .ZN(n9145) );
  INV_X1 U11697 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n15748) );
  OR2_X1 U11698 ( .A1(n14432), .A2(n15748), .ZN(n9144) );
  NAND4_X1 U11699 ( .A1(n9147), .A2(n9146), .A3(n9145), .A4(n9144), .ZN(n15009) );
  XNOR2_X1 U11700 ( .A(n9148), .B(n9380), .ZN(n9158) );
  AND2_X1 U11701 ( .A1(n15009), .A2(n9395), .ZN(n9149) );
  AOI21_X1 U11702 ( .B1(n15144), .B2(n9397), .A(n9149), .ZN(n9156) );
  XNOR2_X1 U11703 ( .A(n9158), .B(n9156), .ZN(n14232) );
  INV_X1 U11704 ( .A(n14232), .ZN(n9155) );
  OR2_X1 U11705 ( .A1(n14169), .A2(n9155), .ZN(n9150) );
  INV_X1 U11706 ( .A(n9151), .ZN(n9154) );
  INV_X1 U11707 ( .A(n9152), .ZN(n9153) );
  NAND2_X1 U11708 ( .A1(n9154), .A2(n9153), .ZN(n14229) );
  INV_X1 U11709 ( .A(n9156), .ZN(n9157) );
  NAND2_X1 U11710 ( .A1(n9158), .A2(n9157), .ZN(n9159) );
  NAND2_X1 U11711 ( .A1(n10763), .A2(n8962), .ZN(n9163) );
  NAND2_X1 U11712 ( .A1(n9160), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9161) );
  AOI22_X1 U11713 ( .A1(n11627), .A2(n10243), .B1(P2_DATAO_REG_14__SCAN_IN), 
        .B2(n9243), .ZN(n9162) );
  NAND2_X2 U11714 ( .A1(n9163), .A2(n9162), .ZN(n15136) );
  NAND2_X1 U11715 ( .A1(n15136), .A2(n9387), .ZN(n9172) );
  NAND2_X1 U11716 ( .A1(n9408), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n9170) );
  NAND2_X1 U11717 ( .A1(n14427), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9169) );
  INV_X1 U11718 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n9164) );
  NAND2_X1 U11719 ( .A1(n9165), .A2(n9164), .ZN(n9166) );
  NAND2_X1 U11720 ( .A1(n9204), .A2(n9166), .ZN(n15007) );
  OR2_X1 U11721 ( .A1(n6438), .A2(n15007), .ZN(n9168) );
  INV_X1 U11722 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11370) );
  OR2_X1 U11723 ( .A1(n14432), .A2(n11370), .ZN(n9167) );
  NAND4_X1 U11724 ( .A1(n9170), .A2(n9169), .A3(n9168), .A4(n9167), .ZN(n14546) );
  NAND2_X1 U11725 ( .A1(n14546), .A2(n9397), .ZN(n9171) );
  NAND2_X1 U11726 ( .A1(n9172), .A2(n9171), .ZN(n9173) );
  XNOR2_X1 U11727 ( .A(n9173), .B(n10810), .ZN(n9177) );
  AND2_X1 U11728 ( .A1(n14546), .A2(n9395), .ZN(n9174) );
  AOI21_X1 U11729 ( .B1(n15136), .B2(n9397), .A(n9174), .ZN(n9176) );
  XNOR2_X1 U11730 ( .A(n9177), .B(n9176), .ZN(n14125) );
  INV_X1 U11731 ( .A(n14125), .ZN(n9175) );
  NAND2_X1 U11732 ( .A1(n9177), .A2(n9176), .ZN(n9178) );
  NAND2_X1 U11733 ( .A1(n10747), .A2(n8962), .ZN(n9181) );
  NAND2_X1 U11734 ( .A1(n9198), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9179) );
  XNOR2_X1 U11735 ( .A(n9179), .B(P1_IR_REG_16__SCAN_IN), .ZN(n14694) );
  AOI22_X1 U11736 ( .A1(n14694), .A2(n10243), .B1(n9243), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n9180) );
  NAND2_X1 U11737 ( .A1(n15122), .A2(n9401), .ZN(n9192) );
  INV_X1 U11738 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9183) );
  NAND2_X1 U11739 ( .A1(n14427), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9182) );
  OAI21_X1 U11740 ( .B1(n14432), .B2(n9183), .A(n9182), .ZN(n9190) );
  INV_X1 U11741 ( .A(n9184), .ZN(n9206) );
  INV_X1 U11742 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9185) );
  NAND2_X1 U11743 ( .A1(n9206), .A2(n9185), .ZN(n9186) );
  NAND2_X1 U11744 ( .A1(n9187), .A2(n9186), .ZN(n14978) );
  NAND2_X1 U11745 ( .A1(n9408), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n9188) );
  OAI21_X1 U11746 ( .B1(n14978), .B2(n6439), .A(n9188), .ZN(n9189) );
  NAND2_X1 U11747 ( .A1(n14954), .A2(n9397), .ZN(n9191) );
  NAND2_X1 U11748 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  XNOR2_X1 U11749 ( .A(n9193), .B(n10810), .ZN(n14188) );
  AND2_X1 U11750 ( .A1(n14954), .A2(n9324), .ZN(n9194) );
  AOI21_X1 U11751 ( .B1(n15122), .B2(n9397), .A(n9194), .ZN(n14187) );
  NAND2_X1 U11752 ( .A1(n10829), .A2(n8962), .ZN(n9202) );
  INV_X1 U11753 ( .A(n9195), .ZN(n9196) );
  NAND2_X1 U11754 ( .A1(n9196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9197) );
  MUX2_X1 U11755 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9197), .S(
        P1_IR_REG_15__SCAN_IN), .Z(n9199) );
  NAND2_X1 U11756 ( .A1(n9199), .A2(n9198), .ZN(n11900) );
  OAI22_X1 U11757 ( .A1(n14476), .A2(n10831), .B1(n11900), .B2(n6434), .ZN(
        n9200) );
  INV_X1 U11758 ( .A(n9200), .ZN(n9201) );
  NAND2_X1 U11759 ( .A1(n15130), .A2(n9401), .ZN(n9213) );
  INV_X1 U11760 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n9203) );
  NAND2_X1 U11761 ( .A1(n9204), .A2(n9203), .ZN(n9205) );
  NAND2_X1 U11762 ( .A1(n9206), .A2(n9205), .ZN(n14986) );
  OR2_X1 U11763 ( .A1(n14986), .A2(n6439), .ZN(n9211) );
  NAND2_X1 U11764 ( .A1(n9408), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n9210) );
  INV_X1 U11765 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n14992) );
  OR2_X1 U11766 ( .A1(n9207), .A2(n14992), .ZN(n9209) );
  INV_X1 U11767 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n11898) );
  OR2_X1 U11768 ( .A1(n14432), .A2(n11898), .ZN(n9208) );
  NAND4_X1 U11769 ( .A1(n9211), .A2(n9210), .A3(n9209), .A4(n9208), .ZN(n15011) );
  NAND2_X1 U11770 ( .A1(n15011), .A2(n9397), .ZN(n9212) );
  NAND2_X1 U11771 ( .A1(n9213), .A2(n9212), .ZN(n9214) );
  XNOR2_X1 U11772 ( .A(n9214), .B(n9380), .ZN(n14190) );
  NAND2_X1 U11773 ( .A1(n15130), .A2(n9397), .ZN(n9216) );
  NAND2_X1 U11774 ( .A1(n15011), .A2(n9324), .ZN(n9215) );
  NAND2_X1 U11775 ( .A1(n9216), .A2(n9215), .ZN(n14275) );
  NAND2_X1 U11776 ( .A1(n7968), .A2(n9217), .ZN(n9222) );
  INV_X1 U11777 ( .A(n14275), .ZN(n9218) );
  NAND2_X1 U11778 ( .A1(n7968), .A2(n9218), .ZN(n9219) );
  NAND2_X1 U11779 ( .A1(n14188), .A2(n14187), .ZN(n14200) );
  OAI21_X1 U11780 ( .B1(n9219), .B2(n14190), .A(n14200), .ZN(n9220) );
  XNOR2_X1 U11781 ( .A(n9224), .B(n9223), .ZN(n14201) );
  NAND2_X1 U11782 ( .A1(n10924), .A2(n8962), .ZN(n9230) );
  NAND2_X1 U11783 ( .A1(n9226), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9227) );
  MUX2_X1 U11784 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9227), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n9228) );
  AND2_X1 U11785 ( .A1(n9228), .A2(n6496), .ZN(n14718) );
  AOI22_X1 U11786 ( .A1(n9243), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10243), 
        .B2(n14718), .ZN(n9229) );
  NAND2_X1 U11787 ( .A1(n15109), .A2(n9387), .ZN(n9238) );
  INV_X1 U11788 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9236) );
  NAND2_X1 U11789 ( .A1(n9232), .A2(n7276), .ZN(n9233) );
  NAND2_X1 U11790 ( .A1(n9246), .A2(n9233), .ZN(n14935) );
  OR2_X1 U11791 ( .A1(n14935), .A2(n6438), .ZN(n9235) );
  AOI22_X1 U11792 ( .A1(n9314), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n14427), 
        .B2(P1_REG2_REG_18__SCAN_IN), .ZN(n9234) );
  OAI211_X1 U11793 ( .C1(n14432), .C2(n9236), .A(n9235), .B(n9234), .ZN(n14956) );
  NAND2_X1 U11794 ( .A1(n14956), .A2(n9397), .ZN(n9237) );
  NAND2_X1 U11795 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  XNOR2_X1 U11796 ( .A(n9239), .B(n9380), .ZN(n9240) );
  AOI22_X1 U11797 ( .A1(n15109), .A2(n9397), .B1(n9324), .B2(n14956), .ZN(
        n9241) );
  XNOR2_X1 U11798 ( .A(n9240), .B(n9241), .ZN(n14251) );
  INV_X1 U11799 ( .A(n9240), .ZN(n9242) );
  NAND2_X1 U11800 ( .A1(n11214), .A2(n8962), .ZN(n9245) );
  AOI22_X1 U11801 ( .A1(n9243), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14738), 
        .B2(n10243), .ZN(n9244) );
  NAND2_X2 U11802 ( .A1(n9245), .A2(n9244), .ZN(n15104) );
  INV_X1 U11803 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14726) );
  NAND2_X1 U11804 ( .A1(n9246), .A2(n7277), .ZN(n9247) );
  NAND2_X1 U11805 ( .A1(n9257), .A2(n9247), .ZN(n14917) );
  OR2_X1 U11806 ( .A1(n14917), .A2(n6438), .ZN(n9249) );
  AOI22_X1 U11807 ( .A1(n9408), .A2(P1_REG0_REG_19__SCAN_IN), .B1(n14427), 
        .B2(P1_REG2_REG_19__SCAN_IN), .ZN(n9248) );
  OAI211_X1 U11808 ( .C1(n14432), .C2(n14726), .A(n9249), .B(n9248), .ZN(
        n14929) );
  AOI22_X1 U11809 ( .A1(n15104), .A2(n9397), .B1(n9324), .B2(n14929), .ZN(
        n9252) );
  AOI22_X1 U11810 ( .A1(n15104), .A2(n9387), .B1(n9397), .B2(n14929), .ZN(
        n9250) );
  XNOR2_X1 U11811 ( .A(n9250), .B(n9380), .ZN(n9251) );
  XOR2_X1 U11812 ( .A(n9252), .B(n9251), .Z(n14153) );
  INV_X1 U11813 ( .A(n9251), .ZN(n9254) );
  NAND2_X1 U11814 ( .A1(n11454), .A2(n8962), .ZN(n9256) );
  INV_X1 U11815 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11455) );
  OR2_X1 U11816 ( .A1(n14476), .A2(n11455), .ZN(n9255) );
  NAND2_X2 U11817 ( .A1(n9256), .A2(n9255), .ZN(n15096) );
  INV_X1 U11818 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U11819 ( .A1(n9257), .A2(n14225), .ZN(n9258) );
  NAND2_X1 U11820 ( .A1(n9274), .A2(n9258), .ZN(n14899) );
  OR2_X1 U11821 ( .A1(n14899), .A2(n6439), .ZN(n9263) );
  INV_X1 U11822 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n15720) );
  NAND2_X1 U11823 ( .A1(n9314), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n9260) );
  NAND2_X1 U11824 ( .A1(n14427), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n9259) );
  OAI211_X1 U11825 ( .C1(n15720), .C2(n14432), .A(n9260), .B(n9259), .ZN(n9261) );
  INV_X1 U11826 ( .A(n9261), .ZN(n9262) );
  NAND2_X1 U11827 ( .A1(n9263), .A2(n9262), .ZN(n14545) );
  AND2_X1 U11828 ( .A1(n14545), .A2(n9395), .ZN(n9264) );
  AOI21_X1 U11829 ( .B1(n15096), .B2(n9397), .A(n9264), .ZN(n9267) );
  AOI22_X1 U11830 ( .A1(n15096), .A2(n9387), .B1(n9397), .B2(n14545), .ZN(
        n9265) );
  XNOR2_X1 U11831 ( .A(n9265), .B(n9380), .ZN(n9266) );
  XOR2_X1 U11832 ( .A(n9267), .B(n9266), .Z(n14222) );
  NAND2_X1 U11833 ( .A1(n9269), .A2(n9268), .ZN(n9270) );
  NAND2_X1 U11834 ( .A1(n11493), .A2(n8962), .ZN(n9272) );
  OR2_X1 U11835 ( .A1(n14476), .A2(n11495), .ZN(n9271) );
  INV_X1 U11836 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9273) );
  NAND2_X1 U11837 ( .A1(n9274), .A2(n9273), .ZN(n9275) );
  AND2_X1 U11838 ( .A1(n9293), .A2(n9275), .ZN(n14890) );
  NAND2_X1 U11839 ( .A1(n14890), .A2(n9388), .ZN(n9281) );
  INV_X1 U11840 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9278) );
  NAND2_X1 U11841 ( .A1(n8925), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n9277) );
  NAND2_X1 U11842 ( .A1(n9314), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n9276) );
  OAI211_X1 U11843 ( .C1(n14432), .C2(n9278), .A(n9277), .B(n9276), .ZN(n9279)
         );
  INV_X1 U11844 ( .A(n9279), .ZN(n9280) );
  AOI22_X1 U11845 ( .A1(n14891), .A2(n9397), .B1(n9395), .B2(n14544), .ZN(
        n9285) );
  NAND2_X1 U11846 ( .A1(n14891), .A2(n9387), .ZN(n9283) );
  NAND2_X1 U11847 ( .A1(n14544), .A2(n9397), .ZN(n9282) );
  NAND2_X1 U11848 ( .A1(n9283), .A2(n9282), .ZN(n9284) );
  XNOR2_X1 U11849 ( .A(n9284), .B(n9380), .ZN(n9287) );
  XOR2_X1 U11850 ( .A(n9285), .B(n9287), .Z(n14160) );
  INV_X1 U11851 ( .A(n9285), .ZN(n9286) );
  OR2_X1 U11852 ( .A1(n9287), .A2(n9286), .ZN(n9288) );
  NAND2_X1 U11853 ( .A1(n9289), .A2(n8209), .ZN(n9290) );
  INV_X1 U11854 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14247) );
  NAND2_X1 U11855 ( .A1(n9293), .A2(n14247), .ZN(n9294) );
  NAND2_X1 U11856 ( .A1(n9312), .A2(n9294), .ZN(n14873) );
  INV_X1 U11857 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n9297) );
  NAND2_X1 U11858 ( .A1(n8925), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n9296) );
  NAND2_X1 U11859 ( .A1(n9314), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n9295) );
  OAI211_X1 U11860 ( .C1(n14432), .C2(n9297), .A(n9296), .B(n9295), .ZN(n9298)
         );
  INV_X1 U11861 ( .A(n9298), .ZN(n9299) );
  OAI22_X1 U11862 ( .A1(n14877), .A2(n9301), .B1(n14852), .B2(n6494), .ZN(
        n9302) );
  XNOR2_X1 U11863 ( .A(n9302), .B(n9380), .ZN(n9304) );
  AND2_X1 U11864 ( .A1(n14543), .A2(n9324), .ZN(n9303) );
  AOI21_X1 U11865 ( .B1(n15084), .B2(n9397), .A(n9303), .ZN(n9305) );
  XNOR2_X1 U11866 ( .A(n9304), .B(n9305), .ZN(n14243) );
  INV_X1 U11867 ( .A(n9304), .ZN(n9306) );
  NAND2_X1 U11868 ( .A1(n14241), .A2(n9307), .ZN(n14132) );
  NAND2_X1 U11869 ( .A1(n11448), .A2(n8962), .ZN(n9309) );
  OR2_X1 U11870 ( .A1(n14476), .A2(n9897), .ZN(n9308) );
  NAND2_X1 U11871 ( .A1(n15078), .A2(n9401), .ZN(n9322) );
  INV_X1 U11872 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9311) );
  NAND2_X1 U11873 ( .A1(n9312), .A2(n9311), .ZN(n9313) );
  NAND2_X1 U11874 ( .A1(n9333), .A2(n9313), .ZN(n14134) );
  INV_X1 U11875 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9317) );
  NAND2_X1 U11876 ( .A1(n9314), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n9316) );
  NAND2_X1 U11877 ( .A1(n8925), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n9315) );
  OAI211_X1 U11878 ( .C1(n9317), .C2(n14432), .A(n9316), .B(n9315), .ZN(n9318)
         );
  INV_X1 U11879 ( .A(n9318), .ZN(n9319) );
  NAND2_X1 U11880 ( .A1(n14832), .A2(n9397), .ZN(n9321) );
  NAND2_X1 U11881 ( .A1(n9322), .A2(n9321), .ZN(n9323) );
  XNOR2_X1 U11882 ( .A(n9323), .B(n9380), .ZN(n9327) );
  AOI22_X1 U11883 ( .A1(n15078), .A2(n9397), .B1(n9324), .B2(n14832), .ZN(
        n9325) );
  XNOR2_X1 U11884 ( .A(n9327), .B(n9325), .ZN(n14133) );
  NAND2_X1 U11885 ( .A1(n14132), .A2(n14133), .ZN(n9329) );
  INV_X1 U11886 ( .A(n9325), .ZN(n9326) );
  NAND2_X1 U11887 ( .A1(n9329), .A2(n9328), .ZN(n14212) );
  INV_X1 U11888 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11566) );
  OR2_X1 U11889 ( .A1(n14476), .A2(n11566), .ZN(n9330) );
  NAND2_X1 U11890 ( .A1(n14840), .A2(n9387), .ZN(n9342) );
  INV_X1 U11891 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9332) );
  NAND2_X1 U11892 ( .A1(n9333), .A2(n9332), .ZN(n9334) );
  NAND2_X1 U11893 ( .A1(n14841), .A2(n9388), .ZN(n9340) );
  INV_X1 U11894 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9337) );
  NAND2_X1 U11895 ( .A1(n9408), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n9336) );
  NAND2_X1 U11896 ( .A1(n8925), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n9335) );
  OAI211_X1 U11897 ( .C1(n9337), .C2(n14432), .A(n9336), .B(n9335), .ZN(n9338)
         );
  INV_X1 U11898 ( .A(n9338), .ZN(n9339) );
  NAND2_X1 U11899 ( .A1(n14542), .A2(n9397), .ZN(n9341) );
  NAND2_X1 U11900 ( .A1(n9342), .A2(n9341), .ZN(n9343) );
  XNOR2_X1 U11901 ( .A(n9343), .B(n9380), .ZN(n9344) );
  AOI22_X1 U11902 ( .A1(n14840), .A2(n9397), .B1(n9395), .B2(n14542), .ZN(
        n9345) );
  XNOR2_X1 U11903 ( .A(n9344), .B(n9345), .ZN(n14213) );
  NAND2_X1 U11904 ( .A1(n14212), .A2(n14213), .ZN(n9348) );
  INV_X1 U11905 ( .A(n9344), .ZN(n9346) );
  NAND2_X1 U11906 ( .A1(n9346), .A2(n9345), .ZN(n9347) );
  NAND2_X1 U11907 ( .A1(n11488), .A2(n8962), .ZN(n9350) );
  OR2_X1 U11908 ( .A1(n14476), .A2(n15767), .ZN(n9349) );
  NAND2_X1 U11909 ( .A1(n15065), .A2(n9387), .ZN(n9361) );
  INV_X1 U11910 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9351) );
  NAND2_X1 U11911 ( .A1(n9352), .A2(n9351), .ZN(n9353) );
  NAND2_X1 U11912 ( .A1(n9370), .A2(n9353), .ZN(n14181) );
  INV_X1 U11913 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U11914 ( .A1(n9408), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n9355) );
  NAND2_X1 U11915 ( .A1(n14427), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n9354) );
  OAI211_X1 U11916 ( .C1(n9356), .C2(n14432), .A(n9355), .B(n9354), .ZN(n9357)
         );
  INV_X1 U11917 ( .A(n9357), .ZN(n9358) );
  NAND2_X1 U11918 ( .A1(n14833), .A2(n9397), .ZN(n9360) );
  NAND2_X1 U11919 ( .A1(n9361), .A2(n9360), .ZN(n9362) );
  XNOR2_X1 U11920 ( .A(n9362), .B(n9380), .ZN(n9363) );
  AOI22_X1 U11921 ( .A1(n15065), .A2(n9397), .B1(n9395), .B2(n14833), .ZN(
        n9364) );
  XNOR2_X1 U11922 ( .A(n9363), .B(n9364), .ZN(n14179) );
  INV_X1 U11923 ( .A(n9363), .ZN(n9365) );
  NAND2_X1 U11924 ( .A1(n9365), .A2(n9364), .ZN(n9366) );
  NAND2_X1 U11925 ( .A1(n11620), .A2(n8962), .ZN(n9368) );
  OR2_X1 U11926 ( .A1(n14476), .A2(n11621), .ZN(n9367) );
  NAND2_X1 U11927 ( .A1(n15060), .A2(n9387), .ZN(n9379) );
  INV_X1 U11928 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9369) );
  NAND2_X1 U11929 ( .A1(n9370), .A2(n9369), .ZN(n9371) );
  NAND2_X1 U11930 ( .A1(n14263), .A2(n9388), .ZN(n9377) );
  INV_X1 U11931 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9374) );
  NAND2_X1 U11932 ( .A1(n9408), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U11933 ( .A1(n8925), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n9372) );
  OAI211_X1 U11934 ( .C1(n9374), .C2(n14432), .A(n9373), .B(n9372), .ZN(n9375)
         );
  INV_X1 U11935 ( .A(n9375), .ZN(n9376) );
  NAND2_X1 U11936 ( .A1(n14753), .A2(n9397), .ZN(n9378) );
  NAND2_X1 U11937 ( .A1(n9379), .A2(n9378), .ZN(n9381) );
  XNOR2_X1 U11938 ( .A(n9381), .B(n9380), .ZN(n9382) );
  AOI22_X1 U11939 ( .A1(n15060), .A2(n9397), .B1(n9395), .B2(n14753), .ZN(
        n9383) );
  XNOR2_X1 U11940 ( .A(n9382), .B(n9383), .ZN(n14261) );
  INV_X1 U11941 ( .A(n9382), .ZN(n9384) );
  NAND2_X1 U11942 ( .A1(n11806), .A2(n8962), .ZN(n9386) );
  OR2_X1 U11943 ( .A1(n14476), .A2(n11807), .ZN(n9385) );
  NAND2_X1 U11944 ( .A1(n14806), .A2(n9387), .ZN(n9393) );
  XNOR2_X1 U11945 ( .A(n9404), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n14805) );
  INV_X1 U11946 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n15056) );
  NAND2_X1 U11947 ( .A1(n8925), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n9390) );
  NAND2_X1 U11948 ( .A1(n9408), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n9389) );
  OAI211_X1 U11949 ( .C1(n15056), .C2(n14432), .A(n9390), .B(n9389), .ZN(n9391) );
  NAND2_X1 U11950 ( .A1(n7796), .A2(n9397), .ZN(n9392) );
  NAND2_X1 U11951 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  XNOR2_X1 U11952 ( .A(n9394), .B(n10810), .ZN(n9423) );
  AND2_X1 U11953 ( .A1(n7796), .A2(n9395), .ZN(n9396) );
  AOI21_X1 U11954 ( .B1(n14806), .B2(n9397), .A(n9396), .ZN(n9422) );
  XNOR2_X1 U11955 ( .A(n9423), .B(n9422), .ZN(n14115) );
  INV_X1 U11956 ( .A(n14115), .ZN(n9398) );
  NAND2_X1 U11957 ( .A1(n14116), .A2(n9398), .ZN(n9448) );
  NAND2_X1 U11958 ( .A1(n11861), .A2(n8962), .ZN(n9400) );
  OR2_X1 U11959 ( .A1(n14476), .A2(n15196), .ZN(n9399) );
  NAND2_X1 U11960 ( .A1(n14787), .A2(n9401), .ZN(n9416) );
  INV_X1 U11961 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9403) );
  INV_X1 U11962 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n9402) );
  OAI21_X1 U11963 ( .B1(n9404), .B2(n9403), .A(n9402), .ZN(n9407) );
  INV_X1 U11964 ( .A(n9404), .ZN(n9406) );
  AND2_X1 U11965 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n9405) );
  NAND2_X1 U11966 ( .A1(n9406), .A2(n9405), .ZN(n14768) );
  NAND2_X1 U11967 ( .A1(n9407), .A2(n14768), .ZN(n9465) );
  INV_X1 U11968 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n9411) );
  NAND2_X1 U11969 ( .A1(n8925), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U11970 ( .A1(n9408), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n9409) );
  OAI211_X1 U11971 ( .C1(n9411), .C2(n14432), .A(n9410), .B(n9409), .ZN(n9412)
         );
  INV_X1 U11972 ( .A(n9412), .ZN(n9413) );
  NAND2_X1 U11973 ( .A1(n14761), .A2(n9397), .ZN(n9415) );
  NAND2_X1 U11974 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  XNOR2_X1 U11975 ( .A(n9417), .B(n10810), .ZN(n9421) );
  NOR2_X1 U11976 ( .A1(n14794), .A2(n9418), .ZN(n9419) );
  AOI21_X1 U11977 ( .B1(n14787), .B2(n9397), .A(n9419), .ZN(n9420) );
  XNOR2_X1 U11978 ( .A(n9421), .B(n9420), .ZN(n9471) );
  NAND2_X1 U11979 ( .A1(n9423), .A2(n9422), .ZN(n9470) );
  INV_X1 U11980 ( .A(n9430), .ZN(n11489) );
  NAND3_X1 U11981 ( .A1(n11489), .A2(P1_B_REG_SCAN_IN), .A3(n11564), .ZN(n9427) );
  INV_X1 U11982 ( .A(P1_B_REG_SCAN_IN), .ZN(n9424) );
  NAND2_X1 U11983 ( .A1(n9425), .A2(n9424), .ZN(n9426) );
  INV_X1 U11984 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U11985 ( .A1(n9439), .A2(n10186), .ZN(n9429) );
  INV_X1 U11986 ( .A(n10182), .ZN(n11622) );
  NAND2_X1 U11987 ( .A1(n11622), .A2(n11564), .ZN(n9428) );
  INV_X1 U11988 ( .A(n11462), .ZN(n15031) );
  OAI22_X1 U11989 ( .A1(n10184), .A2(P1_D_REG_1__SCAN_IN), .B1(n10182), .B2(
        n9430), .ZN(n15029) );
  INV_X1 U11990 ( .A(n15029), .ZN(n9442) );
  NOR4_X1 U11991 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9434) );
  NOR4_X1 U11992 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9433) );
  NOR4_X1 U11993 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9432) );
  NOR4_X1 U11994 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9431) );
  NAND4_X1 U11995 ( .A1(n9434), .A2(n9433), .A3(n9432), .A4(n9431), .ZN(n9441)
         );
  NOR2_X1 U11996 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n9438) );
  NOR4_X1 U11997 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n9437) );
  NOR4_X1 U11998 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9436) );
  NOR4_X1 U11999 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n9435) );
  NAND4_X1 U12000 ( .A1(n9438), .A2(n9437), .A3(n9436), .A4(n9435), .ZN(n9440)
         );
  OAI21_X1 U12001 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9464) );
  NAND3_X1 U12002 ( .A1(n15031), .A2(n9442), .A3(n9464), .ZN(n9451) );
  NAND2_X1 U12003 ( .A1(n9443), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9445) );
  INV_X1 U12004 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9444) );
  NAND2_X1 U12005 ( .A1(n14482), .A2(n14526), .ZN(n9463) );
  INV_X1 U12006 ( .A(n9463), .ZN(n9446) );
  INV_X1 U12007 ( .A(n10245), .ZN(n14481) );
  NAND3_X1 U12008 ( .A1(n10813), .A2(n15344), .A3(n14481), .ZN(n9447) );
  NAND4_X1 U12009 ( .A1(n9448), .A2(n9471), .A3(n9470), .A4(n14273), .ZN(n9475) );
  INV_X1 U12010 ( .A(n9448), .ZN(n9450) );
  INV_X1 U12011 ( .A(n9471), .ZN(n9449) );
  NAND2_X1 U12012 ( .A1(n9451), .A2(n15030), .ZN(n9468) );
  AND2_X1 U12013 ( .A1(n9468), .A2(n10813), .ZN(n14218) );
  NAND2_X1 U12014 ( .A1(n6645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9452) );
  XNOR2_X1 U12015 ( .A(n9452), .B(P1_IR_REG_28__SCAN_IN), .ZN(n14571) );
  NAND2_X1 U12016 ( .A1(n7796), .A2(n15008), .ZN(n9462) );
  OR2_X1 U12017 ( .A1(n14768), .A2(n6438), .ZN(n9460) );
  INV_X1 U12018 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n9457) );
  NAND2_X1 U12019 ( .A1(n8925), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n9456) );
  INV_X1 U12020 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n9454) );
  OR2_X1 U12021 ( .A1(n9079), .A2(n9454), .ZN(n9455) );
  OAI211_X1 U12022 ( .C1(n14432), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9458)
         );
  INV_X1 U12023 ( .A(n9458), .ZN(n9459) );
  NAND2_X1 U12024 ( .A1(n9460), .A2(n9459), .ZN(n14541) );
  INV_X1 U12025 ( .A(n14571), .ZN(n15193) );
  NAND2_X1 U12026 ( .A1(n14541), .A2(n15010), .ZN(n9461) );
  AND2_X1 U12027 ( .A1(n9462), .A2(n9461), .ZN(n15044) );
  NAND2_X1 U12028 ( .A1(n10245), .A2(n9463), .ZN(n9467) );
  NAND3_X1 U12029 ( .A1(n10813), .A2(n9467), .A3(n9464), .ZN(n15033) );
  OR2_X1 U12030 ( .A1(n15033), .A2(n15029), .ZN(n10811) );
  NOR2_X2 U12031 ( .A1(n10811), .A2(n11462), .ZN(n14282) );
  INV_X1 U12032 ( .A(n14282), .ZN(n14183) );
  INV_X1 U12033 ( .A(n9465), .ZN(n14784) );
  AND2_X1 U12034 ( .A1(n10244), .A2(n10106), .ZN(n9466) );
  AND2_X1 U12035 ( .A1(n9467), .A2(n9466), .ZN(n14536) );
  NAND2_X1 U12036 ( .A1(n9468), .A2(n14536), .ZN(n10293) );
  AOI22_X1 U12037 ( .A1(n14784), .A2(n14262), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9469) );
  OAI21_X1 U12038 ( .B1(n15044), .B2(n14183), .A(n9469), .ZN(n9473) );
  NOR3_X1 U12039 ( .A1(n9471), .A2(n14271), .A3(n9470), .ZN(n9472) );
  AOI211_X1 U12040 ( .C1(n14269), .C2(n14787), .A(n9473), .B(n9472), .ZN(n9474) );
  NAND2_X1 U12041 ( .A1(n9487), .A2(n9486), .ZN(n9488) );
  INV_X1 U12042 ( .A(n9501), .ZN(n9490) );
  NAND2_X1 U12043 ( .A1(n9491), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9492) );
  XNOR2_X1 U12044 ( .A(n9525), .B(n9523), .ZN(n10144) );
  NAND2_X1 U12045 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n9495) );
  OAI22_X1 U12046 ( .A1(n9522), .A2(n10144), .B1(n9529), .B2(n10528), .ZN(
        n9498) );
  NAND2_X4 U12047 ( .A1(n6448), .A2(n7875), .ZN(n9989) );
  INV_X1 U12048 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n9503) );
  INV_X1 U12049 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n10595) );
  INV_X1 U12050 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10382) );
  NAND2_X1 U12051 ( .A1(n9577), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n9508) );
  INV_X1 U12052 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10127) );
  OR2_X1 U12053 ( .A1(n10015), .A2(n10127), .ZN(n9507) );
  OR2_X1 U12054 ( .A1(n9846), .A2(n7410), .ZN(n9506) );
  INV_X1 U12055 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10553) );
  OR2_X1 U12056 ( .A1(n9591), .A2(n10553), .ZN(n9505) );
  NAND2_X1 U12057 ( .A1(n9509), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n9510) );
  AND2_X1 U12058 ( .A1(n9523), .A2(n9510), .ZN(n9512) );
  NAND2_X1 U12059 ( .A1(n10589), .A2(n10737), .ZN(n9515) );
  INV_X1 U12060 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9516) );
  INV_X1 U12061 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10400) );
  OR2_X1 U12062 ( .A1(n9846), .A2(n10400), .ZN(n9520) );
  INV_X1 U12063 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n9517) );
  OR2_X1 U12064 ( .A1(n9596), .A2(n9517), .ZN(n9519) );
  INV_X1 U12065 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n15609) );
  OR2_X1 U12066 ( .A1(n9591), .A2(n15609), .ZN(n9518) );
  INV_X1 U12067 ( .A(n9523), .ZN(n9524) );
  NAND2_X1 U12068 ( .A1(n9525), .A2(n9524), .ZN(n9527) );
  NAND2_X1 U12069 ( .A1(n10153), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9526) );
  NAND2_X1 U12070 ( .A1(n9527), .A2(n9526), .ZN(n9542) );
  XNOR2_X1 U12071 ( .A(n10152), .B(P2_DATAO_REG_2__SCAN_IN), .ZN(n9528) );
  XNOR2_X1 U12072 ( .A(n9542), .B(n9528), .ZN(n10151) );
  NAND2_X1 U12073 ( .A1(n9617), .A2(n10151), .ZN(n9532) );
  NAND2_X1 U12074 ( .A1(n9804), .A2(n10634), .ZN(n9531) );
  NOR2_X1 U12075 ( .A1(n12583), .A2(n7169), .ZN(n9534) );
  NAND2_X1 U12076 ( .A1(n6442), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9541) );
  INV_X1 U12077 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10686) );
  NAND2_X1 U12078 ( .A1(n9562), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n9537) );
  AND2_X1 U12079 ( .A1(n9626), .A2(n9537), .ZN(n11001) );
  OR2_X1 U12080 ( .A1(n9591), .A2(n11001), .ZN(n9539) );
  INV_X2 U12081 ( .A(n9596), .ZN(n9577) );
  INV_X1 U12082 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n9538) );
  INV_X1 U12083 ( .A(n9542), .ZN(n9544) );
  NAND2_X1 U12084 ( .A1(n10152), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9543) );
  NAND2_X1 U12085 ( .A1(n9544), .A2(n9543), .ZN(n9546) );
  NAND2_X1 U12086 ( .A1(n10157), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U12087 ( .A1(n10161), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n9549) );
  NAND2_X1 U12088 ( .A1(n9550), .A2(n9549), .ZN(n9583) );
  NAND2_X1 U12089 ( .A1(n10177), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n9551) );
  XNOR2_X1 U12090 ( .A(n15751), .B(P1_DATAO_REG_6__SCAN_IN), .ZN(n9611) );
  XNOR2_X1 U12091 ( .A(n9612), .B(n9611), .ZN(n10154) );
  NAND2_X1 U12092 ( .A1(n10154), .A2(n9617), .ZN(n9559) );
  INV_X1 U12093 ( .A(SI_6_), .ZN(n10156) );
  INV_X1 U12094 ( .A(n9601), .ZN(n9554) );
  INV_X1 U12095 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n9553) );
  NAND2_X1 U12096 ( .A1(n9554), .A2(n9553), .ZN(n9588) );
  NAND2_X1 U12097 ( .A1(n9618), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9556) );
  OAI22_X1 U12098 ( .A1(n9989), .A2(n10156), .B1(n9529), .B2(n15550), .ZN(
        n9557) );
  INV_X1 U12099 ( .A(n9557), .ZN(n9558) );
  NAND2_X2 U12100 ( .A1(n12425), .A2(n12427), .ZN(n12529) );
  NAND2_X1 U12101 ( .A1(n6442), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n9567) );
  INV_X1 U12102 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9560) );
  NAND2_X1 U12103 ( .A1(n9576), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n9561) );
  AND2_X1 U12104 ( .A1(n9562), .A2(n9561), .ZN(n10986) );
  OR2_X1 U12105 ( .A1(n9591), .A2(n10986), .ZN(n9565) );
  INV_X2 U12106 ( .A(n9577), .ZN(n12363) );
  INV_X1 U12107 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n9563) );
  OAI21_X1 U12108 ( .B1(n9570), .B2(n9569), .A(n9568), .ZN(n10148) );
  NAND2_X1 U12109 ( .A1(n9617), .A2(n10148), .ZN(n9574) );
  NAND2_X1 U12110 ( .A1(n9588), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9571) );
  MUX2_X1 U12111 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9571), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n9572) );
  NAND2_X1 U12112 ( .A1(n9572), .A2(n9618), .ZN(n10682) );
  NAND2_X1 U12113 ( .A1(n9804), .A2(n10682), .ZN(n9573) );
  INV_X1 U12114 ( .A(n10985), .ZN(n10805) );
  NAND2_X1 U12115 ( .A1(n10012), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U12116 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n9575) );
  AND2_X1 U12117 ( .A1(n9576), .A2(n9575), .ZN(n10774) );
  OR2_X1 U12118 ( .A1(n9591), .A2(n10774), .ZN(n9580) );
  INV_X1 U12119 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n9578) );
  NAND2_X1 U12120 ( .A1(n9584), .A2(n9583), .ZN(n9585) );
  NAND2_X1 U12121 ( .A1(n9586), .A2(n9585), .ZN(n10145) );
  NAND2_X1 U12122 ( .A1(n9601), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9587) );
  MUX2_X1 U12123 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9587), .S(
        P3_IR_REG_4__SCAN_IN), .Z(n9589) );
  NAND2_X1 U12124 ( .A1(n9589), .A2(n9588), .ZN(n10443) );
  NAND2_X1 U12125 ( .A1(n9804), .A2(n10443), .ZN(n9590) );
  NAND2_X1 U12126 ( .A1(n12582), .A2(n15627), .ZN(n12422) );
  INV_X1 U12127 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n10390) );
  OR2_X1 U12128 ( .A1(n9591), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9593) );
  NAND2_X1 U12129 ( .A1(n6441), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n9592) );
  INV_X1 U12130 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n9595) );
  XNOR2_X1 U12131 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n9598) );
  XNOR2_X1 U12132 ( .A(n9599), .B(n9598), .ZN(n10146) );
  NAND2_X1 U12133 ( .A1(n9637), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9600) );
  MUX2_X1 U12134 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9600), .S(
        P3_IR_REG_3__SCAN_IN), .Z(n9602) );
  NAND2_X1 U12135 ( .A1(n9804), .A2(n10680), .ZN(n9603) );
  NAND2_X1 U12136 ( .A1(n12980), .A2(n10789), .ZN(n12413) );
  AND2_X2 U12137 ( .A1(n12408), .A2(n12413), .ZN(n10783) );
  AND2_X1 U12138 ( .A1(n12980), .A2(n9604), .ZN(n10768) );
  NAND2_X1 U12139 ( .A1(n12582), .A2(n7130), .ZN(n9605) );
  NAND2_X1 U12140 ( .A1(n9606), .A2(n9605), .ZN(n10962) );
  OR2_X1 U12141 ( .A1(n12581), .A2(n10985), .ZN(n12424) );
  NAND2_X1 U12142 ( .A1(n12581), .A2(n10985), .ZN(n12419) );
  NAND2_X1 U12143 ( .A1(n10199), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U12144 ( .A1(n9634), .A2(n9613), .ZN(n9614) );
  NAND2_X1 U12145 ( .A1(n9615), .A2(n9614), .ZN(n9616) );
  NAND2_X1 U12146 ( .A1(n9635), .A2(n9616), .ZN(n10158) );
  NAND2_X1 U12147 ( .A1(n10158), .A2(n9956), .ZN(n9622) );
  OAI21_X1 U12148 ( .B1(n9618), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9619) );
  XNOR2_X1 U12149 ( .A(n9619), .B(P3_IR_REG_7__SCAN_IN), .ZN(n11228) );
  OAI22_X1 U12150 ( .A1(n9989), .A2(SI_7_), .B1(n11228), .B2(n9529), .ZN(n9620) );
  INV_X1 U12151 ( .A(n9620), .ZN(n9621) );
  NAND2_X1 U12152 ( .A1(n10012), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n9632) );
  INV_X1 U12153 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n9623) );
  NAND2_X1 U12154 ( .A1(n9626), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n9627) );
  AND2_X1 U12155 ( .A1(n9646), .A2(n9627), .ZN(n11069) );
  OR2_X1 U12156 ( .A1(n9591), .A2(n11069), .ZN(n9630) );
  INV_X1 U12157 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n9628) );
  OR2_X1 U12158 ( .A1(n6443), .A2(n9628), .ZN(n9629) );
  INV_X1 U12159 ( .A(n12579), .ZN(n10995) );
  OR2_X1 U12160 ( .A1(n10995), .A2(n11096), .ZN(n9633) );
  XNOR2_X1 U12161 ( .A(n10235), .B(P2_DATAO_REG_8__SCAN_IN), .ZN(n9636) );
  XNOR2_X1 U12162 ( .A(n9656), .B(n9636), .ZN(n10171) );
  NAND2_X1 U12163 ( .A1(n10171), .A2(n9956), .ZN(n9645) );
  INV_X1 U12164 ( .A(SI_8_), .ZN(n10173) );
  INV_X1 U12165 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U12166 ( .A1(n10000), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9641) );
  MUX2_X1 U12167 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9641), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n9642) );
  NAND2_X1 U12168 ( .A1(n9642), .A2(n9661), .ZN(n11239) );
  OAI22_X1 U12169 ( .A1(n9989), .A2(n10173), .B1(n9529), .B2(n11239), .ZN(
        n9643) );
  INV_X1 U12170 ( .A(n9643), .ZN(n9644) );
  NAND2_X1 U12171 ( .A1(n6442), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n9652) );
  INV_X1 U12172 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n11223) );
  OR2_X1 U12173 ( .A1(n6443), .A2(n11223), .ZN(n9651) );
  NAND2_X1 U12174 ( .A1(n9646), .A2(P3_REG3_REG_8__SCAN_IN), .ZN(n9647) );
  AND2_X1 U12175 ( .A1(n9669), .A2(n9647), .ZN(n11261) );
  OR2_X1 U12176 ( .A1(n9591), .A2(n11261), .ZN(n9650) );
  INV_X1 U12177 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n9648) );
  OR2_X1 U12178 ( .A1(n12363), .A2(n9648), .ZN(n9649) );
  NAND4_X1 U12179 ( .A1(n9652), .A2(n9651), .A3(n9650), .A4(n9649), .ZN(n12578) );
  OR2_X1 U12180 ( .A1(n12435), .A2(n12578), .ZN(n9653) );
  NAND2_X1 U12181 ( .A1(n12435), .A2(n12578), .ZN(n9654) );
  NAND2_X1 U12182 ( .A1(n10235), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U12183 ( .A1(n9656), .A2(n9655), .ZN(n9658) );
  NAND2_X1 U12184 ( .A1(n10238), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n9657) );
  XNOR2_X1 U12185 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n9659) );
  XNOR2_X1 U12186 ( .A(n9680), .B(n9659), .ZN(n10174) );
  NAND2_X1 U12187 ( .A1(n10174), .A2(n9956), .ZN(n9666) );
  NAND2_X1 U12188 ( .A1(n9661), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9660) );
  MUX2_X1 U12189 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9660), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n9663) );
  INV_X1 U12190 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n9662) );
  NAND2_X1 U12191 ( .A1(n9818), .A2(n9662), .ZN(n9698) );
  NAND2_X1 U12192 ( .A1(n9663), .A2(n9698), .ZN(n11694) );
  INV_X1 U12193 ( .A(n11694), .ZN(n11235) );
  OAI22_X1 U12194 ( .A1(n9989), .A2(SI_9_), .B1(n11235), .B2(n9529), .ZN(n9664) );
  INV_X1 U12195 ( .A(n9664), .ZN(n9665) );
  NAND2_X1 U12196 ( .A1(n9666), .A2(n9665), .ZN(n11272) );
  NAND2_X1 U12197 ( .A1(n10012), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n9675) );
  INV_X1 U12198 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n9667) );
  OR2_X1 U12199 ( .A1(n6443), .A2(n9667), .ZN(n9674) );
  NAND2_X1 U12200 ( .A1(n9669), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n9670) );
  AND2_X1 U12201 ( .A1(n9686), .A2(n9670), .ZN(n10875) );
  OR2_X1 U12202 ( .A1(n9591), .A2(n10875), .ZN(n9673) );
  INV_X1 U12203 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n9671) );
  OR2_X1 U12204 ( .A1(n12363), .A2(n9671), .ZN(n9672) );
  NAND4_X1 U12205 ( .A1(n9675), .A2(n9674), .A3(n9673), .A4(n9672), .ZN(n12577) );
  OR2_X1 U12206 ( .A1(n11272), .A2(n12577), .ZN(n12439) );
  NAND2_X1 U12207 ( .A1(n11266), .A2(n11267), .ZN(n9677) );
  INV_X1 U12208 ( .A(n12577), .ZN(n11294) );
  OR2_X1 U12209 ( .A1(n11272), .A2(n11294), .ZN(n9676) );
  NAND2_X1 U12210 ( .A1(n10240), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n9678) );
  NAND2_X1 U12211 ( .A1(n10286), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n9694) );
  NAND2_X1 U12212 ( .A1(n10289), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n9681) );
  NAND2_X1 U12213 ( .A1(n9694), .A2(n9681), .ZN(n9695) );
  XNOR2_X1 U12214 ( .A(n9696), .B(n9695), .ZN(n10192) );
  NAND2_X1 U12215 ( .A1(n10192), .A2(n9956), .ZN(n9685) );
  NAND2_X1 U12216 ( .A1(n9698), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9682) );
  XNOR2_X1 U12217 ( .A(n9682), .B(P3_IR_REG_10__SCAN_IN), .ZN(n15597) );
  OAI22_X1 U12218 ( .A1(n7167), .A2(SI_10_), .B1(n15597), .B2(n9529), .ZN(
        n9683) );
  INV_X1 U12219 ( .A(n9683), .ZN(n9684) );
  NAND2_X1 U12220 ( .A1(n9685), .A2(n9684), .ZN(n11390) );
  NAND2_X1 U12221 ( .A1(n12360), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n9692) );
  INV_X1 U12222 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n11691) );
  OR2_X1 U12223 ( .A1(n9846), .A2(n11691), .ZN(n9691) );
  NAND2_X1 U12224 ( .A1(n9686), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n9687) );
  AND2_X1 U12225 ( .A1(n9705), .A2(n9687), .ZN(n11392) );
  OR2_X1 U12226 ( .A1(n9591), .A2(n11392), .ZN(n9690) );
  INV_X1 U12227 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n9688) );
  OR2_X1 U12228 ( .A1(n12363), .A2(n9688), .ZN(n9689) );
  NAND4_X1 U12229 ( .A1(n9692), .A2(n9691), .A3(n9690), .A4(n9689), .ZN(n12576) );
  OR2_X1 U12230 ( .A1(n11390), .A2(n12576), .ZN(n12443) );
  NAND2_X1 U12231 ( .A1(n11390), .A2(n12576), .ZN(n12442) );
  INV_X1 U12232 ( .A(n12576), .ZN(n10913) );
  OR2_X1 U12233 ( .A1(n11390), .A2(n10913), .ZN(n9693) );
  XNOR2_X1 U12234 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n9697) );
  XNOR2_X1 U12235 ( .A(n9713), .B(n9697), .ZN(n10200) );
  NAND2_X1 U12236 ( .A1(n10200), .A2(n9956), .ZN(n9704) );
  INV_X1 U12237 ( .A(n9698), .ZN(n9700) );
  NAND2_X1 U12238 ( .A1(n9700), .A2(n9699), .ZN(n9714) );
  NAND2_X1 U12239 ( .A1(n9714), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9701) );
  XNOR2_X1 U12240 ( .A(n9701), .B(P3_IR_REG_11__SCAN_IN), .ZN(n12600) );
  OAI22_X1 U12241 ( .A1(n7167), .A2(SI_11_), .B1(n12600), .B2(n9529), .ZN(
        n9702) );
  INV_X1 U12242 ( .A(n9702), .ZN(n9703) );
  NAND2_X1 U12243 ( .A1(n9704), .A2(n9703), .ZN(n11499) );
  NAND2_X1 U12244 ( .A1(n9705), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n9706) );
  NAND2_X1 U12245 ( .A1(n9722), .A2(n9706), .ZN(n11503) );
  NAND2_X1 U12246 ( .A1(n9991), .A2(n11503), .ZN(n9711) );
  INV_X1 U12247 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n11496) );
  OR2_X1 U12248 ( .A1(n6443), .A2(n11496), .ZN(n9710) );
  INV_X1 U12249 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n11502) );
  OR2_X1 U12250 ( .A1(n9846), .A2(n11502), .ZN(n9709) );
  INV_X1 U12251 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n9707) );
  OR2_X1 U12252 ( .A1(n12363), .A2(n9707), .ZN(n9708) );
  NAND4_X1 U12253 ( .A1(n9711), .A2(n9710), .A3(n9709), .A4(n9708), .ZN(n12575) );
  INV_X1 U12254 ( .A(n12575), .ZN(n10919) );
  NOR2_X1 U12255 ( .A1(n11499), .A2(n10919), .ZN(n9712) );
  XNOR2_X1 U12256 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n9730) );
  XNOR2_X1 U12257 ( .A(n9731), .B(n9730), .ZN(n10232) );
  NAND2_X1 U12258 ( .A1(n10232), .A2(n9956), .ZN(n9721) );
  NAND2_X1 U12259 ( .A1(n9716), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9715) );
  MUX2_X1 U12260 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9715), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n9719) );
  INV_X1 U12261 ( .A(n9716), .ZN(n9718) );
  INV_X1 U12262 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n9717) );
  NAND2_X1 U12263 ( .A1(n9718), .A2(n9717), .ZN(n9734) );
  NAND2_X1 U12264 ( .A1(n9719), .A2(n9734), .ZN(n12612) );
  AOI22_X1 U12265 ( .A1(n12368), .A2(n10233), .B1(n12612), .B2(n9804), .ZN(
        n9720) );
  NAND2_X1 U12266 ( .A1(n9722), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U12267 ( .A1(n9743), .A2(n9723), .ZN(n11517) );
  NAND2_X1 U12268 ( .A1(n9991), .A2(n11517), .ZN(n9728) );
  INV_X1 U12269 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n12596) );
  OR2_X1 U12270 ( .A1(n6443), .A2(n12596), .ZN(n9727) );
  INV_X1 U12271 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n9724) );
  OR2_X1 U12272 ( .A1(n9846), .A2(n9724), .ZN(n9726) );
  INV_X1 U12273 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n11440) );
  OR2_X1 U12274 ( .A1(n12363), .A2(n11440), .ZN(n9725) );
  NAND4_X1 U12275 ( .A1(n9728), .A2(n9727), .A3(n9726), .A4(n9725), .ZN(n12574) );
  NAND2_X1 U12276 ( .A1(n11520), .A2(n12574), .ZN(n12455) );
  INV_X1 U12277 ( .A(n12574), .ZN(n11636) );
  OR2_X1 U12278 ( .A1(n11520), .A2(n11636), .ZN(n9729) );
  NAND2_X1 U12279 ( .A1(n9731), .A2(n9730), .ZN(n9733) );
  NAND2_X1 U12280 ( .A1(n15769), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n9732) );
  XNOR2_X1 U12281 ( .A(n9750), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U12282 ( .A1(n10282), .A2(n9956), .ZN(n9740) );
  NAND2_X1 U12283 ( .A1(n9734), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9735) );
  MUX2_X1 U12284 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9735), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n9737) );
  NAND2_X1 U12285 ( .A1(n9818), .A2(n9736), .ZN(n9769) );
  NAND2_X1 U12286 ( .A1(n9737), .A2(n9769), .ZN(n12637) );
  NOR2_X1 U12287 ( .A1(n7167), .A2(SI_13_), .ZN(n9738) );
  AOI21_X1 U12288 ( .B1(n12637), .B2(n9804), .A(n9738), .ZN(n9739) );
  NAND2_X1 U12289 ( .A1(n9743), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U12290 ( .A1(n9758), .A2(n9744), .ZN(n11647) );
  NAND2_X1 U12291 ( .A1(n11647), .A2(n9991), .ZN(n9748) );
  NAND2_X1 U12292 ( .A1(n10012), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n9747) );
  NAND2_X1 U12293 ( .A1(n12360), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n9746) );
  NAND2_X1 U12294 ( .A1(n9577), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n9745) );
  NAND4_X1 U12295 ( .A1(n9748), .A2(n9747), .A3(n9746), .A4(n9745), .ZN(n12573) );
  NAND2_X1 U12296 ( .A1(n11644), .A2(n12573), .ZN(n12457) );
  INV_X1 U12297 ( .A(n12536), .ZN(n11595) );
  NAND2_X1 U12298 ( .A1(n11596), .A2(n11595), .ZN(n11594) );
  INV_X1 U12299 ( .A(n12573), .ZN(n11674) );
  OR2_X1 U12300 ( .A1(n11644), .A2(n11674), .ZN(n9749) );
  NAND2_X1 U12301 ( .A1(n9750), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n9754) );
  NAND2_X1 U12302 ( .A1(n9752), .A2(n9751), .ZN(n9753) );
  XNOR2_X1 U12303 ( .A(n10767), .B(P2_DATAO_REG_14__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U12304 ( .A(n9766), .B(n9755), .ZN(n10495) );
  NAND2_X1 U12305 ( .A1(n9769), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9756) );
  XNOR2_X1 U12306 ( .A(n9770), .B(n9756), .ZN(n12641) );
  OAI22_X1 U12307 ( .A1(n7167), .A2(n10497), .B1(n9529), .B2(n12641), .ZN(
        n9757) );
  AOI21_X1 U12308 ( .B1(n10495), .B2(n9956), .A(n9757), .ZN(n11675) );
  INV_X1 U12309 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n11783) );
  NAND2_X1 U12310 ( .A1(n9758), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n9759) );
  NAND2_X1 U12311 ( .A1(n9775), .A2(n9759), .ZN(n11786) );
  NAND2_X1 U12312 ( .A1(n11786), .A2(n9991), .ZN(n9763) );
  NAND2_X1 U12313 ( .A1(n12360), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n9761) );
  NAND2_X1 U12314 ( .A1(n6442), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n9760) );
  AND2_X1 U12315 ( .A1(n9761), .A2(n9760), .ZN(n9762) );
  OAI211_X1 U12316 ( .C1(n12363), .C2(n11783), .A(n9763), .B(n9762), .ZN(
        n12572) );
  AND2_X1 U12317 ( .A1(n11675), .A2(n12572), .ZN(n10078) );
  INV_X1 U12318 ( .A(n10078), .ZN(n12462) );
  INV_X1 U12319 ( .A(n11675), .ZN(n11787) );
  INV_X1 U12320 ( .A(n12572), .ZN(n11676) );
  NAND2_X1 U12321 ( .A1(n11787), .A2(n11676), .ZN(n12463) );
  OR2_X1 U12322 ( .A1(n11675), .A2(n11676), .ZN(n9764) );
  NAND2_X1 U12323 ( .A1(n10767), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U12324 ( .A1(n10831), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n9782) );
  NAND2_X1 U12325 ( .A1(n10830), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n9768) );
  XNOR2_X1 U12326 ( .A(n9784), .B(n9781), .ZN(n10635) );
  NAND2_X1 U12327 ( .A1(n10635), .A2(n9956), .ZN(n9774) );
  INV_X1 U12328 ( .A(n9769), .ZN(n9771) );
  NAND2_X1 U12329 ( .A1(n9771), .A2(n9770), .ZN(n9786) );
  NAND2_X1 U12330 ( .A1(n9786), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9772) );
  XNOR2_X1 U12331 ( .A(n9772), .B(P3_IR_REG_15__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U12332 ( .A1(n12368), .A2(SI_15_), .B1(n9804), .B2(n12661), .ZN(
        n9773) );
  NAND2_X1 U12333 ( .A1(n9775), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n9776) );
  NAND2_X1 U12334 ( .A1(n9793), .A2(n9776), .ZN(n11832) );
  NAND2_X1 U12335 ( .A1(n11832), .A2(n9991), .ZN(n9779) );
  AOI22_X1 U12336 ( .A1(n6442), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12360), 
        .B2(P3_REG1_REG_15__SCAN_IN), .ZN(n9778) );
  NAND2_X1 U12337 ( .A1(n9577), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n9777) );
  OR2_X1 U12338 ( .A1(n11826), .A2(n11677), .ZN(n12466) );
  INV_X1 U12339 ( .A(n12538), .ZN(n11764) );
  NAND2_X1 U12340 ( .A1(n11826), .A2(n12918), .ZN(n9780) );
  INV_X1 U12341 ( .A(n9781), .ZN(n9783) );
  NAND2_X1 U12342 ( .A1(n10748), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n9800) );
  NAND2_X1 U12343 ( .A1(n10751), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n9785) );
  NAND2_X1 U12344 ( .A1(n9800), .A2(n9785), .ZN(n9798) );
  NAND2_X1 U12345 ( .A1(n9788), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9787) );
  MUX2_X1 U12346 ( .A(P3_IR_REG_31__SCAN_IN), .B(n9787), .S(
        P3_IR_REG_16__SCAN_IN), .Z(n9791) );
  INV_X1 U12347 ( .A(n9788), .ZN(n9790) );
  NAND2_X1 U12348 ( .A1(n9790), .A2(n9789), .ZN(n9802) );
  NAND2_X1 U12349 ( .A1(n9791), .A2(n9802), .ZN(n12701) );
  OAI22_X1 U12350 ( .A1(n12701), .A2(n9529), .B1(n7167), .B2(n10780), .ZN(
        n9792) );
  INV_X1 U12351 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n15696) );
  NAND2_X1 U12352 ( .A1(n9793), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n9794) );
  NAND2_X1 U12353 ( .A1(n9808), .A2(n9794), .ZN(n12911) );
  NAND2_X1 U12354 ( .A1(n12911), .A2(n9991), .ZN(n9796) );
  AOI22_X1 U12355 ( .A1(n6442), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n12360), 
        .B2(P3_REG1_REG_16__SCAN_IN), .ZN(n9795) );
  INV_X1 U12356 ( .A(n12905), .ZN(n12293) );
  NAND2_X1 U12357 ( .A1(n12286), .A2(n12293), .ZN(n9797) );
  XNOR2_X1 U12358 ( .A(n10900), .B(P2_DATAO_REG_17__SCAN_IN), .ZN(n9801) );
  XNOR2_X1 U12359 ( .A(n9815), .B(n9801), .ZN(n10926) );
  NAND2_X1 U12360 ( .A1(n10926), .A2(n9956), .ZN(n9806) );
  NAND2_X1 U12361 ( .A1(n9802), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9803) );
  XNOR2_X1 U12362 ( .A(n9803), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U12363 ( .A1(n12713), .A2(n9804), .B1(SI_17_), .B2(n12368), .ZN(
        n9805) );
  INV_X1 U12364 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n9807) );
  NAND2_X1 U12365 ( .A1(n9808), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n9809) );
  NAND2_X1 U12366 ( .A1(n9824), .A2(n9809), .ZN(n12901) );
  NAND2_X1 U12367 ( .A1(n12901), .A2(n9991), .ZN(n9814) );
  INV_X1 U12368 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n15723) );
  NAND2_X1 U12369 ( .A1(n9577), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n9811) );
  NAND2_X1 U12370 ( .A1(n10012), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n9810) );
  OAI211_X1 U12371 ( .C1(n6443), .C2(n15723), .A(n9811), .B(n9810), .ZN(n9812)
         );
  INV_X1 U12372 ( .A(n9812), .ZN(n9813) );
  OR2_X1 U12373 ( .A1(n13056), .A2(n12281), .ZN(n12392) );
  NAND2_X1 U12374 ( .A1(n13056), .A2(n12281), .ZN(n12394) );
  NAND2_X1 U12375 ( .A1(n12392), .A2(n12394), .ZN(n12539) );
  XNOR2_X1 U12376 ( .A(n9835), .B(P1_DATAO_REG_18__SCAN_IN), .ZN(n9832) );
  XNOR2_X1 U12377 ( .A(n9834), .B(n9832), .ZN(n11101) );
  NAND2_X1 U12378 ( .A1(n11101), .A2(n9956), .ZN(n9823) );
  NAND2_X1 U12379 ( .A1(n9839), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n9820) );
  XNOR2_X1 U12380 ( .A(n9820), .B(n9819), .ZN(n12746) );
  OAI22_X1 U12381 ( .A1(n7167), .A2(n11103), .B1(n9529), .B2(n12746), .ZN(
        n9821) );
  INV_X1 U12382 ( .A(n9821), .ZN(n9822) );
  NAND2_X1 U12383 ( .A1(n9824), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U12384 ( .A1(n9842), .A2(n9825), .ZN(n12892) );
  NAND2_X1 U12385 ( .A1(n12892), .A2(n9991), .ZN(n9830) );
  INV_X1 U12386 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n13049) );
  NAND2_X1 U12387 ( .A1(n12360), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n9827) );
  NAND2_X1 U12388 ( .A1(n6442), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n9826) );
  OAI211_X1 U12389 ( .C1(n13049), .C2(n12363), .A(n9827), .B(n9826), .ZN(n9828) );
  INV_X1 U12390 ( .A(n9828), .ZN(n9829) );
  NAND2_X1 U12391 ( .A1(n13050), .A2(n12328), .ZN(n12477) );
  NAND2_X1 U12392 ( .A1(n12390), .A2(n12477), .ZN(n12893) );
  OR2_X1 U12393 ( .A1(n13050), .A2(n12903), .ZN(n9831) );
  INV_X1 U12394 ( .A(n9832), .ZN(n9833) );
  NAND2_X1 U12395 ( .A1(n9834), .A2(n9833), .ZN(n9837) );
  NAND2_X1 U12396 ( .A1(n9835), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n9836) );
  INV_X1 U12397 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11217) );
  NAND2_X1 U12398 ( .A1(n11217), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n9852) );
  INV_X1 U12399 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11215) );
  NAND2_X1 U12400 ( .A1(n11215), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n9838) );
  XNOR2_X1 U12401 ( .A(n9853), .B(n9851), .ZN(n11165) );
  OAI21_X1 U12402 ( .B1(n9839), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n9840) );
  OAI22_X1 U12403 ( .A1(n7167), .A2(SI_19_), .B1(n12548), .B2(n9529), .ZN(
        n9841) );
  NAND2_X1 U12404 ( .A1(n9842), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n9843) );
  NAND2_X1 U12405 ( .A1(n9857), .A2(n9843), .ZN(n12884) );
  NAND2_X1 U12406 ( .A1(n12884), .A2(n9991), .ZN(n9849) );
  INV_X1 U12407 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n15693) );
  NAND2_X1 U12408 ( .A1(n9577), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n9845) );
  NAND2_X1 U12409 ( .A1(n12360), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n9844) );
  OAI211_X1 U12410 ( .C1(n9846), .C2(n15693), .A(n9845), .B(n9844), .ZN(n9847)
         );
  INV_X1 U12411 ( .A(n9847), .ZN(n9848) );
  NAND2_X1 U12412 ( .A1(n12249), .A2(n12333), .ZN(n12540) );
  INV_X1 U12413 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n11457) );
  NAND2_X1 U12414 ( .A1(n11457), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n9867) );
  NAND2_X1 U12415 ( .A1(n11455), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n9854) );
  XNOR2_X1 U12416 ( .A(n9866), .B(n9865), .ZN(n11333) );
  NAND2_X1 U12417 ( .A1(n11333), .A2(n9956), .ZN(n9856) );
  NAND2_X1 U12418 ( .A1(n12368), .A2(SI_20_), .ZN(n9855) );
  NAND2_X1 U12419 ( .A1(n9857), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n9858) );
  NAND2_X1 U12420 ( .A1(n9871), .A2(n9858), .ZN(n12874) );
  NAND2_X1 U12421 ( .A1(n12874), .A2(n9991), .ZN(n9863) );
  INV_X1 U12422 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13036) );
  NAND2_X1 U12423 ( .A1(n10012), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n9860) );
  NAND2_X1 U12424 ( .A1(n12360), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n9859) );
  OAI211_X1 U12425 ( .C1(n12363), .C2(n13036), .A(n9860), .B(n9859), .ZN(n9861) );
  INV_X1 U12426 ( .A(n9861), .ZN(n9862) );
  XNOR2_X1 U12427 ( .A(n13038), .B(n12887), .ZN(n12872) );
  INV_X1 U12428 ( .A(n12872), .ZN(n12876) );
  NAND2_X1 U12429 ( .A1(n13038), .A2(n12887), .ZN(n9864) );
  XNOR2_X1 U12430 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .ZN(n9879) );
  XNOR2_X1 U12431 ( .A(n9880), .B(n9879), .ZN(n11458) );
  NAND2_X1 U12432 ( .A1(n11458), .A2(n9956), .ZN(n9869) );
  NAND2_X1 U12433 ( .A1(n12368), .A2(SI_21_), .ZN(n9868) );
  INV_X1 U12434 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12435 ( .A1(n9871), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12436 ( .A1(n9885), .A2(n9872), .ZN(n12863) );
  NAND2_X1 U12437 ( .A1(n12863), .A2(n9991), .ZN(n9877) );
  INV_X1 U12438 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n15799) );
  NAND2_X1 U12439 ( .A1(n12360), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n9874) );
  NAND2_X1 U12440 ( .A1(n6442), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n9873) );
  OAI211_X1 U12441 ( .C1(n15799), .C2(n12363), .A(n9874), .B(n9873), .ZN(n9875) );
  INV_X1 U12442 ( .A(n9875), .ZN(n9876) );
  AND2_X1 U12443 ( .A1(n13032), .A2(n12570), .ZN(n9878) );
  INV_X1 U12444 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11951) );
  NAND2_X1 U12445 ( .A1(n11951), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n9893) );
  INV_X1 U12446 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9881) );
  NAND2_X1 U12447 ( .A1(n9881), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U12448 ( .A1(n9893), .A2(n9882), .ZN(n9894) );
  XNOR2_X1 U12449 ( .A(n9895), .B(n9894), .ZN(n11588) );
  NAND2_X1 U12450 ( .A1(n11588), .A2(n9956), .ZN(n9884) );
  NAND2_X1 U12451 ( .A1(n12368), .A2(SI_22_), .ZN(n9883) );
  NAND2_X1 U12452 ( .A1(n9885), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n9886) );
  NAND2_X1 U12453 ( .A1(n9903), .A2(n9886), .ZN(n12854) );
  NAND2_X1 U12454 ( .A1(n12854), .A2(n9991), .ZN(n9891) );
  INV_X1 U12455 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13026) );
  NAND2_X1 U12456 ( .A1(n6442), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n9888) );
  NAND2_X1 U12457 ( .A1(n12360), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n9887) );
  OAI211_X1 U12458 ( .C1(n13026), .C2(n12363), .A(n9888), .B(n9887), .ZN(n9889) );
  INV_X1 U12459 ( .A(n9889), .ZN(n9890) );
  OR2_X1 U12460 ( .A1(n13027), .A2(n12569), .ZN(n9892) );
  NAND2_X1 U12461 ( .A1(n9896), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n9912) );
  NAND2_X1 U12462 ( .A1(n9897), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n9898) );
  AND2_X1 U12463 ( .A1(n9912), .A2(n9898), .ZN(n9899) );
  OAI21_X1 U12464 ( .B1(n9900), .B2(n9899), .A(n9913), .ZN(n11743) );
  NAND2_X1 U12465 ( .A1(n11743), .A2(n9956), .ZN(n9902) );
  NAND2_X1 U12466 ( .A1(n12368), .A2(SI_23_), .ZN(n9901) );
  NAND2_X1 U12467 ( .A1(n9903), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n9904) );
  NAND2_X1 U12468 ( .A1(n6630), .A2(n9904), .ZN(n12846) );
  NAND2_X1 U12469 ( .A1(n12846), .A2(n9991), .ZN(n9910) );
  INV_X1 U12470 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n9907) );
  NAND2_X1 U12471 ( .A1(n6442), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n9906) );
  NAND2_X1 U12472 ( .A1(n12360), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n9905) );
  OAI211_X1 U12473 ( .C1(n12363), .C2(n9907), .A(n9906), .B(n9905), .ZN(n9908)
         );
  INV_X1 U12474 ( .A(n9908), .ZN(n9909) );
  NAND2_X1 U12475 ( .A1(n12944), .A2(n12821), .ZN(n9911) );
  XNOR2_X1 U12476 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .ZN(n9914) );
  XNOR2_X1 U12477 ( .A(n9925), .B(n9914), .ZN(n9915) );
  INV_X1 U12478 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15691) );
  NAND2_X1 U12479 ( .A1(n6630), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n9916) );
  NAND2_X1 U12480 ( .A1(n9929), .A2(n9916), .ZN(n12826) );
  NAND2_X1 U12481 ( .A1(n12826), .A2(n9991), .ZN(n9921) );
  INV_X1 U12482 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13018) );
  NAND2_X1 U12483 ( .A1(n6441), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U12484 ( .A1(n12360), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n9917) );
  OAI211_X1 U12485 ( .C1(n12363), .C2(n13018), .A(n9918), .B(n9917), .ZN(n9919) );
  INV_X1 U12486 ( .A(n9919), .ZN(n9920) );
  NAND2_X1 U12487 ( .A1(n13020), .A2(n12839), .ZN(n12501) );
  NAND2_X1 U12488 ( .A1(n12941), .A2(n12567), .ZN(n12498) );
  NAND2_X1 U12489 ( .A1(n12501), .A2(n12498), .ZN(n12820) );
  NAND2_X1 U12490 ( .A1(n13020), .A2(n12567), .ZN(n12806) );
  AND2_X1 U12491 ( .A1(n12944), .A2(n12568), .ZN(n12804) );
  NAND2_X1 U12492 ( .A1(n12820), .A2(n12804), .ZN(n9922) );
  NOR2_X1 U12493 ( .A1(n11566), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U12494 ( .A1(n11566), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n9923) );
  XNOR2_X1 U12495 ( .A(n11492), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n9938) );
  XNOR2_X1 U12496 ( .A(n9940), .B(n9938), .ZN(n13092) );
  NAND2_X1 U12497 ( .A1(n13092), .A2(n9956), .ZN(n9927) );
  NAND2_X1 U12498 ( .A1(n12368), .A2(SI_25_), .ZN(n9926) );
  INV_X1 U12499 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n9928) );
  NAND2_X1 U12500 ( .A1(n9929), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n9930) );
  NAND2_X1 U12501 ( .A1(n9945), .A2(n9930), .ZN(n12802) );
  NAND2_X1 U12502 ( .A1(n12802), .A2(n9991), .ZN(n9936) );
  INV_X1 U12503 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n9933) );
  NAND2_X1 U12504 ( .A1(n12360), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n9932) );
  NAND2_X1 U12505 ( .A1(n10012), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n9931) );
  OAI211_X1 U12506 ( .C1(n9933), .C2(n12363), .A(n9932), .B(n9931), .ZN(n9934)
         );
  INV_X1 U12507 ( .A(n9934), .ZN(n9935) );
  NAND2_X1 U12508 ( .A1(n13012), .A2(n12796), .ZN(n12508) );
  INV_X1 U12509 ( .A(n12505), .ZN(n9937) );
  INV_X1 U12510 ( .A(n9938), .ZN(n9939) );
  NAND2_X1 U12511 ( .A1(n15767), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n9941) );
  XNOR2_X1 U12512 ( .A(n15780), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n9952) );
  XNOR2_X1 U12513 ( .A(n9954), .B(n9952), .ZN(n13088) );
  NAND2_X1 U12514 ( .A1(n13088), .A2(n9956), .ZN(n9944) );
  NAND2_X1 U12515 ( .A1(n12368), .A2(SI_26_), .ZN(n9943) );
  NAND2_X1 U12516 ( .A1(n9945), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n9946) );
  NAND2_X1 U12517 ( .A1(n9961), .A2(n9946), .ZN(n12792) );
  INV_X1 U12518 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13007) );
  NAND2_X1 U12519 ( .A1(n10012), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n9948) );
  NAND2_X1 U12520 ( .A1(n12360), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n9947) );
  OAI211_X1 U12521 ( .C1(n12363), .C2(n13007), .A(n9948), .B(n9947), .ZN(n9949) );
  INV_X1 U12522 ( .A(n12269), .ZN(n12566) );
  INV_X1 U12523 ( .A(n13008), .ZN(n9951) );
  INV_X1 U12524 ( .A(n9952), .ZN(n9953) );
  NAND2_X1 U12525 ( .A1(n11621), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n9955) );
  XNOR2_X1 U12526 ( .A(n12206), .B(P2_DATAO_REG_27__SCAN_IN), .ZN(n9970) );
  XNOR2_X1 U12527 ( .A(n9972), .B(n9970), .ZN(n13084) );
  NAND2_X1 U12528 ( .A1(n13084), .A2(n9956), .ZN(n9958) );
  NAND2_X1 U12529 ( .A1(n12368), .A2(SI_27_), .ZN(n9957) );
  INV_X1 U12530 ( .A(n9961), .ZN(n9960) );
  INV_X1 U12531 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n9959) );
  NAND2_X1 U12532 ( .A1(n9961), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n9962) );
  NAND2_X1 U12533 ( .A1(n9976), .A2(n9962), .ZN(n12785) );
  NAND2_X1 U12534 ( .A1(n12785), .A2(n9991), .ZN(n9968) );
  INV_X1 U12535 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n9965) );
  NAND2_X1 U12536 ( .A1(n12360), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U12537 ( .A1(n10012), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n9963) );
  OAI211_X1 U12538 ( .C1(n9965), .C2(n12363), .A(n9964), .B(n9963), .ZN(n9966)
         );
  INV_X1 U12539 ( .A(n9966), .ZN(n9967) );
  NAND2_X1 U12540 ( .A1(n12932), .A2(n12345), .ZN(n12768) );
  INV_X1 U12541 ( .A(n9970), .ZN(n9971) );
  XNOR2_X1 U12542 ( .A(n9973), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n9983) );
  XNOR2_X1 U12543 ( .A(n9985), .B(n9983), .ZN(n13080) );
  NAND2_X1 U12544 ( .A1(n13080), .A2(n9956), .ZN(n9975) );
  NAND2_X1 U12545 ( .A1(n12368), .A2(SI_28_), .ZN(n9974) );
  NAND2_X1 U12546 ( .A1(n9976), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n9977) );
  NAND2_X1 U12547 ( .A1(n12756), .A2(n9977), .ZN(n12771) );
  INV_X1 U12548 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n13000) );
  NAND2_X1 U12549 ( .A1(n12360), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U12550 ( .A1(n6442), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n9978) );
  OAI211_X1 U12551 ( .C1(n13000), .C2(n12363), .A(n9979), .B(n9978), .ZN(n9980) );
  INV_X1 U12552 ( .A(n12230), .ZN(n12565) );
  INV_X1 U12553 ( .A(n9983), .ZN(n9984) );
  NAND2_X1 U12554 ( .A1(n9985), .A2(n9984), .ZN(n9987) );
  NAND2_X1 U12555 ( .A1(n15196), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n9986) );
  XNOR2_X1 U12556 ( .A(n14101), .B(P2_DATAO_REG_29__SCAN_IN), .ZN(n9988) );
  INV_X1 U12557 ( .A(SI_29_), .ZN(n12199) );
  NOR2_X1 U12558 ( .A1(n7167), .A2(n12199), .ZN(n9990) );
  INV_X1 U12559 ( .A(n12756), .ZN(n9992) );
  INV_X1 U12560 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n10089) );
  NAND2_X1 U12561 ( .A1(n10012), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n9994) );
  NAND2_X1 U12562 ( .A1(n9577), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n9993) );
  OAI211_X1 U12563 ( .C1(n10089), .C2(n10015), .A(n9994), .B(n9993), .ZN(n9995) );
  INV_X1 U12564 ( .A(n9995), .ZN(n9996) );
  NAND2_X1 U12565 ( .A1(n12366), .A2(n9996), .ZN(n12564) );
  AND2_X1 U12566 ( .A1(n12387), .A2(n12564), .ZN(n12351) );
  INV_X1 U12567 ( .A(n12387), .ZN(n9997) );
  NAND2_X1 U12568 ( .A1(n10022), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10006) );
  NAND2_X1 U12569 ( .A1(n12560), .A2(n12548), .ZN(n10098) );
  NAND2_X1 U12570 ( .A1(n10009), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10007) );
  NAND2_X1 U12571 ( .A1(n10026), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10008) );
  MUX2_X1 U12572 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10008), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n10010) );
  AND2_X1 U12573 ( .A1(n12400), .A2(n10097), .ZN(n12378) );
  INV_X1 U12574 ( .A(n12378), .ZN(n10011) );
  INV_X1 U12575 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n12928) );
  NAND2_X1 U12576 ( .A1(n9577), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n10014) );
  NAND2_X1 U12577 ( .A1(n6442), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n10013) );
  OAI211_X1 U12578 ( .C1(n6443), .C2(n12928), .A(n10014), .B(n10013), .ZN(
        n10016) );
  INV_X1 U12579 ( .A(n10016), .ZN(n10017) );
  INV_X1 U12580 ( .A(n13081), .ZN(n12556) );
  INV_X1 U12581 ( .A(n7168), .ZN(n12737) );
  NAND2_X1 U12582 ( .A1(n12556), .A2(n12737), .ZN(n10123) );
  INV_X1 U12583 ( .A(n10878), .ZN(n10876) );
  AND2_X2 U12584 ( .A1(n12560), .A2(n12400), .ZN(n12512) );
  INV_X1 U12585 ( .A(P3_B_REG_SCAN_IN), .ZN(n10030) );
  NOR2_X1 U12586 ( .A1(n13081), .A2(n10030), .ZN(n10018) );
  OR2_X1 U12587 ( .A1(n12838), .A2(n10018), .ZN(n12754) );
  NOR2_X1 U12588 ( .A1(n12387), .A2(n15626), .ZN(n12763) );
  NAND2_X1 U12589 ( .A1(n10024), .A2(n10023), .ZN(n10050) );
  INV_X1 U12590 ( .A(n10052), .ZN(n10028) );
  AND2_X1 U12591 ( .A1(n10042), .A2(P3_B_REG_SCAN_IN), .ZN(n10027) );
  NAND2_X1 U12592 ( .A1(n10028), .A2(n10027), .ZN(n10038) );
  XNOR2_X1 U12593 ( .A(n10031), .B(P3_IR_REG_31__SCAN_IN), .ZN(n10029) );
  NAND3_X1 U12594 ( .A1(n10042), .A2(P3_B_REG_SCAN_IN), .A3(n10029), .ZN(
        n10033) );
  NAND3_X1 U12595 ( .A1(n10031), .A2(n10030), .A3(n13074), .ZN(n10032) );
  OAI211_X1 U12596 ( .C1(n10042), .C2(P3_B_REG_SCAN_IN), .A(n10033), .B(n10032), .ZN(n10034) );
  INV_X1 U12597 ( .A(n10034), .ZN(n10035) );
  INV_X1 U12598 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10164) );
  NOR2_X1 U12599 ( .A1(n10048), .A2(n10047), .ZN(n10039) );
  INV_X1 U12600 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10040) );
  NAND2_X1 U12601 ( .A1(n10046), .A2(n10037), .ZN(n10043) );
  NAND2_X1 U12602 ( .A1(n10502), .A2(n10578), .ZN(n10094) );
  INV_X1 U12603 ( .A(n10578), .ZN(n10045) );
  INV_X1 U12604 ( .A(n10502), .ZN(n10070) );
  NAND2_X1 U12605 ( .A1(n10045), .A2(n10070), .ZN(n10505) );
  AND2_X1 U12606 ( .A1(n10094), .A2(n10505), .ZN(n10073) );
  INV_X1 U12607 ( .A(n10046), .ZN(n13097) );
  AND2_X1 U12608 ( .A1(n10047), .A2(n10048), .ZN(n10049) );
  NAND2_X1 U12609 ( .A1(n10050), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n10051) );
  MUX2_X1 U12610 ( .A(P3_IR_REG_31__SCAN_IN), .B(n10051), .S(
        P3_IR_REG_23__SCAN_IN), .Z(n10053) );
  INV_X1 U12611 ( .A(n10202), .ZN(n10064) );
  NOR2_X1 U12612 ( .A1(P3_D_REG_24__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .ZN(
        n15675) );
  NOR4_X1 U12613 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_7__SCAN_IN), .A4(P3_D_REG_17__SCAN_IN), .ZN(n10056) );
  NOR4_X1 U12614 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_29__SCAN_IN), .A4(P3_D_REG_10__SCAN_IN), .ZN(n10055) );
  NOR4_X1 U12615 ( .A1(P3_D_REG_22__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n10054) );
  NAND4_X1 U12616 ( .A1(n15675), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10062) );
  NOR4_X1 U12617 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_26__SCAN_IN), .A3(
        P3_D_REG_9__SCAN_IN), .A4(P3_D_REG_16__SCAN_IN), .ZN(n10060) );
  NOR4_X1 U12618 ( .A1(P3_D_REG_31__SCAN_IN), .A2(P3_D_REG_14__SCAN_IN), .A3(
        P3_D_REG_11__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n10059) );
  NOR4_X1 U12619 ( .A1(P3_D_REG_6__SCAN_IN), .A2(P3_D_REG_3__SCAN_IN), .A3(
        P3_D_REG_5__SCAN_IN), .A4(P3_D_REG_4__SCAN_IN), .ZN(n10058) );
  NOR4_X1 U12620 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_23__SCAN_IN), .A3(
        P3_D_REG_30__SCAN_IN), .A4(P3_D_REG_28__SCAN_IN), .ZN(n10057) );
  NAND4_X1 U12621 ( .A1(n10060), .A2(n10059), .A3(n10058), .A4(n10057), .ZN(
        n10061) );
  NOR2_X1 U12622 ( .A1(n10062), .A2(n10061), .ZN(n10063) );
  NOR2_X1 U12623 ( .A1(n10548), .A2(n10100), .ZN(n10507) );
  NAND3_X1 U12624 ( .A1(n12743), .A2(n12560), .A3(n10097), .ZN(n10087) );
  NAND2_X1 U12625 ( .A1(n10087), .A2(n12513), .ZN(n10504) );
  NAND2_X1 U12626 ( .A1(n12743), .A2(n12560), .ZN(n10065) );
  OAI21_X1 U12627 ( .B1(n15626), .B2(n10097), .A(n10065), .ZN(n10066) );
  NAND2_X1 U12628 ( .A1(n12743), .A2(n11334), .ZN(n12522) );
  NAND2_X1 U12629 ( .A1(n10066), .A2(n12522), .ZN(n10067) );
  NAND2_X1 U12630 ( .A1(n10067), .A2(n12513), .ZN(n10068) );
  NAND2_X1 U12631 ( .A1(n10070), .A2(n10068), .ZN(n10069) );
  INV_X1 U12632 ( .A(n12522), .ZN(n10085) );
  OAI211_X1 U12633 ( .C1(n10070), .C2(n10504), .A(n10069), .B(n10529), .ZN(
        n10071) );
  INV_X1 U12634 ( .A(n10071), .ZN(n10072) );
  NAND2_X1 U12635 ( .A1(n10586), .A2(n12401), .ZN(n12977) );
  NAND2_X1 U12636 ( .A1(n10075), .A2(n12407), .ZN(n10782) );
  INV_X1 U12637 ( .A(n12408), .ZN(n12411) );
  OR2_X1 U12638 ( .A1(n11096), .A2(n12579), .ZN(n12432) );
  NAND2_X1 U12639 ( .A1(n12432), .A2(n12425), .ZN(n10076) );
  XNOR2_X1 U12640 ( .A(n12435), .B(n12578), .ZN(n12530) );
  NAND2_X1 U12641 ( .A1(n11096), .A2(n12579), .ZN(n12431) );
  OAI211_X1 U12642 ( .C1(n11090), .C2(n10076), .A(n12530), .B(n12431), .ZN(
        n10077) );
  INV_X1 U12643 ( .A(n12578), .ZN(n12434) );
  NAND2_X1 U12644 ( .A1(n12435), .A2(n12434), .ZN(n12436) );
  OR2_X1 U12645 ( .A1(n11499), .A2(n12575), .ZN(n12448) );
  NAND2_X1 U12646 ( .A1(n11499), .A2(n12575), .ZN(n12447) );
  NAND2_X1 U12647 ( .A1(n12448), .A2(n12447), .ZN(n12533) );
  AND2_X1 U12648 ( .A1(n12286), .A2(n12905), .ZN(n12465) );
  INV_X1 U12649 ( .A(n12390), .ZN(n10079) );
  NAND2_X1 U12650 ( .A1(n12249), .A2(n12895), .ZN(n12482) );
  OR2_X1 U12651 ( .A1(n13038), .A2(n12485), .ZN(n12487) );
  NAND2_X1 U12652 ( .A1(n13032), .A2(n12320), .ZN(n12491) );
  OR2_X1 U12653 ( .A1(n13032), .A2(n12320), .ZN(n12490) );
  NAND2_X1 U12654 ( .A1(n13027), .A2(n12837), .ZN(n12389) );
  NAND2_X1 U12655 ( .A1(n12946), .A2(n12497), .ZN(n12817) );
  NOR2_X1 U12656 ( .A1(n13008), .A2(n12269), .ZN(n12506) );
  NAND2_X1 U12657 ( .A1(n13008), .A2(n12269), .ZN(n12509) );
  INV_X1 U12658 ( .A(n12768), .ZN(n10080) );
  NAND2_X1 U12659 ( .A1(n11461), .A2(n11334), .ZN(n10082) );
  XNOR2_X1 U12660 ( .A(n12560), .B(n10082), .ZN(n10084) );
  OR2_X1 U12661 ( .A1(n12400), .A2(n12548), .ZN(n10083) );
  NAND2_X1 U12662 ( .A1(n10084), .A2(n10083), .ZN(n10539) );
  AND2_X1 U12663 ( .A1(n15626), .A2(n10085), .ZN(n10086) );
  NAND2_X1 U12664 ( .A1(n10539), .A2(n10086), .ZN(n10088) );
  NAND2_X1 U12665 ( .A1(n12548), .A2(n11334), .ZN(n12521) );
  NAND2_X1 U12666 ( .A1(n15665), .A2(n15630), .ZN(n12971) );
  INV_X1 U12667 ( .A(n10094), .ZN(n10096) );
  INV_X1 U12668 ( .A(n10100), .ZN(n10095) );
  NAND2_X1 U12669 ( .A1(n10096), .A2(n10095), .ZN(n10545) );
  INV_X1 U12670 ( .A(n12549), .ZN(n10099) );
  AND2_X1 U12671 ( .A1(n10541), .A2(n10535), .ZN(n10102) );
  INV_X1 U12672 ( .A(n10539), .ZN(n10101) );
  OAI22_X1 U12673 ( .A1(n10545), .A2(n10102), .B1(n10101), .B2(n10540), .ZN(
        n10103) );
  OR2_X1 U12674 ( .A1(n15654), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n10104) );
  INV_X1 U12675 ( .A(n11449), .ZN(n10724) );
  NOR2_X1 U12676 ( .A1(n10106), .A2(P1_U3086), .ZN(n10107) );
  OAI21_X1 U12677 ( .B1(n10109), .B2(n13542), .A(n10108), .ZN(n10110) );
  INV_X1 U12678 ( .A(n13880), .ZN(n13274) );
  OAI22_X1 U12679 ( .A1(n11183), .A2(n13274), .B1(n13304), .B2(n13273), .ZN(
        n11040) );
  AOI21_X1 U12680 ( .B1(n10110), .B2(n13897), .A(n11040), .ZN(n10111) );
  INV_X1 U12681 ( .A(n10111), .ZN(n10793) );
  MUX2_X1 U12682 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10793), .S(n13913), .Z(
        n10120) );
  OAI21_X1 U12683 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10795) );
  INV_X1 U12684 ( .A(n10795), .ZN(n10115) );
  NOR2_X1 U12685 ( .A1(n13908), .A2(n10115), .ZN(n10119) );
  AOI21_X1 U12686 ( .B1(n11207), .B2(n13286), .A(n6409), .ZN(n10116) );
  AND2_X1 U12687 ( .A1(n11010), .A2(n10116), .ZN(n10794) );
  AND2_X1 U12688 ( .A1(n13919), .A2(n10794), .ZN(n10118) );
  OAI22_X1 U12689 ( .A1(n13904), .A2(n6888), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n13843), .ZN(n10117) );
  OR4_X1 U12690 ( .A1(n10120), .A2(n10119), .A3(n10118), .A4(n10117), .ZN(
        P2_U3262) );
  AND2_X1 U12691 ( .A1(n10121), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12554) );
  INV_X1 U12692 ( .A(n12554), .ZN(n12559) );
  NAND2_X1 U12693 ( .A1(n10548), .A2(n12559), .ZN(n10133) );
  OAI21_X1 U12694 ( .B1(n10121), .B2(n12513), .A(n9529), .ZN(n10132) );
  INV_X1 U12695 ( .A(n10132), .ZN(n10122) );
  NAND2_X1 U12696 ( .A1(n10133), .A2(n10122), .ZN(n10125) );
  MUX2_X1 U12697 ( .A(n10125), .B(n12571), .S(n12556), .Z(n15549) );
  INV_X1 U12698 ( .A(n15549), .ZN(n15598) );
  NOR2_X1 U12699 ( .A1(n15570), .A2(n7410), .ZN(n10124) );
  MUX2_X1 U12700 ( .A(n15598), .B(n10124), .S(n10140), .Z(n10139) );
  INV_X1 U12701 ( .A(n10125), .ZN(n10126) );
  NOR2_X1 U12702 ( .A1(n15591), .A2(n15595), .ZN(n10128) );
  MUX2_X1 U12703 ( .A(n7410), .B(n10127), .S(n13085), .Z(n10130) );
  NAND2_X1 U12704 ( .A1(n10130), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10384) );
  AOI21_X1 U12705 ( .B1(n10128), .B2(n15570), .A(n10384), .ZN(n10138) );
  NAND2_X1 U12706 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n10140), .ZN(n10409) );
  INV_X1 U12707 ( .A(n10409), .ZN(n10129) );
  AND2_X1 U12708 ( .A1(n15591), .A2(n10129), .ZN(n10137) );
  INV_X1 U12709 ( .A(n10130), .ZN(n10131) );
  NAND3_X1 U12710 ( .A1(n15595), .A2(n10131), .A3(n10140), .ZN(n10135) );
  NAND2_X1 U12711 ( .A1(n15539), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n10134) );
  OAI211_X1 U12712 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10553), .A(n10135), .B(
        n10134), .ZN(n10136) );
  OR4_X1 U12713 ( .A1(n10139), .A2(n10138), .A3(n10137), .A4(n10136), .ZN(
        P3_U3182) );
  OR2_X1 U12714 ( .A1(P3_U3151), .A2(n10140), .ZN(n10141) );
  OAI21_X1 U12715 ( .B1(n10142), .B2(P3_STATE_REG_SCAN_IN), .A(n10141), .ZN(
        P3_U3295) );
  AND2_X1 U12716 ( .A1(n8017), .A2(P3_U3151), .ZN(n11742) );
  INV_X2 U12717 ( .A(n11742), .ZN(n13090) );
  NAND2_X2 U12718 ( .A1(n7875), .A2(P3_U3151), .ZN(n13095) );
  OAI222_X1 U12719 ( .A1(n13090), .A2(n10144), .B1(n13095), .B2(n10143), .C1(
        P3_U3151), .C2(n10528), .ZN(P3_U3294) );
  OAI222_X1 U12720 ( .A1(P3_U3151), .A2(n10443), .B1(n13095), .B2(n6424), .C1(
        n13090), .C2(n10145), .ZN(P3_U3291) );
  INV_X1 U12721 ( .A(SI_3_), .ZN(n10147) );
  OAI222_X1 U12722 ( .A1(P3_U3151), .A2(n10680), .B1(n13095), .B2(n10147), 
        .C1(n13090), .C2(n10146), .ZN(P3_U3292) );
  INV_X1 U12723 ( .A(SI_5_), .ZN(n10149) );
  OAI222_X1 U12724 ( .A1(P3_U3151), .A2(n10682), .B1(n13095), .B2(n10149), 
        .C1(n13090), .C2(n10148), .ZN(P3_U3290) );
  OAI222_X1 U12725 ( .A1(n10634), .A2(P3_U3151), .B1(n13090), .B2(n10151), 
        .C1(n10150), .C2(n13095), .ZN(P3_U3293) );
  NOR2_X1 U12726 ( .A1(n7875), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14093) );
  INV_X2 U12727 ( .A(n14093), .ZN(n14102) );
  OAI222_X1 U12728 ( .A1(n14102), .A2(n10152), .B1(n14099), .B2(n10165), .C1(
        P2_U3088), .C2(n10350), .ZN(P2_U3325) );
  OAI222_X1 U12729 ( .A1(n15379), .A2(P2_U3088), .B1(n14099), .B2(n10189), 
        .C1(n10153), .C2(n14102), .ZN(P2_U3326) );
  INV_X1 U12730 ( .A(n10154), .ZN(n10155) );
  OAI222_X1 U12731 ( .A1(P3_U3151), .A2(n15550), .B1(n13095), .B2(n10156), 
        .C1(n13090), .C2(n10155), .ZN(P3_U3289) );
  INV_X1 U12732 ( .A(n10317), .ZN(n15391) );
  OAI222_X1 U12733 ( .A1(n14102), .A2(n10157), .B1(n14099), .B2(n10167), .C1(
        P2_U3088), .C2(n15391), .ZN(P2_U3324) );
  INV_X1 U12734 ( .A(n11228), .ZN(n11219) );
  INV_X1 U12735 ( .A(SI_7_), .ZN(n10159) );
  OAI222_X1 U12736 ( .A1(P3_U3151), .A2(n11219), .B1(n13095), .B2(n10159), 
        .C1(n13090), .C2(n10158), .ZN(P3_U3288) );
  INV_X1 U12737 ( .A(n10160), .ZN(n10169) );
  OAI222_X1 U12738 ( .A1(n14102), .A2(n10161), .B1(n14099), .B2(n10169), .C1(
        P2_U3088), .C2(n15403), .ZN(P2_U3323) );
  NAND2_X1 U12739 ( .A1(n10502), .A2(n10163), .ZN(n10162) );
  OAI21_X1 U12740 ( .B1(n10164), .B2(n10163), .A(n10162), .ZN(P3_U3377) );
  NAND2_X1 U12741 ( .A1(n8209), .A2(P1_U3086), .ZN(n15195) );
  OAI222_X1 U12742 ( .A1(n15189), .A2(n10166), .B1(n15195), .B2(n10165), .C1(
        P1_U3086), .C2(n10267), .ZN(P1_U3353) );
  OAI222_X1 U12743 ( .A1(n15189), .A2(n10168), .B1(n15195), .B2(n10167), .C1(
        P1_U3086), .C2(n14589), .ZN(P1_U3352) );
  OAI222_X1 U12744 ( .A1(n15189), .A2(n10170), .B1(n15195), .B2(n10169), .C1(
        P1_U3086), .C2(n10272), .ZN(P1_U3351) );
  INV_X1 U12745 ( .A(n10171), .ZN(n10172) );
  OAI222_X1 U12746 ( .A1(P3_U3151), .A2(n11239), .B1(n13095), .B2(n10173), 
        .C1(n13090), .C2(n10172), .ZN(P3_U3287) );
  INV_X1 U12747 ( .A(SI_9_), .ZN(n10175) );
  OAI222_X1 U12748 ( .A1(P3_U3151), .A2(n11694), .B1(n13095), .B2(n10175), 
        .C1(n13090), .C2(n10174), .ZN(P3_U3286) );
  INV_X1 U12749 ( .A(n10176), .ZN(n10178) );
  INV_X1 U12750 ( .A(n10362), .ZN(n10330) );
  OAI222_X1 U12751 ( .A1(n14102), .A2(n10177), .B1(n14099), .B2(n10178), .C1(
        P2_U3088), .C2(n10330), .ZN(P2_U3322) );
  INV_X1 U12752 ( .A(n14622), .ZN(n10255) );
  OAI222_X1 U12753 ( .A1(n15189), .A2(n10179), .B1(n15195), .B2(n10178), .C1(
        P1_U3086), .C2(n10255), .ZN(P1_U3350) );
  INV_X1 U12754 ( .A(n10180), .ZN(n10191) );
  AOI22_X1 U12755 ( .A1(n13615), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n14093), .ZN(n10181) );
  OAI21_X1 U12756 ( .B1(n10191), .B2(n14099), .A(n10181), .ZN(P2_U3321) );
  INV_X1 U12757 ( .A(n10244), .ZN(n10183) );
  NOR3_X1 U12758 ( .A1(n10183), .A2(n10182), .A3(P1_U3086), .ZN(n10187) );
  INV_X1 U12759 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U12760 ( .A1(n10187), .A2(n11489), .B1(n10185), .B2(n15666), .ZN(
        P1_U3446) );
  AOI22_X1 U12761 ( .A1(n10187), .A2(n11564), .B1(n10186), .B2(n15666), .ZN(
        P1_U3445) );
  CLKBUF_X1 U12762 ( .A(n15195), .Z(n15192) );
  OAI222_X1 U12763 ( .A1(n10264), .A2(P1_U3086), .B1(n15192), .B2(n10189), 
        .C1(n10188), .C2(n15189), .ZN(P1_U3354) );
  INV_X1 U12764 ( .A(n10481), .ZN(n10190) );
  OAI222_X1 U12765 ( .A1(n15189), .A2(n15751), .B1(n15195), .B2(n10191), .C1(
        P1_U3086), .C2(n10190), .ZN(P1_U3349) );
  INV_X1 U12766 ( .A(n15597), .ZN(n11698) );
  INV_X1 U12767 ( .A(SI_10_), .ZN(n10193) );
  OAI222_X1 U12768 ( .A1(P3_U3151), .A2(n11698), .B1(n13095), .B2(n10193), 
        .C1(n13090), .C2(n10192), .ZN(P3_U3285) );
  INV_X1 U12769 ( .A(n10194), .ZN(n10198) );
  INV_X1 U12770 ( .A(n14636), .ZN(n10195) );
  OAI222_X1 U12771 ( .A1(n15189), .A2(n10196), .B1(n15195), .B2(n10198), .C1(
        P1_U3086), .C2(n10195), .ZN(P1_U3348) );
  INV_X1 U12772 ( .A(n13628), .ZN(n10197) );
  OAI222_X1 U12773 ( .A1(n14102), .A2(n10199), .B1(n14099), .B2(n10198), .C1(
        P2_U3088), .C2(n10197), .ZN(P2_U3320) );
  INV_X1 U12774 ( .A(n12600), .ZN(n11703) );
  OAI222_X1 U12775 ( .A1(P3_U3151), .A2(n11703), .B1(n13095), .B2(n10201), 
        .C1(n13090), .C2(n10200), .ZN(P3_U3284) );
  NOR2_X1 U12776 ( .A1(n13072), .A2(n10202), .ZN(n10207) );
  CLKBUF_X1 U12777 ( .A(n10207), .Z(n10231) );
  INV_X1 U12778 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n10203) );
  NOR2_X1 U12779 ( .A1(n10231), .A2(n10203), .ZN(P3_U3257) );
  INV_X1 U12780 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n10204) );
  NOR2_X1 U12781 ( .A1(n10231), .A2(n10204), .ZN(P3_U3255) );
  INV_X1 U12782 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n10205) );
  NOR2_X1 U12783 ( .A1(n10231), .A2(n10205), .ZN(P3_U3249) );
  INV_X1 U12784 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n10206) );
  NOR2_X1 U12785 ( .A1(n10231), .A2(n10206), .ZN(P3_U3254) );
  INV_X1 U12786 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n10208) );
  NOR2_X1 U12787 ( .A1(n10231), .A2(n10208), .ZN(P3_U3244) );
  INV_X1 U12788 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U12789 ( .A1(n10231), .A2(n10209), .ZN(P3_U3256) );
  INV_X1 U12790 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n10210) );
  NOR2_X1 U12791 ( .A1(n10231), .A2(n10210), .ZN(P3_U3247) );
  INV_X1 U12792 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n15713) );
  NOR2_X1 U12793 ( .A1(n10207), .A2(n15713), .ZN(P3_U3241) );
  INV_X1 U12794 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n10211) );
  NOR2_X1 U12795 ( .A1(n10207), .A2(n10211), .ZN(P3_U3243) );
  INV_X1 U12796 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U12797 ( .A1(n10231), .A2(n10212), .ZN(P3_U3253) );
  INV_X1 U12798 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n15792) );
  NOR2_X1 U12799 ( .A1(n10231), .A2(n15792), .ZN(P3_U3252) );
  INV_X1 U12800 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n10213) );
  NOR2_X1 U12801 ( .A1(n10207), .A2(n10213), .ZN(P3_U3240) );
  INV_X1 U12802 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n10214) );
  NOR2_X1 U12803 ( .A1(n10207), .A2(n10214), .ZN(P3_U3260) );
  INV_X1 U12804 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n10215) );
  NOR2_X1 U12805 ( .A1(n10207), .A2(n10215), .ZN(P3_U3238) );
  INV_X1 U12806 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n10216) );
  NOR2_X1 U12807 ( .A1(n10231), .A2(n10216), .ZN(P3_U3250) );
  INV_X1 U12808 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n10217) );
  NOR2_X1 U12809 ( .A1(n10207), .A2(n10217), .ZN(P3_U3237) );
  INV_X1 U12810 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U12811 ( .A1(n10231), .A2(n10218), .ZN(P3_U3248) );
  INV_X1 U12812 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n10219) );
  NOR2_X1 U12813 ( .A1(n10207), .A2(n10219), .ZN(P3_U3236) );
  INV_X1 U12814 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n10220) );
  NOR2_X1 U12815 ( .A1(n10207), .A2(n10220), .ZN(P3_U3235) );
  INV_X1 U12816 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n10221) );
  NOR2_X1 U12817 ( .A1(n10207), .A2(n10221), .ZN(P3_U3239) );
  INV_X1 U12818 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U12819 ( .A1(n10207), .A2(n10222), .ZN(P3_U3234) );
  INV_X1 U12820 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n10223) );
  NOR2_X1 U12821 ( .A1(n10231), .A2(n10223), .ZN(P3_U3246) );
  INV_X1 U12822 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U12823 ( .A1(n10207), .A2(n10224), .ZN(P3_U3245) );
  INV_X1 U12824 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n15712) );
  NOR2_X1 U12825 ( .A1(n10231), .A2(n15712), .ZN(P3_U3258) );
  INV_X1 U12826 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U12827 ( .A1(n10231), .A2(n10225), .ZN(P3_U3259) );
  INV_X1 U12828 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n10226) );
  NOR2_X1 U12829 ( .A1(n10231), .A2(n10226), .ZN(P3_U3242) );
  INV_X1 U12830 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n10227) );
  NOR2_X1 U12831 ( .A1(n10231), .A2(n10227), .ZN(P3_U3251) );
  INV_X1 U12832 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n10228) );
  NOR2_X1 U12833 ( .A1(n10231), .A2(n10228), .ZN(P3_U3261) );
  INV_X1 U12834 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n10229) );
  NOR2_X1 U12835 ( .A1(n10231), .A2(n10229), .ZN(P3_U3262) );
  INV_X1 U12836 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n10230) );
  NOR2_X1 U12837 ( .A1(n10231), .A2(n10230), .ZN(P3_U3263) );
  OAI222_X1 U12838 ( .A1(P3_U3151), .A2(n12612), .B1(n13095), .B2(n10233), 
        .C1(n13090), .C2(n10232), .ZN(P3_U3283) );
  INV_X1 U12839 ( .A(n10234), .ZN(n10237) );
  INV_X1 U12840 ( .A(n10369), .ZN(n15415) );
  OAI222_X1 U12841 ( .A1(n14102), .A2(n10235), .B1(n14099), .B2(n10237), .C1(
        P2_U3088), .C2(n15415), .ZN(P2_U3319) );
  INV_X1 U12842 ( .A(n14648), .ZN(n10236) );
  OAI222_X1 U12843 ( .A1(n15189), .A2(n10238), .B1(n15195), .B2(n10237), .C1(
        P1_U3086), .C2(n10236), .ZN(P1_U3347) );
  INV_X1 U12844 ( .A(n10239), .ZN(n10241) );
  OAI222_X1 U12845 ( .A1(n14102), .A2(n10240), .B1(n14099), .B2(n10241), .C1(
        P2_U3088), .C2(n10944), .ZN(P2_U3318) );
  INV_X1 U12846 ( .A(n14666), .ZN(n10472) );
  OAI222_X1 U12847 ( .A1(n15189), .A2(n10242), .B1(n15195), .B2(n10241), .C1(
        P1_U3086), .C2(n10472), .ZN(P1_U3346) );
  OR2_X1 U12848 ( .A1(n10244), .A2(P1_U3086), .ZN(n14539) );
  INV_X1 U12849 ( .A(n14539), .ZN(n11451) );
  OR2_X1 U12850 ( .A1(n10813), .A2(n11451), .ZN(n10247) );
  AOI21_X1 U12851 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(n10246) );
  NAND2_X1 U12852 ( .A1(n10247), .A2(n10246), .ZN(n15249) );
  NOR2_X2 U12853 ( .A1(n15249), .A2(n14571), .ZN(n14735) );
  INV_X1 U12854 ( .A(n10246), .ZN(n10248) );
  AND2_X1 U12855 ( .A1(n10248), .A2(n10247), .ZN(n15247) );
  NAND2_X1 U12856 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n10249) );
  OAI21_X1 U12857 ( .B1(n14742), .B2(n15782), .A(n10249), .ZN(n10263) );
  XNOR2_X1 U12858 ( .A(n10481), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n10261) );
  MUX2_X1 U12859 ( .A(n8878), .B(P1_REG1_REG_1__SCAN_IN), .S(n10264), .Z(
        n14561) );
  AND2_X1 U12860 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14560) );
  NAND2_X1 U12861 ( .A1(n14561), .A2(n14560), .ZN(n14559) );
  INV_X1 U12862 ( .A(n10264), .ZN(n14562) );
  NAND2_X1 U12863 ( .A1(n14562), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n10250) );
  NAND2_X1 U12864 ( .A1(n14559), .A2(n10250), .ZN(n14577) );
  MUX2_X1 U12865 ( .A(n8923), .B(P1_REG1_REG_2__SCAN_IN), .S(n10267), .Z(
        n14578) );
  NAND2_X1 U12866 ( .A1(n14577), .A2(n14578), .ZN(n14576) );
  INV_X1 U12867 ( .A(n10267), .ZN(n14585) );
  NAND2_X1 U12868 ( .A1(n14585), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n10251) );
  NAND2_X1 U12869 ( .A1(n14576), .A2(n10251), .ZN(n14595) );
  XNOR2_X1 U12870 ( .A(n14589), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n14596) );
  NAND2_X1 U12871 ( .A1(n14595), .A2(n14596), .ZN(n14594) );
  OR2_X1 U12872 ( .A1(n14589), .A2(n10252), .ZN(n10253) );
  NAND2_X1 U12873 ( .A1(n14594), .A2(n10253), .ZN(n14606) );
  MUX2_X1 U12874 ( .A(n8957), .B(P1_REG1_REG_4__SCAN_IN), .S(n10272), .Z(
        n14607) );
  NAND2_X1 U12875 ( .A1(n14606), .A2(n14607), .ZN(n14605) );
  INV_X1 U12876 ( .A(n10272), .ZN(n14614) );
  NAND2_X1 U12877 ( .A1(n14614), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10254) );
  AND2_X1 U12878 ( .A1(n14605), .A2(n10254), .ZN(n14625) );
  MUX2_X1 U12879 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n15360), .S(n14622), .Z(
        n14624) );
  NAND2_X1 U12880 ( .A1(n14625), .A2(n14624), .ZN(n14623) );
  NAND2_X1 U12881 ( .A1(n10255), .A2(n15360), .ZN(n10256) );
  NAND2_X1 U12882 ( .A1(n14623), .A2(n10256), .ZN(n10260) );
  INV_X1 U12883 ( .A(n10466), .ZN(n10259) );
  INV_X1 U12884 ( .A(n15249), .ZN(n10258) );
  XNOR2_X1 U12885 ( .A(n10257), .B(P1_IR_REG_27__SCAN_IN), .ZN(n15245) );
  INV_X1 U12886 ( .A(n15245), .ZN(n14573) );
  NAND2_X1 U12887 ( .A1(n10258), .A2(n14573), .ZN(n14733) );
  AOI211_X1 U12888 ( .C1(n10261), .C2(n10260), .A(n10259), .B(n14733), .ZN(
        n10262) );
  AOI211_X1 U12889 ( .C1(n14735), .C2(n10481), .A(n10263), .B(n10262), .ZN(
        n10281) );
  INV_X1 U12890 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11353) );
  XNOR2_X1 U12891 ( .A(n10481), .B(n11353), .ZN(n10279) );
  INV_X1 U12892 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n10265) );
  MUX2_X1 U12893 ( .A(n10265), .B(P1_REG2_REG_1__SCAN_IN), .S(n10264), .Z(
        n14564) );
  AND2_X1 U12894 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14574) );
  NAND2_X1 U12895 ( .A1(n14564), .A2(n14574), .ZN(n14563) );
  NAND2_X1 U12896 ( .A1(n14562), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U12897 ( .A1(n14563), .A2(n10266), .ZN(n14580) );
  INV_X1 U12898 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10268) );
  MUX2_X1 U12899 ( .A(n10268), .B(P1_REG2_REG_2__SCAN_IN), .S(n10267), .Z(
        n14581) );
  NAND2_X1 U12900 ( .A1(n14580), .A2(n14581), .ZN(n14579) );
  NAND2_X1 U12901 ( .A1(n14585), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12902 ( .A1(n14579), .A2(n10269), .ZN(n14598) );
  XNOR2_X1 U12903 ( .A(n14589), .B(P1_REG2_REG_3__SCAN_IN), .ZN(n14599) );
  NAND2_X1 U12904 ( .A1(n14598), .A2(n14599), .ZN(n14597) );
  INV_X1 U12905 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10270) );
  OR2_X1 U12906 ( .A1(n14589), .A2(n10270), .ZN(n10271) );
  NAND2_X1 U12907 ( .A1(n14597), .A2(n10271), .ZN(n14609) );
  INV_X1 U12908 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10273) );
  MUX2_X1 U12909 ( .A(n10273), .B(P1_REG2_REG_4__SCAN_IN), .S(n10272), .Z(
        n14610) );
  NAND2_X1 U12910 ( .A1(n14609), .A2(n14610), .ZN(n14608) );
  NAND2_X1 U12911 ( .A1(n14614), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n10274) );
  NAND2_X1 U12912 ( .A1(n14608), .A2(n10274), .ZN(n14628) );
  INV_X1 U12913 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10275) );
  MUX2_X1 U12914 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10275), .S(n14622), .Z(
        n14629) );
  NAND2_X1 U12915 ( .A1(n14628), .A2(n14629), .ZN(n14627) );
  NAND2_X1 U12916 ( .A1(n14622), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10276) );
  NAND2_X1 U12917 ( .A1(n14627), .A2(n10276), .ZN(n10278) );
  NAND2_X1 U12918 ( .A1(n14571), .A2(n15245), .ZN(n10277) );
  NOR2_X2 U12919 ( .A1(n15249), .A2(n10277), .ZN(n14737) );
  NAND2_X1 U12920 ( .A1(n10278), .A2(n10279), .ZN(n10483) );
  OAI211_X1 U12921 ( .C1(n10279), .C2(n10278), .A(n14737), .B(n10483), .ZN(
        n10280) );
  NAND2_X1 U12922 ( .A1(n10281), .A2(n10280), .ZN(P1_U3249) );
  NOR2_X1 U12923 ( .A1(n15247), .A2(P1_U4016), .ZN(P1_U3085) );
  OAI222_X1 U12924 ( .A1(P3_U3151), .A2(n12637), .B1(n13095), .B2(n10283), 
        .C1(n13090), .C2(n10282), .ZN(P3_U3282) );
  INV_X1 U12925 ( .A(n10284), .ZN(n10288) );
  INV_X1 U12926 ( .A(n10841), .ZN(n10285) );
  OAI222_X1 U12927 ( .A1(n15189), .A2(n10286), .B1(n15192), .B2(n10288), .C1(
        P1_U3086), .C2(n10285), .ZN(P1_U3345) );
  INV_X1 U12928 ( .A(n15428), .ZN(n10287) );
  OAI222_X1 U12929 ( .A1(n14102), .A2(n10289), .B1(n14099), .B2(n10288), .C1(
        P2_U3088), .C2(n10287), .ZN(P2_U3317) );
  OAI21_X1 U12930 ( .B1(n10292), .B2(n10291), .A(n10290), .ZN(n14570) );
  AOI22_X1 U12931 ( .A1(n14273), .A2(n14570), .B1(n14269), .B2(n15276), .ZN(
        n10295) );
  NAND2_X1 U12932 ( .A1(n14282), .A2(n15010), .ZN(n14267) );
  INV_X1 U12933 ( .A(n14267), .ZN(n14209) );
  OR2_X1 U12934 ( .A1(n10293), .A2(P1_U3086), .ZN(n10760) );
  AOI22_X1 U12935 ( .A1(n14209), .A2(n8892), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n10760), .ZN(n10294) );
  NAND2_X1 U12936 ( .A1(n10295), .A2(n10294), .ZN(P1_U3232) );
  NAND2_X1 U12937 ( .A1(n11449), .A2(n10563), .ZN(n10297) );
  NAND2_X1 U12938 ( .A1(n10297), .A2(n10296), .ZN(n10298) );
  AND2_X1 U12939 ( .A1(n10299), .A2(n10298), .ZN(n10300) );
  AND2_X1 U12940 ( .A1(n10323), .A2(n10307), .ZN(n15432) );
  AND2_X1 U12941 ( .A1(n10300), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15368) );
  NAND2_X1 U12942 ( .A1(n15368), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n10328) );
  XNOR2_X1 U12943 ( .A(n10362), .B(n10301), .ZN(n10310) );
  AND2_X1 U12944 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n10302) );
  NAND2_X1 U12945 ( .A1(n10312), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10303) );
  NAND2_X1 U12946 ( .A1(n15376), .A2(n10303), .ZN(n10344) );
  MUX2_X1 U12947 ( .A(n8034), .B(P2_REG1_REG_2__SCAN_IN), .S(n10350), .Z(
        n10345) );
  NAND2_X1 U12948 ( .A1(n10314), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U12949 ( .A1(n10343), .A2(n10304), .ZN(n15387) );
  MUX2_X1 U12950 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n8060), .S(n10317), .Z(
        n15388) );
  NAND2_X1 U12951 ( .A1(n15387), .A2(n15388), .ZN(n15386) );
  NAND2_X1 U12952 ( .A1(n10317), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10305) );
  NAND2_X1 U12953 ( .A1(n15386), .A2(n10305), .ZN(n15399) );
  MUX2_X1 U12954 ( .A(n8079), .B(P2_REG1_REG_4__SCAN_IN), .S(n15403), .Z(
        n15400) );
  NAND2_X1 U12955 ( .A1(n15399), .A2(n15400), .ZN(n15398) );
  NAND2_X1 U12956 ( .A1(n10320), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n10306) );
  NAND2_X1 U12957 ( .A1(n15398), .A2(n10306), .ZN(n10309) );
  NOR2_X1 U12958 ( .A1(n10307), .A2(P2_U3088), .ZN(n11862) );
  AND2_X1 U12959 ( .A1(n11862), .A2(n12205), .ZN(n10308) );
  NAND2_X1 U12960 ( .A1(n10323), .A2(n10308), .ZN(n15492) );
  NAND2_X1 U12961 ( .A1(n10309), .A2(n10310), .ZN(n10364) );
  OAI211_X1 U12962 ( .C1(n10310), .C2(n10309), .A(n15460), .B(n10364), .ZN(
        n10327) );
  NAND2_X1 U12963 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n10722) );
  XNOR2_X1 U12964 ( .A(n10362), .B(n10311), .ZN(n10325) );
  INV_X1 U12965 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n15797) );
  MUX2_X1 U12966 ( .A(n15797), .B(P2_REG2_REG_1__SCAN_IN), .S(n15379), .Z(
        n15371) );
  AND2_X1 U12967 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n15370) );
  NAND2_X1 U12968 ( .A1(n15371), .A2(n15370), .ZN(n15369) );
  NAND2_X1 U12969 ( .A1(n10312), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n10313) );
  NAND2_X1 U12970 ( .A1(n15369), .A2(n10313), .ZN(n10340) );
  INV_X1 U12971 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n11209) );
  MUX2_X1 U12972 ( .A(n11209), .B(P2_REG2_REG_2__SCAN_IN), .S(n10350), .Z(
        n10341) );
  NAND2_X1 U12973 ( .A1(n10340), .A2(n10341), .ZN(n10339) );
  NAND2_X1 U12974 ( .A1(n10314), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10315) );
  NAND2_X1 U12975 ( .A1(n10339), .A2(n10315), .ZN(n15384) );
  INV_X1 U12976 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10316) );
  MUX2_X1 U12977 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n10316), .S(n10317), .Z(
        n15385) );
  NAND2_X1 U12978 ( .A1(n15384), .A2(n15385), .ZN(n15383) );
  NAND2_X1 U12979 ( .A1(n10317), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10318) );
  NAND2_X1 U12980 ( .A1(n15383), .A2(n10318), .ZN(n15396) );
  INV_X1 U12981 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U12982 ( .A(n10319), .B(P2_REG2_REG_4__SCAN_IN), .S(n15403), .Z(
        n15397) );
  NAND2_X1 U12983 ( .A1(n15396), .A2(n15397), .ZN(n15395) );
  NAND2_X1 U12984 ( .A1(n10320), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n10321) );
  NAND2_X1 U12985 ( .A1(n15395), .A2(n10321), .ZN(n10324) );
  AND2_X1 U12986 ( .A1(n11862), .A2(n13575), .ZN(n10322) );
  NAND2_X1 U12987 ( .A1(n10324), .A2(n10325), .ZN(n10352) );
  OAI211_X1 U12988 ( .C1(n10325), .C2(n10324), .A(n15486), .B(n10352), .ZN(
        n10326) );
  AND4_X1 U12989 ( .A1(n10328), .A2(n10327), .A3(n10722), .A4(n10326), .ZN(
        n10329) );
  OAI21_X1 U12990 ( .B1(n10330), .B2(n15468), .A(n10329), .ZN(P2_U3219) );
  INV_X1 U12991 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n15735) );
  NAND2_X1 U12992 ( .A1(n12916), .A2(P3_U3897), .ZN(n10331) );
  OAI21_X1 U12993 ( .B1(P3_U3897), .B2(n15735), .A(n10331), .ZN(P3_U3508) );
  AOI22_X1 U12994 ( .A1(n15460), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15486), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10336) );
  INV_X1 U12995 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10332) );
  NAND2_X1 U12996 ( .A1(n15486), .A2(n10332), .ZN(n10333) );
  OAI211_X1 U12997 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n15492), .A(n15468), .B(
        n10333), .ZN(n10334) );
  INV_X1 U12998 ( .A(n10334), .ZN(n10335) );
  MUX2_X1 U12999 ( .A(n10336), .B(n10335), .S(P2_IR_REG_0__SCAN_IN), .Z(n10338) );
  AOI22_X1 U13000 ( .A1(n15368), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n10337) );
  NAND2_X1 U13001 ( .A1(n10338), .A2(n10337), .ZN(P2_U3214) );
  OAI211_X1 U13002 ( .C1(n10341), .C2(n10340), .A(n15486), .B(n10339), .ZN(
        n10342) );
  INV_X1 U13003 ( .A(n10342), .ZN(n10348) );
  OAI211_X1 U13004 ( .C1(n10345), .C2(n10344), .A(n15460), .B(n10343), .ZN(
        n10346) );
  OAI21_X1 U13005 ( .B1(P2_STATE_REG_SCAN_IN), .B2(n11208), .A(n10346), .ZN(
        n10347) );
  AOI211_X1 U13006 ( .C1(n15368), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10348), .B(
        n10347), .ZN(n10349) );
  OAI21_X1 U13007 ( .B1(n10350), .B2(n15468), .A(n10349), .ZN(P2_U3216) );
  MUX2_X1 U13008 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n11612), .S(n10944), .Z(
        n10360) );
  NAND2_X1 U13009 ( .A1(n10362), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10351) );
  NAND2_X1 U13010 ( .A1(n10352), .A2(n10351), .ZN(n13617) );
  XNOR2_X1 U13011 ( .A(n13615), .B(n10353), .ZN(n13618) );
  NAND2_X1 U13012 ( .A1(n13617), .A2(n13618), .ZN(n13616) );
  NAND2_X1 U13013 ( .A1(n13615), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n10354) );
  NAND2_X1 U13014 ( .A1(n13616), .A2(n10354), .ZN(n13633) );
  XNOR2_X1 U13015 ( .A(n13628), .B(n11175), .ZN(n13634) );
  NAND2_X1 U13016 ( .A1(n13633), .A2(n13634), .ZN(n13632) );
  NAND2_X1 U13017 ( .A1(n13628), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10355) );
  NAND2_X1 U13018 ( .A1(n13632), .A2(n10355), .ZN(n15411) );
  INV_X1 U13019 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n10356) );
  MUX2_X1 U13020 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10356), .S(n10369), .Z(
        n15412) );
  NAND2_X1 U13021 ( .A1(n15411), .A2(n15412), .ZN(n15410) );
  NAND2_X1 U13022 ( .A1(n10369), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n10357) );
  NAND2_X1 U13023 ( .A1(n15410), .A2(n10357), .ZN(n10359) );
  INV_X1 U13024 ( .A(n10946), .ZN(n10358) );
  AOI21_X1 U13025 ( .B1(n10360), .B2(n10359), .A(n10358), .ZN(n10374) );
  INV_X1 U13026 ( .A(n15486), .ZN(n15448) );
  INV_X1 U13027 ( .A(n10944), .ZN(n10954) );
  NAND2_X1 U13028 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n12160) );
  OAI21_X1 U13029 ( .B1(n15500), .B2(n7632), .A(n12160), .ZN(n10361) );
  AOI21_X1 U13030 ( .B1(n10954), .B2(n7441), .A(n10361), .ZN(n10373) );
  XNOR2_X1 U13031 ( .A(n10944), .B(P2_REG1_REG_9__SCAN_IN), .ZN(n10370) );
  NAND2_X1 U13032 ( .A1(n10362), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10363) );
  NAND2_X1 U13033 ( .A1(n10364), .A2(n10363), .ZN(n13620) );
  XNOR2_X1 U13034 ( .A(n13615), .B(n10365), .ZN(n13621) );
  NAND2_X1 U13035 ( .A1(n13620), .A2(n13621), .ZN(n13619) );
  NAND2_X1 U13036 ( .A1(n13615), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10366) );
  NAND2_X1 U13037 ( .A1(n13619), .A2(n10366), .ZN(n13630) );
  MUX2_X1 U13038 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8133), .S(n13628), .Z(
        n13631) );
  NAND2_X1 U13039 ( .A1(n13628), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10367) );
  XNOR2_X1 U13040 ( .A(n10369), .B(n10368), .ZN(n15409) );
  OAI21_X1 U13041 ( .B1(n10370), .B2(n6647), .A(n10953), .ZN(n10371) );
  NAND2_X1 U13042 ( .A1(n10371), .A2(n15460), .ZN(n10372) );
  OAI211_X1 U13043 ( .C1(n10374), .C2(n15448), .A(n10373), .B(n10372), .ZN(
        P2_U3223) );
  INV_X1 U13044 ( .A(n13296), .ZN(n10375) );
  NAND2_X1 U13045 ( .A1(n13293), .A2(n10375), .ZN(n10376) );
  NAND2_X1 U13046 ( .A1(n10376), .A2(n12142), .ZN(n13539) );
  NOR2_X1 U13047 ( .A1(n13539), .A2(n13285), .ZN(n10380) );
  OR2_X1 U13048 ( .A1(n13539), .A2(n10377), .ZN(n10379) );
  OR2_X1 U13049 ( .A1(n8651), .A2(n13274), .ZN(n10378) );
  NAND2_X1 U13050 ( .A1(n10379), .A2(n10378), .ZN(n10886) );
  AOI211_X1 U13051 ( .C1(n10884), .C2(n13296), .A(n10380), .B(n10886), .ZN(
        n10513) );
  NAND2_X1 U13052 ( .A1(n15536), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n10381) );
  OAI21_X1 U13053 ( .B1(n15536), .B2(n10513), .A(n10381), .ZN(P2_U3499) );
  INV_X1 U13054 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n10742) );
  NAND2_X1 U13055 ( .A1(n10383), .A2(n10410), .ZN(n10617) );
  INV_X1 U13056 ( .A(n10384), .ZN(n10517) );
  NAND2_X1 U13057 ( .A1(n10516), .A2(n10517), .ZN(n10619) );
  NAND2_X1 U13058 ( .A1(n10619), .A2(n10617), .ZN(n10389) );
  MUX2_X1 U13059 ( .A(n10400), .B(n9516), .S(n13085), .Z(n10386) );
  INV_X1 U13060 ( .A(n10634), .ZN(n10385) );
  NAND2_X1 U13061 ( .A1(n10386), .A2(n10385), .ZN(n10672) );
  INV_X1 U13062 ( .A(n10386), .ZN(n10387) );
  NAND2_X1 U13063 ( .A1(n10387), .A2(n10634), .ZN(n10388) );
  AND2_X1 U13064 ( .A1(n10672), .A2(n10388), .ZN(n10616) );
  NAND2_X1 U13065 ( .A1(n10389), .A2(n10616), .ZN(n10673) );
  NAND2_X1 U13066 ( .A1(n10673), .A2(n10672), .ZN(n10394) );
  MUX2_X1 U13067 ( .A(n7597), .B(n10390), .S(n13085), .Z(n10391) );
  INV_X1 U13068 ( .A(n10680), .ZN(n10414) );
  NAND2_X1 U13069 ( .A1(n10391), .A2(n10414), .ZN(n10395) );
  INV_X1 U13070 ( .A(n10391), .ZN(n10392) );
  NAND2_X1 U13071 ( .A1(n10392), .A2(n10680), .ZN(n10393) );
  AND2_X1 U13072 ( .A1(n10395), .A2(n10393), .ZN(n10670) );
  NAND2_X1 U13073 ( .A1(n10394), .A2(n10670), .ZN(n10675) );
  NAND2_X1 U13074 ( .A1(n10675), .A2(n10395), .ZN(n10397) );
  MUX2_X1 U13075 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n13085), .Z(n10433) );
  INV_X1 U13076 ( .A(n10443), .ZN(n10434) );
  XNOR2_X1 U13077 ( .A(n10433), .B(n10434), .ZN(n10396) );
  NAND2_X1 U13078 ( .A1(n10397), .A2(n10396), .ZN(n10437) );
  OAI21_X1 U13079 ( .B1(n10397), .B2(n10396), .A(n10437), .ZN(n10427) );
  INV_X1 U13080 ( .A(n10398), .ZN(n10399) );
  NAND2_X1 U13081 ( .A1(n10514), .A2(n10399), .ZN(n10625) );
  XNOR2_X1 U13082 ( .A(n10634), .B(n10400), .ZN(n10626) );
  NAND2_X1 U13083 ( .A1(n10634), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n10401) );
  OR2_X1 U13084 ( .A1(n10402), .A2(n10680), .ZN(n10403) );
  INV_X1 U13085 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10404) );
  XNOR2_X1 U13086 ( .A(n10443), .B(n10404), .ZN(n10405) );
  INV_X1 U13087 ( .A(n10405), .ZN(n10407) );
  NAND3_X1 U13088 ( .A1(n10663), .A2(n10407), .A3(n10406), .ZN(n10408) );
  AND2_X1 U13089 ( .A1(n10445), .A2(n10408), .ZN(n10424) );
  MUX2_X1 U13090 ( .A(P3_REG1_REG_4__SCAN_IN), .B(n15657), .S(n10443), .Z(
        n10419) );
  NOR2_X1 U13091 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10409), .ZN(n10411) );
  NAND2_X1 U13092 ( .A1(n10522), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10521) );
  INV_X1 U13093 ( .A(n10411), .ZN(n10412) );
  NAND2_X1 U13094 ( .A1(n10521), .A2(n10412), .ZN(n10628) );
  XNOR2_X1 U13095 ( .A(n10634), .B(n9516), .ZN(n10629) );
  NAND2_X1 U13096 ( .A1(n10628), .A2(n10629), .ZN(n10627) );
  NAND2_X1 U13097 ( .A1(n10634), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U13098 ( .A1(n10665), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10417) );
  NAND2_X1 U13099 ( .A1(n10415), .A2(n10680), .ZN(n10416) );
  NAND2_X1 U13100 ( .A1(n10417), .A2(n10416), .ZN(n10418) );
  OAI21_X1 U13101 ( .B1(n10419), .B2(n10418), .A(n10430), .ZN(n10420) );
  NAND2_X1 U13102 ( .A1(n15591), .A2(n10420), .ZN(n10423) );
  AND2_X1 U13103 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10421) );
  AOI21_X1 U13104 ( .B1(n15539), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10421), .ZN(
        n10422) );
  OAI211_X1 U13105 ( .C1(n10424), .C2(n15570), .A(n10423), .B(n10422), .ZN(
        n10426) );
  NOR2_X1 U13106 ( .A1(n15549), .A2(n10443), .ZN(n10425) );
  AOI211_X1 U13107 ( .C1(n15595), .C2(n10427), .A(n10426), .B(n10425), .ZN(
        n10428) );
  INV_X1 U13108 ( .A(n10428), .ZN(P3_U3186) );
  NAND2_X1 U13109 ( .A1(n10443), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10429) );
  INV_X1 U13110 ( .A(n10682), .ZN(n10431) );
  XOR2_X1 U13111 ( .A(n10681), .B(P3_REG1_REG_5__SCAN_IN), .Z(n10454) );
  MUX2_X1 U13112 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n13085), .Z(n10438) );
  INV_X1 U13113 ( .A(n10438), .ZN(n10432) );
  NAND2_X1 U13114 ( .A1(n10432), .A2(n10431), .ZN(n10688) );
  INV_X1 U13115 ( .A(n10433), .ZN(n10435) );
  NAND2_X1 U13116 ( .A1(n10435), .A2(n10434), .ZN(n10436) );
  NAND2_X1 U13117 ( .A1(n10437), .A2(n10436), .ZN(n10439) );
  NAND2_X1 U13118 ( .A1(n10438), .A2(n10682), .ZN(n10440) );
  AOI21_X1 U13119 ( .B1(n10440), .B2(n10688), .A(n10439), .ZN(n10441) );
  INV_X1 U13120 ( .A(n10441), .ZN(n10442) );
  OAI21_X1 U13121 ( .B1(n7372), .B2(n10689), .A(n10442), .ZN(n10452) );
  AND2_X1 U13122 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10804) );
  AOI21_X1 U13123 ( .B1(n15539), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10804), .ZN(
        n10450) );
  NAND2_X1 U13124 ( .A1(n10443), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n10444) );
  NAND2_X1 U13125 ( .A1(n10446), .A2(n10682), .ZN(n15543) );
  OAI21_X1 U13126 ( .B1(P3_REG2_REG_5__SCAN_IN), .B2(n6644), .A(n15547), .ZN(
        n10448) );
  NAND2_X1 U13127 ( .A1(n15586), .A2(n10448), .ZN(n10449) );
  OAI211_X1 U13128 ( .C1(n15549), .C2(n10682), .A(n10450), .B(n10449), .ZN(
        n10451) );
  AOI21_X1 U13129 ( .B1(n10452), .B2(n15595), .A(n10451), .ZN(n10453) );
  OAI21_X1 U13130 ( .B1(n10454), .B2(n12730), .A(n10453), .ZN(P3_U3187) );
  INV_X1 U13131 ( .A(n10455), .ZN(n10493) );
  INV_X1 U13132 ( .A(n15189), .ZN(n15186) );
  AOI22_X1 U13133 ( .A1(n11377), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n15186), .ZN(n10456) );
  OAI21_X1 U13134 ( .B1(n10493), .B2(n15195), .A(n10456), .ZN(P1_U3342) );
  INV_X1 U13135 ( .A(n10457), .ZN(n10463) );
  INV_X1 U13136 ( .A(n11751), .ZN(n10952) );
  OAI222_X1 U13137 ( .A1(n14102), .A2(n10458), .B1(n14099), .B2(n10463), .C1(
        P2_U3088), .C2(n10952), .ZN(P2_U3316) );
  INV_X1 U13138 ( .A(n12396), .ZN(n10459) );
  NAND2_X1 U13139 ( .A1(n10535), .A2(n15626), .ZN(n10460) );
  OAI22_X1 U13140 ( .A1(n12525), .A2(n10460), .B1(n7152), .B2(n12838), .ZN(
        n10754) );
  NOR2_X1 U13141 ( .A1(n15665), .A2(n10127), .ZN(n10461) );
  AOI21_X1 U13142 ( .B1(n15665), .B2(n10754), .A(n10461), .ZN(n10462) );
  OAI21_X1 U13143 ( .B1(n10756), .B2(n12976), .A(n10462), .ZN(P3_U3459) );
  INV_X1 U13144 ( .A(n14679), .ZN(n10845) );
  OAI222_X1 U13145 ( .A1(n10464), .A2(n15189), .B1(P1_U3086), .B2(n10845), 
        .C1(n15195), .C2(n10463), .ZN(P1_U3344) );
  NAND2_X1 U13146 ( .A1(n10481), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n10465) );
  XNOR2_X1 U13147 ( .A(n14636), .B(n10467), .ZN(n14642) );
  NAND2_X1 U13148 ( .A1(n14641), .A2(n14642), .ZN(n14640) );
  NAND2_X1 U13149 ( .A1(n14636), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n10468) );
  AND2_X1 U13150 ( .A1(n14640), .A2(n10468), .ZN(n14651) );
  MUX2_X1 U13151 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10469), .S(n14648), .Z(
        n14650) );
  NAND2_X1 U13152 ( .A1(n14651), .A2(n14650), .ZN(n14649) );
  OR2_X1 U13153 ( .A1(n14648), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U13154 ( .A1(n14649), .A2(n10470), .ZN(n14660) );
  MUX2_X1 U13155 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10471), .S(n14666), .Z(
        n14661) );
  NAND2_X1 U13156 ( .A1(n14660), .A2(n14661), .ZN(n14659) );
  NAND2_X1 U13157 ( .A1(n10472), .A2(n10471), .ZN(n10473) );
  NAND2_X1 U13158 ( .A1(n14659), .A2(n10473), .ZN(n10476) );
  INV_X1 U13159 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10474) );
  MUX2_X1 U13160 ( .A(n10474), .B(P1_REG1_REG_10__SCAN_IN), .S(n10841), .Z(
        n10475) );
  AOI21_X1 U13161 ( .B1(n10476), .B2(n10475), .A(n14733), .ZN(n10480) );
  NAND2_X1 U13162 ( .A1(n14735), .A2(n10841), .ZN(n10478) );
  NAND2_X1 U13163 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10477)
         );
  OAI211_X1 U13164 ( .C1(n14742), .C2(n15774), .A(n10478), .B(n10477), .ZN(
        n10479) );
  AOI21_X1 U13165 ( .B1(n10480), .B2(n10843), .A(n10479), .ZN(n10491) );
  NAND2_X1 U13166 ( .A1(n10481), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U13167 ( .A1(n10483), .A2(n10482), .ZN(n14638) );
  INV_X1 U13168 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n11417) );
  XNOR2_X1 U13169 ( .A(n14636), .B(n11417), .ZN(n14639) );
  NAND2_X1 U13170 ( .A1(n14638), .A2(n14639), .ZN(n14637) );
  NAND2_X1 U13171 ( .A1(n14636), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n10484) );
  NAND2_X1 U13172 ( .A1(n14637), .A2(n10484), .ZN(n14654) );
  INV_X1 U13173 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10485) );
  MUX2_X1 U13174 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10485), .S(n14648), .Z(
        n14655) );
  NAND2_X1 U13175 ( .A1(n14654), .A2(n14655), .ZN(n14653) );
  NAND2_X1 U13176 ( .A1(n14648), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10486) );
  NAND2_X1 U13177 ( .A1(n14653), .A2(n10486), .ZN(n14669) );
  INV_X1 U13178 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n11532) );
  XNOR2_X1 U13179 ( .A(n14666), .B(n11532), .ZN(n14668) );
  NAND2_X1 U13180 ( .A1(n14669), .A2(n14668), .ZN(n14667) );
  NAND2_X1 U13181 ( .A1(n14666), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n10487) );
  NAND2_X1 U13182 ( .A1(n14667), .A2(n10487), .ZN(n10489) );
  INV_X1 U13183 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11544) );
  XNOR2_X1 U13184 ( .A(n10841), .B(n11544), .ZN(n10488) );
  NAND2_X1 U13185 ( .A1(n10489), .A2(n10488), .ZN(n10834) );
  OAI211_X1 U13186 ( .C1(n10489), .C2(n10488), .A(n10834), .B(n14737), .ZN(
        n10490) );
  NAND2_X1 U13187 ( .A1(n10491), .A2(n10490), .ZN(P1_U3253) );
  INV_X1 U13188 ( .A(n15456), .ZN(n10492) );
  OAI222_X1 U13189 ( .A1(n14102), .A2(n10494), .B1(n14099), .B2(n10493), .C1(
        n10492), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U13190 ( .A(n10495), .ZN(n10496) );
  OAI222_X1 U13191 ( .A1(P3_U3151), .A2(n12641), .B1(n13095), .B2(n10497), 
        .C1(n13090), .C2(n10496), .ZN(P3_U3281) );
  INV_X1 U13192 ( .A(n11305), .ZN(n10850) );
  INV_X1 U13193 ( .A(n10498), .ZN(n10499) );
  OAI222_X1 U13194 ( .A1(P1_U3086), .A2(n10850), .B1(n15192), .B2(n10499), 
        .C1(n15769), .C2(n15189), .ZN(P1_U3343) );
  INV_X1 U13195 ( .A(n11754), .ZN(n15433) );
  OAI222_X1 U13196 ( .A1(n14102), .A2(n10500), .B1(n14099), .B2(n10499), .C1(
        n15433), .C2(P2_U3088), .ZN(P2_U3315) );
  INV_X1 U13197 ( .A(n10504), .ZN(n10501) );
  OR2_X1 U13198 ( .A1(n10502), .A2(n10501), .ZN(n10503) );
  OAI21_X1 U13199 ( .B1(n10578), .B2(n10504), .A(n10503), .ZN(n10506) );
  NAND4_X1 U13200 ( .A1(n10507), .A2(n10506), .A3(n10505), .A4(n10529), .ZN(
        n10509) );
  INV_X1 U13201 ( .A(n12521), .ZN(n15608) );
  NOR2_X1 U13202 ( .A1(n15626), .A2(n12521), .ZN(n10508) );
  AOI21_X1 U13203 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n12912), .A(n10754), .ZN(
        n10510) );
  MUX2_X1 U13204 ( .A(n7410), .B(n10510), .S(n15616), .Z(n10511) );
  OAI21_X1 U13205 ( .B1(n10756), .B2(n12828), .A(n10511), .ZN(P3_U3233) );
  OR2_X1 U13206 ( .A1(n15533), .A2(n8022), .ZN(n10512) );
  OAI21_X1 U13207 ( .B1(n15531), .B2(n10513), .A(n10512), .ZN(P2_U3430) );
  OAI21_X1 U13208 ( .B1(P3_REG2_REG_1__SCAN_IN), .B2(n10515), .A(n10514), .ZN(
        n10526) );
  OAI21_X1 U13209 ( .B1(n10517), .B2(n10516), .A(n10619), .ZN(n10518) );
  NAND2_X1 U13210 ( .A1(n15595), .A2(n10518), .ZN(n10520) );
  NAND2_X1 U13211 ( .A1(n15539), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n10519) );
  OAI211_X1 U13212 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n10595), .A(n10520), .B(
        n10519), .ZN(n10525) );
  OAI21_X1 U13213 ( .B1(P3_REG1_REG_1__SCAN_IN), .B2(n10522), .A(n10521), .ZN(
        n10523) );
  AND2_X1 U13214 ( .A1(n15591), .A2(n10523), .ZN(n10524) );
  AOI211_X1 U13215 ( .C1(n15586), .C2(n10526), .A(n10525), .B(n10524), .ZN(
        n10527) );
  OAI21_X1 U13216 ( .B1(n10528), .B2(n15549), .A(n10527), .ZN(P3_U3183) );
  INV_X1 U13217 ( .A(n10540), .ZN(n10549) );
  NAND2_X1 U13218 ( .A1(n10545), .A2(n10539), .ZN(n10533) );
  AND3_X1 U13219 ( .A1(n10531), .A2(n10530), .A3(n10529), .ZN(n10532) );
  OAI211_X1 U13220 ( .C1(n10549), .C2(n10541), .A(n10533), .B(n10532), .ZN(
        n10534) );
  NAND2_X1 U13221 ( .A1(n10534), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10538) );
  NOR2_X1 U13222 ( .A1(n10548), .A2(n10535), .ZN(n10536) );
  NAND2_X1 U13223 ( .A1(n10540), .A2(n10536), .ZN(n10537) );
  NOR2_X1 U13224 ( .A1(n12340), .A2(P3_U3151), .ZN(n10604) );
  NAND2_X1 U13225 ( .A1(n10539), .A2(n15626), .ZN(n10542) );
  OAI22_X1 U13226 ( .A1(n10545), .A2(n10542), .B1(n10541), .B2(n10540), .ZN(
        n10544) );
  INV_X1 U13227 ( .A(n12525), .ZN(n10551) );
  NAND2_X1 U13228 ( .A1(n10545), .A2(n12521), .ZN(n10547) );
  NOR2_X1 U13229 ( .A1(n10548), .A2(n15626), .ZN(n10546) );
  NOR2_X1 U13230 ( .A1(n10548), .A2(n12522), .ZN(n12557) );
  NAND2_X1 U13231 ( .A1(n10549), .A2(n12557), .ZN(n12313) );
  INV_X1 U13232 ( .A(n12313), .ZN(n12324) );
  NAND2_X1 U13233 ( .A1(n12324), .A2(n12981), .ZN(n12344) );
  OAI22_X1 U13234 ( .A1(n12285), .A2(n10756), .B1(n12344), .B2(n7152), .ZN(
        n10550) );
  AOI21_X1 U13235 ( .B1(n12308), .B2(n10551), .A(n10550), .ZN(n10552) );
  OAI21_X1 U13236 ( .B1(n10604), .B2(n10553), .A(n10552), .ZN(P3_U3172) );
  NOR2_X1 U13237 ( .A1(n8651), .A2(n6406), .ZN(n13238) );
  XNOR2_X1 U13238 ( .A(n10717), .B(n7216), .ZN(n13237) );
  XNOR2_X1 U13239 ( .A(n13238), .B(n13237), .ZN(n10572) );
  INV_X1 U13240 ( .A(n10572), .ZN(n10558) );
  OR2_X1 U13241 ( .A1(n10717), .A2(n13296), .ZN(n10711) );
  INV_X1 U13242 ( .A(n10711), .ZN(n10557) );
  INV_X1 U13243 ( .A(n12142), .ZN(n10555) );
  INV_X1 U13244 ( .A(n10709), .ZN(n10556) );
  NAND2_X1 U13245 ( .A1(n10572), .A2(n10556), .ZN(n13233) );
  INV_X1 U13246 ( .A(n13233), .ZN(n13243) );
  AOI21_X1 U13247 ( .B1(n10558), .B2(n10557), .A(n13243), .ZN(n10576) );
  AND2_X1 U13248 ( .A1(n10559), .A2(n15507), .ZN(n10560) );
  NOR2_X1 U13249 ( .A1(n15524), .A2(n10563), .ZN(n10564) );
  INV_X2 U13250 ( .A(n13270), .ZN(n13250) );
  NAND2_X1 U13251 ( .A1(n10567), .A2(n10565), .ZN(n10566) );
  INV_X1 U13252 ( .A(n13570), .ZN(n13574) );
  AOI22_X1 U13253 ( .A1(n13878), .A2(n13612), .B1(n13610), .B2(n13880), .ZN(
        n12154) );
  OAI21_X1 U13254 ( .B1(n15506), .B2(n10569), .A(n10568), .ZN(n10571) );
  NAND2_X1 U13255 ( .A1(n10571), .A2(n10570), .ZN(n10726) );
  NOR2_X1 U13256 ( .A1(n10726), .A2(n15509), .ZN(n13235) );
  OAI22_X1 U13257 ( .A1(n13263), .A2(n12154), .B1(n13235), .B2(n6948), .ZN(
        n10574) );
  NAND2_X1 U13258 ( .A1(n13270), .A2(n6409), .ZN(n13256) );
  NOR3_X1 U13259 ( .A1(n13256), .A2(n12142), .A3(n10572), .ZN(n10573) );
  AOI211_X1 U13260 ( .C1(n13916), .C2(n13280), .A(n10574), .B(n10573), .ZN(
        n10575) );
  OAI21_X1 U13261 ( .B1(n10576), .B2(n13250), .A(n10575), .ZN(P2_U3194) );
  NOR2_X2 U13262 ( .A1(n12313), .A2(n12836), .ZN(n12341) );
  INV_X1 U13263 ( .A(n12583), .ZN(n10643) );
  OAI22_X1 U13264 ( .A1(n12285), .A2(n10736), .B1(n12344), .B2(n10643), .ZN(
        n10577) );
  AOI21_X1 U13265 ( .B1(n12341), .B2(n12584), .A(n10577), .ZN(n10594) );
  NAND2_X1 U13266 ( .A1(n12548), .A2(n11461), .ZN(n10579) );
  NAND2_X1 U13267 ( .A1(n10579), .A2(n11334), .ZN(n10580) );
  NAND3_X1 U13268 ( .A1(n12220), .A2(n9514), .A3(n7151), .ZN(n10585) );
  AND2_X1 U13269 ( .A1(n10585), .A2(n10596), .ZN(n10591) );
  INV_X1 U13270 ( .A(n10737), .ZN(n10587) );
  OAI21_X1 U13271 ( .B1(n6445), .B2(n10587), .A(n10586), .ZN(n10588) );
  NAND2_X1 U13272 ( .A1(n10591), .A2(n10588), .ZN(n10597) );
  NAND3_X1 U13273 ( .A1(n12399), .A2(n10589), .A3(n6445), .ZN(n10590) );
  OAI211_X1 U13274 ( .C1(n10591), .C2(n10737), .A(n10597), .B(n10590), .ZN(
        n10592) );
  NAND2_X1 U13275 ( .A1(n10592), .A2(n12308), .ZN(n10593) );
  OAI211_X1 U13276 ( .C1(n10604), .C2(n10595), .A(n10594), .B(n10593), .ZN(
        P3_U3162) );
  XNOR2_X1 U13277 ( .A(n6446), .B(n7169), .ZN(n10638) );
  XNOR2_X1 U13278 ( .A(n10638), .B(n12583), .ZN(n10599) );
  NAND2_X1 U13279 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  OAI21_X1 U13280 ( .B1(n10599), .B2(n10598), .A(n10642), .ZN(n10600) );
  NAND2_X1 U13281 ( .A1(n10600), .A2(n12308), .ZN(n10603) );
  OAI22_X1 U13282 ( .A1(n12285), .A2(n12990), .B1(n12344), .B2(n6411), .ZN(
        n10601) );
  AOI21_X1 U13283 ( .B1(n12341), .B2(n9514), .A(n10601), .ZN(n10602) );
  OAI211_X1 U13284 ( .C1(n10604), .C2(n15609), .A(n10603), .B(n10602), .ZN(
        P3_U3177) );
  INV_X1 U13285 ( .A(n10606), .ZN(n10607) );
  AOI21_X1 U13286 ( .B1(n10609), .B2(n10608), .A(n10607), .ZN(n10615) );
  INV_X1 U13287 ( .A(n10760), .ZN(n10612) );
  AOI22_X1 U13288 ( .A1(n14209), .A2(n14557), .B1(n14264), .B2(n14558), .ZN(
        n10610) );
  OAI21_X1 U13289 ( .B1(n10612), .B2(n10611), .A(n10610), .ZN(n10613) );
  AOI21_X1 U13290 ( .B1(n14269), .B2(n14295), .A(n10613), .ZN(n10614) );
  OAI21_X1 U13291 ( .B1(n10615), .B2(n14271), .A(n10614), .ZN(P1_U3222) );
  INV_X1 U13292 ( .A(n10616), .ZN(n10618) );
  NAND3_X1 U13293 ( .A1(n10619), .A2(n10618), .A3(n10617), .ZN(n10620) );
  AOI21_X1 U13294 ( .B1(n10673), .B2(n10620), .A(n15576), .ZN(n10623) );
  OAI22_X1 U13295 ( .A1(n15605), .A2(n10621), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15609), .ZN(n10622) );
  NOR2_X1 U13296 ( .A1(n10623), .A2(n10622), .ZN(n10633) );
  OAI21_X1 U13297 ( .B1(n10626), .B2(n10625), .A(n10624), .ZN(n10631) );
  OAI21_X1 U13298 ( .B1(n10629), .B2(n10628), .A(n10627), .ZN(n10630) );
  AOI22_X1 U13299 ( .A1(n15586), .A2(n10631), .B1(n15591), .B2(n10630), .ZN(
        n10632) );
  OAI211_X1 U13300 ( .C1(n10634), .C2(n15549), .A(n10633), .B(n10632), .ZN(
        P3_U3184) );
  INV_X1 U13301 ( .A(n12661), .ZN(n12683) );
  INV_X1 U13302 ( .A(n10635), .ZN(n10636) );
  OAI222_X1 U13303 ( .A1(P3_U3151), .A2(n12683), .B1(n13095), .B2(n10637), 
        .C1(n13090), .C2(n10636), .ZN(P3_U3280) );
  NAND2_X1 U13304 ( .A1(n10638), .A2(n10643), .ZN(n10639) );
  XNOR2_X1 U13305 ( .A(n10649), .B(n12980), .ZN(n10640) );
  AOI21_X1 U13306 ( .B1(n10642), .B2(n10639), .A(n10640), .ZN(n10648) );
  AND2_X1 U13307 ( .A1(n10640), .A2(n10639), .ZN(n10641) );
  NAND2_X1 U13308 ( .A1(n10652), .A2(n12308), .ZN(n10647) );
  OAI22_X1 U13309 ( .A1(n12285), .A2(n10789), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n9535), .ZN(n10645) );
  INV_X1 U13310 ( .A(n12341), .ZN(n12292) );
  INV_X1 U13311 ( .A(n12582), .ZN(n10980) );
  OAI22_X1 U13312 ( .A1(n12292), .A2(n10643), .B1(n10980), .B2(n12344), .ZN(
        n10644) );
  AOI211_X1 U13313 ( .C1(n9535), .C2(n12340), .A(n10645), .B(n10644), .ZN(
        n10646) );
  OAI21_X1 U13314 ( .B1(n10648), .B2(n10647), .A(n10646), .ZN(P3_U3158) );
  INV_X1 U13315 ( .A(n10649), .ZN(n10650) );
  NAND2_X1 U13316 ( .A1(n10650), .A2(n12980), .ZN(n10651) );
  INV_X1 U13317 ( .A(n10857), .ZN(n10655) );
  INV_X1 U13318 ( .A(n10653), .ZN(n10654) );
  NAND2_X1 U13319 ( .A1(n10654), .A2(n12582), .ZN(n10856) );
  NAND2_X1 U13320 ( .A1(n10655), .A2(n10856), .ZN(n10656) );
  NOR2_X1 U13321 ( .A1(n10863), .A2(n10656), .ZN(n10800) );
  AOI21_X1 U13322 ( .B1(n10863), .B2(n10656), .A(n10800), .ZN(n10662) );
  INV_X1 U13323 ( .A(n10774), .ZN(n10660) );
  OAI22_X1 U13324 ( .A1(n12285), .A2(n15627), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n10657), .ZN(n10659) );
  INV_X1 U13325 ( .A(n12581), .ZN(n10996) );
  OAI22_X1 U13326 ( .A1(n12292), .A2(n6411), .B1(n10996), .B2(n12344), .ZN(
        n10658) );
  AOI211_X1 U13327 ( .C1(n10660), .C2(n12340), .A(n10659), .B(n10658), .ZN(
        n10661) );
  OAI21_X1 U13328 ( .B1(n10662), .B2(n12349), .A(n10661), .ZN(P3_U3170) );
  OAI21_X1 U13329 ( .B1(P3_REG2_REG_3__SCAN_IN), .B2(n10664), .A(n10663), .ZN(
        n10678) );
  XNOR2_X1 U13330 ( .A(n10665), .B(P3_REG1_REG_3__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13331 ( .A1(n15591), .A2(n10666), .ZN(n10669) );
  NOR2_X1 U13332 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n9535), .ZN(n10667) );
  AOI21_X1 U13333 ( .B1(n15539), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10667), .ZN(
        n10668) );
  NAND2_X1 U13334 ( .A1(n10669), .A2(n10668), .ZN(n10677) );
  INV_X1 U13335 ( .A(n10670), .ZN(n10671) );
  NAND3_X1 U13336 ( .A1(n10673), .A2(n10672), .A3(n10671), .ZN(n10674) );
  AOI21_X1 U13337 ( .B1(n10675), .B2(n10674), .A(n15576), .ZN(n10676) );
  AOI211_X1 U13338 ( .C1(n15586), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10679) );
  OAI21_X1 U13339 ( .B1(n10680), .B2(n15549), .A(n10679), .ZN(P3_U3185) );
  NAND2_X1 U13340 ( .A1(n10683), .A2(n10682), .ZN(n10684) );
  NAND2_X1 U13341 ( .A1(n10685), .A2(n10684), .ZN(n15541) );
  MUX2_X1 U13342 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10686), .S(n15550), .Z(
        n15542) );
  NAND2_X1 U13343 ( .A1(n15550), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10687) );
  XOR2_X1 U13344 ( .A(n11218), .B(P3_REG1_REG_7__SCAN_IN), .Z(n10703) );
  MUX2_X1 U13345 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n7168), .Z(n10690) );
  INV_X1 U13346 ( .A(n15550), .ZN(n10691) );
  XNOR2_X1 U13347 ( .A(n10690), .B(n10691), .ZN(n15553) );
  INV_X1 U13348 ( .A(n10690), .ZN(n10692) );
  MUX2_X1 U13349 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n7168), .Z(n11227) );
  XNOR2_X1 U13350 ( .A(n11227), .B(n11228), .ZN(n11225) );
  XNOR2_X1 U13351 ( .A(n11226), .B(n11225), .ZN(n10701) );
  INV_X1 U13352 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n10970) );
  XNOR2_X1 U13353 ( .A(n15550), .B(n10970), .ZN(n15544) );
  NAND2_X1 U13354 ( .A1(n15550), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10693) );
  OAI21_X1 U13355 ( .B1(P3_REG2_REG_7__SCAN_IN), .B2(n10695), .A(n15569), .ZN(
        n10696) );
  NAND2_X1 U13356 ( .A1(n10696), .A2(n15586), .ZN(n10699) );
  NAND2_X1 U13357 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11070) );
  INV_X1 U13358 ( .A(n11070), .ZN(n10697) );
  AOI21_X1 U13359 ( .B1(n15539), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n10697), .ZN(
        n10698) );
  OAI211_X1 U13360 ( .C1(n15549), .C2(n11219), .A(n10699), .B(n10698), .ZN(
        n10700) );
  AOI21_X1 U13361 ( .B1(n15595), .B2(n10701), .A(n10700), .ZN(n10702) );
  OAI21_X1 U13362 ( .B1(n10703), .B2(n12730), .A(n10702), .ZN(P3_U3189) );
  INV_X1 U13363 ( .A(n13256), .ZN(n13269) );
  NAND2_X1 U13364 ( .A1(n13269), .A2(n13612), .ZN(n10706) );
  AOI21_X1 U13365 ( .B1(n13612), .B2(n6409), .A(n13250), .ZN(n10704) );
  NOR2_X1 U13366 ( .A1(n10704), .A2(n13280), .ZN(n10705) );
  MUX2_X1 U13367 ( .A(n10706), .B(n10705), .S(n13296), .Z(n10708) );
  AND2_X1 U13368 ( .A1(n13275), .A2(n13880), .ZN(n13229) );
  OAI211_X1 U13369 ( .C1(n13235), .C2(n10887), .A(n10708), .B(n10707), .ZN(
        P2_U3204) );
  NOR2_X1 U13370 ( .A1(n13304), .A2(n6405), .ZN(n13232) );
  INV_X1 U13371 ( .A(n13238), .ZN(n10712) );
  XNOR2_X1 U13372 ( .A(n13286), .B(n10717), .ZN(n10713) );
  AND2_X1 U13373 ( .A1(n13609), .A2(n6409), .ZN(n10714) );
  NAND2_X1 U13374 ( .A1(n10713), .A2(n10714), .ZN(n10718) );
  INV_X1 U13375 ( .A(n10713), .ZN(n13191) );
  INV_X1 U13376 ( .A(n10714), .ZN(n10715) );
  NAND2_X1 U13377 ( .A1(n13191), .A2(n10715), .ZN(n10716) );
  NAND2_X1 U13378 ( .A1(n10718), .A2(n10716), .ZN(n11043) );
  NAND2_X1 U13379 ( .A1(n13608), .A2(n6409), .ZN(n10720) );
  INV_X1 U13380 ( .A(n10719), .ZN(n10730) );
  NAND2_X1 U13381 ( .A1(n10730), .A2(n10720), .ZN(n10721) );
  XNOR2_X1 U13382 ( .A(n13328), .B(n13139), .ZN(n11112) );
  NOR2_X1 U13383 ( .A1(n13330), .A2(n6406), .ZN(n11113) );
  INV_X1 U13384 ( .A(n11113), .ZN(n10933) );
  XNOR2_X1 U13385 ( .A(n11112), .B(n10933), .ZN(n10731) );
  NAND2_X1 U13386 ( .A1(n11118), .A2(n10731), .ZN(n10935) );
  AND2_X1 U13387 ( .A1(n13275), .A2(n13878), .ZN(n13230) );
  OAI21_X1 U13388 ( .B1(n13227), .B2(n11191), .A(n10722), .ZN(n10729) );
  INV_X1 U13389 ( .A(n13229), .ZN(n13198) );
  INV_X1 U13390 ( .A(n10723), .ZN(n10725) );
  OR3_X1 U13391 ( .A1(n10726), .A2(n10725), .A3(n10724), .ZN(n10727) );
  OAI22_X1 U13392 ( .A1(n13198), .A2(n11182), .B1(n13277), .B2(n11194), .ZN(
        n10728) );
  AOI211_X1 U13393 ( .C1(n13230), .C2(n13608), .A(n10729), .B(n10728), .ZN(
        n10735) );
  OAI22_X1 U13394 ( .A1(n11183), .A2(n13256), .B1(n13250), .B2(n10730), .ZN(
        n10733) );
  INV_X1 U13395 ( .A(n10731), .ZN(n10732) );
  NAND3_X1 U13396 ( .A1(n10733), .A2(n10732), .A3(n13187), .ZN(n10734) );
  OAI211_X1 U13397 ( .C1(n10935), .C2(n13250), .A(n10735), .B(n10734), .ZN(
        P2_U3199) );
  NOR2_X1 U13398 ( .A1(n10736), .A2(n15626), .ZN(n15620) );
  INV_X1 U13399 ( .A(n12978), .ZN(n10981) );
  AOI22_X1 U13400 ( .A1(n12981), .A2(n12583), .B1(n12584), .B2(n12982), .ZN(
        n10740) );
  XNOR2_X1 U13401 ( .A(n10589), .B(n10737), .ZN(n10738) );
  NAND2_X1 U13402 ( .A1(n10738), .A2(n12986), .ZN(n10739) );
  OAI211_X1 U13403 ( .C1(n10744), .C2(n10981), .A(n10740), .B(n10739), .ZN(
        n15619) );
  AOI21_X1 U13404 ( .B1(n15620), .B2(n12521), .A(n15619), .ZN(n10741) );
  MUX2_X1 U13405 ( .A(n10742), .B(n10741), .S(n15616), .Z(n10746) );
  NOR2_X1 U13406 ( .A1(n12521), .A2(n11461), .ZN(n15615) );
  INV_X1 U13407 ( .A(n15615), .ZN(n10743) );
  NOR2_X1 U13408 ( .A1(n15618), .A2(n10743), .ZN(n12789) );
  INV_X1 U13409 ( .A(n10744), .ZN(n15621) );
  AOI22_X1 U13410 ( .A1(n12789), .A2(n15621), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n12912), .ZN(n10745) );
  NAND2_X1 U13411 ( .A1(n10746), .A2(n10745), .ZN(P3_U3232) );
  INV_X1 U13412 ( .A(n14694), .ZN(n10749) );
  INV_X1 U13413 ( .A(n10747), .ZN(n10750) );
  OAI222_X1 U13414 ( .A1(P1_U3086), .A2(n10749), .B1(n15192), .B2(n10750), 
        .C1(n10748), .C2(n15189), .ZN(P1_U3339) );
  OAI222_X1 U13415 ( .A1(n14102), .A2(n10751), .B1(n14099), .B2(n10750), .C1(
        n13643), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U13416 ( .A(n13061), .ZN(n13070) );
  INV_X1 U13417 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10752) );
  NOR2_X1 U13418 ( .A1(n15654), .A2(n10752), .ZN(n10753) );
  AOI21_X1 U13419 ( .B1(n15654), .B2(n10754), .A(n10753), .ZN(n10755) );
  OAI21_X1 U13420 ( .B1(n10756), .B2(n13070), .A(n10755), .ZN(P3_U3390) );
  OAI21_X1 U13421 ( .B1(n10758), .B2(n10757), .A(n14141), .ZN(n10759) );
  NAND2_X1 U13422 ( .A1(n10759), .A2(n14273), .ZN(n10762) );
  OAI22_X1 U13423 ( .A1(n11054), .A2(n14855), .B1(n6853), .B2(n14853), .ZN(
        n15259) );
  AOI22_X1 U13424 ( .A1(n15259), .A2(n14282), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n10760), .ZN(n10761) );
  OAI211_X1 U13425 ( .C1(n15286), .C2(n14285), .A(n10762), .B(n10761), .ZN(
        P1_U3237) );
  INV_X1 U13426 ( .A(n11627), .ZN(n10765) );
  INV_X1 U13427 ( .A(n10763), .ZN(n10766) );
  OAI222_X1 U13428 ( .A1(P1_U3086), .A2(n10765), .B1(n15192), .B2(n10766), 
        .C1(n10764), .C2(n15189), .ZN(P1_U3341) );
  INV_X1 U13429 ( .A(n13649), .ZN(n11759) );
  OAI222_X1 U13430 ( .A1(n14102), .A2(n10767), .B1(n14099), .B2(n10766), .C1(
        n11759), .C2(P2_U3088), .ZN(P2_U3313) );
  INV_X1 U13431 ( .A(n10783), .ZN(n12527) );
  AND2_X1 U13432 ( .A1(n10964), .A2(n12527), .ZN(n10786) );
  NOR2_X1 U13433 ( .A1(n10786), .A2(n10768), .ZN(n10769) );
  XNOR2_X1 U13434 ( .A(n10769), .B(n7416), .ZN(n10771) );
  AOI22_X1 U13435 ( .A1(n12981), .A2(n12581), .B1(n12980), .B2(n12982), .ZN(
        n10770) );
  OAI21_X1 U13436 ( .B1(n10771), .B2(n12834), .A(n10770), .ZN(n15628) );
  INV_X1 U13437 ( .A(n15628), .ZN(n10778) );
  XNOR2_X1 U13438 ( .A(n12414), .B(n10772), .ZN(n15631) );
  OR2_X1 U13439 ( .A1(n12978), .A2(n15615), .ZN(n10773) );
  INV_X1 U13440 ( .A(n12922), .ZN(n12845) );
  OAI22_X1 U13441 ( .A1(n15616), .A2(n10404), .B1(n10774), .B2(n15610), .ZN(
        n10776) );
  NOR2_X1 U13442 ( .A1(n12828), .A2(n15627), .ZN(n10775) );
  AOI211_X1 U13443 ( .C1(n15631), .C2(n12845), .A(n10776), .B(n10775), .ZN(
        n10777) );
  OAI21_X1 U13444 ( .B1(n10778), .B2(n15618), .A(n10777), .ZN(P3_U3229) );
  INV_X1 U13445 ( .A(n10779), .ZN(n10781) );
  OAI222_X1 U13446 ( .A1(n12701), .A2(P3_U3151), .B1(n13090), .B2(n10781), 
        .C1(n10780), .C2(n13095), .ZN(P3_U3279) );
  XNOR2_X1 U13447 ( .A(n10782), .B(n10783), .ZN(n15625) );
  INV_X1 U13448 ( .A(n15625), .ZN(n10792) );
  OAI21_X1 U13449 ( .B1(n10964), .B2(n12527), .A(n12986), .ZN(n10787) );
  NAND2_X1 U13450 ( .A1(n15625), .A2(n12978), .ZN(n10785) );
  AOI22_X1 U13451 ( .A1(n12981), .A2(n12582), .B1(n12583), .B2(n12982), .ZN(
        n10784) );
  OAI211_X1 U13452 ( .C1(n10787), .C2(n10786), .A(n10785), .B(n10784), .ZN(
        n15623) );
  MUX2_X1 U13453 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15623), .S(n15616), .Z(
        n10788) );
  INV_X1 U13454 ( .A(n10788), .ZN(n10791) );
  NOR2_X1 U13455 ( .A1(n10789), .A2(n15626), .ZN(n15624) );
  AOI22_X1 U13456 ( .A1(n12762), .A2(n15624), .B1(n12912), .B2(n9535), .ZN(
        n10790) );
  OAI211_X1 U13457 ( .C1(n10792), .C2(n11276), .A(n10791), .B(n10790), .ZN(
        P3_U3230) );
  AOI211_X1 U13458 ( .C1(n15522), .C2(n10795), .A(n10794), .B(n10793), .ZN(
        n10799) );
  NOR2_X1 U13459 ( .A1(n15533), .A2(n8059), .ZN(n10796) );
  AOI21_X1 U13460 ( .B1(n14086), .B2(n13286), .A(n10796), .ZN(n10797) );
  OAI21_X1 U13461 ( .B1(n10799), .B2(n15531), .A(n10797), .ZN(P2_U3439) );
  AOI22_X1 U13462 ( .A1(n14023), .A2(n13286), .B1(n15536), .B2(
        P2_REG1_REG_3__SCAN_IN), .ZN(n10798) );
  OAI21_X1 U13463 ( .B1(n10799), .B2(n15536), .A(n10798), .ZN(P2_U3502) );
  INV_X1 U13464 ( .A(n12340), .ZN(n12321) );
  XNOR2_X1 U13465 ( .A(n6446), .B(n10805), .ZN(n10859) );
  XNOR2_X1 U13466 ( .A(n10859), .B(n12581), .ZN(n10858) );
  OR2_X1 U13467 ( .A1(n10800), .A2(n10857), .ZN(n10801) );
  NAND2_X1 U13468 ( .A1(n10801), .A2(n10858), .ZN(n10991) );
  OAI21_X1 U13469 ( .B1(n10858), .B2(n10801), .A(n10991), .ZN(n10802) );
  NAND2_X1 U13470 ( .A1(n10802), .A2(n12308), .ZN(n10807) );
  INV_X1 U13471 ( .A(n12580), .ZN(n10979) );
  OAI22_X1 U13472 ( .A1(n12292), .A2(n10980), .B1(n10979), .B2(n12344), .ZN(
        n10803) );
  AOI211_X1 U13473 ( .C1(n12347), .C2(n10805), .A(n10804), .B(n10803), .ZN(
        n10806) );
  OAI211_X1 U13474 ( .C1(n10986), .C2(n12321), .A(n10807), .B(n10806), .ZN(
        P3_U3167) );
  NOR2_X1 U13475 ( .A1(n10808), .A2(n14286), .ZN(n10809) );
  NOR2_X1 U13476 ( .A1(n10810), .A2(n10809), .ZN(n10902) );
  NAND2_X1 U13477 ( .A1(n10902), .A2(n14526), .ZN(n15294) );
  INV_X1 U13478 ( .A(n15294), .ZN(n15348) );
  INV_X1 U13479 ( .A(n10811), .ZN(n10812) );
  NAND2_X1 U13480 ( .A1(n10812), .A2(n11462), .ZN(n14762) );
  INV_X1 U13481 ( .A(n10813), .ZN(n10814) );
  AND2_X1 U13482 ( .A1(n14292), .A2(n14738), .ZN(n14479) );
  AND2_X1 U13483 ( .A1(n14993), .A2(n14479), .ZN(n15269) );
  AOI21_X1 U13484 ( .B1(n15348), .B2(n14993), .A(n15269), .ZN(n11929) );
  XNOR2_X1 U13485 ( .A(n8892), .B(n14295), .ZN(n15253) );
  INV_X1 U13486 ( .A(n15276), .ZN(n10909) );
  OR2_X1 U13487 ( .A1(n10904), .A2(n10909), .ZN(n11024) );
  XNOR2_X1 U13488 ( .A(n15253), .B(n11024), .ZN(n15278) );
  INV_X1 U13489 ( .A(n15018), .ZN(n10822) );
  INV_X1 U13490 ( .A(n14295), .ZN(n15279) );
  OAI21_X1 U13491 ( .B1(n15279), .B2(n10909), .A(n15263), .ZN(n15281) );
  INV_X1 U13492 ( .A(n15281), .ZN(n10821) );
  NAND2_X1 U13493 ( .A1(n15198), .A2(n14738), .ZN(n10816) );
  NAND2_X1 U13494 ( .A1(n14483), .A2(n10825), .ZN(n10815) );
  AOI21_X1 U13495 ( .B1(n15253), .B2(n14558), .A(n15296), .ZN(n10819) );
  XNOR2_X1 U13496 ( .A(n6853), .B(n15281), .ZN(n10817) );
  OAI21_X1 U13497 ( .B1(n10817), .B2(n15296), .A(n10904), .ZN(n10818) );
  OAI21_X1 U13498 ( .B1(n10819), .B2(n15008), .A(n10818), .ZN(n10820) );
  OAI21_X1 U13499 ( .B1(n14298), .B2(n14855), .A(n10820), .ZN(n15282) );
  AOI21_X1 U13500 ( .B1(n10822), .B2(n10821), .A(n15282), .ZN(n10823) );
  MUX2_X1 U13501 ( .A(n10265), .B(n10823), .S(n14993), .Z(n10828) );
  INV_X1 U13502 ( .A(n10824), .ZN(n15277) );
  NAND2_X1 U13503 ( .A1(n15277), .A2(n10825), .ZN(n10826) );
  INV_X1 U13504 ( .A(n14977), .ZN(n15262) );
  AOI22_X1 U13505 ( .A1(n15260), .A2(n14295), .B1(n15262), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n10827) );
  OAI211_X1 U13506 ( .C1(n11929), .C2(n15278), .A(n10828), .B(n10827), .ZN(
        P1_U3292) );
  INV_X1 U13507 ( .A(n10829), .ZN(n10832) );
  INV_X1 U13508 ( .A(n13652), .ZN(n15467) );
  OAI222_X1 U13509 ( .A1(n14102), .A2(n10830), .B1(n14099), .B2(n10832), .C1(
        n15467), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13510 ( .A1(P1_U3086), .A2(n11900), .B1(n15192), .B2(n10832), 
        .C1(n10831), .C2(n15189), .ZN(P1_U3340) );
  MUX2_X1 U13511 ( .A(n9123), .B(P1_REG2_REG_12__SCAN_IN), .S(n11305), .Z(
        n10839) );
  NAND2_X1 U13512 ( .A1(n10841), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10833) );
  NAND2_X1 U13513 ( .A1(n10834), .A2(n10833), .ZN(n14682) );
  INV_X1 U13514 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10835) );
  MUX2_X1 U13515 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10835), .S(n14679), .Z(
        n14681) );
  NAND2_X1 U13516 ( .A1(n14682), .A2(n14681), .ZN(n14680) );
  NAND2_X1 U13517 ( .A1(n14679), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13518 ( .A1(n14680), .A2(n10836), .ZN(n10838) );
  OR2_X1 U13519 ( .A1(n10838), .A2(n10839), .ZN(n11307) );
  INV_X1 U13520 ( .A(n11307), .ZN(n10837) );
  AOI21_X1 U13521 ( .B1(n10839), .B2(n10838), .A(n10837), .ZN(n10855) );
  INV_X1 U13522 ( .A(n14737), .ZN(n14710) );
  INV_X1 U13523 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10840) );
  XNOR2_X1 U13524 ( .A(n11305), .B(n10840), .ZN(n10848) );
  NAND2_X1 U13525 ( .A1(n10841), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n10842) );
  AND2_X1 U13526 ( .A1(n10843), .A2(n10842), .ZN(n14675) );
  XNOR2_X1 U13527 ( .A(n14679), .B(n10844), .ZN(n14674) );
  NAND2_X1 U13528 ( .A1(n14675), .A2(n14674), .ZN(n14673) );
  NAND2_X1 U13529 ( .A1(n10845), .A2(n10844), .ZN(n10846) );
  NAND2_X1 U13530 ( .A1(n14673), .A2(n10846), .ZN(n10847) );
  NAND2_X1 U13531 ( .A1(n10847), .A2(n10848), .ZN(n11301) );
  OAI21_X1 U13532 ( .B1(n10848), .B2(n10847), .A(n11301), .ZN(n10853) );
  INV_X1 U13533 ( .A(n14733), .ZN(n14732) );
  INV_X1 U13534 ( .A(n14735), .ZN(n10851) );
  AND2_X1 U13535 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n14173) );
  AOI21_X1 U13536 ( .B1(n15247), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n14173), 
        .ZN(n10849) );
  OAI21_X1 U13537 ( .B1(n10851), .B2(n10850), .A(n10849), .ZN(n10852) );
  AOI21_X1 U13538 ( .B1(n10853), .B2(n14732), .A(n10852), .ZN(n10854) );
  OAI21_X1 U13539 ( .B1(n10855), .B2(n14710), .A(n10854), .ZN(P1_U3255) );
  XNOR2_X1 U13540 ( .A(n11272), .B(n6445), .ZN(n10911) );
  XNOR2_X1 U13541 ( .A(n10911), .B(n12577), .ZN(n10874) );
  NAND2_X1 U13542 ( .A1(n10858), .A2(n10856), .ZN(n10862) );
  NAND2_X1 U13543 ( .A1(n10858), .A2(n10857), .ZN(n10861) );
  XNOR2_X1 U13544 ( .A(n6446), .B(n7155), .ZN(n10992) );
  NAND2_X1 U13545 ( .A1(n10992), .A2(n10979), .ZN(n10860) );
  NAND2_X1 U13546 ( .A1(n10859), .A2(n10996), .ZN(n10990) );
  XNOR2_X1 U13547 ( .A(n12435), .B(n6445), .ZN(n10869) );
  INV_X1 U13548 ( .A(n11290), .ZN(n10866) );
  INV_X1 U13549 ( .A(n11288), .ZN(n10864) );
  OAI21_X1 U13550 ( .B1(n10866), .B2(n10995), .A(n10864), .ZN(n10868) );
  INV_X1 U13551 ( .A(n10992), .ZN(n10865) );
  NAND2_X1 U13552 ( .A1(n10865), .A2(n12580), .ZN(n11067) );
  OAI21_X1 U13553 ( .B1(n10866), .B2(n11067), .A(n11288), .ZN(n10867) );
  INV_X1 U13554 ( .A(n10869), .ZN(n10870) );
  NAND2_X1 U13555 ( .A1(n10870), .A2(n12578), .ZN(n10871) );
  INV_X1 U13556 ( .A(n10916), .ZN(n10872) );
  AOI21_X1 U13557 ( .B1(n10874), .B2(n10873), .A(n10872), .ZN(n10883) );
  INV_X1 U13558 ( .A(n10875), .ZN(n11273) );
  OR2_X1 U13559 ( .A1(n12578), .A2(n10876), .ZN(n10877) );
  OAI211_X1 U13560 ( .C1(n12576), .C2(n10878), .A(n10877), .B(n12512), .ZN(
        n11268) );
  NAND2_X1 U13561 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11236) );
  OAI21_X1 U13562 ( .B1(n12313), .B2(n11268), .A(n11236), .ZN(n10879) );
  AOI21_X1 U13563 ( .B1(n12340), .B2(n11273), .A(n10879), .ZN(n10882) );
  INV_X1 U13564 ( .A(n11272), .ZN(n10880) );
  NAND2_X1 U13565 ( .A1(n12347), .A2(n10880), .ZN(n10881) );
  OAI211_X1 U13566 ( .C1(n10883), .C2(n12349), .A(n10882), .B(n10881), .ZN(
        P3_U3171) );
  INV_X1 U13567 ( .A(n10884), .ZN(n10885) );
  OAI21_X1 U13568 ( .B1(n13744), .B2(n10885), .A(n13904), .ZN(n10893) );
  INV_X1 U13569 ( .A(n10886), .ZN(n10888) );
  OAI22_X1 U13570 ( .A1(n13894), .A2(n10888), .B1(n10887), .B2(n13843), .ZN(
        n10889) );
  INV_X1 U13571 ( .A(n10889), .ZN(n10891) );
  OR2_X1 U13572 ( .A1(n11724), .A2(n13539), .ZN(n10890) );
  OAI211_X1 U13573 ( .C1(n10332), .C2(n13913), .A(n10891), .B(n10890), .ZN(
        n10892) );
  AOI21_X1 U13574 ( .B1(n13296), .B2(n10893), .A(n10892), .ZN(n10894) );
  INV_X1 U13575 ( .A(n10894), .ZN(P2_U3265) );
  INV_X1 U13576 ( .A(n14715), .ZN(n10897) );
  INV_X1 U13577 ( .A(n10895), .ZN(n10899) );
  OAI222_X1 U13578 ( .A1(P1_U3086), .A2(n10897), .B1(n15192), .B2(n10899), 
        .C1(n10896), .C2(n15189), .ZN(P1_U3338) );
  INV_X1 U13579 ( .A(n15497), .ZN(n10898) );
  OAI222_X1 U13580 ( .A1(n14102), .A2(n10900), .B1(n14099), .B2(n10899), .C1(
        n10898), .C2(P2_U3088), .ZN(P2_U3310) );
  NOR2_X2 U13581 ( .A1(n6408), .A2(n14738), .ZN(n15268) );
  AOI21_X1 U13582 ( .B1(n15268), .B2(n15277), .A(n15260), .ZN(n10910) );
  AND2_X1 U13583 ( .A1(n8892), .A2(n15010), .ZN(n15275) );
  INV_X1 U13584 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n14569) );
  INV_X1 U13585 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10901) );
  OAI22_X1 U13586 ( .A1(n14993), .A2(n14569), .B1(n10901), .B2(n14977), .ZN(
        n10907) );
  INV_X1 U13587 ( .A(n10902), .ZN(n10903) );
  AND2_X1 U13588 ( .A1(n10904), .A2(n15276), .ZN(n14293) );
  OR2_X1 U13589 ( .A1(n10904), .A2(n15276), .ZN(n14291) );
  INV_X1 U13590 ( .A(n14291), .ZN(n10905) );
  NOR2_X1 U13591 ( .A1(n14293), .A2(n10905), .ZN(n15273) );
  AOI21_X1 U13592 ( .B1(n14925), .B2(n15026), .A(n15273), .ZN(n10906) );
  AOI211_X1 U13593 ( .C1(n15275), .C2(n14993), .A(n10907), .B(n10906), .ZN(
        n10908) );
  OAI21_X1 U13594 ( .B1(n10910), .B2(n10909), .A(n10908), .ZN(P1_U3293) );
  INV_X1 U13595 ( .A(n10911), .ZN(n10912) );
  NAND2_X1 U13596 ( .A1(n10912), .A2(n11294), .ZN(n10914) );
  AND2_X1 U13597 ( .A1(n10916), .A2(n10914), .ZN(n10918) );
  XNOR2_X1 U13598 ( .A(n11390), .B(n6446), .ZN(n11423) );
  XNOR2_X1 U13599 ( .A(n11423), .B(n10913), .ZN(n10917) );
  AND2_X1 U13600 ( .A1(n10917), .A2(n10914), .ZN(n10915) );
  OAI211_X1 U13601 ( .C1(n10918), .C2(n10917), .A(n12308), .B(n11424), .ZN(
        n10923) );
  NAND2_X1 U13602 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n15603)
         );
  OAI21_X1 U13603 ( .B1(n12344), .B2(n10919), .A(n15603), .ZN(n10921) );
  NOR2_X1 U13604 ( .A1(n12321), .A2(n11392), .ZN(n10920) );
  AOI211_X1 U13605 ( .C1(n12341), .C2(n12577), .A(n10921), .B(n10920), .ZN(
        n10922) );
  OAI211_X1 U13606 ( .C1(n12285), .C2(n11390), .A(n10923), .B(n10922), .ZN(
        P3_U3157) );
  INV_X1 U13607 ( .A(n10924), .ZN(n11019) );
  AOI22_X1 U13608 ( .A1(n14718), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n15186), .ZN(n10925) );
  OAI21_X1 U13609 ( .B1(n11019), .B2(n15195), .A(n10925), .ZN(P1_U3337) );
  INV_X1 U13610 ( .A(n12713), .ZN(n12724) );
  INV_X1 U13611 ( .A(n10926), .ZN(n10927) );
  OAI222_X1 U13612 ( .A1(P3_U3151), .A2(n12724), .B1(n13095), .B2(n10928), 
        .C1(n13090), .C2(n10927), .ZN(P3_U3278) );
  OR2_X1 U13613 ( .A1(n13343), .A2(n13274), .ZN(n10930) );
  OR2_X1 U13614 ( .A1(n13330), .A2(n13273), .ZN(n10929) );
  NAND2_X1 U13615 ( .A1(n10930), .A2(n10929), .ZN(n11328) );
  AOI22_X1 U13616 ( .A1(n13275), .A2(n11328), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(P2_U3088), .ZN(n10931) );
  OAI21_X1 U13617 ( .B1(n11322), .B2(n13277), .A(n10931), .ZN(n10932) );
  AOI21_X1 U13618 ( .B1(n14036), .B2(n13280), .A(n10932), .ZN(n10943) );
  INV_X1 U13619 ( .A(n11112), .ZN(n10934) );
  NAND2_X1 U13620 ( .A1(n10934), .A2(n10933), .ZN(n11111) );
  AND2_X1 U13621 ( .A1(n10935), .A2(n11111), .ZN(n10941) );
  XNOR2_X1 U13622 ( .A(n14036), .B(n10936), .ZN(n11110) );
  NAND2_X1 U13623 ( .A1(n13606), .A2(n6409), .ZN(n10937) );
  NAND2_X1 U13624 ( .A1(n11110), .A2(n10937), .ZN(n11114) );
  INV_X1 U13625 ( .A(n11110), .ZN(n10939) );
  INV_X1 U13626 ( .A(n10937), .ZN(n10938) );
  NAND2_X1 U13627 ( .A1(n10939), .A2(n10938), .ZN(n11116) );
  AND2_X1 U13628 ( .A1(n11114), .A2(n11116), .ZN(n10940) );
  NAND2_X1 U13629 ( .A1(n10941), .A2(n10940), .ZN(n11109) );
  OAI211_X1 U13630 ( .C1(n10941), .C2(n10940), .A(n11109), .B(n13270), .ZN(
        n10942) );
  NAND2_X1 U13631 ( .A1(n10943), .A2(n10942), .ZN(P2_U3211) );
  NAND2_X1 U13632 ( .A1(n10944), .A2(n11612), .ZN(n10945) );
  XNOR2_X1 U13633 ( .A(n15428), .B(n10947), .ZN(n15420) );
  NAND2_X1 U13634 ( .A1(n15421), .A2(n15420), .ZN(n15419) );
  NAND2_X1 U13635 ( .A1(n15428), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n10948) );
  MUX2_X1 U13636 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11735), .S(n11751), .Z(
        n10949) );
  NAND2_X1 U13637 ( .A1(n10950), .A2(n10949), .ZN(n11753) );
  OAI21_X1 U13638 ( .B1(n10950), .B2(n10949), .A(n11753), .ZN(n10959) );
  NAND2_X1 U13639 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n12173)
         );
  NAND2_X1 U13640 ( .A1(n15368), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n10951) );
  OAI211_X1 U13641 ( .C1(n15468), .C2(n10952), .A(n12173), .B(n10951), .ZN(
        n10958) );
  OAI21_X1 U13642 ( .B1(n10954), .B2(P2_REG1_REG_9__SCAN_IN), .A(n10953), .ZN(
        n15424) );
  XNOR2_X1 U13643 ( .A(n15428), .B(P2_REG1_REG_10__SCAN_IN), .ZN(n15425) );
  NOR2_X1 U13644 ( .A1(n15424), .A2(n15425), .ZN(n15423) );
  XNOR2_X1 U13645 ( .A(n11751), .B(P2_REG1_REG_11__SCAN_IN), .ZN(n10955) );
  AOI211_X1 U13646 ( .C1(n10956), .C2(n10955), .A(n15492), .B(n11746), .ZN(
        n10957) );
  AOI211_X1 U13647 ( .C1(n15486), .C2(n10959), .A(n10958), .B(n10957), .ZN(
        n10960) );
  INV_X1 U13648 ( .A(n10960), .ZN(P2_U3225) );
  XNOR2_X1 U13649 ( .A(n10961), .B(n12529), .ZN(n15640) );
  INV_X1 U13650 ( .A(n15640), .ZN(n10975) );
  AOI21_X1 U13651 ( .B1(n10964), .B2(n10963), .A(n10962), .ZN(n10978) );
  NAND2_X1 U13652 ( .A1(n10978), .A2(n7413), .ZN(n10977) );
  NAND2_X1 U13653 ( .A1(n10977), .A2(n10965), .ZN(n10966) );
  XOR2_X1 U13654 ( .A(n12529), .B(n10966), .Z(n10968) );
  AOI22_X1 U13655 ( .A1(n12981), .A2(n12579), .B1(n12581), .B2(n12982), .ZN(
        n10967) );
  OAI21_X1 U13656 ( .B1(n10968), .B2(n12834), .A(n10967), .ZN(n10969) );
  AOI21_X1 U13657 ( .B1(n15640), .B2(n12978), .A(n10969), .ZN(n15637) );
  MUX2_X1 U13658 ( .A(n10970), .B(n15637), .S(n15616), .Z(n10974) );
  NOR2_X1 U13659 ( .A1(n10971), .A2(n15626), .ZN(n15639) );
  INV_X1 U13660 ( .A(n11001), .ZN(n10972) );
  AOI22_X1 U13661 ( .A1(n12762), .A2(n15639), .B1(n12912), .B2(n10972), .ZN(
        n10973) );
  OAI211_X1 U13662 ( .C1(n10975), .C2(n11276), .A(n10974), .B(n10973), .ZN(
        P3_U3227) );
  XNOR2_X1 U13663 ( .A(n10976), .B(n7413), .ZN(n15632) );
  OAI21_X1 U13664 ( .B1(n10978), .B2(n7413), .A(n10977), .ZN(n10984) );
  OAI22_X1 U13665 ( .A1(n10980), .A2(n12836), .B1(n10979), .B2(n12838), .ZN(
        n10983) );
  NOR2_X1 U13666 ( .A1(n15632), .A2(n10981), .ZN(n10982) );
  AOI211_X1 U13667 ( .C1(n12986), .C2(n10984), .A(n10983), .B(n10982), .ZN(
        n15633) );
  MUX2_X1 U13668 ( .A(n7619), .B(n15633), .S(n15616), .Z(n10989) );
  NOR2_X1 U13669 ( .A1(n10985), .A2(n15626), .ZN(n15635) );
  INV_X1 U13670 ( .A(n10986), .ZN(n10987) );
  AOI22_X1 U13671 ( .A1(n12762), .A2(n15635), .B1(n12912), .B2(n10987), .ZN(
        n10988) );
  OAI211_X1 U13672 ( .C1(n15632), .C2(n11276), .A(n10989), .B(n10988), .ZN(
        P3_U3228) );
  AND2_X1 U13673 ( .A1(n10991), .A2(n10990), .ZN(n10994) );
  XNOR2_X1 U13674 ( .A(n10992), .B(n12580), .ZN(n10993) );
  NAND2_X1 U13675 ( .A1(n10994), .A2(n10993), .ZN(n11068) );
  OAI211_X1 U13676 ( .C1(n10994), .C2(n10993), .A(n11068), .B(n12308), .ZN(
        n11000) );
  NAND2_X1 U13677 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15558) );
  INV_X1 U13678 ( .A(n15558), .ZN(n10998) );
  OAI22_X1 U13679 ( .A1(n12292), .A2(n10996), .B1(n10995), .B2(n12344), .ZN(
        n10997) );
  AOI211_X1 U13680 ( .C1(n12347), .C2(n7155), .A(n10998), .B(n10997), .ZN(
        n10999) );
  OAI211_X1 U13681 ( .C1(n11001), .C2(n12321), .A(n11000), .B(n10999), .ZN(
        P3_U3179) );
  OR2_X1 U13682 ( .A1(n11003), .A2(n11002), .ZN(n11004) );
  AND2_X1 U13683 ( .A1(n11005), .A2(n11004), .ZN(n11012) );
  OAI21_X1 U13684 ( .B1(n11006), .B2(n13543), .A(n11186), .ZN(n11007) );
  NAND2_X1 U13685 ( .A1(n11007), .A2(n13897), .ZN(n11009) );
  AOI22_X1 U13686 ( .A1(n13607), .A2(n13880), .B1(n13878), .B2(n13609), .ZN(
        n11008) );
  MUX2_X1 U13687 ( .A(n15519), .B(P2_REG2_REG_4__SCAN_IN), .S(n13894), .Z(
        n11017) );
  AOI21_X1 U13688 ( .B1(n11010), .B2(n13320), .A(n6409), .ZN(n11011) );
  NAND2_X1 U13689 ( .A1(n6885), .A2(n11011), .ZN(n15517) );
  INV_X1 U13690 ( .A(n11012), .ZN(n15521) );
  INV_X1 U13691 ( .A(n11724), .ZN(n13921) );
  NAND2_X1 U13692 ( .A1(n15521), .A2(n13921), .ZN(n11015) );
  OAI22_X1 U13693 ( .A1(n13904), .A2(n7013), .B1(n13184), .B2(n13843), .ZN(
        n11013) );
  INV_X1 U13694 ( .A(n11013), .ZN(n11014) );
  OAI211_X1 U13695 ( .C1(n13744), .C2(n15517), .A(n11015), .B(n11014), .ZN(
        n11016) );
  OR2_X1 U13696 ( .A1(n11017), .A2(n11016), .ZN(P2_U3261) );
  INV_X1 U13697 ( .A(n13663), .ZN(n13653) );
  INV_X1 U13698 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11018) );
  OAI222_X1 U13699 ( .A1(P2_U3088), .A2(n13653), .B1(n14099), .B2(n11019), 
        .C1(n11018), .C2(n14102), .ZN(P2_U3309) );
  INV_X1 U13700 ( .A(n14502), .ZN(n11022) );
  NAND2_X1 U13701 ( .A1(n8892), .A2(n15279), .ZN(n11020) );
  NAND2_X1 U13702 ( .A1(n11020), .A2(n14293), .ZN(n11021) );
  NAND2_X1 U13703 ( .A1(n11022), .A2(n15255), .ZN(n11023) );
  NAND2_X1 U13704 ( .A1(n11023), .A2(n14289), .ZN(n11049) );
  XNOR2_X1 U13705 ( .A(n11052), .B(n11049), .ZN(n15297) );
  INV_X1 U13706 ( .A(n11929), .ZN(n11536) );
  NAND2_X1 U13707 ( .A1(n11024), .A2(n15279), .ZN(n11025) );
  INV_X1 U13708 ( .A(n11024), .ZN(n15252) );
  AOI22_X1 U13709 ( .A1(n8892), .A2(n11025), .B1(n15252), .B2(n14295), .ZN(
        n11026) );
  NAND2_X1 U13710 ( .A1(n14502), .A2(n11026), .ZN(n11028) );
  NAND2_X1 U13711 ( .A1(n14298), .A2(n15286), .ZN(n11027) );
  NAND2_X1 U13712 ( .A1(n11028), .A2(n11027), .ZN(n11053) );
  XNOR2_X1 U13713 ( .A(n11053), .B(n14503), .ZN(n15295) );
  INV_X1 U13714 ( .A(n15295), .ZN(n15300) );
  INV_X1 U13715 ( .A(n11029), .ZN(n15265) );
  AOI21_X1 U13716 ( .B1(n15265), .B2(n14148), .A(n15280), .ZN(n11031) );
  INV_X1 U13717 ( .A(n11051), .ZN(n11030) );
  NAND2_X1 U13718 ( .A1(n11031), .A2(n11030), .ZN(n15292) );
  NOR2_X1 U13719 ( .A1(n14982), .A2(n15292), .ZN(n11038) );
  INV_X1 U13720 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n14145) );
  AOI22_X1 U13721 ( .A1(n6408), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15262), .B2(
        n14145), .ZN(n11036) );
  NAND2_X1 U13722 ( .A1(n14555), .A2(n15010), .ZN(n11033) );
  NAND2_X1 U13723 ( .A1(n14557), .A2(n15008), .ZN(n11032) );
  AND2_X1 U13724 ( .A1(n11033), .A2(n11032), .ZN(n15291) );
  INV_X1 U13725 ( .A(n15291), .ZN(n11034) );
  NAND2_X1 U13726 ( .A1(n14993), .A2(n11034), .ZN(n11035) );
  OAI211_X1 U13727 ( .C1(n14994), .C2(n15293), .A(n11036), .B(n11035), .ZN(
        n11037) );
  AOI211_X1 U13728 ( .C1(n11536), .C2(n15300), .A(n11038), .B(n11037), .ZN(
        n11039) );
  OAI21_X1 U13729 ( .B1(n15026), .B2(n15297), .A(n11039), .ZN(P1_U3290) );
  INV_X1 U13730 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n11047) );
  AOI22_X1 U13731 ( .A1(n13275), .A2(n11040), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11041) );
  OAI21_X1 U13732 ( .B1(n6888), .B2(n13227), .A(n11041), .ZN(n11046) );
  INV_X1 U13733 ( .A(n13188), .ZN(n11042) );
  AOI211_X1 U13734 ( .C1(n11044), .C2(n11043), .A(n11042), .B(n13250), .ZN(
        n11045) );
  AOI211_X1 U13735 ( .C1(n13261), .C2(n11047), .A(n11046), .B(n11045), .ZN(
        n11048) );
  INV_X1 U13736 ( .A(n11048), .ZN(P2_U3190) );
  INV_X1 U13737 ( .A(n15026), .ZN(n14914) );
  NAND2_X1 U13738 ( .A1(n11049), .A2(n14503), .ZN(n11050) );
  NAND2_X1 U13739 ( .A1(n11050), .A2(n14303), .ZN(n11132) );
  XNOR2_X1 U13740 ( .A(n11132), .B(n14501), .ZN(n15310) );
  INV_X1 U13741 ( .A(n14309), .ZN(n11058) );
  OAI211_X1 U13742 ( .C1(n11051), .C2(n11058), .A(n15264), .B(n11139), .ZN(
        n15306) );
  NAND2_X1 U13743 ( .A1(n11053), .A2(n11052), .ZN(n11056) );
  NAND2_X1 U13744 ( .A1(n11054), .A2(n15293), .ZN(n11055) );
  NAND2_X1 U13745 ( .A1(n11056), .A2(n11055), .ZN(n11057) );
  NAND2_X1 U13746 ( .A1(n11057), .A2(n14501), .ZN(n15302) );
  NAND3_X1 U13747 ( .A1(n15303), .A2(n15024), .A3(n15302), .ZN(n11064) );
  OAI22_X1 U13748 ( .A1(n14994), .A2(n11058), .B1(n14977), .B2(n11151), .ZN(
        n11062) );
  NAND2_X1 U13749 ( .A1(n14554), .A2(n15010), .ZN(n11060) );
  NAND2_X1 U13750 ( .A1(n14556), .A2(n15008), .ZN(n11059) );
  NAND2_X1 U13751 ( .A1(n11060), .A2(n11059), .ZN(n15305) );
  MUX2_X1 U13752 ( .A(n15305), .B(P1_REG2_REG_4__SCAN_IN), .S(n6408), .Z(
        n11061) );
  NOR2_X1 U13753 ( .A1(n11062), .A2(n11061), .ZN(n11063) );
  OAI211_X1 U13754 ( .C1(n15306), .C2(n14982), .A(n11064), .B(n11063), .ZN(
        n11065) );
  AOI21_X1 U13755 ( .B1(n14914), .B2(n15310), .A(n11065), .ZN(n11066) );
  INV_X1 U13756 ( .A(n11066), .ZN(P1_U3289) );
  NAND2_X1 U13757 ( .A1(n11068), .A2(n11067), .ZN(n11289) );
  XNOR2_X1 U13758 ( .A(n11288), .B(n11289), .ZN(n11074) );
  INV_X1 U13759 ( .A(n11069), .ZN(n11097) );
  INV_X1 U13760 ( .A(n12344), .ZN(n12289) );
  AOI22_X1 U13761 ( .A1(n12289), .A2(n12578), .B1(n12341), .B2(n12580), .ZN(
        n11071) );
  OAI211_X1 U13762 ( .C1(n12285), .C2(n11096), .A(n11071), .B(n11070), .ZN(
        n11072) );
  AOI21_X1 U13763 ( .B1(n11097), .B2(n12340), .A(n11072), .ZN(n11073) );
  OAI21_X1 U13764 ( .B1(n11074), .B2(n12349), .A(n11073), .ZN(P3_U3153) );
  AOI21_X1 U13765 ( .B1(n14142), .B2(n11076), .A(n11077), .ZN(n11145) );
  INV_X1 U13766 ( .A(n11148), .ZN(n11078) );
  NAND3_X1 U13767 ( .A1(n14142), .A2(n11077), .A3(n11076), .ZN(n11146) );
  OAI21_X1 U13768 ( .B1(n11145), .B2(n11078), .A(n11146), .ZN(n11082) );
  NAND2_X1 U13769 ( .A1(n11080), .A2(n11079), .ZN(n11081) );
  XNOR2_X1 U13770 ( .A(n11082), .B(n11081), .ZN(n11088) );
  AND2_X1 U13771 ( .A1(n14313), .A2(n15336), .ZN(n15314) );
  NAND2_X1 U13772 ( .A1(n14553), .A2(n15010), .ZN(n11084) );
  NAND2_X1 U13773 ( .A1(n14555), .A2(n15008), .ZN(n11083) );
  NAND2_X1 U13774 ( .A1(n11084), .A2(n11083), .ZN(n11135) );
  AOI22_X1 U13775 ( .A1(n11135), .A2(n14282), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11085) );
  OAI21_X1 U13776 ( .B1(n14279), .B2(n11140), .A(n11085), .ZN(n11086) );
  AOI21_X1 U13777 ( .B1(n14218), .B2(n15314), .A(n11086), .ZN(n11087) );
  OAI21_X1 U13778 ( .B1(n11088), .B2(n14271), .A(n11087), .ZN(P1_U3227) );
  INV_X1 U13779 ( .A(n12425), .ZN(n11089) );
  NOR2_X1 U13780 ( .A1(n11090), .A2(n11089), .ZN(n11254) );
  XNOR2_X1 U13781 ( .A(n11254), .B(n7209), .ZN(n15644) );
  INV_X1 U13782 ( .A(n15644), .ZN(n11100) );
  OAI211_X1 U13783 ( .C1(n11092), .C2(n7209), .A(n11091), .B(n12986), .ZN(
        n11094) );
  AOI22_X1 U13784 ( .A1(n12981), .A2(n12578), .B1(n12580), .B2(n12982), .ZN(
        n11093) );
  NAND2_X1 U13785 ( .A1(n11094), .A2(n11093), .ZN(n11095) );
  AOI21_X1 U13786 ( .B1(n15644), .B2(n12978), .A(n11095), .ZN(n15641) );
  MUX2_X1 U13787 ( .A(n6909), .B(n15641), .S(n15616), .Z(n11099) );
  NOR2_X1 U13788 ( .A1(n11096), .A2(n15626), .ZN(n15643) );
  AOI22_X1 U13789 ( .A1(n12762), .A2(n15643), .B1(n12912), .B2(n11097), .ZN(
        n11098) );
  OAI211_X1 U13790 ( .C1(n11100), .C2(n11276), .A(n11099), .B(n11098), .ZN(
        P3_U3226) );
  INV_X1 U13791 ( .A(n11101), .ZN(n11102) );
  OAI222_X1 U13792 ( .A1(P3_U3151), .A2(n12746), .B1(n13095), .B2(n11103), 
        .C1(n13090), .C2(n11102), .ZN(P3_U3277) );
  INV_X1 U13793 ( .A(n15525), .ZN(n11130) );
  XNOR2_X1 U13794 ( .A(n15525), .B(n13139), .ZN(n12185) );
  NOR2_X1 U13795 ( .A1(n13343), .A2(n6405), .ZN(n11104) );
  NAND2_X1 U13796 ( .A1(n12185), .A2(n11104), .ZN(n11657) );
  INV_X1 U13797 ( .A(n12185), .ZN(n11106) );
  INV_X1 U13798 ( .A(n11104), .ZN(n11105) );
  NAND2_X1 U13799 ( .A1(n11106), .A2(n11105), .ZN(n11107) );
  AND2_X1 U13800 ( .A1(n11657), .A2(n11107), .ZN(n11119) );
  INV_X1 U13801 ( .A(n11119), .ZN(n11108) );
  AOI21_X1 U13802 ( .B1(n11109), .B2(n11108), .A(n13250), .ZN(n11122) );
  NOR3_X1 U13803 ( .A1(n13256), .A2(n11182), .A3(n11110), .ZN(n11121) );
  NAND2_X1 U13804 ( .A1(n11114), .A2(n11111), .ZN(n11117) );
  NAND3_X1 U13805 ( .A1(n11114), .A2(n11113), .A3(n11112), .ZN(n11115) );
  OAI211_X1 U13806 ( .C1(n11118), .C2(n11117), .A(n11116), .B(n11115), .ZN(
        n11120) );
  OAI21_X1 U13807 ( .B1(n11122), .B2(n11121), .A(n12187), .ZN(n11129) );
  INV_X1 U13808 ( .A(n11174), .ZN(n11127) );
  OR2_X1 U13809 ( .A1(n13345), .A2(n13274), .ZN(n11124) );
  NAND2_X1 U13810 ( .A1(n13606), .A2(n13878), .ZN(n11123) );
  AND2_X1 U13811 ( .A1(n11124), .A2(n11123), .ZN(n11168) );
  OAI22_X1 U13812 ( .A1(n13263), .A2(n11168), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11125), .ZN(n11126) );
  AOI21_X1 U13813 ( .B1(n11127), .B2(n13261), .A(n11126), .ZN(n11128) );
  OAI211_X1 U13814 ( .C1(n11130), .C2(n13227), .A(n11129), .B(n11128), .ZN(
        P2_U3185) );
  NAND2_X1 U13815 ( .A1(n14555), .A2(n14309), .ZN(n11401) );
  AND2_X1 U13816 ( .A1(n15303), .A2(n11401), .ZN(n11131) );
  XNOR2_X1 U13817 ( .A(n14554), .B(n11345), .ZN(n14506) );
  NAND2_X1 U13818 ( .A1(n11131), .A2(n14506), .ZN(n11342) );
  OAI21_X1 U13819 ( .B1(n11131), .B2(n14506), .A(n11342), .ZN(n15318) );
  INV_X1 U13820 ( .A(n15318), .ZN(n11144) );
  NAND2_X1 U13821 ( .A1(n11132), .A2(n14501), .ZN(n11134) );
  INV_X1 U13822 ( .A(n14555), .ZN(n14146) );
  NAND2_X1 U13823 ( .A1(n14146), .A2(n14309), .ZN(n11133) );
  XNOR2_X1 U13824 ( .A(n11344), .B(n14506), .ZN(n11137) );
  INV_X1 U13825 ( .A(n11135), .ZN(n11136) );
  OAI21_X1 U13826 ( .B1(n11137), .B2(n15296), .A(n11136), .ZN(n15317) );
  INV_X1 U13827 ( .A(n15317), .ZN(n11138) );
  MUX2_X1 U13828 ( .A(n10275), .B(n11138), .S(n14993), .Z(n11143) );
  AOI211_X1 U13829 ( .C1(n14313), .C2(n11139), .A(n15280), .B(n11350), .ZN(
        n15313) );
  OAI22_X1 U13830 ( .A1(n14994), .A2(n11345), .B1(n14977), .B2(n11140), .ZN(
        n11141) );
  AOI21_X1 U13831 ( .B1(n15313), .B2(n15268), .A(n11141), .ZN(n11142) );
  OAI211_X1 U13832 ( .C1(n11929), .C2(n11144), .A(n11143), .B(n11142), .ZN(
        P1_U3288) );
  INV_X1 U13833 ( .A(n11145), .ZN(n11147) );
  NAND2_X1 U13834 ( .A1(n11147), .A2(n11146), .ZN(n11149) );
  XNOR2_X1 U13835 ( .A(n11149), .B(n11148), .ZN(n11154) );
  AND2_X1 U13836 ( .A1(n14309), .A2(n15336), .ZN(n15304) );
  NAND2_X1 U13837 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n14603) );
  NAND2_X1 U13838 ( .A1(n15305), .A2(n14282), .ZN(n11150) );
  OAI211_X1 U13839 ( .C1(n14279), .C2(n11151), .A(n14603), .B(n11150), .ZN(
        n11152) );
  AOI21_X1 U13840 ( .B1(n14218), .B2(n15304), .A(n11152), .ZN(n11153) );
  OAI21_X1 U13841 ( .B1(n11154), .B2(n14271), .A(n11153), .ZN(P1_U3230) );
  INV_X1 U13842 ( .A(n11155), .ZN(n11157) );
  NOR2_X1 U13843 ( .A1(n11157), .A2(n11156), .ZN(n11158) );
  XNOR2_X1 U13844 ( .A(n11159), .B(n11158), .ZN(n11163) );
  AND2_X1 U13845 ( .A1(n14319), .A2(n15336), .ZN(n15323) );
  OAI22_X1 U13846 ( .A1(n14267), .A2(n11571), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15783), .ZN(n11161) );
  INV_X1 U13847 ( .A(n14264), .ZN(n14255) );
  OAI22_X1 U13848 ( .A1(n14255), .A2(n11402), .B1(n14279), .B2(n11352), .ZN(
        n11160) );
  AOI211_X1 U13849 ( .C1(n14218), .C2(n15323), .A(n11161), .B(n11160), .ZN(
        n11162) );
  OAI21_X1 U13850 ( .B1(n11163), .B2(n14271), .A(n11162), .ZN(P1_U3239) );
  OAI222_X1 U13851 ( .A1(P3_U3151), .A2(n12743), .B1(n13090), .B2(n11165), 
        .C1(n11164), .C2(n13095), .ZN(P3_U3276) );
  INV_X1 U13852 ( .A(n11171), .ZN(n13547) );
  XNOR2_X1 U13853 ( .A(n11166), .B(n13547), .ZN(n11167) );
  NAND2_X1 U13854 ( .A1(n11167), .A2(n13897), .ZN(n11169) );
  NAND2_X1 U13855 ( .A1(n11169), .A2(n11168), .ZN(n15530) );
  INV_X1 U13856 ( .A(n15530), .ZN(n11180) );
  XNOR2_X1 U13857 ( .A(n11170), .B(n11171), .ZN(n15523) );
  INV_X1 U13858 ( .A(n13908), .ZN(n13826) );
  NAND2_X1 U13859 ( .A1(n15525), .A2(n11319), .ZN(n11172) );
  NAND2_X1 U13860 ( .A1(n11172), .A2(n6406), .ZN(n11173) );
  OR2_X1 U13861 ( .A1(n11173), .A2(n11364), .ZN(n15527) );
  OAI22_X1 U13862 ( .A1(n13913), .A2(n11175), .B1(n11174), .B2(n13843), .ZN(
        n11176) );
  AOI21_X1 U13863 ( .B1(n13917), .B2(n15525), .A(n11176), .ZN(n11177) );
  OAI21_X1 U13864 ( .B1(n13744), .B2(n15527), .A(n11177), .ZN(n11178) );
  AOI21_X1 U13865 ( .B1(n15523), .B2(n13826), .A(n11178), .ZN(n11179) );
  OAI21_X1 U13866 ( .B1(n11180), .B2(n13797), .A(n11179), .ZN(P2_U3258) );
  INV_X1 U13867 ( .A(n13545), .ZN(n11184) );
  XNOR2_X1 U13868 ( .A(n11181), .B(n11184), .ZN(n11278) );
  OAI22_X1 U13869 ( .A1(n11183), .A2(n13273), .B1(n11182), .B2(n13274), .ZN(
        n11190) );
  NAND3_X1 U13870 ( .A1(n11186), .A2(n11185), .A3(n11184), .ZN(n11187) );
  AOI21_X1 U13871 ( .B1(n11188), .B2(n11187), .A(n13836), .ZN(n11189) );
  AOI211_X1 U13872 ( .C1(n12152), .C2(n11278), .A(n11190), .B(n11189), .ZN(
        n11280) );
  OAI211_X1 U13873 ( .C1(n11192), .C2(n11191), .A(n6405), .B(n11321), .ZN(
        n11279) );
  NAND2_X1 U13874 ( .A1(n13894), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n11193) );
  OAI21_X1 U13875 ( .B1(n13843), .B2(n11194), .A(n11193), .ZN(n11195) );
  AOI21_X1 U13876 ( .B1(n13917), .B2(n13328), .A(n11195), .ZN(n11196) );
  OAI21_X1 U13877 ( .B1(n13744), .B2(n11279), .A(n11196), .ZN(n11197) );
  AOI21_X1 U13878 ( .B1(n13921), .B2(n11278), .A(n11197), .ZN(n11198) );
  OAI21_X1 U13879 ( .B1(n11280), .B2(n13797), .A(n11198), .ZN(P2_U3260) );
  OAI21_X1 U13880 ( .B1(n13540), .B2(n11200), .A(n11199), .ZN(n11206) );
  OAI22_X1 U13881 ( .A1(n7395), .A2(n13274), .B1(n8651), .B2(n13273), .ZN(
        n11205) );
  NAND2_X1 U13882 ( .A1(n12144), .A2(n7962), .ZN(n11202) );
  INV_X1 U13883 ( .A(n13540), .ZN(n11201) );
  XNOR2_X1 U13884 ( .A(n11202), .B(n11201), .ZN(n15516) );
  INV_X1 U13885 ( .A(n15516), .ZN(n11203) );
  AOI211_X1 U13886 ( .C1(n13897), .C2(n11206), .A(n11205), .B(n11204), .ZN(
        n15513) );
  OAI211_X1 U13887 ( .C1(n12147), .C2(n15512), .A(n11207), .B(n6406), .ZN(
        n15511) );
  OAI22_X1 U13888 ( .A1(n13913), .A2(n11209), .B1(n11208), .B2(n13843), .ZN(
        n11210) );
  AOI21_X1 U13889 ( .B1(n13917), .B2(n6751), .A(n11210), .ZN(n11211) );
  OAI21_X1 U13890 ( .B1(n13744), .B2(n15511), .A(n11211), .ZN(n11212) );
  AOI21_X1 U13891 ( .B1(n13921), .B2(n15516), .A(n11212), .ZN(n11213) );
  OAI21_X1 U13892 ( .B1(n13894), .B2(n15513), .A(n11213), .ZN(P2_U3263) );
  INV_X1 U13893 ( .A(n11214), .ZN(n11216) );
  OAI222_X1 U13894 ( .A1(n15189), .A2(n11215), .B1(n15192), .B2(n11216), .C1(
        P1_U3086), .C2(n14526), .ZN(P1_U3336) );
  OAI222_X1 U13895 ( .A1(n14102), .A2(n11217), .B1(n14099), .B2(n11216), .C1(
        n13568), .C2(P2_U3088), .ZN(P2_U3308) );
  NAND2_X1 U13896 ( .A1(n11220), .A2(n11219), .ZN(n11221) );
  NAND2_X1 U13897 ( .A1(n11222), .A2(n11221), .ZN(n15562) );
  MUX2_X1 U13898 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n11223), .S(n11239), .Z(
        n15563) );
  NAND2_X1 U13899 ( .A1(n15562), .A2(n15563), .ZN(n15561) );
  NAND2_X1 U13900 ( .A1(n11239), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n11224) );
  XNOR2_X1 U13901 ( .A(n11686), .B(n11235), .ZN(n11685) );
  XOR2_X1 U13902 ( .A(n11685), .B(P3_REG1_REG_9__SCAN_IN), .Z(n11248) );
  NAND2_X1 U13903 ( .A1(n11226), .A2(n11225), .ZN(n11231) );
  INV_X1 U13904 ( .A(n11227), .ZN(n11229) );
  NAND2_X1 U13905 ( .A1(n11229), .A2(n11228), .ZN(n11230) );
  NAND2_X1 U13906 ( .A1(n11231), .A2(n11230), .ZN(n15564) );
  MUX2_X1 U13907 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n7168), .Z(n11232) );
  INV_X1 U13908 ( .A(n11239), .ZN(n15574) );
  XNOR2_X1 U13909 ( .A(n11232), .B(n15574), .ZN(n15565) );
  INV_X1 U13910 ( .A(n11232), .ZN(n11233) );
  NAND2_X1 U13911 ( .A1(n11233), .A2(n15574), .ZN(n11234) );
  MUX2_X1 U13912 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n7168), .Z(n11695) );
  XNOR2_X1 U13913 ( .A(n11695), .B(n11235), .ZN(n11696) );
  XNOR2_X1 U13914 ( .A(n11697), .B(n11696), .ZN(n11246) );
  INV_X1 U13915 ( .A(n11236), .ZN(n11237) );
  AOI21_X1 U13916 ( .B1(n15539), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11237), .ZN(
        n11238) );
  OAI21_X1 U13917 ( .B1(n15549), .B2(n11694), .A(n11238), .ZN(n11245) );
  INV_X1 U13918 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n11260) );
  XNOR2_X1 U13919 ( .A(n11239), .B(n11260), .ZN(n15566) );
  NAND2_X1 U13920 ( .A1(n11239), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U13921 ( .A1(n15572), .A2(n11240), .ZN(n11241) );
  INV_X1 U13922 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11271) );
  NAND2_X1 U13923 ( .A1(n11242), .A2(n11271), .ZN(n11243) );
  AOI21_X1 U13924 ( .B1(n15585), .B2(n11243), .A(n15570), .ZN(n11244) );
  AOI211_X1 U13925 ( .C1(n15595), .C2(n11246), .A(n11245), .B(n11244), .ZN(
        n11247) );
  OAI21_X1 U13926 ( .B1(n11248), .B2(n12730), .A(n11247), .ZN(P3_U3191) );
  XNOR2_X1 U13927 ( .A(n11249), .B(n7081), .ZN(n11250) );
  AOI222_X1 U13928 ( .A1(n12577), .A2(n12982), .B1(n12986), .B2(n11250), .C1(
        n12575), .C2(n12981), .ZN(n11395) );
  XNOR2_X1 U13929 ( .A(n11251), .B(n7081), .ZN(n11391) );
  INV_X1 U13930 ( .A(n13065), .ZN(n11605) );
  NAND2_X1 U13931 ( .A1(n11391), .A2(n11605), .ZN(n11253) );
  INV_X1 U13932 ( .A(n11390), .ZN(n11394) );
  AOI22_X1 U13933 ( .A1(n13061), .A2(n11394), .B1(n15653), .B2(
        P3_REG0_REG_10__SCAN_IN), .ZN(n11252) );
  OAI211_X1 U13934 ( .C1(n11395), .C2(n15653), .A(n11253), .B(n11252), .ZN(
        P3_U3420) );
  OAI21_X1 U13935 ( .B1(n11254), .B2(n7209), .A(n12432), .ZN(n11255) );
  XNOR2_X1 U13936 ( .A(n11255), .B(n12530), .ZN(n15648) );
  INV_X1 U13937 ( .A(n15648), .ZN(n11264) );
  XOR2_X1 U13938 ( .A(n11256), .B(n12530), .Z(n11258) );
  AOI22_X1 U13939 ( .A1(n12981), .A2(n12577), .B1(n12579), .B2(n12982), .ZN(
        n11257) );
  OAI21_X1 U13940 ( .B1(n11258), .B2(n12834), .A(n11257), .ZN(n11259) );
  AOI21_X1 U13941 ( .B1(n15648), .B2(n12978), .A(n11259), .ZN(n15645) );
  MUX2_X1 U13942 ( .A(n11260), .B(n15645), .S(n15616), .Z(n11263) );
  AND2_X1 U13943 ( .A1(n12435), .A2(n12933), .ZN(n15647) );
  INV_X1 U13944 ( .A(n11261), .ZN(n11297) );
  AOI22_X1 U13945 ( .A1(n12762), .A2(n15647), .B1(n12912), .B2(n11297), .ZN(
        n11262) );
  OAI211_X1 U13946 ( .C1(n11264), .C2(n11276), .A(n11263), .B(n11262), .ZN(
        P3_U3225) );
  XNOR2_X1 U13947 ( .A(n11265), .B(n11267), .ZN(n15652) );
  INV_X1 U13948 ( .A(n15652), .ZN(n11277) );
  XNOR2_X1 U13949 ( .A(n11266), .B(n11267), .ZN(n11269) );
  OAI21_X1 U13950 ( .B1(n11269), .B2(n12834), .A(n11268), .ZN(n11270) );
  AOI21_X1 U13951 ( .B1(n15652), .B2(n12978), .A(n11270), .ZN(n15649) );
  MUX2_X1 U13952 ( .A(n11271), .B(n15649), .S(n15616), .Z(n11275) );
  NOR2_X1 U13953 ( .A1(n11272), .A2(n15626), .ZN(n15651) );
  AOI22_X1 U13954 ( .A1(n15651), .A2(n12762), .B1(n12912), .B2(n11273), .ZN(
        n11274) );
  OAI211_X1 U13955 ( .C1(n11277), .C2(n11276), .A(n11275), .B(n11274), .ZN(
        P3_U3224) );
  INV_X1 U13956 ( .A(n11278), .ZN(n11281) );
  OAI211_X1 U13957 ( .C1(n11281), .C2(n13285), .A(n11280), .B(n11279), .ZN(
        n11284) );
  NAND2_X1 U13958 ( .A1(n11284), .A2(n15538), .ZN(n11283) );
  NAND2_X1 U13959 ( .A1(n14023), .A2(n13328), .ZN(n11282) );
  OAI211_X1 U13960 ( .C1(n15538), .C2(n10301), .A(n11283), .B(n11282), .ZN(
        P2_U3504) );
  INV_X1 U13961 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11287) );
  NAND2_X1 U13962 ( .A1(n11284), .A2(n15533), .ZN(n11286) );
  NAND2_X1 U13963 ( .A1(n14086), .A2(n13328), .ZN(n11285) );
  OAI211_X1 U13964 ( .C1(n15533), .C2(n11287), .A(n11286), .B(n11285), .ZN(
        P2_U3445) );
  MUX2_X1 U13965 ( .A(n12579), .B(n11289), .S(n11288), .Z(n11291) );
  XNOR2_X1 U13966 ( .A(n11291), .B(n11290), .ZN(n11299) );
  INV_X1 U13967 ( .A(n12435), .ZN(n11292) );
  NOR2_X1 U13968 ( .A1(n12285), .A2(n11292), .ZN(n11296) );
  NAND2_X1 U13969 ( .A1(n12341), .A2(n12579), .ZN(n11293) );
  NAND2_X1 U13970 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15580) );
  OAI211_X1 U13971 ( .C1(n12344), .C2(n11294), .A(n11293), .B(n15580), .ZN(
        n11295) );
  AOI211_X1 U13972 ( .C1(n11297), .C2(n12340), .A(n11296), .B(n11295), .ZN(
        n11298) );
  OAI21_X1 U13973 ( .B1(n11299), .B2(n12349), .A(n11298), .ZN(P3_U3161) );
  XNOR2_X1 U13974 ( .A(n11377), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n11304) );
  OR2_X1 U13975 ( .A1(n11305), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n11300) );
  NAND2_X1 U13976 ( .A1(n11301), .A2(n11300), .ZN(n11303) );
  INV_X1 U13977 ( .A(n11372), .ZN(n11302) );
  AOI211_X1 U13978 ( .C1(n11304), .C2(n11303), .A(n14733), .B(n11302), .ZN(
        n11317) );
  INV_X1 U13979 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11857) );
  MUX2_X1 U13980 ( .A(n11857), .B(P1_REG2_REG_13__SCAN_IN), .S(n11377), .Z(
        n11310) );
  OR2_X1 U13981 ( .A1(n11305), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U13982 ( .A1(n11307), .A2(n11306), .ZN(n11309) );
  OR2_X1 U13983 ( .A1(n11309), .A2(n11310), .ZN(n11379) );
  INV_X1 U13984 ( .A(n11379), .ZN(n11308) );
  AOI211_X1 U13985 ( .C1(n11310), .C2(n11309), .A(n14710), .B(n11308), .ZN(
        n11316) );
  NAND2_X1 U13986 ( .A1(n14735), .A2(n11377), .ZN(n11313) );
  NOR2_X1 U13987 ( .A1(n11311), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14236) );
  INV_X1 U13988 ( .A(n14236), .ZN(n11312) );
  OAI211_X1 U13989 ( .C1(n14742), .C2(n11314), .A(n11313), .B(n11312), .ZN(
        n11315) );
  OR3_X1 U13990 ( .A1(n11317), .A2(n11316), .A3(n11315), .ZN(P1_U3256) );
  XNOR2_X1 U13991 ( .A(n11318), .B(n13546), .ZN(n14039) );
  INV_X1 U13992 ( .A(n11319), .ZN(n11320) );
  AOI211_X1 U13993 ( .C1(n14036), .C2(n11321), .A(n6409), .B(n11320), .ZN(
        n14035) );
  INV_X1 U13994 ( .A(n14036), .ZN(n11325) );
  INV_X1 U13995 ( .A(n11322), .ZN(n11323) );
  AOI22_X1 U13996 ( .A1(n13894), .A2(P2_REG2_REG_6__SCAN_IN), .B1(n11323), 
        .B2(n13915), .ZN(n11324) );
  OAI21_X1 U13997 ( .B1(n11325), .B2(n13904), .A(n11324), .ZN(n11331) );
  OAI21_X1 U13998 ( .B1(n11327), .B2(n13546), .A(n11326), .ZN(n11329) );
  AOI21_X1 U13999 ( .B1(n11329), .B2(n13897), .A(n11328), .ZN(n14038) );
  NOR2_X1 U14000 ( .A1(n14038), .A2(n13894), .ZN(n11330) );
  AOI211_X1 U14001 ( .C1(n14035), .C2(n13919), .A(n11331), .B(n11330), .ZN(
        n11332) );
  OAI21_X1 U14002 ( .B1(n13908), .B2(n14039), .A(n11332), .ZN(P2_U3259) );
  INV_X1 U14003 ( .A(n11333), .ZN(n11336) );
  OAI222_X1 U14004 ( .A1(n13090), .A2(n11336), .B1(n13095), .B2(n11335), .C1(
        P3_U3151), .C2(n11334), .ZN(P3_U3275) );
  XOR2_X1 U14005 ( .A(n11337), .B(n12533), .Z(n11338) );
  AOI222_X1 U14006 ( .A1(n12576), .A2(n12982), .B1(n12986), .B2(n11338), .C1(
        n12574), .C2(n12981), .ZN(n11501) );
  INV_X1 U14007 ( .A(n11499), .ZN(n11504) );
  AOI22_X1 U14008 ( .A1(n11504), .A2(n13061), .B1(P3_REG0_REG_11__SCAN_IN), 
        .B2(n15653), .ZN(n11341) );
  XNOR2_X1 U14009 ( .A(n11339), .B(n12533), .ZN(n11500) );
  NAND2_X1 U14010 ( .A1(n11500), .A2(n11605), .ZN(n11340) );
  OAI211_X1 U14011 ( .C1(n11501), .C2(n15653), .A(n11341), .B(n11340), .ZN(
        P3_U3423) );
  NAND2_X1 U14012 ( .A1(n11402), .A2(n11345), .ZN(n11465) );
  NAND2_X1 U14013 ( .A1(n11342), .A2(n11465), .ZN(n11343) );
  NAND2_X1 U14014 ( .A1(n11406), .A2(n14553), .ZN(n11479) );
  XNOR2_X1 U14015 ( .A(n11343), .B(n11346), .ZN(n15321) );
  INV_X1 U14016 ( .A(n15269), .ZN(n14939) );
  AOI22_X1 U14017 ( .A1(n15008), .A2(n14554), .B1(n14552), .B2(n15010), .ZN(
        n11349) );
  NAND2_X1 U14018 ( .A1(n11480), .A2(n11346), .ZN(n11410) );
  OAI21_X1 U14019 ( .B1(n11480), .B2(n11346), .A(n11410), .ZN(n11347) );
  NAND2_X1 U14020 ( .A1(n11347), .A2(n15311), .ZN(n11348) );
  OAI211_X1 U14021 ( .C1(n15321), .C2(n15294), .A(n11349), .B(n11348), .ZN(
        n15325) );
  NAND2_X1 U14022 ( .A1(n15325), .A2(n14993), .ZN(n11357) );
  INV_X1 U14023 ( .A(n11415), .ZN(n11351) );
  AOI211_X1 U14024 ( .C1(n14319), .C2(n7457), .A(n15280), .B(n11351), .ZN(
        n15322) );
  NOR2_X1 U14025 ( .A1(n14994), .A2(n11406), .ZN(n11355) );
  OAI22_X1 U14026 ( .A1(n14993), .A2(n11353), .B1(n11352), .B2(n14977), .ZN(
        n11354) );
  AOI211_X1 U14027 ( .C1(n15322), .C2(n15268), .A(n11355), .B(n11354), .ZN(
        n11356) );
  OAI211_X1 U14028 ( .C1(n15321), .C2(n14939), .A(n11357), .B(n11356), .ZN(
        P1_U3287) );
  OAI21_X1 U14029 ( .B1(n7964), .B2(n8657), .A(n11358), .ZN(n14034) );
  XNOR2_X1 U14030 ( .A(n11359), .B(n11360), .ZN(n11363) );
  OR2_X1 U14031 ( .A1(n13343), .A2(n13273), .ZN(n11362) );
  NAND2_X1 U14032 ( .A1(n13603), .A2(n13880), .ZN(n11361) );
  NAND2_X1 U14033 ( .A1(n11362), .A2(n11361), .ZN(n12189) );
  AOI21_X1 U14034 ( .B1(n11363), .B2(n13897), .A(n12189), .ZN(n14033) );
  MUX2_X1 U14035 ( .A(n10356), .B(n14033), .S(n13913), .Z(n11369) );
  INV_X1 U14036 ( .A(n11364), .ZN(n11365) );
  AOI211_X1 U14037 ( .C1(n14031), .C2(n11365), .A(n6409), .B(n11583), .ZN(
        n14030) );
  OAI22_X1 U14038 ( .A1(n11366), .A2(n13904), .B1(n12192), .B2(n13843), .ZN(
        n11367) );
  AOI21_X1 U14039 ( .B1(n14030), .B2(n13919), .A(n11367), .ZN(n11368) );
  OAI211_X1 U14040 ( .C1(n13908), .C2(n14034), .A(n11369), .B(n11368), .ZN(
        P2_U3257) );
  XNOR2_X1 U14041 ( .A(n11627), .B(n11370), .ZN(n11374) );
  NAND2_X1 U14042 ( .A1(n11377), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n11371) );
  NAND2_X1 U14043 ( .A1(n11373), .A2(n11374), .ZN(n11629) );
  OAI21_X1 U14044 ( .B1(n11374), .B2(n11373), .A(n11629), .ZN(n11386) );
  INV_X1 U14045 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U14046 ( .A1(n14735), .A2(n11627), .ZN(n11375) );
  NAND2_X1 U14047 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n14126)
         );
  OAI211_X1 U14048 ( .C1(n14742), .C2(n11376), .A(n11375), .B(n14126), .ZN(
        n11385) );
  NAND2_X1 U14049 ( .A1(n11377), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U14050 ( .A1(n11379), .A2(n11378), .ZN(n11382) );
  INV_X1 U14051 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11380) );
  XNOR2_X1 U14052 ( .A(n11627), .B(n11380), .ZN(n11381) );
  NAND2_X1 U14053 ( .A1(n11382), .A2(n11381), .ZN(n11626) );
  OAI211_X1 U14054 ( .C1(n11382), .C2(n11381), .A(n11626), .B(n14737), .ZN(
        n11383) );
  INV_X1 U14055 ( .A(n11383), .ZN(n11384) );
  AOI211_X1 U14056 ( .C1(n11386), .C2(n14732), .A(n11385), .B(n11384), .ZN(
        n11387) );
  INV_X1 U14057 ( .A(n11387), .ZN(P1_U3257) );
  INV_X1 U14058 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n11689) );
  MUX2_X1 U14059 ( .A(n11689), .B(n11395), .S(n15665), .Z(n11389) );
  NAND2_X1 U14060 ( .A1(n11391), .A2(n10091), .ZN(n11388) );
  OAI211_X1 U14061 ( .C1(n12976), .C2(n11390), .A(n11389), .B(n11388), .ZN(
        P3_U3469) );
  INV_X1 U14062 ( .A(n11391), .ZN(n11398) );
  INV_X1 U14063 ( .A(n11392), .ZN(n11393) );
  AOI22_X1 U14064 ( .A1(n12913), .A2(n11394), .B1(n12912), .B2(n11393), .ZN(
        n11397) );
  MUX2_X1 U14065 ( .A(n11691), .B(n11395), .S(n15616), .Z(n11396) );
  OAI211_X1 U14066 ( .C1(n11398), .C2(n12922), .A(n11397), .B(n11396), .ZN(
        P3_U3223) );
  INV_X1 U14067 ( .A(n11465), .ZN(n11404) );
  NAND2_X1 U14068 ( .A1(n11401), .A2(n11402), .ZN(n11399) );
  NAND2_X1 U14069 ( .A1(n11399), .A2(n14313), .ZN(n11400) );
  OAI211_X1 U14070 ( .C1(n11402), .C2(n11401), .A(n14504), .B(n11400), .ZN(
        n11467) );
  INV_X1 U14071 ( .A(n11467), .ZN(n11403) );
  OAI21_X1 U14072 ( .B1(n15303), .B2(n11404), .A(n11403), .ZN(n11407) );
  NAND2_X1 U14073 ( .A1(n11406), .A2(n11405), .ZN(n11466) );
  NAND2_X1 U14074 ( .A1(n11407), .A2(n11466), .ZN(n11408) );
  INV_X1 U14075 ( .A(n14510), .ZN(n11469) );
  XNOR2_X1 U14076 ( .A(n11408), .B(n11469), .ZN(n15328) );
  INV_X1 U14077 ( .A(n15328), .ZN(n11422) );
  NAND2_X1 U14078 ( .A1(n11410), .A2(n11409), .ZN(n11411) );
  NAND2_X1 U14079 ( .A1(n11411), .A2(n14510), .ZN(n11522) );
  OAI21_X1 U14080 ( .B1(n11411), .B2(n14510), .A(n11522), .ZN(n11412) );
  NAND2_X1 U14081 ( .A1(n11412), .A2(n15311), .ZN(n11414) );
  AOI22_X1 U14082 ( .A1(n15008), .A2(n14553), .B1(n14551), .B2(n15010), .ZN(
        n11413) );
  NAND2_X1 U14083 ( .A1(n11414), .A2(n11413), .ZN(n15332) );
  AOI21_X1 U14084 ( .B1(n11415), .B2(n14325), .A(n15280), .ZN(n11416) );
  NAND2_X1 U14085 ( .A1(n11416), .A2(n11558), .ZN(n15329) );
  OAI22_X1 U14086 ( .A1(n14993), .A2(n11417), .B1(n14109), .B2(n14977), .ZN(
        n11418) );
  AOI21_X1 U14087 ( .B1(n15260), .B2(n14325), .A(n11418), .ZN(n11419) );
  OAI21_X1 U14088 ( .B1(n15329), .B2(n14982), .A(n11419), .ZN(n11420) );
  AOI21_X1 U14089 ( .B1(n15332), .B2(n14993), .A(n11420), .ZN(n11421) );
  OAI21_X1 U14090 ( .B1(n11929), .B2(n11422), .A(n11421), .ZN(P1_U3286) );
  XNOR2_X1 U14091 ( .A(n11499), .B(n6445), .ZN(n11639) );
  XOR2_X1 U14092 ( .A(n11637), .B(n11639), .Z(n11510) );
  XNOR2_X1 U14093 ( .A(n11510), .B(n12575), .ZN(n11429) );
  NAND2_X1 U14094 ( .A1(n12341), .A2(n12576), .ZN(n11425) );
  NAND2_X1 U14095 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n11702)
         );
  OAI211_X1 U14096 ( .C1(n12344), .C2(n11636), .A(n11425), .B(n11702), .ZN(
        n11427) );
  NOR2_X1 U14097 ( .A1(n11499), .A2(n12285), .ZN(n11426) );
  AOI211_X1 U14098 ( .C1(n11503), .C2(n12340), .A(n11427), .B(n11426), .ZN(
        n11428) );
  OAI21_X1 U14099 ( .B1(n11429), .B2(n12349), .A(n11428), .ZN(P3_U3176) );
  INV_X1 U14100 ( .A(n11436), .ZN(n12535) );
  XNOR2_X1 U14101 ( .A(n11430), .B(n12535), .ZN(n11434) );
  NAND2_X1 U14102 ( .A1(n12981), .A2(n12573), .ZN(n11432) );
  NAND2_X1 U14103 ( .A1(n12575), .A2(n12982), .ZN(n11431) );
  AND2_X1 U14104 ( .A1(n11432), .A2(n11431), .ZN(n11515) );
  INV_X1 U14105 ( .A(n11515), .ZN(n11433) );
  AOI21_X1 U14106 ( .B1(n11434), .B2(n12986), .A(n11433), .ZN(n11447) );
  OAI21_X1 U14107 ( .B1(n11437), .B2(n11436), .A(n11435), .ZN(n11445) );
  OAI22_X1 U14108 ( .A1(n11520), .A2(n12976), .B1(n15665), .B2(n12596), .ZN(
        n11438) );
  AOI21_X1 U14109 ( .B1(n11445), .B2(n10091), .A(n11438), .ZN(n11439) );
  OAI21_X1 U14110 ( .B1(n11447), .B2(n15663), .A(n11439), .ZN(P3_U3471) );
  OAI22_X1 U14111 ( .A1(n11520), .A2(n13070), .B1(n15654), .B2(n11440), .ZN(
        n11441) );
  AOI21_X1 U14112 ( .B1(n11445), .B2(n11605), .A(n11441), .ZN(n11442) );
  OAI21_X1 U14113 ( .B1(n11447), .B2(n15653), .A(n11442), .ZN(P3_U3426) );
  AOI22_X1 U14114 ( .A1(n15618), .A2(P3_REG2_REG_12__SCAN_IN), .B1(n12912), 
        .B2(n11517), .ZN(n11443) );
  OAI21_X1 U14115 ( .B1(n11520), .B2(n12828), .A(n11443), .ZN(n11444) );
  AOI21_X1 U14116 ( .B1(n11445), .B2(n12845), .A(n11444), .ZN(n11446) );
  OAI21_X1 U14117 ( .B1(n15618), .B2(n11447), .A(n11446), .ZN(P3_U3221) );
  INV_X1 U14118 ( .A(n11448), .ZN(n11453) );
  OR2_X1 U14119 ( .A1(n11449), .A2(P2_U3088), .ZN(n13577) );
  INV_X1 U14120 ( .A(n13577), .ZN(n13582) );
  AOI21_X1 U14121 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n14093), .A(n13582), 
        .ZN(n11450) );
  OAI21_X1 U14122 ( .B1(n11453), .B2(n14099), .A(n11450), .ZN(P2_U3304) );
  AOI21_X1 U14123 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n15186), .A(n11451), 
        .ZN(n11452) );
  OAI21_X1 U14124 ( .B1(n11453), .B2(n15195), .A(n11452), .ZN(P1_U3332) );
  INV_X1 U14125 ( .A(n11454), .ZN(n11456) );
  OAI222_X1 U14126 ( .A1(P1_U3086), .A2(n14482), .B1(n15192), .B2(n11456), 
        .C1(n11455), .C2(n15189), .ZN(P1_U3335) );
  OAI222_X1 U14127 ( .A1(n14102), .A2(n11457), .B1(P2_U3088), .B2(n13578), 
        .C1(n14099), .C2(n11456), .ZN(P2_U3307) );
  INV_X1 U14128 ( .A(n11458), .ZN(n11460) );
  INV_X1 U14129 ( .A(SI_21_), .ZN(n11459) );
  OAI222_X1 U14130 ( .A1(P3_U3151), .A2(n11461), .B1(n13090), .B2(n11460), 
        .C1(n11459), .C2(n13095), .ZN(P3_U3274) );
  NAND3_X1 U14131 ( .A1(n15030), .A2(n15029), .A3(n11462), .ZN(n11463) );
  AND2_X1 U14132 ( .A1(n14482), .A2(n14738), .ZN(n11464) );
  NAND2_X1 U14133 ( .A1(n14286), .A2(n11464), .ZN(n15320) );
  NAND2_X1 U14134 ( .A1(n11466), .A2(n11465), .ZN(n11470) );
  NAND2_X1 U14135 ( .A1(n11467), .A2(n11466), .ZN(n11468) );
  OR2_X1 U14136 ( .A1(n14325), .A2(n14552), .ZN(n11471) );
  INV_X1 U14137 ( .A(n14326), .ZN(n11523) );
  NAND2_X1 U14138 ( .A1(n15335), .A2(n14107), .ZN(n14327) );
  NAND2_X1 U14139 ( .A1(n11523), .A2(n14327), .ZN(n14318) );
  OR2_X1 U14140 ( .A1(n15335), .A2(n14551), .ZN(n14332) );
  NAND2_X1 U14141 ( .A1(n11472), .A2(n14332), .ZN(n11528) );
  XNOR2_X1 U14142 ( .A(n14344), .B(n14343), .ZN(n14508) );
  NAND2_X1 U14143 ( .A1(n11528), .A2(n14508), .ZN(n11474) );
  OR2_X1 U14144 ( .A1(n14344), .A2(n14550), .ZN(n11473) );
  NAND2_X1 U14145 ( .A1(n11474), .A2(n11473), .ZN(n11800) );
  XNOR2_X1 U14146 ( .A(n11800), .B(n11799), .ZN(n11550) );
  NAND2_X1 U14147 ( .A1(n14548), .A2(n15010), .ZN(n11539) );
  NAND2_X1 U14148 ( .A1(n14550), .A2(n15008), .ZN(n11541) );
  NAND2_X1 U14149 ( .A1(n11539), .A2(n11541), .ZN(n11882) );
  INV_X1 U14150 ( .A(n11530), .ZN(n11478) );
  INV_X1 U14151 ( .A(n14350), .ZN(n11543) );
  NAND2_X1 U14152 ( .A1(n11530), .A2(n11543), .ZN(n11796) );
  INV_X1 U14153 ( .A(n11796), .ZN(n11477) );
  AOI211_X1 U14154 ( .C1(n14350), .C2(n11478), .A(n15280), .B(n11477), .ZN(
        n11538) );
  AOI211_X1 U14155 ( .C1(n15336), .C2(n14350), .A(n11882), .B(n11538), .ZN(
        n11486) );
  NAND2_X1 U14156 ( .A1(n14510), .A2(n11481), .ZN(n11482) );
  INV_X1 U14157 ( .A(n14344), .ZN(n15345) );
  NAND2_X1 U14158 ( .A1(n11523), .A2(n14343), .ZN(n11483) );
  AOI22_X1 U14159 ( .A1(n15345), .A2(n11483), .B1(n14326), .B2(n14550), .ZN(
        n11484) );
  OAI211_X1 U14160 ( .C1(n11485), .C2(n11799), .A(n15311), .B(n11794), .ZN(
        n11542) );
  OAI211_X1 U14161 ( .C1(n15340), .C2(n11550), .A(n11486), .B(n11542), .ZN(
        n15158) );
  NAND2_X1 U14162 ( .A1(n15158), .A2(n15354), .ZN(n11487) );
  OAI21_X1 U14163 ( .B1(n15354), .B2(n9080), .A(n11487), .ZN(P1_U3489) );
  INV_X1 U14164 ( .A(n11488), .ZN(n11491) );
  OAI222_X1 U14165 ( .A1(n15189), .A2(n15767), .B1(n15192), .B2(n11491), .C1(
        P1_U3086), .C2(n11489), .ZN(P1_U3330) );
  OAI222_X1 U14166 ( .A1(n14102), .A2(n11492), .B1(n14099), .B2(n11491), .C1(
        P2_U3088), .C2(n11490), .ZN(P2_U3302) );
  INV_X1 U14167 ( .A(n11493), .ZN(n11508) );
  OAI222_X1 U14168 ( .A1(n15189), .A2(n11495), .B1(n15192), .B2(n11508), .C1(
        n11494), .C2(P1_U3086), .ZN(P1_U3334) );
  MUX2_X1 U14169 ( .A(n11496), .B(n11501), .S(n15665), .Z(n11498) );
  NAND2_X1 U14170 ( .A1(n11500), .A2(n10091), .ZN(n11497) );
  OAI211_X1 U14171 ( .C1(n12976), .C2(n11499), .A(n11498), .B(n11497), .ZN(
        P3_U3470) );
  INV_X1 U14172 ( .A(n11500), .ZN(n11507) );
  MUX2_X1 U14173 ( .A(n11502), .B(n11501), .S(n15616), .Z(n11506) );
  AOI22_X1 U14174 ( .A1(n11504), .A2(n12913), .B1(n12912), .B2(n11503), .ZN(
        n11505) );
  OAI211_X1 U14175 ( .C1(n11507), .C2(n12922), .A(n11506), .B(n11505), .ZN(
        P3_U3222) );
  OAI222_X1 U14176 ( .A1(n14102), .A2(n11509), .B1(P2_U3088), .B2(n13284), 
        .C1(n14099), .C2(n11508), .ZN(P2_U3306) );
  AOI22_X1 U14177 ( .A1(n11510), .A2(n12575), .B1(n11637), .B2(n11639), .ZN(
        n11512) );
  XOR2_X1 U14178 ( .A(n6445), .B(n11520), .Z(n11641) );
  XNOR2_X1 U14179 ( .A(n11641), .B(n12574), .ZN(n11511) );
  XNOR2_X1 U14180 ( .A(n11512), .B(n11511), .ZN(n11513) );
  NAND2_X1 U14181 ( .A1(n11513), .A2(n12308), .ZN(n11519) );
  OAI22_X1 U14182 ( .A1(n12313), .A2(n11515), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11514), .ZN(n11516) );
  AOI21_X1 U14183 ( .B1(n12340), .B2(n11517), .A(n11516), .ZN(n11518) );
  OAI211_X1 U14184 ( .C1(n12285), .C2(n11520), .A(n11519), .B(n11518), .ZN(
        P3_U3164) );
  NAND2_X1 U14185 ( .A1(n11522), .A2(n11521), .ZN(n11552) );
  OR2_X1 U14186 ( .A1(n11552), .A2(n14318), .ZN(n11554) );
  NAND2_X1 U14187 ( .A1(n11554), .A2(n11523), .ZN(n11524) );
  XNOR2_X1 U14188 ( .A(n11524), .B(n14508), .ZN(n11527) );
  NAND2_X1 U14189 ( .A1(n14549), .A2(n15010), .ZN(n11526) );
  NAND2_X1 U14190 ( .A1(n14551), .A2(n15008), .ZN(n11525) );
  NAND2_X1 U14191 ( .A1(n11526), .A2(n11525), .ZN(n11895) );
  AOI21_X1 U14192 ( .B1(n11527), .B2(n15311), .A(n11895), .ZN(n15352) );
  XNOR2_X1 U14193 ( .A(n11528), .B(n14508), .ZN(n15349) );
  NAND2_X1 U14194 ( .A1(n11556), .A2(n14344), .ZN(n11529) );
  NAND2_X1 U14195 ( .A1(n11529), .A2(n15264), .ZN(n11531) );
  OR2_X1 U14196 ( .A1(n11531), .A2(n11530), .ZN(n15343) );
  OAI22_X1 U14197 ( .A1(n14993), .A2(n11532), .B1(n11892), .B2(n14977), .ZN(
        n11533) );
  AOI21_X1 U14198 ( .B1(n15260), .B2(n14344), .A(n11533), .ZN(n11534) );
  OAI21_X1 U14199 ( .B1(n15343), .B2(n14982), .A(n11534), .ZN(n11535) );
  AOI21_X1 U14200 ( .B1(n15349), .B2(n11536), .A(n11535), .ZN(n11537) );
  OAI21_X1 U14201 ( .B1(n15352), .B2(n6408), .A(n11537), .ZN(P1_U3284) );
  INV_X1 U14202 ( .A(n11538), .ZN(n11540) );
  AOI21_X1 U14203 ( .B1(n11540), .B2(n11539), .A(n14982), .ZN(n11548) );
  AOI21_X1 U14204 ( .B1(n11542), .B2(n11541), .A(n6408), .ZN(n11547) );
  NOR2_X1 U14205 ( .A1(n11543), .A2(n14994), .ZN(n11546) );
  OAI22_X1 U14206 ( .A1(n14993), .A2(n11544), .B1(n11884), .B2(n14977), .ZN(
        n11545) );
  NOR4_X1 U14207 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11549) );
  OAI21_X1 U14208 ( .B1(n14925), .B2(n11550), .A(n11549), .ZN(P1_U3283) );
  INV_X1 U14209 ( .A(n14318), .ZN(n14511) );
  XNOR2_X1 U14210 ( .A(n11551), .B(n14511), .ZN(n15339) );
  AOI21_X1 U14211 ( .B1(n11552), .B2(n14318), .A(n15296), .ZN(n11555) );
  OAI22_X1 U14212 ( .A1(n11571), .A2(n14853), .B1(n14343), .B2(n14855), .ZN(
        n11553) );
  AOI21_X1 U14213 ( .B1(n11555), .B2(n11554), .A(n11553), .ZN(n15338) );
  MUX2_X1 U14214 ( .A(n15338), .B(n10485), .S(n6408), .Z(n11561) );
  INV_X1 U14215 ( .A(n11556), .ZN(n11557) );
  AOI211_X1 U14216 ( .C1(n15335), .C2(n11558), .A(n15280), .B(n11557), .ZN(
        n15334) );
  OAI22_X1 U14217 ( .A1(n11475), .A2(n14994), .B1(n14977), .B2(n11570), .ZN(
        n11559) );
  AOI21_X1 U14218 ( .B1(n15334), .B2(n15268), .A(n11559), .ZN(n11560) );
  OAI211_X1 U14219 ( .C1(n15339), .C2(n14925), .A(n11561), .B(n11560), .ZN(
        P1_U3285) );
  INV_X1 U14220 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n15731) );
  INV_X1 U14221 ( .A(n11562), .ZN(n11565) );
  OAI222_X1 U14222 ( .A1(n14102), .A2(n15731), .B1(n14099), .B2(n11565), .C1(
        P2_U3088), .C2(n11563), .ZN(P2_U3303) );
  OAI222_X1 U14223 ( .A1(n15189), .A2(n11566), .B1(n15192), .B2(n11565), .C1(
        P1_U3086), .C2(n11564), .ZN(P1_U3331) );
  AOI21_X1 U14224 ( .B1(n11569), .B2(n11568), .A(n11567), .ZN(n11575) );
  NAND2_X1 U14225 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n14646) );
  OAI21_X1 U14226 ( .B1(n14267), .B2(n14343), .A(n14646), .ZN(n11573) );
  OAI22_X1 U14227 ( .A1(n14255), .A2(n11571), .B1(n14279), .B2(n11570), .ZN(
        n11572) );
  AOI211_X1 U14228 ( .C1(n14269), .C2(n15335), .A(n11573), .B(n11572), .ZN(
        n11574) );
  OAI21_X1 U14229 ( .B1(n11575), .B2(n14271), .A(n11574), .ZN(P1_U3221) );
  NAND2_X1 U14230 ( .A1(n11358), .A2(n11576), .ZN(n11577) );
  INV_X1 U14231 ( .A(n13549), .ZN(n11579) );
  NAND2_X1 U14232 ( .A1(n11577), .A2(n11579), .ZN(n11713) );
  OAI21_X1 U14233 ( .B1(n11577), .B2(n11579), .A(n11713), .ZN(n11619) );
  XNOR2_X1 U14234 ( .A(n11578), .B(n11579), .ZN(n11582) );
  OR2_X1 U14235 ( .A1(n13358), .A2(n13274), .ZN(n11581) );
  OR2_X1 U14236 ( .A1(n13345), .A2(n13273), .ZN(n11580) );
  NAND2_X1 U14237 ( .A1(n11581), .A2(n11580), .ZN(n12159) );
  AOI21_X1 U14238 ( .B1(n11582), .B2(n13897), .A(n12159), .ZN(n11611) );
  OAI211_X1 U14239 ( .C1(n11614), .C2(n11583), .A(n6406), .B(n11719), .ZN(
        n11613) );
  OAI211_X1 U14240 ( .C1(n14040), .C2(n11619), .A(n11611), .B(n11613), .ZN(
        n11584) );
  INV_X1 U14241 ( .A(n11584), .ZN(n11587) );
  AOI22_X1 U14242 ( .A1(n14023), .A2(n13352), .B1(n15536), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n11585) );
  OAI21_X1 U14243 ( .B1(n11587), .B2(n15536), .A(n11585), .ZN(P2_U3508) );
  AOI22_X1 U14244 ( .A1(n14086), .A2(n13352), .B1(n15531), .B2(
        P2_REG0_REG_9__SCAN_IN), .ZN(n11586) );
  OAI21_X1 U14245 ( .B1(n11587), .B2(n15531), .A(n11586), .ZN(P2_U3457) );
  INV_X1 U14246 ( .A(n11588), .ZN(n11590) );
  OAI22_X1 U14247 ( .A1(n12560), .A2(P3_U3151), .B1(SI_22_), .B2(n13095), .ZN(
        n11589) );
  AOI21_X1 U14248 ( .B1(n11590), .B2(n11742), .A(n11589), .ZN(P3_U3273) );
  XNOR2_X1 U14249 ( .A(n11591), .B(n12536), .ZN(n11606) );
  INV_X1 U14250 ( .A(n11647), .ZN(n11592) );
  OAI22_X1 U14251 ( .A1(n11644), .A2(n12828), .B1(n11592), .B2(n15610), .ZN(
        n11593) );
  AOI21_X1 U14252 ( .B1(n11606), .B2(n12845), .A(n11593), .ZN(n11601) );
  OAI211_X1 U14253 ( .C1(n11596), .C2(n11595), .A(n11594), .B(n12986), .ZN(
        n11598) );
  AOI22_X1 U14254 ( .A1(n12572), .A2(n12981), .B1(n12982), .B2(n12574), .ZN(
        n11597) );
  AND2_X1 U14255 ( .A1(n11598), .A2(n11597), .ZN(n11608) );
  INV_X1 U14256 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n11599) );
  MUX2_X1 U14257 ( .A(n11608), .B(n11599), .S(n15618), .Z(n11600) );
  NAND2_X1 U14258 ( .A1(n11601), .A2(n11600), .ZN(P3_U3220) );
  NAND2_X1 U14259 ( .A1(n11606), .A2(n10091), .ZN(n11604) );
  INV_X1 U14260 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n11602) );
  MUX2_X1 U14261 ( .A(n11608), .B(n11602), .S(n15663), .Z(n11603) );
  OAI211_X1 U14262 ( .C1(n12976), .C2(n11644), .A(n11604), .B(n11603), .ZN(
        P3_U3472) );
  NAND2_X1 U14263 ( .A1(n11606), .A2(n11605), .ZN(n11610) );
  INV_X1 U14264 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n11607) );
  MUX2_X1 U14265 ( .A(n11608), .B(n11607), .S(n15653), .Z(n11609) );
  OAI211_X1 U14266 ( .C1(n13070), .C2(n11644), .A(n11610), .B(n11609), .ZN(
        P3_U3429) );
  MUX2_X1 U14267 ( .A(n11612), .B(n11611), .S(n13913), .Z(n11618) );
  INV_X1 U14268 ( .A(n11613), .ZN(n11616) );
  OAI22_X1 U14269 ( .A1(n11614), .A2(n13904), .B1(n13843), .B2(n12162), .ZN(
        n11615) );
  AOI21_X1 U14270 ( .B1(n11616), .B2(n13919), .A(n11615), .ZN(n11617) );
  OAI211_X1 U14271 ( .C1(n13908), .C2(n11619), .A(n11618), .B(n11617), .ZN(
        P2_U3256) );
  INV_X1 U14272 ( .A(n11620), .ZN(n11623) );
  OAI222_X1 U14273 ( .A1(P1_U3086), .A2(n11622), .B1(n15192), .B2(n11623), 
        .C1(n11621), .C2(n15189), .ZN(P1_U3329) );
  OAI222_X1 U14274 ( .A1(P2_U3088), .A2(n11624), .B1(n14099), .B2(n11623), 
        .C1(n15780), .C2(n14102), .ZN(P2_U3301) );
  NAND2_X1 U14275 ( .A1(n11627), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n11625) );
  NAND2_X1 U14276 ( .A1(n11626), .A2(n11625), .ZN(n11909) );
  XNOR2_X1 U14277 ( .A(n11909), .B(n11900), .ZN(n11907) );
  XNOR2_X1 U14278 ( .A(n11907), .B(P1_REG2_REG_15__SCAN_IN), .ZN(n11635) );
  OR2_X1 U14279 ( .A1(n11627), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n11628) );
  NAND2_X1 U14280 ( .A1(n11629), .A2(n11628), .ZN(n11901) );
  INV_X1 U14281 ( .A(n11900), .ZN(n11908) );
  XNOR2_X1 U14282 ( .A(n11899), .B(n11898), .ZN(n11630) );
  NAND2_X1 U14283 ( .A1(n11630), .A2(n14732), .ZN(n11634) );
  AND2_X1 U14284 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14281) );
  NOR2_X1 U14285 ( .A1(n14742), .A2(n11631), .ZN(n11632) );
  AOI211_X1 U14286 ( .C1(n14735), .C2(n11908), .A(n14281), .B(n11632), .ZN(
        n11633) );
  OAI211_X1 U14287 ( .C1(n11635), .C2(n14710), .A(n11634), .B(n11633), .ZN(
        P1_U3258) );
  OAI21_X1 U14288 ( .B1(n11639), .B2(n12575), .A(n12574), .ZN(n11640) );
  NOR2_X1 U14289 ( .A1(n11641), .A2(n11636), .ZN(n11638) );
  XNOR2_X1 U14290 ( .A(n11671), .B(n12573), .ZN(n11642) );
  XNOR2_X1 U14291 ( .A(n11644), .B(n6445), .ZN(n11672) );
  INV_X1 U14292 ( .A(n11672), .ZN(n11673) );
  XNOR2_X1 U14293 ( .A(n11642), .B(n11673), .ZN(n11649) );
  AOI22_X1 U14294 ( .A1(n12341), .A2(n12574), .B1(P3_REG3_REG_13__SCAN_IN), 
        .B2(P3_U3151), .ZN(n11643) );
  OAI21_X1 U14295 ( .B1(n11676), .B2(n12344), .A(n11643), .ZN(n11646) );
  NOR2_X1 U14296 ( .A1(n11644), .A2(n12285), .ZN(n11645) );
  AOI211_X1 U14297 ( .C1(n11647), .C2(n12340), .A(n11646), .B(n11645), .ZN(
        n11648) );
  OAI21_X1 U14298 ( .B1(n11649), .B2(n12349), .A(n11648), .ZN(P3_U3174) );
  NAND2_X1 U14299 ( .A1(n13603), .A2(n13878), .ZN(n11651) );
  NAND2_X1 U14300 ( .A1(n13601), .A2(n13880), .ZN(n11650) );
  NAND2_X1 U14301 ( .A1(n11651), .A2(n11650), .ZN(n11716) );
  NAND2_X1 U14302 ( .A1(n13275), .A2(n11716), .ZN(n11652) );
  NAND2_X1 U14303 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n15429)
         );
  OAI211_X1 U14304 ( .C1(n13277), .C2(n11720), .A(n11652), .B(n15429), .ZN(
        n11669) );
  XNOR2_X1 U14305 ( .A(n14026), .B(n13139), .ZN(n11653) );
  NOR2_X1 U14306 ( .A1(n13358), .A2(n6406), .ZN(n11654) );
  NAND2_X1 U14307 ( .A1(n11653), .A2(n11654), .ZN(n11952) );
  INV_X1 U14308 ( .A(n11653), .ZN(n12176) );
  INV_X1 U14309 ( .A(n11654), .ZN(n11655) );
  NAND2_X1 U14310 ( .A1(n12176), .A2(n11655), .ZN(n11656) );
  NAND2_X1 U14311 ( .A1(n11952), .A2(n11656), .ZN(n11667) );
  XNOR2_X1 U14312 ( .A(n14031), .B(n10936), .ZN(n12163) );
  NOR2_X1 U14313 ( .A1(n13345), .A2(n6406), .ZN(n11658) );
  XNOR2_X1 U14314 ( .A(n12163), .B(n11658), .ZN(n12188) );
  INV_X1 U14315 ( .A(n11658), .ZN(n11659) );
  NAND2_X1 U14316 ( .A1(n12163), .A2(n11659), .ZN(n11660) );
  XNOR2_X1 U14317 ( .A(n13352), .B(n13139), .ZN(n11661) );
  NAND2_X1 U14318 ( .A1(n13603), .A2(n6409), .ZN(n11662) );
  XNOR2_X1 U14319 ( .A(n11661), .B(n11662), .ZN(n12166) );
  INV_X1 U14320 ( .A(n11661), .ZN(n11663) );
  NAND2_X1 U14321 ( .A1(n11663), .A2(n11662), .ZN(n11664) );
  NAND2_X1 U14322 ( .A1(n12171), .A2(n11664), .ZN(n11666) );
  INV_X1 U14323 ( .A(n11954), .ZN(n12178) );
  AOI211_X1 U14324 ( .C1(n11667), .C2(n11666), .A(n13250), .B(n12178), .ZN(
        n11668) );
  AOI211_X1 U14325 ( .C1(n14026), .C2(n13280), .A(n11669), .B(n11668), .ZN(
        n11670) );
  INV_X1 U14326 ( .A(n11670), .ZN(P2_U3189) );
  XNOR2_X1 U14327 ( .A(n11675), .B(n6446), .ZN(n11823) );
  XNOR2_X1 U14328 ( .A(n11823), .B(n11676), .ZN(n11824) );
  XNOR2_X1 U14329 ( .A(n11825), .B(n11824), .ZN(n11684) );
  INV_X1 U14330 ( .A(n11786), .ZN(n11681) );
  OR2_X1 U14331 ( .A1(n11677), .A2(n12838), .ZN(n11679) );
  NAND2_X1 U14332 ( .A1(n12573), .A2(n12982), .ZN(n11678) );
  NAND2_X1 U14333 ( .A1(n11679), .A2(n11678), .ZN(n11777) );
  AND2_X1 U14334 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12635) );
  AOI21_X1 U14335 ( .B1(n12324), .B2(n11777), .A(n12635), .ZN(n11680) );
  OAI21_X1 U14336 ( .B1(n12321), .B2(n11681), .A(n11680), .ZN(n11682) );
  AOI21_X1 U14337 ( .B1(n11787), .B2(n12347), .A(n11682), .ZN(n11683) );
  OAI21_X1 U14338 ( .B1(n11684), .B2(n12349), .A(n11683), .ZN(P3_U3155) );
  NAND2_X1 U14339 ( .A1(n11685), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n11688) );
  NAND2_X1 U14340 ( .A1(n11686), .A2(n11694), .ZN(n11687) );
  NAND2_X1 U14341 ( .A1(n11688), .A2(n11687), .ZN(n15590) );
  XNOR2_X1 U14342 ( .A(n15597), .B(P3_REG1_REG_10__SCAN_IN), .ZN(n15589) );
  OR2_X1 U14343 ( .A1(n15597), .A2(n11689), .ZN(n11690) );
  XOR2_X1 U14344 ( .A(P3_REG1_REG_11__SCAN_IN), .B(n12594), .Z(n11708) );
  XNOR2_X1 U14345 ( .A(n15597), .B(n11691), .ZN(n15584) );
  OAI21_X1 U14346 ( .B1(P3_REG2_REG_11__SCAN_IN), .B2(n11693), .A(n12588), 
        .ZN(n11706) );
  MUX2_X1 U14347 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n7168), .Z(n12598) );
  XNOR2_X1 U14348 ( .A(n12598), .B(n12600), .ZN(n12601) );
  MUX2_X1 U14349 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n7168), .Z(n11699) );
  XNOR2_X1 U14350 ( .A(n11699), .B(n11698), .ZN(n15593) );
  XOR2_X1 U14351 ( .A(n12601), .B(n12602), .Z(n11700) );
  NOR2_X1 U14352 ( .A1(n11700), .A2(n15576), .ZN(n11705) );
  NAND2_X1 U14353 ( .A1(n15539), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11701) );
  OAI211_X1 U14354 ( .C1(n15549), .C2(n11703), .A(n11702), .B(n11701), .ZN(
        n11704) );
  AOI211_X1 U14355 ( .C1(n11706), .C2(n15586), .A(n11705), .B(n11704), .ZN(
        n11707) );
  OAI21_X1 U14356 ( .B1(n11708), .B2(n12730), .A(n11707), .ZN(P3_U3193) );
  NAND2_X1 U14357 ( .A1(n11710), .A2(n11709), .ZN(n13551) );
  XOR2_X1 U14358 ( .A(n11711), .B(n13551), .Z(n11717) );
  NAND2_X1 U14359 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  XNOR2_X1 U14360 ( .A(n11714), .B(n13551), .ZN(n14029) );
  AOI211_X1 U14361 ( .C1(n13897), .C2(n11717), .A(n11716), .B(n11715), .ZN(
        n14028) );
  INV_X1 U14362 ( .A(n11733), .ZN(n11718) );
  AOI211_X1 U14363 ( .C1(n14026), .C2(n11719), .A(n6409), .B(n11718), .ZN(
        n14025) );
  INV_X1 U14364 ( .A(n14026), .ZN(n11723) );
  INV_X1 U14365 ( .A(n11720), .ZN(n11721) );
  AOI22_X1 U14366 ( .A1(n13894), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n11721), 
        .B2(n13915), .ZN(n11722) );
  OAI21_X1 U14367 ( .B1(n11723), .B2(n13904), .A(n11722), .ZN(n11726) );
  NOR2_X1 U14368 ( .A1(n14029), .A2(n11724), .ZN(n11725) );
  AOI211_X1 U14369 ( .C1(n14025), .C2(n13919), .A(n11726), .B(n11725), .ZN(
        n11727) );
  OAI21_X1 U14370 ( .B1(n14028), .B2(n13894), .A(n11727), .ZN(P2_U3255) );
  XNOR2_X1 U14371 ( .A(n11728), .B(n11729), .ZN(n11837) );
  INV_X1 U14372 ( .A(n11837), .ZN(n11740) );
  XNOR2_X1 U14373 ( .A(n11730), .B(n6407), .ZN(n11732) );
  OAI22_X1 U14374 ( .A1(n13372), .A2(n13274), .B1(n13358), .B2(n13273), .ZN(
        n12172) );
  INV_X1 U14375 ( .A(n12172), .ZN(n11731) );
  OAI21_X1 U14376 ( .B1(n11732), .B2(n13836), .A(n11731), .ZN(n11835) );
  NAND2_X1 U14377 ( .A1(n11835), .A2(n13913), .ZN(n11739) );
  AOI211_X1 U14378 ( .C1(n13365), .C2(n11733), .A(n6409), .B(n11816), .ZN(
        n11836) );
  INV_X1 U14379 ( .A(n13365), .ZN(n11734) );
  NOR2_X1 U14380 ( .A1(n11734), .A2(n13904), .ZN(n11737) );
  OAI22_X1 U14381 ( .A1(n13913), .A2(n11735), .B1(n12175), .B2(n13843), .ZN(
        n11736) );
  AOI211_X1 U14382 ( .C1(n11836), .C2(n13919), .A(n11737), .B(n11736), .ZN(
        n11738) );
  OAI211_X1 U14383 ( .C1(n13908), .C2(n11740), .A(n11739), .B(n11738), .ZN(
        P2_U3254) );
  NAND2_X1 U14384 ( .A1(n12571), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11741) );
  OAI21_X1 U14385 ( .B1(n12374), .B2(n12571), .A(n11741), .ZN(P3_U3521) );
  NAND2_X1 U14386 ( .A1(n11743), .A2(n11742), .ZN(n11744) );
  OAI211_X1 U14387 ( .C1(n11745), .C2(n13095), .A(n11744), .B(n12559), .ZN(
        P3_U3272) );
  NAND2_X1 U14388 ( .A1(P2_U3088), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n13102)
         );
  OAI21_X1 U14389 ( .B1(n15500), .B2(n8780), .A(n13102), .ZN(n11750) );
  XOR2_X1 U14390 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n11754), .Z(n15438) );
  OAI21_X1 U14391 ( .B1(n11754), .B2(P2_REG1_REG_12__SCAN_IN), .A(n15436), 
        .ZN(n15452) );
  XNOR2_X1 U14392 ( .A(n15456), .B(P2_REG1_REG_13__SCAN_IN), .ZN(n15453) );
  NOR2_X1 U14393 ( .A1(n15452), .A2(n15453), .ZN(n15451) );
  XNOR2_X1 U14394 ( .A(n13649), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n11747) );
  AOI211_X1 U14395 ( .C1(n11748), .C2(n11747), .A(n15492), .B(n13648), .ZN(
        n11749) );
  AOI211_X1 U14396 ( .C1(n7441), .C2(n13649), .A(n11750), .B(n11749), .ZN(
        n11762) );
  OR2_X1 U14397 ( .A1(n11751), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n11752) );
  NAND2_X1 U14398 ( .A1(n11753), .A2(n11752), .ZN(n15440) );
  XNOR2_X1 U14399 ( .A(n11754), .B(n11755), .ZN(n15439) );
  NAND2_X1 U14400 ( .A1(n15440), .A2(n15439), .ZN(n11757) );
  NAND2_X1 U14401 ( .A1(n15433), .A2(n11755), .ZN(n11756) );
  NAND2_X1 U14402 ( .A1(n11757), .A2(n11756), .ZN(n15449) );
  XNOR2_X1 U14403 ( .A(n15456), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n15450) );
  NAND2_X1 U14404 ( .A1(n15456), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n11758) );
  NAND2_X1 U14405 ( .A1(n15446), .A2(n11758), .ZN(n13638) );
  XNOR2_X1 U14406 ( .A(n13638), .B(n11759), .ZN(n11760) );
  NAND2_X1 U14407 ( .A1(n11760), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n13640) );
  OAI211_X1 U14408 ( .C1(n11760), .C2(P2_REG2_REG_14__SCAN_IN), .A(n13640), 
        .B(n15486), .ZN(n11761) );
  NAND2_X1 U14409 ( .A1(n11762), .A2(n11761), .ZN(P2_U3228) );
  OAI211_X1 U14410 ( .C1(n11765), .C2(n11764), .A(n11763), .B(n12986), .ZN(
        n11766) );
  AOI22_X1 U14411 ( .A1(n12905), .A2(n12981), .B1(n12982), .B2(n12572), .ZN(
        n11830) );
  NAND2_X1 U14412 ( .A1(n11766), .A2(n11830), .ZN(n12972) );
  INV_X1 U14413 ( .A(n12972), .ZN(n11772) );
  OAI21_X1 U14414 ( .B1(n11768), .B2(n12538), .A(n11767), .ZN(n12973) );
  INV_X1 U14415 ( .A(n11826), .ZN(n13071) );
  AOI22_X1 U14416 ( .A1(n15618), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n12912), 
        .B2(n11832), .ZN(n11769) );
  OAI21_X1 U14417 ( .B1(n13071), .B2(n12828), .A(n11769), .ZN(n11770) );
  AOI21_X1 U14418 ( .B1(n12973), .B2(n12845), .A(n11770), .ZN(n11771) );
  OAI21_X1 U14419 ( .B1(n15618), .B2(n11772), .A(n11771), .ZN(P3_U3218) );
  INV_X1 U14420 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n15775) );
  NAND2_X1 U14421 ( .A1(n12795), .A2(P3_U3897), .ZN(n11773) );
  OAI21_X1 U14422 ( .B1(P3_U3897), .B2(n15775), .A(n11773), .ZN(P3_U3518) );
  XNOR2_X1 U14423 ( .A(n11774), .B(n12537), .ZN(n11792) );
  INV_X1 U14424 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n11780) );
  INV_X1 U14425 ( .A(n11775), .ZN(n11776) );
  AOI21_X1 U14426 ( .B1(n11776), .B2(n12537), .A(n12834), .ZN(n11779) );
  AOI21_X1 U14427 ( .B1(n11779), .B2(n11778), .A(n11777), .ZN(n11788) );
  MUX2_X1 U14428 ( .A(n11780), .B(n11788), .S(n15665), .Z(n11782) );
  NAND2_X1 U14429 ( .A1(n11787), .A2(n12968), .ZN(n11781) );
  OAI211_X1 U14430 ( .C1(n11792), .C2(n12971), .A(n11782), .B(n11781), .ZN(
        P3_U3473) );
  MUX2_X1 U14431 ( .A(n11783), .B(n11788), .S(n15654), .Z(n11785) );
  NAND2_X1 U14432 ( .A1(n11787), .A2(n13061), .ZN(n11784) );
  OAI211_X1 U14433 ( .C1(n11792), .C2(n13065), .A(n11785), .B(n11784), .ZN(
        P3_U3432) );
  AOI22_X1 U14434 ( .A1(n11787), .A2(n12913), .B1(n12912), .B2(n11786), .ZN(
        n11791) );
  INV_X1 U14435 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n11789) );
  MUX2_X1 U14436 ( .A(n11789), .B(n11788), .S(n15616), .Z(n11790) );
  OAI211_X1 U14437 ( .C1(n11792), .C2(n12922), .A(n11791), .B(n11790), .ZN(
        P3_U3219) );
  INV_X1 U14438 ( .A(n14549), .ZN(n11869) );
  OR2_X1 U14439 ( .A1(n14350), .A2(n11869), .ZN(n11793) );
  INV_X1 U14440 ( .A(n14548), .ZN(n11920) );
  XNOR2_X1 U14441 ( .A(n15154), .B(n11920), .ZN(n14513) );
  XNOR2_X1 U14442 ( .A(n11849), .B(n14513), .ZN(n11795) );
  AOI222_X1 U14443 ( .A1(n14549), .A2(n15008), .B1(n15311), .B2(n11795), .C1(
        n14547), .C2(n15010), .ZN(n15156) );
  AOI211_X1 U14444 ( .C1(n15154), .C2(n11796), .A(n15280), .B(n7459), .ZN(
        n15153) );
  INV_X1 U14445 ( .A(n15154), .ZN(n11873) );
  INV_X1 U14446 ( .A(n11868), .ZN(n11797) );
  AOI22_X1 U14447 ( .A1(n6408), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n11797), 
        .B2(n15262), .ZN(n11798) );
  OAI21_X1 U14448 ( .B1(n11873), .B2(n14994), .A(n11798), .ZN(n11804) );
  INV_X1 U14449 ( .A(n11799), .ZN(n14515) );
  NAND2_X1 U14450 ( .A1(n11800), .A2(n14515), .ZN(n11802) );
  OR2_X1 U14451 ( .A1(n14350), .A2(n14549), .ZN(n11801) );
  XOR2_X1 U14452 ( .A(n14513), .B(n11842), .Z(n15157) );
  NOR2_X1 U14453 ( .A1(n15157), .A2(n14925), .ZN(n11803) );
  AOI211_X1 U14454 ( .C1(n15153), .C2(n15268), .A(n11804), .B(n11803), .ZN(
        n11805) );
  OAI21_X1 U14455 ( .B1(n6408), .B2(n15156), .A(n11805), .ZN(P1_U3282) );
  INV_X1 U14456 ( .A(n11806), .ZN(n12204) );
  OAI222_X1 U14457 ( .A1(P1_U3086), .A2(n14573), .B1(n15195), .B2(n12204), 
        .C1(n11807), .C2(n15189), .ZN(P1_U3328) );
  INV_X1 U14458 ( .A(n13553), .ZN(n11808) );
  XNOR2_X1 U14459 ( .A(n11809), .B(n11808), .ZN(n14018) );
  INV_X1 U14460 ( .A(n14018), .ZN(n11822) );
  NAND2_X1 U14461 ( .A1(n11810), .A2(n13553), .ZN(n11811) );
  NAND3_X1 U14462 ( .A1(n11812), .A2(n13897), .A3(n11811), .ZN(n11815) );
  OR2_X1 U14463 ( .A1(n13552), .A2(n13274), .ZN(n11814) );
  NAND2_X1 U14464 ( .A1(n13601), .A2(n13878), .ZN(n11813) );
  AND2_X1 U14465 ( .A1(n11814), .A2(n11813), .ZN(n12079) );
  NAND2_X1 U14466 ( .A1(n11815), .A2(n12079), .ZN(n14021) );
  OR2_X1 U14467 ( .A1(n12080), .A2(n11816), .ZN(n11817) );
  AND3_X1 U14468 ( .A1(n11817), .A2(n6406), .A3(n13900), .ZN(n14019) );
  NAND2_X1 U14469 ( .A1(n14019), .A2(n13919), .ZN(n11819) );
  AOI22_X1 U14470 ( .A1(n13797), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n12083), 
        .B2(n13915), .ZN(n11818) );
  OAI211_X1 U14471 ( .C1(n12080), .C2(n13904), .A(n11819), .B(n11818), .ZN(
        n11820) );
  AOI21_X1 U14472 ( .B1(n14021), .B2(n13913), .A(n11820), .ZN(n11821) );
  OAI21_X1 U14473 ( .B1(n13908), .B2(n11822), .A(n11821), .ZN(P2_U3253) );
  XNOR2_X1 U14474 ( .A(n11826), .B(n6446), .ZN(n12207) );
  XNOR2_X1 U14475 ( .A(n12207), .B(n12918), .ZN(n11827) );
  OAI21_X1 U14476 ( .B1(n11828), .B2(n11827), .A(n12208), .ZN(n11829) );
  NAND2_X1 U14477 ( .A1(n11829), .A2(n12308), .ZN(n11834) );
  NAND2_X1 U14478 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n12666)
         );
  OAI21_X1 U14479 ( .B1(n11830), .B2(n12313), .A(n12666), .ZN(n11831) );
  AOI21_X1 U14480 ( .B1(n11832), .B2(n12340), .A(n11831), .ZN(n11833) );
  OAI211_X1 U14481 ( .C1(n13071), .C2(n12285), .A(n11834), .B(n11833), .ZN(
        P3_U3181) );
  AOI211_X1 U14482 ( .C1(n15522), .C2(n11837), .A(n11836), .B(n11835), .ZN(
        n11840) );
  AOI22_X1 U14483 ( .A1(n13365), .A2(n14023), .B1(P2_REG1_REG_11__SCAN_IN), 
        .B2(n15536), .ZN(n11838) );
  OAI21_X1 U14484 ( .B1(n11840), .B2(n15536), .A(n11838), .ZN(P2_U3510) );
  AOI22_X1 U14485 ( .A1(n13365), .A2(n14086), .B1(P2_REG0_REG_11__SCAN_IN), 
        .B2(n15531), .ZN(n11839) );
  OAI21_X1 U14486 ( .B1(n11840), .B2(n15531), .A(n11839), .ZN(P2_U3463) );
  NOR2_X1 U14487 ( .A1(n15154), .A2(n14548), .ZN(n11841) );
  NAND2_X1 U14488 ( .A1(n15154), .A2(n14548), .ZN(n11843) );
  XNOR2_X1 U14489 ( .A(n15149), .B(n14547), .ZN(n14516) );
  OR2_X1 U14490 ( .A1(n15149), .A2(n14547), .ZN(n11845) );
  XNOR2_X1 U14491 ( .A(n15144), .B(n15009), .ZN(n11852) );
  OAI21_X1 U14492 ( .B1(n11846), .B2(n7777), .A(n12121), .ZN(n11847) );
  INV_X1 U14493 ( .A(n11847), .ZN(n15147) );
  NAND2_X1 U14494 ( .A1(n15154), .A2(n11920), .ZN(n11848) );
  INV_X1 U14495 ( .A(n14547), .ZN(n11853) );
  AOI21_X1 U14496 ( .B1(n6631), .B2(n7777), .A(n15296), .ZN(n11854) );
  INV_X1 U14497 ( .A(n14546), .ZN(n12093) );
  OAI22_X1 U14498 ( .A1(n11853), .A2(n14853), .B1(n12093), .B2(n14855), .ZN(
        n14237) );
  AOI21_X1 U14499 ( .B1(n11854), .B2(n12092), .A(n14237), .ZN(n15146) );
  OAI21_X1 U14500 ( .B1(n14234), .B2(n14977), .A(n15146), .ZN(n11855) );
  NAND2_X1 U14501 ( .A1(n11855), .A2(n14993), .ZN(n11860) );
  INV_X1 U14502 ( .A(n11923), .ZN(n11856) );
  INV_X1 U14503 ( .A(n15144), .ZN(n14240) );
  AOI211_X1 U14504 ( .C1(n15144), .C2(n11856), .A(n15280), .B(n15015), .ZN(
        n15143) );
  OAI22_X1 U14505 ( .A1(n14240), .A2(n14994), .B1(n14993), .B2(n11857), .ZN(
        n11858) );
  AOI21_X1 U14506 ( .B1(n15143), .B2(n15268), .A(n11858), .ZN(n11859) );
  OAI211_X1 U14507 ( .C1(n15147), .C2(n14925), .A(n11860), .B(n11859), .ZN(
        P1_U3280) );
  INV_X1 U14508 ( .A(n11861), .ZN(n15194) );
  AOI21_X1 U14509 ( .B1(P1_DATAO_REG_28__SCAN_IN), .B2(n14093), .A(n11862), 
        .ZN(n11863) );
  OAI21_X1 U14510 ( .B1(n15194), .B2(n14099), .A(n11863), .ZN(P2_U3299) );
  OAI21_X1 U14511 ( .B1(n11866), .B2(n11865), .A(n11864), .ZN(n11867) );
  NAND2_X1 U14512 ( .A1(n11867), .A2(n14273), .ZN(n11872) );
  AND2_X1 U14513 ( .A1(P1_U3086), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n14678) );
  OAI22_X1 U14514 ( .A1(n14255), .A2(n11869), .B1(n14279), .B2(n11868), .ZN(
        n11870) );
  AOI211_X1 U14515 ( .C1(n14209), .C2(n14547), .A(n14678), .B(n11870), .ZN(
        n11871) );
  OAI211_X1 U14516 ( .C1(n11873), .C2(n14285), .A(n11872), .B(n11871), .ZN(
        P1_U3236) );
  NOR2_X1 U14517 ( .A1(n11875), .A2(n11874), .ZN(n11876) );
  AOI21_X1 U14518 ( .B1(n11875), .B2(n11874), .A(n11876), .ZN(n11889) );
  NAND2_X1 U14519 ( .A1(n11889), .A2(n11890), .ZN(n11888) );
  AOI21_X1 U14520 ( .B1(n11877), .B2(n11879), .A(n11876), .ZN(n11881) );
  INV_X1 U14521 ( .A(n11878), .ZN(n11880) );
  AOI22_X1 U14522 ( .A1(n11888), .A2(n11881), .B1(n11880), .B2(n11879), .ZN(
        n11887) );
  AOI22_X1 U14523 ( .A1(n11882), .A2(n14282), .B1(P1_REG3_REG_10__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11883) );
  OAI21_X1 U14524 ( .B1(n11884), .B2(n14279), .A(n11883), .ZN(n11885) );
  AOI21_X1 U14525 ( .B1(n14350), .B2(n14269), .A(n11885), .ZN(n11886) );
  OAI21_X1 U14526 ( .B1(n11887), .B2(n14271), .A(n11886), .ZN(P1_U3217) );
  OAI21_X1 U14527 ( .B1(n11890), .B2(n11889), .A(n11888), .ZN(n11891) );
  NAND2_X1 U14528 ( .A1(n11891), .A2(n14273), .ZN(n11897) );
  NAND2_X1 U14529 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n14663) );
  INV_X1 U14530 ( .A(n14663), .ZN(n11894) );
  NOR2_X1 U14531 ( .A1(n14279), .A2(n11892), .ZN(n11893) );
  AOI211_X1 U14532 ( .C1(n14282), .C2(n11895), .A(n11894), .B(n11893), .ZN(
        n11896) );
  OAI211_X1 U14533 ( .C1(n15345), .C2(n14285), .A(n11897), .B(n11896), .ZN(
        P1_U3231) );
  XNOR2_X1 U14534 ( .A(n14694), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U14535 ( .A1(n11899), .A2(n11898), .ZN(n11903) );
  NAND2_X1 U14536 ( .A1(n11901), .A2(n11900), .ZN(n11902) );
  NAND2_X1 U14537 ( .A1(n11903), .A2(n11902), .ZN(n11905) );
  INV_X1 U14538 ( .A(n14687), .ZN(n11904) );
  AOI211_X1 U14539 ( .C1(n11906), .C2(n11905), .A(n14733), .B(n11904), .ZN(
        n11919) );
  XNOR2_X1 U14540 ( .A(n14694), .B(P1_REG2_REG_16__SCAN_IN), .ZN(n11914) );
  NAND2_X1 U14541 ( .A1(n11907), .A2(n14992), .ZN(n11911) );
  OR2_X1 U14542 ( .A1(n11909), .A2(n11908), .ZN(n11910) );
  NAND2_X1 U14543 ( .A1(n11911), .A2(n11910), .ZN(n11913) );
  INV_X1 U14544 ( .A(n14696), .ZN(n11912) );
  AOI211_X1 U14545 ( .C1(n11914), .C2(n11913), .A(n14710), .B(n11912), .ZN(
        n11918) );
  NAND2_X1 U14546 ( .A1(n14735), .A2(n14694), .ZN(n11915) );
  NAND2_X1 U14547 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14195)
         );
  OAI211_X1 U14548 ( .C1(n14742), .C2(n11916), .A(n11915), .B(n14195), .ZN(
        n11917) );
  OR3_X1 U14549 ( .A1(n11919), .A2(n11918), .A3(n11917), .ZN(P1_U3259) );
  AOI21_X1 U14550 ( .B1(n11850), .B2(n11844), .A(n15296), .ZN(n11922) );
  INV_X1 U14551 ( .A(n15009), .ZN(n14127) );
  OAI22_X1 U14552 ( .A1(n11920), .A2(n14853), .B1(n14127), .B2(n14855), .ZN(
        n14174) );
  AOI21_X1 U14553 ( .B1(n11922), .B2(n11921), .A(n14174), .ZN(n15151) );
  AOI211_X1 U14554 ( .C1(n15149), .C2(n7953), .A(n15280), .B(n11923), .ZN(
        n15148) );
  INV_X1 U14555 ( .A(n15149), .ZN(n14177) );
  INV_X1 U14556 ( .A(n14171), .ZN(n11924) );
  AOI22_X1 U14557 ( .A1(n6408), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n11924), 
        .B2(n15262), .ZN(n11925) );
  OAI21_X1 U14558 ( .B1(n14177), .B2(n14994), .A(n11925), .ZN(n11931) );
  INV_X1 U14559 ( .A(n11926), .ZN(n11927) );
  AOI21_X1 U14560 ( .B1(n14516), .B2(n11928), .A(n11927), .ZN(n15152) );
  NOR2_X1 U14561 ( .A1(n15152), .A2(n11929), .ZN(n11930) );
  AOI211_X1 U14562 ( .C1(n15148), .C2(n15268), .A(n11931), .B(n11930), .ZN(
        n11932) );
  OAI21_X1 U14563 ( .B1(n6408), .B2(n15151), .A(n11932), .ZN(P1_U3281) );
  INV_X1 U14564 ( .A(SI_30_), .ZN(n11939) );
  AND2_X1 U14565 ( .A1(n15190), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11933) );
  NAND2_X1 U14566 ( .A1(n14101), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11935) );
  XNOR2_X1 U14567 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n11936) );
  INV_X1 U14568 ( .A(n12367), .ZN(n11938) );
  OAI222_X1 U14569 ( .A1(n13095), .A2(n11939), .B1(n13090), .B2(n11938), .C1(
        n11937), .C2(P3_U3151), .ZN(P3_U3265) );
  INV_X1 U14570 ( .A(n11940), .ZN(n11946) );
  INV_X1 U14571 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n11941) );
  OAI22_X1 U14572 ( .A1(n13143), .A2(n13843), .B1(n11941), .B2(n13913), .ZN(
        n11942) );
  AOI21_X1 U14573 ( .B1(n13456), .B2(n13917), .A(n11942), .ZN(n11943) );
  OAI21_X1 U14574 ( .B1(n11944), .B2(n13744), .A(n11943), .ZN(n11945) );
  AOI21_X1 U14575 ( .B1(n11946), .B2(n13913), .A(n11945), .ZN(n11947) );
  OAI21_X1 U14576 ( .B1(n13908), .B2(n11948), .A(n11947), .ZN(P2_U3237) );
  INV_X1 U14577 ( .A(n11949), .ZN(n11950) );
  OAI222_X1 U14578 ( .A1(n14102), .A2(n11951), .B1(n14099), .B2(n11950), .C1(
        n13294), .C2(P2_U3088), .ZN(P2_U3305) );
  NAND2_X1 U14579 ( .A1(n13720), .A2(n6409), .ZN(n12011) );
  INV_X1 U14580 ( .A(n12011), .ZN(n12014) );
  XNOR2_X1 U14581 ( .A(n13940), .B(n13139), .ZN(n12013) );
  XNOR2_X1 U14582 ( .A(n13956), .B(n10936), .ZN(n12000) );
  OR2_X1 U14583 ( .A1(n13437), .A2(n6405), .ZN(n13115) );
  XNOR2_X1 U14584 ( .A(n13365), .B(n13139), .ZN(n11955) );
  NAND2_X1 U14585 ( .A1(n13601), .A2(n6409), .ZN(n11956) );
  XNOR2_X1 U14586 ( .A(n11955), .B(n11956), .ZN(n12179) );
  INV_X1 U14587 ( .A(n11955), .ZN(n12085) );
  NAND2_X1 U14588 ( .A1(n12085), .A2(n11956), .ZN(n11957) );
  XNOR2_X1 U14589 ( .A(n14085), .B(n13139), .ZN(n11959) );
  NAND2_X1 U14590 ( .A1(n13600), .A2(n6409), .ZN(n11960) );
  XNOR2_X1 U14591 ( .A(n11959), .B(n11960), .ZN(n12084) );
  INV_X1 U14592 ( .A(n11959), .ZN(n11961) );
  NAND2_X1 U14593 ( .A1(n11961), .A2(n11960), .ZN(n11962) );
  XNOR2_X1 U14594 ( .A(n14014), .B(n13139), .ZN(n11963) );
  NOR2_X1 U14595 ( .A1(n13552), .A2(n6405), .ZN(n11964) );
  NAND2_X1 U14596 ( .A1(n11963), .A2(n11964), .ZN(n11967) );
  INV_X1 U14597 ( .A(n11963), .ZN(n13100) );
  INV_X1 U14598 ( .A(n11964), .ZN(n11965) );
  NAND2_X1 U14599 ( .A1(n13100), .A2(n11965), .ZN(n11966) );
  NAND2_X1 U14600 ( .A1(n11967), .A2(n11966), .ZN(n13214) );
  XNOR2_X1 U14601 ( .A(n14009), .B(n13139), .ZN(n11969) );
  NAND2_X1 U14602 ( .A1(n13599), .A2(n6409), .ZN(n11970) );
  XNOR2_X1 U14603 ( .A(n11969), .B(n11970), .ZN(n13108) );
  AND2_X1 U14604 ( .A1(n13108), .A2(n11967), .ZN(n11968) );
  INV_X1 U14605 ( .A(n11969), .ZN(n11971) );
  NAND2_X1 U14606 ( .A1(n11971), .A2(n11970), .ZN(n11972) );
  NOR2_X1 U14607 ( .A1(n13392), .A2(n6405), .ZN(n12063) );
  XNOR2_X1 U14608 ( .A(n13996), .B(n10936), .ZN(n12067) );
  NAND2_X1 U14609 ( .A1(n13598), .A2(n6409), .ZN(n12066) );
  NAND2_X1 U14610 ( .A1(n12067), .A2(n12066), .ZN(n11973) );
  OAI21_X1 U14611 ( .B1(n12062), .B2(n12063), .A(n11973), .ZN(n11977) );
  XNOR2_X1 U14612 ( .A(n14073), .B(n13139), .ZN(n11978) );
  NOR2_X1 U14613 ( .A1(n13409), .A2(n6405), .ZN(n11979) );
  XNOR2_X1 U14614 ( .A(n11978), .B(n11979), .ZN(n12069) );
  NAND3_X1 U14615 ( .A1(n12062), .A2(n11973), .A3(n12063), .ZN(n11974) );
  OAI21_X1 U14616 ( .B1(n12067), .B2(n12066), .A(n11974), .ZN(n11975) );
  NOR2_X1 U14617 ( .A1(n12069), .A2(n11975), .ZN(n11976) );
  INV_X1 U14618 ( .A(n11978), .ZN(n11981) );
  INV_X1 U14619 ( .A(n11979), .ZN(n11980) );
  XNOR2_X1 U14620 ( .A(n13821), .B(n13139), .ZN(n11982) );
  NOR2_X1 U14621 ( .A1(n13126), .A2(n6405), .ZN(n11983) );
  NAND2_X1 U14622 ( .A1(n11982), .A2(n11983), .ZN(n11986) );
  INV_X1 U14623 ( .A(n11982), .ZN(n13124) );
  INV_X1 U14624 ( .A(n11983), .ZN(n11984) );
  NAND2_X1 U14625 ( .A1(n13124), .A2(n11984), .ZN(n11985) );
  NAND2_X1 U14626 ( .A1(n11986), .A2(n11985), .ZN(n13251) );
  NAND2_X1 U14627 ( .A1(n13782), .A2(n6409), .ZN(n11989) );
  XNOR2_X1 U14628 ( .A(n11988), .B(n11989), .ZN(n13133) );
  XNOR2_X1 U14629 ( .A(n13972), .B(n10717), .ZN(n11990) );
  NAND2_X1 U14630 ( .A1(n13595), .A2(n6409), .ZN(n11991) );
  XNOR2_X1 U14631 ( .A(n11990), .B(n11991), .ZN(n13202) );
  INV_X1 U14632 ( .A(n11990), .ZN(n11992) );
  XNOR2_X1 U14633 ( .A(n13432), .B(n10717), .ZN(n11994) );
  NOR2_X1 U14634 ( .A1(n13430), .A2(n6406), .ZN(n11993) );
  XNOR2_X1 U14635 ( .A(n11994), .B(n11993), .ZN(n13153) );
  NAND2_X1 U14636 ( .A1(n11994), .A2(n11993), .ZN(n11995) );
  XNOR2_X1 U14637 ( .A(n14058), .B(n10717), .ZN(n11996) );
  NAND2_X1 U14638 ( .A1(n12000), .A2(n13437), .ZN(n11999) );
  NAND2_X1 U14639 ( .A1(n13594), .A2(n6409), .ZN(n13110) );
  INV_X1 U14640 ( .A(n13110), .ZN(n11998) );
  INV_X1 U14641 ( .A(n12000), .ZN(n13112) );
  INV_X1 U14642 ( .A(n13115), .ZN(n12001) );
  XNOR2_X1 U14643 ( .A(n13948), .B(n10717), .ZN(n13161) );
  NOR2_X1 U14644 ( .A1(n13475), .A2(n6406), .ZN(n12004) );
  NAND2_X1 U14645 ( .A1(n13161), .A2(n12004), .ZN(n12005) );
  OAI21_X1 U14646 ( .B1(n13161), .B2(n12004), .A(n12005), .ZN(n13180) );
  INV_X1 U14647 ( .A(n12005), .ZN(n12010) );
  XNOR2_X1 U14648 ( .A(n13722), .B(n10717), .ZN(n12006) );
  AND2_X1 U14649 ( .A1(n13592), .A2(n6409), .ZN(n12007) );
  NAND2_X1 U14650 ( .A1(n12006), .A2(n12007), .ZN(n12012) );
  INV_X1 U14651 ( .A(n12006), .ZN(n13258) );
  INV_X1 U14652 ( .A(n12007), .ZN(n12008) );
  NAND2_X1 U14653 ( .A1(n13258), .A2(n12008), .ZN(n12009) );
  AND2_X1 U14654 ( .A1(n12012), .A2(n12009), .ZN(n13162) );
  XNOR2_X1 U14655 ( .A(n12013), .B(n12011), .ZN(n13267) );
  XNOR2_X1 U14656 ( .A(n13933), .B(n10717), .ZN(n13136) );
  AND2_X1 U14657 ( .A1(n13591), .A2(n6409), .ZN(n12015) );
  NAND2_X1 U14658 ( .A1(n13136), .A2(n12015), .ZN(n13147) );
  OAI21_X1 U14659 ( .B1(n13136), .B2(n12015), .A(n13147), .ZN(n12016) );
  AOI22_X1 U14660 ( .A1(n13590), .A2(n13880), .B1(n13720), .B2(n13878), .ZN(
        n13688) );
  INV_X1 U14661 ( .A(n13692), .ZN(n12018) );
  AOI22_X1 U14662 ( .A1(n12018), .A2(n13261), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12019) );
  OAI21_X1 U14663 ( .B1(n13688), .B2(n13263), .A(n12019), .ZN(n12020) );
  INV_X1 U14664 ( .A(n12025), .ZN(P2_U3186) );
  INV_X1 U14665 ( .A(n15136), .ZN(n15014) );
  INV_X1 U14666 ( .A(n15109), .ZN(n14938) );
  AND2_X2 U14667 ( .A1(n14933), .A2(n14938), .ZN(n14934) );
  INV_X1 U14668 ( .A(n15104), .ZN(n14921) );
  INV_X1 U14669 ( .A(n15096), .ZN(n14903) );
  INV_X1 U14670 ( .A(n15078), .ZN(n14859) );
  INV_X1 U14671 ( .A(n14840), .ZN(n14843) );
  NAND2_X1 U14672 ( .A1(n14098), .A2(n8962), .ZN(n12027) );
  OR2_X1 U14673 ( .A1(n14476), .A2(n15190), .ZN(n12026) );
  INV_X1 U14674 ( .A(n14759), .ZN(n12040) );
  NAND2_X1 U14675 ( .A1(n12030), .A2(n12199), .ZN(n12031) );
  MUX2_X1 U14676 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n7875), .Z(n12032) );
  NAND2_X1 U14677 ( .A1(n12032), .A2(SI_30_), .ZN(n13445) );
  OAI21_X1 U14678 ( .B1(SI_30_), .B2(n12032), .A(n13445), .ZN(n12033) );
  NAND2_X1 U14679 ( .A1(n12034), .A2(n12033), .ZN(n12035) );
  INV_X1 U14680 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12203) );
  OR2_X1 U14681 ( .A1(n14476), .A2(n12203), .ZN(n12037) );
  INV_X1 U14682 ( .A(n14744), .ZN(n12039) );
  OAI211_X1 U14683 ( .C1(n12040), .C2(n15036), .A(n12039), .B(n15264), .ZN(
        n15035) );
  INV_X1 U14684 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n12044) );
  NAND2_X1 U14685 ( .A1(n14427), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n12043) );
  INV_X1 U14686 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n12041) );
  OR2_X1 U14687 ( .A1(n9079), .A2(n12041), .ZN(n12042) );
  OAI211_X1 U14688 ( .C1(n14432), .C2(n12044), .A(n12043), .B(n12042), .ZN(
        n14540) );
  NAND2_X1 U14689 ( .A1(n15245), .A2(P1_B_REG_SCAN_IN), .ZN(n12045) );
  AND2_X1 U14690 ( .A1(n15010), .A2(n12045), .ZN(n14763) );
  NAND2_X1 U14691 ( .A1(n14540), .A2(n14763), .ZN(n15034) );
  NOR2_X1 U14692 ( .A1(n6408), .A2(n15034), .ZN(n14747) );
  NOR2_X1 U14693 ( .A1(n15036), .A2(n14994), .ZN(n12046) );
  AOI211_X1 U14694 ( .C1(n6408), .C2(P1_REG2_REG_30__SCAN_IN), .A(n14747), .B(
        n12046), .ZN(n12047) );
  OAI21_X1 U14695 ( .B1(n15035), .B2(n14982), .A(n12047), .ZN(P1_U3264) );
  OAI21_X1 U14696 ( .B1(n12049), .B2(n13558), .A(n12048), .ZN(n13959) );
  NAND2_X1 U14697 ( .A1(n12050), .A2(n13558), .ZN(n12051) );
  NAND3_X1 U14698 ( .A1(n12052), .A2(n13897), .A3(n12051), .ZN(n12055) );
  OR2_X1 U14699 ( .A1(n13437), .A2(n13274), .ZN(n12054) );
  NAND2_X1 U14700 ( .A1(n13783), .A2(n13878), .ZN(n12053) );
  AND2_X1 U14701 ( .A1(n12054), .A2(n12053), .ZN(n13222) );
  NAND2_X1 U14702 ( .A1(n12055), .A2(n13222), .ZN(n13961) );
  OAI21_X1 U14703 ( .B1(n13770), .B2(n13228), .A(n6406), .ZN(n12056) );
  OR2_X1 U14704 ( .A1(n13753), .A2(n12056), .ZN(n13960) );
  INV_X1 U14705 ( .A(n12057), .ZN(n13224) );
  AOI22_X1 U14706 ( .A1(n13224), .A2(n13915), .B1(P2_REG2_REG_22__SCAN_IN), 
        .B2(n13797), .ZN(n12059) );
  NAND2_X1 U14707 ( .A1(n14058), .A2(n13917), .ZN(n12058) );
  OAI211_X1 U14708 ( .C1(n13960), .C2(n13744), .A(n12059), .B(n12058), .ZN(
        n12060) );
  AOI21_X1 U14709 ( .B1(n13961), .B2(n13913), .A(n12060), .ZN(n12061) );
  OAI21_X1 U14710 ( .B1(n13908), .B2(n13959), .A(n12061), .ZN(P2_U3243) );
  INV_X1 U14711 ( .A(n12062), .ZN(n12065) );
  XNOR2_X1 U14712 ( .A(n12064), .B(n12062), .ZN(n13271) );
  NAND2_X1 U14713 ( .A1(n13271), .A2(n12063), .ZN(n13272) );
  OAI21_X1 U14714 ( .B1(n12065), .B2(n12064), .A(n13272), .ZN(n13170) );
  XNOR2_X1 U14715 ( .A(n12067), .B(n12066), .ZN(n13171) );
  NOR2_X1 U14716 ( .A1(n13170), .A2(n13171), .ZN(n13169) );
  INV_X1 U14717 ( .A(n13169), .ZN(n12070) );
  OAI22_X1 U14718 ( .A1(n12067), .A2(n13250), .B1(n13397), .B2(n13256), .ZN(
        n12068) );
  NAND3_X1 U14719 ( .A1(n12070), .A2(n12069), .A3(n12068), .ZN(n12076) );
  NOR2_X1 U14720 ( .A1(n13397), .A2(n13273), .ZN(n12071) );
  AOI21_X1 U14721 ( .B1(n13596), .B2(n13880), .A(n12071), .ZN(n13838) );
  INV_X1 U14722 ( .A(n13838), .ZN(n12072) );
  AOI22_X1 U14723 ( .A1(n12072), .A2(n13275), .B1(P2_REG3_REG_17__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12073) );
  OAI21_X1 U14724 ( .B1(n13844), .B2(n13277), .A(n12073), .ZN(n12074) );
  AOI21_X1 U14725 ( .B1(n14073), .B2(n13280), .A(n12074), .ZN(n12075) );
  OAI211_X1 U14726 ( .C1(n12077), .C2(n13250), .A(n12076), .B(n12075), .ZN(
        P2_U3200) );
  OAI22_X1 U14727 ( .A1(n13263), .A2(n12079), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12078), .ZN(n12082) );
  NOR2_X1 U14728 ( .A1(n12080), .A2(n13227), .ZN(n12081) );
  AOI211_X1 U14729 ( .C1(n13261), .C2(n12083), .A(n12082), .B(n12081), .ZN(
        n12089) );
  INV_X1 U14730 ( .A(n12084), .ZN(n12087) );
  OAI22_X1 U14731 ( .A1(n12085), .A2(n13250), .B1(n13367), .B2(n13256), .ZN(
        n12086) );
  NAND3_X1 U14732 ( .A1(n12184), .A2(n12087), .A3(n12086), .ZN(n12088) );
  OAI211_X1 U14733 ( .C1(n12090), .C2(n13250), .A(n12089), .B(n12088), .ZN(
        P2_U3196) );
  OR2_X1 U14734 ( .A1(n15144), .A2(n14127), .ZN(n12091) );
  NAND2_X1 U14735 ( .A1(n15136), .A2(n12093), .ZN(n14362) );
  NAND2_X1 U14736 ( .A1(n15130), .A2(n14370), .ZN(n14368) );
  NAND2_X1 U14737 ( .A1(n15122), .A2(n14384), .ZN(n12096) );
  OR2_X1 U14738 ( .A1(n15122), .A2(n14384), .ZN(n12094) );
  NAND2_X1 U14739 ( .A1(n12096), .A2(n12094), .ZN(n14973) );
  INV_X1 U14740 ( .A(n14969), .ZN(n14254) );
  OR2_X1 U14741 ( .A1(n14960), .A2(n14254), .ZN(n14390) );
  NAND2_X1 U14742 ( .A1(n14960), .A2(n14254), .ZN(n14943) );
  OR2_X1 U14743 ( .A1(n15109), .A2(n14956), .ZN(n12129) );
  NAND2_X1 U14744 ( .A1(n15109), .A2(n14956), .ZN(n12128) );
  INV_X1 U14745 ( .A(n14956), .ZN(n14155) );
  OR2_X1 U14746 ( .A1(n15109), .A2(n14155), .ZN(n12097) );
  INV_X1 U14747 ( .A(n14929), .ZN(n14253) );
  OR2_X1 U14748 ( .A1(n15104), .A2(n14253), .ZN(n14401) );
  NAND2_X1 U14749 ( .A1(n15104), .A2(n14253), .ZN(n14402) );
  NAND2_X1 U14750 ( .A1(n14401), .A2(n14402), .ZN(n14912) );
  INV_X1 U14751 ( .A(n14545), .ZN(n14405) );
  OR2_X1 U14752 ( .A1(n15096), .A2(n14405), .ZN(n12098) );
  XNOR2_X1 U14753 ( .A(n14891), .B(n14544), .ZN(n12132) );
  NAND2_X1 U14754 ( .A1(n14880), .A2(n12132), .ZN(n12100) );
  INV_X1 U14755 ( .A(n14544), .ZN(n14224) );
  OR2_X1 U14756 ( .A1(n14891), .A2(n14224), .ZN(n12099) );
  NAND2_X1 U14757 ( .A1(n14877), .A2(n14543), .ZN(n12101) );
  INV_X1 U14758 ( .A(n14869), .ZN(n12102) );
  XNOR2_X1 U14759 ( .A(n15078), .B(n14832), .ZN(n14860) );
  INV_X1 U14760 ( .A(n14832), .ZN(n12103) );
  NAND2_X1 U14761 ( .A1(n15078), .A2(n12103), .ZN(n12107) );
  INV_X1 U14762 ( .A(n14542), .ZN(n14854) );
  OR2_X1 U14763 ( .A1(n14840), .A2(n14854), .ZN(n12104) );
  NOR2_X1 U14764 ( .A1(n15065), .A2(n14216), .ZN(n12112) );
  INV_X1 U14765 ( .A(n12112), .ZN(n12105) );
  NAND2_X1 U14766 ( .A1(n15065), .A2(n14216), .ZN(n12110) );
  NAND2_X1 U14767 ( .A1(n12105), .A2(n12110), .ZN(n14812) );
  NAND2_X1 U14768 ( .A1(n15060), .A2(n14793), .ZN(n14796) );
  OR2_X1 U14769 ( .A1(n15060), .A2(n14793), .ZN(n12106) );
  NAND2_X1 U14770 ( .A1(n14755), .A2(n12110), .ZN(n12114) );
  NAND2_X1 U14771 ( .A1(n14840), .A2(n14854), .ZN(n12108) );
  AND3_X1 U14772 ( .A1(n12108), .A2(n12110), .A3(n12107), .ZN(n12109) );
  NAND2_X1 U14773 ( .A1(n12110), .A2(n14542), .ZN(n12111) );
  NOR2_X1 U14774 ( .A1(n14840), .A2(n12111), .ZN(n12113) );
  OAI21_X1 U14775 ( .B1(n14814), .B2(n12114), .A(n14749), .ZN(n12118) );
  AOI211_X1 U14776 ( .C1(n15060), .C2(n14819), .A(n15280), .B(n6497), .ZN(
        n15059) );
  AOI22_X1 U14777 ( .A1(n14263), .A2(n15262), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n6408), .ZN(n12119) );
  OAI21_X1 U14778 ( .B1(n7470), .B2(n14994), .A(n12119), .ZN(n12140) );
  OR2_X1 U14779 ( .A1(n15144), .A2(n15009), .ZN(n12120) );
  NAND2_X1 U14780 ( .A1(n15136), .A2(n14546), .ZN(n12122) );
  NAND3_X1 U14781 ( .A1(n15005), .A2(n14998), .A3(n12122), .ZN(n12125) );
  NAND2_X1 U14782 ( .A1(n14371), .A2(n14362), .ZN(n14361) );
  INV_X1 U14783 ( .A(n12122), .ZN(n14997) );
  NOR2_X1 U14784 ( .A1(n14361), .A2(n14997), .ZN(n12123) );
  INV_X1 U14785 ( .A(n15130), .ZN(n14995) );
  AOI22_X1 U14786 ( .A1(n14998), .A2(n12123), .B1(n14995), .B2(n14370), .ZN(
        n12124) );
  NAND2_X1 U14787 ( .A1(n12125), .A2(n12124), .ZN(n14972) );
  NAND2_X1 U14788 ( .A1(n15122), .A2(n14954), .ZN(n12126) );
  OR2_X1 U14789 ( .A1(n15122), .A2(n14954), .ZN(n12127) );
  NOR2_X1 U14790 ( .A1(n14960), .A2(n14969), .ZN(n14382) );
  NAND2_X1 U14791 ( .A1(n14960), .A2(n14969), .ZN(n14380) );
  INV_X1 U14792 ( .A(n12128), .ZN(n12130) );
  OR2_X1 U14793 ( .A1(n15104), .A2(n14929), .ZN(n12131) );
  INV_X1 U14794 ( .A(n12132), .ZN(n14887) );
  NAND2_X1 U14795 ( .A1(n15096), .A2(n14545), .ZN(n14884) );
  NAND2_X1 U14796 ( .A1(n14877), .A2(n14852), .ZN(n12134) );
  NOR2_X1 U14797 ( .A1(n15078), .A2(n14832), .ZN(n12137) );
  NAND2_X1 U14798 ( .A1(n15078), .A2(n14832), .ZN(n12136) );
  INV_X1 U14799 ( .A(n14812), .ZN(n14815) );
  AND2_X1 U14800 ( .A1(n15065), .A2(n14833), .ZN(n14754) );
  NOR2_X1 U14801 ( .A1(n14818), .A2(n14754), .ZN(n12138) );
  XOR2_X1 U14802 ( .A(n12138), .B(n14755), .Z(n15058) );
  NOR2_X1 U14803 ( .A1(n15058), .A2(n14925), .ZN(n12139) );
  AOI211_X1 U14804 ( .C1(n15059), .C2(n15268), .A(n12140), .B(n12139), .ZN(
        n12141) );
  OAI21_X1 U14805 ( .B1(n6408), .B2(n15063), .A(n12141), .ZN(P1_U3267) );
  INV_X1 U14806 ( .A(n14086), .ZN(n14079) );
  OR2_X1 U14807 ( .A1(n12151), .A2(n12142), .ZN(n12143) );
  NAND2_X1 U14808 ( .A1(n12144), .A2(n12143), .ZN(n13920) );
  NAND2_X1 U14809 ( .A1(n13916), .A2(n13296), .ZN(n12145) );
  NAND2_X1 U14810 ( .A1(n12145), .A2(n6405), .ZN(n12146) );
  NOR2_X1 U14811 ( .A1(n12147), .A2(n12146), .ZN(n13918) );
  INV_X1 U14812 ( .A(n12148), .ZN(n12149) );
  AOI21_X1 U14813 ( .B1(n12151), .B2(n12150), .A(n12149), .ZN(n12155) );
  NAND2_X1 U14814 ( .A1(n13920), .A2(n12152), .ZN(n12153) );
  OAI211_X1 U14815 ( .C1(n12155), .C2(n13836), .A(n12154), .B(n12153), .ZN(
        n13912) );
  AOI211_X1 U14816 ( .C1(n7492), .C2(n13920), .A(n13918), .B(n13912), .ZN(
        n12157) );
  MUX2_X1 U14817 ( .A(n7991), .B(n12157), .S(n15533), .Z(n12156) );
  OAI21_X1 U14818 ( .B1(n7216), .B2(n14079), .A(n12156), .ZN(P2_U3433) );
  INV_X1 U14819 ( .A(n14023), .ZN(n14007) );
  MUX2_X1 U14820 ( .A(n7995), .B(n12157), .S(n15538), .Z(n12158) );
  OAI21_X1 U14821 ( .B1(n7216), .B2(n14007), .A(n12158), .ZN(P2_U3500) );
  NAND2_X1 U14822 ( .A1(n13275), .A2(n12159), .ZN(n12161) );
  OAI211_X1 U14823 ( .C1(n13277), .C2(n12162), .A(n12161), .B(n12160), .ZN(
        n12169) );
  INV_X1 U14824 ( .A(n12197), .ZN(n12167) );
  INV_X1 U14825 ( .A(n12163), .ZN(n12164) );
  AOI22_X1 U14826 ( .A1(n13269), .A2(n13604), .B1(n13270), .B2(n12164), .ZN(
        n12165) );
  NOR3_X1 U14827 ( .A1(n12167), .A2(n12166), .A3(n12165), .ZN(n12168) );
  AOI211_X1 U14828 ( .C1(n13352), .C2(n13280), .A(n12169), .B(n12168), .ZN(
        n12170) );
  OAI21_X1 U14829 ( .B1(n13250), .B2(n12171), .A(n12170), .ZN(P2_U3203) );
  NAND2_X1 U14830 ( .A1(n13275), .A2(n12172), .ZN(n12174) );
  OAI211_X1 U14831 ( .C1(n13277), .C2(n12175), .A(n12174), .B(n12173), .ZN(
        n12182) );
  NOR3_X1 U14832 ( .A1(n12176), .A2(n13358), .A3(n13256), .ZN(n12177) );
  AOI21_X1 U14833 ( .B1(n12178), .B2(n13270), .A(n12177), .ZN(n12180) );
  NOR2_X1 U14834 ( .A1(n12180), .A2(n12179), .ZN(n12181) );
  AOI211_X1 U14835 ( .C1(n13365), .C2(n13280), .A(n12182), .B(n12181), .ZN(
        n12183) );
  OAI21_X1 U14836 ( .B1(n13250), .B2(n12184), .A(n12183), .ZN(P2_U3208) );
  NAND3_X1 U14837 ( .A1(n13269), .A2(n13605), .A3(n12185), .ZN(n12186) );
  OAI21_X1 U14838 ( .B1(n12187), .B2(n13250), .A(n12186), .ZN(n12195) );
  INV_X1 U14839 ( .A(n12188), .ZN(n12194) );
  NAND2_X1 U14840 ( .A1(n13280), .A2(n14031), .ZN(n12191) );
  AOI22_X1 U14841 ( .A1(n13275), .A2(n12189), .B1(P2_REG3_REG_8__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12190) );
  OAI211_X1 U14842 ( .C1(n13277), .C2(n12192), .A(n12191), .B(n12190), .ZN(
        n12193) );
  AOI21_X1 U14843 ( .B1(n12195), .B2(n12194), .A(n12193), .ZN(n12196) );
  OAI21_X1 U14844 ( .B1(n13250), .B2(n12197), .A(n12196), .ZN(P2_U3193) );
  INV_X1 U14845 ( .A(n12198), .ZN(n12200) );
  OAI222_X1 U14846 ( .A1(n15189), .A2(n12203), .B1(P1_U3086), .B2(n12202), 
        .C1(n15192), .C2(n14095), .ZN(P1_U3325) );
  OAI222_X1 U14847 ( .A1(n14102), .A2(n12206), .B1(P2_U3088), .B2(n12205), 
        .C1(n14099), .C2(n12204), .ZN(P2_U3300) );
  XNOR2_X1 U14848 ( .A(n12932), .B(n6445), .ZN(n12250) );
  XNOR2_X1 U14849 ( .A(n12250), .B(n12795), .ZN(n12251) );
  XNOR2_X1 U14850 ( .A(n13008), .B(n6446), .ZN(n12227) );
  INV_X1 U14851 ( .A(n12227), .ZN(n12229) );
  XNOR2_X1 U14852 ( .A(n13044), .B(n6446), .ZN(n12214) );
  XNOR2_X1 U14853 ( .A(n12286), .B(n6445), .ZN(n12210) );
  INV_X1 U14854 ( .A(n12207), .ZN(n12209) );
  XNOR2_X1 U14855 ( .A(n12210), .B(n12905), .ZN(n12278) );
  XNOR2_X1 U14856 ( .A(n13056), .B(n6446), .ZN(n12211) );
  XNOR2_X1 U14857 ( .A(n12211), .B(n12281), .ZN(n12287) );
  XOR2_X1 U14858 ( .A(n6445), .B(n13050), .Z(n12329) );
  INV_X1 U14859 ( .A(n12329), .ZN(n12212) );
  NOR2_X1 U14860 ( .A1(n12212), .A2(n12328), .ZN(n12213) );
  XNOR2_X1 U14861 ( .A(n12214), .B(n12333), .ZN(n12241) );
  XNOR2_X1 U14862 ( .A(n13038), .B(n6446), .ZN(n12215) );
  XNOR2_X1 U14863 ( .A(n12215), .B(n12887), .ZN(n12310) );
  XNOR2_X1 U14864 ( .A(n13032), .B(n6445), .ZN(n12217) );
  XNOR2_X1 U14865 ( .A(n12217), .B(n12320), .ZN(n12261) );
  INV_X1 U14866 ( .A(n12217), .ZN(n12218) );
  XOR2_X1 U14867 ( .A(n6445), .B(n13027), .Z(n12317) );
  XNOR2_X1 U14868 ( .A(n12941), .B(n6446), .ZN(n12300) );
  XNOR2_X1 U14869 ( .A(n12944), .B(n12220), .ZN(n12235) );
  AOI22_X1 U14870 ( .A1(n12300), .A2(n12567), .B1(n12235), .B2(n12568), .ZN(
        n12224) );
  INV_X1 U14871 ( .A(n12235), .ZN(n12297) );
  AOI21_X1 U14872 ( .B1(n12297), .B2(n12821), .A(n12839), .ZN(n12222) );
  NAND3_X1 U14873 ( .A1(n12297), .A2(n12821), .A3(n12839), .ZN(n12221) );
  OAI21_X1 U14874 ( .B1(n12300), .B2(n12222), .A(n12221), .ZN(n12223) );
  XNOR2_X1 U14875 ( .A(n12803), .B(n6445), .ZN(n12226) );
  XNOR2_X1 U14876 ( .A(n12226), .B(n12822), .ZN(n12268) );
  XNOR2_X1 U14877 ( .A(n12227), .B(n12566), .ZN(n12339) );
  OAI21_X1 U14878 ( .B1(n12229), .B2(n12566), .A(n12228), .ZN(n12252) );
  XOR2_X1 U14879 ( .A(n12251), .B(n12252), .Z(n12234) );
  OAI22_X1 U14880 ( .A1(n12230), .A2(n12838), .B1(n12269), .B2(n12836), .ZN(
        n12784) );
  AOI22_X1 U14881 ( .A1(n12785), .A2(n12340), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12231) );
  OAI21_X1 U14882 ( .B1(n7227), .B2(n12313), .A(n12231), .ZN(n12232) );
  AOI21_X1 U14883 ( .B1(n12932), .B2(n12347), .A(n12232), .ZN(n12233) );
  OAI21_X1 U14884 ( .B1(n12234), .B2(n12349), .A(n12233), .ZN(P3_U3154) );
  XNOR2_X1 U14885 ( .A(n12299), .B(n12568), .ZN(n12240) );
  AOI22_X1 U14886 ( .A1(n12569), .A2(n12341), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12237) );
  NAND2_X1 U14887 ( .A1(n12846), .A2(n12340), .ZN(n12236) );
  OAI211_X1 U14888 ( .C1(n12839), .C2(n12344), .A(n12237), .B(n12236), .ZN(
        n12238) );
  AOI21_X1 U14889 ( .B1(n12944), .B2(n12347), .A(n12238), .ZN(n12239) );
  OAI21_X1 U14890 ( .B1(n12240), .B2(n12349), .A(n12239), .ZN(P3_U3156) );
  AOI21_X1 U14891 ( .B1(n12242), .B2(n12241), .A(n12349), .ZN(n12244) );
  NAND2_X1 U14892 ( .A1(n12244), .A2(n12243), .ZN(n12248) );
  NAND2_X1 U14893 ( .A1(n12903), .A2(n12341), .ZN(n12245) );
  NAND2_X1 U14894 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12742)
         );
  OAI211_X1 U14895 ( .C1(n12485), .C2(n12344), .A(n12245), .B(n12742), .ZN(
        n12246) );
  AOI21_X1 U14896 ( .B1(n12884), .B2(n12340), .A(n12246), .ZN(n12247) );
  OAI211_X1 U14897 ( .C1(n12285), .C2(n12249), .A(n12248), .B(n12247), .ZN(
        P3_U3159) );
  AOI22_X1 U14898 ( .A1(n12252), .A2(n12251), .B1(n12345), .B2(n12250), .ZN(
        n12254) );
  XNOR2_X1 U14899 ( .A(n6818), .B(n6446), .ZN(n12253) );
  XNOR2_X1 U14900 ( .A(n12254), .B(n12253), .ZN(n12259) );
  OAI22_X1 U14901 ( .A1(n12385), .A2(n12838), .B1(n12345), .B2(n12836), .ZN(
        n12774) );
  INV_X1 U14902 ( .A(n12774), .ZN(n12256) );
  AOI22_X1 U14903 ( .A1(n12771), .A2(n12340), .B1(P3_REG3_REG_28__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12255) );
  OAI21_X1 U14904 ( .B1(n12256), .B2(n12313), .A(n12255), .ZN(n12257) );
  AOI21_X1 U14905 ( .B1(n13001), .B2(n12347), .A(n12257), .ZN(n12258) );
  OAI21_X1 U14906 ( .B1(n12259), .B2(n12349), .A(n12258), .ZN(P3_U3160) );
  AOI21_X1 U14907 ( .B1(n12261), .B2(n12260), .A(n6565), .ZN(n12266) );
  OAI22_X1 U14908 ( .A1(n12837), .A2(n12838), .B1(n12485), .B2(n12836), .ZN(
        n12866) );
  INV_X1 U14909 ( .A(n12866), .ZN(n12263) );
  AOI22_X1 U14910 ( .A1(n12863), .A2(n12340), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12262) );
  OAI21_X1 U14911 ( .B1(n12263), .B2(n12313), .A(n12262), .ZN(n12264) );
  AOI21_X1 U14912 ( .B1(n13032), .B2(n12347), .A(n12264), .ZN(n12265) );
  OAI21_X1 U14913 ( .B1(n12266), .B2(n12349), .A(n12265), .ZN(P3_U3163) );
  XOR2_X1 U14914 ( .A(n12268), .B(n12267), .Z(n12275) );
  OR2_X1 U14915 ( .A1(n12269), .A2(n12838), .ZN(n12271) );
  OR2_X1 U14916 ( .A1(n12839), .A2(n12836), .ZN(n12270) );
  AND2_X1 U14917 ( .A1(n12271), .A2(n12270), .ZN(n12810) );
  AOI22_X1 U14918 ( .A1(n12802), .A2(n12340), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12272) );
  OAI21_X1 U14919 ( .B1(n12810), .B2(n12313), .A(n12272), .ZN(n12273) );
  AOI21_X1 U14920 ( .B1(n12803), .B2(n12347), .A(n12273), .ZN(n12274) );
  OAI21_X1 U14921 ( .B1(n12275), .B2(n12349), .A(n12274), .ZN(P3_U3165) );
  AOI211_X1 U14922 ( .C1(n12278), .C2(n12277), .A(n12349), .B(n12276), .ZN(
        n12279) );
  INV_X1 U14923 ( .A(n12279), .ZN(n12284) );
  NAND2_X1 U14924 ( .A1(n12341), .A2(n12918), .ZN(n12280) );
  NAND2_X1 U14925 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12681)
         );
  OAI211_X1 U14926 ( .C1(n12344), .C2(n12281), .A(n12280), .B(n12681), .ZN(
        n12282) );
  AOI21_X1 U14927 ( .B1(n12911), .B2(n12340), .A(n12282), .ZN(n12283) );
  OAI211_X1 U14928 ( .C1(n12286), .C2(n12285), .A(n12284), .B(n12283), .ZN(
        P3_U3166) );
  XNOR2_X1 U14929 ( .A(n12288), .B(n12287), .ZN(n12296) );
  AND2_X1 U14930 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n12705) );
  AOI21_X1 U14931 ( .B1(n12903), .B2(n12289), .A(n12705), .ZN(n12291) );
  NAND2_X1 U14932 ( .A1(n12340), .A2(n12901), .ZN(n12290) );
  OAI211_X1 U14933 ( .C1(n12293), .C2(n12292), .A(n12291), .B(n12290), .ZN(
        n12294) );
  AOI21_X1 U14934 ( .B1(n13056), .B2(n12347), .A(n12294), .ZN(n12295) );
  OAI21_X1 U14935 ( .B1(n12296), .B2(n12349), .A(n12295), .ZN(P3_U3168) );
  XNOR2_X1 U14936 ( .A(n12300), .B(n12839), .ZN(n12301) );
  XNOR2_X1 U14937 ( .A(n12302), .B(n12301), .ZN(n12307) );
  AOI22_X1 U14938 ( .A1(n12826), .A2(n12340), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12304) );
  NAND2_X1 U14939 ( .A1(n12568), .A2(n12341), .ZN(n12303) );
  OAI211_X1 U14940 ( .C1(n12822), .C2(n12344), .A(n12304), .B(n12303), .ZN(
        n12305) );
  AOI21_X1 U14941 ( .B1(n13020), .B2(n12347), .A(n12305), .ZN(n12306) );
  OAI21_X1 U14942 ( .B1(n12307), .B2(n12349), .A(n12306), .ZN(P3_U3169) );
  OAI211_X1 U14943 ( .C1(n12311), .C2(n12310), .A(n12309), .B(n12308), .ZN(
        n12316) );
  AOI22_X1 U14944 ( .A1(n12570), .A2(n12981), .B1(n12982), .B2(n12895), .ZN(
        n12878) );
  AOI22_X1 U14945 ( .A1(n12874), .A2(n12340), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12312) );
  OAI21_X1 U14946 ( .B1(n12878), .B2(n12313), .A(n12312), .ZN(n12314) );
  AOI21_X1 U14947 ( .B1(n13038), .B2(n12347), .A(n12314), .ZN(n12315) );
  NAND2_X1 U14948 ( .A1(n12316), .A2(n12315), .ZN(P3_U3173) );
  XNOR2_X1 U14949 ( .A(n12317), .B(n12569), .ZN(n12318) );
  XNOR2_X1 U14950 ( .A(n12319), .B(n12318), .ZN(n12327) );
  OAI22_X1 U14951 ( .A1(n12821), .A2(n12838), .B1(n12320), .B2(n12836), .ZN(
        n12857) );
  INV_X1 U14952 ( .A(n12854), .ZN(n12322) );
  OAI22_X1 U14953 ( .A1(n12322), .A2(n12321), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n6920), .ZN(n12323) );
  AOI21_X1 U14954 ( .B1(n12857), .B2(n12324), .A(n12323), .ZN(n12326) );
  NAND2_X1 U14955 ( .A1(n13027), .A2(n12347), .ZN(n12325) );
  OAI211_X1 U14956 ( .C1(n12327), .C2(n12349), .A(n12326), .B(n12325), .ZN(
        P3_U3175) );
  XNOR2_X1 U14957 ( .A(n12329), .B(n12328), .ZN(n12330) );
  XNOR2_X1 U14958 ( .A(n12331), .B(n12330), .ZN(n12337) );
  NAND2_X1 U14959 ( .A1(n12341), .A2(n12916), .ZN(n12332) );
  NAND2_X1 U14960 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12722)
         );
  OAI211_X1 U14961 ( .C1(n12333), .C2(n12344), .A(n12332), .B(n12722), .ZN(
        n12334) );
  AOI21_X1 U14962 ( .B1(n12892), .B2(n12340), .A(n12334), .ZN(n12336) );
  NAND2_X1 U14963 ( .A1(n13050), .A2(n12347), .ZN(n12335) );
  OAI211_X1 U14964 ( .C1(n12337), .C2(n12349), .A(n12336), .B(n12335), .ZN(
        P3_U3178) );
  XOR2_X1 U14965 ( .A(n12339), .B(n12338), .Z(n12350) );
  AOI22_X1 U14966 ( .A1(n12792), .A2(n12340), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12343) );
  NAND2_X1 U14967 ( .A1(n12796), .A2(n12341), .ZN(n12342) );
  OAI211_X1 U14968 ( .C1(n12345), .C2(n12344), .A(n12343), .B(n12342), .ZN(
        n12346) );
  AOI21_X1 U14969 ( .B1(n13008), .B2(n12347), .A(n12346), .ZN(n12348) );
  OAI21_X1 U14970 ( .B1(n12350), .B2(n12349), .A(n12348), .ZN(P3_U3180) );
  INV_X1 U14971 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n14097) );
  AND2_X1 U14972 ( .A1(n14097), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12353) );
  OAI22_X1 U14973 ( .A1(n12354), .A2(n12353), .B1(P2_DATAO_REG_30__SCAN_IN), 
        .B2(n14097), .ZN(n12357) );
  INV_X1 U14974 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n12355) );
  XNOR2_X1 U14975 ( .A(n12355), .B(P2_DATAO_REG_31__SCAN_IN), .ZN(n12356) );
  XNOR2_X1 U14976 ( .A(n12357), .B(n12356), .ZN(n13073) );
  NAND2_X1 U14977 ( .A1(n13073), .A2(n9956), .ZN(n12359) );
  NAND2_X1 U14978 ( .A1(n12368), .A2(SI_31_), .ZN(n12358) );
  INV_X1 U14979 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n12995) );
  NAND2_X1 U14980 ( .A1(n12360), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12362) );
  NAND2_X1 U14981 ( .A1(n10012), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12361) );
  OAI211_X1 U14982 ( .C1(n12995), .C2(n12363), .A(n12362), .B(n12361), .ZN(
        n12364) );
  INV_X1 U14983 ( .A(n12364), .ZN(n12365) );
  OR2_X1 U14984 ( .A1(n12375), .A2(n12755), .ZN(n12372) );
  NAND2_X1 U14985 ( .A1(n12367), .A2(n9956), .ZN(n12370) );
  NAND2_X1 U14986 ( .A1(n12368), .A2(SI_30_), .ZN(n12369) );
  NAND2_X1 U14987 ( .A1(n12925), .A2(n12374), .ZN(n12371) );
  AOI211_X1 U14988 ( .C1(n12755), .C2(n12925), .A(n12548), .B(n12377), .ZN(
        n12373) );
  OR2_X1 U14989 ( .A1(n12925), .A2(n12374), .ZN(n12546) );
  INV_X1 U14990 ( .A(n12546), .ZN(n12516) );
  NOR3_X1 U14991 ( .A1(n12516), .A2(n12755), .A3(n12743), .ZN(n12382) );
  INV_X1 U14992 ( .A(n12755), .ZN(n12563) );
  AOI211_X1 U14993 ( .C1(n12563), .C2(n12546), .A(n12548), .B(n12924), .ZN(
        n12376) );
  AOI21_X1 U14994 ( .B1(n12382), .B2(n12377), .A(n12376), .ZN(n12380) );
  OAI211_X1 U14995 ( .C1(n12377), .C2(n12925), .A(n12924), .B(n12548), .ZN(
        n12379) );
  NAND2_X1 U14996 ( .A1(n12381), .A2(n7967), .ZN(n12553) );
  AOI21_X1 U14997 ( .B1(n12924), .B2(n12548), .A(n12382), .ZN(n12383) );
  AOI21_X1 U14998 ( .B1(n12384), .B2(n12547), .A(n12383), .ZN(n12552) );
  AOI21_X1 U14999 ( .B1(n6502), .B2(n12515), .A(n12385), .ZN(n12388) );
  NAND3_X1 U15000 ( .A1(n12515), .A2(n12385), .A3(n6502), .ZN(n12386) );
  OAI21_X1 U15001 ( .B1(n12388), .B2(n12387), .A(n12386), .ZN(n12518) );
  MUX2_X1 U15002 ( .A(n6467), .B(n12389), .S(n12513), .Z(n12495) );
  INV_X1 U15003 ( .A(n12477), .ZN(n12393) );
  AND2_X1 U15004 ( .A1(n12390), .A2(n12512), .ZN(n12391) );
  OAI211_X1 U15005 ( .C1(n12393), .C2(n12392), .A(n12482), .B(n12391), .ZN(
        n12479) );
  INV_X1 U15006 ( .A(n12394), .ZN(n12476) );
  NAND2_X1 U15007 ( .A1(n12395), .A2(n12513), .ZN(n12398) );
  NAND3_X1 U15008 ( .A1(n12402), .A2(n12396), .A3(n12560), .ZN(n12397) );
  NOR2_X1 U15009 ( .A1(n12402), .A2(n12512), .ZN(n12403) );
  NOR2_X1 U15010 ( .A1(n12403), .A2(n12979), .ZN(n12406) );
  AOI21_X1 U15011 ( .B1(n12413), .B2(n12404), .A(n12513), .ZN(n12405) );
  NAND2_X1 U15012 ( .A1(n12408), .A2(n12407), .ZN(n12409) );
  NAND2_X1 U15013 ( .A1(n12409), .A2(n12513), .ZN(n12410) );
  OAI21_X1 U15014 ( .B1(n12412), .B2(n12411), .A(n12410), .ZN(n12417) );
  NOR2_X1 U15015 ( .A1(n12413), .A2(n12512), .ZN(n12415) );
  NOR2_X1 U15016 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  NAND2_X1 U15017 ( .A1(n12417), .A2(n12416), .ZN(n12423) );
  NAND3_X1 U15018 ( .A1(n12423), .A2(n12526), .A3(n12418), .ZN(n12420) );
  NAND3_X1 U15019 ( .A1(n12420), .A2(n12427), .A3(n12419), .ZN(n12421) );
  NAND2_X1 U15020 ( .A1(n12421), .A2(n12425), .ZN(n12430) );
  NAND3_X1 U15021 ( .A1(n12423), .A2(n12526), .A3(n12422), .ZN(n12426) );
  NAND3_X1 U15022 ( .A1(n12426), .A2(n12425), .A3(n12424), .ZN(n12428) );
  NAND2_X1 U15023 ( .A1(n12428), .A2(n12427), .ZN(n12429) );
  MUX2_X1 U15024 ( .A(n12432), .B(n12431), .S(n12513), .Z(n12433) );
  OR2_X1 U15025 ( .A1(n12435), .A2(n12434), .ZN(n12437) );
  MUX2_X1 U15026 ( .A(n12437), .B(n12436), .S(n12513), .Z(n12438) );
  MUX2_X1 U15027 ( .A(n12439), .B(n6461), .S(n12513), .Z(n12440) );
  NAND2_X1 U15028 ( .A1(n12441), .A2(n7081), .ZN(n12453) );
  INV_X1 U15029 ( .A(n12442), .ZN(n12445) );
  INV_X1 U15030 ( .A(n12443), .ZN(n12444) );
  MUX2_X1 U15031 ( .A(n12445), .B(n12444), .S(n12512), .Z(n12446) );
  NOR2_X1 U15032 ( .A1(n12533), .A2(n12446), .ZN(n12452) );
  NAND2_X1 U15033 ( .A1(n12455), .A2(n12447), .ZN(n12450) );
  NAND2_X1 U15034 ( .A1(n12454), .A2(n12448), .ZN(n12449) );
  MUX2_X1 U15035 ( .A(n12450), .B(n12449), .S(n12513), .Z(n12451) );
  AOI21_X1 U15036 ( .B1(n12453), .B2(n12452), .A(n12451), .ZN(n12460) );
  MUX2_X1 U15037 ( .A(n12455), .B(n12454), .S(n12512), .Z(n12456) );
  NAND2_X1 U15038 ( .A1(n12536), .A2(n12456), .ZN(n12459) );
  MUX2_X1 U15039 ( .A(n12457), .B(n6509), .S(n12513), .Z(n12458) );
  OAI21_X1 U15040 ( .B1(n12460), .B2(n12459), .A(n12458), .ZN(n12461) );
  MUX2_X1 U15041 ( .A(n12463), .B(n12462), .S(n12512), .Z(n12464) );
  INV_X1 U15042 ( .A(n12465), .ZN(n12467) );
  NAND2_X1 U15043 ( .A1(n12467), .A2(n12466), .ZN(n12468) );
  NAND2_X1 U15044 ( .A1(n12468), .A2(n12513), .ZN(n12469) );
  INV_X1 U15045 ( .A(n12470), .ZN(n12472) );
  NAND2_X1 U15046 ( .A1(n12905), .A2(n12512), .ZN(n12473) );
  AOI22_X1 U15047 ( .A1(n12479), .A2(n12476), .B1(n7062), .B2(n12475), .ZN(
        n12481) );
  NAND3_X1 U15048 ( .A1(n6528), .A2(n12477), .A3(n12513), .ZN(n12478) );
  NAND2_X1 U15049 ( .A1(n12479), .A2(n12478), .ZN(n12480) );
  OAI21_X1 U15050 ( .B1(n12481), .B2(n12893), .A(n12480), .ZN(n12484) );
  MUX2_X1 U15051 ( .A(n12482), .B(n6528), .S(n12512), .Z(n12483) );
  NAND3_X1 U15052 ( .A1(n12484), .A2(n12872), .A3(n12483), .ZN(n12489) );
  XNOR2_X1 U15053 ( .A(n13032), .B(n12570), .ZN(n12864) );
  NAND2_X1 U15054 ( .A1(n13038), .A2(n12485), .ZN(n12486) );
  MUX2_X1 U15055 ( .A(n12487), .B(n12486), .S(n12513), .Z(n12488) );
  MUX2_X1 U15056 ( .A(n12491), .B(n12490), .S(n12513), .Z(n12492) );
  NAND3_X1 U15057 ( .A1(n12852), .A2(n12493), .A3(n12492), .ZN(n12494) );
  NAND3_X1 U15058 ( .A1(n12944), .A2(n12821), .A3(n12512), .ZN(n12496) );
  NAND2_X1 U15059 ( .A1(n12498), .A2(n12497), .ZN(n12499) );
  NAND2_X1 U15060 ( .A1(n12501), .A2(n12499), .ZN(n12500) );
  MUX2_X1 U15061 ( .A(n12501), .B(n12500), .S(n12513), .Z(n12502) );
  INV_X1 U15062 ( .A(n12506), .ZN(n12504) );
  NAND2_X1 U15063 ( .A1(n12504), .A2(n12509), .ZN(n12523) );
  NOR2_X1 U15064 ( .A1(n12523), .A2(n12505), .ZN(n12507) );
  NOR2_X1 U15065 ( .A1(n12523), .A2(n6709), .ZN(n12510) );
  NOR2_X1 U15066 ( .A1(n12769), .A2(n12513), .ZN(n12520) );
  INV_X1 U15067 ( .A(n12523), .ZN(n12793) );
  INV_X1 U15068 ( .A(n12914), .ZN(n12909) );
  NAND4_X1 U15069 ( .A1(n10074), .A2(n7416), .A3(n12526), .A4(n12525), .ZN(
        n12528) );
  NOR4_X1 U15070 ( .A1(n12529), .A2(n10589), .A3(n12528), .A4(n12527), .ZN(
        n12531) );
  NAND2_X1 U15071 ( .A1(n12541), .A2(n12540), .ZN(n12885) );
  INV_X1 U15072 ( .A(n12852), .ZN(n12855) );
  NOR4_X1 U15073 ( .A1(n12801), .A2(n7181), .A3(n12542), .A4(n12855), .ZN(
        n12543) );
  NAND2_X1 U15074 ( .A1(n12550), .A2(n12549), .ZN(n12551) );
  NAND2_X1 U15075 ( .A1(n12555), .A2(n12554), .ZN(n12562) );
  NAND3_X1 U15076 ( .A1(n12557), .A2(n12556), .A3(n12982), .ZN(n12558) );
  OAI211_X1 U15077 ( .C1(n12560), .C2(n12559), .A(n12558), .B(P3_B_REG_SCAN_IN), .ZN(n12561) );
  NAND2_X1 U15078 ( .A1(n12562), .A2(n12561), .ZN(P3_U3296) );
  MUX2_X1 U15079 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n12563), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U15080 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12564), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U15081 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12565), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U15082 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12566), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U15083 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12796), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U15084 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12567), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U15085 ( .A(n12568), .B(P3_DATAO_REG_23__SCAN_IN), .S(n12571), .Z(
        P3_U3514) );
  MUX2_X1 U15086 ( .A(n12569), .B(P3_DATAO_REG_22__SCAN_IN), .S(n12571), .Z(
        P3_U3513) );
  MUX2_X1 U15087 ( .A(n12570), .B(P3_DATAO_REG_21__SCAN_IN), .S(n12571), .Z(
        P3_U3512) );
  MUX2_X1 U15088 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12887), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15089 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12895), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U15090 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12903), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U15091 ( .A(n12905), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12571), .Z(
        P3_U3507) );
  MUX2_X1 U15092 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12918), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U15093 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12572), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U15094 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12573), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U15095 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12574), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15096 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12575), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U15097 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12576), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15098 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12577), .S(P3_U3897), .Z(
        P3_U3500) );
  MUX2_X1 U15099 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12578), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U15100 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12579), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U15101 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12580), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15102 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12581), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U15103 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12582), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U15104 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12980), .S(P3_U3897), .Z(
        P3_U3494) );
  MUX2_X1 U15105 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12583), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15106 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n9514), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15107 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n12584), .S(P3_U3897), .Z(
        P3_U3491) );
  XNOR2_X1 U15108 ( .A(n12612), .B(P3_REG2_REG_12__SCAN_IN), .ZN(n12587) );
  AND3_X1 U15109 ( .A1(n12588), .A2(n12587), .A3(n12586), .ZN(n12589) );
  OAI21_X1 U15110 ( .B1(n6641), .B2(n12589), .A(n15586), .ZN(n12608) );
  INV_X1 U15111 ( .A(n12612), .ZN(n12617) );
  INV_X1 U15112 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n12591) );
  NAND2_X1 U15113 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n12590)
         );
  OAI21_X1 U15114 ( .B1(n15605), .B2(n12591), .A(n12590), .ZN(n12592) );
  AOI21_X1 U15115 ( .B1(n15598), .B2(n12617), .A(n12592), .ZN(n12607) );
  INV_X1 U15116 ( .A(n12593), .ZN(n12595) );
  XNOR2_X1 U15117 ( .A(n12612), .B(n12596), .ZN(n12609) );
  XNOR2_X1 U15118 ( .A(n12610), .B(n12609), .ZN(n12597) );
  NAND2_X1 U15119 ( .A1(n12597), .A2(n15591), .ZN(n12606) );
  INV_X1 U15120 ( .A(n12598), .ZN(n12599) );
  AOI22_X1 U15121 ( .A1(n12602), .A2(n12601), .B1(n12600), .B2(n12599), .ZN(
        n12604) );
  MUX2_X1 U15122 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n7168), .Z(n12614) );
  XOR2_X1 U15123 ( .A(n12612), .B(n12614), .Z(n12603) );
  OAI211_X1 U15124 ( .C1(n12604), .C2(n12603), .A(n12615), .B(n15595), .ZN(
        n12605) );
  NAND4_X1 U15125 ( .A1(n12608), .A2(n12607), .A3(n12606), .A4(n12605), .ZN(
        P3_U3194) );
  NAND2_X1 U15126 ( .A1(n12612), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12611) );
  INV_X1 U15127 ( .A(n12637), .ZN(n12646) );
  XOR2_X1 U15128 ( .A(P3_REG1_REG_13__SCAN_IN), .B(n12636), .Z(n12627) );
  OAI21_X1 U15129 ( .B1(P3_REG2_REG_13__SCAN_IN), .B2(n12613), .A(n12632), 
        .ZN(n12625) );
  MUX2_X1 U15130 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n7168), .Z(n12644) );
  XNOR2_X1 U15131 ( .A(n12637), .B(n12644), .ZN(n12619) );
  INV_X1 U15132 ( .A(n12614), .ZN(n12616) );
  AOI21_X1 U15133 ( .B1(n12619), .B2(n12618), .A(n6629), .ZN(n12620) );
  NOR2_X1 U15134 ( .A1(n12620), .A2(n15576), .ZN(n12624) );
  NAND2_X1 U15135 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(P3_U3151), .ZN(n12622)
         );
  NAND2_X1 U15136 ( .A1(n15539), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n12621) );
  OAI211_X1 U15137 ( .C1(n15549), .C2(n12637), .A(n12622), .B(n12621), .ZN(
        n12623) );
  AOI211_X1 U15138 ( .C1(n12625), .C2(n15586), .A(n12624), .B(n12623), .ZN(
        n12626) );
  OAI21_X1 U15139 ( .B1(n12627), .B2(n12730), .A(n12626), .ZN(P3_U3195) );
  INV_X1 U15140 ( .A(n12632), .ZN(n12629) );
  NAND2_X1 U15141 ( .A1(n12641), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12657) );
  OR2_X1 U15142 ( .A1(n12641), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12628) );
  NOR3_X1 U15143 ( .A1(n12629), .A2(n6623), .A3(n12630), .ZN(n12633) );
  INV_X1 U15144 ( .A(n12630), .ZN(n12631) );
  OAI21_X1 U15145 ( .B1(n12633), .B2(n6642), .A(n15586), .ZN(n12652) );
  NOR2_X1 U15146 ( .A1(n15549), .A2(n12641), .ZN(n12634) );
  AOI211_X1 U15147 ( .C1(n15539), .C2(P3_ADDR_REG_14__SCAN_IN), .A(n12635), 
        .B(n12634), .ZN(n12651) );
  NAND2_X1 U15148 ( .A1(n12636), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n12640) );
  NAND2_X1 U15149 ( .A1(n12638), .A2(n12637), .ZN(n12639) );
  NAND2_X1 U15150 ( .A1(n12641), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12658) );
  OR2_X1 U15151 ( .A1(n12641), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12642) );
  AND2_X1 U15152 ( .A1(n12658), .A2(n12642), .ZN(n12653) );
  XNOR2_X1 U15153 ( .A(n12654), .B(n12653), .ZN(n12643) );
  NAND2_X1 U15154 ( .A1(n12643), .A2(n15591), .ZN(n12650) );
  INV_X1 U15155 ( .A(n12644), .ZN(n12645) );
  MUX2_X1 U15156 ( .A(n12653), .B(n6623), .S(n12737), .Z(n12647) );
  OAI211_X1 U15157 ( .C1(n12648), .C2(n12647), .A(n12660), .B(n15595), .ZN(
        n12649) );
  NAND4_X1 U15158 ( .A1(n12652), .A2(n12651), .A3(n12650), .A4(n12649), .ZN(
        P3_U3196) );
  INV_X1 U15159 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12974) );
  XNOR2_X1 U15160 ( .A(n12672), .B(n12974), .ZN(n12671) );
  NOR2_X1 U15161 ( .A1(n12655), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n12656) );
  OAI21_X1 U15162 ( .B1(n12656), .B2(n12678), .A(n15586), .ZN(n12670) );
  MUX2_X1 U15163 ( .A(n12658), .B(n12657), .S(n12737), .Z(n12659) );
  INV_X1 U15164 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12662) );
  MUX2_X1 U15165 ( .A(n12662), .B(n12974), .S(n7168), .Z(n12663) );
  NAND2_X1 U15166 ( .A1(n12664), .A2(n12663), .ZN(n12682) );
  OAI21_X1 U15167 ( .B1(n12664), .B2(n12663), .A(n12682), .ZN(n12668) );
  NAND2_X1 U15168 ( .A1(n15539), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n12665) );
  OAI211_X1 U15169 ( .C1(n15549), .C2(n12683), .A(n12666), .B(n12665), .ZN(
        n12667) );
  AOI21_X1 U15170 ( .B1(n12668), .B2(n15595), .A(n12667), .ZN(n12669) );
  OAI211_X1 U15171 ( .C1(n12671), .C2(n12730), .A(n12670), .B(n12669), .ZN(
        P3_U3197) );
  INV_X1 U15172 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12967) );
  XNOR2_X1 U15173 ( .A(n12701), .B(n12967), .ZN(n12692) );
  NAND2_X1 U15174 ( .A1(n12672), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U15175 ( .A1(n12673), .A2(n12683), .ZN(n12674) );
  XOR2_X1 U15176 ( .A(n12692), .B(n12693), .Z(n12691) );
  INV_X1 U15177 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12919) );
  XNOR2_X1 U15178 ( .A(n12701), .B(n12919), .ZN(n12676) );
  INV_X1 U15179 ( .A(n12694), .ZN(n12680) );
  NOR3_X1 U15180 ( .A1(n12678), .A2(n12677), .A3(n12676), .ZN(n12679) );
  OAI21_X1 U15181 ( .B1(n12680), .B2(n12679), .A(n15586), .ZN(n12690) );
  INV_X1 U15182 ( .A(n12701), .ZN(n12695) );
  OAI21_X1 U15183 ( .B1(n15605), .B2(n15734), .A(n12681), .ZN(n12688) );
  MUX2_X1 U15184 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n7168), .Z(n12702) );
  XNOR2_X1 U15185 ( .A(n12701), .B(n12702), .ZN(n12686) );
  OAI21_X1 U15186 ( .B1(n12684), .B2(n12683), .A(n12682), .ZN(n12685) );
  AOI211_X1 U15187 ( .C1(n12686), .C2(n12685), .A(n15576), .B(n12700), .ZN(
        n12687) );
  AOI211_X1 U15188 ( .C1(n15598), .C2(n12695), .A(n12688), .B(n12687), .ZN(
        n12689) );
  OAI211_X1 U15189 ( .C1(n12691), .C2(n12730), .A(n12690), .B(n12689), .ZN(
        P3_U3198) );
  XNOR2_X1 U15190 ( .A(n12714), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n12711) );
  NAND2_X1 U15191 ( .A1(n12696), .A2(n12724), .ZN(n12715) );
  OAI21_X1 U15192 ( .B1(n12696), .B2(n12724), .A(n12715), .ZN(n12697) );
  INV_X1 U15193 ( .A(n12697), .ZN(n12699) );
  INV_X1 U15194 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12906) );
  NOR2_X1 U15195 ( .A1(n12697), .A2(n12906), .ZN(n12719) );
  INV_X1 U15196 ( .A(n12719), .ZN(n12698) );
  OAI21_X1 U15197 ( .B1(P3_REG2_REG_17__SCAN_IN), .B2(n12699), .A(n12698), 
        .ZN(n12709) );
  MUX2_X1 U15198 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n7168), .Z(n12725) );
  XOR2_X1 U15199 ( .A(n12725), .B(n12713), .Z(n12703) );
  AOI211_X1 U15200 ( .C1(n12704), .C2(n12703), .A(n15576), .B(n12723), .ZN(
        n12708) );
  AOI21_X1 U15201 ( .B1(n15539), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12705), 
        .ZN(n12706) );
  OAI21_X1 U15202 ( .B1(n15549), .B2(n12724), .A(n12706), .ZN(n12707) );
  AOI211_X1 U15203 ( .C1(n12709), .C2(n15586), .A(n12708), .B(n12707), .ZN(
        n12710) );
  OAI21_X1 U15204 ( .B1(n12711), .B2(n12730), .A(n12710), .ZN(P3_U3199) );
  XOR2_X1 U15205 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n12746), .Z(n12747) );
  XOR2_X1 U15206 ( .A(n12747), .B(n12748), .Z(n12731) );
  INV_X1 U15207 ( .A(n12715), .ZN(n12718) );
  NAND2_X1 U15208 ( .A1(n12746), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12732) );
  OR2_X1 U15209 ( .A1(n12746), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12716) );
  AND2_X1 U15210 ( .A1(n12732), .A2(n12716), .ZN(n12717) );
  OAI21_X1 U15211 ( .B1(n12719), .B2(n12718), .A(n12717), .ZN(n12733) );
  INV_X1 U15212 ( .A(n12733), .ZN(n12721) );
  NOR3_X1 U15213 ( .A1(n12719), .A2(n12718), .A3(n12717), .ZN(n12720) );
  OAI21_X1 U15214 ( .B1(n12721), .B2(n12720), .A(n15586), .ZN(n12729) );
  OAI21_X1 U15215 ( .B1(n15605), .B2(n8795), .A(n12722), .ZN(n12728) );
  MUX2_X1 U15216 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n7168), .Z(n12727) );
  NOR2_X1 U15217 ( .A1(n12726), .A2(n12727), .ZN(n12735) );
  NAND2_X1 U15218 ( .A1(n12733), .A2(n12732), .ZN(n12734) );
  XNOR2_X1 U15219 ( .A(n12743), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12738) );
  XNOR2_X1 U15220 ( .A(n12734), .B(n12738), .ZN(n12753) );
  AOI21_X1 U15221 ( .B1(n12736), .B2(n6986), .A(n12735), .ZN(n12740) );
  XNOR2_X1 U15222 ( .A(n12743), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12749) );
  MUX2_X1 U15223 ( .A(n12749), .B(n12738), .S(n12737), .Z(n12739) );
  XNOR2_X1 U15224 ( .A(n12740), .B(n12739), .ZN(n12745) );
  NAND2_X1 U15225 ( .A1(n15539), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n12741) );
  OAI211_X1 U15226 ( .C1(n15549), .C2(n12743), .A(n12742), .B(n12741), .ZN(
        n12744) );
  AOI21_X1 U15227 ( .B1(n12745), .B2(n15595), .A(n12744), .ZN(n12752) );
  NAND2_X1 U15228 ( .A1(n12750), .A2(n15591), .ZN(n12751) );
  NAND2_X1 U15229 ( .A1(n15618), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n12757) );
  NOR2_X1 U15230 ( .A1(n12756), .A2(n15610), .ZN(n12761) );
  OAI21_X1 U15231 ( .B1(n12993), .B2(n12761), .A(n15616), .ZN(n12758) );
  OAI211_X1 U15232 ( .C1(n12924), .C2(n12828), .A(n12757), .B(n12758), .ZN(
        P3_U3202) );
  INV_X1 U15233 ( .A(n12925), .ZN(n12998) );
  NAND2_X1 U15234 ( .A1(n15618), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n12759) );
  OAI211_X1 U15235 ( .C1(n12998), .C2(n12828), .A(n12759), .B(n12758), .ZN(
        P3_U3203) );
  AND2_X1 U15236 ( .A1(n15618), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n12760) );
  AOI211_X1 U15237 ( .C1(n12763), .C2(n12762), .A(n12761), .B(n12760), .ZN(
        n12766) );
  NAND2_X1 U15238 ( .A1(n12764), .A2(n15616), .ZN(n12765) );
  NAND2_X1 U15239 ( .A1(n12778), .A2(n12768), .ZN(n12770) );
  AOI22_X1 U15240 ( .A1(n13001), .A2(n12913), .B1(n12912), .B2(n12771), .ZN(
        n12777) );
  INV_X1 U15241 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12775) );
  OAI211_X1 U15242 ( .C1(n13004), .C2(n12922), .A(n12777), .B(n12776), .ZN(
        P3_U3205) );
  XNOR2_X1 U15243 ( .A(n12782), .B(n12781), .ZN(n12783) );
  INV_X1 U15244 ( .A(n12932), .ZN(n12787) );
  AOI22_X1 U15245 ( .A1(n12785), .A2(n12912), .B1(n15618), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12786) );
  OAI21_X1 U15246 ( .B1(n12787), .B2(n12828), .A(n12786), .ZN(n12788) );
  AOI21_X1 U15247 ( .B1(n12934), .B2(n12789), .A(n12788), .ZN(n12790) );
  OAI21_X1 U15248 ( .B1(n12935), .B2(n15618), .A(n12790), .ZN(P3_U3206) );
  XNOR2_X1 U15249 ( .A(n12791), .B(n12793), .ZN(n13011) );
  AOI22_X1 U15250 ( .A1(n13008), .A2(n12913), .B1(n12912), .B2(n12792), .ZN(
        n12799) );
  INV_X1 U15251 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n12797) );
  MUX2_X1 U15252 ( .A(n12797), .B(n13006), .S(n15616), .Z(n12798) );
  OAI211_X1 U15253 ( .C1(n13011), .C2(n12922), .A(n12799), .B(n12798), .ZN(
        P3_U3207) );
  XNOR2_X1 U15254 ( .A(n12800), .B(n12801), .ZN(n13013) );
  AOI22_X1 U15255 ( .A1(n12803), .A2(n12913), .B1(n12912), .B2(n12802), .ZN(
        n12814) );
  INV_X1 U15256 ( .A(n12804), .ZN(n12805) );
  NAND2_X1 U15257 ( .A1(n12841), .A2(n12805), .ZN(n12819) );
  NAND2_X1 U15258 ( .A1(n12819), .A2(n12820), .ZN(n12818) );
  NAND3_X1 U15259 ( .A1(n12818), .A2(n12807), .A3(n12806), .ZN(n12808) );
  NAND3_X1 U15260 ( .A1(n12809), .A2(n12986), .A3(n12808), .ZN(n12811) );
  NAND2_X1 U15261 ( .A1(n12811), .A2(n12810), .ZN(n13014) );
  MUX2_X1 U15262 ( .A(P3_REG2_REG_25__SCAN_IN), .B(n13014), .S(n15616), .Z(
        n12812) );
  INV_X1 U15263 ( .A(n12812), .ZN(n12813) );
  OAI211_X1 U15264 ( .C1(n13013), .C2(n12922), .A(n12814), .B(n12813), .ZN(
        P3_U3208) );
  INV_X1 U15265 ( .A(n12815), .ZN(n12816) );
  AOI21_X1 U15266 ( .B1(n12820), .B2(n12817), .A(n12816), .ZN(n13023) );
  INV_X1 U15267 ( .A(n13023), .ZN(n12831) );
  OAI211_X1 U15268 ( .C1(n12820), .C2(n12819), .A(n12818), .B(n12986), .ZN(
        n12825) );
  OAI22_X1 U15269 ( .A1(n12822), .A2(n12838), .B1(n12821), .B2(n12836), .ZN(
        n12823) );
  INV_X1 U15270 ( .A(n12823), .ZN(n12824) );
  NAND2_X1 U15271 ( .A1(n12825), .A2(n12824), .ZN(n13017) );
  MUX2_X1 U15272 ( .A(n13017), .B(P3_REG2_REG_24__SCAN_IN), .S(n15618), .Z(
        n12830) );
  INV_X1 U15273 ( .A(n12826), .ZN(n12827) );
  OAI22_X1 U15274 ( .A1(n12941), .A2(n12828), .B1(n12827), .B2(n15610), .ZN(
        n12829) );
  AOI211_X1 U15275 ( .C1(n12831), .C2(n12845), .A(n12830), .B(n12829), .ZN(
        n12832) );
  INV_X1 U15276 ( .A(n12832), .ZN(P3_U3209) );
  AOI21_X1 U15277 ( .B1(n12833), .B2(n12835), .A(n12834), .ZN(n12842) );
  OAI22_X1 U15278 ( .A1(n12839), .A2(n12838), .B1(n12837), .B2(n12836), .ZN(
        n12840) );
  AOI21_X1 U15279 ( .B1(n12842), .B2(n12841), .A(n12840), .ZN(n12947) );
  NAND2_X1 U15280 ( .A1(n12844), .A2(n12843), .ZN(n12945) );
  NAND3_X1 U15281 ( .A1(n12946), .A2(n12945), .A3(n12845), .ZN(n12851) );
  INV_X1 U15282 ( .A(n12846), .ZN(n12848) );
  INV_X1 U15283 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n12847) );
  OAI22_X1 U15284 ( .A1(n12848), .A2(n15610), .B1(n15616), .B2(n12847), .ZN(
        n12849) );
  AOI21_X1 U15285 ( .B1(n12944), .B2(n12913), .A(n12849), .ZN(n12850) );
  OAI211_X1 U15286 ( .C1(n15618), .C2(n12947), .A(n12851), .B(n12850), .ZN(
        P3_U3210) );
  XNOR2_X1 U15287 ( .A(n12853), .B(n12852), .ZN(n13030) );
  AOI22_X1 U15288 ( .A1(n13027), .A2(n12913), .B1(n12912), .B2(n12854), .ZN(
        n12861) );
  INV_X1 U15289 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n12859) );
  XNOR2_X1 U15290 ( .A(n12856), .B(n12855), .ZN(n12858) );
  AOI21_X1 U15291 ( .B1(n12858), .B2(n12986), .A(n12857), .ZN(n13025) );
  MUX2_X1 U15292 ( .A(n12859), .B(n13025), .S(n15616), .Z(n12860) );
  OAI211_X1 U15293 ( .C1(n13030), .C2(n12922), .A(n12861), .B(n12860), .ZN(
        P3_U3211) );
  XNOR2_X1 U15294 ( .A(n12862), .B(n12864), .ZN(n13035) );
  AOI22_X1 U15295 ( .A1(n13032), .A2(n12913), .B1(n12912), .B2(n12863), .ZN(
        n12870) );
  INV_X1 U15296 ( .A(P3_REG2_REG_21__SCAN_IN), .ZN(n12868) );
  XNOR2_X1 U15297 ( .A(n12865), .B(n12864), .ZN(n12867) );
  AOI21_X1 U15298 ( .B1(n12867), .B2(n12986), .A(n12866), .ZN(n13031) );
  MUX2_X1 U15299 ( .A(n12868), .B(n13031), .S(n15616), .Z(n12869) );
  OAI211_X1 U15300 ( .C1(n13035), .C2(n12922), .A(n12870), .B(n12869), .ZN(
        P3_U3212) );
  OAI21_X1 U15301 ( .B1(n12873), .B2(n12872), .A(n12871), .ZN(n13041) );
  AOI22_X1 U15302 ( .A1(n13038), .A2(n12913), .B1(n12912), .B2(n12874), .ZN(
        n12882) );
  OAI211_X1 U15303 ( .C1(n12877), .C2(n12876), .A(n12875), .B(n12986), .ZN(
        n12879) );
  INV_X1 U15304 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12880) );
  MUX2_X1 U15305 ( .A(n13037), .B(n12880), .S(n15618), .Z(n12881) );
  OAI211_X1 U15306 ( .C1(n13041), .C2(n12922), .A(n12882), .B(n12881), .ZN(
        P3_U3213) );
  XOR2_X1 U15307 ( .A(n12883), .B(n12885), .Z(n13047) );
  AOI22_X1 U15308 ( .A1(n13044), .A2(n12913), .B1(n12912), .B2(n12884), .ZN(
        n12890) );
  XOR2_X1 U15309 ( .A(n12886), .B(n12885), .Z(n12888) );
  AOI222_X1 U15310 ( .A1(n12903), .A2(n12982), .B1(n12986), .B2(n12888), .C1(
        n12887), .C2(n12981), .ZN(n13042) );
  MUX2_X1 U15311 ( .A(n15693), .B(n13042), .S(n15616), .Z(n12889) );
  OAI211_X1 U15312 ( .C1(n13047), .C2(n12922), .A(n12890), .B(n12889), .ZN(
        P3_U3214) );
  OAI21_X1 U15313 ( .B1(n6627), .B2(n6701), .A(n12891), .ZN(n13053) );
  AOI22_X1 U15314 ( .A1(n13050), .A2(n12913), .B1(n12912), .B2(n12892), .ZN(
        n12899) );
  INV_X1 U15315 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12897) );
  OAI21_X1 U15316 ( .B1(n12894), .B2(n12893), .A(n7952), .ZN(n12896) );
  AOI222_X1 U15317 ( .A1(n12896), .A2(n12986), .B1(n12895), .B2(n12981), .C1(
        n12916), .C2(n12982), .ZN(n13048) );
  MUX2_X1 U15318 ( .A(n12897), .B(n13048), .S(n15616), .Z(n12898) );
  OAI211_X1 U15319 ( .C1(n13053), .C2(n12922), .A(n12899), .B(n12898), .ZN(
        P3_U3215) );
  XNOR2_X1 U15320 ( .A(n12900), .B(n7062), .ZN(n13059) );
  AOI22_X1 U15321 ( .A1(n13056), .A2(n12913), .B1(n12912), .B2(n12901), .ZN(
        n12908) );
  XNOR2_X1 U15322 ( .A(n12902), .B(n7062), .ZN(n12904) );
  AOI222_X1 U15323 ( .A1(n12905), .A2(n12982), .B1(n12986), .B2(n12904), .C1(
        n12903), .C2(n12981), .ZN(n13054) );
  MUX2_X1 U15324 ( .A(n12906), .B(n13054), .S(n15616), .Z(n12907) );
  OAI211_X1 U15325 ( .C1(n13059), .C2(n12922), .A(n12908), .B(n12907), .ZN(
        P3_U3216) );
  XNOR2_X1 U15326 ( .A(n12910), .B(n12909), .ZN(n13066) );
  AOI22_X1 U15327 ( .A1(n13062), .A2(n12913), .B1(n12912), .B2(n12911), .ZN(
        n12921) );
  XNOR2_X1 U15328 ( .A(n12915), .B(n12914), .ZN(n12917) );
  AOI222_X1 U15329 ( .A1(n12918), .A2(n12982), .B1(n12986), .B2(n12917), .C1(
        n12916), .C2(n12981), .ZN(n13060) );
  MUX2_X1 U15330 ( .A(n12919), .B(n13060), .S(n15616), .Z(n12920) );
  OAI211_X1 U15331 ( .C1(n13066), .C2(n12922), .A(n12921), .B(n12920), .ZN(
        P3_U3217) );
  NAND2_X1 U15332 ( .A1(n12993), .A2(n15665), .ZN(n12926) );
  NAND2_X1 U15333 ( .A1(n15663), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n12923) );
  OAI211_X1 U15334 ( .C1(n12924), .C2(n12976), .A(n12926), .B(n12923), .ZN(
        P3_U3490) );
  NAND2_X1 U15335 ( .A1(n12925), .A2(n12968), .ZN(n12927) );
  OAI211_X1 U15336 ( .C1(n15665), .C2(n12928), .A(n12927), .B(n12926), .ZN(
        P3_U3489) );
  INV_X1 U15337 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n12929) );
  MUX2_X1 U15338 ( .A(n12929), .B(n12999), .S(n15665), .Z(n12931) );
  NAND2_X1 U15339 ( .A1(n13001), .A2(n12968), .ZN(n12930) );
  OAI211_X1 U15340 ( .C1(n13004), .C2(n12971), .A(n12931), .B(n12930), .ZN(
        P3_U3487) );
  INV_X1 U15341 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12936) );
  MUX2_X1 U15342 ( .A(n12936), .B(n13006), .S(n15665), .Z(n12938) );
  NAND2_X1 U15343 ( .A1(n13008), .A2(n12968), .ZN(n12937) );
  OAI211_X1 U15344 ( .C1(n13011), .C2(n12971), .A(n12938), .B(n12937), .ZN(
        P3_U3485) );
  OAI22_X1 U15345 ( .A1(n13013), .A2(n12971), .B1(n13012), .B2(n12976), .ZN(
        n12940) );
  MUX2_X1 U15346 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n13014), .S(n15665), .Z(
        n12939) );
  OR2_X1 U15347 ( .A1(n12940), .A2(n12939), .ZN(P3_U3484) );
  OAI22_X1 U15348 ( .A1(n13023), .A2(n12971), .B1(n12941), .B2(n12976), .ZN(
        n12943) );
  MUX2_X1 U15349 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n13017), .S(n15665), .Z(
        n12942) );
  OR2_X1 U15350 ( .A1(n12943), .A2(n12942), .ZN(P3_U3483) );
  INV_X1 U15351 ( .A(n12944), .ZN(n12949) );
  NAND3_X1 U15352 ( .A1(n12946), .A2(n12945), .A3(n15630), .ZN(n12948) );
  OAI211_X1 U15353 ( .C1(n12949), .C2(n15626), .A(n12948), .B(n12947), .ZN(
        n13024) );
  MUX2_X1 U15354 ( .A(P3_REG1_REG_23__SCAN_IN), .B(n13024), .S(n15665), .Z(
        P3_U3482) );
  INV_X1 U15355 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12950) );
  MUX2_X1 U15356 ( .A(n12950), .B(n13025), .S(n15665), .Z(n12952) );
  NAND2_X1 U15357 ( .A1(n13027), .A2(n12968), .ZN(n12951) );
  OAI211_X1 U15358 ( .C1(n13030), .C2(n12971), .A(n12952), .B(n12951), .ZN(
        P3_U3481) );
  INV_X1 U15359 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12953) );
  MUX2_X1 U15360 ( .A(n12953), .B(n13031), .S(n15665), .Z(n12955) );
  NAND2_X1 U15361 ( .A1(n13032), .A2(n12968), .ZN(n12954) );
  OAI211_X1 U15362 ( .C1(n13035), .C2(n12971), .A(n12955), .B(n12954), .ZN(
        P3_U3480) );
  INV_X1 U15363 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12956) );
  MUX2_X1 U15364 ( .A(n13037), .B(n12956), .S(n15663), .Z(n12958) );
  NAND2_X1 U15365 ( .A1(n13038), .A2(n12968), .ZN(n12957) );
  OAI211_X1 U15366 ( .C1(n13041), .C2(n12971), .A(n12958), .B(n12957), .ZN(
        P3_U3479) );
  INV_X1 U15367 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12959) );
  MUX2_X1 U15368 ( .A(n12959), .B(n13042), .S(n15665), .Z(n12961) );
  NAND2_X1 U15369 ( .A1(n13044), .A2(n12968), .ZN(n12960) );
  OAI211_X1 U15370 ( .C1(n13047), .C2(n12971), .A(n12961), .B(n12960), .ZN(
        P3_U3478) );
  INV_X1 U15371 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12962) );
  MUX2_X1 U15372 ( .A(n12962), .B(n13048), .S(n15665), .Z(n12964) );
  NAND2_X1 U15373 ( .A1(n13050), .A2(n12968), .ZN(n12963) );
  OAI211_X1 U15374 ( .C1(n13053), .C2(n12971), .A(n12964), .B(n12963), .ZN(
        P3_U3477) );
  MUX2_X1 U15375 ( .A(n15723), .B(n13054), .S(n15665), .Z(n12966) );
  NAND2_X1 U15376 ( .A1(n13056), .A2(n12968), .ZN(n12965) );
  OAI211_X1 U15377 ( .C1(n13059), .C2(n12971), .A(n12966), .B(n12965), .ZN(
        P3_U3476) );
  MUX2_X1 U15378 ( .A(n12967), .B(n13060), .S(n15665), .Z(n12970) );
  NAND2_X1 U15379 ( .A1(n13062), .A2(n12968), .ZN(n12969) );
  OAI211_X1 U15380 ( .C1(n13066), .C2(n12971), .A(n12970), .B(n12969), .ZN(
        P3_U3475) );
  AOI21_X1 U15381 ( .B1(n12973), .B2(n15630), .A(n12972), .ZN(n13067) );
  MUX2_X1 U15382 ( .A(n12974), .B(n13067), .S(n15665), .Z(n12975) );
  OAI21_X1 U15383 ( .B1(n13071), .B2(n12976), .A(n12975), .ZN(P3_U3474) );
  XNOR2_X1 U15384 ( .A(n10074), .B(n12977), .ZN(n15614) );
  NAND2_X1 U15385 ( .A1(n15614), .A2(n12978), .ZN(n12989) );
  NAND2_X1 U15386 ( .A1(n12981), .A2(n12980), .ZN(n12984) );
  NAND2_X1 U15387 ( .A1(n9514), .A2(n12982), .ZN(n12983) );
  NAND2_X1 U15388 ( .A1(n12984), .A2(n12983), .ZN(n12985) );
  AOI21_X1 U15389 ( .B1(n12987), .B2(n12986), .A(n12985), .ZN(n12988) );
  AND2_X1 U15390 ( .A1(n12989), .A2(n12988), .ZN(n15611) );
  NOR2_X1 U15391 ( .A1(n12990), .A2(n15626), .ZN(n15606) );
  AOI21_X1 U15392 ( .B1(n15614), .B2(n6643), .A(n15606), .ZN(n12991) );
  AND2_X1 U15393 ( .A1(n15611), .A2(n12991), .ZN(n15622) );
  INV_X1 U15394 ( .A(n15622), .ZN(n12992) );
  MUX2_X1 U15395 ( .A(n12992), .B(P3_REG1_REG_2__SCAN_IN), .S(n15663), .Z(
        P3_U3461) );
  NAND2_X1 U15396 ( .A1(n12375), .A2(n13061), .ZN(n12994) );
  NAND2_X1 U15397 ( .A1(n12993), .A2(n15654), .ZN(n12996) );
  OAI211_X1 U15398 ( .C1(n15654), .C2(n12995), .A(n12994), .B(n12996), .ZN(
        P3_U3458) );
  NAND2_X1 U15399 ( .A1(n15653), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n12997) );
  OAI211_X1 U15400 ( .C1(n12998), .C2(n13070), .A(n12997), .B(n12996), .ZN(
        P3_U3457) );
  MUX2_X1 U15401 ( .A(n13000), .B(n12999), .S(n15654), .Z(n13003) );
  NAND2_X1 U15402 ( .A1(n13001), .A2(n13061), .ZN(n13002) );
  OAI211_X1 U15403 ( .C1(n13004), .C2(n13065), .A(n13003), .B(n13002), .ZN(
        P3_U3455) );
  MUX2_X1 U15404 ( .A(n13007), .B(n13006), .S(n15654), .Z(n13010) );
  NAND2_X1 U15405 ( .A1(n13008), .A2(n13061), .ZN(n13009) );
  OAI211_X1 U15406 ( .C1(n13011), .C2(n13065), .A(n13010), .B(n13009), .ZN(
        P3_U3453) );
  OAI22_X1 U15407 ( .A1(n13013), .A2(n13065), .B1(n13012), .B2(n13070), .ZN(
        n13016) );
  MUX2_X1 U15408 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n13014), .S(n15654), .Z(
        n13015) );
  OR2_X1 U15409 ( .A1(n13016), .A2(n13015), .ZN(P3_U3452) );
  INV_X1 U15410 ( .A(n13017), .ZN(n13019) );
  MUX2_X1 U15411 ( .A(n13019), .B(n13018), .S(n15653), .Z(n13022) );
  NAND2_X1 U15412 ( .A1(n13020), .A2(n13061), .ZN(n13021) );
  OAI211_X1 U15413 ( .C1(n13023), .C2(n13065), .A(n13022), .B(n13021), .ZN(
        P3_U3451) );
  MUX2_X1 U15414 ( .A(P3_REG0_REG_23__SCAN_IN), .B(n13024), .S(n15654), .Z(
        P3_U3450) );
  MUX2_X1 U15415 ( .A(n13026), .B(n13025), .S(n15654), .Z(n13029) );
  NAND2_X1 U15416 ( .A1(n13027), .A2(n13061), .ZN(n13028) );
  OAI211_X1 U15417 ( .C1(n13030), .C2(n13065), .A(n13029), .B(n13028), .ZN(
        P3_U3449) );
  MUX2_X1 U15418 ( .A(n15799), .B(n13031), .S(n15654), .Z(n13034) );
  NAND2_X1 U15419 ( .A1(n13032), .A2(n13061), .ZN(n13033) );
  OAI211_X1 U15420 ( .C1(n13035), .C2(n13065), .A(n13034), .B(n13033), .ZN(
        P3_U3448) );
  MUX2_X1 U15421 ( .A(n13037), .B(n13036), .S(n15653), .Z(n13040) );
  NAND2_X1 U15422 ( .A1(n13038), .A2(n13061), .ZN(n13039) );
  OAI211_X1 U15423 ( .C1(n13041), .C2(n13065), .A(n13040), .B(n13039), .ZN(
        P3_U3447) );
  INV_X1 U15424 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13043) );
  MUX2_X1 U15425 ( .A(n13043), .B(n13042), .S(n15654), .Z(n13046) );
  NAND2_X1 U15426 ( .A1(n13044), .A2(n13061), .ZN(n13045) );
  OAI211_X1 U15427 ( .C1(n13047), .C2(n13065), .A(n13046), .B(n13045), .ZN(
        P3_U3446) );
  MUX2_X1 U15428 ( .A(n13049), .B(n13048), .S(n15654), .Z(n13052) );
  NAND2_X1 U15429 ( .A1(n13050), .A2(n13061), .ZN(n13051) );
  OAI211_X1 U15430 ( .C1(n13053), .C2(n13065), .A(n13052), .B(n13051), .ZN(
        P3_U3444) );
  INV_X1 U15431 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13055) );
  MUX2_X1 U15432 ( .A(n13055), .B(n13054), .S(n15654), .Z(n13058) );
  NAND2_X1 U15433 ( .A1(n13056), .A2(n13061), .ZN(n13057) );
  OAI211_X1 U15434 ( .C1(n13059), .C2(n13065), .A(n13058), .B(n13057), .ZN(
        P3_U3441) );
  MUX2_X1 U15435 ( .A(n15696), .B(n13060), .S(n15654), .Z(n13064) );
  NAND2_X1 U15436 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  OAI211_X1 U15437 ( .C1(n13066), .C2(n13065), .A(n13064), .B(n13063), .ZN(
        P3_U3438) );
  INV_X1 U15438 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n13068) );
  MUX2_X1 U15439 ( .A(n13068), .B(n13067), .S(n15654), .Z(n13069) );
  OAI21_X1 U15440 ( .B1(n13071), .B2(n13070), .A(n13069), .ZN(P3_U3435) );
  MUX2_X1 U15441 ( .A(n10578), .B(P3_D_REG_0__SCAN_IN), .S(n13072), .Z(
        P3_U3376) );
  INV_X1 U15442 ( .A(n13073), .ZN(n13079) );
  INV_X1 U15443 ( .A(n13095), .ZN(n13077) );
  NOR4_X1 U15444 ( .A1(n13075), .A2(P3_IR_REG_30__SCAN_IN), .A3(n13074), .A4(
        P3_U3151), .ZN(n13076) );
  AOI21_X1 U15445 ( .B1(SI_31_), .B2(n13077), .A(n13076), .ZN(n13078) );
  OAI21_X1 U15446 ( .B1(n13079), .B2(n13090), .A(n13078), .ZN(P3_U3264) );
  INV_X1 U15447 ( .A(n13080), .ZN(n13083) );
  OAI222_X1 U15448 ( .A1(n13090), .A2(n13083), .B1(n13095), .B2(n13082), .C1(
        P3_U3151), .C2(n13081), .ZN(P3_U3267) );
  INV_X1 U15449 ( .A(n13084), .ZN(n13087) );
  INV_X1 U15450 ( .A(SI_27_), .ZN(n13086) );
  OAI222_X1 U15451 ( .A1(n13090), .A2(n13087), .B1(n13095), .B2(n13086), .C1(
        P3_U3151), .C2(n7168), .ZN(P3_U3268) );
  INV_X1 U15452 ( .A(n13088), .ZN(n13089) );
  OAI222_X1 U15453 ( .A1(P3_U3151), .A2(n10037), .B1(n13095), .B2(n13091), 
        .C1(n13090), .C2(n13089), .ZN(P3_U3269) );
  INV_X1 U15454 ( .A(n13092), .ZN(n13093) );
  OAI222_X1 U15455 ( .A1(P3_U3151), .A2(n13096), .B1(n13095), .B2(n13094), 
        .C1(n13090), .C2(n13093), .ZN(P3_U3270) );
  MUX2_X1 U15456 ( .A(n13098), .B(n13097), .S(P3_STATE_REG_SCAN_IN), .Z(
        P3_U3271) );
  INV_X1 U15457 ( .A(n13099), .ZN(n13212) );
  NOR3_X1 U15458 ( .A1(n13100), .A2(n13552), .A3(n13256), .ZN(n13101) );
  AOI21_X1 U15459 ( .B1(n13212), .B2(n13270), .A(n13101), .ZN(n13109) );
  AOI22_X1 U15460 ( .A1(n13230), .A2(n13879), .B1(n13229), .B2(n13881), .ZN(
        n13103) );
  OAI211_X1 U15461 ( .C1(n13277), .C2(n13886), .A(n13103), .B(n13102), .ZN(
        n13106) );
  NOR2_X1 U15462 ( .A1(n13104), .A2(n13250), .ZN(n13105) );
  AOI211_X1 U15463 ( .C1(n14009), .C2(n13280), .A(n13106), .B(n13105), .ZN(
        n13107) );
  OAI21_X1 U15464 ( .B1(n13109), .B2(n13108), .A(n13107), .ZN(P2_U3187) );
  NAND2_X1 U15465 ( .A1(n13219), .A2(n13111), .ZN(n13113) );
  XNOR2_X1 U15466 ( .A(n13113), .B(n13112), .ZN(n13116) );
  OAI22_X1 U15467 ( .A1(n13116), .A2(n13250), .B1(n13437), .B2(n13256), .ZN(
        n13114) );
  OAI21_X1 U15468 ( .B1(n13116), .B2(n13115), .A(n13114), .ZN(n13122) );
  AOI22_X1 U15469 ( .A1(n13719), .A2(n13880), .B1(n13878), .B2(n13594), .ZN(
        n13750) );
  INV_X1 U15470 ( .A(n13750), .ZN(n13120) );
  INV_X1 U15471 ( .A(n13752), .ZN(n13118) );
  OAI22_X1 U15472 ( .A1(n13118), .A2(n13277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13117), .ZN(n13119) );
  AOI21_X1 U15473 ( .B1(n13120), .B2(n13275), .A(n13119), .ZN(n13121) );
  OAI211_X1 U15474 ( .C1(n13758), .C2(n13227), .A(n13122), .B(n13121), .ZN(
        P2_U3188) );
  INV_X1 U15475 ( .A(n13123), .ZN(n13249) );
  NOR3_X1 U15476 ( .A1(n13124), .A2(n13126), .A3(n13256), .ZN(n13125) );
  AOI21_X1 U15477 ( .B1(n13249), .B2(n13270), .A(n13125), .ZN(n13134) );
  NOR2_X1 U15478 ( .A1(n13126), .A2(n13273), .ZN(n13127) );
  AOI21_X1 U15479 ( .B1(n13595), .B2(n13880), .A(n13127), .ZN(n13976) );
  NAND2_X1 U15480 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13674)
         );
  INV_X1 U15481 ( .A(n13128), .ZN(n13798) );
  NAND2_X1 U15482 ( .A1(n13261), .A2(n13798), .ZN(n13129) );
  OAI211_X1 U15483 ( .C1(n13976), .C2(n13263), .A(n13674), .B(n13129), .ZN(
        n13131) );
  NOR2_X1 U15484 ( .A1(n13206), .A2(n13250), .ZN(n13130) );
  AOI211_X1 U15485 ( .C1(n14065), .C2(n13280), .A(n13131), .B(n13130), .ZN(
        n13132) );
  OAI21_X1 U15486 ( .B1(n13134), .B2(n13133), .A(n13132), .ZN(P2_U3191) );
  NOR2_X1 U15487 ( .A1(n13135), .A2(n13256), .ZN(n13137) );
  AOI22_X1 U15488 ( .A1(n13138), .A2(n13270), .B1(n13137), .B2(n13136), .ZN(
        n13152) );
  NAND2_X1 U15489 ( .A1(n13590), .A2(n6409), .ZN(n13140) );
  XNOR2_X1 U15490 ( .A(n13140), .B(n13139), .ZN(n13141) );
  XNOR2_X1 U15491 ( .A(n13456), .B(n13141), .ZN(n13151) );
  OAI22_X1 U15492 ( .A1(n13143), .A2(n13277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13142), .ZN(n13145) );
  NOR2_X1 U15493 ( .A1(n6880), .A2(n13227), .ZN(n13144) );
  AOI211_X1 U15494 ( .C1(n13275), .C2(n13146), .A(n13145), .B(n13144), .ZN(
        n13150) );
  NAND4_X1 U15495 ( .A1(n13148), .A2(n13270), .A3(n13147), .A4(n13151), .ZN(
        n13149) );
  OAI211_X1 U15496 ( .C1(n13152), .C2(n13151), .A(n13150), .B(n13149), .ZN(
        P2_U3192) );
  AOI21_X1 U15497 ( .B1(n13154), .B2(n13153), .A(n13250), .ZN(n13156) );
  NAND2_X1 U15498 ( .A1(n13156), .A2(n13155), .ZN(n13160) );
  AOI22_X1 U15499 ( .A1(n13594), .A2(n13880), .B1(n13878), .B2(n13595), .ZN(
        n13768) );
  OAI22_X1 U15500 ( .A1(n13768), .A2(n13263), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13157), .ZN(n13158) );
  AOI21_X1 U15501 ( .B1(n13772), .B2(n13261), .A(n13158), .ZN(n13159) );
  OAI211_X1 U15502 ( .C1(n6876), .C2(n13227), .A(n13160), .B(n13159), .ZN(
        P2_U3195) );
  NAND3_X1 U15503 ( .A1(n13161), .A2(n13269), .A3(n13719), .ZN(n13164) );
  OAI21_X1 U15504 ( .B1(n13179), .B2(n13162), .A(n13270), .ZN(n13163) );
  AOI21_X1 U15505 ( .B1(n13164), .B2(n13163), .A(n6498), .ZN(n13168) );
  INV_X1 U15506 ( .A(n13722), .ZN(n14053) );
  AOI22_X1 U15507 ( .A1(n13726), .A2(n13261), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13166) );
  AOI22_X1 U15508 ( .A1(n13720), .A2(n13229), .B1(n13230), .B2(n13719), .ZN(
        n13165) );
  OAI211_X1 U15509 ( .C1(n14053), .C2(n13227), .A(n13166), .B(n13165), .ZN(
        n13167) );
  OR2_X1 U15510 ( .A1(n13168), .A2(n13167), .ZN(P2_U3197) );
  AOI21_X1 U15511 ( .B1(n13171), .B2(n13170), .A(n13169), .ZN(n13175) );
  OAI22_X1 U15512 ( .A1(n13409), .A2(n13274), .B1(n13392), .B2(n13273), .ZN(
        n13852) );
  NAND2_X1 U15513 ( .A1(n13275), .A2(n13852), .ZN(n13172) );
  NAND2_X1 U15514 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n15483)
         );
  OAI211_X1 U15515 ( .C1(n13277), .C2(n13854), .A(n13172), .B(n15483), .ZN(
        n13173) );
  AOI21_X1 U15516 ( .B1(n13996), .B2(n13280), .A(n13173), .ZN(n13174) );
  OAI21_X1 U15517 ( .B1(n13175), .B2(n13250), .A(n13174), .ZN(P2_U3198) );
  NOR2_X1 U15518 ( .A1(n13437), .A2(n13273), .ZN(n13176) );
  AOI21_X1 U15519 ( .B1(n13592), .B2(n13880), .A(n13176), .ZN(n13738) );
  INV_X1 U15520 ( .A(n13741), .ZN(n13177) );
  AOI22_X1 U15521 ( .A1(n13177), .A2(n13261), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13178) );
  OAI21_X1 U15522 ( .B1(n13738), .B2(n13263), .A(n13178), .ZN(n13182) );
  AOI211_X1 U15523 ( .C1(n6605), .C2(n13180), .A(n13250), .B(n13179), .ZN(
        n13181) );
  AOI211_X1 U15524 ( .C1(n13948), .C2(n13280), .A(n13182), .B(n13181), .ZN(
        n13183) );
  INV_X1 U15525 ( .A(n13183), .ZN(P2_U3201) );
  NOR2_X1 U15526 ( .A1(n13277), .A2(n13184), .ZN(n13186) );
  NAND2_X1 U15527 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n15405) );
  OAI21_X1 U15528 ( .B1(n13227), .B2(n7013), .A(n15405), .ZN(n13185) );
  AOI211_X1 U15529 ( .C1(n13229), .C2(n13607), .A(n13186), .B(n13185), .ZN(
        n13195) );
  OAI21_X1 U15530 ( .B1(n13188), .B2(n13190), .A(n13187), .ZN(n13189) );
  NAND2_X1 U15531 ( .A1(n13270), .A2(n13189), .ZN(n13194) );
  NOR3_X1 U15532 ( .A1(n13256), .A2(n13191), .A3(n13190), .ZN(n13192) );
  OAI21_X1 U15533 ( .B1(n13192), .B2(n13230), .A(n13609), .ZN(n13193) );
  NAND3_X1 U15534 ( .A1(n13195), .A2(n13194), .A3(n13193), .ZN(P2_U3202) );
  INV_X1 U15535 ( .A(n13788), .ZN(n13197) );
  OAI22_X1 U15536 ( .A1(n13197), .A2(n13277), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13196), .ZN(n13201) );
  INV_X1 U15537 ( .A(n13230), .ZN(n13199) );
  OAI22_X1 U15538 ( .A1(n13203), .A2(n13199), .B1(n13198), .B2(n13430), .ZN(
        n13200) );
  AOI211_X1 U15539 ( .C1(n13972), .C2(n13280), .A(n13201), .B(n13200), .ZN(
        n13209) );
  INV_X1 U15540 ( .A(n13202), .ZN(n13207) );
  OAI22_X1 U15541 ( .A1(n13204), .A2(n13250), .B1(n13203), .B2(n13256), .ZN(
        n13205) );
  NAND3_X1 U15542 ( .A1(n13207), .A2(n13206), .A3(n13205), .ZN(n13208) );
  OAI211_X1 U15543 ( .C1(n13210), .C2(n13250), .A(n13209), .B(n13208), .ZN(
        P2_U3205) );
  OAI22_X1 U15544 ( .A1(n13386), .A2(n13274), .B1(n13372), .B2(n13273), .ZN(
        n13896) );
  AOI22_X1 U15545 ( .A1(n13275), .A2(n13896), .B1(P2_REG3_REG_13__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13211) );
  OAI21_X1 U15546 ( .B1(n13901), .B2(n13277), .A(n13211), .ZN(n13216) );
  AOI211_X1 U15547 ( .C1(n13214), .C2(n13213), .A(n13250), .B(n13212), .ZN(
        n13215) );
  AOI211_X1 U15548 ( .C1(n14014), .C2(n13280), .A(n13216), .B(n13215), .ZN(
        n13217) );
  INV_X1 U15549 ( .A(n13217), .ZN(P2_U3206) );
  OAI22_X1 U15550 ( .A1(n13218), .A2(n13250), .B1(n13426), .B2(n13256), .ZN(
        n13220) );
  NAND2_X1 U15551 ( .A1(n13220), .A2(n13219), .ZN(n13226) );
  OAI22_X1 U15552 ( .A1(n13222), .A2(n13263), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13221), .ZN(n13223) );
  AOI21_X1 U15553 ( .B1(n13224), .B2(n13261), .A(n13223), .ZN(n13225) );
  OAI211_X1 U15554 ( .C1(n13228), .C2(n13227), .A(n13226), .B(n13225), .ZN(
        P2_U3207) );
  OAI22_X1 U15555 ( .A1(n8651), .A2(n13256), .B1(n13250), .B2(n13237), .ZN(
        n13234) );
  XNOR2_X1 U15556 ( .A(n13232), .B(n13231), .ZN(n13240) );
  NAND3_X1 U15557 ( .A1(n13234), .A2(n13240), .A3(n13233), .ZN(n13246) );
  INV_X1 U15558 ( .A(n13235), .ZN(n13236) );
  AOI22_X1 U15559 ( .A1(n13280), .A2(n6751), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n13236), .ZN(n13245) );
  INV_X1 U15560 ( .A(n13237), .ZN(n13239) );
  NOR2_X1 U15561 ( .A1(n13239), .A2(n13238), .ZN(n13242) );
  INV_X1 U15562 ( .A(n13240), .ZN(n13241) );
  OAI211_X1 U15563 ( .C1(n13243), .C2(n13242), .A(n13270), .B(n13241), .ZN(
        n13244) );
  NAND4_X1 U15564 ( .A1(n13247), .A2(n13246), .A3(n13245), .A4(n13244), .ZN(
        P2_U3209) );
  AOI22_X1 U15565 ( .A1(n13782), .A2(n13880), .B1(n13878), .B2(n13597), .ZN(
        n13814) );
  NAND2_X1 U15566 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13646)
         );
  NAND2_X1 U15567 ( .A1(n13261), .A2(n13822), .ZN(n13248) );
  OAI211_X1 U15568 ( .C1(n13814), .C2(n13263), .A(n13646), .B(n13248), .ZN(
        n13254) );
  AOI211_X1 U15569 ( .C1(n13252), .C2(n13251), .A(n13250), .B(n13249), .ZN(
        n13253) );
  AOI211_X1 U15570 ( .C1(n13821), .C2(n13280), .A(n13254), .B(n13253), .ZN(
        n13255) );
  INV_X1 U15571 ( .A(n13255), .ZN(P2_U3210) );
  NOR3_X1 U15572 ( .A1(n13258), .A2(n13257), .A3(n13256), .ZN(n13259) );
  AOI21_X1 U15573 ( .B1(n6498), .B2(n13270), .A(n13259), .ZN(n13268) );
  AOI22_X1 U15574 ( .A1(n13591), .A2(n13880), .B1(n13878), .B2(n13592), .ZN(
        n13705) );
  INV_X1 U15575 ( .A(n13260), .ZN(n13709) );
  AOI22_X1 U15576 ( .A1(n13709), .A2(n13261), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13262) );
  OAI21_X1 U15577 ( .B1(n13705), .B2(n13263), .A(n13262), .ZN(n13265) );
  AOI211_X1 U15578 ( .C1(n13940), .C2(n13280), .A(n13265), .B(n13264), .ZN(
        n13266) );
  OAI21_X1 U15579 ( .B1(n13268), .B2(n13267), .A(n13266), .ZN(P2_U3212) );
  AOI22_X1 U15580 ( .A1(n13271), .A2(n13270), .B1(n13269), .B2(n13881), .ZN(
        n13283) );
  INV_X1 U15581 ( .A(n13272), .ZN(n13282) );
  INV_X1 U15582 ( .A(n13872), .ZN(n13278) );
  OAI22_X1 U15583 ( .A1(n13397), .A2(n13274), .B1(n13386), .B2(n13273), .ZN(
        n14001) );
  AOI22_X1 U15584 ( .A1(n13275), .A2(n14001), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13276) );
  OAI21_X1 U15585 ( .B1(n13278), .B2(n13277), .A(n13276), .ZN(n13279) );
  AOI21_X1 U15586 ( .B1(n13866), .B2(n13280), .A(n13279), .ZN(n13281) );
  OAI21_X1 U15587 ( .B1(n13283), .B2(n13282), .A(n13281), .ZN(P2_U3213) );
  AOI22_X1 U15588 ( .A1(n13286), .A2(n13474), .B1(n13609), .B2(n6440), .ZN(
        n13317) );
  NAND2_X1 U15589 ( .A1(n13286), .A2(n6440), .ZN(n13288) );
  NAND2_X1 U15590 ( .A1(n13609), .A2(n13474), .ZN(n13287) );
  NAND2_X1 U15591 ( .A1(n13288), .A2(n13287), .ZN(n13316) );
  OR2_X1 U15592 ( .A1(n8651), .A2(n13474), .ZN(n13290) );
  NAND2_X1 U15593 ( .A1(n13474), .A2(n13916), .ZN(n13289) );
  OR2_X1 U15594 ( .A1(n8651), .A2(n6440), .ZN(n13292) );
  NAND2_X1 U15595 ( .A1(n6440), .A2(n13916), .ZN(n13291) );
  NAND2_X1 U15596 ( .A1(n13292), .A2(n13291), .ZN(n13307) );
  OR2_X1 U15597 ( .A1(n13293), .A2(n13474), .ZN(n13297) );
  INV_X1 U15598 ( .A(n13297), .ZN(n13300) );
  MUX2_X1 U15599 ( .A(n13293), .B(n13474), .S(n13296), .Z(n13299) );
  AOI21_X1 U15600 ( .B1(n13672), .B2(n13294), .A(n13571), .ZN(n13295) );
  OAI21_X1 U15601 ( .B1(n13297), .B2(n13296), .A(n13295), .ZN(n13298) );
  OAI21_X1 U15602 ( .B1(n13300), .B2(n13299), .A(n13298), .ZN(n13301) );
  OAI21_X1 U15603 ( .B1(n13308), .B2(n13307), .A(n13301), .ZN(n13311) );
  OR2_X1 U15604 ( .A1(n13304), .A2(n13474), .ZN(n13303) );
  NAND2_X1 U15605 ( .A1(n13474), .A2(n6751), .ZN(n13302) );
  OR2_X1 U15606 ( .A1(n13304), .A2(n6440), .ZN(n13306) );
  NAND2_X1 U15607 ( .A1(n6751), .A2(n6440), .ZN(n13305) );
  NAND2_X1 U15608 ( .A1(n13306), .A2(n13305), .ZN(n13312) );
  NAND2_X1 U15609 ( .A1(n13313), .A2(n13312), .ZN(n13310) );
  NAND2_X1 U15610 ( .A1(n13308), .A2(n13307), .ZN(n13309) );
  INV_X1 U15611 ( .A(n13312), .ZN(n13315) );
  INV_X1 U15612 ( .A(n13313), .ZN(n13314) );
  NAND2_X1 U15613 ( .A1(n13320), .A2(n6440), .ZN(n13319) );
  NAND2_X1 U15614 ( .A1(n13608), .A2(n13492), .ZN(n13318) );
  NAND2_X1 U15615 ( .A1(n13319), .A2(n13318), .ZN(n13321) );
  AOI22_X1 U15616 ( .A1(n13320), .A2(n13492), .B1(n13608), .B2(n6440), .ZN(
        n13322) );
  INV_X1 U15617 ( .A(n13321), .ZN(n13324) );
  INV_X1 U15618 ( .A(n13322), .ZN(n13323) );
  NAND2_X1 U15619 ( .A1(n13324), .A2(n13323), .ZN(n13325) );
  NAND2_X1 U15620 ( .A1(n13328), .A2(n13492), .ZN(n13327) );
  OR2_X1 U15621 ( .A1(n13330), .A2(n13492), .ZN(n13326) );
  NAND2_X1 U15622 ( .A1(n13328), .A2(n6440), .ZN(n13329) );
  OAI21_X1 U15623 ( .B1(n13330), .B2(n6440), .A(n13329), .ZN(n13331) );
  NAND2_X1 U15624 ( .A1(n14036), .A2(n6440), .ZN(n13333) );
  NAND2_X1 U15625 ( .A1(n13606), .A2(n13492), .ZN(n13332) );
  NAND2_X1 U15626 ( .A1(n13333), .A2(n13332), .ZN(n13335) );
  NAND2_X1 U15627 ( .A1(n13336), .A2(n13335), .ZN(n13334) );
  INV_X1 U15628 ( .A(n13335), .ZN(n13338) );
  INV_X1 U15629 ( .A(n13336), .ZN(n13337) );
  NAND2_X1 U15630 ( .A1(n15525), .A2(n13474), .ZN(n13341) );
  OR2_X1 U15631 ( .A1(n13343), .A2(n13492), .ZN(n13340) );
  NAND2_X1 U15632 ( .A1(n15525), .A2(n6440), .ZN(n13342) );
  OAI21_X1 U15633 ( .B1(n13343), .B2(n6440), .A(n13342), .ZN(n13344) );
  NAND2_X1 U15634 ( .A1(n14031), .A2(n6440), .ZN(n13347) );
  OR2_X1 U15635 ( .A1(n13345), .A2(n6440), .ZN(n13346) );
  NAND2_X1 U15636 ( .A1(n13347), .A2(n13346), .ZN(n13349) );
  AOI22_X1 U15637 ( .A1(n14031), .A2(n13474), .B1(n13604), .B2(n6440), .ZN(
        n13348) );
  NAND2_X1 U15638 ( .A1(n13352), .A2(n13492), .ZN(n13351) );
  NAND2_X1 U15639 ( .A1(n13603), .A2(n6440), .ZN(n13350) );
  NAND2_X1 U15640 ( .A1(n13351), .A2(n13350), .ZN(n13354) );
  AOI22_X1 U15641 ( .A1(n13352), .A2(n6440), .B1(n13474), .B2(n13603), .ZN(
        n13353) );
  AOI21_X1 U15642 ( .B1(n13355), .B2(n13354), .A(n13353), .ZN(n13357) );
  NOR2_X1 U15643 ( .A1(n13355), .A2(n13354), .ZN(n13356) );
  NAND2_X1 U15644 ( .A1(n14026), .A2(n6440), .ZN(n13360) );
  OR2_X1 U15645 ( .A1(n13358), .A2(n6440), .ZN(n13359) );
  AOI22_X1 U15646 ( .A1(n14026), .A2(n13492), .B1(n13602), .B2(n6440), .ZN(
        n13361) );
  NAND2_X1 U15647 ( .A1(n13365), .A2(n13492), .ZN(n13364) );
  NAND2_X1 U15648 ( .A1(n13601), .A2(n6440), .ZN(n13363) );
  NAND2_X1 U15649 ( .A1(n13365), .A2(n6440), .ZN(n13366) );
  OAI21_X1 U15650 ( .B1(n13367), .B2(n6440), .A(n13366), .ZN(n13368) );
  NAND2_X1 U15651 ( .A1(n14085), .A2(n6440), .ZN(n13371) );
  NAND2_X1 U15652 ( .A1(n13600), .A2(n13474), .ZN(n13370) );
  NAND2_X1 U15653 ( .A1(n13371), .A2(n13370), .ZN(n13375) );
  NOR2_X1 U15654 ( .A1(n13372), .A2(n13492), .ZN(n13373) );
  AOI21_X1 U15655 ( .B1(n14085), .B2(n13492), .A(n13373), .ZN(n13374) );
  NAND2_X1 U15656 ( .A1(n14014), .A2(n6402), .ZN(n13377) );
  NAND2_X1 U15657 ( .A1(n13879), .A2(n6440), .ZN(n13376) );
  NAND2_X1 U15658 ( .A1(n13377), .A2(n13376), .ZN(n13379) );
  AOI22_X1 U15659 ( .A1(n14014), .A2(n6440), .B1(n13474), .B2(n13879), .ZN(
        n13378) );
  AOI21_X1 U15660 ( .B1(n13380), .B2(n13379), .A(n13378), .ZN(n13382) );
  NOR2_X1 U15661 ( .A1(n13380), .A2(n13379), .ZN(n13381) );
  NAND2_X1 U15662 ( .A1(n14009), .A2(n6440), .ZN(n13384) );
  NAND2_X1 U15663 ( .A1(n13599), .A2(n6402), .ZN(n13383) );
  NAND2_X1 U15664 ( .A1(n13384), .A2(n13383), .ZN(n13388) );
  NAND2_X1 U15665 ( .A1(n14009), .A2(n13492), .ZN(n13385) );
  OAI21_X1 U15666 ( .B1(n13386), .B2(n13492), .A(n13385), .ZN(n13387) );
  NAND2_X1 U15667 ( .A1(n13866), .A2(n13492), .ZN(n13390) );
  NAND2_X1 U15668 ( .A1(n13881), .A2(n6440), .ZN(n13389) );
  NAND2_X1 U15669 ( .A1(n13866), .A2(n6440), .ZN(n13391) );
  OAI21_X1 U15670 ( .B1(n13392), .B2(n6440), .A(n13391), .ZN(n13393) );
  NAND2_X1 U15671 ( .A1(n13996), .A2(n6440), .ZN(n13395) );
  NAND2_X1 U15672 ( .A1(n13598), .A2(n13492), .ZN(n13394) );
  NAND2_X1 U15673 ( .A1(n13395), .A2(n13394), .ZN(n13401) );
  NAND2_X1 U15674 ( .A1(n13400), .A2(n13401), .ZN(n13399) );
  NAND2_X1 U15675 ( .A1(n13996), .A2(n13492), .ZN(n13396) );
  OAI21_X1 U15676 ( .B1(n13397), .B2(n13492), .A(n13396), .ZN(n13398) );
  NAND2_X1 U15677 ( .A1(n13399), .A2(n13398), .ZN(n13405) );
  INV_X1 U15678 ( .A(n13400), .ZN(n13403) );
  INV_X1 U15679 ( .A(n13401), .ZN(n13402) );
  NAND2_X1 U15680 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  NAND2_X1 U15681 ( .A1(n14073), .A2(n13492), .ZN(n13407) );
  NAND2_X1 U15682 ( .A1(n13597), .A2(n6440), .ZN(n13406) );
  NAND2_X1 U15683 ( .A1(n14073), .A2(n6440), .ZN(n13408) );
  OAI21_X1 U15684 ( .B1(n13409), .B2(n6440), .A(n13408), .ZN(n13410) );
  NAND2_X1 U15685 ( .A1(n13821), .A2(n6440), .ZN(n13412) );
  NAND2_X1 U15686 ( .A1(n13596), .A2(n13492), .ZN(n13411) );
  AOI22_X1 U15687 ( .A1(n13821), .A2(n13474), .B1(n13596), .B2(n6440), .ZN(
        n13413) );
  NAND2_X1 U15688 ( .A1(n14065), .A2(n13492), .ZN(n13415) );
  NAND2_X1 U15689 ( .A1(n13782), .A2(n6440), .ZN(n13414) );
  NAND2_X1 U15690 ( .A1(n13415), .A2(n13414), .ZN(n13417) );
  AOI22_X1 U15691 ( .A1(n14065), .A2(n6440), .B1(n13474), .B2(n13782), .ZN(
        n13416) );
  NAND2_X1 U15692 ( .A1(n13972), .A2(n6440), .ZN(n13419) );
  NAND2_X1 U15693 ( .A1(n13595), .A2(n13492), .ZN(n13418) );
  NAND2_X1 U15694 ( .A1(n13419), .A2(n13418), .ZN(n13423) );
  NAND2_X1 U15695 ( .A1(n13972), .A2(n13492), .ZN(n13420) );
  OAI21_X1 U15696 ( .B1(n13421), .B2(n13492), .A(n13420), .ZN(n13422) );
  NAND2_X1 U15697 ( .A1(n13432), .A2(n13492), .ZN(n13425) );
  NAND2_X1 U15698 ( .A1(n13783), .A2(n6440), .ZN(n13424) );
  NAND2_X1 U15699 ( .A1(n13425), .A2(n13424), .ZN(n13434) );
  NOR2_X1 U15700 ( .A1(n13426), .A2(n6440), .ZN(n13427) );
  AOI21_X1 U15701 ( .B1(n14058), .B2(n6440), .A(n13427), .ZN(n13441) );
  NAND2_X1 U15702 ( .A1(n14058), .A2(n13492), .ZN(n13429) );
  NAND2_X1 U15703 ( .A1(n13594), .A2(n6440), .ZN(n13428) );
  NAND2_X1 U15704 ( .A1(n13429), .A2(n13428), .ZN(n13440) );
  NOR2_X1 U15705 ( .A1(n13430), .A2(n6440), .ZN(n13431) );
  AOI21_X1 U15706 ( .B1(n13432), .B2(n6440), .A(n13431), .ZN(n13433) );
  AOI21_X1 U15707 ( .B1(n13435), .B2(n13434), .A(n13433), .ZN(n13443) );
  NOR2_X1 U15708 ( .A1(n13437), .A2(n6440), .ZN(n13436) );
  AOI21_X1 U15709 ( .B1(n13956), .B2(n6440), .A(n13436), .ZN(n13480) );
  NAND2_X1 U15710 ( .A1(n13956), .A2(n13492), .ZN(n13439) );
  OR2_X1 U15711 ( .A1(n13437), .A2(n6402), .ZN(n13438) );
  NAND2_X1 U15712 ( .A1(n13439), .A2(n13438), .ZN(n13479) );
  AOI22_X1 U15713 ( .A1(n13441), .A2(n13440), .B1(n13480), .B2(n13479), .ZN(
        n13442) );
  OAI21_X1 U15714 ( .B1(n13444), .B2(n13443), .A(n13442), .ZN(n13485) );
  MUX2_X1 U15715 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n7875), .Z(n13447) );
  XNOR2_X1 U15716 ( .A(n13447), .B(SI_31_), .ZN(n13448) );
  NAND2_X1 U15717 ( .A1(n14474), .A2(n8146), .ZN(n13450) );
  NAND2_X1 U15718 ( .A1(n13496), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n13449) );
  NAND2_X1 U15719 ( .A1(n8596), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13454) );
  INV_X1 U15720 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n15695) );
  OR2_X1 U15721 ( .A1(n8239), .A2(n15695), .ZN(n13453) );
  INV_X1 U15722 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n14041) );
  OR2_X1 U15723 ( .A1(n8077), .A2(n14041), .ZN(n13452) );
  AND3_X1 U15724 ( .A1(n13454), .A2(n13453), .A3(n13452), .ZN(n13530) );
  AND2_X1 U15725 ( .A1(n13590), .A2(n13474), .ZN(n13455) );
  NAND2_X1 U15726 ( .A1(n13456), .A2(n13492), .ZN(n13458) );
  NAND2_X1 U15727 ( .A1(n13590), .A2(n6440), .ZN(n13457) );
  NAND2_X1 U15728 ( .A1(n13458), .A2(n13457), .ZN(n13510) );
  AND2_X1 U15729 ( .A1(n13589), .A2(n6440), .ZN(n13459) );
  AOI21_X1 U15730 ( .B1(n13460), .B2(n13492), .A(n13459), .ZN(n13507) );
  NAND2_X1 U15731 ( .A1(n13460), .A2(n6440), .ZN(n13462) );
  NAND2_X1 U15732 ( .A1(n13589), .A2(n13492), .ZN(n13461) );
  NAND2_X1 U15733 ( .A1(n13462), .A2(n13461), .ZN(n13506) );
  NAND2_X1 U15734 ( .A1(n13507), .A2(n13506), .ZN(n13511) );
  AND2_X1 U15735 ( .A1(n13591), .A2(n6440), .ZN(n13463) );
  AOI21_X1 U15736 ( .B1(n13933), .B2(n13492), .A(n13463), .ZN(n13490) );
  NAND2_X1 U15737 ( .A1(n13933), .A2(n6440), .ZN(n13465) );
  NAND2_X1 U15738 ( .A1(n13591), .A2(n13492), .ZN(n13464) );
  NAND2_X1 U15739 ( .A1(n13465), .A2(n13464), .ZN(n13489) );
  NOR2_X1 U15740 ( .A1(n13466), .A2(n13492), .ZN(n13467) );
  AOI21_X1 U15741 ( .B1(n13940), .B2(n13492), .A(n13467), .ZN(n13487) );
  NAND2_X1 U15742 ( .A1(n13940), .A2(n6440), .ZN(n13469) );
  NAND2_X1 U15743 ( .A1(n13720), .A2(n13492), .ZN(n13468) );
  NAND2_X1 U15744 ( .A1(n13469), .A2(n13468), .ZN(n13486) );
  AND2_X1 U15745 ( .A1(n13592), .A2(n6440), .ZN(n13470) );
  AOI21_X1 U15746 ( .B1(n13722), .B2(n13492), .A(n13470), .ZN(n13523) );
  NAND2_X1 U15747 ( .A1(n13722), .A2(n6440), .ZN(n13472) );
  NAND2_X1 U15748 ( .A1(n13592), .A2(n13492), .ZN(n13471) );
  NAND2_X1 U15749 ( .A1(n13472), .A2(n13471), .ZN(n13522) );
  AND2_X1 U15750 ( .A1(n13523), .A2(n13522), .ZN(n13473) );
  NOR2_X1 U15751 ( .A1(n13475), .A2(n13474), .ZN(n13476) );
  AOI21_X1 U15752 ( .B1(n13948), .B2(n13474), .A(n13476), .ZN(n13518) );
  NAND2_X1 U15753 ( .A1(n13948), .A2(n6440), .ZN(n13478) );
  NAND2_X1 U15754 ( .A1(n13719), .A2(n13492), .ZN(n13477) );
  NAND2_X1 U15755 ( .A1(n13478), .A2(n13477), .ZN(n13517) );
  INV_X1 U15756 ( .A(n13479), .ZN(n13482) );
  INV_X1 U15757 ( .A(n13480), .ZN(n13481) );
  AOI22_X1 U15758 ( .A1(n13518), .A2(n13517), .B1(n13482), .B2(n13481), .ZN(
        n13483) );
  OR3_X1 U15759 ( .A1(n13491), .A2(n13490), .A3(n13489), .ZN(n13515) );
  MUX2_X1 U15760 ( .A(n13679), .B(n13492), .S(n13676), .Z(n13494) );
  NAND2_X1 U15761 ( .A1(n13679), .A2(n13492), .ZN(n13493) );
  NAND2_X1 U15762 ( .A1(n13494), .A2(n13493), .ZN(n13509) );
  NAND2_X1 U15763 ( .A1(n13496), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13497) );
  OAI211_X1 U15764 ( .C1(n13499), .C2(n7902), .A(n13580), .B(n13570), .ZN(
        n13500) );
  AOI21_X1 U15765 ( .B1(n13679), .B2(n6440), .A(n13500), .ZN(n13502) );
  INV_X1 U15766 ( .A(n13588), .ZN(n13501) );
  NOR2_X1 U15767 ( .A1(n13502), .A2(n13501), .ZN(n13503) );
  AOI21_X1 U15768 ( .B1(n13675), .B2(n13492), .A(n13503), .ZN(n13529) );
  NAND2_X1 U15769 ( .A1(n13675), .A2(n6440), .ZN(n13505) );
  NAND2_X1 U15770 ( .A1(n13588), .A2(n13492), .ZN(n13504) );
  NAND2_X1 U15771 ( .A1(n13505), .A2(n13504), .ZN(n13528) );
  OAI22_X1 U15772 ( .A1(n13529), .A2(n13528), .B1(n13507), .B2(n13506), .ZN(
        n13508) );
  NAND2_X1 U15773 ( .A1(n13509), .A2(n13508), .ZN(n13514) );
  NAND4_X1 U15774 ( .A1(n7161), .A2(n13512), .A3(n13511), .A4(n13510), .ZN(
        n13513) );
  AND4_X1 U15775 ( .A1(n13516), .A2(n13515), .A3(n13514), .A4(n13513), .ZN(
        n13527) );
  INV_X1 U15776 ( .A(n13517), .ZN(n13520) );
  INV_X1 U15777 ( .A(n13518), .ZN(n13519) );
  NAND3_X1 U15778 ( .A1(n13521), .A2(n13520), .A3(n13519), .ZN(n13526) );
  OR3_X1 U15779 ( .A1(n13676), .A2(n13530), .A3(n6440), .ZN(n13532) );
  NAND3_X1 U15780 ( .A1(n13676), .A2(n13530), .A3(n6440), .ZN(n13531) );
  AND2_X1 U15781 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  XNOR2_X1 U15782 ( .A(n13675), .B(n13588), .ZN(n13563) );
  INV_X1 U15783 ( .A(n13534), .ZN(n13536) );
  NAND2_X1 U15784 ( .A1(n13538), .A2(n13537), .ZN(n13704) );
  AND4_X1 U15785 ( .A1(n13541), .A2(n13540), .A3(n7902), .A4(n13539), .ZN(
        n13544) );
  AND4_X1 U15786 ( .A1(n13545), .A2(n13544), .A3(n13543), .A4(n13542), .ZN(
        n13548) );
  NAND4_X1 U15787 ( .A1(n13549), .A2(n13548), .A3(n13547), .A4(n13546), .ZN(
        n13550) );
  OR3_X1 U15788 ( .A1(n13551), .A2(n8657), .A3(n13550), .ZN(n13554) );
  XNOR2_X1 U15789 ( .A(n14014), .B(n13552), .ZN(n13907) );
  NOR2_X1 U15790 ( .A1(n13889), .A2(n13555), .ZN(n13556) );
  XNOR2_X1 U15791 ( .A(n13996), .B(n13598), .ZN(n13858) );
  INV_X1 U15792 ( .A(n13718), .ZN(n13559) );
  NAND4_X1 U15793 ( .A1(n13563), .A2(n7973), .A3(n13562), .A4(n8503), .ZN(
        n13564) );
  NOR3_X1 U15794 ( .A1(n13566), .A2(n13565), .A3(n13564), .ZN(n13567) );
  INV_X1 U15795 ( .A(n13583), .ZN(n13573) );
  NAND2_X1 U15796 ( .A1(n13568), .A2(n13580), .ZN(n13569) );
  OAI211_X1 U15797 ( .C1(n13579), .C2(n13571), .A(n13570), .B(n13569), .ZN(
        n13572) );
  NAND3_X1 U15798 ( .A1(n13573), .A2(n13582), .A3(n13572), .ZN(n13586) );
  NAND4_X1 U15799 ( .A1(n15507), .A2(n13575), .A3(n13878), .A4(n13574), .ZN(
        n13576) );
  OAI211_X1 U15800 ( .C1(n13579), .C2(n13577), .A(n13576), .B(P2_B_REG_SCAN_IN), .ZN(n13585) );
  MUX2_X1 U15801 ( .A(n13580), .B(n13579), .S(n13578), .Z(n13581) );
  NAND4_X1 U15802 ( .A1(n13583), .A2(n13672), .A3(n13582), .A4(n13581), .ZN(
        n13584) );
  NAND4_X1 U15803 ( .A1(n13587), .A2(n13586), .A3(n13585), .A4(n13584), .ZN(
        P2_U3328) );
  MUX2_X1 U15804 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n13679), .S(n13611), .Z(
        P2_U3562) );
  MUX2_X1 U15805 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13588), .S(P2_U3947), .Z(
        P2_U3561) );
  MUX2_X1 U15806 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13589), .S(P2_U3947), .Z(
        P2_U3560) );
  MUX2_X1 U15807 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13590), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15808 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13591), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15809 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13720), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15810 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13592), .S(P2_U3947), .Z(
        P2_U3556) );
  MUX2_X1 U15811 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13719), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15812 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13593), .S(P2_U3947), .Z(
        P2_U3554) );
  MUX2_X1 U15813 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13594), .S(n13611), .Z(
        P2_U3553) );
  MUX2_X1 U15814 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13783), .S(n13611), .Z(
        P2_U3552) );
  MUX2_X1 U15815 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13595), .S(n13611), .Z(
        P2_U3551) );
  CLKBUF_X2 U15816 ( .A(P2_U3947), .Z(n13611) );
  MUX2_X1 U15817 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13782), .S(n13611), .Z(
        P2_U3550) );
  MUX2_X1 U15818 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13596), .S(n13611), .Z(
        P2_U3549) );
  MUX2_X1 U15819 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13597), .S(n13611), .Z(
        P2_U3548) );
  MUX2_X1 U15820 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13598), .S(n13611), .Z(
        P2_U3547) );
  MUX2_X1 U15821 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13881), .S(n13611), .Z(
        P2_U3546) );
  MUX2_X1 U15822 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13599), .S(n13611), .Z(
        P2_U3545) );
  MUX2_X1 U15823 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13879), .S(n13611), .Z(
        P2_U3544) );
  MUX2_X1 U15824 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13600), .S(n13611), .Z(
        P2_U3543) );
  MUX2_X1 U15825 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13601), .S(n13611), .Z(
        P2_U3542) );
  MUX2_X1 U15826 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13602), .S(n13611), .Z(
        P2_U3541) );
  MUX2_X1 U15827 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13603), .S(n13611), .Z(
        P2_U3540) );
  MUX2_X1 U15828 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13604), .S(n13611), .Z(
        P2_U3539) );
  MUX2_X1 U15829 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13605), .S(n13611), .Z(
        P2_U3538) );
  MUX2_X1 U15830 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13606), .S(n13611), .Z(
        P2_U3537) );
  MUX2_X1 U15831 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13607), .S(n13611), .Z(
        P2_U3536) );
  MUX2_X1 U15832 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13608), .S(n13611), .Z(
        P2_U3535) );
  MUX2_X1 U15833 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13609), .S(n13611), .Z(
        P2_U3534) );
  MUX2_X1 U15834 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13610), .S(n13611), .Z(
        P2_U3533) );
  MUX2_X1 U15835 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n13612), .S(n13611), .Z(
        P2_U3531) );
  NAND2_X1 U15836 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n13613) );
  OAI21_X1 U15837 ( .B1(n15500), .B2(n8759), .A(n13613), .ZN(n13614) );
  AOI21_X1 U15838 ( .B1(n13615), .B2(n7441), .A(n13614), .ZN(n13624) );
  OAI211_X1 U15839 ( .C1(n13618), .C2(n13617), .A(n15486), .B(n13616), .ZN(
        n13623) );
  OAI211_X1 U15840 ( .C1(n13621), .C2(n13620), .A(n15460), .B(n13619), .ZN(
        n13622) );
  NAND3_X1 U15841 ( .A1(n13624), .A2(n13623), .A3(n13622), .ZN(P2_U3220) );
  NAND2_X1 U15842 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3088), .ZN(n13625) );
  OAI21_X1 U15843 ( .B1(n15500), .B2(n13626), .A(n13625), .ZN(n13627) );
  AOI21_X1 U15844 ( .B1(n13628), .B2(n7441), .A(n13627), .ZN(n13637) );
  OAI211_X1 U15845 ( .C1(n13631), .C2(n13630), .A(n15460), .B(n13629), .ZN(
        n13636) );
  OAI211_X1 U15846 ( .C1(n13634), .C2(n13633), .A(n15486), .B(n13632), .ZN(
        n13635) );
  NAND3_X1 U15847 ( .A1(n13637), .A2(n13636), .A3(n13635), .ZN(P2_U3221) );
  NAND2_X1 U15848 ( .A1(n13638), .A2(n13649), .ZN(n13639) );
  NAND2_X1 U15849 ( .A1(n13640), .A2(n13639), .ZN(n13641) );
  XNOR2_X1 U15850 ( .A(n13641), .B(n15467), .ZN(n15464) );
  NAND2_X1 U15851 ( .A1(n15464), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n15463) );
  NAND2_X1 U15852 ( .A1(n13641), .A2(n13652), .ZN(n13642) );
  NAND2_X1 U15853 ( .A1(n15463), .A2(n13642), .ZN(n15475) );
  XNOR2_X1 U15854 ( .A(n13643), .B(P2_REG2_REG_16__SCAN_IN), .ZN(n15474) );
  NAND2_X1 U15855 ( .A1(n15475), .A2(n15474), .ZN(n15473) );
  NAND2_X1 U15856 ( .A1(n15482), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n13644) );
  NAND2_X1 U15857 ( .A1(n15473), .A2(n13644), .ZN(n15489) );
  INV_X1 U15858 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13845) );
  XNOR2_X1 U15859 ( .A(n15497), .B(n13845), .ZN(n15488) );
  NAND2_X1 U15860 ( .A1(n15489), .A2(n15488), .ZN(n15487) );
  NAND2_X1 U15861 ( .A1(n15497), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n13645) );
  NAND2_X1 U15862 ( .A1(n15487), .A2(n13645), .ZN(n13664) );
  XNOR2_X1 U15863 ( .A(n13664), .B(n13653), .ZN(n13662) );
  XOR2_X1 U15864 ( .A(n8354), .B(n13662), .Z(n13658) );
  INV_X1 U15865 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n13647) );
  OAI21_X1 U15866 ( .B1(n15500), .B2(n13647), .A(n13646), .ZN(n13656) );
  INV_X1 U15867 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n13987) );
  INV_X1 U15868 ( .A(n13650), .ZN(n13651) );
  XNOR2_X1 U15869 ( .A(n15482), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n15478) );
  XNOR2_X1 U15870 ( .A(n15497), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n15493) );
  AOI211_X1 U15871 ( .C1(n13987), .C2(n13654), .A(n15492), .B(n13659), .ZN(
        n13655) );
  AOI211_X1 U15872 ( .C1(n7441), .C2(n13663), .A(n13656), .B(n13655), .ZN(
        n13657) );
  OAI21_X1 U15873 ( .B1(n15448), .B2(n13658), .A(n13657), .ZN(P2_U3232) );
  NOR2_X1 U15874 ( .A1(n13660), .A2(n13659), .ZN(n13661) );
  XNOR2_X1 U15875 ( .A(n13661), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n13670) );
  NAND2_X1 U15876 ( .A1(n13662), .A2(n8354), .ZN(n13666) );
  OR2_X1 U15877 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  NAND2_X1 U15878 ( .A1(n13666), .A2(n13665), .ZN(n13668) );
  XNOR2_X1 U15879 ( .A(n13668), .B(n13667), .ZN(n13671) );
  INV_X1 U15880 ( .A(n13671), .ZN(n13669) );
  AOI22_X1 U15881 ( .A1(n13670), .A2(n15460), .B1(n15486), .B2(n13669), .ZN(
        n13673) );
  XNOR2_X1 U15882 ( .A(n13682), .B(n14043), .ZN(n13677) );
  NAND2_X1 U15883 ( .A1(n13677), .A2(n6405), .ZN(n13925) );
  NAND2_X1 U15884 ( .A1(n13679), .A2(n13678), .ZN(n13927) );
  NOR2_X1 U15885 ( .A1(n13797), .A2(n13927), .ZN(n13685) );
  NOR2_X1 U15886 ( .A1(n14043), .A2(n13904), .ZN(n13680) );
  AOI211_X1 U15887 ( .C1(n13797), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13685), 
        .B(n13680), .ZN(n13681) );
  OAI21_X1 U15888 ( .B1(n13925), .B2(n13744), .A(n13681), .ZN(P2_U3234) );
  OAI211_X1 U15889 ( .C1(n13683), .C2(n14047), .A(n6406), .B(n13682), .ZN(
        n13928) );
  NOR2_X1 U15890 ( .A1(n14047), .A2(n13904), .ZN(n13684) );
  AOI211_X1 U15891 ( .C1(n13894), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13685), 
        .B(n13684), .ZN(n13686) );
  OAI21_X1 U15892 ( .B1(n13928), .B2(n13744), .A(n13686), .ZN(P2_U3235) );
  XNOR2_X1 U15893 ( .A(n13687), .B(n13697), .ZN(n13689) );
  OAI21_X1 U15894 ( .B1(n13689), .B2(n13836), .A(n13688), .ZN(n13690) );
  INV_X1 U15895 ( .A(n13690), .ZN(n13936) );
  INV_X1 U15896 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n13691) );
  OAI22_X1 U15897 ( .A1(n13692), .A2(n13843), .B1(n13691), .B2(n13913), .ZN(
        n13696) );
  OAI211_X1 U15898 ( .C1(n13694), .C2(n13707), .A(n13693), .B(n6405), .ZN(
        n13935) );
  NOR2_X1 U15899 ( .A1(n13935), .A2(n13744), .ZN(n13695) );
  AOI211_X1 U15900 ( .C1(n13917), .C2(n13933), .A(n13696), .B(n13695), .ZN(
        n13701) );
  NAND3_X1 U15901 ( .A1(n13932), .A2(n13699), .A3(n13826), .ZN(n13700) );
  OAI211_X1 U15902 ( .C1(n13936), .C2(n13894), .A(n13701), .B(n13700), .ZN(
        P2_U3238) );
  XNOR2_X1 U15903 ( .A(n13702), .B(n13704), .ZN(n13941) );
  XNOR2_X1 U15904 ( .A(n13703), .B(n13704), .ZN(n13706) );
  OAI21_X1 U15905 ( .B1(n13706), .B2(n13836), .A(n13705), .ZN(n13938) );
  OAI21_X1 U15906 ( .B1(n13725), .B2(n13712), .A(n6406), .ZN(n13708) );
  NOR2_X1 U15907 ( .A1(n13708), .A2(n13707), .ZN(n13939) );
  NAND2_X1 U15908 ( .A1(n13939), .A2(n13919), .ZN(n13711) );
  AOI22_X1 U15909 ( .A1(n13709), .A2(n13915), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n13797), .ZN(n13710) );
  OAI211_X1 U15910 ( .C1(n13712), .C2(n13904), .A(n13711), .B(n13710), .ZN(
        n13713) );
  AOI21_X1 U15911 ( .B1(n13938), .B2(n13913), .A(n13713), .ZN(n13714) );
  OAI21_X1 U15912 ( .B1(n13908), .B2(n13941), .A(n13714), .ZN(P2_U3239) );
  XNOR2_X1 U15913 ( .A(n13715), .B(n13718), .ZN(n13944) );
  INV_X1 U15914 ( .A(n13944), .ZN(n13731) );
  INV_X1 U15915 ( .A(n13721), .ZN(n13942) );
  NAND2_X1 U15916 ( .A1(n13742), .A2(n13722), .ZN(n13723) );
  NAND2_X1 U15917 ( .A1(n13723), .A2(n6405), .ZN(n13724) );
  NOR2_X1 U15918 ( .A1(n13725), .A2(n13724), .ZN(n13943) );
  NAND2_X1 U15919 ( .A1(n13943), .A2(n13919), .ZN(n13728) );
  AOI22_X1 U15920 ( .A1(n13726), .A2(n13915), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n13797), .ZN(n13727) );
  OAI211_X1 U15921 ( .C1(n14053), .C2(n13904), .A(n13728), .B(n13727), .ZN(
        n13729) );
  AOI21_X1 U15922 ( .B1(n13942), .B2(n13913), .A(n13729), .ZN(n13730) );
  OAI21_X1 U15923 ( .B1(n13908), .B2(n13731), .A(n13730), .ZN(P2_U3240) );
  NAND2_X1 U15924 ( .A1(n13732), .A2(n8503), .ZN(n13733) );
  NAND2_X1 U15925 ( .A1(n13734), .A2(n13733), .ZN(n13947) );
  XNOR2_X1 U15926 ( .A(n13735), .B(n13736), .ZN(n13737) );
  NAND2_X1 U15927 ( .A1(n13737), .A2(n13897), .ZN(n13739) );
  NAND2_X1 U15928 ( .A1(n13739), .A2(n13738), .ZN(n13952) );
  NAND2_X1 U15929 ( .A1(n13952), .A2(n13913), .ZN(n13748) );
  INV_X1 U15930 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13740) );
  OAI22_X1 U15931 ( .A1(n13741), .A2(n13843), .B1(n13740), .B2(n13913), .ZN(
        n13746) );
  AOI21_X1 U15932 ( .B1(n13754), .B2(n13948), .A(n6409), .ZN(n13743) );
  NAND2_X1 U15933 ( .A1(n13743), .A2(n13742), .ZN(n13950) );
  NOR2_X1 U15934 ( .A1(n13950), .A2(n13744), .ZN(n13745) );
  AOI211_X1 U15935 ( .C1(n13917), .C2(n13948), .A(n13746), .B(n13745), .ZN(
        n13747) );
  OAI211_X1 U15936 ( .C1(n13908), .C2(n13947), .A(n13748), .B(n13747), .ZN(
        P2_U3241) );
  XOR2_X1 U15937 ( .A(n13760), .B(n13749), .Z(n13751) );
  OAI21_X1 U15938 ( .B1(n13751), .B2(n13836), .A(n13750), .ZN(n13954) );
  AOI21_X1 U15939 ( .B1(n13752), .B2(n13915), .A(n13954), .ZN(n13764) );
  INV_X1 U15940 ( .A(n13753), .ZN(n13756) );
  INV_X1 U15941 ( .A(n13754), .ZN(n13755) );
  AOI211_X1 U15942 ( .C1(n13956), .C2(n13756), .A(n6409), .B(n13755), .ZN(
        n13955) );
  INV_X1 U15943 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13757) );
  OAI22_X1 U15944 ( .A1(n13758), .A2(n13904), .B1(n13757), .B2(n13913), .ZN(
        n13762) );
  XNOR2_X1 U15945 ( .A(n13759), .B(n13760), .ZN(n13958) );
  NOR2_X1 U15946 ( .A1(n13958), .A2(n13908), .ZN(n13761) );
  AOI211_X1 U15947 ( .C1(n13955), .C2(n13919), .A(n13762), .B(n13761), .ZN(
        n13763) );
  OAI21_X1 U15948 ( .B1(n13764), .B2(n13894), .A(n13763), .ZN(P2_U3242) );
  XNOR2_X1 U15949 ( .A(n13765), .B(n13766), .ZN(n13968) );
  INV_X1 U15950 ( .A(n13968), .ZN(n13777) );
  XNOR2_X1 U15951 ( .A(n13767), .B(n8677), .ZN(n13769) );
  OAI21_X1 U15952 ( .B1(n13769), .B2(n13836), .A(n13768), .ZN(n13966) );
  OAI21_X1 U15953 ( .B1(n13787), .B2(n6876), .A(n6406), .ZN(n13771) );
  NOR2_X1 U15954 ( .A1(n13771), .A2(n13770), .ZN(n13967) );
  NAND2_X1 U15955 ( .A1(n13967), .A2(n13919), .ZN(n13774) );
  AOI22_X1 U15956 ( .A1(n13772), .A2(n13915), .B1(P2_REG2_REG_21__SCAN_IN), 
        .B2(n13797), .ZN(n13773) );
  OAI211_X1 U15957 ( .C1(n6876), .C2(n13904), .A(n13774), .B(n13773), .ZN(
        n13775) );
  AOI21_X1 U15958 ( .B1(n13966), .B2(n13913), .A(n13775), .ZN(n13776) );
  OAI21_X1 U15959 ( .B1(n13908), .B2(n13777), .A(n13776), .ZN(P2_U3244) );
  XNOR2_X1 U15960 ( .A(n13778), .B(n13781), .ZN(n13975) );
  OAI21_X1 U15961 ( .B1(n13781), .B2(n13780), .A(n13779), .ZN(n13784) );
  AOI222_X1 U15962 ( .A1(n13897), .A2(n13784), .B1(n13783), .B2(n13880), .C1(
        n13782), .C2(n13878), .ZN(n13974) );
  INV_X1 U15963 ( .A(n13974), .ZN(n13793) );
  NAND2_X1 U15964 ( .A1(n6527), .A2(n13972), .ZN(n13785) );
  NAND2_X1 U15965 ( .A1(n13785), .A2(n6405), .ZN(n13786) );
  NOR2_X1 U15966 ( .A1(n13787), .A2(n13786), .ZN(n13971) );
  NAND2_X1 U15967 ( .A1(n13971), .A2(n13919), .ZN(n13790) );
  AOI22_X1 U15968 ( .A1(n13788), .A2(n13915), .B1(P2_REG2_REG_20__SCAN_IN), 
        .B2(n13797), .ZN(n13789) );
  OAI211_X1 U15969 ( .C1(n13791), .C2(n13904), .A(n13790), .B(n13789), .ZN(
        n13792) );
  AOI21_X1 U15970 ( .B1(n13793), .B2(n13913), .A(n13792), .ZN(n13794) );
  OAI21_X1 U15971 ( .B1(n13908), .B2(n13975), .A(n13794), .ZN(P2_U3245) );
  XNOR2_X1 U15972 ( .A(n13795), .B(n8403), .ZN(n13980) );
  AOI21_X1 U15973 ( .B1(n13820), .B2(n14065), .A(n6409), .ZN(n13796) );
  NAND2_X1 U15974 ( .A1(n13796), .A2(n6527), .ZN(n13977) );
  INV_X1 U15975 ( .A(n13977), .ZN(n13807) );
  AOI22_X1 U15976 ( .A1(n13798), .A2(n13915), .B1(P2_REG2_REG_19__SCAN_IN), 
        .B2(n13797), .ZN(n13799) );
  OAI21_X1 U15977 ( .B1(n6879), .B2(n13904), .A(n13799), .ZN(n13806) );
  NAND2_X1 U15978 ( .A1(n13800), .A2(n13801), .ZN(n13802) );
  NAND2_X1 U15979 ( .A1(n13803), .A2(n13802), .ZN(n13804) );
  NAND2_X1 U15980 ( .A1(n13804), .A2(n13897), .ZN(n13979) );
  AOI21_X1 U15981 ( .B1(n13979), .B2(n13976), .A(n13894), .ZN(n13805) );
  AOI211_X1 U15982 ( .C1(n13807), .C2(n13919), .A(n13806), .B(n13805), .ZN(
        n13808) );
  OAI21_X1 U15983 ( .B1(n13908), .B2(n13980), .A(n13808), .ZN(P2_U3246) );
  NAND2_X1 U15984 ( .A1(n13870), .A2(n13869), .ZN(n13868) );
  INV_X1 U15985 ( .A(n13809), .ZN(n13810) );
  NAND2_X1 U15986 ( .A1(n13868), .A2(n13810), .ZN(n13851) );
  AOI21_X1 U15987 ( .B1(n13851), .B2(n13811), .A(n7970), .ZN(n13834) );
  AND2_X1 U15988 ( .A1(n13834), .A2(n13833), .ZN(n13835) );
  NOR2_X1 U15989 ( .A1(n13835), .A2(n13812), .ZN(n13813) );
  XOR2_X1 U15990 ( .A(n13817), .B(n13813), .Z(n13815) );
  OAI21_X1 U15991 ( .B1(n13815), .B2(n13836), .A(n13814), .ZN(n13984) );
  INV_X1 U15992 ( .A(n13984), .ZN(n13828) );
  INV_X1 U15993 ( .A(n13816), .ZN(n13819) );
  INV_X1 U15994 ( .A(n13817), .ZN(n13818) );
  OAI21_X1 U15995 ( .B1(n13819), .B2(n13818), .A(n6510), .ZN(n13986) );
  AOI211_X1 U15996 ( .C1(n13821), .C2(n13841), .A(n6409), .B(n6875), .ZN(
        n13985) );
  NAND2_X1 U15997 ( .A1(n13985), .A2(n13919), .ZN(n13824) );
  AOI22_X1 U15998 ( .A1(n13894), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13822), 
        .B2(n13915), .ZN(n13823) );
  OAI211_X1 U15999 ( .C1(n14070), .C2(n13904), .A(n13824), .B(n13823), .ZN(
        n13825) );
  AOI21_X1 U16000 ( .B1(n13826), .B2(n13986), .A(n13825), .ZN(n13827) );
  OAI21_X1 U16001 ( .B1(n13828), .B2(n13894), .A(n13827), .ZN(P2_U3247) );
  INV_X1 U16002 ( .A(n13830), .ZN(n13831) );
  NAND2_X1 U16003 ( .A1(n13860), .A2(n13831), .ZN(n13832) );
  XNOR2_X1 U16004 ( .A(n13832), .B(n13833), .ZN(n13989) );
  INV_X1 U16005 ( .A(n13989), .ZN(n13850) );
  NOR2_X1 U16006 ( .A1(n13834), .A2(n13833), .ZN(n13837) );
  OR3_X1 U16007 ( .A1(n13837), .A2(n13836), .A3(n13835), .ZN(n13839) );
  NAND2_X1 U16008 ( .A1(n13839), .A2(n13838), .ZN(n13992) );
  NAND2_X1 U16009 ( .A1(n13992), .A2(n13913), .ZN(n13849) );
  OR2_X1 U16010 ( .A1(n6463), .A2(n13842), .ZN(n13840) );
  AND3_X1 U16011 ( .A1(n13841), .A2(n13840), .A3(n6406), .ZN(n13990) );
  NOR2_X1 U16012 ( .A1(n13842), .A2(n13904), .ZN(n13847) );
  OAI22_X1 U16013 ( .A1(n13913), .A2(n13845), .B1(n13844), .B2(n13843), .ZN(
        n13846) );
  AOI211_X1 U16014 ( .C1(n13990), .C2(n13919), .A(n13847), .B(n13846), .ZN(
        n13848) );
  OAI211_X1 U16015 ( .C1(n13908), .C2(n13850), .A(n13849), .B(n13848), .ZN(
        P2_U3248) );
  XNOR2_X1 U16016 ( .A(n13851), .B(n13858), .ZN(n13853) );
  AOI21_X1 U16017 ( .B1(n13853), .B2(n13897), .A(n13852), .ZN(n13998) );
  AOI211_X1 U16018 ( .C1(n13996), .C2(n7760), .A(n6409), .B(n6463), .ZN(n13995) );
  INV_X1 U16019 ( .A(n13854), .ZN(n13855) );
  AOI22_X1 U16020 ( .A1(n13894), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n13855), 
        .B2(n13915), .ZN(n13856) );
  OAI21_X1 U16021 ( .B1(n13857), .B2(n13904), .A(n13856), .ZN(n13862) );
  NAND2_X1 U16022 ( .A1(n13829), .A2(n13858), .ZN(n13859) );
  NAND2_X1 U16023 ( .A1(n13860), .A2(n13859), .ZN(n13999) );
  NOR2_X1 U16024 ( .A1(n13999), .A2(n13908), .ZN(n13861) );
  AOI211_X1 U16025 ( .C1(n13995), .C2(n13919), .A(n13862), .B(n13861), .ZN(
        n13863) );
  OAI21_X1 U16026 ( .B1(n13998), .B2(n13894), .A(n13863), .ZN(P2_U3249) );
  XOR2_X1 U16027 ( .A(n13869), .B(n13864), .Z(n14000) );
  AOI211_X1 U16028 ( .C1(n13866), .C2(n13884), .A(n6409), .B(n13865), .ZN(
        n14002) );
  INV_X1 U16029 ( .A(n13866), .ZN(n14080) );
  INV_X1 U16030 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n13867) );
  OAI22_X1 U16031 ( .A1(n14080), .A2(n13904), .B1(n13867), .B2(n13913), .ZN(
        n13875) );
  OAI21_X1 U16032 ( .B1(n13870), .B2(n13869), .A(n13868), .ZN(n13871) );
  AND2_X1 U16033 ( .A1(n13871), .A2(n13897), .ZN(n14004) );
  AOI211_X1 U16034 ( .C1(n13915), .C2(n13872), .A(n14001), .B(n14004), .ZN(
        n13873) );
  NOR2_X1 U16035 ( .A1(n13873), .A2(n13894), .ZN(n13874) );
  AOI211_X1 U16036 ( .C1(n14002), .C2(n13919), .A(n13875), .B(n13874), .ZN(
        n13876) );
  OAI21_X1 U16037 ( .B1(n13908), .B2(n14000), .A(n13876), .ZN(P2_U3250) );
  XNOR2_X1 U16038 ( .A(n13877), .B(n13889), .ZN(n13882) );
  AOI222_X1 U16039 ( .A1(n13897), .A2(n13882), .B1(n13881), .B2(n13880), .C1(
        n13879), .C2(n13878), .ZN(n14011) );
  INV_X1 U16040 ( .A(n13884), .ZN(n13885) );
  AOI211_X1 U16041 ( .C1(n14009), .C2(n13899), .A(n6409), .B(n13885), .ZN(
        n14008) );
  INV_X1 U16042 ( .A(n13886), .ZN(n13887) );
  AOI22_X1 U16043 ( .A1(n13894), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n13887), 
        .B2(n13915), .ZN(n13888) );
  OAI21_X1 U16044 ( .B1(n8688), .B2(n13904), .A(n13888), .ZN(n13892) );
  XNOR2_X1 U16045 ( .A(n13890), .B(n13889), .ZN(n14012) );
  NOR2_X1 U16046 ( .A1(n14012), .A2(n13908), .ZN(n13891) );
  AOI211_X1 U16047 ( .C1(n14008), .C2(n13919), .A(n13892), .B(n13891), .ZN(
        n13893) );
  OAI21_X1 U16048 ( .B1(n14011), .B2(n13894), .A(n13893), .ZN(P2_U3251) );
  XNOR2_X1 U16049 ( .A(n13895), .B(n13907), .ZN(n13898) );
  AOI21_X1 U16050 ( .B1(n13898), .B2(n13897), .A(n13896), .ZN(n14016) );
  AOI211_X1 U16051 ( .C1(n14014), .C2(n13900), .A(n6409), .B(n13883), .ZN(
        n14013) );
  INV_X1 U16052 ( .A(n13901), .ZN(n13902) );
  AOI22_X1 U16053 ( .A1(n13797), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n13902), 
        .B2(n13915), .ZN(n13903) );
  OAI21_X1 U16054 ( .B1(n13905), .B2(n13904), .A(n13903), .ZN(n13910) );
  XOR2_X1 U16055 ( .A(n13906), .B(n13907), .Z(n14017) );
  NOR2_X1 U16056 ( .A1(n14017), .A2(n13908), .ZN(n13909) );
  AOI211_X1 U16057 ( .C1(n14013), .C2(n13919), .A(n13910), .B(n13909), .ZN(
        n13911) );
  OAI21_X1 U16058 ( .B1(n13797), .B2(n14016), .A(n13911), .ZN(P2_U3252) );
  INV_X1 U16059 ( .A(n13912), .ZN(n13914) );
  MUX2_X1 U16060 ( .A(n15797), .B(n13914), .S(n13913), .Z(n13924) );
  AOI22_X1 U16061 ( .A1(n13917), .A2(n13916), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n13915), .ZN(n13923) );
  AOI22_X1 U16062 ( .A1(n13921), .A2(n13920), .B1(n13919), .B2(n13918), .ZN(
        n13922) );
  NAND3_X1 U16063 ( .A1(n13924), .A2(n13923), .A3(n13922), .ZN(P2_U3264) );
  OAI21_X1 U16064 ( .B1(n14043), .B2(n14007), .A(n13926), .ZN(P2_U3530) );
  AND2_X1 U16065 ( .A1(n13928), .A2(n13927), .ZN(n14044) );
  MUX2_X1 U16066 ( .A(n13929), .B(n14044), .S(n15538), .Z(n13930) );
  OAI21_X1 U16067 ( .B1(n14047), .B2(n14007), .A(n13930), .ZN(P2_U3529) );
  NAND3_X1 U16068 ( .A1(n13932), .A2(n15522), .A3(n13699), .ZN(n13937) );
  NAND2_X1 U16069 ( .A1(n13933), .A2(n15524), .ZN(n13934) );
  NAND4_X1 U16070 ( .A1(n13937), .A2(n13936), .A3(n13935), .A4(n13934), .ZN(
        n14048) );
  MUX2_X1 U16071 ( .A(n14048), .B(P2_REG1_REG_27__SCAN_IN), .S(n15536), .Z(
        P2_U3526) );
  MUX2_X1 U16072 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14049), .S(n15538), .Z(
        P2_U3525) );
  OAI21_X1 U16073 ( .B1(n14053), .B2(n14007), .A(n13946), .ZN(P2_U3524) );
  NOR2_X1 U16074 ( .A1(n13947), .A2(n14040), .ZN(n13953) );
  NAND2_X1 U16075 ( .A1(n13948), .A2(n15524), .ZN(n13949) );
  NAND2_X1 U16076 ( .A1(n13950), .A2(n13949), .ZN(n13951) );
  OR3_X2 U16077 ( .A1(n13953), .A2(n13952), .A3(n13951), .ZN(n14054) );
  MUX2_X1 U16078 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14054), .S(n15538), .Z(
        P2_U3523) );
  AOI211_X1 U16079 ( .C1(n15524), .C2(n13956), .A(n13955), .B(n13954), .ZN(
        n13957) );
  OAI21_X1 U16080 ( .B1(n14040), .B2(n13958), .A(n13957), .ZN(n14055) );
  MUX2_X1 U16081 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14055), .S(n15538), .Z(
        P2_U3522) );
  NOR2_X1 U16082 ( .A1(n13959), .A2(n14040), .ZN(n13963) );
  INV_X1 U16083 ( .A(n13960), .ZN(n13962) );
  MUX2_X1 U16084 ( .A(n14056), .B(P2_REG1_REG_22__SCAN_IN), .S(n15536), .Z(
        n13964) );
  AOI21_X1 U16085 ( .B1(n14023), .B2(n14058), .A(n13964), .ZN(n13965) );
  INV_X1 U16086 ( .A(n13965), .ZN(P2_U3521) );
  INV_X1 U16087 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n13969) );
  AOI211_X1 U16088 ( .C1(n15522), .C2(n13968), .A(n13967), .B(n13966), .ZN(
        n14060) );
  MUX2_X1 U16089 ( .A(n13969), .B(n14060), .S(n15538), .Z(n13970) );
  OAI21_X1 U16090 ( .B1(n6876), .B2(n14007), .A(n13970), .ZN(P2_U3520) );
  AOI21_X1 U16091 ( .B1(n15524), .B2(n13972), .A(n13971), .ZN(n13973) );
  OAI211_X1 U16092 ( .C1(n14040), .C2(n13975), .A(n13974), .B(n13973), .ZN(
        n14062) );
  MUX2_X1 U16093 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14062), .S(n15538), .Z(
        P2_U3519) );
  AND2_X1 U16094 ( .A1(n13977), .A2(n13976), .ZN(n13978) );
  OAI211_X1 U16095 ( .C1(n14040), .C2(n13980), .A(n13979), .B(n13978), .ZN(
        n14063) );
  INV_X1 U16096 ( .A(n14063), .ZN(n13982) );
  INV_X1 U16097 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n13981) );
  MUX2_X1 U16098 ( .A(n13982), .B(n13981), .S(n15536), .Z(n13983) );
  OAI21_X1 U16099 ( .B1(n6879), .B2(n14007), .A(n13983), .ZN(P2_U3518) );
  AOI211_X1 U16100 ( .C1(n15522), .C2(n13986), .A(n13985), .B(n13984), .ZN(
        n14067) );
  MUX2_X1 U16101 ( .A(n13987), .B(n14067), .S(n15538), .Z(n13988) );
  OAI21_X1 U16102 ( .B1(n14070), .B2(n14007), .A(n13988), .ZN(P2_U3517) );
  AND2_X1 U16103 ( .A1(n13989), .A2(n15522), .ZN(n13991) );
  MUX2_X1 U16104 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14071), .S(n15538), .Z(
        n13993) );
  AOI21_X1 U16105 ( .B1(n14023), .B2(n14073), .A(n13993), .ZN(n13994) );
  INV_X1 U16106 ( .A(n13994), .ZN(P2_U3516) );
  AOI21_X1 U16107 ( .B1(n15524), .B2(n13996), .A(n13995), .ZN(n13997) );
  OAI211_X1 U16108 ( .C1(n14040), .C2(n13999), .A(n13998), .B(n13997), .ZN(
        n14075) );
  MUX2_X1 U16109 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n14075), .S(n15538), .Z(
        P2_U3515) );
  INV_X1 U16110 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14005) );
  NOR2_X1 U16111 ( .A1(n14000), .A2(n14040), .ZN(n14003) );
  NOR4_X1 U16112 ( .A1(n14004), .A2(n14003), .A3(n14002), .A4(n14001), .ZN(
        n14076) );
  MUX2_X1 U16113 ( .A(n14005), .B(n14076), .S(n15538), .Z(n14006) );
  OAI21_X1 U16114 ( .B1(n14080), .B2(n14007), .A(n14006), .ZN(P2_U3514) );
  AOI21_X1 U16115 ( .B1(n15524), .B2(n14009), .A(n14008), .ZN(n14010) );
  OAI211_X1 U16116 ( .C1(n14040), .C2(n14012), .A(n14011), .B(n14010), .ZN(
        n14081) );
  MUX2_X1 U16117 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n14081), .S(n15538), .Z(
        P2_U3513) );
  AOI21_X1 U16118 ( .B1(n15524), .B2(n14014), .A(n14013), .ZN(n14015) );
  OAI211_X1 U16119 ( .C1(n14040), .C2(n14017), .A(n14016), .B(n14015), .ZN(
        n14082) );
  MUX2_X1 U16120 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n14082), .S(n15538), .Z(
        P2_U3512) );
  AND2_X1 U16121 ( .A1(n14018), .A2(n15522), .ZN(n14020) );
  MUX2_X1 U16122 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14083), .S(n15538), .Z(
        n14022) );
  AOI21_X1 U16123 ( .B1(n14023), .B2(n14085), .A(n14022), .ZN(n14024) );
  INV_X1 U16124 ( .A(n14024), .ZN(P2_U3511) );
  AOI21_X1 U16125 ( .B1(n15524), .B2(n14026), .A(n14025), .ZN(n14027) );
  OAI211_X1 U16126 ( .C1(n13285), .C2(n14029), .A(n14028), .B(n14027), .ZN(
        n14088) );
  MUX2_X1 U16127 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n14088), .S(n15538), .Z(
        P2_U3509) );
  AOI21_X1 U16128 ( .B1(n15524), .B2(n14031), .A(n14030), .ZN(n14032) );
  OAI211_X1 U16129 ( .C1(n14040), .C2(n14034), .A(n14033), .B(n14032), .ZN(
        n14089) );
  MUX2_X1 U16130 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n14089), .S(n15538), .Z(
        P2_U3507) );
  AOI21_X1 U16131 ( .B1(n15524), .B2(n14036), .A(n14035), .ZN(n14037) );
  OAI211_X1 U16132 ( .C1(n14040), .C2(n14039), .A(n14038), .B(n14037), .ZN(
        n14090) );
  MUX2_X1 U16133 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n14090), .S(n15538), .Z(
        P2_U3505) );
  OAI21_X1 U16134 ( .B1(n14043), .B2(n14079), .A(n14042), .ZN(P2_U3498) );
  MUX2_X1 U16135 ( .A(n14045), .B(n14044), .S(n15533), .Z(n14046) );
  OAI21_X1 U16136 ( .B1(n14047), .B2(n14079), .A(n14046), .ZN(P2_U3497) );
  MUX2_X1 U16137 ( .A(n14048), .B(P2_REG0_REG_27__SCAN_IN), .S(n15531), .Z(
        P2_U3494) );
  MUX2_X1 U16138 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14049), .S(n15533), .Z(
        P2_U3493) );
  INV_X1 U16139 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n14051) );
  MUX2_X1 U16140 ( .A(n14051), .B(n14050), .S(n15533), .Z(n14052) );
  MUX2_X1 U16141 ( .A(n14054), .B(P2_REG0_REG_24__SCAN_IN), .S(n15531), .Z(
        P2_U3491) );
  MUX2_X1 U16142 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14055), .S(n15533), .Z(
        P2_U3490) );
  MUX2_X1 U16143 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n14056), .S(n15533), .Z(
        n14057) );
  AOI21_X1 U16144 ( .B1(n14086), .B2(n14058), .A(n14057), .ZN(n14059) );
  INV_X1 U16145 ( .A(n14059), .ZN(P2_U3489) );
  MUX2_X1 U16146 ( .A(n15733), .B(n14060), .S(n15533), .Z(n14061) );
  OAI21_X1 U16147 ( .B1(n6876), .B2(n14079), .A(n14061), .ZN(P2_U3488) );
  MUX2_X1 U16148 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14062), .S(n15533), .Z(
        P2_U3487) );
  MUX2_X1 U16149 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14063), .S(n15533), .Z(
        n14064) );
  AOI21_X1 U16150 ( .B1(n14086), .B2(n14065), .A(n14064), .ZN(n14066) );
  INV_X1 U16151 ( .A(n14066), .ZN(P2_U3486) );
  INV_X1 U16152 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n14068) );
  MUX2_X1 U16153 ( .A(n14068), .B(n14067), .S(n15533), .Z(n14069) );
  OAI21_X1 U16154 ( .B1(n14070), .B2(n14079), .A(n14069), .ZN(P2_U3484) );
  MUX2_X1 U16155 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n14071), .S(n15533), .Z(
        n14072) );
  AOI21_X1 U16156 ( .B1(n14086), .B2(n14073), .A(n14072), .ZN(n14074) );
  INV_X1 U16157 ( .A(n14074), .ZN(P2_U3481) );
  MUX2_X1 U16158 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n14075), .S(n15533), .Z(
        P2_U3478) );
  INV_X1 U16159 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14077) );
  MUX2_X1 U16160 ( .A(n14077), .B(n14076), .S(n15533), .Z(n14078) );
  OAI21_X1 U16161 ( .B1(n14080), .B2(n14079), .A(n14078), .ZN(P2_U3475) );
  MUX2_X1 U16162 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n14081), .S(n15533), .Z(
        P2_U3472) );
  MUX2_X1 U16163 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n14082), .S(n15533), .Z(
        P2_U3469) );
  MUX2_X1 U16164 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n14083), .S(n15533), .Z(
        n14084) );
  AOI21_X1 U16165 ( .B1(n14086), .B2(n14085), .A(n14084), .ZN(n14087) );
  INV_X1 U16166 ( .A(n14087), .ZN(P2_U3466) );
  MUX2_X1 U16167 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n14088), .S(n15533), .Z(
        P2_U3460) );
  MUX2_X1 U16168 ( .A(P2_REG0_REG_8__SCAN_IN), .B(n14089), .S(n15533), .Z(
        P2_U3454) );
  MUX2_X1 U16169 ( .A(P2_REG0_REG_6__SCAN_IN), .B(n14090), .S(n15533), .Z(
        P2_U3448) );
  INV_X1 U16170 ( .A(n14474), .ZN(n15188) );
  NOR4_X1 U16171 ( .A1(n14091), .A2(P2_IR_REG_30__SCAN_IN), .A3(n7989), .A4(
        P2_U3088), .ZN(n14092) );
  AOI21_X1 U16172 ( .B1(n14093), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n14092), 
        .ZN(n14094) );
  OAI21_X1 U16173 ( .B1(n15188), .B2(n14099), .A(n14094), .ZN(P2_U3296) );
  OAI222_X1 U16174 ( .A1(n14102), .A2(n14097), .B1(P2_U3088), .B2(n14096), 
        .C1(n14099), .C2(n14095), .ZN(P2_U3297) );
  INV_X1 U16175 ( .A(n14098), .ZN(n15191) );
  OAI222_X1 U16176 ( .A1(n14102), .A2(n14101), .B1(P2_U3088), .B2(n7993), .C1(
        n14099), .C2(n15191), .ZN(P2_U3298) );
  MUX2_X1 U16177 ( .A(n14103), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  XOR2_X1 U16178 ( .A(n14105), .B(n14104), .Z(n14106) );
  NAND2_X1 U16179 ( .A1(n14106), .A2(n14273), .ZN(n14114) );
  NAND2_X1 U16180 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n14633) );
  OAI21_X1 U16181 ( .B1(n14267), .B2(n14107), .A(n14633), .ZN(n14108) );
  INV_X1 U16182 ( .A(n14108), .ZN(n14113) );
  INV_X1 U16183 ( .A(n14109), .ZN(n14110) );
  AOI22_X1 U16184 ( .A1(n14264), .A2(n14553), .B1(n14262), .B2(n14110), .ZN(
        n14112) );
  NAND2_X1 U16185 ( .A1(n14269), .A2(n14325), .ZN(n14111) );
  NAND4_X1 U16186 ( .A1(n14114), .A2(n14113), .A3(n14112), .A4(n14111), .ZN(
        P1_U3213) );
  XNOR2_X1 U16187 ( .A(n14116), .B(n14115), .ZN(n14121) );
  AOI22_X1 U16188 ( .A1(n14753), .A2(n14264), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14118) );
  NAND2_X1 U16189 ( .A1(n14805), .A2(n14262), .ZN(n14117) );
  OAI211_X1 U16190 ( .C1(n14794), .C2(n14267), .A(n14118), .B(n14117), .ZN(
        n14119) );
  AOI21_X1 U16191 ( .B1(n14806), .B2(n14269), .A(n14119), .ZN(n14120) );
  OAI21_X1 U16192 ( .B1(n14121), .B2(n14271), .A(n14120), .ZN(P1_U3214) );
  INV_X1 U16193 ( .A(n14122), .ZN(n14123) );
  AOI21_X1 U16194 ( .B1(n14125), .B2(n14124), .A(n14123), .ZN(n14131) );
  OAI21_X1 U16195 ( .B1(n14267), .B2(n14370), .A(n14126), .ZN(n14129) );
  OAI22_X1 U16196 ( .A1(n14255), .A2(n14127), .B1(n14279), .B2(n15007), .ZN(
        n14128) );
  AOI211_X1 U16197 ( .C1(n15136), .C2(n14269), .A(n14129), .B(n14128), .ZN(
        n14130) );
  OAI21_X1 U16198 ( .B1(n14131), .B2(n14271), .A(n14130), .ZN(P1_U3215) );
  XOR2_X1 U16199 ( .A(n14133), .B(n14132), .Z(n14139) );
  INV_X1 U16200 ( .A(n14134), .ZN(n14857) );
  AOI22_X1 U16201 ( .A1(n14857), .A2(n14262), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14136) );
  NAND2_X1 U16202 ( .A1(n14543), .A2(n14264), .ZN(n14135) );
  OAI211_X1 U16203 ( .C1(n14854), .C2(n14267), .A(n14136), .B(n14135), .ZN(
        n14137) );
  AOI21_X1 U16204 ( .B1(n15078), .B2(n14269), .A(n14137), .ZN(n14138) );
  OAI21_X1 U16205 ( .B1(n14139), .B2(n14271), .A(n14138), .ZN(P1_U3216) );
  AND2_X1 U16206 ( .A1(n14141), .A2(n14140), .ZN(n14143) );
  OAI211_X1 U16207 ( .C1(n14144), .C2(n14143), .A(n14142), .B(n14273), .ZN(
        n14151) );
  AOI22_X1 U16208 ( .A1(n14264), .A2(n14557), .B1(n14262), .B2(n14145), .ZN(
        n14150) );
  OAI22_X1 U16209 ( .A1(n14267), .A2(n14146), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14145), .ZN(n14147) );
  AOI21_X1 U16210 ( .B1(n14269), .B2(n14148), .A(n14147), .ZN(n14149) );
  NAND3_X1 U16211 ( .A1(n14151), .A2(n14150), .A3(n14149), .ZN(P1_U3218) );
  OAI211_X1 U16212 ( .C1(n14154), .C2(n14153), .A(n14152), .B(n14273), .ZN(
        n14158) );
  OAI22_X1 U16213 ( .A1(n14405), .A2(n14855), .B1(n14155), .B2(n14853), .ZN(
        n15103) );
  NAND2_X1 U16214 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14740)
         );
  OAI21_X1 U16215 ( .B1(n14279), .B2(n14917), .A(n14740), .ZN(n14156) );
  AOI21_X1 U16216 ( .B1(n15103), .B2(n14282), .A(n14156), .ZN(n14157) );
  OAI211_X1 U16217 ( .C1(n14921), .C2(n14285), .A(n14158), .B(n14157), .ZN(
        P1_U3219) );
  NAND2_X1 U16218 ( .A1(n14161), .A2(n14160), .ZN(n14162) );
  AOI21_X1 U16219 ( .B1(n14159), .B2(n14162), .A(n14271), .ZN(n14167) );
  NAND2_X1 U16220 ( .A1(n14891), .A2(n15336), .ZN(n15092) );
  INV_X1 U16221 ( .A(n14218), .ZN(n14165) );
  AOI22_X1 U16222 ( .A1(n14890), .A2(n14262), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14164) );
  OAI22_X1 U16223 ( .A1(n14852), .A2(n14855), .B1(n14405), .B2(n14853), .ZN(
        n14881) );
  NAND2_X1 U16224 ( .A1(n14881), .A2(n14282), .ZN(n14163) );
  OAI211_X1 U16225 ( .C1(n15092), .C2(n14165), .A(n14164), .B(n14163), .ZN(
        n14166) );
  OR2_X1 U16226 ( .A1(n14167), .A2(n14166), .ZN(P1_U3223) );
  AOI21_X1 U16227 ( .B1(n14168), .B2(n14169), .A(n14271), .ZN(n14170) );
  OR2_X1 U16228 ( .A1(n14168), .A2(n14169), .ZN(n14230) );
  NAND2_X1 U16229 ( .A1(n14170), .A2(n14230), .ZN(n14176) );
  NOR2_X1 U16230 ( .A1(n14279), .A2(n14171), .ZN(n14172) );
  AOI211_X1 U16231 ( .C1(n14282), .C2(n14174), .A(n14173), .B(n14172), .ZN(
        n14175) );
  OAI211_X1 U16232 ( .C1(n14177), .C2(n14285), .A(n14176), .B(n14175), .ZN(
        P1_U3224) );
  XOR2_X1 U16233 ( .A(n14179), .B(n14178), .Z(n14186) );
  AND2_X1 U16234 ( .A1(n14542), .A2(n15008), .ZN(n14180) );
  AOI21_X1 U16235 ( .B1(n14753), .B2(n15010), .A(n14180), .ZN(n15066) );
  INV_X1 U16236 ( .A(n14181), .ZN(n14821) );
  AOI22_X1 U16237 ( .A1(n14821), .A2(n14262), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14182) );
  OAI21_X1 U16238 ( .B1(n15066), .B2(n14183), .A(n14182), .ZN(n14184) );
  AOI21_X1 U16239 ( .B1(n15065), .B2(n14269), .A(n14184), .ZN(n14185) );
  OAI21_X1 U16240 ( .B1(n14186), .B2(n14271), .A(n14185), .ZN(P1_U3225) );
  XNOR2_X1 U16241 ( .A(n14188), .B(n14187), .ZN(n14194) );
  INV_X1 U16242 ( .A(n14190), .ZN(n14192) );
  INV_X1 U16243 ( .A(n14189), .ZN(n14191) );
  XOR2_X1 U16244 ( .A(n14190), .B(n14189), .Z(n14276) );
  NAND2_X1 U16245 ( .A1(n14276), .A2(n14275), .ZN(n14274) );
  OAI21_X1 U16246 ( .B1(n14192), .B2(n14191), .A(n14274), .ZN(n14193) );
  NOR2_X1 U16247 ( .A1(n14193), .A2(n14194), .ZN(n14203) );
  AOI21_X1 U16248 ( .B1(n14194), .B2(n14193), .A(n14203), .ZN(n14199) );
  OAI21_X1 U16249 ( .B1(n14254), .B2(n14267), .A(n14195), .ZN(n14197) );
  OAI22_X1 U16250 ( .A1(n14255), .A2(n14370), .B1(n14279), .B2(n14978), .ZN(
        n14196) );
  AOI211_X1 U16251 ( .C1(n15122), .C2(n14269), .A(n14197), .B(n14196), .ZN(
        n14198) );
  OAI21_X1 U16252 ( .B1(n14199), .B2(n14271), .A(n14198), .ZN(P1_U3226) );
  INV_X1 U16253 ( .A(n14960), .ZN(n15116) );
  INV_X1 U16254 ( .A(n14200), .ZN(n14202) );
  NOR3_X1 U16255 ( .A1(n14203), .A2(n14202), .A3(n14201), .ZN(n14206) );
  INV_X1 U16256 ( .A(n14204), .ZN(n14205) );
  OAI21_X1 U16257 ( .B1(n14206), .B2(n14205), .A(n14273), .ZN(n14211) );
  NOR2_X1 U16258 ( .A1(n14207), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14693) );
  OAI22_X1 U16259 ( .A1(n14255), .A2(n14384), .B1(n14279), .B2(n14957), .ZN(
        n14208) );
  AOI211_X1 U16260 ( .C1(n14209), .C2(n14956), .A(n14693), .B(n14208), .ZN(
        n14210) );
  OAI211_X1 U16261 ( .C1(n15116), .C2(n14285), .A(n14211), .B(n14210), .ZN(
        P1_U3228) );
  XOR2_X1 U16262 ( .A(n14213), .B(n14212), .Z(n14220) );
  AOI22_X1 U16263 ( .A1(n14841), .A2(n14262), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14215) );
  NAND2_X1 U16264 ( .A1(n14832), .A2(n14264), .ZN(n14214) );
  OAI211_X1 U16265 ( .C1(n14216), .C2(n14267), .A(n14215), .B(n14214), .ZN(
        n14217) );
  AOI21_X1 U16266 ( .B1(n15073), .B2(n14218), .A(n14217), .ZN(n14219) );
  OAI21_X1 U16267 ( .B1(n14220), .B2(n14271), .A(n14219), .ZN(P1_U3229) );
  OAI211_X1 U16268 ( .C1(n14223), .C2(n14222), .A(n14221), .B(n14273), .ZN(
        n14228) );
  OAI22_X1 U16269 ( .A1(n14224), .A2(n14855), .B1(n14253), .B2(n14853), .ZN(
        n15095) );
  OAI22_X1 U16270 ( .A1(n14279), .A2(n14899), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14225), .ZN(n14226) );
  AOI21_X1 U16271 ( .B1(n15095), .B2(n14282), .A(n14226), .ZN(n14227) );
  OAI211_X1 U16272 ( .C1(n14903), .C2(n14285), .A(n14228), .B(n14227), .ZN(
        P1_U3233) );
  NAND2_X1 U16273 ( .A1(n14230), .A2(n14229), .ZN(n14233) );
  OAI211_X1 U16274 ( .C1(n14233), .C2(n14232), .A(n14231), .B(n14273), .ZN(
        n14239) );
  NOR2_X1 U16275 ( .A1(n14279), .A2(n14234), .ZN(n14235) );
  AOI211_X1 U16276 ( .C1(n14282), .C2(n14237), .A(n14236), .B(n14235), .ZN(
        n14238) );
  OAI211_X1 U16277 ( .C1(n14240), .C2(n14285), .A(n14239), .B(n14238), .ZN(
        P1_U3234) );
  OAI21_X1 U16278 ( .B1(n14243), .B2(n14242), .A(n14241), .ZN(n14244) );
  NAND2_X1 U16279 ( .A1(n14244), .A2(n14273), .ZN(n14250) );
  NAND2_X1 U16280 ( .A1(n14832), .A2(n15010), .ZN(n14246) );
  NAND2_X1 U16281 ( .A1(n14544), .A2(n15008), .ZN(n14245) );
  NAND2_X1 U16282 ( .A1(n14246), .A2(n14245), .ZN(n15083) );
  OAI22_X1 U16283 ( .A1(n14873), .A2(n14279), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14247), .ZN(n14248) );
  AOI21_X1 U16284 ( .B1(n15083), .B2(n14282), .A(n14248), .ZN(n14249) );
  OAI211_X1 U16285 ( .C1(n14285), .C2(n14877), .A(n14250), .B(n14249), .ZN(
        P1_U3235) );
  XOR2_X1 U16286 ( .A(n14252), .B(n14251), .Z(n14259) );
  NAND2_X1 U16287 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n14703)
         );
  OAI21_X1 U16288 ( .B1(n14253), .B2(n14267), .A(n14703), .ZN(n14257) );
  OAI22_X1 U16289 ( .A1(n14255), .A2(n14254), .B1(n14279), .B2(n14935), .ZN(
        n14256) );
  AOI211_X1 U16290 ( .C1(n15109), .C2(n14269), .A(n14257), .B(n14256), .ZN(
        n14258) );
  OAI21_X1 U16291 ( .B1(n14259), .B2(n14271), .A(n14258), .ZN(P1_U3238) );
  XOR2_X1 U16292 ( .A(n14261), .B(n14260), .Z(n14272) );
  AOI22_X1 U16293 ( .A1(n14263), .A2(n14262), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14266) );
  NAND2_X1 U16294 ( .A1(n14833), .A2(n14264), .ZN(n14265) );
  OAI211_X1 U16295 ( .C1(n14750), .C2(n14267), .A(n14266), .B(n14265), .ZN(
        n14268) );
  AOI21_X1 U16296 ( .B1(n15060), .B2(n14269), .A(n14268), .ZN(n14270) );
  OAI21_X1 U16297 ( .B1(n14272), .B2(n14271), .A(n14270), .ZN(P1_U3240) );
  OAI211_X1 U16298 ( .C1(n14276), .C2(n14275), .A(n14274), .B(n14273), .ZN(
        n14284) );
  NAND2_X1 U16299 ( .A1(n14954), .A2(n15010), .ZN(n14278) );
  NAND2_X1 U16300 ( .A1(n14546), .A2(n15008), .ZN(n14277) );
  NAND2_X1 U16301 ( .A1(n14278), .A2(n14277), .ZN(n15129) );
  NOR2_X1 U16302 ( .A1(n14279), .A2(n14986), .ZN(n14280) );
  AOI211_X1 U16303 ( .C1(n14282), .C2(n15129), .A(n14281), .B(n14280), .ZN(
        n14283) );
  OAI211_X1 U16304 ( .C1(n14995), .C2(n14285), .A(n14284), .B(n14283), .ZN(
        P1_U3241) );
  XNOR2_X1 U16305 ( .A(n14286), .B(n14738), .ZN(n14424) );
  MUX2_X1 U16306 ( .A(n14555), .B(n14309), .S(n14436), .Z(n14311) );
  INV_X2 U16307 ( .A(n14441), .ZN(n14484) );
  AOI21_X1 U16308 ( .B1(n14302), .B2(n14287), .A(n14484), .ZN(n14288) );
  AND2_X1 U16309 ( .A1(n14302), .A2(n14436), .ZN(n14290) );
  AOI21_X1 U16310 ( .B1(n14303), .B2(n14288), .A(n14290), .ZN(n14308) );
  OAI21_X1 U16311 ( .B1(n14293), .B2(n14292), .A(n14291), .ZN(n14294) );
  NAND2_X1 U16312 ( .A1(n6853), .A2(n15279), .ZN(n15251) );
  NAND3_X1 U16313 ( .A1(n14296), .A2(n14295), .A3(n8892), .ZN(n14297) );
  NAND3_X1 U16314 ( .A1(n14303), .A2(n15286), .A3(n6412), .ZN(n14300) );
  NAND3_X1 U16315 ( .A1(n14302), .A2(n14298), .A3(n14436), .ZN(n14299) );
  NAND2_X1 U16316 ( .A1(n14300), .A2(n14299), .ZN(n14301) );
  NAND2_X1 U16317 ( .A1(n14305), .A2(n14301), .ZN(n14307) );
  AND4_X1 U16318 ( .A1(n14303), .A2(n14302), .A3(n15261), .A4(n14557), .ZN(
        n14304) );
  NAND2_X1 U16319 ( .A1(n14305), .A2(n14304), .ZN(n14306) );
  MUX2_X1 U16320 ( .A(n14555), .B(n14309), .S(n6412), .Z(n14310) );
  MUX2_X1 U16321 ( .A(n14554), .B(n14313), .S(n6412), .Z(n14321) );
  INV_X1 U16322 ( .A(n14321), .ZN(n14314) );
  MUX2_X1 U16323 ( .A(n14554), .B(n14313), .S(n14436), .Z(n14320) );
  NAND2_X1 U16324 ( .A1(n14314), .A2(n14320), .ZN(n14315) );
  MUX2_X1 U16325 ( .A(n14552), .B(n14325), .S(n14441), .Z(n14328) );
  NAND2_X1 U16326 ( .A1(n14325), .A2(n14552), .ZN(n14316) );
  AND2_X1 U16327 ( .A1(n14328), .A2(n14316), .ZN(n14317) );
  NOR2_X1 U16328 ( .A1(n14318), .A2(n14317), .ZN(n14338) );
  MUX2_X1 U16329 ( .A(n14553), .B(n14319), .S(n14436), .Z(n14336) );
  INV_X1 U16330 ( .A(n14336), .ZN(n14323) );
  MUX2_X1 U16331 ( .A(n14553), .B(n14319), .S(n6412), .Z(n14335) );
  INV_X1 U16332 ( .A(n14320), .ZN(n14322) );
  AOI22_X1 U16333 ( .A1(n14323), .A2(n14335), .B1(n14322), .B2(n14321), .ZN(
        n14324) );
  NOR2_X1 U16334 ( .A1(n14326), .A2(n6410), .ZN(n14331) );
  AND2_X1 U16335 ( .A1(n14327), .A2(n14552), .ZN(n14330) );
  INV_X1 U16336 ( .A(n14328), .ZN(n14329) );
  OAI21_X1 U16337 ( .B1(n14331), .B2(n14330), .A(n14329), .ZN(n14341) );
  INV_X1 U16338 ( .A(n14332), .ZN(n14334) );
  MUX2_X1 U16339 ( .A(n14551), .B(n15335), .S(n6412), .Z(n14333) );
  OR2_X1 U16340 ( .A1(n14334), .A2(n14333), .ZN(n14340) );
  INV_X1 U16341 ( .A(n14335), .ZN(n14337) );
  NAND3_X1 U16342 ( .A1(n14338), .A2(n14337), .A3(n14336), .ZN(n14339) );
  NAND4_X1 U16343 ( .A1(n14342), .A2(n14341), .A3(n14340), .A4(n14339), .ZN(
        n14347) );
  MUX2_X1 U16344 ( .A(n14343), .B(n15345), .S(n6412), .Z(n14346) );
  MUX2_X1 U16345 ( .A(n14550), .B(n14344), .S(n14436), .Z(n14345) );
  OAI21_X1 U16346 ( .B1(n14347), .B2(n14346), .A(n14345), .ZN(n14349) );
  NAND2_X1 U16347 ( .A1(n14347), .A2(n14346), .ZN(n14348) );
  MUX2_X1 U16348 ( .A(n14549), .B(n14350), .S(n14436), .Z(n14352) );
  MUX2_X1 U16349 ( .A(n14549), .B(n14350), .S(n14441), .Z(n14351) );
  MUX2_X1 U16350 ( .A(n14548), .B(n15154), .S(n6412), .Z(n14354) );
  MUX2_X1 U16351 ( .A(n14548), .B(n15154), .S(n14436), .Z(n14353) );
  MUX2_X1 U16352 ( .A(n14547), .B(n15149), .S(n14436), .Z(n14358) );
  MUX2_X1 U16353 ( .A(n14547), .B(n15149), .S(n6412), .Z(n14356) );
  NAND2_X1 U16354 ( .A1(n14357), .A2(n14356), .ZN(n14360) );
  MUX2_X1 U16355 ( .A(n15009), .B(n15144), .S(n6412), .Z(n14367) );
  NAND3_X1 U16356 ( .A1(n14365), .A2(n15006), .A3(n15144), .ZN(n14363) );
  NAND3_X1 U16357 ( .A1(n14363), .A2(n14368), .A3(n14362), .ZN(n14364) );
  NAND2_X1 U16358 ( .A1(n14364), .A2(n14484), .ZN(n14379) );
  INV_X1 U16359 ( .A(n14366), .ZN(n14375) );
  INV_X1 U16360 ( .A(n14367), .ZN(n14369) );
  AND3_X1 U16361 ( .A1(n15006), .A2(n14369), .A3(n14368), .ZN(n14374) );
  AOI21_X1 U16362 ( .B1(n14371), .B2(n14370), .A(n14484), .ZN(n14373) );
  OAI21_X1 U16363 ( .B1(n14371), .B2(n14370), .A(n15130), .ZN(n14372) );
  NAND2_X1 U16364 ( .A1(n14379), .A2(n14378), .ZN(n14389) );
  INV_X1 U16365 ( .A(n14380), .ZN(n14381) );
  OR2_X1 U16366 ( .A1(n14382), .A2(n14381), .ZN(n14946) );
  MUX2_X1 U16367 ( .A(n14954), .B(n15122), .S(n6412), .Z(n14391) );
  NAND2_X1 U16368 ( .A1(n15122), .A2(n14484), .ZN(n14383) );
  OAI211_X1 U16369 ( .C1(n14384), .C2(n14484), .A(n14391), .B(n14383), .ZN(
        n14385) );
  OAI211_X1 U16370 ( .C1(n14441), .C2(n14386), .A(n14946), .B(n14385), .ZN(
        n14387) );
  INV_X1 U16371 ( .A(n14387), .ZN(n14388) );
  NAND2_X1 U16372 ( .A1(n14389), .A2(n14388), .ZN(n14396) );
  MUX2_X1 U16373 ( .A(n14943), .B(n14390), .S(n6412), .Z(n14395) );
  INV_X1 U16374 ( .A(n14391), .ZN(n14393) );
  MUX2_X1 U16375 ( .A(n14954), .B(n15122), .S(n14436), .Z(n14392) );
  NAND3_X1 U16376 ( .A1(n14946), .A2(n14393), .A3(n14392), .ZN(n14394) );
  NAND4_X1 U16377 ( .A1(n14396), .A2(n14395), .A3(n7803), .A4(n14394), .ZN(
        n14400) );
  INV_X1 U16378 ( .A(n14912), .ZN(n14910) );
  NAND2_X1 U16379 ( .A1(n15109), .A2(n6412), .ZN(n14398) );
  OR2_X1 U16380 ( .A1(n15109), .A2(n6412), .ZN(n14397) );
  MUX2_X1 U16381 ( .A(n14398), .B(n14397), .S(n14956), .Z(n14399) );
  NAND3_X1 U16382 ( .A1(n14400), .A2(n14910), .A3(n14399), .ZN(n14404) );
  MUX2_X1 U16383 ( .A(n14402), .B(n14401), .S(n6412), .Z(n14403) );
  MUX2_X1 U16384 ( .A(n14405), .B(n14903), .S(n6412), .Z(n14407) );
  MUX2_X1 U16385 ( .A(n14545), .B(n15096), .S(n14436), .Z(n14406) );
  MUX2_X1 U16386 ( .A(n14544), .B(n14891), .S(n14436), .Z(n14409) );
  MUX2_X1 U16387 ( .A(n14544), .B(n14891), .S(n6412), .Z(n14408) );
  MUX2_X1 U16388 ( .A(n14543), .B(n15084), .S(n6412), .Z(n14411) );
  MUX2_X1 U16389 ( .A(n14852), .B(n14877), .S(n14436), .Z(n14410) );
  MUX2_X1 U16390 ( .A(n14832), .B(n15078), .S(n14436), .Z(n14412) );
  MUX2_X1 U16391 ( .A(n14832), .B(n15078), .S(n6412), .Z(n14413) );
  MUX2_X1 U16392 ( .A(n14542), .B(n14840), .S(n14441), .Z(n14416) );
  NAND2_X1 U16393 ( .A1(n14417), .A2(n14416), .ZN(n14415) );
  MUX2_X1 U16394 ( .A(n14542), .B(n14840), .S(n14484), .Z(n14414) );
  NAND2_X1 U16395 ( .A1(n14415), .A2(n14414), .ZN(n14419) );
  OR2_X1 U16396 ( .A1(n14417), .A2(n14416), .ZN(n14418) );
  NAND2_X1 U16397 ( .A1(n14419), .A2(n14418), .ZN(n14423) );
  MUX2_X1 U16398 ( .A(n14833), .B(n15065), .S(n14484), .Z(n14422) );
  NAND2_X1 U16399 ( .A1(n14423), .A2(n14422), .ZN(n14421) );
  MUX2_X1 U16400 ( .A(n14833), .B(n15065), .S(n14441), .Z(n14420) );
  INV_X1 U16401 ( .A(n14424), .ZN(n14426) );
  NAND2_X1 U16402 ( .A1(n14540), .A2(n14484), .ZN(n14425) );
  OAI21_X1 U16403 ( .B1(n14483), .B2(n14426), .A(n14425), .ZN(n14433) );
  INV_X1 U16404 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14431) );
  NAND2_X1 U16405 ( .A1(n14427), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n14430) );
  INV_X1 U16406 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14428) );
  OR2_X1 U16407 ( .A1(n9079), .A2(n14428), .ZN(n14429) );
  OAI211_X1 U16408 ( .C1(n14432), .C2(n14431), .A(n14430), .B(n14429), .ZN(
        n14764) );
  AND2_X1 U16409 ( .A1(n14433), .A2(n14764), .ZN(n14434) );
  AOI21_X1 U16410 ( .B1(n14499), .B2(n6412), .A(n14434), .ZN(n14464) );
  OAI21_X1 U16411 ( .B1(n14540), .B2(n14482), .A(n14764), .ZN(n14435) );
  INV_X1 U16412 ( .A(n14435), .ZN(n14437) );
  MUX2_X1 U16413 ( .A(n14437), .B(n14499), .S(n14436), .Z(n14458) );
  NAND2_X1 U16414 ( .A1(n14464), .A2(n14458), .ZN(n14440) );
  INV_X1 U16415 ( .A(n14541), .ZN(n14438) );
  INV_X1 U16416 ( .A(n14758), .ZN(n15039) );
  MUX2_X1 U16417 ( .A(n14438), .B(n15039), .S(n14441), .Z(n14452) );
  MUX2_X1 U16418 ( .A(n14541), .B(n14758), .S(n14484), .Z(n14451) );
  NAND2_X1 U16419 ( .A1(n14452), .A2(n14451), .ZN(n14439) );
  NAND2_X1 U16420 ( .A1(n14440), .A2(n14439), .ZN(n14457) );
  MUX2_X1 U16421 ( .A(n14794), .B(n15046), .S(n14441), .Z(n14456) );
  MUX2_X1 U16422 ( .A(n14761), .B(n14787), .S(n14484), .Z(n14455) );
  MUX2_X1 U16423 ( .A(n14750), .B(n7795), .S(n14441), .Z(n14467) );
  MUX2_X1 U16424 ( .A(n7796), .B(n14806), .S(n14484), .Z(n14466) );
  AND2_X1 U16425 ( .A1(n14467), .A2(n14466), .ZN(n14442) );
  NOR2_X1 U16426 ( .A1(n14468), .A2(n14442), .ZN(n14446) );
  MUX2_X1 U16427 ( .A(n14793), .B(n7470), .S(n14441), .Z(n14448) );
  MUX2_X1 U16428 ( .A(n14753), .B(n15060), .S(n14484), .Z(n14447) );
  NAND2_X1 U16429 ( .A1(n14448), .A2(n14447), .ZN(n14443) );
  INV_X1 U16430 ( .A(n14446), .ZN(n14472) );
  INV_X1 U16431 ( .A(n14447), .ZN(n14450) );
  INV_X1 U16432 ( .A(n14448), .ZN(n14449) );
  NAND2_X1 U16433 ( .A1(n14450), .A2(n14449), .ZN(n14471) );
  INV_X1 U16434 ( .A(n14451), .ZN(n14454) );
  INV_X1 U16435 ( .A(n14452), .ZN(n14453) );
  NAND2_X1 U16436 ( .A1(n14454), .A2(n14453), .ZN(n14463) );
  OR3_X1 U16437 ( .A1(n14457), .A2(n14456), .A3(n14455), .ZN(n14462) );
  NAND2_X1 U16438 ( .A1(n14463), .A2(n14464), .ZN(n14460) );
  INV_X1 U16439 ( .A(n14458), .ZN(n14459) );
  NAND2_X1 U16440 ( .A1(n14460), .A2(n14459), .ZN(n14461) );
  OAI211_X1 U16441 ( .C1(n14464), .C2(n14463), .A(n14462), .B(n14461), .ZN(
        n14465) );
  INV_X1 U16442 ( .A(n14465), .ZN(n14470) );
  OR3_X1 U16443 ( .A1(n14468), .A2(n14467), .A3(n14466), .ZN(n14469) );
  OAI211_X1 U16444 ( .C1(n14472), .C2(n14471), .A(n14470), .B(n14469), .ZN(
        n14473) );
  INV_X1 U16445 ( .A(n14487), .ZN(n14534) );
  NAND2_X1 U16446 ( .A1(n14474), .A2(n8962), .ZN(n14478) );
  INV_X1 U16447 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14475) );
  OR2_X1 U16448 ( .A1(n14476), .A2(n14475), .ZN(n14477) );
  NOR2_X1 U16449 ( .A1(n14743), .A2(n14484), .ZN(n14490) );
  NAND2_X1 U16450 ( .A1(n14286), .A2(n14482), .ZN(n14480) );
  AOI21_X1 U16451 ( .B1(n14481), .B2(n14480), .A(n14479), .ZN(n14491) );
  INV_X1 U16452 ( .A(n14491), .ZN(n14489) );
  OR2_X1 U16453 ( .A1(n14483), .A2(n14482), .ZN(n14528) );
  NAND2_X1 U16454 ( .A1(n14489), .A2(n14528), .ZN(n14488) );
  NAND2_X1 U16455 ( .A1(n14743), .A2(n14484), .ZN(n14497) );
  NOR2_X1 U16456 ( .A1(n14497), .A2(n14540), .ZN(n14485) );
  AOI211_X1 U16457 ( .C1(n14490), .C2(n14540), .A(n14488), .B(n14485), .ZN(
        n14533) );
  XNOR2_X1 U16458 ( .A(n14743), .B(n14540), .ZN(n14524) );
  AND2_X1 U16459 ( .A1(n14524), .A2(n14491), .ZN(n14486) );
  NOR3_X1 U16460 ( .A1(n15028), .A2(n14540), .A3(n14488), .ZN(n14498) );
  NOR3_X1 U16461 ( .A1(n14497), .A2(n14540), .A3(n14489), .ZN(n14496) );
  XOR2_X1 U16462 ( .A(n14491), .B(n14490), .Z(n14494) );
  INV_X1 U16463 ( .A(n14540), .ZN(n14493) );
  INV_X1 U16464 ( .A(n14528), .ZN(n14492) );
  NOR4_X1 U16465 ( .A1(n14494), .A2(n14493), .A3(n14492), .A4(n14743), .ZN(
        n14495) );
  AOI211_X1 U16466 ( .C1(n14498), .C2(n14497), .A(n14496), .B(n14495), .ZN(
        n14531) );
  XOR2_X1 U16467 ( .A(n14764), .B(n14499), .Z(n14523) );
  NAND2_X1 U16468 ( .A1(n14787), .A2(n14794), .ZN(n14751) );
  OR2_X1 U16469 ( .A1(n14787), .A2(n14794), .ZN(n14500) );
  NAND2_X1 U16470 ( .A1(n14751), .A2(n14500), .ZN(n14776) );
  INV_X1 U16471 ( .A(n14776), .ZN(n14780) );
  INV_X1 U16472 ( .A(n14946), .ZN(n14950) );
  INV_X1 U16473 ( .A(n14501), .ZN(n14507) );
  NAND4_X1 U16474 ( .A1(n14503), .A2(n11022), .A3(n15273), .A4(n15253), .ZN(
        n14505) );
  INV_X1 U16475 ( .A(n14508), .ZN(n14509) );
  NAND4_X1 U16476 ( .A1(n14512), .A2(n14511), .A3(n14510), .A4(n14509), .ZN(
        n14514) );
  NOR4_X1 U16477 ( .A1(n7777), .A2(n14515), .A3(n14514), .A4(n14513), .ZN(
        n14517) );
  NAND4_X1 U16478 ( .A1(n14517), .A2(n12095), .A3(n15006), .A4(n14516), .ZN(
        n14518) );
  NAND4_X1 U16479 ( .A1(n14815), .A2(n14910), .A3(n14519), .A4(n14907), .ZN(
        n14520) );
  NAND4_X1 U16480 ( .A1(n14780), .A2(n14521), .A3(n14830), .A4(n14860), .ZN(
        n14522) );
  NOR3_X1 U16481 ( .A1(n14523), .A2(n14797), .A3(n14522), .ZN(n14525) );
  XNOR2_X1 U16482 ( .A(n14758), .B(n14541), .ZN(n14757) );
  NAND3_X1 U16483 ( .A1(n14525), .A2(n14757), .A3(n14524), .ZN(n14527) );
  AND2_X1 U16484 ( .A1(n15245), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14535) );
  NAND3_X1 U16485 ( .A1(n14536), .A2(n15008), .A3(n14535), .ZN(n14537) );
  OAI211_X1 U16486 ( .C1(n15198), .C2(n14539), .A(n14537), .B(P1_B_REG_SCAN_IN), .ZN(n14538) );
  MUX2_X1 U16487 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14540), .S(P1_U4016), .Z(
        P1_U3591) );
  MUX2_X1 U16488 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14764), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16489 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14541), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16490 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14761), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16491 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n7796), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16492 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14753), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16493 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14833), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16494 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14542), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16495 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14832), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16496 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14543), .S(P1_U4016), .Z(
        P1_U3582) );
  MUX2_X1 U16497 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14544), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U16498 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14545), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U16499 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14929), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U16500 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14956), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U16501 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14969), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16502 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14954), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16503 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n15011), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16504 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14546), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16505 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n15009), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16506 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14547), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16507 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14548), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16508 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14549), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16509 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14550), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U16510 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14551), .S(P1_U4016), .Z(
        P1_U3568) );
  MUX2_X1 U16511 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14552), .S(P1_U4016), .Z(
        P1_U3567) );
  MUX2_X1 U16512 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14553), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16513 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14554), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U16514 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14555), .S(P1_U4016), .Z(
        P1_U3564) );
  MUX2_X1 U16515 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14556), .S(P1_U4016), .Z(
        P1_U3563) );
  MUX2_X1 U16516 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14557), .S(P1_U4016), .Z(
        P1_U3562) );
  MUX2_X1 U16517 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n8892), .S(P1_U4016), .Z(
        P1_U3561) );
  MUX2_X1 U16518 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14558), .S(P1_U4016), .Z(
        P1_U3560) );
  OAI211_X1 U16519 ( .C1(n14561), .C2(n14560), .A(n14732), .B(n14559), .ZN(
        n14568) );
  AOI22_X1 U16520 ( .A1(n15247), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14567) );
  NAND2_X1 U16521 ( .A1(n14735), .A2(n14562), .ZN(n14566) );
  OAI211_X1 U16522 ( .C1(n14564), .C2(n14574), .A(n14737), .B(n14563), .ZN(
        n14565) );
  NAND4_X1 U16523 ( .A1(n14568), .A2(n14567), .A3(n14566), .A4(n14565), .ZN(
        P1_U3244) );
  AOI21_X1 U16524 ( .B1(n15245), .B2(n14569), .A(n15193), .ZN(n15244) );
  NAND2_X1 U16525 ( .A1(n14570), .A2(n14573), .ZN(n14572) );
  OAI211_X1 U16526 ( .C1(n14574), .C2(n14573), .A(n14572), .B(n14571), .ZN(
        n14575) );
  OAI211_X1 U16527 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n15244), .A(n14575), .B(
        P1_U4016), .ZN(n14618) );
  AOI22_X1 U16528 ( .A1(n15247), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n14588) );
  OAI21_X1 U16529 ( .B1(n14578), .B2(n14577), .A(n14576), .ZN(n14583) );
  OAI211_X1 U16530 ( .C1(n14581), .C2(n14580), .A(n14737), .B(n14579), .ZN(
        n14582) );
  OAI21_X1 U16531 ( .B1(n14583), .B2(n14733), .A(n14582), .ZN(n14584) );
  INV_X1 U16532 ( .A(n14584), .ZN(n14587) );
  NAND2_X1 U16533 ( .A1(n14735), .A2(n14585), .ZN(n14586) );
  NAND4_X1 U16534 ( .A1(n14618), .A2(n14588), .A3(n14587), .A4(n14586), .ZN(
        P1_U3245) );
  INV_X1 U16535 ( .A(n14589), .ZN(n14593) );
  NAND2_X1 U16536 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n14590) );
  OAI21_X1 U16537 ( .B1(n14742), .B2(n14591), .A(n14590), .ZN(n14592) );
  AOI21_X1 U16538 ( .B1(n14593), .B2(n14735), .A(n14592), .ZN(n14602) );
  OAI211_X1 U16539 ( .C1(n14596), .C2(n14595), .A(n14732), .B(n14594), .ZN(
        n14601) );
  OAI211_X1 U16540 ( .C1(n14599), .C2(n14598), .A(n14737), .B(n14597), .ZN(
        n14600) );
  NAND3_X1 U16541 ( .A1(n14602), .A2(n14601), .A3(n14600), .ZN(P1_U3246) );
  INV_X1 U16542 ( .A(n14603), .ZN(n14604) );
  AOI21_X1 U16543 ( .B1(n15247), .B2(P1_ADDR_REG_4__SCAN_IN), .A(n14604), .ZN(
        n14617) );
  OAI21_X1 U16544 ( .B1(n14607), .B2(n14606), .A(n14605), .ZN(n14612) );
  OAI211_X1 U16545 ( .C1(n14610), .C2(n14609), .A(n14737), .B(n14608), .ZN(
        n14611) );
  OAI21_X1 U16546 ( .B1(n14733), .B2(n14612), .A(n14611), .ZN(n14613) );
  INV_X1 U16547 ( .A(n14613), .ZN(n14616) );
  NAND2_X1 U16548 ( .A1(n14735), .A2(n14614), .ZN(n14615) );
  NAND4_X1 U16549 ( .A1(n14618), .A2(n14617), .A3(n14616), .A4(n14615), .ZN(
        P1_U3247) );
  NAND2_X1 U16550 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n14619) );
  OAI21_X1 U16551 ( .B1(n14742), .B2(n14620), .A(n14619), .ZN(n14621) );
  AOI21_X1 U16552 ( .B1(n14622), .B2(n14735), .A(n14621), .ZN(n14632) );
  OAI21_X1 U16553 ( .B1(n14625), .B2(n14624), .A(n14623), .ZN(n14626) );
  NAND2_X1 U16554 ( .A1(n14732), .A2(n14626), .ZN(n14631) );
  OAI211_X1 U16555 ( .C1(n14629), .C2(n14628), .A(n14737), .B(n14627), .ZN(
        n14630) );
  NAND3_X1 U16556 ( .A1(n14632), .A2(n14631), .A3(n14630), .ZN(P1_U3248) );
  INV_X1 U16557 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14634) );
  OAI21_X1 U16558 ( .B1(n14742), .B2(n14634), .A(n14633), .ZN(n14635) );
  AOI21_X1 U16559 ( .B1(n14636), .B2(n14735), .A(n14635), .ZN(n14645) );
  OAI211_X1 U16560 ( .C1(n14639), .C2(n14638), .A(n14737), .B(n14637), .ZN(
        n14644) );
  OAI211_X1 U16561 ( .C1(n14642), .C2(n14641), .A(n14732), .B(n14640), .ZN(
        n14643) );
  NAND3_X1 U16562 ( .A1(n14645), .A2(n14644), .A3(n14643), .ZN(P1_U3250) );
  OAI21_X1 U16563 ( .B1(n14742), .B2(n8719), .A(n14646), .ZN(n14647) );
  AOI21_X1 U16564 ( .B1(n14648), .B2(n14735), .A(n14647), .ZN(n14658) );
  OAI21_X1 U16565 ( .B1(n14651), .B2(n14650), .A(n14649), .ZN(n14652) );
  NAND2_X1 U16566 ( .A1(n14652), .A2(n14732), .ZN(n14657) );
  OAI211_X1 U16567 ( .C1(n14655), .C2(n14654), .A(n14737), .B(n14653), .ZN(
        n14656) );
  NAND3_X1 U16568 ( .A1(n14658), .A2(n14657), .A3(n14656), .ZN(P1_U3251) );
  OAI21_X1 U16569 ( .B1(n14661), .B2(n14660), .A(n14659), .ZN(n14662) );
  NAND2_X1 U16570 ( .A1(n14662), .A2(n14732), .ZN(n14672) );
  OAI21_X1 U16571 ( .B1(n14742), .B2(n14664), .A(n14663), .ZN(n14665) );
  AOI21_X1 U16572 ( .B1(n14666), .B2(n14735), .A(n14665), .ZN(n14671) );
  OAI211_X1 U16573 ( .C1(n14669), .C2(n14668), .A(n14667), .B(n14737), .ZN(
        n14670) );
  NAND3_X1 U16574 ( .A1(n14672), .A2(n14671), .A3(n14670), .ZN(P1_U3252) );
  OAI21_X1 U16575 ( .B1(n14675), .B2(n14674), .A(n14673), .ZN(n14676) );
  NAND2_X1 U16576 ( .A1(n14676), .A2(n14732), .ZN(n14685) );
  NOR2_X1 U16577 ( .A1(n14742), .A2(n15749), .ZN(n14677) );
  AOI211_X1 U16578 ( .C1(n14735), .C2(n14679), .A(n14678), .B(n14677), .ZN(
        n14684) );
  OAI211_X1 U16579 ( .C1(n14682), .C2(n14681), .A(n14680), .B(n14737), .ZN(
        n14683) );
  NAND3_X1 U16580 ( .A1(n14685), .A2(n14684), .A3(n14683), .ZN(P1_U3254) );
  NAND2_X1 U16581 ( .A1(n14694), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n14686) );
  NAND2_X1 U16582 ( .A1(n14687), .A2(n14686), .ZN(n14690) );
  INV_X1 U16583 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14688) );
  XNOR2_X1 U16584 ( .A(n14715), .B(n14688), .ZN(n14689) );
  NAND2_X1 U16585 ( .A1(n14690), .A2(n14689), .ZN(n14717) );
  OAI211_X1 U16586 ( .C1(n14690), .C2(n14689), .A(n14717), .B(n14732), .ZN(
        n14702) );
  NOR2_X1 U16587 ( .A1(n14742), .A2(n14691), .ZN(n14692) );
  AOI211_X1 U16588 ( .C1(n14715), .C2(n14735), .A(n14693), .B(n14692), .ZN(
        n14701) );
  NAND2_X1 U16589 ( .A1(n14694), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n14695) );
  NAND2_X1 U16590 ( .A1(n14696), .A2(n14695), .ZN(n14699) );
  INV_X1 U16591 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14697) );
  XNOR2_X1 U16592 ( .A(n14715), .B(n14697), .ZN(n14698) );
  NAND2_X1 U16593 ( .A1(n14699), .A2(n14698), .ZN(n14706) );
  OAI211_X1 U16594 ( .C1(n14699), .C2(n14698), .A(n14706), .B(n14737), .ZN(
        n14700) );
  NAND3_X1 U16595 ( .A1(n14702), .A2(n14701), .A3(n14700), .ZN(P1_U3260) );
  INV_X1 U16596 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n14704) );
  OAI21_X1 U16597 ( .B1(n14742), .B2(n14704), .A(n14703), .ZN(n14714) );
  INV_X1 U16598 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14712) );
  NAND2_X1 U16599 ( .A1(n14715), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14705) );
  NAND2_X1 U16600 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  NAND2_X1 U16601 ( .A1(n14707), .A2(n14718), .ZN(n14728) );
  OR2_X1 U16602 ( .A1(n14707), .A2(n14718), .ZN(n14708) );
  NAND2_X1 U16603 ( .A1(n14728), .A2(n14708), .ZN(n14711) );
  INV_X1 U16604 ( .A(n14729), .ZN(n14709) );
  AOI211_X1 U16605 ( .C1(n14712), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        n14713) );
  AOI211_X1 U16606 ( .C1(n14735), .C2(n14718), .A(n14714), .B(n14713), .ZN(
        n14723) );
  NAND2_X1 U16607 ( .A1(n14715), .A2(P1_REG1_REG_17__SCAN_IN), .ZN(n14716) );
  NAND2_X1 U16608 ( .A1(n14717), .A2(n14716), .ZN(n14719) );
  NAND2_X1 U16609 ( .A1(n14719), .A2(n14718), .ZN(n14724) );
  OR2_X1 U16610 ( .A1(n14719), .A2(n14718), .ZN(n14720) );
  AND2_X1 U16611 ( .A1(n14724), .A2(n14720), .ZN(n14721) );
  NAND2_X1 U16612 ( .A1(n14721), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n14725) );
  OAI211_X1 U16613 ( .C1(n14721), .C2(P1_REG1_REG_18__SCAN_IN), .A(n14725), 
        .B(n14732), .ZN(n14722) );
  NAND2_X1 U16614 ( .A1(n14723), .A2(n14722), .ZN(P1_U3261) );
  NAND2_X1 U16615 ( .A1(n14725), .A2(n14724), .ZN(n14727) );
  NAND2_X1 U16616 ( .A1(n14729), .A2(n14728), .ZN(n14730) );
  XNOR2_X1 U16617 ( .A(n14730), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n14736) );
  INV_X1 U16618 ( .A(n14736), .ZN(n14731) );
  AOI22_X1 U16619 ( .A1(n14734), .A2(n14732), .B1(n14737), .B2(n14731), .ZN(
        n14739) );
  OAI211_X1 U16620 ( .C1(n7553), .C2(n14742), .A(n14741), .B(n14740), .ZN(
        P1_U3262) );
  XNOR2_X1 U16621 ( .A(n14744), .B(n14743), .ZN(n14745) );
  NAND2_X1 U16622 ( .A1(n14745), .A2(n15264), .ZN(n15027) );
  NOR2_X1 U16623 ( .A1(n15028), .A2(n14994), .ZN(n14746) );
  AOI211_X1 U16624 ( .C1(P1_REG2_REG_31__SCAN_IN), .C2(n6408), .A(n14747), .B(
        n14746), .ZN(n14748) );
  OAI21_X1 U16625 ( .B1(n15027), .B2(n14982), .A(n14748), .ZN(P1_U3263) );
  AOI22_X1 U16626 ( .A1(n14755), .A2(n14754), .B1(n15060), .B2(n14753), .ZN(
        n14756) );
  AOI21_X1 U16627 ( .B1(n14783), .B2(n14758), .A(n15280), .ZN(n14760) );
  NAND2_X1 U16628 ( .A1(n15041), .A2(n15268), .ZN(n14772) );
  NAND2_X1 U16629 ( .A1(n14761), .A2(n15008), .ZN(n15038) );
  INV_X1 U16630 ( .A(n15038), .ZN(n14770) );
  INV_X1 U16631 ( .A(n14762), .ZN(n14766) );
  NAND2_X1 U16632 ( .A1(n14764), .A2(n14763), .ZN(n15037) );
  INV_X1 U16633 ( .A(n15037), .ZN(n14765) );
  AOI22_X1 U16634 ( .A1(n6408), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n14766), 
        .B2(n14765), .ZN(n14767) );
  OAI21_X1 U16635 ( .B1(n14768), .B2(n14977), .A(n14767), .ZN(n14769) );
  AOI21_X1 U16636 ( .B1(n14770), .B2(n14993), .A(n14769), .ZN(n14771) );
  OAI211_X1 U16637 ( .C1(n15039), .C2(n14994), .A(n14772), .B(n14771), .ZN(
        n14773) );
  AOI21_X1 U16638 ( .B1(n15042), .B2(n15024), .A(n14773), .ZN(n14774) );
  OAI21_X1 U16639 ( .B1(n15043), .B2(n15026), .A(n14774), .ZN(P1_U3356) );
  AOI21_X1 U16640 ( .B1(n14777), .B2(n14776), .A(n14775), .ZN(n15050) );
  AOI21_X1 U16641 ( .B1(n14780), .B2(n14779), .A(n14778), .ZN(n15048) );
  INV_X1 U16642 ( .A(n14803), .ZN(n14781) );
  AOI21_X1 U16643 ( .B1(n14781), .B2(n14787), .A(n15280), .ZN(n14782) );
  NAND2_X1 U16644 ( .A1(n14783), .A2(n14782), .ZN(n15045) );
  AOI22_X1 U16645 ( .A1(n14784), .A2(n15262), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n6408), .ZN(n14785) );
  OAI21_X1 U16646 ( .B1(n15044), .B2(n6408), .A(n14785), .ZN(n14786) );
  AOI21_X1 U16647 ( .B1(n14787), .B2(n15260), .A(n14786), .ZN(n14788) );
  OAI21_X1 U16648 ( .B1(n15045), .B2(n14982), .A(n14788), .ZN(n14789) );
  AOI21_X1 U16649 ( .B1(n15048), .B2(n15024), .A(n14789), .ZN(n14790) );
  OAI21_X1 U16650 ( .B1(n15050), .B2(n15026), .A(n14790), .ZN(P1_U3265) );
  OAI21_X1 U16651 ( .B1(n14792), .B2(n14797), .A(n14791), .ZN(n15051) );
  NAND2_X1 U16652 ( .A1(n15051), .A2(n15348), .ZN(n14802) );
  OAI22_X1 U16653 ( .A1(n14794), .A2(n14855), .B1(n14793), .B2(n14853), .ZN(
        n14795) );
  INV_X1 U16654 ( .A(n14795), .ZN(n14801) );
  AND3_X1 U16655 ( .A1(n14749), .A2(n14797), .A3(n14796), .ZN(n14798) );
  OAI21_X1 U16656 ( .B1(n14799), .B2(n14798), .A(n15311), .ZN(n14800) );
  NAND3_X1 U16657 ( .A1(n14802), .A2(n14801), .A3(n14800), .ZN(n15055) );
  INV_X1 U16658 ( .A(n15055), .ZN(n14811) );
  OAI21_X1 U16659 ( .B1(n6497), .B2(n7795), .A(n15264), .ZN(n14804) );
  OR2_X1 U16660 ( .A1(n14804), .A2(n14803), .ZN(n15052) );
  AOI22_X1 U16661 ( .A1(n14805), .A2(n15262), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n6408), .ZN(n14808) );
  NAND2_X1 U16662 ( .A1(n14806), .A2(n15260), .ZN(n14807) );
  OAI211_X1 U16663 ( .C1(n15052), .C2(n14982), .A(n14808), .B(n14807), .ZN(
        n14809) );
  AOI21_X1 U16664 ( .B1(n15051), .B2(n15269), .A(n14809), .ZN(n14810) );
  OAI21_X1 U16665 ( .B1(n14811), .B2(n6408), .A(n14810), .ZN(P1_U3266) );
  INV_X1 U16666 ( .A(n15064), .ZN(n14827) );
  AND2_X1 U16667 ( .A1(n14816), .A2(n14815), .ZN(n14817) );
  NOR2_X1 U16668 ( .A1(n14818), .A2(n14817), .ZN(n15069) );
  AOI21_X1 U16669 ( .B1(n14837), .B2(n15065), .A(n15280), .ZN(n14820) );
  NAND2_X1 U16670 ( .A1(n14820), .A2(n14819), .ZN(n15067) );
  AOI22_X1 U16671 ( .A1(n14821), .A2(n15262), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n6408), .ZN(n14822) );
  OAI21_X1 U16672 ( .B1(n15066), .B2(n6408), .A(n14822), .ZN(n14823) );
  AOI21_X1 U16673 ( .B1(n15065), .B2(n15260), .A(n14823), .ZN(n14824) );
  OAI21_X1 U16674 ( .B1(n15067), .B2(n14982), .A(n14824), .ZN(n14825) );
  AOI21_X1 U16675 ( .B1(n15069), .B2(n15024), .A(n14825), .ZN(n14826) );
  OAI21_X1 U16676 ( .B1(n14827), .B2(n15026), .A(n14826), .ZN(P1_U3268) );
  OAI211_X1 U16677 ( .C1(n14831), .C2(n14830), .A(n14829), .B(n15311), .ZN(
        n14835) );
  AOI22_X1 U16678 ( .A1(n14833), .A2(n15010), .B1(n15008), .B2(n14832), .ZN(
        n14834) );
  OAI211_X1 U16679 ( .C1(n15072), .C2(n15294), .A(n14835), .B(n14834), .ZN(
        n15076) );
  NAND2_X1 U16680 ( .A1(n15076), .A2(n14993), .ZN(n14846) );
  INV_X1 U16681 ( .A(n14836), .ZN(n14839) );
  INV_X1 U16682 ( .A(n14837), .ZN(n14838) );
  AOI211_X1 U16683 ( .C1(n14840), .C2(n14839), .A(n15280), .B(n14838), .ZN(
        n15074) );
  AOI22_X1 U16684 ( .A1(n14841), .A2(n15262), .B1(P1_REG2_REG_24__SCAN_IN), 
        .B2(n6408), .ZN(n14842) );
  OAI21_X1 U16685 ( .B1(n14843), .B2(n14994), .A(n14842), .ZN(n14844) );
  AOI21_X1 U16686 ( .B1(n15074), .B2(n15268), .A(n14844), .ZN(n14845) );
  OAI211_X1 U16687 ( .C1(n15072), .C2(n14939), .A(n14846), .B(n14845), .ZN(
        P1_U3269) );
  INV_X1 U16688 ( .A(n14847), .ZN(n14865) );
  NOR3_X1 U16689 ( .A1(n14865), .A2(n7779), .A3(n14860), .ZN(n14851) );
  INV_X1 U16690 ( .A(n14849), .ZN(n14850) );
  OAI21_X1 U16691 ( .B1(n14851), .B2(n14850), .A(n15311), .ZN(n15080) );
  XNOR2_X1 U16692 ( .A(n14871), .B(n14859), .ZN(n14856) );
  OAI222_X1 U16693 ( .A1(n15280), .A2(n14856), .B1(n14855), .B2(n14854), .C1(
        n14853), .C2(n14852), .ZN(n15077) );
  AOI22_X1 U16694 ( .A1(n14857), .A2(n15262), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n6408), .ZN(n14858) );
  OAI21_X1 U16695 ( .B1(n14859), .B2(n14994), .A(n14858), .ZN(n14863) );
  XNOR2_X1 U16696 ( .A(n14861), .B(n14860), .ZN(n15081) );
  NOR2_X1 U16697 ( .A1(n15081), .A2(n14925), .ZN(n14862) );
  AOI211_X1 U16698 ( .C1(n15268), .C2(n15077), .A(n14863), .B(n14862), .ZN(
        n14864) );
  OAI21_X1 U16699 ( .B1(n15080), .B2(n6408), .A(n14864), .ZN(P1_U3270) );
  AOI21_X1 U16700 ( .B1(n14869), .B2(n14866), .A(n14865), .ZN(n15088) );
  AND2_X1 U16701 ( .A1(n14868), .A2(n14867), .ZN(n14870) );
  XNOR2_X1 U16702 ( .A(n14870), .B(n14869), .ZN(n15085) );
  AOI211_X1 U16703 ( .C1(n15084), .C2(n14889), .A(n15280), .B(n14871), .ZN(
        n15082) );
  NAND2_X1 U16704 ( .A1(n15082), .A2(n15268), .ZN(n14876) );
  INV_X1 U16705 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n14872) );
  OAI22_X1 U16706 ( .A1(n14873), .A2(n14977), .B1(n14872), .B2(n14993), .ZN(
        n14874) );
  AOI21_X1 U16707 ( .B1(n15083), .B2(n14993), .A(n14874), .ZN(n14875) );
  OAI211_X1 U16708 ( .C1(n14994), .C2(n14877), .A(n14876), .B(n14875), .ZN(
        n14878) );
  AOI21_X1 U16709 ( .B1(n15085), .B2(n15024), .A(n14878), .ZN(n14879) );
  OAI21_X1 U16710 ( .B1(n15088), .B2(n15026), .A(n14879), .ZN(P1_U3271) );
  XNOR2_X1 U16711 ( .A(n14880), .B(n14887), .ZN(n14882) );
  AOI21_X1 U16712 ( .B1(n14882), .B2(n15311), .A(n14881), .ZN(n15093) );
  OR2_X1 U16713 ( .A1(n14883), .A2(n14907), .ZN(n14905) );
  AND2_X1 U16714 ( .A1(n14905), .A2(n14884), .ZN(n14888) );
  NAND2_X1 U16715 ( .A1(n14905), .A2(n14885), .ZN(n14886) );
  OAI21_X1 U16716 ( .B1(n14888), .B2(n14887), .A(n14886), .ZN(n15089) );
  OAI211_X1 U16717 ( .C1(n6499), .C2(n7466), .A(n15264), .B(n14889), .ZN(
        n15090) );
  AOI22_X1 U16718 ( .A1(n14890), .A2(n15262), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n6408), .ZN(n14893) );
  NAND2_X1 U16719 ( .A1(n14891), .A2(n15260), .ZN(n14892) );
  OAI211_X1 U16720 ( .C1(n15090), .C2(n14982), .A(n14893), .B(n14892), .ZN(
        n14894) );
  AOI21_X1 U16721 ( .B1(n15089), .B2(n15024), .A(n14894), .ZN(n14895) );
  OAI21_X1 U16722 ( .B1(n15093), .B2(n6408), .A(n14895), .ZN(P1_U3272) );
  OAI21_X1 U16723 ( .B1(n14897), .B2(n14907), .A(n14896), .ZN(n15100) );
  INV_X1 U16724 ( .A(n14915), .ZN(n14898) );
  AOI211_X1 U16725 ( .C1(n15096), .C2(n14898), .A(n15280), .B(n6499), .ZN(
        n15094) );
  NAND2_X1 U16726 ( .A1(n6408), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14902) );
  NOR2_X1 U16727 ( .A1(n14899), .A2(n14977), .ZN(n14900) );
  OAI21_X1 U16728 ( .B1(n15095), .B2(n14900), .A(n14993), .ZN(n14901) );
  OAI211_X1 U16729 ( .C1(n14903), .C2(n14994), .A(n14902), .B(n14901), .ZN(
        n14904) );
  AOI21_X1 U16730 ( .B1(n15094), .B2(n15268), .A(n14904), .ZN(n14909) );
  INV_X1 U16731 ( .A(n14905), .ZN(n14906) );
  AOI21_X1 U16732 ( .B1(n14907), .B2(n14883), .A(n14906), .ZN(n15097) );
  NAND2_X1 U16733 ( .A1(n15097), .A2(n15024), .ZN(n14908) );
  OAI211_X1 U16734 ( .C1(n15100), .C2(n15026), .A(n14909), .B(n14908), .ZN(
        P1_U3273) );
  XNOR2_X1 U16735 ( .A(n14911), .B(n14910), .ZN(n15107) );
  XNOR2_X1 U16736 ( .A(n14913), .B(n14912), .ZN(n15101) );
  NAND2_X1 U16737 ( .A1(n15101), .A2(n14914), .ZN(n14924) );
  INV_X1 U16738 ( .A(n14934), .ZN(n14916) );
  AOI211_X1 U16739 ( .C1(n15104), .C2(n14916), .A(n15280), .B(n14915), .ZN(
        n15102) );
  INV_X1 U16740 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14918) );
  OAI22_X1 U16741 ( .A1(n14993), .A2(n14918), .B1(n14917), .B2(n14977), .ZN(
        n14919) );
  AOI21_X1 U16742 ( .B1(n15103), .B2(n14993), .A(n14919), .ZN(n14920) );
  OAI21_X1 U16743 ( .B1(n14921), .B2(n14994), .A(n14920), .ZN(n14922) );
  AOI21_X1 U16744 ( .B1(n15102), .B2(n15268), .A(n14922), .ZN(n14923) );
  OAI211_X1 U16745 ( .C1(n15107), .C2(n14925), .A(n14924), .B(n14923), .ZN(
        P1_U3274) );
  XNOR2_X1 U16746 ( .A(n14926), .B(n7803), .ZN(n14932) );
  XNOR2_X1 U16747 ( .A(n14928), .B(n14927), .ZN(n15112) );
  AOI22_X1 U16748 ( .A1(n14929), .A2(n15010), .B1(n15008), .B2(n14969), .ZN(
        n14930) );
  OAI21_X1 U16749 ( .B1(n15112), .B2(n15294), .A(n14930), .ZN(n14931) );
  AOI21_X1 U16750 ( .B1(n15311), .B2(n14932), .A(n14931), .ZN(n15111) );
  INV_X1 U16751 ( .A(n14933), .ZN(n14953) );
  AOI211_X1 U16752 ( .C1(n15109), .C2(n14953), .A(n15280), .B(n14934), .ZN(
        n15108) );
  INV_X1 U16753 ( .A(n14935), .ZN(n14936) );
  AOI22_X1 U16754 ( .A1(n6408), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14936), 
        .B2(n15262), .ZN(n14937) );
  OAI21_X1 U16755 ( .B1(n14938), .B2(n14994), .A(n14937), .ZN(n14941) );
  NOR2_X1 U16756 ( .A1(n15112), .A2(n14939), .ZN(n14940) );
  AOI211_X1 U16757 ( .C1(n15108), .C2(n15268), .A(n14941), .B(n14940), .ZN(
        n14942) );
  OAI21_X1 U16758 ( .B1(n6408), .B2(n15111), .A(n14942), .ZN(P1_U3275) );
  INV_X1 U16759 ( .A(n14943), .ZN(n14944) );
  OR2_X1 U16760 ( .A1(n14945), .A2(n14944), .ZN(n14949) );
  OR2_X1 U16761 ( .A1(n14947), .A2(n14946), .ZN(n14948) );
  NAND2_X1 U16762 ( .A1(n14949), .A2(n14948), .ZN(n15113) );
  INV_X1 U16763 ( .A(n15113), .ZN(n14964) );
  XNOR2_X1 U16764 ( .A(n14951), .B(n14950), .ZN(n15118) );
  AOI21_X1 U16765 ( .B1(n14975), .B2(n14960), .A(n15280), .ZN(n14952) );
  NAND2_X1 U16766 ( .A1(n14953), .A2(n14952), .ZN(n15115) );
  AND2_X1 U16767 ( .A1(n14954), .A2(n15008), .ZN(n14955) );
  AOI21_X1 U16768 ( .B1(n14956), .B2(n15010), .A(n14955), .ZN(n15114) );
  OAI21_X1 U16769 ( .B1(n14957), .B2(n14977), .A(n15114), .ZN(n14958) );
  MUX2_X1 U16770 ( .A(P1_REG2_REG_17__SCAN_IN), .B(n14958), .S(n14993), .Z(
        n14959) );
  AOI21_X1 U16771 ( .B1(n14960), .B2(n15260), .A(n14959), .ZN(n14961) );
  OAI21_X1 U16772 ( .B1(n15115), .B2(n14982), .A(n14961), .ZN(n14962) );
  AOI21_X1 U16773 ( .B1(n15118), .B2(n15024), .A(n14962), .ZN(n14963) );
  OAI21_X1 U16774 ( .B1(n14964), .B2(n15026), .A(n14963), .ZN(P1_U3276) );
  NAND2_X1 U16775 ( .A1(n14965), .A2(n14973), .ZN(n14966) );
  NAND2_X1 U16776 ( .A1(n14967), .A2(n14966), .ZN(n14968) );
  NAND2_X1 U16777 ( .A1(n14968), .A2(n15311), .ZN(n14971) );
  AOI22_X1 U16778 ( .A1(n14969), .A2(n15010), .B1(n15008), .B2(n15011), .ZN(
        n14970) );
  NAND2_X1 U16779 ( .A1(n14971), .A2(n14970), .ZN(n15127) );
  INV_X1 U16780 ( .A(n15127), .ZN(n14985) );
  XNOR2_X1 U16781 ( .A(n14972), .B(n14973), .ZN(n15121) );
  AOI21_X1 U16782 ( .B1(n14991), .B2(n15122), .A(n15280), .ZN(n14976) );
  NAND2_X1 U16783 ( .A1(n14976), .A2(n14975), .ZN(n15123) );
  INV_X1 U16784 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n14979) );
  OAI22_X1 U16785 ( .A1(n14993), .A2(n14979), .B1(n14978), .B2(n14977), .ZN(
        n14980) );
  AOI21_X1 U16786 ( .B1(n15122), .B2(n15260), .A(n14980), .ZN(n14981) );
  OAI21_X1 U16787 ( .B1(n15123), .B2(n14982), .A(n14981), .ZN(n14983) );
  AOI21_X1 U16788 ( .B1(n15121), .B2(n15024), .A(n14983), .ZN(n14984) );
  OAI21_X1 U16789 ( .B1(n14985), .B2(n6408), .A(n14984), .ZN(P1_U3277) );
  INV_X1 U16790 ( .A(n14986), .ZN(n14990) );
  XNOR2_X1 U16791 ( .A(n14988), .B(n14987), .ZN(n15134) );
  NOR2_X1 U16792 ( .A1(n15134), .A2(n15026), .ZN(n14989) );
  AOI211_X1 U16793 ( .C1(n15262), .C2(n14990), .A(n15129), .B(n14989), .ZN(
        n15002) );
  AOI211_X1 U16794 ( .C1(n15130), .C2(n15017), .A(n15280), .B(n14974), .ZN(
        n15128) );
  OAI22_X1 U16795 ( .A1(n14995), .A2(n14994), .B1(n14993), .B2(n14992), .ZN(
        n14996) );
  AOI21_X1 U16796 ( .B1(n15128), .B2(n15268), .A(n14996), .ZN(n15001) );
  NOR2_X1 U16797 ( .A1(n15005), .A2(n15006), .ZN(n15004) );
  NOR2_X1 U16798 ( .A1(n15004), .A2(n14997), .ZN(n14999) );
  XNOR2_X1 U16799 ( .A(n14999), .B(n14998), .ZN(n15131) );
  NAND2_X1 U16800 ( .A1(n15131), .A2(n15024), .ZN(n15000) );
  OAI211_X1 U16801 ( .C1(n15002), .C2(n6408), .A(n15001), .B(n15000), .ZN(
        P1_U3278) );
  XNOR2_X1 U16802 ( .A(n15003), .B(n15006), .ZN(n15142) );
  AOI21_X1 U16803 ( .B1(n15006), .B2(n15005), .A(n15004), .ZN(n15140) );
  INV_X1 U16804 ( .A(n15007), .ZN(n15020) );
  NAND2_X1 U16805 ( .A1(n15009), .A2(n15008), .ZN(n15013) );
  NAND2_X1 U16806 ( .A1(n15011), .A2(n15010), .ZN(n15012) );
  NAND2_X1 U16807 ( .A1(n15013), .A2(n15012), .ZN(n15135) );
  OR2_X1 U16808 ( .A1(n15015), .A2(n15014), .ZN(n15016) );
  NAND2_X1 U16809 ( .A1(n15017), .A2(n15016), .ZN(n15138) );
  NOR2_X1 U16810 ( .A1(n15138), .A2(n15018), .ZN(n15019) );
  AOI211_X1 U16811 ( .C1(n15262), .C2(n15020), .A(n15135), .B(n15019), .ZN(
        n15022) );
  AOI22_X1 U16812 ( .A1(n15136), .A2(n15260), .B1(n6408), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n15021) );
  OAI21_X1 U16813 ( .B1(n15022), .B2(n6408), .A(n15021), .ZN(n15023) );
  AOI21_X1 U16814 ( .B1(n15140), .B2(n15024), .A(n15023), .ZN(n15025) );
  OAI21_X1 U16815 ( .B1(n15142), .B2(n15026), .A(n15025), .ZN(P1_U3279) );
  OAI211_X1 U16816 ( .C1(n15028), .C2(n15344), .A(n15027), .B(n15034), .ZN(
        n15159) );
  NAND3_X1 U16817 ( .A1(n15031), .A2(n15030), .A3(n15029), .ZN(n15032) );
  MUX2_X1 U16818 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n15159), .S(n15367), .Z(
        P1_U3559) );
  OAI211_X1 U16819 ( .C1(n15036), .C2(n15344), .A(n15035), .B(n15034), .ZN(
        n15160) );
  MUX2_X1 U16820 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n15160), .S(n15367), .Z(
        P1_U3558) );
  OAI211_X1 U16821 ( .C1(n15039), .C2(n15344), .A(n15038), .B(n15037), .ZN(
        n15040) );
  OAI211_X1 U16822 ( .C1(n15046), .C2(n15344), .A(n15045), .B(n15044), .ZN(
        n15047) );
  AOI21_X1 U16823 ( .B1(n15048), .B2(n15327), .A(n15047), .ZN(n15049) );
  OAI21_X1 U16824 ( .B1(n15050), .B2(n15296), .A(n15049), .ZN(n15162) );
  MUX2_X1 U16825 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n15162), .S(n15367), .Z(
        P1_U3556) );
  INV_X1 U16826 ( .A(n15320), .ZN(n15347) );
  NAND2_X1 U16827 ( .A1(n15051), .A2(n15347), .ZN(n15053) );
  OAI211_X1 U16828 ( .C1(n7795), .C2(n15344), .A(n15053), .B(n15052), .ZN(
        n15054) );
  NOR2_X1 U16829 ( .A1(n15055), .A2(n15054), .ZN(n15163) );
  MUX2_X1 U16830 ( .A(n15056), .B(n15163), .S(n15367), .Z(n15057) );
  INV_X1 U16831 ( .A(n15057), .ZN(P1_U3555) );
  AOI21_X1 U16832 ( .B1(n15336), .B2(n15060), .A(n15059), .ZN(n15061) );
  MUX2_X1 U16833 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n15166), .S(n15367), .Z(
        P1_U3554) );
  OAI211_X1 U16834 ( .C1(n7471), .C2(n15344), .A(n15067), .B(n15066), .ZN(
        n15068) );
  AOI21_X1 U16835 ( .B1(n15069), .B2(n15327), .A(n15068), .ZN(n15070) );
  NAND2_X1 U16836 ( .A1(n15071), .A2(n15070), .ZN(n15167) );
  MUX2_X1 U16837 ( .A(n15167), .B(P1_REG1_REG_25__SCAN_IN), .S(n15365), .Z(
        P1_U3553) );
  NOR2_X1 U16838 ( .A1(n15072), .A2(n15320), .ZN(n15075) );
  MUX2_X1 U16839 ( .A(n15168), .B(P1_REG1_REG_24__SCAN_IN), .S(n15365), .Z(
        P1_U3552) );
  AOI21_X1 U16840 ( .B1(n15336), .B2(n15078), .A(n15077), .ZN(n15079) );
  OAI211_X1 U16841 ( .C1(n15340), .C2(n15081), .A(n15080), .B(n15079), .ZN(
        n15169) );
  MUX2_X1 U16842 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n15169), .S(n15367), .Z(
        P1_U3551) );
  AOI211_X1 U16843 ( .C1(n15336), .C2(n15084), .A(n15083), .B(n15082), .ZN(
        n15087) );
  NAND2_X1 U16844 ( .A1(n15085), .A2(n15327), .ZN(n15086) );
  OAI211_X1 U16845 ( .C1(n15088), .C2(n15296), .A(n15087), .B(n15086), .ZN(
        n15170) );
  MUX2_X1 U16846 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n15170), .S(n15367), .Z(
        P1_U3550) );
  NAND2_X1 U16847 ( .A1(n15089), .A2(n15327), .ZN(n15091) );
  NAND4_X1 U16848 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15171) );
  MUX2_X1 U16849 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n15171), .S(n15367), .Z(
        P1_U3549) );
  AOI211_X1 U16850 ( .C1(n15336), .C2(n15096), .A(n15095), .B(n15094), .ZN(
        n15099) );
  NAND2_X1 U16851 ( .A1(n15097), .A2(n15327), .ZN(n15098) );
  OAI211_X1 U16852 ( .C1(n15100), .C2(n15296), .A(n15099), .B(n15098), .ZN(
        n15172) );
  MUX2_X1 U16853 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n15172), .S(n15367), .Z(
        P1_U3548) );
  NAND2_X1 U16854 ( .A1(n15101), .A2(n15311), .ZN(n15106) );
  AOI211_X1 U16855 ( .C1(n15336), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15105) );
  OAI211_X1 U16856 ( .C1(n15340), .C2(n15107), .A(n15106), .B(n15105), .ZN(
        n15173) );
  MUX2_X1 U16857 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n15173), .S(n15367), .Z(
        P1_U3547) );
  AOI21_X1 U16858 ( .B1(n15336), .B2(n15109), .A(n15108), .ZN(n15110) );
  OAI211_X1 U16859 ( .C1(n15112), .C2(n15320), .A(n15111), .B(n15110), .ZN(
        n15174) );
  MUX2_X1 U16860 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n15174), .S(n15367), .Z(
        P1_U3546) );
  NAND2_X1 U16861 ( .A1(n15113), .A2(n15311), .ZN(n15120) );
  OAI211_X1 U16862 ( .C1(n15116), .C2(n15344), .A(n15115), .B(n15114), .ZN(
        n15117) );
  AOI21_X1 U16863 ( .B1(n15118), .B2(n15327), .A(n15117), .ZN(n15119) );
  NAND2_X1 U16864 ( .A1(n15120), .A2(n15119), .ZN(n15175) );
  MUX2_X1 U16865 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n15175), .S(n15367), .Z(
        P1_U3545) );
  AND2_X1 U16866 ( .A1(n15121), .A2(n15327), .ZN(n15126) );
  INV_X1 U16867 ( .A(n15122), .ZN(n15124) );
  OAI21_X1 U16868 ( .B1(n15124), .B2(n15344), .A(n15123), .ZN(n15125) );
  MUX2_X1 U16869 ( .A(n15176), .B(P1_REG1_REG_16__SCAN_IN), .S(n15365), .Z(
        P1_U3544) );
  AOI211_X1 U16870 ( .C1(n15336), .C2(n15130), .A(n15129), .B(n15128), .ZN(
        n15133) );
  NAND2_X1 U16871 ( .A1(n15131), .A2(n15327), .ZN(n15132) );
  OAI211_X1 U16872 ( .C1(n15296), .C2(n15134), .A(n15133), .B(n15132), .ZN(
        n15177) );
  MUX2_X1 U16873 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n15177), .S(n15367), .Z(
        P1_U3543) );
  AOI21_X1 U16874 ( .B1(n15136), .B2(n15336), .A(n15135), .ZN(n15137) );
  OAI21_X1 U16875 ( .B1(n15138), .B2(n15280), .A(n15137), .ZN(n15139) );
  AOI21_X1 U16876 ( .B1(n15140), .B2(n15327), .A(n15139), .ZN(n15141) );
  OAI21_X1 U16877 ( .B1(n15296), .B2(n15142), .A(n15141), .ZN(n15178) );
  MUX2_X1 U16878 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15178), .S(n15367), .Z(
        P1_U3542) );
  AOI21_X1 U16879 ( .B1(n15336), .B2(n15144), .A(n15143), .ZN(n15145) );
  OAI211_X1 U16880 ( .C1(n15340), .C2(n15147), .A(n15146), .B(n15145), .ZN(
        n15179) );
  MUX2_X1 U16881 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n15179), .S(n15367), .Z(
        P1_U3541) );
  AOI21_X1 U16882 ( .B1(n15336), .B2(n15149), .A(n15148), .ZN(n15150) );
  OAI211_X1 U16883 ( .C1(n15152), .C2(n15340), .A(n15151), .B(n15150), .ZN(
        n15180) );
  MUX2_X1 U16884 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n15180), .S(n15367), .Z(
        P1_U3540) );
  AOI21_X1 U16885 ( .B1(n15336), .B2(n15154), .A(n15153), .ZN(n15155) );
  OAI211_X1 U16886 ( .C1(n15340), .C2(n15157), .A(n15156), .B(n15155), .ZN(
        n15181) );
  MUX2_X1 U16887 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n15181), .S(n15367), .Z(
        P1_U3539) );
  MUX2_X1 U16888 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n15158), .S(n15367), .Z(
        P1_U3538) );
  MUX2_X1 U16889 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n15159), .S(n15354), .Z(
        P1_U3527) );
  MUX2_X1 U16890 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n15160), .S(n15354), .Z(
        P1_U3526) );
  MUX2_X1 U16891 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n15162), .S(n15354), .Z(
        P1_U3524) );
  INV_X1 U16892 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n15164) );
  MUX2_X1 U16893 ( .A(n15164), .B(n15163), .S(n15354), .Z(n15165) );
  INV_X1 U16894 ( .A(n15165), .ZN(P1_U3523) );
  MUX2_X1 U16895 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n15166), .S(n15354), .Z(
        P1_U3522) );
  MUX2_X1 U16896 ( .A(n15167), .B(P1_REG0_REG_25__SCAN_IN), .S(n15353), .Z(
        P1_U3521) );
  MUX2_X1 U16897 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n15169), .S(n15354), .Z(
        P1_U3519) );
  MUX2_X1 U16898 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n15170), .S(n15354), .Z(
        P1_U3518) );
  MUX2_X1 U16899 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n15171), .S(n15354), .Z(
        P1_U3517) );
  MUX2_X1 U16900 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n15172), .S(n15354), .Z(
        P1_U3516) );
  MUX2_X1 U16901 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n15173), .S(n15354), .Z(
        P1_U3515) );
  MUX2_X1 U16902 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n15174), .S(n15354), .Z(
        P1_U3513) );
  MUX2_X1 U16903 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n15175), .S(n15354), .Z(
        P1_U3510) );
  MUX2_X1 U16904 ( .A(n15176), .B(P1_REG0_REG_16__SCAN_IN), .S(n15353), .Z(
        P1_U3507) );
  MUX2_X1 U16905 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n15177), .S(n15354), .Z(
        P1_U3504) );
  MUX2_X1 U16906 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n15178), .S(n15354), .Z(
        P1_U3501) );
  MUX2_X1 U16907 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n15179), .S(n15354), .Z(
        P1_U3498) );
  MUX2_X1 U16908 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n15180), .S(n15354), .Z(
        P1_U3495) );
  MUX2_X1 U16909 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n15181), .S(n15354), .Z(
        P1_U3492) );
  NOR4_X1 U16910 ( .A1(n15182), .A2(P1_IR_REG_30__SCAN_IN), .A3(n15184), .A4(
        P1_U3086), .ZN(n15185) );
  AOI21_X1 U16911 ( .B1(n15186), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n15185), 
        .ZN(n15187) );
  OAI21_X1 U16912 ( .B1(n15188), .B2(n15195), .A(n15187), .ZN(P1_U3324) );
  OAI222_X1 U16913 ( .A1(P1_U3086), .A2(n8871), .B1(n15192), .B2(n15191), .C1(
        n15190), .C2(n15189), .ZN(P1_U3326) );
  OAI222_X1 U16914 ( .A1(n15189), .A2(n15196), .B1(n15195), .B2(n15194), .C1(
        P1_U3086), .C2(n15193), .ZN(P1_U3327) );
  MUX2_X1 U16915 ( .A(n15198), .B(n15197), .S(P1_U3086), .Z(P1_U3333) );
  MUX2_X1 U16916 ( .A(n15199), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  AOI21_X1 U16917 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n15203) );
  OAI21_X1 U16918 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n15203), 
        .ZN(U28) );
  AOI21_X1 U16919 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n15204) );
  OAI21_X1 U16920 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n15204), 
        .ZN(U29) );
  OAI21_X1 U16921 ( .B1(n15207), .B2(n15206), .A(n15205), .ZN(n15208) );
  XNOR2_X1 U16922 ( .A(n15208), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16923 ( .B1(n15211), .B2(n15210), .A(n15209), .ZN(SUB_1596_U57) );
  OAI21_X1 U16924 ( .B1(n15213), .B2(n15801), .A(n15212), .ZN(SUB_1596_U55) );
  OAI21_X1 U16925 ( .B1(n15216), .B2(n15215), .A(n15214), .ZN(n15217) );
  XNOR2_X1 U16926 ( .A(n15217), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(SUB_1596_U54)
         );
  OAI222_X1 U16927 ( .A1(n15431), .A2(n15220), .B1(n15431), .B2(n7624), .C1(
        n15219), .C2(n15218), .ZN(SUB_1596_U70) );
  OAI222_X1 U16928 ( .A1(n15501), .A2(n15222), .B1(n15501), .B2(n8790), .C1(
        n6826), .C2(n15221), .ZN(SUB_1596_U63) );
  OAI21_X1 U16929 ( .B1(n15225), .B2(n15224), .A(n15223), .ZN(n15226) );
  XNOR2_X1 U16930 ( .A(n15226), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI21_X1 U16931 ( .B1(n15228), .B2(n15445), .A(n15227), .ZN(SUB_1596_U68) );
  AOI21_X1 U16932 ( .B1(n15231), .B2(n15230), .A(n15229), .ZN(n15232) );
  XOR2_X1 U16933 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n15232), .Z(SUB_1596_U67)
         );
  OAI21_X1 U16934 ( .B1(n15234), .B2(n6580), .A(n15233), .ZN(n15235) );
  XNOR2_X1 U16935 ( .A(n15235), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  OAI222_X1 U16936 ( .A1(n15472), .A2(n15239), .B1(n15472), .B2(n15238), .C1(
        n15237), .C2(n15236), .ZN(SUB_1596_U65) );
  INV_X1 U16937 ( .A(n15242), .ZN(n15241) );
  OAI222_X1 U16938 ( .A1(n15485), .A2(n15243), .B1(n15485), .B2(n15242), .C1(
        n15241), .C2(n15240), .ZN(SUB_1596_U64) );
  OAI21_X1 U16939 ( .B1(P1_REG1_REG_0__SCAN_IN), .B2(n15245), .A(n15244), .ZN(
        n15246) );
  XOR2_X1 U16940 ( .A(P1_IR_REG_0__SCAN_IN), .B(n15246), .Z(n15250) );
  AOI22_X1 U16941 ( .A1(n15247), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n15248) );
  OAI21_X1 U16942 ( .B1(n15250), .B2(n15249), .A(n15248), .ZN(P1_U3243) );
  OAI21_X1 U16943 ( .B1(n15253), .B2(n15252), .A(n15251), .ZN(n15254) );
  XNOR2_X1 U16944 ( .A(n15256), .B(n15254), .ZN(n15290) );
  XNOR2_X1 U16945 ( .A(n15256), .B(n15255), .ZN(n15257) );
  NOR2_X1 U16946 ( .A1(n15257), .A2(n15296), .ZN(n15258) );
  AOI211_X1 U16947 ( .C1(n15348), .C2(n15290), .A(n15259), .B(n15258), .ZN(
        n15287) );
  AOI222_X1 U16948 ( .A1(P1_REG2_REG_2__SCAN_IN), .A2(n6408), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n15262), .C1(n15261), .C2(n15260), .ZN(
        n15271) );
  INV_X1 U16949 ( .A(n15263), .ZN(n15266) );
  OAI211_X1 U16950 ( .C1(n15286), .C2(n15266), .A(n15265), .B(n15264), .ZN(
        n15285) );
  INV_X1 U16951 ( .A(n15285), .ZN(n15267) );
  AOI22_X1 U16952 ( .A1(n15290), .A2(n15269), .B1(n15268), .B2(n15267), .ZN(
        n15270) );
  OAI211_X1 U16953 ( .C1(n6408), .C2(n15287), .A(n15271), .B(n15270), .ZN(
        P1_U3291) );
  AND2_X1 U16954 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15666), .ZN(P1_U3294) );
  AND2_X1 U16955 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15666), .ZN(P1_U3296) );
  AND2_X1 U16956 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15666), .ZN(P1_U3297) );
  AND2_X1 U16957 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15666), .ZN(P1_U3298) );
  AND2_X1 U16958 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15666), .ZN(P1_U3299) );
  AND2_X1 U16959 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15666), .ZN(P1_U3300) );
  INV_X1 U16960 ( .A(n15666), .ZN(n15272) );
  INV_X1 U16961 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n15802) );
  NOR2_X1 U16962 ( .A1(n15272), .A2(n15802), .ZN(P1_U3301) );
  INV_X1 U16963 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n15768) );
  NOR2_X1 U16964 ( .A1(n15272), .A2(n15768), .ZN(P1_U3302) );
  AND2_X1 U16965 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15666), .ZN(P1_U3303) );
  AND2_X1 U16966 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15666), .ZN(P1_U3304) );
  AND2_X1 U16967 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15666), .ZN(P1_U3305) );
  AND2_X1 U16968 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15666), .ZN(P1_U3306) );
  AND2_X1 U16969 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15666), .ZN(P1_U3307) );
  AND2_X1 U16970 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15666), .ZN(P1_U3308) );
  AND2_X1 U16971 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15666), .ZN(P1_U3309) );
  AND2_X1 U16972 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15666), .ZN(P1_U3310) );
  AND2_X1 U16973 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15666), .ZN(P1_U3311) );
  AND2_X1 U16974 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15666), .ZN(P1_U3312) );
  INV_X1 U16975 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n15805) );
  NOR2_X1 U16976 ( .A1(n15272), .A2(n15805), .ZN(P1_U3313) );
  AND2_X1 U16977 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15666), .ZN(P1_U3314) );
  AND2_X1 U16978 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15666), .ZN(P1_U3315) );
  AND2_X1 U16979 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15666), .ZN(P1_U3316) );
  AND2_X1 U16980 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15666), .ZN(P1_U3317) );
  INV_X1 U16981 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n15759) );
  NOR2_X1 U16982 ( .A1(n15272), .A2(n15759), .ZN(P1_U3318) );
  AND2_X1 U16983 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15666), .ZN(P1_U3319) );
  AND2_X1 U16984 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15666), .ZN(P1_U3320) );
  AND2_X1 U16985 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15666), .ZN(P1_U3321) );
  AND2_X1 U16986 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15666), .ZN(P1_U3322) );
  AND2_X1 U16987 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15666), .ZN(P1_U3323) );
  AOI21_X1 U16988 ( .B1(n15340), .B2(n15296), .A(n15273), .ZN(n15274) );
  AOI211_X1 U16989 ( .C1(n15277), .C2(n15276), .A(n15275), .B(n15274), .ZN(
        n15355) );
  AOI22_X1 U16990 ( .A1(n15354), .A2(n15355), .B1(n8899), .B2(n15353), .ZN(
        P1_U3459) );
  INV_X1 U16991 ( .A(n15278), .ZN(n15284) );
  OAI22_X1 U16992 ( .A1(n15281), .A2(n15280), .B1(n15279), .B2(n15344), .ZN(
        n15283) );
  AOI211_X1 U16993 ( .C1(n15284), .C2(n15327), .A(n15283), .B(n15282), .ZN(
        n15356) );
  AOI22_X1 U16994 ( .A1(n15354), .A2(n15356), .B1(n8879), .B2(n15353), .ZN(
        P1_U3462) );
  OAI21_X1 U16995 ( .B1(n15286), .B2(n15344), .A(n15285), .ZN(n15289) );
  INV_X1 U16996 ( .A(n15287), .ZN(n15288) );
  AOI211_X1 U16997 ( .C1(n15347), .C2(n15290), .A(n15289), .B(n15288), .ZN(
        n15357) );
  AOI22_X1 U16998 ( .A1(n15354), .A2(n15357), .B1(n8926), .B2(n15353), .ZN(
        P1_U3465) );
  OAI211_X1 U16999 ( .C1(n15293), .C2(n15344), .A(n15292), .B(n15291), .ZN(
        n15299) );
  OAI22_X1 U17000 ( .A1(n15297), .A2(n15296), .B1(n15295), .B2(n15294), .ZN(
        n15298) );
  AOI211_X1 U17001 ( .C1(n15347), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        n15358) );
  INV_X1 U17002 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n15301) );
  AOI22_X1 U17003 ( .A1(n15354), .A2(n15358), .B1(n15301), .B2(n15353), .ZN(
        P1_U3468) );
  NAND3_X1 U17004 ( .A1(n15303), .A2(n15327), .A3(n15302), .ZN(n15308) );
  NOR2_X1 U17005 ( .A1(n15305), .A2(n15304), .ZN(n15307) );
  NAND3_X1 U17006 ( .A1(n15308), .A2(n15307), .A3(n15306), .ZN(n15309) );
  AOI21_X1 U17007 ( .B1(n15311), .B2(n15310), .A(n15309), .ZN(n15359) );
  INV_X1 U17008 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n15312) );
  AOI22_X1 U17009 ( .A1(n15354), .A2(n15359), .B1(n15312), .B2(n15353), .ZN(
        P1_U3471) );
  AOI211_X1 U17010 ( .C1(n15318), .C2(n15348), .A(n15314), .B(n15313), .ZN(
        n15315) );
  INV_X1 U17011 ( .A(n15315), .ZN(n15316) );
  AOI211_X1 U17012 ( .C1(n15347), .C2(n15318), .A(n15317), .B(n15316), .ZN(
        n15361) );
  INV_X1 U17013 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n15319) );
  AOI22_X1 U17014 ( .A1(n15354), .A2(n15361), .B1(n15319), .B2(n15353), .ZN(
        P1_U3474) );
  NOR2_X1 U17015 ( .A1(n15321), .A2(n15320), .ZN(n15324) );
  NOR4_X1 U17016 ( .A1(n15325), .A2(n15324), .A3(n15323), .A4(n15322), .ZN(
        n15362) );
  INV_X1 U17017 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n15326) );
  AOI22_X1 U17018 ( .A1(n15354), .A2(n15362), .B1(n15326), .B2(n15353), .ZN(
        P1_U3477) );
  AND2_X1 U17019 ( .A1(n15328), .A2(n15327), .ZN(n15331) );
  OAI21_X1 U17020 ( .B1(n6410), .B2(n15344), .A(n15329), .ZN(n15330) );
  NOR3_X1 U17021 ( .A1(n15332), .A2(n15331), .A3(n15330), .ZN(n15363) );
  INV_X1 U17022 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n15333) );
  AOI22_X1 U17023 ( .A1(n15354), .A2(n15363), .B1(n15333), .B2(n15353), .ZN(
        P1_U3480) );
  AOI21_X1 U17024 ( .B1(n15336), .B2(n15335), .A(n15334), .ZN(n15337) );
  OAI211_X1 U17025 ( .C1(n15340), .C2(n15339), .A(n15338), .B(n15337), .ZN(
        n15341) );
  INV_X1 U17026 ( .A(n15341), .ZN(n15364) );
  INV_X1 U17027 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15342) );
  AOI22_X1 U17028 ( .A1(n15354), .A2(n15364), .B1(n15342), .B2(n15353), .ZN(
        P1_U3483) );
  OAI21_X1 U17029 ( .B1(n15345), .B2(n15344), .A(n15343), .ZN(n15346) );
  AOI21_X1 U17030 ( .B1(n15349), .B2(n15347), .A(n15346), .ZN(n15351) );
  NAND2_X1 U17031 ( .A1(n15349), .A2(n15348), .ZN(n15350) );
  INV_X1 U17032 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n15764) );
  AOI22_X1 U17033 ( .A1(n15354), .A2(n15366), .B1(n15764), .B2(n15353), .ZN(
        P1_U3486) );
  AOI22_X1 U17034 ( .A1(n15367), .A2(n15355), .B1(n8917), .B2(n15365), .ZN(
        P1_U3528) );
  AOI22_X1 U17035 ( .A1(n15367), .A2(n15356), .B1(n8878), .B2(n15365), .ZN(
        P1_U3529) );
  AOI22_X1 U17036 ( .A1(n15367), .A2(n15357), .B1(n8923), .B2(n15365), .ZN(
        P1_U3530) );
  AOI22_X1 U17037 ( .A1(n15367), .A2(n15358), .B1(n10252), .B2(n15365), .ZN(
        P1_U3531) );
  AOI22_X1 U17038 ( .A1(n15367), .A2(n15359), .B1(n8957), .B2(n15365), .ZN(
        P1_U3532) );
  INV_X1 U17039 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n15360) );
  AOI22_X1 U17040 ( .A1(n15367), .A2(n15361), .B1(n15360), .B2(n15365), .ZN(
        P1_U3533) );
  AOI22_X1 U17041 ( .A1(n15367), .A2(n15362), .B1(n9003), .B2(n15365), .ZN(
        P1_U3534) );
  AOI22_X1 U17042 ( .A1(n15367), .A2(n15363), .B1(n10467), .B2(n15365), .ZN(
        P1_U3535) );
  AOI22_X1 U17043 ( .A1(n15367), .A2(n15364), .B1(n10469), .B2(n15365), .ZN(
        P1_U3536) );
  AOI22_X1 U17044 ( .A1(n15367), .A2(n15366), .B1(n10471), .B2(n15365), .ZN(
        P1_U3537) );
  NOR2_X1 U17045 ( .A1(n15368), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U17046 ( .A1(n15368), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n15382) );
  OAI211_X1 U17047 ( .C1(n15371), .C2(n15370), .A(n15486), .B(n15369), .ZN(
        n15378) );
  INV_X1 U17048 ( .A(n15372), .ZN(n15374) );
  NAND2_X1 U17049 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15373) );
  NAND2_X1 U17050 ( .A1(n15374), .A2(n15373), .ZN(n15375) );
  NAND3_X1 U17051 ( .A1(n15460), .A2(n15376), .A3(n15375), .ZN(n15377) );
  OAI211_X1 U17052 ( .C1(n15468), .C2(n15379), .A(n15378), .B(n15377), .ZN(
        n15380) );
  INV_X1 U17053 ( .A(n15380), .ZN(n15381) );
  NAND2_X1 U17054 ( .A1(n15382), .A2(n15381), .ZN(P2_U3215) );
  INV_X1 U17055 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n15833) );
  OAI211_X1 U17056 ( .C1(n15385), .C2(n15384), .A(n15486), .B(n15383), .ZN(
        n15390) );
  OAI211_X1 U17057 ( .C1(n15388), .C2(n15387), .A(n15460), .B(n15386), .ZN(
        n15389) );
  OAI211_X1 U17058 ( .C1(n15468), .C2(n15391), .A(n15390), .B(n15389), .ZN(
        n15392) );
  INV_X1 U17059 ( .A(n15392), .ZN(n15394) );
  NAND2_X1 U17060 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3088), .ZN(n15393) );
  OAI211_X1 U17061 ( .C1(n15500), .C2(n15833), .A(n15394), .B(n15393), .ZN(
        P2_U3217) );
  OAI211_X1 U17062 ( .C1(n15397), .C2(n15396), .A(n15486), .B(n15395), .ZN(
        n15402) );
  OAI211_X1 U17063 ( .C1(n15400), .C2(n15399), .A(n15460), .B(n15398), .ZN(
        n15401) );
  OAI211_X1 U17064 ( .C1(n15468), .C2(n15403), .A(n15402), .B(n15401), .ZN(
        n15404) );
  INV_X1 U17065 ( .A(n15404), .ZN(n15406) );
  OAI211_X1 U17066 ( .C1(n15500), .C2(n15407), .A(n15406), .B(n15405), .ZN(
        P2_U3218) );
  OAI211_X1 U17067 ( .C1(n15409), .C2(n15408), .A(n6646), .B(n15460), .ZN(
        n15414) );
  OAI211_X1 U17068 ( .C1(n15412), .C2(n15411), .A(n15486), .B(n15410), .ZN(
        n15413) );
  OAI211_X1 U17069 ( .C1(n15468), .C2(n15415), .A(n15414), .B(n15413), .ZN(
        n15416) );
  INV_X1 U17070 ( .A(n15416), .ZN(n15418) );
  NAND2_X1 U17071 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n15417) );
  OAI211_X1 U17072 ( .C1(n15801), .C2(n15500), .A(n15418), .B(n15417), .ZN(
        P2_U3222) );
  OAI211_X1 U17073 ( .C1(n15421), .C2(n15420), .A(n15419), .B(n15486), .ZN(
        n15422) );
  INV_X1 U17074 ( .A(n15422), .ZN(n15427) );
  AOI211_X1 U17075 ( .C1(n15425), .C2(n15424), .A(n15492), .B(n15423), .ZN(
        n15426) );
  AOI211_X1 U17076 ( .C1(n7441), .C2(n15428), .A(n15427), .B(n15426), .ZN(
        n15430) );
  OAI211_X1 U17077 ( .C1(n15431), .C2(n15500), .A(n15430), .B(n15429), .ZN(
        P2_U3224) );
  INV_X1 U17078 ( .A(n15432), .ZN(n15434) );
  OAI21_X1 U17079 ( .B1(n15434), .B2(n15433), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15435) );
  OAI21_X1 U17080 ( .B1(P2_REG3_REG_12__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15435), .ZN(n15444) );
  OAI21_X1 U17081 ( .B1(n15438), .B2(n15437), .A(n15436), .ZN(n15442) );
  XNOR2_X1 U17082 ( .A(n15440), .B(n15439), .ZN(n15441) );
  AOI22_X1 U17083 ( .A1(n15442), .A2(n15460), .B1(n15486), .B2(n15441), .ZN(
        n15443) );
  OAI211_X1 U17084 ( .C1(n15445), .C2(n15500), .A(n15444), .B(n15443), .ZN(
        P2_U3226) );
  INV_X1 U17085 ( .A(n15446), .ZN(n15447) );
  AOI211_X1 U17086 ( .C1(n15450), .C2(n15449), .A(n15448), .B(n15447), .ZN(
        n15455) );
  AOI211_X1 U17087 ( .C1(n15453), .C2(n15452), .A(n15492), .B(n15451), .ZN(
        n15454) );
  AOI211_X1 U17088 ( .C1(n7441), .C2(n15456), .A(n15455), .B(n15454), .ZN(
        n15458) );
  NAND2_X1 U17089 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_U3088), .ZN(n15457)
         );
  OAI211_X1 U17090 ( .C1(n7313), .C2(n15500), .A(n15458), .B(n15457), .ZN(
        P2_U3227) );
  INV_X1 U17091 ( .A(n15459), .ZN(n15461) );
  OAI211_X1 U17092 ( .C1(P2_REG1_REG_15__SCAN_IN), .C2(n15462), .A(n15461), 
        .B(n15460), .ZN(n15466) );
  OAI211_X1 U17093 ( .C1(n15464), .C2(P2_REG2_REG_15__SCAN_IN), .A(n15463), 
        .B(n15486), .ZN(n15465) );
  OAI211_X1 U17094 ( .C1(n15468), .C2(n15467), .A(n15466), .B(n15465), .ZN(
        n15469) );
  INV_X1 U17095 ( .A(n15469), .ZN(n15471) );
  NAND2_X1 U17096 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3088), .ZN(n15470)
         );
  OAI211_X1 U17097 ( .C1(n15472), .C2(n15500), .A(n15471), .B(n15470), .ZN(
        P2_U3229) );
  OAI211_X1 U17098 ( .C1(n15475), .C2(n15474), .A(n15473), .B(n15486), .ZN(
        n15476) );
  INV_X1 U17099 ( .A(n15476), .ZN(n15481) );
  AOI211_X1 U17100 ( .C1(n15479), .C2(n15478), .A(n15492), .B(n15477), .ZN(
        n15480) );
  AOI211_X1 U17101 ( .C1(n7441), .C2(n15482), .A(n15481), .B(n15480), .ZN(
        n15484) );
  OAI211_X1 U17102 ( .C1(n15485), .C2(n15500), .A(n15484), .B(n15483), .ZN(
        P2_U3230) );
  OAI211_X1 U17103 ( .C1(n15489), .C2(n15488), .A(n15487), .B(n15486), .ZN(
        n15490) );
  INV_X1 U17104 ( .A(n15490), .ZN(n15496) );
  AOI211_X1 U17105 ( .C1(n15494), .C2(n15493), .A(n15492), .B(n15491), .ZN(
        n15495) );
  AOI211_X1 U17106 ( .C1(n7441), .C2(n15497), .A(n15496), .B(n15495), .ZN(
        n15499) );
  NAND2_X1 U17107 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3088), .ZN(n15498)
         );
  OAI211_X1 U17108 ( .C1(n15501), .C2(n15500), .A(n15499), .B(n15498), .ZN(
        P2_U3231) );
  AND2_X1 U17109 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15504), .ZN(P2_U3266) );
  INV_X1 U17110 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n15758) );
  NOR2_X1 U17111 ( .A1(n15503), .A2(n15758), .ZN(P2_U3267) );
  AND2_X1 U17112 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15504), .ZN(P2_U3268) );
  AND2_X1 U17113 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15504), .ZN(P2_U3269) );
  AND2_X1 U17114 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15504), .ZN(P2_U3270) );
  AND2_X1 U17115 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15504), .ZN(P2_U3271) );
  AND2_X1 U17116 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15504), .ZN(P2_U3272) );
  AND2_X1 U17117 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15504), .ZN(P2_U3273) );
  AND2_X1 U17118 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15504), .ZN(P2_U3274) );
  AND2_X1 U17119 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15504), .ZN(P2_U3275) );
  AND2_X1 U17120 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15504), .ZN(P2_U3276) );
  AND2_X1 U17121 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15504), .ZN(P2_U3277) );
  AND2_X1 U17122 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15504), .ZN(P2_U3278) );
  AND2_X1 U17123 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15504), .ZN(P2_U3279) );
  AND2_X1 U17124 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15504), .ZN(P2_U3280) );
  AND2_X1 U17125 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15504), .ZN(P2_U3281) );
  AND2_X1 U17126 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15504), .ZN(P2_U3282) );
  AND2_X1 U17127 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15504), .ZN(P2_U3283) );
  AND2_X1 U17128 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15504), .ZN(P2_U3284) );
  AND2_X1 U17129 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15504), .ZN(P2_U3285) );
  INV_X1 U17130 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n15750) );
  NOR2_X1 U17131 ( .A1(n15503), .A2(n15750), .ZN(P2_U3286) );
  AND2_X1 U17132 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15504), .ZN(P2_U3287) );
  AND2_X1 U17133 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15504), .ZN(P2_U3288) );
  AND2_X1 U17134 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15504), .ZN(P2_U3289) );
  AND2_X1 U17135 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15504), .ZN(P2_U3290) );
  AND2_X1 U17136 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15504), .ZN(P2_U3291) );
  AND2_X1 U17137 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15504), .ZN(P2_U3292) );
  AND2_X1 U17138 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15504), .ZN(P2_U3293) );
  AND2_X1 U17139 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15504), .ZN(P2_U3294) );
  AND2_X1 U17140 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15504), .ZN(P2_U3295) );
  AOI22_X1 U17141 ( .A1(n15507), .A2(n15506), .B1(n15505), .B2(n15509), .ZN(
        P2_U3416) );
  AOI21_X1 U17142 ( .B1(n15510), .B2(n15509), .A(n15508), .ZN(P2_U3417) );
  INV_X1 U17143 ( .A(n15524), .ZN(n15518) );
  OAI21_X1 U17144 ( .B1(n15512), .B2(n15518), .A(n15511), .ZN(n15515) );
  INV_X1 U17145 ( .A(n15513), .ZN(n15514) );
  AOI211_X1 U17146 ( .C1(n7492), .C2(n15516), .A(n15515), .B(n15514), .ZN(
        n15534) );
  AOI22_X1 U17147 ( .A1(n15533), .A2(n15534), .B1(n8033), .B2(n15531), .ZN(
        P2_U3436) );
  OAI21_X1 U17148 ( .B1(n7013), .B2(n15518), .A(n15517), .ZN(n15520) );
  AOI211_X1 U17149 ( .C1(n7492), .C2(n15521), .A(n15520), .B(n15519), .ZN(
        n15535) );
  AOI22_X1 U17150 ( .A1(n15533), .A2(n15535), .B1(n8078), .B2(n15531), .ZN(
        P2_U3442) );
  AND2_X1 U17151 ( .A1(n15523), .A2(n15522), .ZN(n15529) );
  NAND2_X1 U17152 ( .A1(n15525), .A2(n15524), .ZN(n15526) );
  NAND2_X1 U17153 ( .A1(n15527), .A2(n15526), .ZN(n15528) );
  NOR3_X1 U17154 ( .A1(n15530), .A2(n15529), .A3(n15528), .ZN(n15537) );
  INV_X1 U17155 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U17156 ( .A1(n15533), .A2(n15537), .B1(n15532), .B2(n15531), .ZN(
        P2_U3451) );
  AOI22_X1 U17157 ( .A1(n15538), .A2(n15534), .B1(n8034), .B2(n15536), .ZN(
        P2_U3501) );
  AOI22_X1 U17158 ( .A1(n15538), .A2(n15535), .B1(n8079), .B2(n15536), .ZN(
        P2_U3503) );
  AOI22_X1 U17159 ( .A1(n15538), .A2(n15537), .B1(n8133), .B2(n15536), .ZN(
        P2_U3506) );
  NOR2_X1 U17160 ( .A1(P3_U3897), .A2(n15539), .ZN(P3_U3150) );
  OAI21_X1 U17161 ( .B1(n15542), .B2(n15541), .A(n15540), .ZN(n15557) );
  NOR2_X1 U17162 ( .A1(n7617), .A2(n15544), .ZN(n15548) );
  INV_X1 U17163 ( .A(n15545), .ZN(n15546) );
  AOI21_X1 U17164 ( .B1(n15548), .B2(n15547), .A(n15546), .ZN(n15551) );
  OAI22_X1 U17165 ( .A1(n15551), .A2(n15570), .B1(n15550), .B2(n15549), .ZN(
        n15556) );
  XOR2_X1 U17166 ( .A(n15553), .B(n15552), .Z(n15554) );
  NOR2_X1 U17167 ( .A1(n15554), .A2(n15576), .ZN(n15555) );
  AOI211_X1 U17168 ( .C1(n15591), .C2(n15557), .A(n15556), .B(n15555), .ZN(
        n15559) );
  OAI211_X1 U17169 ( .C1(n15560), .C2(n15605), .A(n15559), .B(n15558), .ZN(
        P3_U3188) );
  INV_X1 U17170 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15582) );
  OAI21_X1 U17171 ( .B1(n15563), .B2(n15562), .A(n15561), .ZN(n15579) );
  XOR2_X1 U17172 ( .A(n15565), .B(n15564), .Z(n15577) );
  INV_X1 U17173 ( .A(n15566), .ZN(n15568) );
  NAND3_X1 U17174 ( .A1(n15569), .A2(n15568), .A3(n15567), .ZN(n15571) );
  AOI21_X1 U17175 ( .B1(n15572), .B2(n15571), .A(n15570), .ZN(n15573) );
  AOI21_X1 U17176 ( .B1(n15598), .B2(n15574), .A(n15573), .ZN(n15575) );
  OAI21_X1 U17177 ( .B1(n15577), .B2(n15576), .A(n15575), .ZN(n15578) );
  AOI21_X1 U17178 ( .B1(n15591), .B2(n15579), .A(n15578), .ZN(n15581) );
  OAI211_X1 U17179 ( .C1(n15582), .C2(n15605), .A(n15581), .B(n15580), .ZN(
        P3_U3190) );
  AND3_X1 U17180 ( .A1(n15585), .A2(n15584), .A3(n15583), .ZN(n15587) );
  OAI21_X1 U17181 ( .B1(n15588), .B2(n15587), .A(n15586), .ZN(n15602) );
  XNOR2_X1 U17182 ( .A(n15590), .B(n15589), .ZN(n15592) );
  NAND2_X1 U17183 ( .A1(n15592), .A2(n15591), .ZN(n15601) );
  XNOR2_X1 U17184 ( .A(n15594), .B(n15593), .ZN(n15596) );
  NAND2_X1 U17185 ( .A1(n15596), .A2(n15595), .ZN(n15600) );
  NAND2_X1 U17186 ( .A1(n15598), .A2(n15597), .ZN(n15599) );
  AND4_X1 U17187 ( .A1(n15602), .A2(n15601), .A3(n15600), .A4(n15599), .ZN(
        n15604) );
  OAI211_X1 U17188 ( .C1(n6684), .C2(n15605), .A(n15604), .B(n15603), .ZN(
        P3_U3192) );
  INV_X1 U17189 ( .A(n15606), .ZN(n15607) );
  OAI22_X1 U17190 ( .A1(n15610), .A2(n15609), .B1(n15608), .B2(n15607), .ZN(
        n15613) );
  INV_X1 U17191 ( .A(n15611), .ZN(n15612) );
  AOI211_X1 U17192 ( .C1(n15615), .C2(n15614), .A(n15613), .B(n15612), .ZN(
        n15617) );
  AOI22_X1 U17193 ( .A1(n15618), .A2(n10400), .B1(n15617), .B2(n15616), .ZN(
        P3_U3231) );
  AOI211_X1 U17194 ( .C1(n6643), .C2(n15621), .A(n15620), .B(n15619), .ZN(
        n15655) );
  AOI22_X1 U17195 ( .A1(n15654), .A2(n15655), .B1(n9503), .B2(n15653), .ZN(
        P3_U3393) );
  AOI22_X1 U17196 ( .A1(n15654), .A2(n15622), .B1(n9517), .B2(n15653), .ZN(
        P3_U3396) );
  AOI211_X1 U17197 ( .C1(n15625), .C2(n6643), .A(n15624), .B(n15623), .ZN(
        n15656) );
  AOI22_X1 U17198 ( .A1(n15654), .A2(n15656), .B1(n9595), .B2(n15653), .ZN(
        P3_U3399) );
  NOR2_X1 U17199 ( .A1(n15627), .A2(n15626), .ZN(n15629) );
  AOI211_X1 U17200 ( .C1(n15631), .C2(n15630), .A(n15629), .B(n15628), .ZN(
        n15658) );
  AOI22_X1 U17201 ( .A1(n15654), .A2(n15658), .B1(n9578), .B2(n15653), .ZN(
        P3_U3402) );
  INV_X1 U17202 ( .A(n15632), .ZN(n15636) );
  INV_X1 U17203 ( .A(n15633), .ZN(n15634) );
  AOI211_X1 U17204 ( .C1(n15636), .C2(n6643), .A(n15635), .B(n15634), .ZN(
        n15659) );
  AOI22_X1 U17205 ( .A1(n15654), .A2(n15659), .B1(n9563), .B2(n15653), .ZN(
        P3_U3405) );
  INV_X1 U17206 ( .A(n15637), .ZN(n15638) );
  AOI211_X1 U17207 ( .C1(n15640), .C2(n6643), .A(n15639), .B(n15638), .ZN(
        n15660) );
  AOI22_X1 U17208 ( .A1(n15654), .A2(n15660), .B1(n9538), .B2(n15653), .ZN(
        P3_U3408) );
  INV_X1 U17209 ( .A(n15641), .ZN(n15642) );
  AOI211_X1 U17210 ( .C1(n15644), .C2(n6643), .A(n15643), .B(n15642), .ZN(
        n15661) );
  AOI22_X1 U17211 ( .A1(n15654), .A2(n15661), .B1(n9623), .B2(n15653), .ZN(
        P3_U3411) );
  INV_X1 U17212 ( .A(n15645), .ZN(n15646) );
  AOI211_X1 U17213 ( .C1(n6643), .C2(n15648), .A(n15647), .B(n15646), .ZN(
        n15662) );
  AOI22_X1 U17214 ( .A1(n15654), .A2(n15662), .B1(n9648), .B2(n15653), .ZN(
        P3_U3414) );
  INV_X1 U17215 ( .A(n15649), .ZN(n15650) );
  AOI211_X1 U17216 ( .C1(n15652), .C2(n6643), .A(n15651), .B(n15650), .ZN(
        n15664) );
  AOI22_X1 U17217 ( .A1(n15654), .A2(n15664), .B1(n9671), .B2(n15653), .ZN(
        P3_U3417) );
  AOI22_X1 U17218 ( .A1(n15665), .A2(n15655), .B1(n10382), .B2(n15663), .ZN(
        P3_U3460) );
  AOI22_X1 U17219 ( .A1(n15665), .A2(n15656), .B1(n10390), .B2(n15663), .ZN(
        P3_U3462) );
  INV_X1 U17220 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15657) );
  AOI22_X1 U17221 ( .A1(n15665), .A2(n15658), .B1(n15657), .B2(n15663), .ZN(
        P3_U3463) );
  AOI22_X1 U17222 ( .A1(n15665), .A2(n15659), .B1(n9560), .B2(n15663), .ZN(
        P3_U3464) );
  AOI22_X1 U17223 ( .A1(n15665), .A2(n15660), .B1(n10686), .B2(n15663), .ZN(
        P3_U3465) );
  AOI22_X1 U17224 ( .A1(n15665), .A2(n15661), .B1(n9628), .B2(n15663), .ZN(
        P3_U3466) );
  AOI22_X1 U17225 ( .A1(n15665), .A2(n15662), .B1(n11223), .B2(n15663), .ZN(
        P3_U3467) );
  AOI22_X1 U17226 ( .A1(n15665), .A2(n15664), .B1(n9667), .B2(n15663), .ZN(
        P3_U3468) );
  NAND2_X1 U17227 ( .A1(n15666), .A2(P1_D_REG_30__SCAN_IN), .ZN(n15819) );
  NAND4_X1 U17228 ( .A1(P2_REG0_REG_21__SCAN_IN), .A2(n15765), .A3(n15667), 
        .A4(n15734), .ZN(n15672) );
  AND4_X1 U17229 ( .A1(n15751), .A2(n15769), .A3(P1_DATAO_REG_24__SCAN_IN), 
        .A4(P3_IR_REG_29__SCAN_IN), .ZN(n15669) );
  NAND4_X1 U17230 ( .A1(n15669), .A2(n15749), .A3(P3_DATAO_REG_17__SCAN_IN), 
        .A4(n15668), .ZN(n15671) );
  NAND4_X1 U17231 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P2_DATAO_REG_25__SCAN_IN), 
        .A3(n15764), .A4(n15775), .ZN(n15670) );
  NOR4_X1 U17232 ( .A1(n15672), .A2(n15671), .A3(P1_ADDR_REG_10__SCAN_IN), 
        .A4(n15670), .ZN(n15817) );
  NAND4_X1 U17233 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P3_ADDR_REG_4__SCAN_IN), 
        .A3(n15781), .A4(n15782), .ZN(n15689) );
  NOR4_X1 U17234 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), 
        .A3(P1_IR_REG_26__SCAN_IN), .A4(n8836), .ZN(n15676) );
  AND4_X1 U17235 ( .A1(n15695), .A2(n15696), .A3(SI_6_), .A4(
        P2_REG1_REG_4__SCAN_IN), .ZN(n15673) );
  NAND4_X1 U17236 ( .A1(n15676), .A2(n15675), .A3(n15674), .A4(n15673), .ZN(
        n15688) );
  NOR4_X1 U17237 ( .A1(P2_REG1_REG_0__SCAN_IN), .A2(P3_REG0_REG_9__SCAN_IN), 
        .A3(n15720), .A4(n8926), .ZN(n15681) );
  NOR4_X1 U17238 ( .A1(P3_IR_REG_30__SCAN_IN), .A2(P2_REG0_REG_9__SCAN_IN), 
        .A3(P3_REG1_REG_17__SCAN_IN), .A4(n15722), .ZN(n15677) );
  NAND4_X1 U17239 ( .A1(n15703), .A2(P3_REG1_REG_30__SCAN_IN), .A3(n15677), 
        .A4(P3_ADDR_REG_18__SCAN_IN), .ZN(n15679) );
  NAND4_X1 U17240 ( .A1(n15693), .A2(P2_REG1_REG_28__SCAN_IN), .A3(
        P2_DATAO_REG_0__SCAN_IN), .A4(P2_DATAO_REG_4__SCAN_IN), .ZN(n15678) );
  NOR3_X1 U17241 ( .A1(n15712), .A2(n15679), .A3(n15678), .ZN(n15680) );
  NAND2_X1 U17242 ( .A1(n15681), .A2(n15680), .ZN(n15687) );
  NAND4_X1 U17243 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15799), .A3(n9560), .A4(
        n15748), .ZN(n15685) );
  NAND4_X1 U17244 ( .A1(P2_REG2_REG_19__SCAN_IN), .A2(P2_REG2_REG_1__SCAN_IN), 
        .A3(P3_REG3_REG_22__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n15684)
         );
  NAND4_X1 U17245 ( .A1(P2_REG0_REG_20__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), 
        .A3(P1_D_REG_24__SCAN_IN), .A4(n15801), .ZN(n15683) );
  INV_X1 U17246 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n15790) );
  NAND4_X1 U17247 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(n15791), .A3(n15780), 
        .A4(n15790), .ZN(n15682) );
  OR4_X1 U17248 ( .A1(n15685), .A2(n15684), .A3(n15683), .A4(n15682), .ZN(
        n15686) );
  NOR4_X1 U17249 ( .A1(n15689), .A2(n15688), .A3(n15687), .A4(n15686), .ZN(
        n15816) );
  AOI22_X1 U17250 ( .A1(n15691), .A2(keyinput58), .B1(keyinput28), .B2(n8836), 
        .ZN(n15690) );
  OAI221_X1 U17251 ( .B1(n15691), .B2(keyinput58), .C1(n8836), .C2(keyinput28), 
        .A(n15690), .ZN(n15702) );
  AOI22_X1 U17252 ( .A1(n15693), .A2(keyinput43), .B1(keyinput30), .B2(n8821), 
        .ZN(n15692) );
  OAI221_X1 U17253 ( .B1(n15693), .B2(keyinput43), .C1(n8821), .C2(keyinput30), 
        .A(n15692), .ZN(n15701) );
  AOI22_X1 U17254 ( .A1(n15696), .A2(keyinput3), .B1(keyinput7), .B2(n15695), 
        .ZN(n15694) );
  OAI221_X1 U17255 ( .B1(n15696), .B2(keyinput3), .C1(n15695), .C2(keyinput7), 
        .A(n15694), .ZN(n15700) );
  XNOR2_X1 U17256 ( .A(SI_6_), .B(keyinput46), .ZN(n15698) );
  XNOR2_X1 U17257 ( .A(keyinput25), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n15697) );
  NAND2_X1 U17258 ( .A1(n15698), .A2(n15697), .ZN(n15699) );
  NOR4_X1 U17259 ( .A1(n15702), .A2(n15701), .A3(n15700), .A4(n15699), .ZN(
        n15746) );
  XOR2_X1 U17260 ( .A(P3_REG1_REG_30__SCAN_IN), .B(keyinput16), .Z(n15705) );
  XNOR2_X1 U17261 ( .A(n15703), .B(keyinput5), .ZN(n15704) );
  NOR2_X1 U17262 ( .A1(n15705), .A2(n15704), .ZN(n15709) );
  XNOR2_X1 U17263 ( .A(keyinput8), .B(P3_ADDR_REG_18__SCAN_IN), .ZN(n15708) );
  XNOR2_X1 U17264 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(keyinput20), .ZN(n15707)
         );
  XNOR2_X1 U17265 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput37), .ZN(n15706)
         );
  NAND4_X1 U17266 ( .A1(n15709), .A2(n15708), .A3(n15707), .A4(n15706), .ZN(
        n15716) );
  AOI22_X1 U17267 ( .A1(n15712), .A2(keyinput49), .B1(n15711), .B2(keyinput2), 
        .ZN(n15710) );
  OAI221_X1 U17268 ( .B1(n15712), .B2(keyinput49), .C1(n15711), .C2(keyinput2), 
        .A(n15710), .ZN(n15715) );
  XNOR2_X1 U17269 ( .A(n15713), .B(keyinput55), .ZN(n15714) );
  NOR3_X1 U17270 ( .A1(n15716), .A2(n15715), .A3(n15714), .ZN(n15745) );
  AOI22_X1 U17271 ( .A1(n9499), .A2(keyinput6), .B1(n15718), .B2(keyinput14), 
        .ZN(n15717) );
  OAI221_X1 U17272 ( .B1(n9499), .B2(keyinput6), .C1(n15718), .C2(keyinput14), 
        .A(n15717), .ZN(n15729) );
  AOI22_X1 U17273 ( .A1(n8926), .A2(keyinput4), .B1(n15720), .B2(keyinput0), 
        .ZN(n15719) );
  OAI221_X1 U17274 ( .B1(n8926), .B2(keyinput4), .C1(n15720), .C2(keyinput0), 
        .A(n15719), .ZN(n15728) );
  AOI22_X1 U17275 ( .A1(n15723), .A2(keyinput61), .B1(n15722), .B2(keyinput32), 
        .ZN(n15721) );
  OAI221_X1 U17276 ( .B1(n15723), .B2(keyinput61), .C1(n15722), .C2(keyinput32), .A(n15721), .ZN(n15727) );
  XOR2_X1 U17277 ( .A(n9671), .B(keyinput34), .Z(n15725) );
  XNOR2_X1 U17278 ( .A(P2_REG1_REG_0__SCAN_IN), .B(keyinput19), .ZN(n15724) );
  NAND2_X1 U17279 ( .A1(n15725), .A2(n15724), .ZN(n15726) );
  NOR4_X1 U17280 ( .A1(n15729), .A2(n15728), .A3(n15727), .A4(n15726), .ZN(
        n15744) );
  AOI22_X1 U17281 ( .A1(n15731), .A2(keyinput41), .B1(keyinput36), .B2(n8945), 
        .ZN(n15730) );
  OAI221_X1 U17282 ( .B1(n15731), .B2(keyinput41), .C1(n8945), .C2(keyinput36), 
        .A(n15730), .ZN(n15742) );
  AOI22_X1 U17283 ( .A1(n15734), .A2(keyinput52), .B1(n15733), .B2(keyinput35), 
        .ZN(n15732) );
  OAI221_X1 U17284 ( .B1(n15734), .B2(keyinput52), .C1(n15733), .C2(keyinput35), .A(n15732), .ZN(n15741) );
  XOR2_X1 U17285 ( .A(n15735), .B(keyinput40), .Z(n15739) );
  XNOR2_X1 U17286 ( .A(P2_REG3_REG_13__SCAN_IN), .B(keyinput9), .ZN(n15738) );
  XNOR2_X1 U17287 ( .A(P2_REG1_REG_12__SCAN_IN), .B(keyinput11), .ZN(n15737)
         );
  XNOR2_X1 U17288 ( .A(P3_IR_REG_29__SCAN_IN), .B(keyinput29), .ZN(n15736) );
  NAND4_X1 U17289 ( .A1(n15739), .A2(n15738), .A3(n15737), .A4(n15736), .ZN(
        n15740) );
  NOR3_X1 U17290 ( .A1(n15742), .A2(n15741), .A3(n15740), .ZN(n15743) );
  NAND4_X1 U17291 ( .A1(n15746), .A2(n15745), .A3(n15744), .A4(n15743), .ZN(
        n15815) );
  AOI22_X1 U17292 ( .A1(n15749), .A2(keyinput15), .B1(n15748), .B2(keyinput24), 
        .ZN(n15747) );
  OAI221_X1 U17293 ( .B1(n15749), .B2(keyinput15), .C1(n15748), .C2(keyinput24), .A(n15747), .ZN(n15754) );
  XNOR2_X1 U17294 ( .A(n15750), .B(keyinput1), .ZN(n15753) );
  XNOR2_X1 U17295 ( .A(n15751), .B(keyinput57), .ZN(n15752) );
  OR3_X1 U17296 ( .A1(n15754), .A2(n15753), .A3(n15752), .ZN(n15762) );
  AOI22_X1 U17297 ( .A1(n9560), .A2(keyinput60), .B1(keyinput21), .B2(n15756), 
        .ZN(n15755) );
  OAI221_X1 U17298 ( .B1(n9560), .B2(keyinput60), .C1(n15756), .C2(keyinput21), 
        .A(n15755), .ZN(n15761) );
  AOI22_X1 U17299 ( .A1(n15759), .A2(keyinput45), .B1(n15758), .B2(keyinput48), 
        .ZN(n15757) );
  OAI221_X1 U17300 ( .B1(n15759), .B2(keyinput45), .C1(n15758), .C2(keyinput48), .A(n15757), .ZN(n15760) );
  NOR3_X1 U17301 ( .A1(n15762), .A2(n15761), .A3(n15760), .ZN(n15813) );
  AOI22_X1 U17302 ( .A1(n15765), .A2(keyinput13), .B1(keyinput17), .B2(n15764), 
        .ZN(n15763) );
  OAI221_X1 U17303 ( .B1(n15765), .B2(keyinput13), .C1(n15764), .C2(keyinput17), .A(n15763), .ZN(n15773) );
  AOI22_X1 U17304 ( .A1(n15768), .A2(keyinput53), .B1(n15767), .B2(keyinput54), 
        .ZN(n15766) );
  OAI221_X1 U17305 ( .B1(n15768), .B2(keyinput53), .C1(n15767), .C2(keyinput54), .A(n15766), .ZN(n15772) );
  XNOR2_X1 U17306 ( .A(n15769), .B(keyinput18), .ZN(n15771) );
  XOR2_X1 U17307 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput51), .Z(n15770) );
  OR4_X1 U17308 ( .A1(n15773), .A2(n15772), .A3(n15771), .A4(n15770), .ZN(
        n15778) );
  XNOR2_X1 U17309 ( .A(n15774), .B(keyinput62), .ZN(n15777) );
  XNOR2_X1 U17310 ( .A(n15775), .B(keyinput31), .ZN(n15776) );
  NOR3_X1 U17311 ( .A1(n15778), .A2(n15777), .A3(n15776), .ZN(n15812) );
  AOI22_X1 U17312 ( .A1(n15781), .A2(keyinput39), .B1(n15780), .B2(keyinput63), 
        .ZN(n15779) );
  OAI221_X1 U17313 ( .B1(n15781), .B2(keyinput39), .C1(n15780), .C2(keyinput63), .A(n15779), .ZN(n15788) );
  XNOR2_X1 U17314 ( .A(n15782), .B(keyinput38), .ZN(n15787) );
  XNOR2_X1 U17315 ( .A(n15783), .B(keyinput47), .ZN(n15786) );
  XNOR2_X1 U17316 ( .A(n15784), .B(keyinput59), .ZN(n15785) );
  OR4_X1 U17317 ( .A1(n15788), .A2(n15787), .A3(n15786), .A4(n15785), .ZN(
        n15795) );
  AOI22_X1 U17318 ( .A1(n15791), .A2(keyinput23), .B1(keyinput12), .B2(n15790), 
        .ZN(n15789) );
  OAI221_X1 U17319 ( .B1(n15791), .B2(keyinput23), .C1(n15790), .C2(keyinput12), .A(n15789), .ZN(n15794) );
  XNOR2_X1 U17320 ( .A(n15792), .B(keyinput33), .ZN(n15793) );
  NOR3_X1 U17321 ( .A1(n15795), .A2(n15794), .A3(n15793), .ZN(n15811) );
  AOI22_X1 U17322 ( .A1(n15797), .A2(keyinput22), .B1(n13667), .B2(keyinput10), 
        .ZN(n15796) );
  OAI221_X1 U17323 ( .B1(n15797), .B2(keyinput22), .C1(n13667), .C2(keyinput10), .A(n15796), .ZN(n15809) );
  AOI22_X1 U17324 ( .A1(n15799), .A2(keyinput44), .B1(n6920), .B2(keyinput27), 
        .ZN(n15798) );
  OAI221_X1 U17325 ( .B1(n15799), .B2(keyinput44), .C1(n6920), .C2(keyinput27), 
        .A(n15798), .ZN(n15808) );
  AOI22_X1 U17326 ( .A1(n15802), .A2(keyinput56), .B1(keyinput50), .B2(n15801), 
        .ZN(n15800) );
  OAI221_X1 U17327 ( .B1(n15802), .B2(keyinput56), .C1(n15801), .C2(keyinput50), .A(n15800), .ZN(n15807) );
  AOI22_X1 U17328 ( .A1(n15805), .A2(keyinput26), .B1(n15804), .B2(keyinput42), 
        .ZN(n15803) );
  OAI221_X1 U17329 ( .B1(n15805), .B2(keyinput26), .C1(n15804), .C2(keyinput42), .A(n15803), .ZN(n15806) );
  NOR4_X1 U17330 ( .A1(n15809), .A2(n15808), .A3(n15807), .A4(n15806), .ZN(
        n15810) );
  NAND4_X1 U17331 ( .A1(n15813), .A2(n15812), .A3(n15811), .A4(n15810), .ZN(
        n15814) );
  AOI211_X1 U17332 ( .C1(n15817), .C2(n15816), .A(n15815), .B(n15814), .ZN(
        n15818) );
  XNOR2_X1 U17333 ( .A(n15819), .B(n15818), .ZN(P1_U3295) );
  AOI21_X1 U17334 ( .B1(n15822), .B2(n15821), .A(n15820), .ZN(SUB_1596_U59) );
  OAI21_X1 U17335 ( .B1(n15825), .B2(n15824), .A(n15823), .ZN(SUB_1596_U58) );
  XOR2_X1 U17336 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15826), .Z(SUB_1596_U53) );
  AOI21_X1 U17337 ( .B1(n15829), .B2(n15828), .A(n15827), .ZN(SUB_1596_U56) );
  AOI21_X1 U17338 ( .B1(n15832), .B2(n15831), .A(n15830), .ZN(n15834) );
  XNOR2_X1 U17339 ( .A(n15834), .B(n15833), .ZN(SUB_1596_U60) );
  AOI21_X1 U17340 ( .B1(n15837), .B2(n15836), .A(n15835), .ZN(SUB_1596_U5) );
  INV_X1 U7599 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n15784) );
  INV_X2 U7259 ( .A(n14526), .ZN(n14738) );
  CLKBUF_X1 U7157 ( .A(n6402), .Z(n13474) );
  CLKBUF_X1 U7161 ( .A(n9989), .Z(n7167) );
  NAND2_X2 U7176 ( .A1(n10307), .A2(n12205), .ZN(n10296) );
  NOR2_X2 U7224 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n7218) );
  CLKBUF_X1 U7256 ( .A(n9314), .Z(n9408) );
  CLKBUF_X1 U7850 ( .A(n9453), .Z(n6438) );
  AND4_X1 U9912 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(n13304)
         );
endmodule

