

module b20_C_AntiSAT_k_128_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, 
        ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, 
        ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, 
        ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, 
        ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, 
        U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, 
        P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, 
        P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, 
        P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, 
        P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, 
        P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, 
        P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, 
        P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, 
        P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, 
        P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, 
        P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, 
        P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, 
        P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, 
        P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, 
        P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, 
        P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, 
        P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, 
        P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, 
        P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, 
        P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, 
        P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, 
        P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, 
        P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, 
        P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, 
        P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, 
        P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, 
        P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, 
        P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, 
        P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, 
        P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, 
        P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, 
        P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, 
        P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, 
        P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, 
        P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, 
        P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, 
        P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, 
        P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, 
        P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, 
        P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, 
        P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, 
        P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285;

  AOI211_X1 U4832 ( .C1(n9862), .C2(n7871), .A(n9627), .B(n8235), .ZN(n7932)
         );
  CLKBUF_X2 U4833 ( .A(n8552), .Z(n4342) );
  AND4_X1 U4834 ( .A1(n6099), .A2(n6098), .A3(n6097), .A4(n6096), .ZN(n10154)
         );
  AND3_X2 U4835 ( .A1(n5215), .A2(n5214), .A3(n5213), .ZN(n7582) );
  CLKBUF_X2 U4836 ( .A(n6102), .Z(n6445) );
  CLKBUF_X2 U4837 ( .A(n5688), .Z(n4327) );
  INV_X1 U4838 ( .A(n6131), .ZN(n6110) );
  AND2_X1 U4839 ( .A1(n5511), .A2(n5510), .ZN(n5519) );
  XOR2_X1 U4840 ( .A(n6959), .B(n5551), .Z(n10100) );
  OR2_X1 U4841 ( .A1(n6350), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6362) );
  AND2_X1 U4842 ( .A1(n5459), .A2(n5447), .ZN(n5457) );
  INV_X2 U4843 ( .A(n6601), .ZN(n6746) );
  OR2_X1 U4844 ( .A1(n6522), .A2(n6969), .ZN(n6523) );
  AND2_X1 U4845 ( .A1(n8633), .A2(n8545), .ZN(n8548) );
  INV_X2 U4846 ( .A(n7213), .ZN(n8558) );
  BUF_X1 U4847 ( .A(n6133), .Z(n6442) );
  INV_X1 U4848 ( .A(n6139), .ZN(n6265) );
  INV_X1 U4849 ( .A(n8457), .ZN(n8458) );
  CLKBUF_X2 U4850 ( .A(n5182), .Z(n5343) );
  AND3_X1 U4851 ( .A1(n5190), .A2(n5189), .A3(n5188), .ZN(n10050) );
  AND2_X1 U4852 ( .A1(n8437), .A2(n8438), .ZN(n8830) );
  XNOR2_X1 U4853 ( .A(n5376), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6969) );
  BUF_X1 U4854 ( .A(n5531), .Z(n4329) );
  INV_X1 U4855 ( .A(n8558), .ZN(n8552) );
  AND2_X1 U4856 ( .A1(n7442), .A2(n7332), .ZN(n4326) );
  NOR2_X4 U4857 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P2_ADDR_REG_19__SCAN_IN), 
        .ZN(n9796) );
  NAND2_X2 U4858 ( .A1(n5017), .A2(n5016), .ZN(n5253) );
  OR2_X2 U4859 ( .A1(n5480), .A2(n4945), .ZN(n5461) );
  NAND3_X2 U4860 ( .A1(n7852), .A2(n7855), .A3(n7851), .ZN(n8029) );
  XNOR2_X2 U4861 ( .A(n5544), .B(n7550), .ZN(n7549) );
  NAND4_X2 U4862 ( .A1(n5681), .A2(n5680), .A3(n5679), .A4(n5678), .ZN(n9321)
         );
  NAND2_X2 U4863 ( .A1(n5261), .A2(n5260), .ZN(n9886) );
  AND2_X2 U4864 ( .A1(n4944), .A2(n4360), .ZN(n4687) );
  AND2_X2 U4865 ( .A1(n4944), .A2(n4941), .ZN(n5434) );
  INV_X2 U4866 ( .A(n5480), .ZN(n4944) );
  NOR2_X2 U4867 ( .A1(n8019), .A2(n4452), .ZN(n5494) );
  NOR2_X2 U4868 ( .A1(n9324), .A2(n7264), .ZN(n7258) );
  NAND2_X2 U4869 ( .A1(n6623), .A2(n6622), .ZN(n9856) );
  OAI211_X2 U4870 ( .C1(n6215), .C2(n6857), .A(n6123), .B(n6122), .ZN(n10145)
         );
  AND2_X2 U4871 ( .A1(n5457), .A2(n5448), .ZN(n5511) );
  NAND2_X2 U4873 ( .A1(n5239), .A2(n5238), .ZN(n5017) );
  OAI21_X2 U4874 ( .B1(n5233), .B2(n5232), .A(n5010), .ZN(n5239) );
  INV_X1 U4875 ( .A(n9322), .ZN(n4461) );
  NAND4_X2 U4876 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(n9322)
         );
  NAND2_X2 U4878 ( .A1(n8663), .A2(n8533), .ZN(n8583) );
  NAND2_X2 U4879 ( .A1(n7773), .A2(n7774), .ZN(n7852) );
  NAND2_X2 U4880 ( .A1(n4613), .A2(n5005), .ZN(n5233) );
  NAND2_X2 U4881 ( .A1(n9318), .A2(n7582), .ZN(n6036) );
  NAND2_X2 U4882 ( .A1(n5526), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5528) );
  OAI211_X1 U4883 ( .C1(n7210), .C2(n8504), .A(n7209), .B(n7208), .ZN(n4328)
         );
  AOI21_X2 U4884 ( .B1(n8606), .B2(n8607), .A(n8551), .ZN(n8555) );
  XNOR2_X2 U4885 ( .A(n5253), .B(n5244), .ZN(n6883) );
  NOR2_X2 U4886 ( .A1(n6788), .A2(n6789), .ZN(n6787) );
  XNOR2_X1 U4887 ( .A(n4826), .B(n5399), .ZN(n5531) );
  XNOR2_X1 U4888 ( .A(n6626), .B(n9186), .ZN(n9857) );
  AOI21_X1 U4889 ( .B1(P2_REG1_REG_10__SCAN_IN), .B2(n7898), .A(n7892), .ZN(
        n5548) );
  NAND2_X1 U4890 ( .A1(n5266), .A2(n5265), .ZN(n9872) );
  NAND2_X1 U4891 ( .A1(n9317), .A2(n7610), .ZN(n7605) );
  INV_X1 U4892 ( .A(n6075), .ZN(n5932) );
  NAND4_X1 U4893 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(n9318)
         );
  INV_X4 U4894 ( .A(n6545), .ZN(n4330) );
  CLKBUF_X2 U4895 ( .A(n5693), .Z(n5898) );
  INV_X2 U4896 ( .A(n7572), .ZN(n7264) );
  NAND2_X2 U4897 ( .A1(n6092), .A2(n6093), .ZN(n6149) );
  CLKBUF_X2 U4898 ( .A(n5756), .Z(n4338) );
  NAND2_X1 U4899 ( .A1(n5634), .A2(n5633), .ZN(n5693) );
  INV_X1 U4900 ( .A(n5442), .ZN(n5420) );
  INV_X1 U4901 ( .A(n4992), .ZN(n6100) );
  CLKBUF_X2 U4902 ( .A(n5533), .Z(n7425) );
  INV_X1 U4903 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7025) );
  INV_X2 U4904 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U4905 ( .A(n6718), .ZN(n9163) );
  NAND2_X1 U4906 ( .A1(n8577), .A2(n8865), .ZN(n8632) );
  AOI22_X1 U4907 ( .A1(n8777), .A2(n8776), .B1(n5610), .B2(n8775), .ZN(n8779)
         );
  OR2_X1 U4908 ( .A1(n8771), .A2(n8770), .ZN(n8776) );
  NAND2_X1 U4909 ( .A1(n4844), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4843) );
  INV_X1 U4910 ( .A(n5560), .ZN(n4842) );
  AND2_X1 U4911 ( .A1(n5558), .A2(n5557), .ZN(n5560) );
  AOI21_X1 U4912 ( .B1(n8223), .B2(n7985), .A(n7984), .ZN(n8090) );
  OAI21_X1 U4913 ( .B1(n8715), .B2(n4836), .A(n4835), .ZN(n8009) );
  AOI21_X1 U4914 ( .B1(n9899), .B2(P1_REG1_REG_11__SCAN_IN), .A(n9894), .ZN(
        n9906) );
  NAND2_X1 U4915 ( .A1(n5300), .A2(n5299), .ZN(n9628) );
  NAND2_X2 U4916 ( .A1(n5251), .A2(n5250), .ZN(n9862) );
  OR2_X1 U4917 ( .A1(n7952), .A2(n7881), .ZN(n7791) );
  NAND2_X1 U4918 ( .A1(n5243), .A2(n5242), .ZN(n7952) );
  NAND2_X1 U4919 ( .A1(n5683), .A2(n5682), .ZN(n7309) );
  AND2_X1 U4920 ( .A1(n7362), .A2(n5485), .ZN(n4952) );
  NOR2_X2 U4921 ( .A1(n8705), .A2(n6436), .ZN(n5610) );
  NAND2_X2 U4922 ( .A1(n7561), .A2(n10021), .ZN(n10023) );
  AND2_X1 U4923 ( .A1(n7367), .A2(n4395), .ZN(n5544) );
  NOR2_X1 U4924 ( .A1(n7377), .A2(n5479), .ZN(n7378) );
  AND2_X2 U4925 ( .A1(n4337), .A2(n8258), .ZN(n6557) );
  NAND2_X2 U4926 ( .A1(n7570), .A2(n7891), .ZN(n6075) );
  XNOR2_X1 U4927 ( .A(n4461), .B(n7436), .ZN(n5953) );
  NAND2_X2 U4928 ( .A1(n6524), .A2(n6523), .ZN(n6601) );
  AND2_X1 U4929 ( .A1(n7644), .A2(n6768), .ZN(n6524) );
  NAND4_X1 U4930 ( .A1(n5717), .A2(n5716), .A3(n5715), .A4(n5714), .ZN(n9317)
         );
  NAND2_X2 U4931 ( .A1(n6967), .A2(n6526), .ZN(n8258) );
  NAND4_X1 U4932 ( .A1(n5687), .A2(n5686), .A3(n5685), .A4(n5684), .ZN(n9320)
         );
  AOI21_X1 U4933 ( .B1(n7392), .B2(n7390), .A(n7391), .ZN(n7394) );
  INV_X2 U4934 ( .A(n6445), .ZN(n6318) );
  NAND2_X1 U4935 ( .A1(n6445), .A2(n6100), .ZN(n6215) );
  INV_X1 U4936 ( .A(n6484), .ZN(n8065) );
  AND2_X1 U4937 ( .A1(n6768), .A2(n6520), .ZN(n6549) );
  NAND2_X1 U4938 ( .A1(n5427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5425) );
  INV_X2 U4939 ( .A(n5688), .ZN(n5664) );
  CLKBUF_X2 U4940 ( .A(n5832), .Z(n4341) );
  AND2_X1 U4941 ( .A1(n6102), .A2(n6846), .ZN(n6139) );
  NAND2_X1 U4942 ( .A1(n5422), .A2(n5421), .ZN(n6484) );
  CLKBUF_X2 U4943 ( .A(n5832), .Z(n4340) );
  XNOR2_X1 U4944 ( .A(n5452), .B(n5451), .ZN(n8015) );
  NAND2_X1 U4945 ( .A1(n8510), .A2(n5612), .ZN(n6102) );
  BUF_X2 U4946 ( .A(n5756), .Z(n4339) );
  AND2_X1 U4947 ( .A1(n4743), .A2(n4742), .ZN(n5474) );
  NAND2_X1 U4948 ( .A1(n5520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U4949 ( .A1(n5444), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5441) );
  INV_X1 U4950 ( .A(n6092), .ZN(n8219) );
  NAND2_X1 U4951 ( .A1(n9153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6089) );
  MUX2_X1 U4952 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5138), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5140) );
  NAND2_X1 U4953 ( .A1(n5420), .A2(n5440), .ZN(n5444) );
  NOR2_X1 U4954 ( .A1(n6790), .A2(n4963), .ZN(n5536) );
  XNOR2_X1 U4955 ( .A(n5352), .B(n5351), .ZN(n7624) );
  OAI21_X1 U4956 ( .B1(n5367), .B2(n4462), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5138) );
  NAND2_X2 U4957 ( .A1(n6846), .A2(P1_U3086), .ZN(n9792) );
  NOR2_X1 U4958 ( .A1(n6791), .A2(n6792), .ZN(n6790) );
  OR2_X2 U4959 ( .A1(n6846), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9158) );
  AND2_X1 U4960 ( .A1(n5365), .A2(n4906), .ZN(n5356) );
  NOR2_X1 U4961 ( .A1(n5409), .A2(n4945), .ZN(n4940) );
  AND2_X1 U4962 ( .A1(n4904), .A2(n4903), .ZN(n4905) );
  NAND2_X1 U4963 ( .A1(n5476), .A2(n5401), .ZN(n5480) );
  NAND2_X2 U4964 ( .A1(n4974), .A2(n4973), .ZN(n4992) );
  AND3_X1 U4965 ( .A1(n5129), .A2(n5125), .A3(n5128), .ZN(n4904) );
  AND2_X2 U4966 ( .A1(n5173), .A2(n5124), .ZN(n5126) );
  NAND2_X1 U4967 ( .A1(n5451), .A2(n5450), .ZN(n5505) );
  INV_X1 U4968 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5351) );
  INV_X1 U4969 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5125) );
  INV_X1 U4970 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n7040) );
  AND2_X1 U4971 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n9795) );
  INV_X1 U4972 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5451) );
  NOR2_X1 U4973 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5130) );
  INV_X1 U4974 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5450) );
  NOR2_X1 U4975 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5128) );
  NOR2_X1 U4976 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5129) );
  INV_X2 U4977 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X2 U4978 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5173) );
  NOR2_X1 U4979 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n4519) );
  CLKBUF_X1 U4980 ( .A(n7227), .Z(n4331) );
  NAND3_X1 U4981 ( .A1(n7333), .A2(n4326), .A3(n4909), .ZN(n7443) );
  CLKBUF_X1 U4982 ( .A(n7773), .Z(n4332) );
  XNOR2_X1 U4983 ( .A(n5425), .B(P2_IR_REG_25__SCAN_IN), .ZN(n4333) );
  AOI21_X2 U4984 ( .B1(n8649), .B2(n8541), .A(n8540), .ZN(n4334) );
  NAND2_X1 U4986 ( .A1(n7335), .A2(n10133), .ZN(n4909) );
  NAND2_X2 U4987 ( .A1(n7334), .A2(n7482), .ZN(n7442) );
  XNOR2_X1 U4988 ( .A(n5425), .B(P2_IR_REG_25__SCAN_IN), .ZN(n6479) );
  AOI21_X1 U4989 ( .B1(n8649), .B2(n8541), .A(n8540), .ZN(n8542) );
  CLKBUF_X1 U4990 ( .A(n9328), .Z(n4336) );
  XNOR2_X1 U4991 ( .A(n10145), .B(n7213), .ZN(n7219) );
  NAND2_X2 U4992 ( .A1(n7772), .A2(n7771), .ZN(n7848) );
  NAND2_X2 U4993 ( .A1(n7672), .A2(n4925), .ZN(n7772) );
  NAND2_X2 U4994 ( .A1(n7520), .A2(n4926), .ZN(n7672) );
  NAND2_X2 U4995 ( .A1(n7445), .A2(n7444), .ZN(n7520) );
  XNOR2_X2 U4996 ( .A(n5187), .B(P1_IR_REG_2__SCAN_IN), .ZN(n9341) );
  NAND2_X1 U4997 ( .A1(n6524), .A2(n6523), .ZN(n4337) );
  NAND2_X2 U4998 ( .A1(n6477), .A2(n6476), .ZN(n6483) );
  AND2_X1 U4999 ( .A1(n5359), .A2(n8567), .ZN(n5756) );
  XNOR2_X2 U5000 ( .A(n7848), .B(n7849), .ZN(n7773) );
  NAND2_X1 U5001 ( .A1(n8567), .A2(n5634), .ZN(n5832) );
  OAI211_X2 U5002 ( .C1(n7210), .C2(n8504), .A(n7209), .B(n7208), .ZN(n7213)
         );
  NAND2_X2 U5003 ( .A1(n6485), .A2(n6897), .ZN(n7210) );
  AND2_X1 U5004 ( .A1(n5405), .A2(n4519), .ZN(n4518) );
  INV_X1 U5005 ( .A(n5023), .ZN(n5027) );
  OR2_X1 U5006 ( .A1(n9650), .A2(n9655), .ZN(n4599) );
  NAND2_X1 U5007 ( .A1(n4465), .A2(n5089), .ZN(n5152) );
  AOI21_X1 U5008 ( .B1(n4497), .B2(n4499), .A(n4375), .ZN(n4495) );
  AOI21_X1 U5009 ( .B1(n8467), .B2(n8466), .A(n8465), .ZN(n8470) );
  AND2_X1 U5010 ( .A1(n4577), .A2(n4394), .ZN(n4567) );
  NAND2_X1 U5011 ( .A1(n4545), .A2(n4368), .ZN(n8396) );
  AND2_X1 U5012 ( .A1(n4563), .A2(n8474), .ZN(n4557) );
  OR2_X1 U5013 ( .A1(n9650), .A2(n9196), .ZN(n6029) );
  NAND2_X1 U5014 ( .A1(n9437), .A2(n5941), .ZN(n4610) );
  AND2_X1 U5015 ( .A1(n4482), .A2(n4481), .ZN(n4480) );
  AND2_X1 U5016 ( .A1(n8642), .A2(n8535), .ZN(n4913) );
  AND2_X1 U5017 ( .A1(n4759), .A2(n4756), .ZN(n8459) );
  AOI21_X1 U5018 ( .B1(n4511), .B2(n8457), .A(n4760), .ZN(n4759) );
  NAND2_X1 U5019 ( .A1(n8501), .A2(n8466), .ZN(n4757) );
  OAI21_X1 U5020 ( .B1(n4707), .B2(n4706), .A(n6250), .ZN(n4705) );
  AND2_X1 U5021 ( .A1(n8074), .A2(n6227), .ZN(n4707) );
  OR2_X1 U5022 ( .A1(n7861), .A2(n7963), .ZN(n8373) );
  OR2_X1 U5023 ( .A1(n7776), .A2(n7774), .ZN(n8352) );
  AOI21_X1 U5024 ( .B1(n4712), .B2(n4711), .A(n4378), .ZN(n4710) );
  INV_X1 U5025 ( .A(n6394), .ZN(n4711) );
  OR2_X1 U5026 ( .A1(n9076), .A2(n8698), .ZN(n6404) );
  AOI21_X1 U5027 ( .B1(n4666), .B2(n4669), .A(n4664), .ZN(n4663) );
  INV_X1 U5028 ( .A(n8438), .ZN(n4664) );
  OR2_X1 U5029 ( .A1(n9076), .A2(n8855), .ZN(n8434) );
  OR2_X1 U5030 ( .A1(n9090), .A2(n8854), .ZN(n8427) );
  OAI21_X1 U5031 ( .B1(n7704), .B2(n6180), .A(n6179), .ZN(n7730) );
  XNOR2_X1 U5032 ( .A(n4825), .B(n9186), .ZN(n6533) );
  OAI21_X1 U5033 ( .B1(n6557), .B2(n7436), .A(n6527), .ZN(n4825) );
  INV_X1 U5034 ( .A(n6067), .ZN(n6074) );
  OR2_X1 U5035 ( .A1(n9493), .A2(n9252), .ZN(n8312) );
  NAND2_X1 U5036 ( .A1(n9762), .A2(n8286), .ZN(n4862) );
  OR2_X1 U5037 ( .A1(n9697), .A2(n9177), .ZN(n5862) );
  INV_X1 U5038 ( .A(n4898), .ZN(n4897) );
  NAND2_X1 U5039 ( .A1(n8192), .A2(n8193), .ZN(n4902) );
  AND2_X1 U5040 ( .A1(n8129), .A2(n6045), .ZN(n4635) );
  NAND2_X1 U5041 ( .A1(n4500), .A2(n4410), .ZN(n5078) );
  OAI21_X1 U5042 ( .B1(n5324), .B2(n5321), .A(n5059), .ZN(n5061) );
  AOI21_X1 U5043 ( .B1(n4489), .B2(n4353), .A(n4488), .ZN(n4487) );
  INV_X1 U5044 ( .A(n5048), .ZN(n4488) );
  OAI21_X1 U5045 ( .B1(n5284), .B2(n4405), .A(n5038), .ZN(n5291) );
  XNOR2_X1 U5046 ( .A(n5032), .B(SI_13_), .ZN(n5267) );
  AOI21_X1 U5047 ( .B1(n4763), .B2(n4343), .A(n4379), .ZN(n4761) );
  NAND2_X1 U5048 ( .A1(n9795), .A2(n4972), .ZN(n4973) );
  NAND2_X1 U5049 ( .A1(n9796), .A2(n4439), .ZN(n4974) );
  INV_X1 U5050 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4972) );
  AND2_X1 U5051 ( .A1(n7673), .A2(n7671), .ZN(n4925) );
  AND2_X1 U5052 ( .A1(n8662), .A2(n8532), .ZN(n8533) );
  OAI21_X1 U5053 ( .B1(n4352), .B2(n4922), .A(n4921), .ZN(n4920) );
  AND2_X1 U5054 ( .A1(n8570), .A2(n8560), .ZN(n4922) );
  NAND2_X1 U5055 ( .A1(n4352), .A2(n8560), .ZN(n4921) );
  INV_X1 U5056 ( .A(n10145), .ZN(n7225) );
  AND2_X1 U5057 ( .A1(n8173), .A2(n8070), .ZN(n8071) );
  NAND3_X1 U5058 ( .A1(n6136), .A2(n4354), .A3(n6135), .ZN(n4530) );
  NAND2_X1 U5059 ( .A1(n8452), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6127) );
  AOI21_X1 U5060 ( .B1(n8821), .B2(n6466), .A(n6465), .ZN(n8467) );
  OR2_X1 U5061 ( .A1(n8706), .A2(n10184), .ZN(n8368) );
  XNOR2_X1 U5062 ( .A(n9064), .B(n8697), .ZN(n8822) );
  INV_X1 U5063 ( .A(n10130), .ZN(n10155) );
  INV_X1 U5064 ( .A(n10135), .ZN(n10153) );
  OR2_X1 U5065 ( .A1(n8657), .A2(n8959), .ZN(n8924) );
  NAND2_X1 U5066 ( .A1(n6510), .A2(n8471), .ZN(n10135) );
  NAND2_X1 U5067 ( .A1(n4565), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6091) );
  MUX2_X1 U5068 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5443), .S(
        P2_IR_REG_27__SCAN_IN), .Z(n5445) );
  OR2_X1 U5069 ( .A1(n5348), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n5347) );
  INV_X1 U5070 ( .A(n4341), .ZN(n5934) );
  NAND2_X1 U5071 ( .A1(n5359), .A2(n5633), .ZN(n5688) );
  NOR2_X1 U5072 ( .A1(n4597), .A2(n9432), .ZN(n4596) );
  NAND2_X1 U5073 ( .A1(n4598), .A2(n9741), .ZN(n4597) );
  INV_X1 U5074 ( .A(n4599), .ZN(n4598) );
  NAND2_X1 U5075 ( .A1(n4873), .A2(n4871), .ZN(n9450) );
  AND2_X1 U5076 ( .A1(n4872), .A2(n4399), .ZN(n4871) );
  AOI21_X1 U5077 ( .B1(n4344), .B2(n4625), .A(n4620), .ZN(n4619) );
  INV_X1 U5078 ( .A(n8313), .ZN(n4620) );
  AND2_X1 U5079 ( .A1(n5979), .A2(n8314), .ZN(n9453) );
  NAND2_X1 U5080 ( .A1(n4874), .A2(n4878), .ZN(n9485) );
  OR2_X1 U5081 ( .A1(n8306), .A2(n9568), .ZN(n8308) );
  NAND2_X1 U5082 ( .A1(n9635), .A2(n9634), .ZN(n4630) );
  NAND2_X1 U5083 ( .A1(n5305), .A2(n5304), .ZN(n9610) );
  XNOR2_X1 U5084 ( .A(n5340), .B(n5341), .ZN(n8212) );
  INV_X1 U5085 ( .A(n8697), .ZN(n8837) );
  CLKBUF_X1 U5086 ( .A(n6467), .Z(n5529) );
  OAI21_X1 U5087 ( .B1(n5777), .B2(n5776), .A(n7791), .ZN(n5778) );
  AND2_X1 U5088 ( .A1(n6042), .A2(n6000), .ZN(n4445) );
  INV_X1 U5089 ( .A(n5946), .ZN(n4443) );
  NAND2_X1 U5090 ( .A1(n4550), .A2(n4549), .ZN(n4548) );
  NOR2_X1 U5091 ( .A1(n8358), .A2(n8457), .ZN(n4549) );
  NAND2_X1 U5092 ( .A1(n8359), .A2(n8375), .ZN(n4550) );
  NAND2_X1 U5093 ( .A1(n4553), .A2(n4552), .ZN(n4551) );
  NOR2_X1 U5094 ( .A1(n8374), .A2(n8458), .ZN(n4552) );
  NAND2_X1 U5095 ( .A1(n8376), .A2(n8375), .ZN(n4553) );
  AND2_X1 U5096 ( .A1(n4568), .A2(n8406), .ZN(n4573) );
  OAI21_X1 U5097 ( .B1(n4571), .B2(n4570), .A(n4566), .ZN(n4569) );
  NOR2_X1 U5098 ( .A1(n4577), .A2(n8408), .ZN(n4571) );
  OAI21_X1 U5099 ( .B1(n4567), .B2(n4575), .A(n4753), .ZN(n4566) );
  NOR2_X1 U5100 ( .A1(n8405), .A2(n8457), .ZN(n4750) );
  NAND2_X1 U5101 ( .A1(n4771), .A2(n8457), .ZN(n4770) );
  AOI21_X1 U5102 ( .B1(n8414), .B2(n4532), .A(n4531), .ZN(n4771) );
  NOR2_X1 U5103 ( .A1(n4534), .A2(n4533), .ZN(n4532) );
  NAND2_X1 U5104 ( .A1(n8914), .A2(n8409), .ZN(n4531) );
  OAI21_X1 U5105 ( .B1(n4355), .B2(n4560), .A(n4556), .ZN(n4555) );
  NOR2_X1 U5106 ( .A1(n4563), .A2(n4561), .ZN(n4560) );
  NOR2_X1 U5107 ( .A1(n4558), .A2(n4557), .ZN(n4556) );
  AND2_X1 U5108 ( .A1(n8842), .A2(n8433), .ZN(n4754) );
  INV_X1 U5109 ( .A(n8439), .ZN(n4450) );
  AOI21_X1 U5110 ( .B1(n4507), .B2(n4510), .A(n4506), .ZN(n4505) );
  INV_X1 U5111 ( .A(n5341), .ZN(n4506) );
  OAI21_X1 U5112 ( .B1(n8447), .B2(n8697), .A(n8464), .ZN(n4511) );
  INV_X1 U5113 ( .A(n5552), .ZN(n4829) );
  NAND2_X1 U5114 ( .A1(n4718), .A2(n8954), .ZN(n4716) );
  NOR2_X1 U5115 ( .A1(n4676), .A2(n6456), .ZN(n4675) );
  INV_X1 U5116 ( .A(n8382), .ZN(n4676) );
  AND2_X1 U5117 ( .A1(n5977), .A2(n5976), .ZN(n6027) );
  NAND2_X1 U5118 ( .A1(n9432), .A2(n5932), .ZN(n4471) );
  NAND2_X1 U5119 ( .A1(n4470), .A2(n4469), .ZN(n4475) );
  NAND2_X1 U5120 ( .A1(n4472), .A2(n6075), .ZN(n4469) );
  NAND2_X1 U5121 ( .A1(n5939), .A2(n9432), .ZN(n4470) );
  INV_X1 U5122 ( .A(n4794), .ZN(n4789) );
  NAND2_X1 U5123 ( .A1(n4610), .A2(n4612), .ZN(n4609) );
  NAND2_X1 U5124 ( .A1(n8316), .A2(n4610), .ZN(n4607) );
  AND2_X1 U5125 ( .A1(n4764), .A2(n5262), .ZN(n4763) );
  OR2_X1 U5126 ( .A1(n4343), .A2(n4765), .ZN(n4764) );
  NAND2_X1 U5127 ( .A1(n5020), .A2(n5019), .ZN(n5023) );
  NAND2_X1 U5128 ( .A1(n5013), .A2(n5012), .ZN(n5016) );
  OR2_X1 U5129 ( .A1(n8057), .A2(n8174), .ZN(n8381) );
  NOR2_X1 U5130 ( .A1(n8483), .A2(n4685), .ZN(n4684) );
  INV_X1 U5131 ( .A(n8368), .ZN(n4685) );
  INV_X1 U5132 ( .A(n7478), .ZN(n4695) );
  INV_X1 U5133 ( .A(n4699), .ZN(n4696) );
  NAND2_X1 U5134 ( .A1(n7482), .A2(n4700), .ZN(n4699) );
  INV_X1 U5135 ( .A(n10177), .ZN(n4700) );
  NAND2_X1 U5136 ( .A1(n10133), .A2(n10177), .ZN(n4698) );
  NAND2_X1 U5137 ( .A1(n7352), .A2(n10154), .ZN(n8333) );
  INV_X1 U5138 ( .A(n4666), .ZN(n4665) );
  OR2_X1 U5139 ( .A1(n9070), .A2(n8826), .ZN(n8437) );
  INV_X1 U5140 ( .A(n8431), .ZN(n4670) );
  OR2_X1 U5141 ( .A1(n9103), .A2(n6346), .ZN(n8420) );
  AND2_X1 U5142 ( .A1(n8944), .A2(n6307), .ZN(n4718) );
  NOR2_X1 U5143 ( .A1(n4649), .A2(n8403), .ZN(n4648) );
  INV_X1 U5144 ( .A(n4651), .ZN(n4649) );
  NOR2_X1 U5145 ( .A1(n6457), .A2(n4655), .ZN(n4654) );
  INV_X1 U5146 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5415) );
  AND2_X1 U5147 ( .A1(n5407), .A2(n5406), .ZN(n4521) );
  INV_X1 U5148 ( .A(n5505), .ZN(n4523) );
  INV_X1 U5149 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4946) );
  AND2_X1 U5150 ( .A1(n6698), .A2(n6697), .ZN(n6706) );
  INV_X1 U5151 ( .A(n8567), .ZN(n5633) );
  OR2_X1 U5152 ( .A1(n9655), .A2(n9189), .ZN(n6023) );
  NOR2_X1 U5153 ( .A1(n4882), .A2(n8291), .ZN(n4881) );
  NOR2_X1 U5154 ( .A1(n9502), .A2(n9299), .ZN(n8291) );
  INV_X1 U5155 ( .A(n4891), .ZN(n4882) );
  INV_X1 U5156 ( .A(n8309), .ZN(n4639) );
  AND2_X1 U5157 ( .A1(n9540), .A2(n8307), .ZN(n4640) );
  INV_X1 U5158 ( .A(n4860), .ZN(n4858) );
  INV_X1 U5159 ( .A(n5658), .ZN(n5628) );
  INV_X1 U5160 ( .A(n4629), .ZN(n4628) );
  INV_X1 U5161 ( .A(n4896), .ZN(n4895) );
  OAI21_X1 U5162 ( .B1(n4899), .B2(n4897), .A(n8275), .ZN(n4896) );
  NOR2_X1 U5163 ( .A1(n4595), .A2(n9872), .ZN(n4594) );
  OR2_X1 U5164 ( .A1(n9862), .A2(n8230), .ZN(n6000) );
  NAND2_X1 U5165 ( .A1(n7582), .A2(n7610), .ZN(n4592) );
  OR2_X1 U5166 ( .A1(n9317), .A2(n7610), .ZN(n7633) );
  OR2_X1 U5167 ( .A1(n9655), .A2(n9295), .ZN(n8295) );
  INV_X1 U5168 ( .A(n9749), .ZN(n9493) );
  NAND2_X1 U5169 ( .A1(n5113), .A2(n5112), .ZN(n5146) );
  OR2_X1 U5170 ( .A1(n5111), .A2(n5110), .ZN(n5112) );
  OR2_X1 U5171 ( .A1(n5149), .A2(n5109), .ZN(n5113) );
  NAND2_X1 U5172 ( .A1(n5137), .A2(n4584), .ZN(n4583) );
  INV_X1 U5173 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4584) );
  NAND2_X1 U5174 ( .A1(n4466), .A2(n5083), .ZN(n5157) );
  AND2_X1 U5175 ( .A1(n5077), .A2(n5076), .ZN(n5160) );
  NAND2_X1 U5176 ( .A1(n4479), .A2(n4477), .ZN(n5324) );
  AND2_X1 U5177 ( .A1(n4478), .A2(n5058), .ZN(n4477) );
  NOR2_X1 U5178 ( .A1(n5301), .A2(n4490), .ZN(n4489) );
  INV_X1 U5179 ( .A(n5041), .ZN(n4490) );
  NAND2_X1 U5180 ( .A1(n5010), .A2(n5009), .ZN(n5232) );
  INV_X1 U5181 ( .A(SI_4_), .ZN(n7058) );
  OAI21_X1 U5182 ( .B1(n4992), .B2(P1_DATAO_REG_1__SCAN_IN), .A(n4978), .ZN(
        n4979) );
  NAND2_X1 U5183 ( .A1(n4992), .A2(n4977), .ZN(n4978) );
  INV_X1 U5184 ( .A(n10193), .ZN(n7776) );
  XNOR2_X1 U5185 ( .A(n7352), .B(n4328), .ZN(n7211) );
  NAND2_X1 U5186 ( .A1(n8534), .A2(n8918), .ZN(n8535) );
  OR2_X1 U5187 ( .A1(n8583), .A2(n4948), .ZN(n4914) );
  OR2_X1 U5188 ( .A1(n6149), .A2(n4537), .ZN(n6364) );
  OR2_X1 U5189 ( .A1(n6149), .A2(n4543), .ZN(n6421) );
  OR2_X1 U5190 ( .A1(n6149), .A2(n4539), .ZN(n6389) );
  INV_X1 U5191 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n4539) );
  AND4_X1 U5192 ( .A1(n6225), .A2(n6224), .A3(n6223), .A4(n6222), .ZN(n8075)
         );
  NAND2_X1 U5193 ( .A1(n7361), .A2(n4730), .ZN(n7377) );
  NAND2_X1 U5194 ( .A1(n7830), .A2(n7831), .ZN(n7829) );
  OR2_X1 U5195 ( .A1(n7827), .A2(n10237), .ZN(n4833) );
  OAI21_X1 U5196 ( .B1(n7824), .B2(n4739), .A(n4738), .ZN(n7902) );
  NAND2_X1 U5197 ( .A1(n4740), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U5198 ( .A1(n5488), .A2(n4740), .ZN(n4738) );
  XNOR2_X1 U5199 ( .A(n5548), .B(n8714), .ZN(n8715) );
  NAND2_X1 U5200 ( .A1(n10113), .A2(n10114), .ZN(n10112) );
  OR2_X1 U5201 ( .A1(n8727), .A2(n8728), .ZN(n4737) );
  NAND2_X1 U5202 ( .A1(n8752), .A2(n8753), .ZN(n8751) );
  NAND2_X1 U5203 ( .A1(n8783), .A2(n8782), .ZN(n8787) );
  OR2_X1 U5204 ( .A1(n6418), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8807) );
  NAND2_X1 U5205 ( .A1(n6386), .A2(n6385), .ZN(n6397) );
  INV_X1 U5206 ( .A(n6387), .ZN(n6386) );
  OR2_X1 U5207 ( .A1(n6362), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6375) );
  OR2_X1 U5208 ( .A1(n6333), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6342) );
  OR2_X1 U5209 ( .A1(n6311), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U5210 ( .A1(n8957), .A2(n4575), .ZN(n4719) );
  OR2_X1 U5211 ( .A1(n6288), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U5212 ( .B1(n6228), .B2(n4706), .A(n4704), .ZN(n6252) );
  INV_X1 U5213 ( .A(n4705), .ZN(n4704) );
  INV_X1 U5214 ( .A(n8378), .ZN(n4678) );
  NAND2_X1 U5215 ( .A1(n6228), .A2(n4707), .ZN(n7973) );
  OAI21_X1 U5216 ( .B1(n6193), .B2(n4722), .A(n4720), .ZN(n7962) );
  INV_X1 U5217 ( .A(n4721), .ZN(n4720) );
  OAI22_X1 U5218 ( .A1(n4723), .A2(n4722), .B1(n7861), .B2(n8702), .ZN(n4721)
         );
  NAND2_X1 U5219 ( .A1(n4382), .A2(n6204), .ZN(n4722) );
  NAND2_X1 U5220 ( .A1(n7702), .A2(n7701), .ZN(n4686) );
  NAND2_X1 U5221 ( .A1(n8350), .A2(n7685), .ZN(n8483) );
  NAND2_X1 U5222 ( .A1(n4686), .A2(n4684), .ZN(n7729) );
  NAND2_X1 U5223 ( .A1(n6144), .A2(n6143), .ZN(n7492) );
  NAND2_X1 U5224 ( .A1(n10151), .A2(n8335), .ZN(n4688) );
  OR2_X1 U5225 ( .A1(n6445), .A2(n4329), .ZN(n6123) );
  NAND2_X1 U5226 ( .A1(n4709), .A2(n4708), .ZN(n8823) );
  AOI21_X1 U5227 ( .B1(n4710), .B2(n4713), .A(n4370), .ZN(n4708) );
  AOI21_X1 U5228 ( .B1(n4668), .B2(n6463), .A(n4667), .ZN(n4666) );
  INV_X1 U5229 ( .A(n8434), .ZN(n4667) );
  NAND2_X1 U5230 ( .A1(n6462), .A2(n8427), .ZN(n8858) );
  INV_X1 U5231 ( .A(n4691), .ZN(n4690) );
  OAI21_X1 U5232 ( .B1(n6359), .B2(n4692), .A(n6370), .ZN(n4691) );
  NAND2_X1 U5233 ( .A1(n6358), .A2(n8496), .ZN(n8887) );
  NAND2_X1 U5234 ( .A1(n4681), .A2(n8415), .ZN(n8912) );
  NAND2_X1 U5235 ( .A1(n4971), .A2(n8412), .ZN(n4681) );
  NAND2_X1 U5236 ( .A1(n4719), .A2(n4718), .ZN(n8937) );
  NAND2_X1 U5237 ( .A1(n6309), .A2(n6308), .ZN(n8657) );
  AND2_X1 U5238 ( .A1(n8401), .A2(n6458), .ZN(n8493) );
  AOI21_X1 U5239 ( .B1(n4654), .B2(n8393), .A(n4652), .ZN(n4651) );
  INV_X1 U5240 ( .A(n8398), .ZN(n4652) );
  INV_X1 U5241 ( .A(n4654), .ZN(n4653) );
  INV_X1 U5242 ( .A(n9149), .ZN(n7010) );
  AND2_X1 U5243 ( .A1(n4523), .A2(n4521), .ZN(n4520) );
  INV_X1 U5244 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5503) );
  INV_X1 U5245 ( .A(n6583), .ZN(n4798) );
  NAND2_X1 U5246 ( .A1(n6583), .A2(n6582), .ZN(n7529) );
  OR2_X1 U5247 ( .A1(n5875), .A2(n5630), .ZN(n5888) );
  INV_X1 U5248 ( .A(n9248), .ZN(n6735) );
  XNOR2_X1 U5249 ( .A(n6560), .B(n9186), .ZN(n6570) );
  AOI21_X1 U5250 ( .B1(n4810), .B2(n4812), .A(n4813), .ZN(n4805) );
  NAND2_X1 U5251 ( .A1(n9170), .A2(n4814), .ZN(n4813) );
  INV_X1 U5252 ( .A(n9869), .ZN(n4784) );
  NAND2_X1 U5253 ( .A1(n5626), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5844) );
  INV_X1 U5254 ( .A(n5834), .ZN(n5626) );
  INV_X1 U5255 ( .A(n8166), .ZN(n4803) );
  AND2_X1 U5256 ( .A1(n5940), .A2(n5933), .ZN(n6067) );
  NAND2_X1 U5257 ( .A1(n6072), .A2(n7624), .ZN(n6034) );
  AND2_X1 U5258 ( .A1(n5903), .A2(n5902), .ZN(n9197) );
  AOI21_X1 U5259 ( .B1(n9494), .B2(n5919), .A(n5893), .ZN(n9252) );
  AND4_X1 U5260 ( .A1(n5790), .A2(n5789), .A3(n5788), .A4(n5787), .ZN(n8105)
         );
  NAND2_X1 U5261 ( .A1(n9996), .A2(n9393), .ZN(n9997) );
  NOR2_X1 U5262 ( .A1(n9458), .A2(n4599), .ZN(n9428) );
  OR2_X1 U5263 ( .A1(n9493), .A2(n9298), .ZN(n4890) );
  NAND2_X1 U5264 ( .A1(n9510), .A2(n8311), .ZN(n9488) );
  NOR2_X1 U5265 ( .A1(n9757), .A2(n9276), .ZN(n8289) );
  NAND2_X1 U5266 ( .A1(n9757), .A2(n9276), .ZN(n4891) );
  OR2_X1 U5267 ( .A1(n9508), .A2(n9507), .ZN(n9510) );
  OR2_X1 U5268 ( .A1(n9539), .A2(n8287), .ZN(n4955) );
  AOI21_X1 U5269 ( .B1(n4853), .B2(n4855), .A(n4413), .ZN(n4851) );
  NAND2_X1 U5270 ( .A1(n8308), .A2(n4640), .ZN(n9543) );
  NOR2_X1 U5271 ( .A1(n8285), .A2(n4865), .ZN(n4860) );
  NAND2_X1 U5272 ( .A1(n4864), .A2(n4404), .ZN(n4861) );
  AND2_X1 U5273 ( .A1(n6057), .A2(n6056), .ZN(n9568) );
  NAND2_X1 U5274 ( .A1(n5862), .A2(n9550), .ZN(n9565) );
  NOR2_X1 U5275 ( .A1(n6052), .A2(n6015), .ZN(n4629) );
  AOI22_X1 U5276 ( .A1(n9624), .A2(n8278), .B1(n9307), .B2(n9628), .ZN(n9608)
         );
  INV_X1 U5277 ( .A(n4635), .ZN(n4634) );
  AND2_X1 U5278 ( .A1(n4632), .A2(n6048), .ZN(n4631) );
  AND2_X1 U5279 ( .A1(n4902), .A2(n8127), .ZN(n4899) );
  NAND2_X1 U5280 ( .A1(n4383), .A2(n4902), .ZN(n4898) );
  NAND2_X1 U5281 ( .A1(n8095), .A2(n6044), .ZN(n4636) );
  NAND2_X1 U5282 ( .A1(n4636), .A2(n4635), .ZN(n8203) );
  NAND2_X1 U5283 ( .A1(n8093), .A2(n4954), .ZN(n8128) );
  OR2_X1 U5284 ( .A1(n9872), .A2(n9311), .ZN(n8089) );
  NAND2_X1 U5285 ( .A1(n6009), .A2(n6045), .ZN(n8127) );
  AOI21_X1 U5286 ( .B1(n7869), .B2(n4870), .A(n4371), .ZN(n4869) );
  NAND2_X1 U5287 ( .A1(n9862), .A2(n8230), .ZN(n8226) );
  NOR2_X2 U5288 ( .A1(n7871), .A2(n9862), .ZN(n8235) );
  INV_X1 U5289 ( .A(n4849), .ZN(n4848) );
  OAI21_X1 U5290 ( .B1(n7612), .B2(n4850), .A(n7636), .ZN(n4849) );
  INV_X1 U5291 ( .A(n4957), .ZN(n4850) );
  OR2_X1 U5292 ( .A1(n9318), .A2(n7602), .ZN(n7603) );
  NAND2_X1 U5293 ( .A1(n7606), .A2(n7612), .ZN(n7625) );
  INV_X1 U5294 ( .A(n9320), .ZN(n7458) );
  NAND2_X1 U5295 ( .A1(n5151), .A2(n5150), .ZN(n9650) );
  AOI21_X1 U5296 ( .B1(n9451), .B2(n4606), .A(n4604), .ZN(n4603) );
  NAND2_X1 U5297 ( .A1(n4348), .A2(n9636), .ZN(n4602) );
  NAND2_X1 U5298 ( .A1(n5339), .A2(n5338), .ZN(n9461) );
  NAND2_X1 U5299 ( .A1(n5167), .A2(n5166), .ZN(n9685) );
  NAND2_X1 U5300 ( .A1(n5331), .A2(n5330), .ZN(n9558) );
  AND2_X1 U5301 ( .A1(n7577), .A2(n10069), .ZN(n10062) );
  OR2_X1 U5302 ( .A1(n6075), .A2(n6758), .ZN(n10069) );
  XNOR2_X1 U5303 ( .A(n5146), .B(n5145), .ZN(n8442) );
  INV_X1 U5304 ( .A(n4583), .ZN(n4582) );
  AND2_X1 U5305 ( .A1(n5127), .A2(n5130), .ZN(n4903) );
  NOR2_X1 U5306 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5127) );
  XNOR2_X1 U5307 ( .A(n5337), .B(n5336), .ZN(n8145) );
  NAND2_X1 U5308 ( .A1(n5096), .A2(n5095), .ZN(n5337) );
  XNOR2_X1 U5309 ( .A(n5161), .B(n5160), .ZN(n7956) );
  AND2_X1 U5310 ( .A1(n4500), .A2(n4501), .ZN(n5161) );
  OAI21_X1 U5311 ( .B1(n5291), .B2(n4485), .A(n4482), .ZN(n5316) );
  OAI21_X1 U5312 ( .B1(n5291), .B2(n4353), .A(n5041), .ZN(n5302) );
  AND2_X1 U5313 ( .A1(n4387), .A2(n5297), .ZN(n4796) );
  INV_X1 U5314 ( .A(n5294), .ZN(n4797) );
  NAND2_X1 U5315 ( .A1(n4496), .A2(n5033), .ZN(n5275) );
  NAND2_X1 U5316 ( .A1(n5268), .A2(n5031), .ZN(n4496) );
  NAND2_X1 U5317 ( .A1(n4998), .A2(n4997), .ZN(n5217) );
  XNOR2_X1 U5318 ( .A(n4993), .B(n7058), .ZN(n5201) );
  NAND2_X1 U5319 ( .A1(n4987), .A2(n4986), .ZN(n5192) );
  AND2_X1 U5320 ( .A1(n7672), .A2(n7671), .ZN(n7674) );
  NOR2_X1 U5321 ( .A1(n4347), .A2(n8688), .ZN(n4916) );
  INV_X1 U5322 ( .A(n8560), .ZN(n4919) );
  NAND2_X1 U5323 ( .A1(n4920), .A2(n4923), .ZN(n4918) );
  NAND2_X1 U5324 ( .A1(n4352), .A2(n4924), .ZN(n4923) );
  INV_X1 U5325 ( .A(n8570), .ZN(n4924) );
  AND4_X1 U5326 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n7774)
         );
  AND4_X1 U5327 ( .A1(n6212), .A2(n6211), .A3(n6210), .A4(n6209), .ZN(n7963)
         );
  XNOR2_X1 U5328 ( .A(n8549), .B(n8844), .ZN(n8607) );
  INV_X1 U5329 ( .A(n4929), .ZN(n4928) );
  OAI22_X1 U5330 ( .A1(n4930), .A2(n4934), .B1(n8518), .B2(n8519), .ZN(n4929)
         );
  NAND2_X1 U5331 ( .A1(n4932), .A2(n4931), .ZN(n4930) );
  OAI21_X1 U5332 ( .B1(n4516), .B2(n8461), .A(n4373), .ZN(n4515) );
  NAND2_X1 U5333 ( .A1(n6381), .A2(n6380), .ZN(n8877) );
  NAND2_X1 U5334 ( .A1(n6356), .A2(n6355), .ZN(n8905) );
  NAND4_X1 U5335 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n8706)
         );
  OR2_X1 U5336 ( .A1(n6149), .A2(n4536), .ZN(n6126) );
  AOI21_X1 U5337 ( .B1(n5584), .B2(n4329), .A(n6795), .ZN(n7253) );
  OAI21_X1 U5338 ( .B1(n8787), .B2(n4726), .A(n4724), .ZN(n4438) );
  NAND2_X1 U5339 ( .A1(n4727), .A2(n5568), .ZN(n4726) );
  NAND2_X1 U5340 ( .A1(n8787), .A2(n4725), .ZN(n4724) );
  AND2_X1 U5341 ( .A1(n4727), .A2(n4428), .ZN(n4725) );
  OAI21_X1 U5342 ( .B1(n5620), .B2(n7406), .A(n5619), .ZN(n5621) );
  NAND2_X1 U5343 ( .A1(n6349), .A2(n6348), .ZN(n9019) );
  NAND2_X1 U5344 ( .A1(n7010), .A2(n7009), .ZN(n10149) );
  NAND2_X1 U5345 ( .A1(n4714), .A2(n4712), .ZN(n8833) );
  AND2_X1 U5346 ( .A1(n8812), .A2(n10207), .ZN(n6472) );
  NAND2_X1 U5347 ( .A1(n6417), .A2(n6416), .ZN(n9064) );
  NAND2_X1 U5348 ( .A1(n8212), .A2(n8451), .ZN(n6417) );
  AND2_X1 U5349 ( .A1(n4714), .A2(n8430), .ZN(n8843) );
  INV_X1 U5350 ( .A(n9194), .ZN(n9195) );
  INV_X1 U5351 ( .A(n7610), .ZN(n10056) );
  NAND2_X1 U5352 ( .A1(n6752), .A2(n6751), .ZN(n8266) );
  AND2_X1 U5353 ( .A1(n6757), .A2(n6764), .ZN(n9885) );
  NAND2_X1 U5354 ( .A1(n4958), .A2(n6079), .ZN(n6081) );
  AND2_X1 U5355 ( .A1(n5926), .A2(n5925), .ZN(n9196) );
  INV_X1 U5356 ( .A(n9197), .ZN(n9296) );
  NAND4_X1 U5357 ( .A1(n5731), .A2(n5730), .A3(n5729), .A4(n5728), .ZN(n9316)
         );
  OR2_X1 U5358 ( .A1(n5898), .A2(n7665), .ZN(n5729) );
  OR2_X1 U5359 ( .A1(n4340), .A2(n5727), .ZN(n5728) );
  OR2_X1 U5360 ( .A1(n9968), .A2(n9967), .ZN(n9970) );
  NAND2_X1 U5361 ( .A1(n4454), .A2(n7570), .ZN(n4453) );
  INV_X1 U5362 ( .A(n4456), .ZN(n4455) );
  NOR2_X1 U5363 ( .A1(n5353), .A2(n9627), .ZN(n9424) );
  INV_X1 U5364 ( .A(n9654), .ZN(n4617) );
  OR2_X1 U5365 ( .A1(n10045), .A2(n7578), .ZN(n10020) );
  INV_X1 U5366 ( .A(n9478), .ZN(n9745) );
  AND3_X2 U5367 ( .A1(n5177), .A2(n5175), .A3(n5176), .ZN(n7436) );
  CLKBUF_X1 U5368 ( .A(n6521), .Z(n9418) );
  NOR2_X1 U5369 ( .A1(n4443), .A2(n4442), .ZN(n4441) );
  INV_X1 U5370 ( .A(n6006), .ZN(n4442) );
  INV_X1 U5371 ( .A(n8385), .ZN(n4547) );
  NAND2_X1 U5372 ( .A1(n8404), .A2(n8457), .ZN(n4448) );
  AND2_X1 U5373 ( .A1(n8129), .A2(n6045), .ZN(n4458) );
  INV_X1 U5374 ( .A(n8415), .ZN(n4534) );
  INV_X1 U5375 ( .A(n8411), .ZN(n4533) );
  NAND2_X1 U5376 ( .A1(n4751), .A2(n4749), .ZN(n8414) );
  NAND2_X1 U5377 ( .A1(n4752), .A2(n8457), .ZN(n4751) );
  NAND2_X1 U5378 ( .A1(n4377), .A2(n4750), .ZN(n4749) );
  NAND2_X1 U5379 ( .A1(n4356), .A2(n6075), .ZN(n4440) );
  AND2_X1 U5380 ( .A1(n8885), .A2(n8422), .ZN(n4767) );
  NAND2_X1 U5381 ( .A1(n8859), .A2(n4559), .ZN(n4558) );
  NAND2_X1 U5382 ( .A1(n8475), .A2(n8458), .ZN(n4559) );
  INV_X1 U5383 ( .A(n4564), .ZN(n4563) );
  OAI21_X1 U5384 ( .B1(n8426), .B2(n8474), .A(n8457), .ZN(n4564) );
  NOR2_X1 U5385 ( .A1(n4562), .A2(n8457), .ZN(n4561) );
  INV_X1 U5386 ( .A(n8428), .ZN(n4562) );
  NAND2_X1 U5387 ( .A1(n8440), .A2(n4449), .ZN(n4513) );
  NOR2_X1 U5388 ( .A1(n8500), .A2(n4450), .ZN(n4449) );
  AND2_X1 U5389 ( .A1(n4513), .A2(n4512), .ZN(n8447) );
  NAND2_X1 U5390 ( .A1(n8441), .A2(n8448), .ZN(n4512) );
  AND2_X1 U5391 ( .A1(n8502), .A2(n8446), .ZN(n8464) );
  AND2_X1 U5392 ( .A1(n8449), .A2(n8448), .ZN(n4760) );
  INV_X1 U5393 ( .A(n4513), .ZN(n8449) );
  NOR2_X1 U5394 ( .A1(n8447), .A2(n9064), .ZN(n4758) );
  NAND2_X1 U5395 ( .A1(n7225), .A2(n10131), .ZN(n8339) );
  NOR2_X1 U5396 ( .A1(n4950), .A2(n4818), .ZN(n4815) );
  AOI21_X1 U5397 ( .B1(n4820), .B2(n4817), .A(n9173), .ZN(n4816) );
  INV_X1 U5398 ( .A(n4881), .ZN(n4877) );
  NAND2_X1 U5399 ( .A1(n4881), .A2(n8289), .ZN(n4880) );
  OR2_X1 U5400 ( .A1(n9628), .A2(n9240), .ZN(n5944) );
  AND2_X1 U5401 ( .A1(n6036), .A2(n7605), .ZN(n5719) );
  NAND2_X1 U5402 ( .A1(n4588), .A2(n9767), .ZN(n4587) );
  NOR2_X1 U5403 ( .A1(n9708), .A2(n9610), .ZN(n4588) );
  NAND2_X1 U5404 ( .A1(n5107), .A2(n5106), .ZN(n5111) );
  INV_X1 U5405 ( .A(n5315), .ZN(n4481) );
  INV_X1 U5406 ( .A(n4498), .ZN(n4497) );
  OAI21_X1 U5407 ( .B1(n5031), .B2(n4499), .A(n5034), .ZN(n4498) );
  INV_X1 U5408 ( .A(n5274), .ZN(n5034) );
  INV_X1 U5409 ( .A(n5033), .ZN(n4499) );
  OAI21_X1 U5410 ( .B1(n6846), .B2(P1_DATAO_REG_11__SCAN_IN), .A(n4446), .ZN(
        n5020) );
  NAND2_X1 U5411 ( .A1(n6846), .A2(n5018), .ZN(n4446) );
  NAND2_X1 U5412 ( .A1(n5007), .A2(n5006), .ZN(n5010) );
  INV_X1 U5413 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4439) );
  OR2_X1 U5414 ( .A1(n6504), .A2(n8825), .ZN(n8466) );
  AND2_X1 U5415 ( .A1(n8015), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4452) );
  NAND2_X1 U5416 ( .A1(n10116), .A2(n4421), .ZN(n4827) );
  NAND2_X1 U5417 ( .A1(n4829), .A2(n4421), .ZN(n4828) );
  NOR2_X1 U5418 ( .A1(n5603), .A2(n5604), .ZN(n8795) );
  NAND2_X1 U5419 ( .A1(n8466), .A2(n8446), .ZN(n8500) );
  INV_X1 U5420 ( .A(n6238), .ZN(n4706) );
  AND2_X1 U5421 ( .A1(n8481), .A2(n6192), .ZN(n4723) );
  NAND2_X1 U5422 ( .A1(n10145), .A2(n6129), .ZN(n8338) );
  OR2_X1 U5423 ( .A1(n6149), .A2(n4540), .ZN(n6399) );
  INV_X1 U5424 ( .A(n4718), .ZN(n4717) );
  AND2_X1 U5425 ( .A1(n6330), .A2(n4716), .ZN(n4715) );
  NAND2_X1 U5426 ( .A1(n4773), .A2(n4772), .ZN(n8402) );
  AND2_X1 U5427 ( .A1(n8699), .A2(n6287), .ZN(n4772) );
  AND2_X1 U5428 ( .A1(n8392), .A2(n8391), .ZN(n8390) );
  NAND2_X1 U5429 ( .A1(n4674), .A2(n4672), .ZN(n8043) );
  AOI21_X1 U5430 ( .B1(n4675), .B2(n4678), .A(n4673), .ZN(n4672) );
  INV_X1 U5431 ( .A(n8381), .ZN(n4673) );
  NOR2_X1 U5432 ( .A1(n5409), .A2(n4942), .ZN(n4941) );
  NAND2_X1 U5433 ( .A1(n4943), .A2(n5410), .ZN(n4942) );
  CLKBUF_X1 U5434 ( .A(n5480), .Z(n5481) );
  INV_X1 U5435 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4910) );
  AND2_X1 U5436 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5689) );
  NAND2_X1 U5437 ( .A1(n4820), .A2(n4815), .ZN(n4814) );
  NAND2_X1 U5438 ( .A1(n4809), .A2(n4808), .ZN(n4807) );
  INV_X1 U5439 ( .A(n4815), .ZN(n4808) );
  INV_X1 U5440 ( .A(n4810), .ZN(n4809) );
  AOI21_X1 U5441 ( .B1(n4816), .B2(n4950), .A(n4811), .ZN(n4810) );
  INV_X1 U5442 ( .A(n9172), .ZN(n4811) );
  INV_X1 U5443 ( .A(n4816), .ZN(n4812) );
  OR2_X1 U5444 ( .A1(n6614), .A2(n7662), .ZN(n7812) );
  OR2_X1 U5445 ( .A1(n6557), .A2(n10050), .ZN(n6546) );
  NAND2_X1 U5446 ( .A1(n4475), .A2(n4474), .ZN(n4473) );
  OAI21_X1 U5447 ( .B1(n4467), .B2(n6067), .A(n5938), .ZN(n4476) );
  AND2_X1 U5448 ( .A1(n5940), .A2(n9294), .ZN(n4474) );
  NAND2_X1 U5449 ( .A1(n4887), .A2(n4886), .ZN(n4885) );
  INV_X1 U5450 ( .A(n8294), .ZN(n4887) );
  AND2_X1 U5451 ( .A1(n4890), .A2(n8292), .ZN(n4886) );
  AND2_X1 U5452 ( .A1(n4888), .A2(n4876), .ZN(n4875) );
  NOR2_X1 U5453 ( .A1(n4889), .A2(n8294), .ZN(n4888) );
  NAND2_X1 U5454 ( .A1(n4878), .A2(n4877), .ZN(n4876) );
  INV_X1 U5455 ( .A(n4890), .ZN(n4889) );
  NAND2_X1 U5456 ( .A1(n4875), .A2(n4879), .ZN(n4872) );
  OR2_X1 U5457 ( .A1(n9461), .A2(n9197), .ZN(n5979) );
  AOI21_X1 U5458 ( .B1(n9487), .B2(n5885), .A(n4624), .ZN(n4623) );
  INV_X1 U5459 ( .A(n8312), .ZN(n4624) );
  NAND2_X1 U5460 ( .A1(n4633), .A2(n4635), .ZN(n4632) );
  INV_X1 U5461 ( .A(n6044), .ZN(n4633) );
  NOR2_X1 U5462 ( .A1(n7876), .A2(n4868), .ZN(n4867) );
  INV_X1 U5463 ( .A(n7798), .ZN(n4868) );
  INV_X1 U5464 ( .A(n7867), .ZN(n4870) );
  NOR2_X1 U5465 ( .A1(n4592), .A2(n7784), .ZN(n4591) );
  AND2_X1 U5466 ( .A1(n5689), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5700) );
  OR2_X1 U5467 ( .A1(n7505), .A2(n7504), .ZN(n7632) );
  NAND2_X1 U5468 ( .A1(n4605), .A2(n8318), .ZN(n4604) );
  NAND2_X1 U5469 ( .A1(n4384), .A2(n4608), .ZN(n4605) );
  NAND2_X1 U5470 ( .A1(n8297), .A2(n4609), .ZN(n4608) );
  AND2_X1 U5471 ( .A1(n4396), .A2(n9636), .ZN(n4606) );
  NOR2_X1 U5472 ( .A1(n9501), .A2(n9493), .ZN(n9492) );
  NOR2_X1 U5473 ( .A1(n9625), .A2(n4586), .ZN(n9598) );
  INV_X1 U5474 ( .A(n4588), .ZN(n4586) );
  XNOR2_X1 U5475 ( .A(n5111), .B(n5110), .ZN(n5149) );
  AOI21_X1 U5476 ( .B1(n5336), .B2(n4509), .A(n4508), .ZN(n4507) );
  INV_X1 U5477 ( .A(n5102), .ZN(n4508) );
  INV_X1 U5478 ( .A(n5095), .ZN(n4509) );
  INV_X1 U5479 ( .A(n5336), .ZN(n4510) );
  NAND2_X1 U5480 ( .A1(n4416), .A2(n5070), .ZN(n4501) );
  INV_X1 U5481 ( .A(n5064), .ZN(n4502) );
  AND2_X1 U5482 ( .A1(n7177), .A2(n5318), .ZN(n4794) );
  NAND2_X1 U5483 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n4795) );
  OAI21_X1 U5484 ( .B1(n5318), .B2(P1_IR_REG_31__SCAN_IN), .A(n4793), .ZN(
        n4792) );
  OAI21_X1 U5485 ( .B1(n5318), .B2(n7177), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4793) );
  AOI21_X1 U5486 ( .B1(n4484), .B2(n4483), .A(n4415), .ZN(n4482) );
  INV_X1 U5487 ( .A(n4489), .ZN(n4483) );
  INV_X1 U5488 ( .A(n5267), .ZN(n5031) );
  NOR2_X1 U5489 ( .A1(n4361), .A2(n4766), .ZN(n4765) );
  INV_X1 U5490 ( .A(n5016), .ZN(n4766) );
  AND2_X1 U5491 ( .A1(n5025), .A2(n5254), .ZN(n5026) );
  NAND2_X1 U5492 ( .A1(n4614), .A2(n5002), .ZN(n5225) );
  OAI21_X1 U5493 ( .B1(n6846), .B2(P1_DATAO_REG_5__SCAN_IN), .A(n4994), .ZN(
        n4995) );
  OR2_X1 U5494 ( .A1(n6100), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n4994) );
  CLKBUF_X1 U5495 ( .A(n8622), .Z(n8623) );
  AOI21_X1 U5496 ( .B1(n4913), .B2(n4948), .A(n8595), .ZN(n4912) );
  XNOR2_X1 U5497 ( .A(n9019), .B(n8558), .ZN(n8650) );
  OR2_X1 U5498 ( .A1(n8530), .A2(n8529), .ZN(n8662) );
  OR2_X1 U5499 ( .A1(n4935), .A2(n4933), .ZN(n4932) );
  INV_X1 U5500 ( .A(n4938), .ZN(n4933) );
  NOR2_X1 U5501 ( .A1(n4936), .A2(n8176), .ZN(n4935) );
  INV_X1 U5502 ( .A(n8149), .ZN(n4936) );
  INV_X1 U5503 ( .A(n8520), .ZN(n4931) );
  AND2_X1 U5504 ( .A1(n8082), .A2(n4938), .ZN(n4934) );
  OR2_X1 U5505 ( .A1(n9055), .A2(n8468), .ZN(n4964) );
  NAND2_X1 U5506 ( .A1(n4517), .A2(n4359), .ZN(n4516) );
  NAND2_X1 U5507 ( .A1(n8459), .A2(n8457), .ZN(n4517) );
  NOR2_X1 U5508 ( .A1(n8459), .A2(n4755), .ZN(n8461) );
  AND2_X1 U5509 ( .A1(n8460), .A2(n8501), .ZN(n4755) );
  INV_X1 U5510 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n4544) );
  OR2_X1 U5511 ( .A1(n6149), .A2(n4542), .ZN(n6429) );
  INV_X1 U5512 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n4542) );
  OR2_X1 U5513 ( .A1(n6149), .A2(n4541), .ZN(n6411) );
  OR2_X1 U5514 ( .A1(n6149), .A2(n4538), .ZN(n6378) );
  INV_X1 U5515 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n4538) );
  INV_X2 U5516 ( .A(n6442), .ZN(n8453) );
  XNOR2_X1 U5517 ( .A(n5582), .B(n7425), .ZN(n7417) );
  NOR2_X1 U5518 ( .A1(n5474), .A2(n4741), .ZN(n7244) );
  NAND2_X1 U5519 ( .A1(n7245), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7397) );
  NAND2_X1 U5520 ( .A1(n7244), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7392) );
  NAND2_X1 U5521 ( .A1(n4731), .A2(n5478), .ZN(n7361) );
  AOI21_X1 U5522 ( .B1(n5588), .B2(n5478), .A(n7384), .ZN(n7357) );
  XNOR2_X1 U5523 ( .A(n4952), .B(n7550), .ZN(n7545) );
  NOR2_X1 U5524 ( .A1(n7545), .A2(n7546), .ZN(n7544) );
  NOR2_X1 U5525 ( .A1(n7740), .A2(n4451), .ZN(n5487) );
  NOR2_X1 U5526 ( .A1(n6194), .A2(n7687), .ZN(n4451) );
  NAND2_X1 U5527 ( .A1(n7829), .A2(n5593), .ZN(n7895) );
  OR2_X1 U5528 ( .A1(n5511), .A2(n9152), .ZN(n5453) );
  NOR2_X1 U5529 ( .A1(n5491), .A2(n8709), .ZN(n8021) );
  XNOR2_X1 U5530 ( .A(n5494), .B(n10091), .ZN(n10093) );
  OAI21_X1 U5531 ( .B1(n10093), .B2(n4747), .A(n4746), .ZN(n10110) );
  NAND2_X1 U5532 ( .A1(n4748), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4747) );
  NAND2_X1 U5533 ( .A1(n5495), .A2(n4748), .ZN(n4746) );
  INV_X1 U5534 ( .A(n10111), .ZN(n4748) );
  NOR2_X1 U5535 ( .A1(n10093), .A2(n10094), .ZN(n10092) );
  NAND2_X1 U5536 ( .A1(n10112), .A2(n5598), .ZN(n8734) );
  OR2_X1 U5537 ( .A1(n8747), .A2(n8746), .ZN(n8748) );
  OR2_X1 U5538 ( .A1(n8727), .A2(n4735), .ZN(n4732) );
  OR2_X1 U5539 ( .A1(n8745), .A2(n8728), .ZN(n4735) );
  NAND2_X1 U5540 ( .A1(n5501), .A2(n4734), .ZN(n4733) );
  INV_X1 U5541 ( .A(n8745), .ZN(n4734) );
  NAND2_X1 U5542 ( .A1(n8751), .A2(n5600), .ZN(n8773) );
  NAND2_X1 U5543 ( .A1(n4844), .A2(n4842), .ZN(n8769) );
  NOR2_X1 U5544 ( .A1(n4843), .A2(n5560), .ZN(n8771) );
  NAND2_X1 U5545 ( .A1(n4845), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n4841) );
  AND2_X1 U5546 ( .A1(n8764), .A2(n4426), .ZN(n4727) );
  INV_X1 U5547 ( .A(n5525), .ZN(n4728) );
  INV_X1 U5548 ( .A(n5568), .ZN(n4729) );
  INV_X1 U5549 ( .A(n8500), .ZN(n8441) );
  NAND2_X1 U5550 ( .A1(n6408), .A2(n6407), .ZN(n6418) );
  INV_X1 U5551 ( .A(n6409), .ZN(n6408) );
  OR2_X1 U5552 ( .A1(n6397), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6409) );
  NAND2_X1 U5553 ( .A1(n4658), .A2(n4657), .ZN(n8868) );
  NOR2_X1 U5554 ( .A1(n8425), .A2(n8323), .ZN(n4657) );
  NAND2_X1 U5555 ( .A1(n6374), .A2(n6373), .ZN(n6387) );
  INV_X1 U5556 ( .A(n6375), .ZN(n6374) );
  AND2_X1 U5557 ( .A1(n6460), .A2(n8322), .ZN(n8885) );
  AOI21_X1 U5558 ( .B1(n8912), .B2(n8417), .A(n4956), .ZN(n8882) );
  NAND2_X1 U5559 ( .A1(n6341), .A2(n6340), .ZN(n6350) );
  INV_X1 U5560 ( .A(n6342), .ZN(n6341) );
  NAND2_X1 U5561 ( .A1(n6324), .A2(n6323), .ZN(n6333) );
  INV_X1 U5562 ( .A(n6325), .ZN(n6324) );
  NAND2_X1 U5563 ( .A1(n6300), .A2(n6299), .ZN(n6311) );
  INV_X1 U5564 ( .A(n6301), .ZN(n6300) );
  NAND2_X1 U5565 ( .A1(n6278), .A2(n6277), .ZN(n6288) );
  INV_X1 U5566 ( .A(n6279), .ZN(n6278) );
  OR2_X1 U5567 ( .A1(n6267), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6279) );
  NAND2_X1 U5568 ( .A1(n6256), .A2(n6255), .ZN(n6267) );
  INV_X1 U5569 ( .A(n6257), .ZN(n6256) );
  NAND2_X1 U5570 ( .A1(n6243), .A2(n8014), .ZN(n6257) );
  INV_X1 U5571 ( .A(n6244), .ZN(n6243) );
  OR2_X1 U5572 ( .A1(n6232), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6244) );
  OR2_X1 U5573 ( .A1(n6220), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U5574 ( .A1(n6206), .A2(n6205), .ZN(n6220) );
  INV_X1 U5575 ( .A(n6207), .ZN(n6206) );
  OAI21_X1 U5576 ( .B1(n4684), .B2(n4683), .A(n8353), .ZN(n4682) );
  INV_X1 U5577 ( .A(n8371), .ZN(n4683) );
  AND2_X1 U5578 ( .A1(n8373), .A2(n8357), .ZN(n8487) );
  NAND2_X1 U5579 ( .A1(n4966), .A2(n6204), .ZN(n7761) );
  OR2_X1 U5580 ( .A1(n6198), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U5581 ( .A1(n6193), .A2(n4723), .ZN(n4966) );
  NAND2_X1 U5582 ( .A1(n6193), .A2(n6192), .ZN(n7682) );
  NAND2_X1 U5583 ( .A1(n6183), .A2(n6182), .ZN(n6198) );
  INV_X1 U5584 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6182) );
  INV_X1 U5585 ( .A(n6184), .ZN(n6183) );
  NAND2_X1 U5586 ( .A1(n4701), .A2(n7477), .ZN(n7704) );
  AOI21_X1 U5587 ( .B1(n4696), .B2(n4698), .A(n4695), .ZN(n4694) );
  INV_X1 U5588 ( .A(n4698), .ZN(n4697) );
  OR2_X1 U5589 ( .A1(n6169), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6184) );
  NAND2_X1 U5590 ( .A1(n10141), .A2(n6147), .ZN(n6159) );
  INV_X1 U5591 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U5592 ( .A1(n6158), .A2(n6157), .ZN(n6169) );
  INV_X1 U5593 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n6157) );
  INV_X1 U5594 ( .A(n6159), .ZN(n6158) );
  NOR2_X1 U5595 ( .A1(n4643), .A2(n4642), .ZN(n4641) );
  INV_X1 U5596 ( .A(n8361), .ZN(n4642) );
  NAND2_X1 U5597 ( .A1(n4693), .A2(n4698), .ZN(n7481) );
  NAND2_X1 U5598 ( .A1(n7492), .A2(n4699), .ZN(n4693) );
  NAND2_X1 U5599 ( .A1(n10136), .A2(n10137), .ZN(n4644) );
  INV_X1 U5600 ( .A(n8335), .ZN(n10150) );
  INV_X1 U5601 ( .A(n8830), .ZN(n8834) );
  AND2_X1 U5602 ( .A1(n10147), .A2(n10221), .ZN(n7009) );
  NAND2_X1 U5603 ( .A1(n4661), .A2(n4659), .ZN(n8821) );
  AOI21_X1 U5604 ( .B1(n4663), .B2(n4665), .A(n4660), .ZN(n4659) );
  INV_X1 U5605 ( .A(n8437), .ZN(n4660) );
  AND2_X1 U5606 ( .A1(n8896), .A2(n8897), .ZN(n8914) );
  NOR2_X1 U5607 ( .A1(n8944), .A2(n4680), .ZN(n4679) );
  INV_X1 U5608 ( .A(n8410), .ZN(n4680) );
  AND2_X1 U5609 ( .A1(n8402), .A2(n8406), .ZN(n8968) );
  NAND2_X1 U5610 ( .A1(n4647), .A2(n4645), .ZN(n8966) );
  AOI21_X1 U5611 ( .B1(n4648), .B2(n4653), .A(n4646), .ZN(n4645) );
  INV_X1 U5612 ( .A(n8401), .ZN(n4646) );
  INV_X1 U5613 ( .A(n8390), .ZN(n8489) );
  AND2_X1 U5614 ( .A1(n5440), .A2(n4703), .ZN(n4702) );
  NOR2_X1 U5615 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  OR2_X1 U5616 ( .A1(n5416), .A2(n5415), .ZN(n5422) );
  XNOR2_X1 U5617 ( .A(n5465), .B(P2_IR_REG_4__SCAN_IN), .ZN(n7400) );
  XNOR2_X1 U5618 ( .A(n5468), .B(n5467), .ZN(n5533) );
  INV_X1 U5619 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U5620 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5468) );
  OR2_X1 U5621 ( .A1(n5785), .A2(n5624), .ZN(n5792) );
  AND2_X1 U5622 ( .A1(n9249), .A2(n6725), .ZN(n9162) );
  AND2_X1 U5623 ( .A1(n5747), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5757) );
  NAND2_X1 U5624 ( .A1(n5726), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5736) );
  NOR2_X1 U5625 ( .A1(n9237), .A2(n4820), .ZN(n9234) );
  AND2_X1 U5626 ( .A1(n9261), .A2(n9262), .ZN(n6705) );
  INV_X1 U5627 ( .A(n5854), .ZN(n5629) );
  AND2_X1 U5628 ( .A1(n6805), .A2(n6810), .ZN(n9286) );
  INV_X1 U5629 ( .A(n4775), .ZN(n4774) );
  NAND2_X1 U5630 ( .A1(n6579), .A2(n7533), .ZN(n4799) );
  NOR2_X1 U5631 ( .A1(n6579), .A2(n7533), .ZN(n4800) );
  NAND2_X1 U5632 ( .A1(n5625), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5807) );
  INV_X1 U5633 ( .A(n5792), .ZN(n5625) );
  OR2_X1 U5634 ( .A1(n5807), .A2(n5806), .ZN(n5809) );
  AOI211_X1 U5635 ( .C1(n6032), .C2(n6031), .A(n6063), .B(n6062), .ZN(n6033)
         );
  AND3_X1 U5636 ( .A1(n5655), .A2(n5654), .A3(n5653), .ZN(n9177) );
  INV_X1 U5637 ( .A(n4339), .ZN(n5909) );
  AND4_X1 U5638 ( .A1(n5762), .A2(n5761), .A3(n5760), .A4(n5759), .ZN(n8230)
         );
  NAND2_X1 U5639 ( .A1(n6835), .A2(n6836), .ZN(n6905) );
  NOR2_X1 U5640 ( .A1(n9365), .A2(n4435), .ZN(n9366) );
  AND2_X1 U5641 ( .A1(n9370), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n4435) );
  AOI21_X1 U5642 ( .B1(n9370), .B2(P1_REG1_REG_8__SCAN_IN), .A(n9369), .ZN(
        n9373) );
  AND2_X1 U5643 ( .A1(n9404), .A2(n9904), .ZN(n9928) );
  AND2_X1 U5644 ( .A1(n9943), .A2(n9944), .ZN(n9941) );
  AND2_X1 U5645 ( .A1(n9924), .A2(n9386), .ZN(n9939) );
  NOR2_X1 U5646 ( .A1(n9939), .A2(n9938), .ZN(n9937) );
  AOI21_X1 U5647 ( .B1(n9407), .B2(P1_REG1_REG_14__SCAN_IN), .A(n9941), .ZN(
        n9408) );
  AOI21_X1 U5648 ( .B1(n9407), .B2(P1_REG2_REG_14__SCAN_IN), .A(n9937), .ZN(
        n9388) );
  AND2_X1 U5649 ( .A1(n9979), .A2(n9392), .ZN(n9996) );
  NAND2_X1 U5650 ( .A1(n4621), .A2(n4623), .ZN(n9471) );
  NAND2_X1 U5651 ( .A1(n4622), .A2(n9487), .ZN(n4621) );
  INV_X1 U5652 ( .A(n9510), .ZN(n4622) );
  INV_X1 U5653 ( .A(n4638), .ZN(n4637) );
  OAI21_X1 U5654 ( .B1(n4640), .B2(n4358), .A(n8310), .ZN(n4638) );
  NAND2_X1 U5655 ( .A1(n9535), .A2(n9757), .ZN(n9524) );
  OR2_X1 U5656 ( .A1(n9571), .A2(n9558), .ZN(n9556) );
  NOR2_X1 U5657 ( .A1(n9685), .A2(n9556), .ZN(n9535) );
  NAND2_X1 U5658 ( .A1(n4854), .A2(n4862), .ZN(n4853) );
  INV_X1 U5659 ( .A(n4857), .ZN(n4854) );
  AOI21_X1 U5660 ( .B1(n4859), .B2(n4858), .A(n4406), .ZN(n4857) );
  NAND2_X1 U5661 ( .A1(n4859), .A2(n4862), .ZN(n4855) );
  INV_X1 U5662 ( .A(n4627), .ZN(n4626) );
  OAI21_X1 U5663 ( .B1(n4628), .B2(n9634), .A(n6053), .ZN(n4627) );
  NAND2_X1 U5664 ( .A1(n5627), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5846) );
  AND2_X1 U5665 ( .A1(n5942), .A2(n6056), .ZN(n9581) );
  NOR2_X1 U5666 ( .A1(n9625), .A2(n9610), .ZN(n9609) );
  NAND2_X1 U5667 ( .A1(n4630), .A2(n6051), .ZN(n9616) );
  OR2_X1 U5668 ( .A1(n8195), .A2(n9628), .ZN(n9625) );
  NAND2_X1 U5669 ( .A1(n4893), .A2(n4892), .ZN(n9624) );
  AOI21_X1 U5670 ( .B1(n4895), .B2(n4897), .A(n4381), .ZN(n4892) );
  NAND2_X1 U5671 ( .A1(n8128), .A2(n4895), .ZN(n4893) );
  AND2_X1 U5672 ( .A1(n8235), .A2(n4398), .ZN(n8194) );
  NOR2_X1 U5673 ( .A1(n4595), .A2(n9312), .ZN(n7984) );
  AND2_X1 U5674 ( .A1(n8094), .A2(n6006), .ZN(n7991) );
  NAND2_X1 U5675 ( .A1(n8235), .A2(n4594), .ZN(n4968) );
  NAND2_X1 U5676 ( .A1(n7878), .A2(n6038), .ZN(n8227) );
  AND2_X1 U5677 ( .A1(n7877), .A2(n7876), .ZN(n6038) );
  NAND2_X1 U5678 ( .A1(n8235), .A2(n10068), .ZN(n8234) );
  OR2_X1 U5679 ( .A1(n7915), .A2(n7952), .ZN(n7871) );
  NAND3_X1 U5680 ( .A1(n4590), .A2(n4589), .A3(n4591), .ZN(n7915) );
  NAND2_X1 U5681 ( .A1(n4847), .A2(n4846), .ZN(n7909) );
  AOI21_X1 U5682 ( .B1(n4848), .B2(n4850), .A(n4367), .ZN(n4846) );
  NOR2_X1 U5683 ( .A1(n7503), .A2(n4592), .ZN(n7627) );
  AND2_X1 U5684 ( .A1(n5700), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5726) );
  NOR2_X1 U5685 ( .A1(n7503), .A2(n7602), .ZN(n7608) );
  NAND2_X1 U5686 ( .A1(n10050), .A2(n7304), .ZN(n7305) );
  INV_X1 U5687 ( .A(n5953), .ZN(n7259) );
  AND2_X1 U5688 ( .A1(n7436), .A2(n7264), .ZN(n7649) );
  NAND2_X1 U5689 ( .A1(n5155), .A2(n5154), .ZN(n9478) );
  NAND2_X1 U5690 ( .A1(n5335), .A2(n5334), .ZN(n9502) );
  NAND2_X1 U5691 ( .A1(n5326), .A2(n5325), .ZN(n9697) );
  XNOR2_X1 U5692 ( .A(n5123), .B(n5122), .ZN(n9151) );
  OAI21_X1 U5693 ( .B1(n5146), .B2(n5145), .A(n5118), .ZN(n5123) );
  XNOR2_X1 U5694 ( .A(n5149), .B(SI_29_), .ZN(n8218) );
  NOR2_X1 U5695 ( .A1(n4907), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n4906) );
  NAND2_X1 U5696 ( .A1(n4908), .A2(n5141), .ZN(n4907) );
  NOR2_X1 U5697 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_26__SCAN_IN), .ZN(
        n4908) );
  NAND2_X1 U5698 ( .A1(n5141), .A2(n4463), .ZN(n4462) );
  INV_X1 U5699 ( .A(n5365), .ZN(n5371) );
  NAND2_X1 U5700 ( .A1(n4503), .A2(n5064), .ZN(n5165) );
  NAND2_X1 U5701 ( .A1(n4486), .A2(n4487), .ZN(n5307) );
  NAND2_X1 U5702 ( .A1(n5291), .A2(n4489), .ZN(n4486) );
  XNOR2_X1 U5703 ( .A(n5291), .B(n5290), .ZN(n7197) );
  AND2_X1 U5704 ( .A1(n5270), .A2(n5269), .ZN(n5277) );
  AND2_X1 U5705 ( .A1(n4905), .A2(n5126), .ZN(n5270) );
  OR3_X1 U5706 ( .A1(n5234), .A2(P1_IR_REG_7__SCAN_IN), .A3(
        P1_IR_REG_6__SCAN_IN), .ZN(n5240) );
  INV_X1 U5707 ( .A(n5201), .ZN(n4493) );
  AOI21_X1 U5708 ( .B1(n5201), .B2(n4492), .A(n4372), .ZN(n4491) );
  INV_X1 U5709 ( .A(n4991), .ZN(n4492) );
  XNOR2_X1 U5710 ( .A(n4995), .B(SI_5_), .ZN(n5209) );
  NAND2_X1 U5711 ( .A1(n4982), .A2(n4981), .ZN(n5184) );
  XNOR2_X1 U5712 ( .A(n4979), .B(SI_1_), .ZN(n5169) );
  INV_X4 U5713 ( .A(n6100), .ZN(n6846) );
  NAND2_X1 U5714 ( .A1(n4927), .A2(n4932), .ZN(n8521) );
  NAND2_X1 U5715 ( .A1(n8083), .A2(n4934), .ZN(n4927) );
  INV_X1 U5716 ( .A(n8877), .ZN(n8854) );
  INV_X1 U5717 ( .A(n8672), .ZN(n8681) );
  NAND2_X1 U5718 ( .A1(n4909), .A2(n7442), .ZN(n7338) );
  NAND2_X1 U5719 ( .A1(n7852), .A2(n7851), .ZN(n7853) );
  AND2_X1 U5720 ( .A1(n4914), .A2(n8535), .ZN(n8641) );
  AND2_X1 U5721 ( .A1(n4937), .A2(n4939), .ZN(n8150) );
  NAND2_X1 U5722 ( .A1(n8083), .A2(n8082), .ZN(n4937) );
  AND2_X1 U5723 ( .A1(n6368), .A2(n6367), .ZN(n8865) );
  OR2_X1 U5724 ( .A1(n7002), .A2(n7001), .ZN(n8673) );
  AND2_X1 U5725 ( .A1(n7521), .A2(n7519), .ZN(n4926) );
  AND2_X1 U5726 ( .A1(n7520), .A2(n7519), .ZN(n7522) );
  NAND2_X1 U5727 ( .A1(n6424), .A2(n6423), .ZN(n8697) );
  NAND2_X1 U5728 ( .A1(n6393), .A2(n6392), .ZN(n8844) );
  INV_X1 U5729 ( .A(n8865), .ZN(n8888) );
  INV_X1 U5730 ( .A(n8075), .ZN(n8068) );
  INV_X1 U5731 ( .A(n7963), .ZN(n8702) );
  OR2_X1 U5732 ( .A1(n6145), .A2(n6111), .ZN(n6112) );
  AOI21_X1 U5733 ( .B1(n5586), .B2(n6849), .A(n7405), .ZN(n7385) );
  NOR2_X1 U5734 ( .A1(n7742), .A2(n7741), .ZN(n7740) );
  NOR2_X1 U5735 ( .A1(n7824), .A2(n7825), .ZN(n7823) );
  INV_X1 U5736 ( .A(n4833), .ZN(n7826) );
  OAI21_X1 U5737 ( .B1(n7827), .B2(n4831), .A(n4830), .ZN(n7892) );
  NAND2_X1 U5738 ( .A1(n4834), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4831) );
  INV_X1 U5739 ( .A(n7893), .ZN(n4834) );
  INV_X1 U5740 ( .A(n5547), .ZN(n4832) );
  NAND2_X1 U5741 ( .A1(n4839), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4836) );
  INV_X1 U5742 ( .A(n8010), .ZN(n4839) );
  INV_X1 U5743 ( .A(n5549), .ZN(n4837) );
  NOR2_X1 U5744 ( .A1(n10099), .A2(n5552), .ZN(n10117) );
  NOR2_X1 U5745 ( .A1(n8729), .A2(n8249), .ZN(n8731) );
  NAND2_X1 U5746 ( .A1(n4733), .A2(n4732), .ZN(n8744) );
  INV_X1 U5747 ( .A(n5501), .ZN(n4736) );
  NOR2_X1 U5748 ( .A1(n8762), .A2(n8962), .ZN(n8765) );
  AOI22_X1 U5749 ( .A1(n9151), .A2(n8451), .B1(n8450), .B2(
        P1_DATAO_REG_31__SCAN_IN), .ZN(n8809) );
  XNOR2_X1 U5750 ( .A(n8467), .B(n8441), .ZN(n8812) );
  NAND2_X1 U5751 ( .A1(n8953), .A2(n8410), .ZN(n8945) );
  NAND2_X1 U5752 ( .A1(n4719), .A2(n6307), .ZN(n8939) );
  NAND2_X1 U5753 ( .A1(n6298), .A2(n6297), .ZN(n9039) );
  AOI21_X1 U5754 ( .B1(n6962), .B2(n8451), .A(n6266), .ZN(n8982) );
  NAND2_X1 U5755 ( .A1(n6241), .A2(n6240), .ZN(n10220) );
  NAND2_X1 U5756 ( .A1(n7973), .A2(n6238), .ZN(n8040) );
  AND2_X1 U5757 ( .A1(n4677), .A2(n8377), .ZN(n7972) );
  OR2_X1 U5758 ( .A1(n7961), .A2(n4678), .ZN(n4677) );
  NAND2_X1 U5759 ( .A1(n6218), .A2(n6217), .ZN(n8076) );
  NAND2_X1 U5760 ( .A1(n6214), .A2(n6213), .ZN(n7861) );
  AND2_X1 U5761 ( .A1(n6196), .A2(n6195), .ZN(n10193) );
  NAND2_X1 U5762 ( .A1(n4686), .A2(n8368), .ZN(n7727) );
  AOI21_X1 U5763 ( .B1(n7493), .B2(n10135), .A(n4526), .ZN(n10174) );
  NAND2_X1 U5764 ( .A1(n4528), .A2(n4527), .ZN(n4526) );
  NAND2_X1 U5765 ( .A1(n8707), .A2(n10132), .ZN(n4527) );
  INV_X1 U5766 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10141) );
  NAND2_X1 U5767 ( .A1(n4688), .A2(n6130), .ZN(n10129) );
  NAND2_X1 U5768 ( .A1(n6102), .A2(n4362), .ZN(n6104) );
  AND2_X1 U5769 ( .A1(n8444), .A2(n8443), .ZN(n8996) );
  INV_X1 U5770 ( .A(n8809), .ZN(n9055) );
  INV_X1 U5771 ( .A(n8996), .ZN(n9059) );
  XNOR2_X1 U5772 ( .A(n8821), .B(n8822), .ZN(n9067) );
  NAND2_X1 U5773 ( .A1(n6406), .A2(n6405), .ZN(n9070) );
  NAND2_X1 U5774 ( .A1(n4662), .A2(n4666), .ZN(n8831) );
  NAND2_X1 U5775 ( .A1(n8858), .A2(n4668), .ZN(n4662) );
  NAND2_X1 U5776 ( .A1(n6396), .A2(n6395), .ZN(n9076) );
  NAND2_X1 U5777 ( .A1(n4671), .A2(n8431), .ZN(n8841) );
  OR2_X1 U5778 ( .A1(n8858), .A2(n6463), .ZN(n4671) );
  NAND2_X1 U5779 ( .A1(n6384), .A2(n6383), .ZN(n9083) );
  NAND2_X1 U5780 ( .A1(n6372), .A2(n6371), .ZN(n9090) );
  NAND2_X1 U5781 ( .A1(n6361), .A2(n6360), .ZN(n9096) );
  NAND2_X1 U5782 ( .A1(n8887), .A2(n6359), .ZN(n8876) );
  NAND2_X1 U5783 ( .A1(n6339), .A2(n6338), .ZN(n9103) );
  NAND2_X1 U5784 ( .A1(n6332), .A2(n6331), .ZN(n9109) );
  NAND2_X1 U5785 ( .A1(n6320), .A2(n6319), .ZN(n9115) );
  NAND2_X1 U5786 ( .A1(n4773), .A2(n6287), .ZN(n9130) );
  NAND2_X1 U5787 ( .A1(n6276), .A2(n6275), .ZN(n8694) );
  NAND2_X1 U5788 ( .A1(n4650), .A2(n4651), .ZN(n8243) );
  OR2_X1 U5789 ( .A1(n8121), .A2(n4653), .ZN(n4650) );
  NAND2_X1 U5790 ( .A1(n8121), .A2(n8391), .ZN(n4656) );
  NAND2_X1 U5791 ( .A1(n6254), .A2(n6253), .ZN(n9143) );
  INV_X1 U5792 ( .A(n9122), .ZN(n9144) );
  INV_X2 U5793 ( .A(n10224), .ZN(n10222) );
  INV_X1 U5794 ( .A(n7348), .ZN(n8326) );
  NAND2_X1 U5795 ( .A1(n4520), .A2(n4522), .ZN(n6434) );
  INV_X1 U5796 ( .A(n6176), .ZN(n7364) );
  OR2_X1 U5797 ( .A1(n5466), .A2(n9152), .ZN(n4826) );
  INV_X1 U5798 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10089) );
  AND2_X1 U5799 ( .A1(n4970), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U5800 ( .A1(n5345), .A2(n5344), .ZN(n9655) );
  NAND2_X1 U5801 ( .A1(n8212), .A2(n5342), .ZN(n5345) );
  NAND2_X1 U5802 ( .A1(n6544), .A2(n6543), .ZN(n6979) );
  NAND2_X1 U5803 ( .A1(n6534), .A2(n7236), .ZN(n6980) );
  AND2_X1 U5804 ( .A1(n6648), .A2(n6647), .ZN(n9869) );
  NAND2_X1 U5805 ( .A1(n4424), .A2(n7530), .ZN(n7531) );
  NAND2_X1 U5806 ( .A1(n4798), .A2(n6579), .ZN(n7530) );
  OR2_X1 U5807 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  INV_X1 U5808 ( .A(n10068), .ZN(n4595) );
  AND2_X1 U5809 ( .A1(n6764), .A2(n6763), .ZN(n9882) );
  INV_X1 U5810 ( .A(n4802), .ZN(n4801) );
  NAND2_X1 U5811 ( .A1(n4804), .A2(n6673), .ZN(n8167) );
  NAND2_X1 U5812 ( .A1(n5288), .A2(n5287), .ZN(n8274) );
  INV_X1 U5813 ( .A(n9280), .ZN(n9887) );
  NAND4_X2 U5814 ( .A1(n5673), .A2(n5672), .A3(n5671), .A4(n5670), .ZN(n9324)
         );
  AND2_X1 U5815 ( .A1(n6905), .A2(n4433), .ZN(n6948) );
  NAND2_X1 U5816 ( .A1(n6911), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4433) );
  AOI21_X1 U5817 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n6911), .A(n6910), .ZN(
        n6945) );
  AOI21_X1 U5818 ( .B1(n6949), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6943), .ZN(
        n6914) );
  AOI21_X1 U5819 ( .B1(n6949), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6946), .ZN(
        n6908) );
  NOR2_X1 U5820 ( .A1(n6920), .A2(n4432), .ZN(n6933) );
  AND2_X1 U5821 ( .A1(n6924), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4432) );
  AOI21_X1 U5822 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n6937), .A(n6934), .ZN(
        n6926) );
  NOR2_X1 U5823 ( .A1(n6931), .A2(n4434), .ZN(n6922) );
  AND2_X1 U5824 ( .A1(n6937), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4434) );
  AOI21_X1 U5825 ( .B1(n9853), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9845), .ZN(
        n9896) );
  NOR2_X1 U5826 ( .A1(n9848), .A2(n4436), .ZN(n9893) );
  AND2_X1 U5827 ( .A1(n9853), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4436) );
  NOR2_X1 U5828 ( .A1(n9954), .A2(n9955), .ZN(n9953) );
  AND2_X1 U5829 ( .A1(n9970), .A2(n9391), .ZN(n9980) );
  AOI211_X1 U5830 ( .C1(n9432), .C2(n9431), .A(n9627), .B(n9430), .ZN(n9648)
         );
  AOI21_X1 U5831 ( .B1(n9446), .B2(n9636), .A(n9445), .ZN(n9658) );
  AND2_X1 U5832 ( .A1(n9436), .A2(n4967), .ZN(n9659) );
  NAND2_X1 U5833 ( .A1(n4884), .A2(n4890), .ZN(n9469) );
  OR2_X1 U5834 ( .A1(n9485), .A2(n8292), .ZN(n4884) );
  NAND2_X1 U5835 ( .A1(n9488), .A2(n9487), .ZN(n9486) );
  NAND2_X1 U5836 ( .A1(n4883), .A2(n4891), .ZN(n9500) );
  OR2_X1 U5837 ( .A1(n9518), .A2(n8289), .ZN(n4883) );
  NAND2_X1 U5838 ( .A1(n9543), .A2(n8309), .ZN(n9520) );
  INV_X1 U5839 ( .A(n9685), .ZN(n9539) );
  NAND2_X1 U5840 ( .A1(n4856), .A2(n4859), .ZN(n9549) );
  NAND2_X1 U5841 ( .A1(n8284), .A2(n4860), .ZN(n4856) );
  OAI21_X1 U5842 ( .B1(n8284), .B2(n4404), .A(n4864), .ZN(n9566) );
  NAND2_X1 U5843 ( .A1(n5320), .A2(n5319), .ZN(n9587) );
  NAND2_X1 U5844 ( .A1(n4630), .A2(n4629), .ZN(n9592) );
  NAND2_X1 U5845 ( .A1(n4894), .A2(n4898), .ZN(n8276) );
  NAND2_X1 U5846 ( .A1(n8128), .A2(n4899), .ZN(n4894) );
  NAND2_X1 U5847 ( .A1(n4636), .A2(n6045), .ZN(n8131) );
  INV_X1 U5848 ( .A(n8126), .ZN(n4900) );
  NAND2_X1 U5849 ( .A1(n8128), .A2(n8127), .ZN(n4901) );
  NAND2_X1 U5850 ( .A1(n7870), .A2(n7869), .ZN(n7982) );
  NAND2_X1 U5851 ( .A1(n7868), .A2(n7867), .ZN(n7870) );
  NAND2_X1 U5852 ( .A1(n7625), .A2(n4957), .ZN(n7626) );
  OAI21_X1 U5853 ( .B1(n7606), .B2(n4850), .A(n4848), .ZN(n7785) );
  AND3_X1 U5854 ( .A1(n5223), .A2(n5222), .A3(n5221), .ZN(n7610) );
  AND2_X1 U5855 ( .A1(n9652), .A2(n4345), .ZN(n9653) );
  INV_X1 U5856 ( .A(n9461), .ZN(n9741) );
  AOI211_X1 U5857 ( .C1(n9667), .C2(n9723), .A(n9666), .B(n9665), .ZN(n9742)
         );
  AND2_X1 U5858 ( .A1(n5159), .A2(n5158), .ZN(n9749) );
  NAND2_X1 U5859 ( .A1(n7999), .A2(n5342), .ZN(n5159) );
  AOI211_X1 U5860 ( .C1(n9672), .C2(n9723), .A(n9671), .B(n9670), .ZN(n9746)
         );
  INV_X1 U5861 ( .A(n9502), .ZN(n9753) );
  INV_X1 U5862 ( .A(n9558), .ZN(n9762) );
  INV_X1 U5863 ( .A(n9610), .ZN(n9772) );
  INV_X1 U5864 ( .A(n8274), .ZN(n9781) );
  NAND2_X1 U5865 ( .A1(n6883), .A2(n5342), .ZN(n5251) );
  XNOR2_X1 U5866 ( .A(n5142), .B(n5141), .ZN(n8191) );
  NAND2_X1 U5867 ( .A1(n4346), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5142) );
  NAND2_X1 U5868 ( .A1(n5311), .A2(n7177), .ZN(n5317) );
  NAND2_X1 U5869 ( .A1(n4797), .A2(n4387), .ZN(n5295) );
  INV_X1 U5870 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7166) );
  NAND2_X1 U5871 ( .A1(n4601), .A2(n4991), .ZN(n5202) );
  OR2_X1 U5872 ( .A1(n5173), .A2(n9788), .ZN(n5187) );
  NOR2_X1 U5873 ( .A1(n5174), .A2(n5173), .ZN(n9328) );
  NAND2_X1 U5874 ( .A1(n4918), .A2(n8664), .ZN(n4917) );
  CLKBUF_X1 U5875 ( .A(n7291), .Z(n7292) );
  NOR2_X1 U5876 ( .A1(n7226), .A2(n4529), .ZN(n7232) );
  XNOR2_X1 U5877 ( .A(n4514), .B(n5529), .ZN(n8517) );
  NAND2_X1 U5878 ( .A1(n8705), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4524) );
  INV_X1 U5879 ( .A(n4438), .ZN(n4437) );
  MUX2_X1 U5880 ( .A(n6518), .B(n6517), .S(n10222), .Z(n6519) );
  NOR2_X1 U5881 ( .A1(n6748), .A2(n6750), .ZN(n6783) );
  OAI21_X1 U5882 ( .B1(n6082), .B2(n6081), .A(n6080), .ZN(n6088) );
  NAND2_X1 U5883 ( .A1(n9419), .A2(n9418), .ZN(n4457) );
  NAND2_X1 U5884 ( .A1(n4617), .A2(n4616), .ZN(n4615) );
  MUX2_X1 U5885 ( .A(n5363), .B(n9644), .S(n10082), .Z(n9645) );
  NAND2_X1 U5886 ( .A1(n5940), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U5887 ( .A1(n5237), .A2(n5236), .ZN(n10012) );
  INV_X1 U5888 ( .A(n10012), .ZN(n4589) );
  INV_X2 U5889 ( .A(n6549), .ZN(n6545) );
  INV_X1 U5890 ( .A(n4530), .ZN(n10156) );
  NOR2_X1 U5891 ( .A1(n5027), .A2(n5026), .ZN(n4343) );
  AND2_X1 U5892 ( .A1(n4623), .A2(n5966), .ZN(n4344) );
  AND2_X1 U5893 ( .A1(n4603), .A2(n4393), .ZN(n4345) );
  NAND2_X1 U5894 ( .A1(n8339), .A2(n8338), .ZN(n8335) );
  AND2_X1 U5895 ( .A1(n8312), .A2(n5987), .ZN(n9487) );
  INV_X1 U5896 ( .A(n4329), .ZN(n5583) );
  NAND4_X1 U5897 ( .A1(n4580), .A2(n4953), .A3(n4905), .A4(n4402), .ZN(n4346)
         );
  AND2_X1 U5898 ( .A1(n4920), .A2(n4369), .ZN(n4347) );
  INV_X1 U5899 ( .A(n4713), .ZN(n4712) );
  NAND2_X1 U5900 ( .A1(n8430), .A2(n6404), .ZN(n4713) );
  NAND2_X1 U5901 ( .A1(n9655), .A2(n9189), .ZN(n5941) );
  NAND2_X1 U5902 ( .A1(n8330), .A2(n8333), .ZN(n7345) );
  AND2_X1 U5903 ( .A1(n8297), .A2(n4610), .ZN(n4348) );
  INV_X1 U5904 ( .A(n4865), .ZN(n4864) );
  NOR2_X1 U5905 ( .A1(n9767), .A2(n8283), .ZN(n4865) );
  INV_X1 U5906 ( .A(n4577), .ZN(n4576) );
  AND3_X1 U5907 ( .A1(n4448), .A2(n8406), .A3(n4447), .ZN(n4577) );
  NAND2_X1 U5908 ( .A1(n4385), .A2(n4863), .ZN(n4859) );
  AND2_X1 U5909 ( .A1(n4594), .A2(n4593), .ZN(n4349) );
  OR2_X1 U5910 ( .A1(n9625), .A2(n4587), .ZN(n4350) );
  AND2_X1 U5911 ( .A1(n4590), .A2(n4591), .ZN(n4351) );
  INV_X1 U5912 ( .A(n8764), .ZN(n10122) );
  AND2_X2 U5913 ( .A1(n6812), .A2(n6100), .ZN(n5182) );
  XOR2_X1 U5914 ( .A(n8822), .B(n8552), .Z(n4352) );
  NAND2_X1 U5915 ( .A1(n5126), .A2(n5125), .ZN(n5196) );
  OAI211_X1 U5916 ( .C1(n6215), .C2(n6859), .A(n6142), .B(n6141), .ZN(n10139)
         );
  INV_X2 U5917 ( .A(n6812), .ZN(n5204) );
  NAND4_X1 U5918 ( .A1(n6128), .A2(n6127), .A3(n6126), .A4(n6125), .ZN(n10131)
         );
  NAND2_X1 U5919 ( .A1(n4914), .A2(n4913), .ZN(n8593) );
  AND3_X1 U5920 ( .A1(n4905), .A2(n4953), .A3(n5126), .ZN(n5346) );
  OR2_X1 U5921 ( .A1(n4581), .A2(n4583), .ZN(n5367) );
  NAND2_X1 U5922 ( .A1(n8913), .A2(n6337), .ZN(n8900) );
  XNOR2_X1 U5923 ( .A(n6091), .B(n6090), .ZN(n6092) );
  INV_X1 U5924 ( .A(n5186), .ZN(n5218) );
  NOR2_X1 U5925 ( .A1(n5040), .A2(SI_16_), .ZN(n4353) );
  AND2_X1 U5926 ( .A1(n6137), .A2(n6138), .ZN(n4354) );
  AND2_X1 U5927 ( .A1(n8424), .A2(n8423), .ZN(n4355) );
  INV_X1 U5928 ( .A(n8297), .ZN(n8316) );
  AND2_X1 U5929 ( .A1(n6029), .A2(n5976), .ZN(n8297) );
  AND2_X1 U5930 ( .A1(n5867), .A2(n5866), .ZN(n4356) );
  OR2_X1 U5931 ( .A1(n5481), .A2(P2_IR_REG_6__SCAN_IN), .ZN(n4357) );
  OR2_X1 U5932 ( .A1(n9519), .A2(n4639), .ZN(n4358) );
  INV_X1 U5933 ( .A(n4485), .ZN(n4484) );
  NAND2_X1 U5934 ( .A1(n4487), .A2(n5306), .ZN(n4485) );
  OR2_X1 U5935 ( .A1(n9234), .A2(n4950), .ZN(n4819) );
  OR2_X1 U5936 ( .A1(n8809), .A2(n8806), .ZN(n4359) );
  AND4_X1 U5937 ( .A1(n5418), .A2(n5417), .A3(n5431), .A4(n5424), .ZN(n4360)
         );
  OR2_X1 U5938 ( .A1(n5252), .A2(n5027), .ZN(n4361) );
  NAND2_X1 U5939 ( .A1(n5148), .A2(n5147), .ZN(n9432) );
  INV_X1 U5940 ( .A(n9432), .ZN(n4472) );
  AND2_X1 U5941 ( .A1(n6100), .A2(n6847), .ZN(n4362) );
  INV_X1 U5942 ( .A(n8074), .ZN(n8486) );
  INV_X1 U5943 ( .A(n4950), .ZN(n4817) );
  NAND2_X1 U5944 ( .A1(n5466), .A2(n5399), .ZN(n5472) );
  AND2_X1 U5945 ( .A1(n5231), .A2(n5230), .ZN(n7697) );
  NOR2_X1 U5946 ( .A1(n5369), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n5365) );
  AND2_X1 U5947 ( .A1(n9728), .A2(n9309), .ZN(n4363) );
  INV_X1 U5948 ( .A(n9708), .ZN(n9604) );
  NAND2_X1 U5949 ( .A1(n5314), .A2(n5313), .ZN(n9708) );
  INV_X1 U5950 ( .A(n4578), .ZN(n9501) );
  NOR2_X1 U5951 ( .A1(n9524), .A2(n9502), .ZN(n4578) );
  OR2_X1 U5952 ( .A1(n4530), .A2(n4525), .ZN(n8346) );
  INV_X1 U5953 ( .A(n8346), .ZN(n4643) );
  NOR2_X1 U5954 ( .A1(n10117), .A2(n10116), .ZN(n4364) );
  OR2_X1 U5955 ( .A1(n9753), .A2(n8290), .ZN(n4365) );
  INV_X1 U5956 ( .A(n4669), .ZN(n4668) );
  OR2_X1 U5957 ( .A1(n6464), .A2(n4670), .ZN(n4669) );
  AND2_X1 U5958 ( .A1(n8407), .A2(n8410), .ZN(n8954) );
  AND2_X1 U5959 ( .A1(n4843), .A2(n4842), .ZN(n4366) );
  NAND2_X1 U5960 ( .A1(n5281), .A2(n5280), .ZN(n9728) );
  AND2_X1 U5961 ( .A1(n7697), .A2(n5744), .ZN(n4367) );
  AND3_X1 U5962 ( .A1(n5200), .A2(n5199), .A3(n5198), .ZN(n7431) );
  INV_X1 U5963 ( .A(n9487), .ZN(n4625) );
  AND2_X1 U5964 ( .A1(n8389), .A2(n8390), .ZN(n4368) );
  INV_X1 U5965 ( .A(n7876), .ZN(n7869) );
  AND2_X1 U5966 ( .A1(n6000), .A2(n8226), .ZN(n7876) );
  OR2_X1 U5967 ( .A1(n4352), .A2(n4919), .ZN(n4369) );
  INV_X1 U5968 ( .A(n7593), .ZN(n7498) );
  AND3_X1 U5969 ( .A1(n5208), .A2(n5207), .A3(n5206), .ZN(n7593) );
  INV_X1 U5970 ( .A(n6369), .ZN(n4692) );
  INV_X1 U5971 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4463) );
  INV_X1 U5972 ( .A(n4879), .ZN(n4878) );
  NAND2_X1 U5973 ( .A1(n4880), .A2(n4365), .ZN(n4879) );
  NOR2_X1 U5974 ( .A1(n9070), .A2(n8845), .ZN(n4370) );
  NOR2_X1 U5975 ( .A1(n9313), .A2(n9862), .ZN(n4371) );
  INV_X1 U5976 ( .A(n4600), .ZN(n9439) );
  NOR2_X1 U5977 ( .A1(n9458), .A2(n9655), .ZN(n4600) );
  INV_X1 U5978 ( .A(n4612), .ZN(n4611) );
  OR2_X1 U5979 ( .A1(n8315), .A2(n5989), .ZN(n4612) );
  AND2_X1 U5980 ( .A1(n4993), .A2(SI_4_), .ZN(n4372) );
  AND2_X1 U5981 ( .A1(n4964), .A2(n8463), .ZN(n4373) );
  INV_X1 U5982 ( .A(n4945), .ZN(n4943) );
  NAND2_X1 U5983 ( .A1(n5402), .A2(n4946), .ZN(n4945) );
  INV_X1 U5984 ( .A(n7482), .ZN(n10133) );
  AND4_X1 U5985 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n7482)
         );
  NAND2_X1 U5986 ( .A1(n4940), .A2(n4944), .ZN(n4374) );
  INV_X1 U5987 ( .A(n7582), .ZN(n7602) );
  AND2_X1 U5988 ( .A1(n5035), .A2(SI_14_), .ZN(n4375) );
  OR2_X1 U5989 ( .A1(n5461), .A2(n6434), .ZN(n4376) );
  NOR2_X1 U5990 ( .A1(n8536), .A2(n8933), .ZN(n8595) );
  AND2_X1 U5991 ( .A1(n4574), .A2(n4568), .ZN(n4377) );
  NAND2_X1 U5992 ( .A1(n4969), .A2(n8832), .ZN(n4378) );
  INV_X1 U5993 ( .A(n4753), .ZN(n4570) );
  AND2_X1 U5994 ( .A1(n8924), .A2(n8407), .ZN(n4753) );
  AND2_X1 U5995 ( .A1(n5030), .A2(SI_12_), .ZN(n4379) );
  OR2_X1 U5996 ( .A1(n9745), .A2(n8293), .ZN(n4380) );
  NOR2_X1 U5997 ( .A1(n8277), .A2(n9781), .ZN(n4381) );
  INV_X1 U5998 ( .A(n9757), .ZN(n9527) );
  AND2_X1 U5999 ( .A1(n5163), .A2(n5162), .ZN(n9757) );
  NAND2_X1 U6000 ( .A1(n8702), .A2(n7861), .ZN(n4382) );
  OR2_X1 U6001 ( .A1(n8126), .A2(n4363), .ZN(n4383) );
  AND2_X1 U6002 ( .A1(n4607), .A2(n9636), .ZN(n4384) );
  NAND2_X1 U6003 ( .A1(n9565), .A2(n4861), .ZN(n4385) );
  INV_X1 U6004 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5141) );
  INV_X1 U6005 ( .A(n8699), .ZN(n8960) );
  AND4_X1 U6006 ( .A1(n5404), .A2(n5503), .A3(n7025), .A4(n5403), .ZN(n4386)
         );
  OR2_X1 U6007 ( .A1(n9502), .A2(n8290), .ZN(n8311) );
  OR2_X1 U6008 ( .A1(n9143), .A2(n8182), .ZN(n8392) );
  INV_X1 U6009 ( .A(n8392), .ZN(n4655) );
  AND2_X1 U6010 ( .A1(n5293), .A2(n5292), .ZN(n4387) );
  AND3_X1 U6011 ( .A1(n5404), .A2(n7025), .A3(n5408), .ZN(n4388) );
  AND2_X1 U6012 ( .A1(n5719), .A2(n5932), .ZN(n4389) );
  AND2_X1 U6013 ( .A1(n7701), .A2(n8371), .ZN(n4390) );
  AND2_X1 U6014 ( .A1(n8496), .A2(n6369), .ZN(n4391) );
  NOR2_X1 U6015 ( .A1(n8508), .A2(n8507), .ZN(n4392) );
  OR2_X1 U6016 ( .A1(n9451), .A2(n4602), .ZN(n4393) );
  XNOR2_X1 U6017 ( .A(n5029), .B(SI_12_), .ZN(n5262) );
  NAND2_X1 U6018 ( .A1(n8493), .A2(n8399), .ZN(n4394) );
  NAND2_X1 U6019 ( .A1(n7364), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n4395) );
  AND2_X1 U6020 ( .A1(n8316), .A2(n4611), .ZN(n4396) );
  AND3_X1 U6021 ( .A1(n6105), .A2(n6104), .A3(n6103), .ZN(n7352) );
  INV_X1 U6022 ( .A(n7352), .ZN(n6106) );
  AND2_X1 U6023 ( .A1(n4702), .A2(n6090), .ZN(n4397) );
  AND2_X1 U6024 ( .A1(n4349), .A2(n8192), .ZN(n4398) );
  AND2_X1 U6025 ( .A1(n4380), .A2(n4885), .ZN(n4399) );
  AND2_X1 U6026 ( .A1(n8436), .A2(n8830), .ZN(n4400) );
  AND2_X1 U6027 ( .A1(n4737), .A2(n4736), .ZN(n4401) );
  AND2_X1 U6028 ( .A1(n4582), .A2(n4463), .ZN(n4402) );
  INV_X1 U6029 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9152) );
  BUF_X1 U6030 ( .A(n6131), .Z(n6310) );
  XNOR2_X1 U6031 ( .A(n5473), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6140) );
  INV_X1 U6032 ( .A(n6140), .ZN(n4742) );
  OR2_X1 U6033 ( .A1(n5063), .A2(SI_21_), .ZN(n4403) );
  INV_X1 U6034 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4703) );
  NOR2_X1 U6035 ( .A1(n9587), .A2(n9304), .ZN(n4404) );
  INV_X1 U6036 ( .A(n9312), .ZN(n7983) );
  AND2_X1 U6037 ( .A1(n5282), .A2(SI_15_), .ZN(n4405) );
  NAND2_X1 U6038 ( .A1(n4866), .A2(n4869), .ZN(n8223) );
  NAND2_X1 U6039 ( .A1(n4656), .A2(n8392), .ZN(n8985) );
  NAND2_X1 U6040 ( .A1(n4658), .A2(n6460), .ZN(n8874) );
  AND2_X1 U6041 ( .A1(n9558), .A2(n9302), .ZN(n4406) );
  NOR3_X1 U6042 ( .A1(n9625), .A2(n4587), .A3(n9697), .ZN(n4585) );
  NOR2_X1 U6043 ( .A1(n10092), .A2(n5495), .ZN(n4407) );
  NAND2_X1 U6044 ( .A1(n8308), .A2(n8307), .ZN(n4408) );
  AND2_X1 U6045 ( .A1(n4838), .A2(n4837), .ZN(n4409) );
  AND2_X1 U6046 ( .A1(n4501), .A2(n5160), .ZN(n4410) );
  NAND2_X1 U6047 ( .A1(n6669), .A2(n6670), .ZN(n6673) );
  OR2_X1 U6048 ( .A1(n8715), .A2(n10240), .ZN(n4838) );
  OR2_X1 U6049 ( .A1(n9741), .A2(n9280), .ZN(n4411) );
  AND4_X1 U6050 ( .A1(n5742), .A2(n5741), .A3(n5740), .A4(n5739), .ZN(n7788)
         );
  AND2_X1 U6051 ( .A1(n4801), .A2(n6673), .ZN(n4412) );
  AND4_X1 U6052 ( .A1(n5752), .A2(n5751), .A3(n5750), .A4(n5749), .ZN(n7881)
         );
  INV_X1 U6053 ( .A(n8285), .ZN(n4863) );
  AND2_X1 U6054 ( .A1(n9697), .A2(n9303), .ZN(n8285) );
  NOR2_X1 U6055 ( .A1(n9685), .A2(n9301), .ZN(n4413) );
  NAND2_X1 U6056 ( .A1(n8663), .A2(n8662), .ZN(n4414) );
  AND2_X1 U6057 ( .A1(n5144), .A2(n5143), .ZN(n9646) );
  INV_X1 U6058 ( .A(n9646), .ZN(n5940) );
  AND2_X1 U6059 ( .A1(n5052), .A2(SI_18_), .ZN(n4415) );
  OR2_X1 U6060 ( .A1(n5164), .A2(n4502), .ZN(n4416) );
  OR2_X1 U6061 ( .A1(n9090), .A2(n8877), .ZN(n4417) );
  AND2_X1 U6062 ( .A1(n4901), .A2(n4900), .ZN(n4418) );
  AND2_X1 U6063 ( .A1(n4403), .A2(n5070), .ZN(n4419) );
  INV_X1 U6064 ( .A(n10023), .ZN(n10045) );
  INV_X1 U6065 ( .A(n10020), .ZN(n4616) );
  INV_X1 U6066 ( .A(n9173), .ZN(n4818) );
  NAND2_X1 U6067 ( .A1(n4774), .A2(n7236), .ZN(n6981) );
  AND2_X1 U6068 ( .A1(n8235), .A2(n4349), .ZN(n4420) );
  NAND2_X1 U6069 ( .A1(n10127), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n4421) );
  INV_X1 U6070 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5292) );
  NAND2_X1 U6071 ( .A1(n4644), .A2(n8346), .ZN(n7490) );
  AND2_X1 U6072 ( .A1(n5456), .A2(n5455), .ZN(n8714) );
  NAND2_X1 U6073 ( .A1(n7792), .A2(n7798), .ZN(n7868) );
  NOR2_X1 U6074 ( .A1(n7823), .A2(n5488), .ZN(n4422) );
  AND2_X1 U6075 ( .A1(n4833), .A2(n4832), .ZN(n4423) );
  INV_X1 U6076 ( .A(n9596), .ZN(n9636) );
  AND2_X1 U6077 ( .A1(n7529), .A2(n7533), .ZN(n4424) );
  AND2_X1 U6078 ( .A1(n6228), .A2(n6227), .ZN(n4425) );
  INV_X1 U6079 ( .A(n8176), .ZN(n4939) );
  NAND2_X1 U6080 ( .A1(n5273), .A2(n5272), .ZN(n8163) );
  INV_X1 U6081 ( .A(n8163), .ZN(n4593) );
  INV_X1 U6082 ( .A(n5529), .ZN(n8509) );
  NAND2_X1 U6083 ( .A1(n7333), .A2(n7332), .ZN(n7336) );
  OR2_X1 U6084 ( .A1(n7463), .A2(n7498), .ZN(n7503) );
  INV_X1 U6085 ( .A(n7503), .ZN(n4590) );
  INV_X1 U6086 ( .A(n8789), .ZN(n4845) );
  INV_X1 U6087 ( .A(n7216), .ZN(n8329) );
  INV_X1 U6088 ( .A(n4579), .ZN(n7648) );
  NAND2_X1 U6089 ( .A1(n10050), .A2(n7649), .ZN(n4579) );
  OR2_X1 U6090 ( .A1(n5568), .A2(n5525), .ZN(n4426) );
  NAND2_X1 U6091 ( .A1(n8755), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4427) );
  OR2_X1 U6092 ( .A1(n4729), .A2(n4728), .ZN(n4428) );
  INV_X1 U6093 ( .A(n9418), .ZN(n7570) );
  INV_X1 U6094 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n4536) );
  INV_X1 U6095 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n4543) );
  INV_X1 U6096 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n4541) );
  INV_X1 U6097 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n4540) );
  INV_X1 U6098 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n4537) );
  XNOR2_X1 U6099 ( .A(n5487), .B(n7828), .ZN(n7824) );
  XNOR2_X1 U6100 ( .A(n5554), .B(n6977), .ZN(n8729) );
  XNOR2_X1 U6101 ( .A(n5500), .B(n6977), .ZN(n8727) );
  AOI21_X1 U6102 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n10127), .A(n10110), .ZN(
        n5500) );
  NAND2_X1 U6103 ( .A1(n8403), .A2(n8458), .ZN(n4447) );
  NAND2_X1 U6104 ( .A1(n4429), .A2(n5746), .ZN(n5755) );
  NAND3_X1 U6105 ( .A1(n5732), .A2(n5733), .A3(n7795), .ZN(n4429) );
  MUX2_X2 U6106 ( .A(n5827), .B(n5826), .S(n6075), .Z(n5831) );
  INV_X1 U6107 ( .A(n5719), .ZN(n7634) );
  OR2_X1 U6108 ( .A1(n5975), .A2(n5974), .ZN(n6035) );
  NOR2_X1 U6109 ( .A1(n5887), .A2(n5886), .ZN(n5908) );
  OAI211_X1 U6110 ( .C1(n5868), .C2(n6075), .A(n5869), .B(n4440), .ZN(n5883)
         );
  NAND2_X1 U6111 ( .A1(n4804), .A2(n4803), .ZN(n4802) );
  AOI21_X1 U6112 ( .B1(n5017), .B2(n4765), .A(n4343), .ZN(n5263) );
  NAND2_X1 U6113 ( .A1(n9263), .A2(n6705), .ZN(n9260) );
  NAND2_X1 U6114 ( .A1(n4778), .A2(n4430), .ZN(n7923) );
  INV_X1 U6115 ( .A(n4431), .ZN(n4430) );
  OAI21_X1 U6116 ( .B1(n4783), .B2(n4781), .A(n7925), .ZN(n4431) );
  NOR2_X1 U6117 ( .A1(n9957), .A2(n8199), .ZN(n9956) );
  XNOR2_X1 U6118 ( .A(n9388), .B(n9409), .ZN(n9957) );
  NAND2_X1 U6119 ( .A1(n9414), .A2(n4455), .ZN(n4454) );
  NAND2_X1 U6120 ( .A1(n4457), .A2(n4453), .ZN(n9420) );
  OAI21_X1 U6121 ( .B1(n9415), .B2(n9999), .A(n9974), .ZN(n4456) );
  NAND3_X1 U6122 ( .A1(n5622), .A2(n5623), .A3(n4437), .ZN(P2_U3201) );
  AOI22_X2 U6123 ( .A1(n8526), .A2(n8699), .B1(n8525), .B2(n8524), .ZN(n8622)
         );
  NOR2_X1 U6124 ( .A1(n8689), .A2(n8690), .ZN(n8687) );
  NAND2_X1 U6125 ( .A1(n4806), .A2(n4805), .ZN(n9263) );
  INV_X1 U6126 ( .A(n5253), .ZN(n4464) );
  NAND2_X1 U6127 ( .A1(n4464), .A2(n5244), .ZN(n5255) );
  NOR2_X2 U6128 ( .A1(n9227), .A2(n9226), .ZN(n9237) );
  AOI21_X2 U6129 ( .B1(n6638), .B2(n6637), .A(n4784), .ZN(n4783) );
  NAND2_X1 U6130 ( .A1(n5953), .A2(n7258), .ZN(n5675) );
  NAND2_X1 U6131 ( .A1(n7465), .A2(n5698), .ZN(n5724) );
  NAND2_X1 U6132 ( .A1(n7505), .A2(n4389), .ZN(n5733) );
  NAND2_X1 U6133 ( .A1(n5779), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U6134 ( .A1(n4444), .A2(n4441), .ZN(n5780) );
  NAND2_X2 U6135 ( .A1(n5724), .A2(n5950), .ZN(n7505) );
  NAND2_X1 U6136 ( .A1(n4460), .A2(n5951), .ZN(n7465) );
  INV_X1 U6137 ( .A(n5126), .ZN(n5194) );
  AND2_X2 U6138 ( .A1(n5136), .A2(n5126), .ZN(n4580) );
  OR2_X1 U6139 ( .A1(n5859), .A2(n5858), .ZN(n5868) );
  MUX2_X2 U6140 ( .A(n6071), .B(n6070), .S(n9418), .Z(n6082) );
  NAND2_X1 U6141 ( .A1(n4762), .A2(n4761), .ZN(n5268) );
  NOR2_X1 U6142 ( .A1(n4567), .A2(n4575), .ZN(n4568) );
  NAND2_X1 U6143 ( .A1(n4515), .A2(n4392), .ZN(n4514) );
  NAND2_X1 U6144 ( .A1(n4572), .A2(n4569), .ZN(n4752) );
  NAND2_X1 U6145 ( .A1(n4768), .A2(n4767), .ZN(n8423) );
  NAND2_X1 U6146 ( .A1(n4555), .A2(n4754), .ZN(n4554) );
  OAI21_X1 U6147 ( .B1(n4758), .B2(n4757), .A(n8458), .ZN(n4756) );
  NOR2_X2 U6148 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  OAI21_X2 U6149 ( .B1(n10099), .B2(n4828), .A(n4827), .ZN(n5554) );
  NAND2_X1 U6150 ( .A1(n5560), .A2(n4845), .ZN(n4840) );
  NAND2_X1 U6151 ( .A1(n5543), .A2(n5542), .ZN(n7367) );
  NAND2_X1 U6152 ( .A1(n5549), .A2(n4839), .ZN(n4835) );
  NAND2_X1 U6153 ( .A1(n5547), .A2(n4834), .ZN(n4830) );
  NOR2_X1 U6154 ( .A1(n5539), .A2(n6165), .ZN(n7365) );
  AOI21_X2 U6155 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n7898), .A(n7902), .ZN(
        n5490) );
  NAND2_X1 U6156 ( .A1(n7293), .A2(n7218), .ZN(n7228) );
  AOI21_X2 U6157 ( .B1(n8632), .B2(n8548), .A(n4959), .ZN(n8606) );
  INV_X1 U6158 ( .A(n7309), .ZN(n4460) );
  NAND2_X1 U6159 ( .A1(n5823), .A2(n4458), .ZN(n5825) );
  AOI21_X1 U6160 ( .B1(n4459), .B2(n5857), .A(n5984), .ZN(n5859) );
  NAND2_X1 U6161 ( .A1(n5755), .A2(n5754), .ZN(n5777) );
  NAND2_X2 U6162 ( .A1(n5140), .A2(n5139), .ZN(n8217) );
  NAND3_X1 U6163 ( .A1(n5851), .A2(n6054), .A3(n6056), .ZN(n4459) );
  NAND2_X2 U6164 ( .A1(n8597), .A2(n4951), .ZN(n8649) );
  NAND3_X1 U6165 ( .A1(n8273), .A2(n8272), .A3(n4411), .ZN(P1_U3214) );
  NAND2_X1 U6166 ( .A1(n6671), .A2(n6672), .ZN(n4804) );
  OR2_X1 U6167 ( .A1(n7211), .A2(n10154), .ZN(n7212) );
  NAND2_X1 U6168 ( .A1(n7923), .A2(n6656), .ZN(n6662) );
  AOI22_X2 U6169 ( .A1(n6636), .A2(n6635), .B1(n6634), .B2(n9857), .ZN(n6637)
         );
  INV_X1 U6170 ( .A(n6662), .ZN(n6665) );
  NAND2_X1 U6171 ( .A1(n6736), .A2(n6735), .ZN(n9247) );
  MUX2_X2 U6172 ( .A(n5782), .B(n5781), .S(n5932), .Z(n5822) );
  AOI21_X1 U6173 ( .B1(n6073), .B2(n6969), .A(n7726), .ZN(n5975) );
  NOR2_X1 U6174 ( .A1(n9956), .A2(n9389), .ZN(n9968) );
  NAND2_X1 U6175 ( .A1(n5157), .A2(n5156), .ZN(n4465) );
  NAND2_X1 U6176 ( .A1(n5333), .A2(n5332), .ZN(n4466) );
  NAND2_X1 U6177 ( .A1(n4468), .A2(n4471), .ZN(n4467) );
  NAND2_X1 U6178 ( .A1(n5939), .A2(n4472), .ZN(n4468) );
  NAND2_X1 U6179 ( .A1(n4476), .A2(n4473), .ZN(n6073) );
  NAND2_X1 U6180 ( .A1(n5291), .A2(n4480), .ZN(n4479) );
  NAND3_X1 U6181 ( .A1(n4482), .A2(n4485), .A3(n4481), .ZN(n4478) );
  NAND2_X1 U6182 ( .A1(n5210), .A2(n5209), .ZN(n4998) );
  OAI21_X2 U6183 ( .B1(n4601), .B2(n4493), .A(n4491), .ZN(n5210) );
  NAND2_X1 U6184 ( .A1(n5268), .A2(n4497), .ZN(n4494) );
  NAND2_X1 U6185 ( .A1(n4494), .A2(n4495), .ZN(n5284) );
  NAND3_X1 U6186 ( .A1(n5061), .A2(n5060), .A3(n4419), .ZN(n4500) );
  NAND3_X1 U6187 ( .A1(n5061), .A2(n5060), .A3(n4403), .ZN(n4503) );
  NAND2_X1 U6188 ( .A1(n5061), .A2(n5060), .ZN(n5329) );
  NAND2_X1 U6189 ( .A1(n5096), .A2(n4507), .ZN(n4504) );
  OAI21_X1 U6190 ( .B1(n5096), .B2(n4510), .A(n4507), .ZN(n5340) );
  NAND2_X1 U6191 ( .A1(n4504), .A2(n4505), .ZN(n5107) );
  AND2_X1 U6192 ( .A1(n4386), .A2(n5405), .ZN(n4522) );
  NAND4_X1 U6193 ( .A1(n4523), .A2(n4521), .A3(n4518), .A4(n4388), .ZN(n5409)
         );
  NAND2_X1 U6194 ( .A1(n4525), .A2(n10156), .ZN(n4965) );
  NAND2_X1 U6195 ( .A1(n4530), .A2(n10139), .ZN(n6143) );
  OAI21_X1 U6196 ( .B1(n10156), .B2(n8705), .A(n4524), .ZN(P2_U3494) );
  XNOR2_X1 U6197 ( .A(n4525), .B(n10156), .ZN(n10137) );
  INV_X1 U6198 ( .A(n10139), .ZN(n4525) );
  NAND2_X1 U6199 ( .A1(n4525), .A2(n4530), .ZN(n8360) );
  NAND2_X1 U6200 ( .A1(n7331), .A2(n4530), .ZN(n7332) );
  XNOR2_X1 U6201 ( .A(n7330), .B(n4530), .ZN(n7221) );
  NAND2_X1 U6202 ( .A1(n10130), .A2(n4530), .ZN(n4528) );
  AND2_X1 U6203 ( .A1(n8683), .A2(n4530), .ZN(n4529) );
  NAND2_X1 U6204 ( .A1(n4535), .A2(n6092), .ZN(n6115) );
  AND2_X1 U6205 ( .A1(n6093), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4535) );
  OR2_X1 U6206 ( .A1(n6149), .A2(n7424), .ZN(n6099) );
  OR2_X1 U6207 ( .A1(n6149), .A2(n4544), .ZN(n6440) );
  NAND3_X1 U6208 ( .A1(n4546), .A2(n8384), .A3(n8383), .ZN(n4545) );
  NAND3_X1 U6209 ( .A1(n4551), .A2(n4548), .A3(n4547), .ZN(n4546) );
  NAND2_X1 U6210 ( .A1(n4400), .A2(n4554), .ZN(n8440) );
  NAND2_X1 U6211 ( .A1(n4940), .A2(n4687), .ZN(n5442) );
  NAND3_X1 U6212 ( .A1(n4940), .A2(n4687), .A3(n4702), .ZN(n4565) );
  OR2_X1 U6213 ( .A1(n8400), .A2(n4576), .ZN(n4574) );
  INV_X1 U6214 ( .A(n8954), .ZN(n4575) );
  NAND2_X1 U6215 ( .A1(n8400), .A2(n4573), .ZN(n4572) );
  INV_X1 U6216 ( .A(n7436), .ZN(n10034) );
  NAND3_X1 U6217 ( .A1(n4580), .A2(n4953), .A3(n4905), .ZN(n5369) );
  CLKBUF_X1 U6218 ( .A(n5369), .Z(n4581) );
  INV_X1 U6219 ( .A(n4585), .ZN(n9571) );
  NAND2_X1 U6220 ( .A1(n9476), .A2(n4596), .ZN(n9429) );
  NAND2_X1 U6221 ( .A1(n9476), .A2(n9741), .ZN(n9458) );
  NAND2_X1 U6222 ( .A1(n5192), .A2(n5191), .ZN(n4601) );
  NAND2_X1 U6223 ( .A1(n9451), .A2(n8314), .ZN(n9444) );
  NAND2_X1 U6224 ( .A1(n5225), .A2(n5003), .ZN(n4613) );
  NAND2_X1 U6225 ( .A1(n5217), .A2(n5216), .ZN(n4614) );
  NAND2_X1 U6226 ( .A1(n8321), .A2(n4615), .ZN(P1_U3356) );
  NAND2_X1 U6227 ( .A1(n9510), .A2(n4344), .ZN(n4618) );
  NAND2_X1 U6228 ( .A1(n4618), .A2(n4619), .ZN(n9452) );
  OAI21_X1 U6229 ( .B1(n9635), .B2(n4628), .A(n4626), .ZN(n6055) );
  OAI21_X1 U6230 ( .B1(n8095), .B2(n4634), .A(n4631), .ZN(n6050) );
  OAI21_X1 U6231 ( .B1(n8308), .B2(n4358), .A(n4637), .ZN(n9508) );
  NAND2_X1 U6232 ( .A1(n4641), .A2(n4644), .ZN(n7476) );
  NAND2_X1 U6233 ( .A1(n8121), .A2(n4648), .ZN(n4647) );
  NAND2_X1 U6234 ( .A1(n8882), .A2(n8322), .ZN(n4658) );
  NAND2_X1 U6235 ( .A1(n8858), .A2(n4663), .ZN(n4661) );
  NAND2_X1 U6236 ( .A1(n7961), .A2(n4675), .ZN(n4674) );
  NAND2_X1 U6237 ( .A1(n8953), .A2(n4679), .ZN(n4971) );
  AOI21_X1 U6238 ( .B1(n7702), .B2(n4390), .A(n4682), .ZN(n7760) );
  NAND2_X1 U6239 ( .A1(n5442), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5443) );
  NAND3_X1 U6240 ( .A1(n4688), .A2(n4965), .A3(n6130), .ZN(n6144) );
  NAND2_X1 U6241 ( .A1(n6358), .A2(n4391), .ZN(n4689) );
  NAND2_X1 U6242 ( .A1(n4689), .A2(n4690), .ZN(n8862) );
  OAI21_X1 U6243 ( .B1(n7492), .B2(n4697), .A(n4694), .ZN(n4701) );
  NAND2_X1 U6244 ( .A1(n5420), .A2(n4397), .ZN(n9153) );
  NAND2_X1 U6245 ( .A1(n8851), .A2(n4710), .ZN(n4709) );
  NAND2_X1 U6246 ( .A1(n8851), .A2(n6394), .ZN(n4714) );
  OAI21_X2 U6247 ( .B1(n8957), .B2(n4717), .A(n4715), .ZN(n8913) );
  NAND2_X1 U6248 ( .A1(n6471), .A2(n6470), .ZN(n8813) );
  XNOR2_X1 U6249 ( .A(n9321), .B(n10050), .ZN(n7652) );
  NAND2_X1 U6250 ( .A1(n6382), .A2(n4417), .ZN(n8851) );
  AOI21_X1 U6251 ( .B1(n6450), .B2(n10135), .A(n6449), .ZN(n6471) );
  NAND2_X1 U6252 ( .A1(n5475), .A2(n6165), .ZN(n4730) );
  INV_X1 U6253 ( .A(n5475), .ZN(n4731) );
  NAND3_X1 U6254 ( .A1(n4733), .A2(n4732), .A3(n4427), .ZN(n5514) );
  INV_X1 U6255 ( .A(n4737), .ZN(n8726) );
  INV_X1 U6256 ( .A(n7903), .ZN(n4740) );
  NOR2_X1 U6257 ( .A1(n4743), .A2(n4742), .ZN(n4741) );
  NAND2_X1 U6258 ( .A1(n4745), .A2(n4744), .ZN(n4743) );
  NAND2_X1 U6259 ( .A1(n4329), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4744) );
  INV_X1 U6260 ( .A(n6787), .ZN(n4745) );
  NAND2_X1 U6261 ( .A1(n5017), .A2(n4763), .ZN(n4762) );
  NAND3_X1 U6262 ( .A1(n8419), .A2(n4770), .A3(n4769), .ZN(n4768) );
  NAND4_X1 U6263 ( .A1(n8416), .A2(n8458), .A3(n8897), .A4(n8415), .ZN(n4769)
         );
  NAND2_X1 U6264 ( .A1(n8402), .A2(n8401), .ZN(n8404) );
  NAND2_X1 U6265 ( .A1(n7197), .A2(n8451), .ZN(n4773) );
  NAND2_X1 U6266 ( .A1(n4775), .A2(n7236), .ZN(n6555) );
  NAND3_X1 U6267 ( .A1(n6534), .A2(n6543), .A3(n6544), .ZN(n4775) );
  NAND2_X1 U6268 ( .A1(n4779), .A2(n9856), .ZN(n4778) );
  OAI21_X1 U6269 ( .B1(n9856), .B2(n4777), .A(n4776), .ZN(n7924) );
  AOI21_X1 U6270 ( .B1(n4783), .B2(n4782), .A(n4781), .ZN(n4776) );
  INV_X1 U6271 ( .A(n4783), .ZN(n4777) );
  NOR2_X1 U6272 ( .A1(n4782), .A2(n4781), .ZN(n4779) );
  NAND2_X1 U6273 ( .A1(n4780), .A2(n4783), .ZN(n9867) );
  NAND2_X1 U6274 ( .A1(n9856), .A2(n6637), .ZN(n4780) );
  INV_X1 U6275 ( .A(n6648), .ZN(n4781) );
  INV_X1 U6276 ( .A(n6637), .ZN(n4782) );
  OAI21_X1 U6277 ( .B1(n9856), .B2(n6638), .A(n6637), .ZN(n9868) );
  NAND2_X1 U6278 ( .A1(n5311), .A2(n4794), .ZN(n4785) );
  OR2_X1 U6279 ( .A1(n5311), .A2(n4795), .ZN(n4786) );
  NAND3_X1 U6280 ( .A1(n4786), .A2(n4785), .A3(n4792), .ZN(n6521) );
  NAND2_X1 U6281 ( .A1(n5311), .A2(n4788), .ZN(n4787) );
  AND2_X1 U6282 ( .A1(n4792), .A2(n4789), .ZN(n4788) );
  OR2_X1 U6283 ( .A1(n5311), .A2(n4791), .ZN(n4790) );
  NAND2_X1 U6284 ( .A1(n4792), .A2(n4795), .ZN(n4791) );
  NAND2_X1 U6285 ( .A1(n4797), .A2(n4796), .ZN(n5303) );
  OAI21_X1 U6286 ( .B1(n6583), .B2(n4800), .A(n4799), .ZN(n7715) );
  AND2_X2 U6287 ( .A1(n4802), .A2(n6673), .ZN(n9227) );
  NAND2_X1 U6288 ( .A1(n9237), .A2(n4807), .ZN(n4806) );
  INV_X1 U6289 ( .A(n4819), .ZN(n9171) );
  OR2_X1 U6290 ( .A1(n9235), .A2(n9236), .ZN(n4820) );
  NAND2_X1 U6291 ( .A1(n9216), .A2(n9217), .ZN(n6752) );
  OAI21_X1 U6292 ( .B1(n9216), .B2(n4824), .A(n4821), .ZN(n9194) );
  NAND2_X1 U6293 ( .A1(n6751), .A2(n4823), .ZN(n4822) );
  INV_X1 U6294 ( .A(n9217), .ZN(n4823) );
  INV_X1 U6295 ( .A(n6751), .ZN(n4824) );
  XNOR2_X1 U6296 ( .A(n5546), .B(n7828), .ZN(n7827) );
  OAI21_X1 U6297 ( .B1(n5559), .B2(n4841), .A(n4840), .ZN(n8788) );
  INV_X1 U6298 ( .A(n5559), .ZN(n4844) );
  NAND2_X1 U6299 ( .A1(n7606), .A2(n4848), .ZN(n4847) );
  OAI21_X1 U6300 ( .B1(n8284), .B2(n4855), .A(n4853), .ZN(n9534) );
  NAND2_X1 U6301 ( .A1(n4852), .A2(n4851), .ZN(n8288) );
  NAND2_X1 U6302 ( .A1(n8284), .A2(n4853), .ZN(n4852) );
  NAND2_X1 U6303 ( .A1(n7792), .A2(n4867), .ZN(n4866) );
  NAND2_X1 U6304 ( .A1(n9518), .A2(n4875), .ZN(n4873) );
  NAND2_X1 U6305 ( .A1(n9518), .A2(n4881), .ZN(n4874) );
  NAND2_X2 U6306 ( .A1(n7222), .A2(n7221), .ZN(n7333) );
  AND4_X2 U6307 ( .A1(n5466), .A2(n5400), .A3(n5399), .A4(n4910), .ZN(n5476)
         );
  NAND3_X1 U6308 ( .A1(n5400), .A2(n5466), .A3(n5399), .ZN(n5464) );
  NAND2_X1 U6309 ( .A1(n4911), .A2(n4912), .ZN(n8537) );
  NAND2_X1 U6310 ( .A1(n8583), .A2(n4913), .ZN(n4911) );
  NAND2_X1 U6311 ( .A1(n8569), .A2(n4916), .ZN(n4915) );
  OAI211_X1 U6312 ( .C1(n8569), .C2(n4917), .A(n8564), .B(n4915), .ZN(P2_U3160) );
  OR2_X2 U6313 ( .A1(n8569), .A2(n8570), .ZN(n8571) );
  OAI21_X2 U6314 ( .B1(n8083), .B2(n4930), .A(n4928), .ZN(n8689) );
  NAND2_X1 U6315 ( .A1(n8148), .A2(n8182), .ZN(n4938) );
  AND2_X1 U6316 ( .A1(n5536), .A2(n6140), .ZN(n5537) );
  CLKBUF_X1 U6317 ( .A(n7443), .Z(n7337) );
  NAND2_X1 U6318 ( .A1(n8090), .A2(n8089), .ZN(n8093) );
  NAND2_X2 U6319 ( .A1(n6467), .A2(n7207), .ZN(n7209) );
  INV_X1 U6320 ( .A(n5359), .ZN(n5634) );
  XNOR2_X2 U6321 ( .A(n4334), .B(n8543), .ZN(n8577) );
  NAND2_X2 U6322 ( .A1(n8072), .A2(n8071), .ZN(n8083) );
  NOR2_X1 U6323 ( .A1(n6615), .A2(n7812), .ZN(n4947) );
  AND2_X1 U6324 ( .A1(n8584), .A2(n8943), .ZN(n4948) );
  INV_X1 U6325 ( .A(n6771), .ZN(n6080) );
  AND2_X1 U6326 ( .A1(n8523), .A2(n8978), .ZN(n4949) );
  AND2_X1 U6327 ( .A1(n6687), .A2(n6686), .ZN(n4950) );
  OR2_X1 U6328 ( .A1(n8539), .A2(n8917), .ZN(n4951) );
  INV_X1 U6329 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5402) );
  AND4_X1 U6330 ( .A1(n5134), .A2(n5133), .A3(n5132), .A4(n5131), .ZN(n4953)
         );
  OR2_X1 U6331 ( .A1(n8092), .A2(n8091), .ZN(n4954) );
  NOR2_X1 U6332 ( .A1(n6459), .A2(n8418), .ZN(n4956) );
  OR2_X1 U6333 ( .A1(n9317), .A2(n10056), .ZN(n4957) );
  OR2_X1 U6334 ( .A1(n6072), .A2(n6522), .ZN(n4958) );
  NOR2_X1 U6335 ( .A1(n8547), .A2(n8635), .ZN(n4959) );
  OR2_X1 U6336 ( .A1(n8814), .A2(n9122), .ZN(n4960) );
  OR2_X1 U6337 ( .A1(n8814), .A2(n9037), .ZN(n4961) );
  AND2_X1 U6338 ( .A1(n4961), .A2(n6506), .ZN(n4962) );
  AND2_X1 U6339 ( .A1(n4329), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n4963) );
  NAND2_X1 U6340 ( .A1(n6264), .A2(n6263), .ZN(n8976) );
  INV_X1 U6341 ( .A(n7365), .ZN(n5540) );
  INV_X1 U6342 ( .A(n9886), .ZN(n10068) );
  INV_X1 U6343 ( .A(n9321), .ZN(n7304) );
  OR2_X1 U6344 ( .A1(n9438), .A2(n9437), .ZN(n4967) );
  INV_X1 U6345 ( .A(n7697), .ZN(n7784) );
  NAND2_X1 U6346 ( .A1(n9070), .A2(n8845), .ZN(n4969) );
  AND2_X1 U6347 ( .A1(n8264), .A2(n8265), .ZN(n4970) );
  NAND2_X1 U6348 ( .A1(n6274), .A2(n6273), .ZN(n8244) );
  INV_X1 U6349 ( .A(n10243), .ZN(n6505) );
  INV_X1 U6350 ( .A(n8330), .ZN(n8331) );
  OAI211_X1 U6351 ( .C1(n5929), .C2(n5928), .A(n8297), .B(n5927), .ZN(n5931)
         );
  INV_X1 U6352 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5401) );
  INV_X1 U6353 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5124) );
  INV_X1 U6354 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5399) );
  NAND2_X1 U6355 ( .A1(n7364), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5485) );
  INV_X1 U6356 ( .A(n10131), .ZN(n6129) );
  INV_X1 U6357 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5400) );
  INV_X1 U6358 ( .A(n6620), .ZN(n6621) );
  AND4_X1 U6359 ( .A1(n5135), .A2(n7040), .A3(n5351), .A4(n5375), .ZN(n5136)
         );
  NAND2_X1 U6360 ( .A1(n4359), .A2(n8462), .ZN(n8463) );
  INV_X1 U6361 ( .A(n6165), .ZN(n5478) );
  INV_X1 U6362 ( .A(n8885), .ZN(n8496) );
  NOR2_X1 U6363 ( .A1(P2_IR_REG_26__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5419) );
  INV_X1 U6364 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5375) );
  NOR2_X1 U6365 ( .A1(n4947), .A2(n6621), .ZN(n6622) );
  NAND2_X1 U6366 ( .A1(n5973), .A2(n6758), .ZN(n5974) );
  INV_X1 U6367 ( .A(n5844), .ZN(n5627) );
  OR2_X1 U6368 ( .A1(n9708), .A2(n9305), .ZN(n8281) );
  OR2_X1 U6369 ( .A1(n8274), .A2(n9308), .ZN(n8275) );
  INV_X1 U6370 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5137) );
  INV_X1 U6371 ( .A(n5289), .ZN(n5040) );
  INV_X1 U6372 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5293) );
  INV_X1 U6373 ( .A(n5224), .ZN(n5003) );
  AND2_X1 U6374 ( .A1(n7204), .A2(n7203), .ZN(n8672) );
  INV_X1 U6375 ( .A(n6093), .ZN(n6094) );
  AOI21_X1 U6376 ( .B1(n7397), .B2(n7395), .A(n7396), .ZN(n7399) );
  INV_X1 U6377 ( .A(n7361), .ZN(n5484) );
  INV_X1 U6378 ( .A(n6663), .ZN(n6664) );
  OR2_X1 U6379 ( .A1(n5888), .A2(n9221), .ZN(n5890) );
  NAND2_X1 U6380 ( .A1(n5628), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n5852) );
  NOR2_X1 U6381 ( .A1(n9749), .A2(n9252), .ZN(n8292) );
  OR2_X1 U6382 ( .A1(n5846), .A2(n9178), .ZN(n5658) );
  OR2_X1 U6383 ( .A1(n5809), .A2(n5800), .ZN(n5834) );
  INV_X1 U6384 ( .A(n9728), .ZN(n8192) );
  NOR2_X1 U6385 ( .A1(n5736), .A2(n5735), .ZN(n5747) );
  NAND2_X1 U6386 ( .A1(n7593), .A2(n7499), .ZN(n7500) );
  NAND2_X1 U6387 ( .A1(n7431), .A2(n7458), .ZN(n7459) );
  NAND2_X1 U6388 ( .A1(n5356), .A2(n5357), .ZN(n9787) );
  XNOR2_X1 U6389 ( .A(n5024), .B(SI_10_), .ZN(n5252) );
  NAND2_X1 U6390 ( .A1(n5001), .A2(SI_6_), .ZN(n5002) );
  AND2_X1 U6391 ( .A1(n8506), .A2(n8505), .ZN(n8507) );
  NOR2_X1 U6392 ( .A1(n8710), .A2(n8711), .ZN(n8709) );
  INV_X1 U6393 ( .A(n8926), .ZN(n8959) );
  INV_X1 U6394 ( .A(n8377), .ZN(n6456) );
  INV_X1 U6395 ( .A(n8845), .ZN(n8826) );
  INV_X1 U6396 ( .A(n8977), .ZN(n8182) );
  INV_X1 U6397 ( .A(n10132), .ZN(n10157) );
  NAND2_X1 U6398 ( .A1(n6665), .A2(n6664), .ZN(n8113) );
  NAND2_X1 U6399 ( .A1(n5629), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5875) );
  AND2_X1 U6400 ( .A1(n6750), .A2(n6749), .ZN(n6751) );
  NAND2_X1 U6401 ( .A1(n6078), .A2(n6077), .ZN(n6079) );
  INV_X1 U6402 ( .A(n5898), .ZN(n5919) );
  OR2_X1 U6403 ( .A1(n5852), .A2(n9212), .ZN(n5854) );
  NAND2_X1 U6404 ( .A1(n5978), .A2(n8313), .ZN(n9470) );
  NAND2_X1 U6405 ( .A1(n8311), .A2(n5986), .ZN(n9507) );
  AOI22_X1 U6406 ( .A1(n9608), .A2(n8280), .B1(n9772), .B2(n8279), .ZN(n9590)
         );
  AND2_X1 U6407 ( .A1(n8163), .A2(n9310), .ZN(n8126) );
  NAND2_X1 U6408 ( .A1(n7259), .A2(n7257), .ZN(n7303) );
  INV_X1 U6409 ( .A(n9275), .ZN(n9287) );
  AND2_X1 U6410 ( .A1(n6971), .A2(n6970), .ZN(n9596) );
  XNOR2_X1 U6411 ( .A(n5035), .B(SI_14_), .ZN(n5274) );
  AND2_X1 U6412 ( .A1(n5016), .A2(n5015), .ZN(n5238) );
  XNOR2_X1 U6413 ( .A(n5004), .B(SI_7_), .ZN(n5224) );
  INV_X1 U6414 ( .A(n8688), .ZN(n8664) );
  AND2_X1 U6415 ( .A1(n6403), .A2(n6402), .ZN(n8855) );
  AND3_X1 U6416 ( .A1(n6329), .A2(n6328), .A3(n6327), .ZN(n8943) );
  AND4_X1 U6417 ( .A1(n6237), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(n8174)
         );
  INV_X4 U6418 ( .A(n6265), .ZN(n8450) );
  AND2_X1 U6419 ( .A1(n7203), .A2(n8458), .ZN(n10130) );
  INV_X1 U6420 ( .A(n8949), .ZN(n10138) );
  INV_X1 U6421 ( .A(n8493), .ZN(n8242) );
  INV_X1 U6422 ( .A(n10210), .ZN(n10221) );
  AND2_X1 U6423 ( .A1(n6486), .A2(n6896), .ZN(n6995) );
  AND2_X1 U6424 ( .A1(n5757), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5764) );
  OR2_X1 U6425 ( .A1(n10069), .A2(n6761), .ZN(n10021) );
  NAND2_X1 U6426 ( .A1(n5764), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5785) );
  OAI21_X1 U6427 ( .B1(n9745), .B2(n9280), .A(n6779), .ZN(n6780) );
  AND2_X1 U6428 ( .A1(n5644), .A2(n5643), .ZN(n9276) );
  AND4_X1 U6429 ( .A1(n5805), .A2(n5804), .A3(n5803), .A4(n5802), .ZN(n9240)
         );
  NAND2_X1 U6430 ( .A1(n5664), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5667) );
  AND2_X1 U6431 ( .A1(n8309), .A2(n5871), .ZN(n9540) );
  INV_X1 U6432 ( .A(n10038), .ZN(n10015) );
  INV_X1 U6433 ( .A(n9780), .ZN(n5396) );
  AOI211_X1 U6434 ( .C1(n9662), .C2(n9723), .A(n9661), .B(n9660), .ZN(n9738)
         );
  INV_X1 U6435 ( .A(n10062), .ZN(n9723) );
  INV_X1 U6436 ( .A(n5356), .ZN(n5139) );
  AND2_X1 U6437 ( .A1(n5258), .A2(n5249), .ZN(n9853) );
  XNOR2_X1 U6438 ( .A(n5000), .B(SI_6_), .ZN(n5216) );
  AND2_X1 U6439 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10247), .ZN(n10244) );
  AND2_X1 U6440 ( .A1(n7007), .A2(n7006), .ZN(n8688) );
  AND2_X1 U6441 ( .A1(n8455), .A2(n6432), .ZN(n8825) );
  INV_X1 U6442 ( .A(n8855), .ZN(n8698) );
  INV_X1 U6443 ( .A(n10090), .ZN(n10128) );
  AND2_X1 U6444 ( .A1(n7319), .A2(n10149), .ZN(n10162) );
  XNOR2_X1 U6445 ( .A(n8831), .B(n8830), .ZN(n9073) );
  AND2_X1 U6446 ( .A1(n6516), .A2(n6515), .ZN(n10224) );
  INV_X1 U6447 ( .A(n6194), .ZN(n7750) );
  AND2_X1 U6448 ( .A1(n6762), .A2(n10021), .ZN(n9280) );
  AND2_X1 U6449 ( .A1(n6775), .A2(n6774), .ZN(n9890) );
  OR2_X1 U6450 ( .A1(n6086), .A2(n6085), .ZN(n6087) );
  OR2_X1 U6451 ( .A1(n5661), .A2(n5660), .ZN(n9304) );
  OR2_X1 U6452 ( .A1(n10045), .A2(n7571), .ZN(n9629) );
  INV_X1 U6453 ( .A(n10023), .ZN(n10033) );
  OR2_X1 U6454 ( .A1(n7266), .A2(n7558), .ZN(n10080) );
  INV_X1 U6455 ( .A(n9587), .ZN(n9767) );
  OR2_X1 U6456 ( .A1(n7266), .A2(n6756), .ZN(n10075) );
  INV_X1 U6457 ( .A(n10047), .ZN(n10048) );
  INV_X1 U6458 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7152) );
  INV_X1 U6459 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n10248) );
  AND2_X1 U6460 ( .A1(n6785), .A2(n6784), .ZN(P1_U3973) );
  NAND2_X1 U6461 ( .A1(n6088), .A2(n6087), .ZN(P1_U3242) );
  INV_X1 U6462 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5395) );
  AND2_X1 U6463 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4975) );
  NAND2_X1 U6464 ( .A1(n6100), .A2(n4975), .ZN(n6118) );
  AND2_X1 U6465 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4976) );
  NAND2_X1 U6466 ( .A1(n4992), .A2(n4976), .ZN(n5180) );
  NAND2_X1 U6467 ( .A1(n6118), .A2(n5180), .ZN(n5168) );
  INV_X1 U6468 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6848) );
  INV_X1 U6469 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n4977) );
  NAND2_X1 U6470 ( .A1(n5168), .A2(n5169), .ZN(n4982) );
  INV_X1 U6471 ( .A(n4979), .ZN(n4980) );
  NAND2_X1 U6472 ( .A1(n4980), .A2(SI_1_), .ZN(n4981) );
  INV_X1 U6473 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6858) );
  INV_X1 U6474 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n4983) );
  MUX2_X1 U6475 ( .A(n6858), .B(n4983), .S(n4992), .Z(n4984) );
  XNOR2_X1 U6476 ( .A(n4984), .B(SI_2_), .ZN(n5183) );
  NAND2_X1 U6477 ( .A1(n5184), .A2(n5183), .ZN(n4987) );
  INV_X1 U6478 ( .A(n4984), .ZN(n4985) );
  NAND2_X1 U6479 ( .A1(n4985), .A2(SI_2_), .ZN(n4986) );
  INV_X1 U6480 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6860) );
  INV_X1 U6481 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4988) );
  MUX2_X1 U6482 ( .A(n6860), .B(n4988), .S(n4992), .Z(n4989) );
  XNOR2_X1 U6483 ( .A(n4989), .B(SI_3_), .ZN(n5191) );
  INV_X1 U6484 ( .A(n4989), .ZN(n4990) );
  NAND2_X1 U6485 ( .A1(n4990), .A2(SI_3_), .ZN(n4991) );
  MUX2_X1 U6486 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n4992), .Z(n4993) );
  INV_X1 U6487 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6856) );
  INV_X1 U6488 ( .A(n4995), .ZN(n4996) );
  NAND2_X1 U6489 ( .A1(n4996), .A2(SI_5_), .ZN(n4997) );
  INV_X1 U6490 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6863) );
  INV_X1 U6491 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n4999) );
  MUX2_X1 U6492 ( .A(n6863), .B(n4999), .S(n6846), .Z(n5000) );
  INV_X1 U6493 ( .A(n5000), .ZN(n5001) );
  MUX2_X1 U6494 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6846), .Z(n5004) );
  NAND2_X1 U6495 ( .A1(n5004), .A2(SI_7_), .ZN(n5005) );
  INV_X1 U6496 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6869) );
  MUX2_X1 U6497 ( .A(n6869), .B(n7166), .S(n6846), .Z(n5007) );
  INV_X1 U6498 ( .A(SI_8_), .ZN(n5006) );
  INV_X1 U6499 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6500 ( .A1(n5008), .A2(SI_8_), .ZN(n5009) );
  INV_X1 U6501 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5011) );
  MUX2_X1 U6502 ( .A(n5011), .B(n7152), .S(n6846), .Z(n5013) );
  INV_X1 U6503 ( .A(SI_9_), .ZN(n5012) );
  INV_X1 U6504 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6505 ( .A1(n5014), .A2(SI_9_), .ZN(n5015) );
  MUX2_X1 U6506 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6846), .Z(n5024) );
  INV_X1 U6507 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6902) );
  INV_X1 U6508 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n5018) );
  INV_X1 U6509 ( .A(SI_11_), .ZN(n5019) );
  INV_X1 U6510 ( .A(n5020), .ZN(n5021) );
  NAND2_X1 U6511 ( .A1(n5021), .A2(SI_11_), .ZN(n5022) );
  NAND2_X1 U6512 ( .A1(n5023), .A2(n5022), .ZN(n5256) );
  INV_X1 U6513 ( .A(n5256), .ZN(n5025) );
  NAND2_X1 U6514 ( .A1(n5024), .A2(SI_10_), .ZN(n5254) );
  INV_X1 U6515 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6893) );
  INV_X1 U6516 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5028) );
  MUX2_X1 U6517 ( .A(n6893), .B(n5028), .S(n6846), .Z(n5029) );
  INV_X1 U6518 ( .A(n5029), .ZN(n5030) );
  MUX2_X1 U6519 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6846), .Z(n5032) );
  NAND2_X1 U6520 ( .A1(n5032), .A2(SI_13_), .ZN(n5033) );
  MUX2_X1 U6521 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n6846), .Z(n5035) );
  MUX2_X1 U6522 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6846), .Z(n5282) );
  INV_X1 U6523 ( .A(n5282), .ZN(n5037) );
  INV_X1 U6524 ( .A(SI_15_), .ZN(n5036) );
  NAND2_X1 U6525 ( .A1(n5037), .A2(n5036), .ZN(n5038) );
  INV_X1 U6526 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5039) );
  INV_X1 U6527 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7202) );
  MUX2_X1 U6528 ( .A(n5039), .B(n7202), .S(n6846), .Z(n5289) );
  NAND2_X1 U6529 ( .A1(n5040), .A2(SI_16_), .ZN(n5041) );
  INV_X1 U6530 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n5043) );
  INV_X1 U6531 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5042) );
  MUX2_X1 U6532 ( .A(n5043), .B(n5042), .S(n6846), .Z(n5045) );
  INV_X1 U6533 ( .A(SI_17_), .ZN(n5044) );
  NAND2_X1 U6534 ( .A1(n5045), .A2(n5044), .ZN(n5048) );
  INV_X1 U6535 ( .A(n5045), .ZN(n5046) );
  NAND2_X1 U6536 ( .A1(n5046), .A2(SI_17_), .ZN(n5047) );
  NAND2_X1 U6537 ( .A1(n5048), .A2(n5047), .ZN(n5301) );
  INV_X1 U6538 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n5050) );
  INV_X1 U6539 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n5049) );
  MUX2_X1 U6540 ( .A(n5050), .B(n5049), .S(n6846), .Z(n5051) );
  XNOR2_X1 U6541 ( .A(n5051), .B(SI_18_), .ZN(n5306) );
  INV_X1 U6542 ( .A(n5051), .ZN(n5052) );
  INV_X1 U6543 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n5053) );
  INV_X1 U6544 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7620) );
  MUX2_X1 U6545 ( .A(n5053), .B(n7620), .S(n6846), .Z(n5055) );
  INV_X1 U6546 ( .A(SI_19_), .ZN(n5054) );
  NAND2_X1 U6547 ( .A1(n5055), .A2(n5054), .ZN(n5058) );
  INV_X1 U6548 ( .A(n5055), .ZN(n5056) );
  NAND2_X1 U6549 ( .A1(n5056), .A2(SI_19_), .ZN(n5057) );
  NAND2_X1 U6550 ( .A1(n5058), .A2(n5057), .ZN(n5315) );
  INV_X1 U6551 ( .A(SI_20_), .ZN(n5321) );
  MUX2_X1 U6552 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n6846), .Z(n5322) );
  INV_X1 U6553 ( .A(n5322), .ZN(n5059) );
  NAND2_X1 U6554 ( .A1(n5324), .A2(n5321), .ZN(n5060) );
  INV_X1 U6555 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n5062) );
  INV_X1 U6556 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7724) );
  MUX2_X1 U6557 ( .A(n5062), .B(n7724), .S(n6846), .Z(n5327) );
  INV_X1 U6558 ( .A(n5327), .ZN(n5063) );
  NAND2_X1 U6559 ( .A1(n5063), .A2(SI_21_), .ZN(n5064) );
  INV_X1 U6560 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5065) );
  INV_X1 U6561 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7889) );
  MUX2_X1 U6562 ( .A(n5065), .B(n7889), .S(n6846), .Z(n5067) );
  INV_X1 U6563 ( .A(SI_22_), .ZN(n5066) );
  NAND2_X1 U6564 ( .A1(n5067), .A2(n5066), .ZN(n5070) );
  INV_X1 U6565 ( .A(n5067), .ZN(n5068) );
  NAND2_X1 U6566 ( .A1(n5068), .A2(SI_22_), .ZN(n5069) );
  NAND2_X1 U6567 ( .A1(n5070), .A2(n5069), .ZN(n5164) );
  INV_X1 U6568 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5072) );
  INV_X1 U6569 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5071) );
  MUX2_X1 U6570 ( .A(n5072), .B(n5071), .S(n6846), .Z(n5074) );
  INV_X1 U6571 ( .A(SI_23_), .ZN(n5073) );
  NAND2_X1 U6572 ( .A1(n5074), .A2(n5073), .ZN(n5077) );
  INV_X1 U6573 ( .A(n5074), .ZN(n5075) );
  NAND2_X1 U6574 ( .A1(n5075), .A2(SI_23_), .ZN(n5076) );
  NAND2_X1 U6575 ( .A1(n5078), .A2(n5077), .ZN(n5333) );
  INV_X1 U6576 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5079) );
  INV_X1 U6577 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7996) );
  MUX2_X1 U6578 ( .A(n5079), .B(n7996), .S(n6846), .Z(n5080) );
  INV_X1 U6579 ( .A(SI_24_), .ZN(n7086) );
  NAND2_X1 U6580 ( .A1(n5080), .A2(n7086), .ZN(n5083) );
  INV_X1 U6581 ( .A(n5080), .ZN(n5081) );
  NAND2_X1 U6582 ( .A1(n5081), .A2(SI_24_), .ZN(n5082) );
  AND2_X1 U6583 ( .A1(n5083), .A2(n5082), .ZN(n5332) );
  INV_X1 U6584 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5084) );
  INV_X1 U6585 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8049) );
  MUX2_X1 U6586 ( .A(n5084), .B(n8049), .S(n6846), .Z(n5086) );
  INV_X1 U6587 ( .A(SI_25_), .ZN(n5085) );
  NAND2_X1 U6588 ( .A1(n5086), .A2(n5085), .ZN(n5089) );
  INV_X1 U6589 ( .A(n5086), .ZN(n5087) );
  NAND2_X1 U6590 ( .A1(n5087), .A2(SI_25_), .ZN(n5088) );
  AND2_X1 U6591 ( .A1(n5089), .A2(n5088), .ZN(n5156) );
  INV_X1 U6592 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5090) );
  INV_X1 U6593 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8142) );
  MUX2_X1 U6594 ( .A(n5090), .B(n8142), .S(n6846), .Z(n5092) );
  INV_X1 U6595 ( .A(SI_26_), .ZN(n5091) );
  NAND2_X1 U6596 ( .A1(n5092), .A2(n5091), .ZN(n5095) );
  INV_X1 U6597 ( .A(n5092), .ZN(n5093) );
  NAND2_X1 U6598 ( .A1(n5093), .A2(SI_26_), .ZN(n5094) );
  AND2_X1 U6599 ( .A1(n5095), .A2(n5094), .ZN(n5153) );
  NAND2_X1 U6600 ( .A1(n5152), .A2(n5153), .ZN(n5096) );
  INV_X1 U6601 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5097) );
  INV_X1 U6602 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8189) );
  MUX2_X1 U6603 ( .A(n5097), .B(n8189), .S(n6846), .Z(n5099) );
  INV_X1 U6604 ( .A(SI_27_), .ZN(n5098) );
  NAND2_X1 U6605 ( .A1(n5099), .A2(n5098), .ZN(n5102) );
  INV_X1 U6606 ( .A(n5099), .ZN(n5100) );
  NAND2_X1 U6607 ( .A1(n5100), .A2(SI_27_), .ZN(n5101) );
  AND2_X1 U6608 ( .A1(n5102), .A2(n5101), .ZN(n5336) );
  INV_X1 U6609 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5103) );
  INV_X1 U6610 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n8215) );
  MUX2_X1 U6611 ( .A(n5103), .B(n8215), .S(n6846), .Z(n5105) );
  XNOR2_X1 U6612 ( .A(n5105), .B(SI_28_), .ZN(n5341) );
  INV_X1 U6613 ( .A(SI_28_), .ZN(n5104) );
  NAND2_X1 U6614 ( .A1(n5105), .A2(n5104), .ZN(n5106) );
  INV_X1 U6615 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n5108) );
  INV_X1 U6616 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8566) );
  MUX2_X1 U6617 ( .A(n5108), .B(n8566), .S(n6846), .Z(n5110) );
  INV_X1 U6618 ( .A(SI_29_), .ZN(n5109) );
  INV_X1 U6619 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n5114) );
  INV_X1 U6620 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8222) );
  MUX2_X1 U6621 ( .A(n5114), .B(n8222), .S(n6846), .Z(n5115) );
  INV_X1 U6622 ( .A(SI_30_), .ZN(n7053) );
  NAND2_X1 U6623 ( .A1(n5115), .A2(n7053), .ZN(n5118) );
  INV_X1 U6624 ( .A(n5115), .ZN(n5116) );
  NAND2_X1 U6625 ( .A1(n5116), .A2(SI_30_), .ZN(n5117) );
  NAND2_X1 U6626 ( .A1(n5118), .A2(n5117), .ZN(n5145) );
  INV_X1 U6627 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5120) );
  INV_X1 U6628 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5119) );
  MUX2_X1 U6629 ( .A(n5120), .B(n5119), .S(n6846), .Z(n5121) );
  XNOR2_X1 U6630 ( .A(n5121), .B(SI_31_), .ZN(n5122) );
  NOR2_X1 U6631 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5134) );
  NOR2_X1 U6632 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5133) );
  NOR2_X1 U6633 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5132) );
  NOR2_X1 U6634 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5131) );
  INV_X1 U6635 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5135) );
  NAND2_X2 U6636 ( .A1(n8217), .A2(n8191), .ZN(n6812) );
  AND2_X2 U6637 ( .A1(n6812), .A2(n6846), .ZN(n5186) );
  NAND2_X1 U6638 ( .A1(n9151), .A2(n5342), .ZN(n5144) );
  NAND2_X1 U6639 ( .A1(n5343), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n5143) );
  INV_X4 U6640 ( .A(n5218), .ZN(n5342) );
  NAND2_X1 U6641 ( .A1(n8442), .A2(n5342), .ZN(n5148) );
  NAND2_X1 U6642 ( .A1(n5343), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5147) );
  NAND2_X1 U6643 ( .A1(n8218), .A2(n5342), .ZN(n5151) );
  NAND2_X1 U6644 ( .A1(n5343), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5150) );
  XNOR2_X1 U6645 ( .A(n5152), .B(n5153), .ZN(n8064) );
  NAND2_X1 U6646 ( .A1(n8064), .A2(n5342), .ZN(n5155) );
  NAND2_X1 U6647 ( .A1(n5343), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5154) );
  XNOR2_X1 U6648 ( .A(n5157), .B(n5156), .ZN(n7999) );
  NAND2_X1 U6649 ( .A1(n5343), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5158) );
  NAND2_X1 U6650 ( .A1(n7956), .A2(n5342), .ZN(n5163) );
  NAND2_X1 U6651 ( .A1(n5343), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5162) );
  XNOR2_X1 U6652 ( .A(n5165), .B(n5164), .ZN(n7809) );
  NAND2_X1 U6653 ( .A1(n7809), .A2(n5342), .ZN(n5167) );
  NAND2_X1 U6654 ( .A1(n5343), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U6655 ( .A1(n5182), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5177) );
  XNOR2_X1 U6656 ( .A(n5169), .B(n5168), .ZN(n6847) );
  INV_X1 U6657 ( .A(n6847), .ZN(n5170) );
  NAND2_X1 U6658 ( .A1(n5186), .A2(n5170), .ZN(n5176) );
  NAND2_X1 U6659 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5171) );
  MUX2_X1 U6660 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5171), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5172) );
  INV_X1 U6661 ( .A(n5172), .ZN(n5174) );
  NAND2_X1 U6662 ( .A1(n5204), .A2(n4336), .ZN(n5175) );
  NAND2_X1 U6663 ( .A1(n6846), .A2(SI_0_), .ZN(n5179) );
  INV_X1 U6664 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5178) );
  NAND2_X1 U6665 ( .A1(n5179), .A2(n5178), .ZN(n5181) );
  AND2_X1 U6666 ( .A1(n5181), .A2(n5180), .ZN(n9794) );
  MUX2_X1 U6667 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9794), .S(n6812), .Z(n7572) );
  NAND2_X1 U6668 ( .A1(n5182), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5190) );
  XNOR2_X1 U6669 ( .A(n5184), .B(n5183), .ZN(n6857) );
  INV_X1 U6670 ( .A(n6857), .ZN(n5185) );
  NAND2_X1 U6671 ( .A1(n5186), .A2(n5185), .ZN(n5189) );
  NAND2_X1 U6672 ( .A1(n5204), .A2(n9341), .ZN(n5188) );
  XNOR2_X1 U6673 ( .A(n5192), .B(n5191), .ZN(n6859) );
  INV_X1 U6674 ( .A(n6859), .ZN(n5193) );
  NAND2_X1 U6675 ( .A1(n5186), .A2(n5193), .ZN(n5200) );
  NAND2_X1 U6676 ( .A1(n5182), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5199) );
  NAND2_X1 U6677 ( .A1(n5194), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5195) );
  MUX2_X1 U6678 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5195), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n5197) );
  AND2_X1 U6679 ( .A1(n5197), .A2(n5196), .ZN(n9354) );
  NAND2_X1 U6680 ( .A1(n5204), .A2(n9354), .ZN(n5198) );
  NAND2_X1 U6681 ( .A1(n7648), .A2(n7431), .ZN(n7463) );
  XNOR2_X1 U6682 ( .A(n5202), .B(n5201), .ZN(n6853) );
  INV_X1 U6683 ( .A(n6853), .ZN(n5203) );
  NAND2_X1 U6684 ( .A1(n5342), .A2(n5203), .ZN(n5208) );
  NAND2_X1 U6685 ( .A1(n5182), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5207) );
  NAND2_X1 U6686 ( .A1(n5196), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5205) );
  XNOR2_X1 U6687 ( .A(n5205), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U6688 ( .A1(n5204), .A2(n6911), .ZN(n5206) );
  XNOR2_X1 U6689 ( .A(n5210), .B(n5209), .ZN(n6855) );
  INV_X1 U6690 ( .A(n6855), .ZN(n5211) );
  NAND2_X1 U6691 ( .A1(n5342), .A2(n5211), .ZN(n5215) );
  NAND2_X1 U6692 ( .A1(n5182), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5214) );
  NOR2_X1 U6693 ( .A1(n5196), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5220) );
  OR2_X1 U6694 ( .A1(n5220), .A2(n9788), .ZN(n5212) );
  XNOR2_X1 U6695 ( .A(n5212), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6949) );
  NAND2_X1 U6696 ( .A1(n5204), .A2(n6949), .ZN(n5213) );
  XNOR2_X1 U6697 ( .A(n5217), .B(n5216), .ZN(n6862) );
  OR2_X1 U6698 ( .A1(n5218), .A2(n6862), .ZN(n5223) );
  INV_X1 U6699 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5219) );
  NAND2_X1 U6700 ( .A1(n5220), .A2(n5219), .ZN(n5234) );
  NAND2_X1 U6701 ( .A1(n5234), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5227) );
  XNOR2_X1 U6702 ( .A(n5227), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6924) );
  NAND2_X1 U6703 ( .A1(n5204), .A2(n6924), .ZN(n5222) );
  NAND2_X1 U6704 ( .A1(n5182), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5221) );
  XNOR2_X1 U6705 ( .A(n5225), .B(n5224), .ZN(n6864) );
  NAND2_X1 U6706 ( .A1(n6864), .A2(n5342), .ZN(n5231) );
  INV_X1 U6707 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U6708 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  NAND2_X1 U6709 ( .A1(n5228), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5229) );
  XNOR2_X1 U6710 ( .A(n5229), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6937) );
  AOI22_X1 U6711 ( .A1(n5343), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5204), .B2(
        n6937), .ZN(n5230) );
  XNOR2_X1 U6712 ( .A(n5233), .B(n5232), .ZN(n6868) );
  NAND2_X1 U6713 ( .A1(n6868), .A2(n5342), .ZN(n5237) );
  NAND2_X1 U6714 ( .A1(n5240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5235) );
  XNOR2_X1 U6715 ( .A(n5235), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9370) );
  AOI22_X1 U6716 ( .A1(n5343), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5204), .B2(
        n9370), .ZN(n5236) );
  XNOR2_X1 U6717 ( .A(n5239), .B(n5238), .ZN(n6872) );
  NAND2_X1 U6718 ( .A1(n6872), .A2(n5342), .ZN(n5243) );
  NOR2_X1 U6719 ( .A1(n5240), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n5245) );
  OR2_X1 U6720 ( .A1(n5245), .A2(n9788), .ZN(n5241) );
  XNOR2_X1 U6721 ( .A(n5241), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9400) );
  AOI22_X1 U6722 ( .A1(n5343), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5204), .B2(
        n9400), .ZN(n5242) );
  INV_X1 U6723 ( .A(n5252), .ZN(n5244) );
  INV_X1 U6724 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U6725 ( .A1(n5245), .A2(n7020), .ZN(n5246) );
  NAND2_X1 U6726 ( .A1(n5246), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5248) );
  INV_X1 U6727 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5247) );
  NAND2_X1 U6728 ( .A1(n5248), .A2(n5247), .ZN(n5258) );
  OR2_X1 U6729 ( .A1(n5248), .A2(n5247), .ZN(n5249) );
  AOI22_X1 U6730 ( .A1(n5343), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5204), .B2(
        n9853), .ZN(n5250) );
  NAND2_X1 U6731 ( .A1(n5255), .A2(n5254), .ZN(n5257) );
  XNOR2_X1 U6732 ( .A(n5256), .B(n5257), .ZN(n6887) );
  NAND2_X1 U6733 ( .A1(n6887), .A2(n5342), .ZN(n5261) );
  NAND2_X1 U6734 ( .A1(n5258), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5259) );
  XNOR2_X1 U6735 ( .A(n5259), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9899) );
  AOI22_X1 U6736 ( .A1(n5343), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5204), .B2(
        n9899), .ZN(n5260) );
  XNOR2_X1 U6737 ( .A(n5263), .B(n5262), .ZN(n6889) );
  NAND2_X1 U6738 ( .A1(n6889), .A2(n5342), .ZN(n5266) );
  INV_X1 U6739 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9788) );
  OR2_X1 U6740 ( .A1(n5270), .A2(n9788), .ZN(n5264) );
  XNOR2_X1 U6741 ( .A(n5264), .B(P1_IR_REG_12__SCAN_IN), .ZN(n9903) );
  AOI22_X1 U6742 ( .A1(n5343), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5204), .B2(
        n9903), .ZN(n5265) );
  XNOR2_X1 U6743 ( .A(n5268), .B(n5267), .ZN(n6954) );
  NAND2_X1 U6744 ( .A1(n6954), .A2(n5342), .ZN(n5273) );
  INV_X1 U6745 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5269) );
  OR2_X1 U6746 ( .A1(n5277), .A2(n9788), .ZN(n5271) );
  XNOR2_X1 U6747 ( .A(n5271), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9919) );
  AOI22_X1 U6748 ( .A1(n5343), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5204), .B2(
        n9919), .ZN(n5272) );
  XNOR2_X1 U6749 ( .A(n5275), .B(n5274), .ZN(n6962) );
  NAND2_X1 U6750 ( .A1(n6962), .A2(n5342), .ZN(n5281) );
  INV_X1 U6751 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5276) );
  NAND2_X1 U6752 ( .A1(n5277), .A2(n5276), .ZN(n5294) );
  NAND2_X1 U6753 ( .A1(n5294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6754 ( .A1(n5278), .A2(n5292), .ZN(n5285) );
  OR2_X1 U6755 ( .A1(n5278), .A2(n5292), .ZN(n5279) );
  AND2_X1 U6756 ( .A1(n5285), .A2(n5279), .ZN(n9407) );
  AOI22_X1 U6757 ( .A1(n5343), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5204), .B2(
        n9407), .ZN(n5280) );
  XNOR2_X1 U6758 ( .A(n5282), .B(SI_15_), .ZN(n5283) );
  XNOR2_X1 U6759 ( .A(n5284), .B(n5283), .ZN(n6976) );
  NAND2_X1 U6760 ( .A1(n6976), .A2(n5342), .ZN(n5288) );
  NAND2_X1 U6761 ( .A1(n5285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5286) );
  XNOR2_X1 U6762 ( .A(n5286), .B(n5293), .ZN(n9409) );
  INV_X1 U6763 ( .A(n9409), .ZN(n9960) );
  AOI22_X1 U6764 ( .A1(n5343), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5204), .B2(
        n9960), .ZN(n5287) );
  NAND2_X1 U6765 ( .A1(n8194), .A2(n9781), .ZN(n8195) );
  XNOR2_X1 U6766 ( .A(n5289), .B(SI_16_), .ZN(n5290) );
  NAND2_X1 U6767 ( .A1(n7197), .A2(n5342), .ZN(n5300) );
  NAND2_X1 U6768 ( .A1(n5295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5296) );
  MUX2_X1 U6769 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5296), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n5298) );
  INV_X1 U6770 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5297) );
  NAND2_X1 U6771 ( .A1(n5298), .A2(n5303), .ZN(n9973) );
  INV_X1 U6772 ( .A(n9973), .ZN(n9390) );
  AOI22_X1 U6773 ( .A1(n5343), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5204), .B2(
        n9390), .ZN(n5299) );
  XNOR2_X1 U6774 ( .A(n5302), .B(n5301), .ZN(n7326) );
  NAND2_X1 U6775 ( .A1(n7326), .A2(n5342), .ZN(n5305) );
  NAND2_X1 U6776 ( .A1(n5303), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5309) );
  XNOR2_X1 U6777 ( .A(n5309), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U6778 ( .A1(n5343), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5204), .B2(
        n9984), .ZN(n5304) );
  XNOR2_X1 U6779 ( .A(n5307), .B(n5306), .ZN(n7454) );
  NAND2_X1 U6780 ( .A1(n7454), .A2(n5342), .ZN(n5314) );
  INV_X1 U6781 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5308) );
  NAND2_X1 U6782 ( .A1(n5309), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U6783 ( .A1(n5310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5311) );
  INV_X1 U6784 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7177) );
  OR2_X1 U6785 ( .A1(n5311), .A2(n7177), .ZN(n5312) );
  AND2_X1 U6786 ( .A1(n5317), .A2(n5312), .ZN(n10004) );
  AOI22_X1 U6787 ( .A1(n5343), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5204), .B2(
        n10004), .ZN(n5313) );
  XNOR2_X1 U6788 ( .A(n5316), .B(n5315), .ZN(n7516) );
  NAND2_X1 U6789 ( .A1(n7516), .A2(n5342), .ZN(n5320) );
  INV_X1 U6790 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5318) );
  AOI22_X1 U6791 ( .A1(n5343), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7570), .B2(
        n5204), .ZN(n5319) );
  XNOR2_X1 U6792 ( .A(n5322), .B(n5321), .ZN(n5323) );
  XNOR2_X1 U6793 ( .A(n5324), .B(n5323), .ZN(n7600) );
  NAND2_X1 U6794 ( .A1(n7600), .A2(n5342), .ZN(n5326) );
  NAND2_X1 U6795 ( .A1(n5343), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5325) );
  XNOR2_X1 U6796 ( .A(n5327), .B(SI_21_), .ZN(n5328) );
  XNOR2_X1 U6797 ( .A(n5329), .B(n5328), .ZN(n7710) );
  NAND2_X1 U6798 ( .A1(n7710), .A2(n5342), .ZN(n5331) );
  NAND2_X1 U6799 ( .A1(n5182), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5330) );
  XNOR2_X1 U6800 ( .A(n5333), .B(n5332), .ZN(n7979) );
  NAND2_X1 U6801 ( .A1(n7979), .A2(n5342), .ZN(n5335) );
  NAND2_X1 U6802 ( .A1(n5343), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5334) );
  AND2_X2 U6803 ( .A1(n9745), .A2(n9492), .ZN(n9476) );
  NAND2_X1 U6804 ( .A1(n8145), .A2(n5342), .ZN(n5339) );
  NAND2_X1 U6805 ( .A1(n5182), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5338) );
  NAND2_X1 U6806 ( .A1(n5343), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5344) );
  XNOR2_X1 U6807 ( .A(n5940), .B(n9429), .ZN(n5353) );
  NAND2_X1 U6808 ( .A1(n5346), .A2(n5351), .ZN(n5348) );
  NAND2_X1 U6809 ( .A1(n5347), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5376) );
  INV_X1 U6810 ( .A(n6969), .ZN(n7891) );
  NAND2_X1 U6811 ( .A1(n5348), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U6812 ( .A(n5349), .B(P1_IR_REG_21__SCAN_IN), .ZN(n6083) );
  INV_X1 U6813 ( .A(n6083), .ZN(n7726) );
  AND2_X1 U6814 ( .A1(n7891), .A2(n7726), .ZN(n7563) );
  INV_X1 U6815 ( .A(n5346), .ZN(n5350) );
  NAND2_X1 U6816 ( .A1(n5350), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5352) );
  AND2_X1 U6817 ( .A1(n7563), .A2(n7624), .ZN(n10058) );
  INV_X1 U6818 ( .A(n10058), .ZN(n9627) );
  INV_X1 U6819 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5357) );
  INV_X1 U6820 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5354) );
  XNOR2_X2 U6821 ( .A(n5355), .B(n5354), .ZN(n5359) );
  XNOR2_X2 U6823 ( .A(n5358), .B(n5357), .ZN(n8567) );
  INV_X1 U6824 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6825 ( .A1(n4338), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n5362) );
  INV_X1 U6826 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5360) );
  OR2_X1 U6827 ( .A1(n4340), .A2(n5360), .ZN(n5361) );
  OAI211_X1 U6828 ( .C1(n4327), .C2(n5363), .A(n5362), .B(n5361), .ZN(n6891)
         );
  AND2_X1 U6829 ( .A1(n6969), .A2(n6083), .ZN(n6810) );
  NAND2_X1 U6830 ( .A1(n8217), .A2(n6810), .ZN(n9275) );
  INV_X1 U6831 ( .A(n8191), .ZN(n6084) );
  AND2_X1 U6832 ( .A1(n6084), .A2(P1_B_REG_SCAN_IN), .ZN(n5364) );
  NOR2_X1 U6833 ( .A1(n9275), .A2(n5364), .ZN(n8317) );
  AND2_X1 U6834 ( .A1(n6891), .A2(n8317), .ZN(n9647) );
  NOR2_X1 U6835 ( .A1(n9424), .A2(n9647), .ZN(n9644) );
  INV_X1 U6836 ( .A(n7624), .ZN(n6758) );
  NAND2_X1 U6837 ( .A1(n6521), .A2(n7624), .ZN(n6522) );
  NAND2_X1 U6838 ( .A1(n6522), .A2(n6810), .ZN(n6767) );
  NAND2_X1 U6839 ( .A1(n5371), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5366) );
  MUX2_X1 U6840 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5366), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5368) );
  NAND2_X1 U6841 ( .A1(n5368), .A2(n5367), .ZN(n8051) );
  NAND2_X1 U6842 ( .A1(n4581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5370) );
  MUX2_X1 U6843 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5370), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n5372) );
  NAND2_X1 U6844 ( .A1(n5372), .A2(n5371), .ZN(n7998) );
  NOR2_X1 U6845 ( .A1(n8051), .A2(n7998), .ZN(n5374) );
  NAND2_X1 U6846 ( .A1(n5367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5373) );
  XNOR2_X1 U6847 ( .A(n5373), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6848 ( .A1(n5374), .A2(n5381), .ZN(n6768) );
  NAND2_X1 U6849 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  NAND2_X1 U6850 ( .A1(n5377), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5378) );
  XNOR2_X1 U6851 ( .A(n5378), .B(n7040), .ZN(n6809) );
  AND2_X1 U6852 ( .A1(n6809), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6784) );
  AND2_X1 U6853 ( .A1(n6768), .A2(n6784), .ZN(n6813) );
  AND2_X1 U6854 ( .A1(n6767), .A2(n6813), .ZN(n7560) );
  NAND2_X1 U6855 ( .A1(n8051), .A2(P1_B_REG_SCAN_IN), .ZN(n5379) );
  MUX2_X1 U6856 ( .A(P1_B_REG_SCAN_IN), .B(n5379), .S(n7998), .Z(n5380) );
  INV_X1 U6857 ( .A(n5380), .ZN(n5382) );
  INV_X1 U6858 ( .A(n5381), .ZN(n8144) );
  NOR2_X1 U6859 ( .A1(n5382), .A2(n8144), .ZN(n9784) );
  NOR4_X1 U6860 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n5391) );
  NOR4_X1 U6861 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n5390) );
  OR4_X1 U6862 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .A3(
        P1_D_REG_3__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n5388) );
  NOR4_X1 U6863 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_19__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n5386) );
  NOR4_X1 U6864 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5385) );
  NOR4_X1 U6865 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5384) );
  NOR4_X1 U6866 ( .A1(P1_D_REG_21__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n5383) );
  NAND4_X1 U6867 ( .A1(n5386), .A2(n5385), .A3(n5384), .A4(n5383), .ZN(n5387)
         );
  NOR4_X1 U6868 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        n5388), .A4(n5387), .ZN(n5389) );
  NAND3_X1 U6869 ( .A1(n5391), .A2(n5390), .A3(n5389), .ZN(n5392) );
  NAND2_X1 U6870 ( .A1(n9784), .A2(n5392), .ZN(n6754) );
  INV_X1 U6871 ( .A(n9784), .ZN(n5394) );
  NAND2_X1 U6872 ( .A1(n8144), .A2(n8051), .ZN(n9785) );
  OAI21_X1 U6873 ( .B1(n5394), .B2(P1_D_REG_1__SCAN_IN), .A(n9785), .ZN(n6753)
         );
  AND2_X1 U6874 ( .A1(n6754), .A2(n6753), .ZN(n5393) );
  OAI211_X1 U6875 ( .C1(n10069), .C2(n6083), .A(n7560), .B(n5393), .ZN(n7266)
         );
  NAND2_X1 U6876 ( .A1(n8144), .A2(n7998), .ZN(n9786) );
  OAI21_X1 U6877 ( .B1(n5394), .B2(P1_D_REG_0__SCAN_IN), .A(n9786), .ZN(n7558)
         );
  INV_X1 U6878 ( .A(n7558), .ZN(n6756) );
  INV_X2 U6879 ( .A(n10075), .ZN(n10077) );
  MUX2_X1 U6880 ( .A(n5395), .B(n9644), .S(n10077), .Z(n5398) );
  AND2_X1 U6881 ( .A1(n6522), .A2(n7563), .ZN(n10057) );
  NAND2_X1 U6882 ( .A1(n10077), .A2(n10057), .ZN(n9780) );
  NAND2_X1 U6883 ( .A1(n5398), .A2(n5397), .ZN(P1_U3521) );
  NOR2_X4 U6884 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5466) );
  INV_X1 U6885 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5408) );
  INV_X1 U6886 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5404) );
  INV_X1 U6887 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n5403) );
  NOR2_X1 U6888 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5406) );
  NOR2_X1 U6889 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5405) );
  NOR2_X1 U6890 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5407) );
  INV_X1 U6891 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5410) );
  INV_X1 U6892 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5411) );
  NAND2_X1 U6893 ( .A1(n5434), .A2(n5411), .ZN(n5430) );
  INV_X1 U6894 ( .A(n5430), .ZN(n5412) );
  NAND2_X1 U6895 ( .A1(n5412), .A2(n5431), .ZN(n5423) );
  INV_X1 U6896 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5424) );
  INV_X1 U6897 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5413) );
  NAND2_X1 U6898 ( .A1(n5424), .A2(n5413), .ZN(n5414) );
  OAI21_X1 U6899 ( .B1(n5423), .B2(n5414), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5416) );
  NOR2_X1 U6900 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n5418) );
  NOR2_X1 U6901 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5417) );
  INV_X1 U6902 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6903 ( .A1(n5423), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5426) );
  NAND2_X1 U6904 ( .A1(n5426), .A2(n5424), .ZN(n5427) );
  NAND2_X1 U6905 ( .A1(n8065), .A2(n6479), .ZN(n6476) );
  INV_X1 U6906 ( .A(n6476), .ZN(n5429) );
  OR2_X1 U6907 ( .A1(n5426), .A2(n5424), .ZN(n5428) );
  NAND2_X1 U6908 ( .A1(n5428), .A2(n5427), .ZN(n6474) );
  INV_X1 U6909 ( .A(n6474), .ZN(n7980) );
  NAND2_X1 U6910 ( .A1(n5429), .A2(n7980), .ZN(n6486) );
  INV_X1 U6911 ( .A(n6486), .ZN(n5433) );
  NAND2_X1 U6912 ( .A1(n5430), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5432) );
  XNOR2_X1 U6913 ( .A(n5432), .B(n5431), .ZN(n6896) );
  NAND2_X1 U6914 ( .A1(n5433), .A2(n6896), .ZN(n5615) );
  INV_X1 U6915 ( .A(n5434), .ZN(n5437) );
  NAND2_X1 U6916 ( .A1(n5437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5435) );
  XNOR2_X1 U6917 ( .A(n5435), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8513) );
  NAND2_X1 U6918 ( .A1(n4374), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5436) );
  MUX2_X1 U6919 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5436), .S(
        P2_IR_REG_21__SCAN_IN), .Z(n5438) );
  NAND2_X1 U6920 ( .A1(n5438), .A2(n5437), .ZN(n7348) );
  NAND2_X2 U6921 ( .A1(n8513), .A2(n8326), .ZN(n8457) );
  NAND2_X1 U6922 ( .A1(n8458), .A2(n6896), .ZN(n5439) );
  NAND2_X1 U6923 ( .A1(n5615), .A2(n5439), .ZN(n5614) );
  INV_X1 U6924 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5440) );
  XNOR2_X2 U6925 ( .A(n5441), .B(n4703), .ZN(n8510) );
  NAND2_X4 U6926 ( .A1(n5445), .A2(n5444), .ZN(n5612) );
  OR2_X1 U6927 ( .A1(n5614), .A2(n6318), .ZN(n5446) );
  NAND2_X1 U6928 ( .A1(n5446), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X2 U6929 ( .A1(n5461), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5459) );
  INV_X1 U6930 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5447) );
  INV_X1 U6931 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U6932 ( .A1(n5505), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5449) );
  NAND2_X1 U6933 ( .A1(n5453), .A2(n5449), .ZN(n5493) );
  OAI21_X1 U6934 ( .B1(n5493), .B2(P2_IR_REG_13__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5497) );
  XNOR2_X1 U6935 ( .A(n5497), .B(n5503), .ZN(n10127) );
  NAND2_X1 U6936 ( .A1(n5453), .A2(n5450), .ZN(n5455) );
  NAND2_X1 U6937 ( .A1(n5455), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5452) );
  INV_X1 U6938 ( .A(n5453), .ZN(n5454) );
  NAND2_X1 U6939 ( .A1(n5454), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n5456) );
  OR2_X1 U6940 ( .A1(n5457), .A2(n9152), .ZN(n5458) );
  XNOR2_X1 U6941 ( .A(n5458), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6216) );
  INV_X1 U6942 ( .A(n6216), .ZN(n7898) );
  OR2_X1 U6943 ( .A1(n5459), .A2(n9152), .ZN(n5460) );
  XNOR2_X1 U6944 ( .A(n5460), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U6945 ( .A1(n5461), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U6946 ( .A(n5462), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6194) );
  INV_X1 U6947 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7546) );
  NAND2_X1 U6948 ( .A1(n4357), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5463) );
  XNOR2_X1 U6949 ( .A(n5463), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7550) );
  INV_X1 U6950 ( .A(n7550), .ZN(n6866) );
  NAND2_X1 U6951 ( .A1(n5464), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5465) );
  INV_X1 U6952 ( .A(n7400), .ZN(n6849) );
  INV_X1 U6953 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6108) );
  NOR2_X1 U6954 ( .A1(n6108), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n5469) );
  NAND2_X1 U6955 ( .A1(n5466), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5470) );
  OAI21_X1 U6956 ( .B1(n7425), .B2(n5469), .A(n5470), .ZN(n7423) );
  INV_X1 U6957 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7424) );
  NOR2_X1 U6958 ( .A1(n7423), .A2(n7424), .ZN(n7422) );
  INV_X1 U6959 ( .A(n5470), .ZN(n5471) );
  NOR2_X1 U6960 ( .A1(n7422), .A2(n5471), .ZN(n6788) );
  XNOR2_X1 U6961 ( .A(n5531), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U6962 ( .A1(n5472), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5473) );
  INV_X1 U6963 ( .A(n5474), .ZN(n7390) );
  INV_X1 U6964 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7494) );
  MUX2_X1 U6965 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7494), .S(n7400), .Z(n7391)
         );
  AOI21_X1 U6966 ( .B1(P2_REG2_REG_4__SCAN_IN), .B2(n6849), .A(n7394), .ZN(
        n5475) );
  OR2_X1 U6967 ( .A1(n5476), .A2(n9152), .ZN(n5477) );
  XNOR2_X1 U6968 ( .A(n5477), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6165) );
  INV_X1 U6969 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6970 ( .A1(n5481), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5482) );
  MUX2_X1 U6971 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5482), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5483) );
  AND2_X1 U6972 ( .A1(n5483), .A2(n4357), .ZN(n6176) );
  XNOR2_X1 U6973 ( .A(n6176), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n7359) );
  OAI21_X1 U6974 ( .B1(n7378), .B2(n5484), .A(n7359), .ZN(n7362) );
  NOR2_X1 U6975 ( .A1(n7550), .A2(n4952), .ZN(n5486) );
  NOR2_X1 U6976 ( .A1(n7544), .A2(n5486), .ZN(n7742) );
  INV_X1 U6977 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7687) );
  AOI22_X1 U6978 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(n6194), .B1(n7750), .B2(
        n7687), .ZN(n7741) );
  NOR2_X1 U6979 ( .A1(n7828), .A2(n5487), .ZN(n5488) );
  INV_X1 U6980 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7825) );
  INV_X1 U6981 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n5489) );
  AOI22_X1 U6982 ( .A1(n6216), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n5489), .B2(
        n7898), .ZN(n7903) );
  NOR2_X1 U6983 ( .A1(n8714), .A2(n5490), .ZN(n5491) );
  INV_X1 U6984 ( .A(n8714), .ZN(n6900) );
  XNOR2_X1 U6985 ( .A(n5490), .B(n8714), .ZN(n8710) );
  INV_X1 U6986 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8711) );
  NAND2_X1 U6987 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8015), .ZN(n5492) );
  OAI21_X1 U6988 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n8015), .A(n5492), .ZN(
        n8020) );
  NOR2_X1 U6989 ( .A1(n8021), .A2(n8020), .ZN(n8019) );
  INV_X1 U6990 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5504) );
  XNOR2_X1 U6991 ( .A(n5493), .B(n5504), .ZN(n10091) );
  INV_X1 U6992 ( .A(n10091), .ZN(n6959) );
  INV_X1 U6993 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10094) );
  NOR2_X1 U6994 ( .A1(n10091), .A2(n5494), .ZN(n5495) );
  NAND2_X1 U6995 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10127), .ZN(n5496) );
  OAI21_X1 U6996 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n10127), .A(n5496), .ZN(
        n10111) );
  NAND2_X1 U6997 ( .A1(n5497), .A2(n5503), .ZN(n5498) );
  NAND2_X1 U6998 ( .A1(n5498), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5499) );
  XNOR2_X1 U6999 ( .A(n5499), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6977) );
  INV_X1 U7000 ( .A(n6977), .ZN(n8737) );
  INV_X1 U7001 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8728) );
  NOR2_X1 U7002 ( .A1(n6977), .A2(n5500), .ZN(n5501) );
  INV_X1 U7003 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5502) );
  NAND3_X1 U7004 ( .A1(n5504), .A2(n5503), .A3(n5502), .ZN(n5506) );
  NOR2_X1 U7005 ( .A1(n5506), .A2(n5505), .ZN(n5510) );
  NAND2_X1 U7006 ( .A1(n5511), .A2(n5510), .ZN(n5507) );
  NAND2_X1 U7007 ( .A1(n5507), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5508) );
  INV_X1 U7008 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5517) );
  XNOR2_X1 U7009 ( .A(n5508), .B(n5517), .ZN(n8755) );
  NAND2_X1 U7010 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8755), .ZN(n5509) );
  OAI21_X1 U7011 ( .B1(P2_REG2_REG_16__SCAN_IN), .B2(n8755), .A(n5509), .ZN(
        n8745) );
  NAND2_X1 U7012 ( .A1(n5519), .A2(n5517), .ZN(n5512) );
  NAND2_X1 U7013 ( .A1(n5512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  XNOR2_X1 U7014 ( .A(n5513), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8768) );
  INV_X1 U7015 ( .A(n8768), .ZN(n5558) );
  NAND2_X1 U7016 ( .A1(n5514), .A2(n5558), .ZN(n5515) );
  OAI21_X1 U7017 ( .B1(n5514), .B2(n5558), .A(n5515), .ZN(n8762) );
  INV_X1 U7018 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8962) );
  INV_X1 U7019 ( .A(n8765), .ZN(n5516) );
  NAND2_X1 U7020 ( .A1(n5516), .A2(n5515), .ZN(n8783) );
  AND2_X1 U7021 ( .A1(n5404), .A2(n5517), .ZN(n5518) );
  NAND2_X1 U7022 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  NAND2_X1 U7023 ( .A1(n5521), .A2(n7025), .ZN(n5526) );
  INV_X1 U7024 ( .A(n5521), .ZN(n5522) );
  NAND2_X1 U7025 ( .A1(n5522), .A2(P2_IR_REG_18__SCAN_IN), .ZN(n5523) );
  AND2_X1 U7026 ( .A1(n5526), .A2(n5523), .ZN(n8798) );
  INV_X1 U7027 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n6313) );
  OR2_X1 U7028 ( .A1(n8798), .A2(n6313), .ZN(n5525) );
  NAND2_X1 U7029 ( .A1(n8798), .A2(n6313), .ZN(n5524) );
  AND2_X1 U7030 ( .A1(n5525), .A2(n5524), .ZN(n8782) );
  INV_X1 U7031 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n5530) );
  INV_X1 U7032 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5527) );
  XNOR2_X2 U7033 ( .A(n5528), .B(n5527), .ZN(n6467) );
  MUX2_X1 U7034 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n5530), .S(n5529), .Z(n5568)
         );
  OR2_X1 U7035 ( .A1(n8510), .A2(P2_U3151), .ZN(n8214) );
  OR2_X1 U7036 ( .A1(n5614), .A2(n8214), .ZN(n10083) );
  NOR2_X1 U7037 ( .A1(n10083), .A2(n5612), .ZN(n8764) );
  XNOR2_X1 U7038 ( .A(n5531), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n6792) );
  AND2_X1 U7039 ( .A1(n10089), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U7040 ( .A1(n5466), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5534) );
  OAI21_X1 U7041 ( .B1(n5533), .B2(n5532), .A(n5534), .ZN(n7412) );
  INV_X1 U7042 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10225) );
  NOR2_X1 U7043 ( .A1(n7412), .A2(n10225), .ZN(n7414) );
  INV_X1 U7044 ( .A(n5534), .ZN(n5535) );
  NOR2_X1 U7045 ( .A1(n7414), .A2(n5535), .ZN(n6791) );
  NOR2_X1 U7046 ( .A1(n5536), .A2(n6140), .ZN(n5538) );
  NOR2_X1 U7047 ( .A1(n5538), .A2(n5537), .ZN(n7245) );
  INV_X1 U7048 ( .A(n5538), .ZN(n7395) );
  INV_X1 U7049 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6146) );
  MUX2_X1 U7050 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6146), .S(n7400), .Z(n7396)
         );
  AOI21_X1 U7051 ( .B1(P2_REG1_REG_4__SCAN_IN), .B2(n6849), .A(n7399), .ZN(
        n5539) );
  AOI21_X1 U7052 ( .B1(n5539), .B2(n6165), .A(n7365), .ZN(n7376) );
  NAND2_X1 U7053 ( .A1(n7376), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U7054 ( .A1(n7375), .A2(n5540), .ZN(n5543) );
  INV_X1 U7055 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n5541) );
  XNOR2_X1 U7056 ( .A(n6176), .B(n5541), .ZN(n7366) );
  INV_X1 U7057 ( .A(n7366), .ZN(n5542) );
  NOR2_X1 U7058 ( .A1(n7550), .A2(n5544), .ZN(n5545) );
  INV_X1 U7059 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10234) );
  NOR2_X1 U7060 ( .A1(n10234), .A2(n7549), .ZN(n7548) );
  NOR2_X1 U7061 ( .A1(n5545), .A2(n7548), .ZN(n7753) );
  INV_X1 U7062 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6197) );
  MUX2_X1 U7063 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6197), .S(n6194), .Z(n7752)
         );
  NOR2_X1 U7064 ( .A1(n7753), .A2(n7752), .ZN(n7751) );
  AOI21_X1 U7065 ( .B1(P2_REG1_REG_8__SCAN_IN), .B2(n7750), .A(n7751), .ZN(
        n5546) );
  NOR2_X1 U7066 ( .A1(n7828), .A2(n5546), .ZN(n5547) );
  INV_X1 U7067 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10237) );
  INV_X1 U7068 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6219) );
  MUX2_X1 U7069 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6219), .S(n6216), .Z(n7893)
         );
  NOR2_X1 U7070 ( .A1(n8714), .A2(n5548), .ZN(n5549) );
  INV_X1 U7071 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U7072 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8015), .ZN(n5550) );
  OAI21_X1 U7073 ( .B1(n8015), .B2(P2_REG1_REG_12__SCAN_IN), .A(n5550), .ZN(
        n8010) );
  AOI21_X2 U7074 ( .B1(P2_REG1_REG_12__SCAN_IN), .B2(n8015), .A(n8009), .ZN(
        n5551) );
  NOR2_X1 U7075 ( .A1(n10091), .A2(n5551), .ZN(n5552) );
  INV_X1 U7076 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10101) );
  NAND2_X1 U7077 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n10127), .ZN(n5553) );
  OAI21_X1 U7078 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n10127), .A(n5553), .ZN(
        n10116) );
  INV_X1 U7079 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8249) );
  NOR2_X1 U7080 ( .A1(n6977), .A2(n5554), .ZN(n5555) );
  NOR2_X1 U7081 ( .A1(n8731), .A2(n5555), .ZN(n8747) );
  XNOR2_X1 U7082 ( .A(n8755), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n8746) );
  NAND2_X1 U7083 ( .A1(n8755), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5556) );
  NAND2_X1 U7084 ( .A1(n8748), .A2(n5556), .ZN(n5557) );
  NOR2_X1 U7085 ( .A1(n5558), .A2(n5557), .ZN(n5559) );
  INV_X1 U7086 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9040) );
  INV_X1 U7087 ( .A(n8798), .ZN(n5561) );
  NAND2_X1 U7088 ( .A1(n5561), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n5562) );
  OAI21_X1 U7089 ( .B1(n5561), .B2(P2_REG1_REG_18__SCAN_IN), .A(n5562), .ZN(
        n8789) );
  INV_X1 U7090 ( .A(n5562), .ZN(n5563) );
  NOR2_X1 U7091 ( .A1(n8788), .A2(n5563), .ZN(n5564) );
  XNOR2_X1 U7092 ( .A(n5529), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n5566) );
  XNOR2_X1 U7093 ( .A(n5564), .B(n5566), .ZN(n5565) );
  INV_X1 U7094 ( .A(n5612), .ZN(n8511) );
  NOR2_X1 U7095 ( .A1(n10083), .A2(n8511), .ZN(n8777) );
  NAND2_X1 U7096 ( .A1(n5565), .A2(n8777), .ZN(n5623) );
  INV_X1 U7097 ( .A(n5566), .ZN(n5567) );
  MUX2_X1 U7098 ( .A(n5568), .B(n5567), .S(n5612), .Z(n5609) );
  MUX2_X1 U7099 ( .A(P2_REG2_REG_17__SCAN_IN), .B(P2_REG1_REG_17__SCAN_IN), 
        .S(n5612), .Z(n5569) );
  INV_X1 U7100 ( .A(n5569), .ZN(n5602) );
  XNOR2_X1 U7101 ( .A(n5569), .B(n8768), .ZN(n8774) );
  MUX2_X1 U7102 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n5612), .Z(n5570) );
  OR2_X1 U7103 ( .A1(n5570), .A2(n8755), .ZN(n5600) );
  INV_X1 U7104 ( .A(n8755), .ZN(n7198) );
  XNOR2_X1 U7105 ( .A(n5570), .B(n7198), .ZN(n8753) );
  MUX2_X1 U7106 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n5612), .Z(n5571) );
  OR2_X1 U7107 ( .A1(n5571), .A2(n8737), .ZN(n5599) );
  XNOR2_X1 U7108 ( .A(n6977), .B(n5571), .ZN(n8735) );
  INV_X1 U7109 ( .A(n10127), .ZN(n5572) );
  INV_X1 U7110 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8991) );
  INV_X1 U7111 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n9045) );
  MUX2_X1 U7112 ( .A(n8991), .B(n9045), .S(n5612), .Z(n5573) );
  NAND2_X1 U7113 ( .A1(n5572), .A2(n5573), .ZN(n5598) );
  XNOR2_X1 U7114 ( .A(n10127), .B(n5573), .ZN(n10114) );
  MUX2_X1 U7115 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n5612), .Z(n5574) );
  OR2_X1 U7116 ( .A1(n6959), .A2(n5574), .ZN(n5597) );
  XNOR2_X1 U7117 ( .A(n5574), .B(n10091), .ZN(n10097) );
  INV_X1 U7118 ( .A(n8015), .ZN(n5575) );
  INV_X1 U7119 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8042) );
  INV_X1 U7120 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6242) );
  MUX2_X1 U7121 ( .A(n8042), .B(n6242), .S(n5612), .Z(n5576) );
  NAND2_X1 U7122 ( .A1(n5575), .A2(n5576), .ZN(n5596) );
  XNOR2_X1 U7123 ( .A(n5576), .B(n8015), .ZN(n8013) );
  MUX2_X1 U7124 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n5612), .Z(n5577) );
  OR2_X1 U7125 ( .A1(n5577), .A2(n6900), .ZN(n5595) );
  XNOR2_X1 U7126 ( .A(n5577), .B(n8714), .ZN(n8719) );
  MUX2_X1 U7127 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n5612), .Z(n5578) );
  OR2_X1 U7128 ( .A1(n5578), .A2(n7898), .ZN(n5594) );
  XNOR2_X1 U7129 ( .A(n5578), .B(n6216), .ZN(n7896) );
  MUX2_X1 U7130 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n5612), .Z(n5580) );
  INV_X1 U7131 ( .A(n7828), .ZN(n5579) );
  OR2_X1 U7132 ( .A1(n5580), .A2(n5579), .ZN(n5593) );
  XNOR2_X1 U7133 ( .A(n5580), .B(n7828), .ZN(n7831) );
  MUX2_X1 U7134 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n5612), .Z(n5581) );
  OR2_X1 U7135 ( .A1(n5581), .A2(n7750), .ZN(n5592) );
  XNOR2_X1 U7136 ( .A(n5581), .B(n6194), .ZN(n7746) );
  MUX2_X1 U7137 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n5612), .Z(n5590) );
  OR2_X1 U7138 ( .A1(n5590), .A2(n6866), .ZN(n5591) );
  MUX2_X1 U7139 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n5612), .Z(n5589) );
  INV_X1 U7140 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6156) );
  MUX2_X1 U7141 ( .A(n5479), .B(n6156), .S(n5612), .Z(n5587) );
  INV_X1 U7142 ( .A(n5587), .ZN(n5588) );
  MUX2_X1 U7143 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n5612), .Z(n5586) );
  MUX2_X1 U7144 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n5612), .Z(n5585) );
  MUX2_X1 U7145 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n5612), .Z(n5584) );
  MUX2_X1 U7146 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n5612), .Z(n5582) );
  MUX2_X1 U7147 ( .A(P2_REG2_REG_0__SCAN_IN), .B(P2_REG1_REG_0__SCAN_IN), .S(
        n5612), .Z(n10084) );
  NOR2_X1 U7148 ( .A1(n10084), .A2(n10089), .ZN(n7416) );
  NOR2_X1 U7149 ( .A1(n7417), .A2(n7416), .ZN(n7415) );
  AOI21_X1 U7150 ( .B1(n5582), .B2(n7425), .A(n7415), .ZN(n6796) );
  XOR2_X1 U7151 ( .A(n5583), .B(n5584), .Z(n6797) );
  NOR2_X1 U7152 ( .A1(n6796), .A2(n6797), .ZN(n6795) );
  XNOR2_X1 U7153 ( .A(n5585), .B(n6140), .ZN(n7252) );
  NAND2_X1 U7154 ( .A1(n7253), .A2(n7252), .ZN(n7251) );
  OAI21_X1 U7155 ( .B1(n5585), .B2(n4742), .A(n7251), .ZN(n7407) );
  XOR2_X1 U7156 ( .A(n7400), .B(n5586), .Z(n7408) );
  NOR2_X1 U7157 ( .A1(n7407), .A2(n7408), .ZN(n7405) );
  XNOR2_X1 U7158 ( .A(n5587), .B(n6165), .ZN(n7386) );
  NOR2_X1 U7159 ( .A1(n7385), .A2(n7386), .ZN(n7384) );
  XNOR2_X1 U7160 ( .A(n5589), .B(n6176), .ZN(n7356) );
  NAND2_X1 U7161 ( .A1(n7357), .A2(n7356), .ZN(n7355) );
  OAI21_X1 U7162 ( .B1(n5589), .B2(n7364), .A(n7355), .ZN(n7543) );
  XNOR2_X1 U7163 ( .A(n5590), .B(n7550), .ZN(n7542) );
  NAND2_X1 U7164 ( .A1(n7543), .A2(n7542), .ZN(n7541) );
  NAND2_X1 U7165 ( .A1(n5591), .A2(n7541), .ZN(n7745) );
  NAND2_X1 U7166 ( .A1(n7746), .A2(n7745), .ZN(n7744) );
  NAND2_X1 U7167 ( .A1(n5592), .A2(n7744), .ZN(n7830) );
  NAND2_X1 U7168 ( .A1(n7896), .A2(n7895), .ZN(n7894) );
  NAND2_X1 U7169 ( .A1(n5594), .A2(n7894), .ZN(n8718) );
  NAND2_X1 U7170 ( .A1(n8719), .A2(n8718), .ZN(n8717) );
  NAND2_X1 U7171 ( .A1(n5595), .A2(n8717), .ZN(n8012) );
  NAND2_X1 U7172 ( .A1(n8013), .A2(n8012), .ZN(n8011) );
  NAND2_X1 U7173 ( .A1(n5596), .A2(n8011), .ZN(n10096) );
  NAND2_X1 U7174 ( .A1(n10097), .A2(n10096), .ZN(n10095) );
  NAND2_X1 U7175 ( .A1(n5597), .A2(n10095), .ZN(n10113) );
  NAND2_X1 U7176 ( .A1(n8735), .A2(n8734), .ZN(n8733) );
  NAND2_X1 U7177 ( .A1(n5599), .A2(n8733), .ZN(n8752) );
  NAND2_X1 U7178 ( .A1(n8774), .A2(n8773), .ZN(n8772) );
  INV_X1 U7179 ( .A(n8772), .ZN(n5601) );
  AOI21_X1 U7180 ( .B1(n5602), .B2(n8768), .A(n5601), .ZN(n5603) );
  MUX2_X1 U7181 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n5612), .Z(n5604) );
  INV_X1 U7182 ( .A(n5603), .ZN(n5606) );
  INV_X1 U7183 ( .A(n5604), .ZN(n5605) );
  NOR2_X1 U7184 ( .A1(n5606), .A2(n5605), .ZN(n8794) );
  INV_X1 U7185 ( .A(n8794), .ZN(n5607) );
  OAI21_X1 U7186 ( .B1(n8795), .B2(n8798), .A(n5607), .ZN(n5608) );
  XNOR2_X1 U7187 ( .A(n5609), .B(n5608), .ZN(n5620) );
  OR2_X2 U7188 ( .A1(n5615), .A2(P2_U3151), .ZN(n8705) );
  INV_X1 U7189 ( .A(n8510), .ZN(n6436) );
  INV_X1 U7190 ( .A(n5610), .ZN(n7406) );
  INV_X1 U7191 ( .A(n5615), .ZN(n5611) );
  NOR2_X2 U7192 ( .A1(P2_U3150), .A2(n5611), .ZN(n10109) );
  NOR2_X1 U7193 ( .A1(n5612), .A2(P2_U3151), .ZN(n8146) );
  NAND2_X1 U7194 ( .A1(n8146), .A2(n8510), .ZN(n5613) );
  OR2_X1 U7195 ( .A1(n5614), .A2(n5613), .ZN(n5617) );
  OR2_X1 U7196 ( .A1(n5615), .A2(n8214), .ZN(n5616) );
  NAND2_X1 U7197 ( .A1(n5617), .A2(n5616), .ZN(n10090) );
  NAND2_X1 U7198 ( .A1(P2_U3151), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8587) );
  OAI21_X1 U7199 ( .B1(n10128), .B2(n5529), .A(n8587), .ZN(n5618) );
  AOI21_X1 U7200 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n10109), .A(n5618), .ZN(
        n5619) );
  INV_X1 U7201 ( .A(n5621), .ZN(n5622) );
  INV_X1 U7202 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7203 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_REG3_REG_13__SCAN_IN), 
        .ZN(n5624) );
  INV_X1 U7204 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5806) );
  INV_X1 U7205 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5800) );
  INV_X1 U7206 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n9178) );
  INV_X1 U7207 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U7208 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5630) );
  INV_X1 U7209 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n9221) );
  INV_X1 U7210 ( .A(n5890), .ZN(n5631) );
  NAND2_X1 U7211 ( .A1(n5631), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n5896) );
  INV_X1 U7212 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6776) );
  NAND2_X1 U7213 ( .A1(n5890), .A2(n6776), .ZN(n5632) );
  AND2_X1 U7214 ( .A1(n5896), .A2(n5632), .ZN(n9479) );
  NAND2_X1 U7215 ( .A1(n9479), .A2(n5919), .ZN(n5639) );
  INV_X1 U7216 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9668) );
  NAND2_X1 U7217 ( .A1(n5934), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U7218 ( .A1(n4338), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5635) );
  OAI211_X1 U7219 ( .C1(n4327), .C2(n9668), .A(n5636), .B(n5635), .ZN(n5637)
         );
  INV_X1 U7220 ( .A(n5637), .ZN(n5638) );
  NAND2_X1 U7221 ( .A1(n5639), .A2(n5638), .ZN(n9297) );
  INV_X1 U7222 ( .A(n9297), .ZN(n8293) );
  NAND2_X1 U7223 ( .A1(n9478), .A2(n8293), .ZN(n8313) );
  XNOR2_X1 U7224 ( .A(n5875), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n9528) );
  NAND2_X1 U7225 ( .A1(n9528), .A2(n5919), .ZN(n5644) );
  INV_X1 U7226 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9683) );
  NAND2_X1 U7227 ( .A1(n5934), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U7228 ( .A1(n4338), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5640) );
  OAI211_X1 U7229 ( .C1(n4327), .C2(n9683), .A(n5641), .B(n5640), .ZN(n5642)
         );
  INV_X1 U7230 ( .A(n5642), .ZN(n5643) );
  OR2_X1 U7231 ( .A1(n9527), .A2(n9276), .ZN(n5872) );
  NAND2_X1 U7232 ( .A1(n9527), .A2(n9276), .ZN(n8310) );
  NAND2_X1 U7233 ( .A1(n5872), .A2(n8310), .ZN(n9519) );
  INV_X1 U7234 ( .A(n9519), .ZN(n9517) );
  INV_X1 U7235 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9279) );
  NAND2_X1 U7236 ( .A1(n5854), .A2(n9279), .ZN(n5645) );
  NAND2_X1 U7237 ( .A1(n5875), .A2(n5645), .ZN(n9536) );
  OR2_X1 U7238 ( .A1(n9536), .A2(n5898), .ZN(n5651) );
  INV_X1 U7239 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U7240 ( .A1(n5934), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5647) );
  NAND2_X1 U7241 ( .A1(n4339), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5646) );
  OAI211_X1 U7242 ( .C1(n4327), .C2(n5648), .A(n5647), .B(n5646), .ZN(n5649)
         );
  INV_X1 U7243 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7244 ( .A1(n5651), .A2(n5650), .ZN(n9301) );
  INV_X1 U7245 ( .A(n9301), .ZN(n8287) );
  OR2_X1 U7246 ( .A1(n9685), .A2(n8287), .ZN(n8309) );
  NAND2_X1 U7247 ( .A1(n9685), .A2(n8287), .ZN(n5871) );
  NAND2_X1 U7248 ( .A1(n9517), .A2(n9540), .ZN(n5964) );
  INV_X1 U7249 ( .A(n5964), .ZN(n5869) );
  INV_X1 U7250 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9268) );
  NAND2_X1 U7251 ( .A1(n5658), .A2(n9268), .ZN(n5652) );
  NAND2_X1 U7252 ( .A1(n5852), .A2(n5652), .ZN(n9266) );
  OR2_X1 U7253 ( .A1(n9266), .A2(n5898), .ZN(n5655) );
  AOI22_X1 U7254 ( .A1(n5934), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n4338), .B2(
        P1_REG0_REG_20__SCAN_IN), .ZN(n5654) );
  NAND2_X1 U7255 ( .A1(n5664), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U7256 ( .A1(n9697), .A2(n9177), .ZN(n9550) );
  NAND2_X1 U7257 ( .A1(n5862), .A2(n5932), .ZN(n5656) );
  OAI21_X1 U7258 ( .B1(n9565), .B2(n9587), .A(n5656), .ZN(n5663) );
  NAND2_X1 U7259 ( .A1(n5846), .A2(n9178), .ZN(n5657) );
  NAND2_X1 U7260 ( .A1(n5658), .A2(n5657), .ZN(n9583) );
  INV_X1 U7261 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9584) );
  OAI22_X1 U7262 ( .A1(n9583), .A2(n5898), .B1(n4341), .B2(n9584), .ZN(n5661)
         );
  INV_X1 U7263 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9704) );
  NAND2_X1 U7264 ( .A1(n4339), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5659) );
  OAI21_X1 U7265 ( .B1(n9704), .B2(n4327), .A(n5659), .ZN(n5660) );
  INV_X1 U7266 ( .A(n9304), .ZN(n8283) );
  OR2_X1 U7267 ( .A1(n9587), .A2(n8283), .ZN(n5942) );
  AND3_X1 U7268 ( .A1(n9550), .A2(n9304), .A3(n6075), .ZN(n5662) );
  AOI21_X1 U7269 ( .B1(n5663), .B2(n5942), .A(n5662), .ZN(n5865) );
  INV_X1 U7270 ( .A(n5865), .ZN(n5857) );
  INV_X1 U7271 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6830) );
  OR2_X1 U7272 ( .A1(n5832), .A2(n6830), .ZN(n5668) );
  NAND2_X1 U7273 ( .A1(n5756), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5666) );
  INV_X1 U7274 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9325) );
  OR2_X1 U7275 ( .A1(n5693), .A2(n9325), .ZN(n5665) );
  NAND2_X1 U7276 ( .A1(n4339), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5673) );
  INV_X1 U7277 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7567) );
  OR2_X1 U7278 ( .A1(n5693), .A2(n7567), .ZN(n5672) );
  INV_X1 U7279 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5669) );
  OR2_X1 U7280 ( .A1(n4340), .A2(n5669), .ZN(n5671) );
  INV_X1 U7281 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6875) );
  OR2_X1 U7282 ( .A1(n5688), .A2(n6875), .ZN(n5670) );
  NAND2_X1 U7283 ( .A1(n4461), .A2(n10034), .ZN(n5674) );
  NAND2_X1 U7284 ( .A1(n5675), .A2(n5674), .ZN(n7653) );
  INV_X1 U7285 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n5676) );
  OR2_X1 U7286 ( .A1(n4341), .A2(n5676), .ZN(n5681) );
  INV_X1 U7287 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9338) );
  OR2_X1 U7288 ( .A1(n5693), .A2(n9338), .ZN(n5680) );
  NAND2_X1 U7289 ( .A1(n4338), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5679) );
  INV_X1 U7290 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5677) );
  OR2_X1 U7291 ( .A1(n5688), .A2(n5677), .ZN(n5678) );
  INV_X1 U7292 ( .A(n7652), .ZN(n5954) );
  NAND2_X1 U7293 ( .A1(n7653), .A2(n5954), .ZN(n5683) );
  INV_X1 U7294 ( .A(n10050), .ZN(n7650) );
  NAND2_X1 U7295 ( .A1(n7304), .A2(n7650), .ZN(n5682) );
  NAND2_X1 U7296 ( .A1(n4339), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n5687) );
  INV_X1 U7297 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6819) );
  OR2_X1 U7298 ( .A1(n4327), .A2(n6819), .ZN(n5686) );
  INV_X1 U7299 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10022) );
  OR2_X1 U7300 ( .A1(n4341), .A2(n10022), .ZN(n5685) );
  OR2_X1 U7301 ( .A1(n5898), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5684) );
  OR2_X1 U7302 ( .A1(n9320), .A2(n7431), .ZN(n5951) );
  NAND2_X1 U7303 ( .A1(n9320), .A2(n7431), .ZN(n7464) );
  NAND2_X1 U7304 ( .A1(n4338), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5697) );
  INV_X1 U7305 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6815) );
  OR2_X1 U7306 ( .A1(n4327), .A2(n6815), .ZN(n5696) );
  INV_X1 U7307 ( .A(n5689), .ZN(n5702) );
  INV_X1 U7308 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5691) );
  INV_X1 U7309 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U7310 ( .A1(n5691), .A2(n5690), .ZN(n5692) );
  NAND2_X1 U7311 ( .A1(n5702), .A2(n5692), .ZN(n7590) );
  OR2_X1 U7312 ( .A1(n5898), .A2(n7590), .ZN(n5695) );
  INV_X1 U7313 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6829) );
  OR2_X1 U7314 ( .A1(n4340), .A2(n6829), .ZN(n5694) );
  NAND4_X1 U7315 ( .A1(n5697), .A2(n5696), .A3(n5695), .A4(n5694), .ZN(n9319)
         );
  NAND2_X1 U7316 ( .A1(n9319), .A2(n7593), .ZN(n5992) );
  AND2_X1 U7317 ( .A1(n7464), .A2(n5992), .ZN(n5698) );
  OR2_X1 U7318 ( .A1(n9319), .A2(n7593), .ZN(n5950) );
  NAND2_X1 U7319 ( .A1(n5664), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5708) );
  INV_X1 U7320 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5699) );
  OR2_X1 U7321 ( .A1(n5909), .A2(n5699), .ZN(n5707) );
  INV_X1 U7322 ( .A(n5700), .ZN(n5711) );
  INV_X1 U7323 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U7324 ( .A1(n5702), .A2(n5701), .ZN(n5703) );
  NAND2_X1 U7325 ( .A1(n5711), .A2(n5703), .ZN(n7579) );
  OR2_X1 U7326 ( .A1(n5693), .A2(n7579), .ZN(n5706) );
  INV_X1 U7327 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5704) );
  OR2_X1 U7328 ( .A1(n4340), .A2(n5704), .ZN(n5705) );
  NAND2_X1 U7329 ( .A1(n5664), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5717) );
  INV_X1 U7330 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5709) );
  OR2_X1 U7331 ( .A1(n5909), .A2(n5709), .ZN(n5716) );
  INV_X1 U7332 ( .A(n5726), .ZN(n5713) );
  INV_X1 U7333 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5710) );
  NAND2_X1 U7334 ( .A1(n5711), .A2(n5710), .ZN(n5712) );
  NAND2_X1 U7335 ( .A1(n5713), .A2(n5712), .ZN(n7714) );
  OR2_X1 U7336 ( .A1(n5693), .A2(n7714), .ZN(n5715) );
  INV_X1 U7337 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7617) );
  OR2_X1 U7338 ( .A1(n4341), .A2(n7617), .ZN(n5714) );
  OR2_X1 U7339 ( .A1(n9318), .A2(n7582), .ZN(n5994) );
  AND4_X1 U7340 ( .A1(n7633), .A2(n5994), .A3(n5950), .A4(n6075), .ZN(n5723)
         );
  INV_X1 U7341 ( .A(n5994), .ZN(n5718) );
  NAND3_X1 U7342 ( .A1(n5719), .A2(n5718), .A3(n5932), .ZN(n5721) );
  NAND3_X1 U7343 ( .A1(n7634), .A2(n7633), .A3(n6075), .ZN(n5720) );
  OAI211_X1 U7344 ( .C1(n6075), .C2(n7633), .A(n5721), .B(n5720), .ZN(n5722)
         );
  AOI21_X1 U7345 ( .B1(n5724), .B2(n5723), .A(n5722), .ZN(n5732) );
  NAND2_X1 U7346 ( .A1(n5664), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5731) );
  INV_X1 U7347 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5725) );
  OR2_X1 U7348 ( .A1(n5909), .A2(n5725), .ZN(n5730) );
  OAI21_X1 U7349 ( .B1(n5726), .B2(P1_REG3_REG_7__SCAN_IN), .A(n5736), .ZN(
        n7665) );
  INV_X1 U7350 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n5727) );
  XNOR2_X1 U7351 ( .A(n9316), .B(n7697), .ZN(n7636) );
  INV_X1 U7352 ( .A(n7636), .ZN(n7795) );
  NAND2_X1 U7353 ( .A1(n4339), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5742) );
  INV_X1 U7354 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5734) );
  OR2_X1 U7355 ( .A1(n4327), .A2(n5734), .ZN(n5741) );
  AND2_X1 U7356 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  OR2_X1 U7357 ( .A1(n5737), .A2(n5747), .ZN(n10010) );
  OR2_X1 U7358 ( .A1(n5898), .A2(n10010), .ZN(n5740) );
  INV_X1 U7359 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5738) );
  OR2_X1 U7360 ( .A1(n4341), .A2(n5738), .ZN(n5739) );
  OR2_X1 U7361 ( .A1(n10012), .A2(n7788), .ZN(n7787) );
  NAND2_X1 U7362 ( .A1(n7697), .A2(n9316), .ZN(n5743) );
  AND2_X1 U7363 ( .A1(n7787), .A2(n5743), .ZN(n5949) );
  NAND2_X1 U7364 ( .A1(n10012), .A2(n7788), .ZN(n7786) );
  INV_X1 U7365 ( .A(n9316), .ZN(n5744) );
  NAND2_X1 U7366 ( .A1(n5744), .A2(n7784), .ZN(n7793) );
  NAND2_X1 U7367 ( .A1(n7786), .A2(n7793), .ZN(n5947) );
  INV_X1 U7368 ( .A(n5947), .ZN(n5745) );
  MUX2_X1 U7369 ( .A(n5949), .B(n5745), .S(n6075), .Z(n5746) );
  NAND2_X1 U7370 ( .A1(n4339), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5752) );
  INV_X1 U7371 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n9371) );
  OR2_X1 U7372 ( .A1(n4327), .A2(n9371), .ZN(n5751) );
  NOR2_X1 U7373 ( .A1(n5747), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5748) );
  OR2_X1 U7374 ( .A1(n5757), .A2(n5748), .ZN(n7803) );
  OR2_X1 U7375 ( .A1(n5898), .A2(n7803), .ZN(n5750) );
  INV_X1 U7376 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9364) );
  OR2_X1 U7377 ( .A1(n4340), .A2(n9364), .ZN(n5749) );
  AND2_X1 U7378 ( .A1(n7791), .A2(n7787), .ZN(n5753) );
  MUX2_X1 U7379 ( .A(n7786), .B(n5753), .S(n6075), .Z(n5754) );
  NAND2_X1 U7380 ( .A1(n7952), .A2(n7881), .ZN(n7790) );
  NAND2_X1 U7381 ( .A1(n5777), .A2(n7790), .ZN(n5770) );
  NAND2_X1 U7382 ( .A1(n4339), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5762) );
  NOR2_X1 U7383 ( .A1(n5757), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5758) );
  OR2_X1 U7384 ( .A1(n5764), .A2(n5758), .ZN(n9865) );
  OR2_X1 U7385 ( .A1(n5898), .A2(n9865), .ZN(n5761) );
  INV_X1 U7386 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7873) );
  OR2_X1 U7387 ( .A1(n4341), .A2(n7873), .ZN(n5760) );
  INV_X1 U7388 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9401) );
  OR2_X1 U7389 ( .A1(n4327), .A2(n9401), .ZN(n5759) );
  NAND2_X1 U7390 ( .A1(n4338), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5769) );
  INV_X1 U7391 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n9402) );
  OR2_X1 U7392 ( .A1(n4327), .A2(n9402), .ZN(n5768) );
  INV_X1 U7393 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n5763) );
  OR2_X1 U7394 ( .A1(n4340), .A2(n5763), .ZN(n5767) );
  OR2_X1 U7395 ( .A1(n5764), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5765) );
  NAND2_X1 U7396 ( .A1(n5785), .A2(n5765), .ZN(n9889) );
  OR2_X1 U7397 ( .A1(n5898), .A2(n9889), .ZN(n5766) );
  NAND4_X1 U7398 ( .A1(n5769), .A2(n5768), .A3(n5767), .A4(n5766), .ZN(n9312)
         );
  NAND2_X1 U7399 ( .A1(n9886), .A2(n7983), .ZN(n5946) );
  NAND2_X1 U7400 ( .A1(n5946), .A2(n8226), .ZN(n6004) );
  AOI21_X1 U7401 ( .B1(n5770), .B2(n6000), .A(n6004), .ZN(n5775) );
  NAND2_X1 U7402 ( .A1(n4338), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5774) );
  INV_X1 U7403 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5784) );
  XNOR2_X1 U7404 ( .A(n5785), .B(n5784), .ZN(n9874) );
  OR2_X1 U7405 ( .A1(n5898), .A2(n9874), .ZN(n5773) );
  INV_X1 U7406 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7987) );
  OR2_X1 U7407 ( .A1(n4341), .A2(n7987), .ZN(n5772) );
  INV_X1 U7408 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9403) );
  OR2_X1 U7409 ( .A1(n4327), .A2(n9403), .ZN(n5771) );
  NAND4_X1 U7410 ( .A1(n5774), .A2(n5773), .A3(n5772), .A4(n5771), .ZN(n9311)
         );
  INV_X1 U7411 ( .A(n9311), .ZN(n8091) );
  OR2_X1 U7412 ( .A1(n9872), .A2(n8091), .ZN(n8094) );
  OR2_X1 U7413 ( .A1(n9886), .A2(n7983), .ZN(n6042) );
  NAND2_X1 U7414 ( .A1(n8094), .A2(n6042), .ZN(n6007) );
  NAND2_X1 U7415 ( .A1(n9872), .A2(n8091), .ZN(n6006) );
  OAI21_X1 U7416 ( .B1(n5775), .B2(n6007), .A(n6006), .ZN(n5782) );
  INV_X1 U7417 ( .A(n7790), .ZN(n5776) );
  NAND2_X1 U7418 ( .A1(n5778), .A2(n8226), .ZN(n5779) );
  NAND2_X1 U7419 ( .A1(n5780), .A2(n8094), .ZN(n5781) );
  NAND2_X1 U7420 ( .A1(n4338), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n5790) );
  INV_X1 U7421 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9396) );
  OR2_X1 U7422 ( .A1(n4327), .A2(n9396), .ZN(n5789) );
  INV_X1 U7423 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5783) );
  OAI21_X1 U7424 ( .B1(n5785), .B2(n5784), .A(n5783), .ZN(n5786) );
  NAND2_X1 U7425 ( .A1(n5786), .A2(n5792), .ZN(n7927) );
  OR2_X1 U7426 ( .A1(n5898), .A2(n7927), .ZN(n5788) );
  INV_X1 U7427 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9380) );
  OR2_X1 U7428 ( .A1(n4340), .A2(n9380), .ZN(n5787) );
  NAND2_X1 U7429 ( .A1(n8163), .A2(n8105), .ZN(n6045) );
  NAND2_X1 U7430 ( .A1(n5822), .A2(n6045), .ZN(n5799) );
  NAND2_X1 U7431 ( .A1(n4339), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n5798) );
  INV_X1 U7432 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9406) );
  OR2_X1 U7433 ( .A1(n4327), .A2(n9406), .ZN(n5797) );
  INV_X1 U7434 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7435 ( .A1(n5792), .A2(n5791), .ZN(n5793) );
  NAND2_X1 U7436 ( .A1(n5807), .A2(n5793), .ZN(n8135) );
  OR2_X1 U7437 ( .A1(n5898), .A2(n8135), .ZN(n5796) );
  INV_X1 U7438 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n5794) );
  OR2_X1 U7439 ( .A1(n4341), .A2(n5794), .ZN(n5795) );
  NAND4_X1 U7440 ( .A1(n5798), .A2(n5797), .A3(n5796), .A4(n5795), .ZN(n9309)
         );
  INV_X1 U7441 ( .A(n9309), .ZN(n8193) );
  OR2_X1 U7442 ( .A1(n9728), .A2(n8193), .ZN(n8202) );
  NAND2_X1 U7443 ( .A1(n9728), .A2(n8193), .ZN(n5814) );
  NAND2_X1 U7444 ( .A1(n8202), .A2(n5814), .ZN(n8130) );
  INV_X1 U7445 ( .A(n8130), .ZN(n8129) );
  NAND2_X1 U7446 ( .A1(n5799), .A2(n8129), .ZN(n5821) );
  NAND2_X1 U7447 ( .A1(n4339), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5805) );
  INV_X1 U7448 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9719) );
  OR2_X1 U7449 ( .A1(n4327), .A2(n9719), .ZN(n5804) );
  NAND2_X1 U7450 ( .A1(n5809), .A2(n5800), .ZN(n5801) );
  NAND2_X1 U7451 ( .A1(n5834), .A2(n5801), .ZN(n9630) );
  OR2_X1 U7452 ( .A1(n5898), .A2(n9630), .ZN(n5803) );
  INV_X1 U7453 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9631) );
  OR2_X1 U7454 ( .A1(n4341), .A2(n9631), .ZN(n5802) );
  NAND2_X1 U7455 ( .A1(n9628), .A2(n9240), .ZN(n6051) );
  NAND2_X1 U7456 ( .A1(n4338), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5813) );
  INV_X1 U7457 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9954) );
  OR2_X1 U7458 ( .A1(n4327), .A2(n9954), .ZN(n5812) );
  NAND2_X1 U7459 ( .A1(n5807), .A2(n5806), .ZN(n5808) );
  NAND2_X1 U7460 ( .A1(n5809), .A2(n5808), .ZN(n8198) );
  OR2_X1 U7461 ( .A1(n5898), .A2(n8198), .ZN(n5811) );
  INV_X1 U7462 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8199) );
  OR2_X1 U7463 ( .A1(n4340), .A2(n8199), .ZN(n5810) );
  NAND4_X1 U7464 ( .A1(n5813), .A2(n5812), .A3(n5811), .A4(n5810), .ZN(n9308)
         );
  INV_X1 U7465 ( .A(n9308), .ZN(n8277) );
  NAND2_X1 U7466 ( .A1(n8274), .A2(n8277), .ZN(n6049) );
  AND2_X1 U7467 ( .A1(n6049), .A2(n5814), .ZN(n6013) );
  AND2_X1 U7468 ( .A1(n6051), .A2(n6013), .ZN(n5820) );
  NAND2_X1 U7469 ( .A1(n6051), .A2(n9308), .ZN(n5815) );
  NAND2_X1 U7470 ( .A1(n5815), .A2(n5932), .ZN(n5829) );
  NAND2_X1 U7471 ( .A1(n5829), .A2(n9781), .ZN(n5818) );
  OR2_X1 U7472 ( .A1(n8163), .A2(n8105), .ZN(n6009) );
  INV_X1 U7473 ( .A(n6009), .ZN(n5816) );
  NAND3_X1 U7474 ( .A1(n6051), .A2(n5816), .A3(n6013), .ZN(n5817) );
  NAND3_X1 U7475 ( .A1(n5818), .A2(n5944), .A3(n5817), .ZN(n5819) );
  AOI21_X1 U7476 ( .B1(n5821), .B2(n5820), .A(n5819), .ZN(n5827) );
  NAND2_X1 U7477 ( .A1(n5822), .A2(n6009), .ZN(n5823) );
  OR2_X1 U7478 ( .A1(n8274), .A2(n8277), .ZN(n5945) );
  NAND2_X1 U7479 ( .A1(n5944), .A2(n5945), .ZN(n6011) );
  INV_X1 U7480 ( .A(n8202), .ZN(n6046) );
  NOR2_X1 U7481 ( .A1(n6011), .A2(n6046), .ZN(n5824) );
  INV_X1 U7482 ( .A(n6051), .ZN(n6015) );
  AOI21_X1 U7483 ( .B1(n5825), .B2(n5824), .A(n6015), .ZN(n5826) );
  INV_X1 U7484 ( .A(n6049), .ZN(n5828) );
  NAND3_X1 U7485 ( .A1(n5829), .A2(n5828), .A3(n5944), .ZN(n5830) );
  NAND2_X1 U7486 ( .A1(n5831), .A2(n5830), .ZN(n5841) );
  INV_X1 U7487 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n9770) );
  OR2_X1 U7488 ( .A1(n5909), .A2(n9770), .ZN(n5839) );
  INV_X1 U7489 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9612) );
  OR2_X1 U7490 ( .A1(n4340), .A2(n9612), .ZN(n5838) );
  INV_X1 U7491 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7492 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  NAND2_X1 U7493 ( .A1(n5844), .A2(n5835), .ZN(n9611) );
  OR2_X1 U7494 ( .A1(n5898), .A2(n9611), .ZN(n5837) );
  INV_X1 U7495 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9714) );
  OR2_X1 U7496 ( .A1(n4327), .A2(n9714), .ZN(n5836) );
  NAND4_X1 U7497 ( .A1(n5839), .A2(n5838), .A3(n5837), .A4(n5836), .ZN(n9306)
         );
  INV_X1 U7498 ( .A(n9306), .ZN(n8279) );
  OR2_X1 U7499 ( .A1(n9610), .A2(n8279), .ZN(n9591) );
  INV_X1 U7500 ( .A(n9591), .ZN(n5840) );
  AND2_X1 U7501 ( .A1(n9610), .A2(n8279), .ZN(n6052) );
  OR2_X1 U7502 ( .A1(n5840), .A2(n6052), .ZN(n9607) );
  INV_X1 U7503 ( .A(n9607), .ZN(n9615) );
  NAND2_X1 U7504 ( .A1(n5841), .A2(n9615), .ZN(n5861) );
  NAND2_X1 U7505 ( .A1(n4339), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5850) );
  INV_X1 U7506 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n5842) );
  OR2_X1 U7507 ( .A1(n4340), .A2(n5842), .ZN(n5849) );
  INV_X1 U7508 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5843) );
  NAND2_X1 U7509 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  NAND2_X1 U7510 ( .A1(n5846), .A2(n5845), .ZN(n9600) );
  OR2_X1 U7511 ( .A1(n5898), .A2(n9600), .ZN(n5848) );
  INV_X1 U7512 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n7155) );
  OR2_X1 U7513 ( .A1(n4327), .A2(n7155), .ZN(n5847) );
  NAND4_X1 U7514 ( .A1(n5850), .A2(n5849), .A3(n5848), .A4(n5847), .ZN(n9305)
         );
  INV_X1 U7515 ( .A(n9305), .ZN(n9176) );
  OR2_X1 U7516 ( .A1(n9708), .A2(n9176), .ZN(n5943) );
  AND2_X1 U7517 ( .A1(n5943), .A2(n9591), .ZN(n6053) );
  NAND2_X1 U7518 ( .A1(n5861), .A2(n6053), .ZN(n5851) );
  NAND2_X1 U7519 ( .A1(n9587), .A2(n8283), .ZN(n6056) );
  NAND2_X1 U7520 ( .A1(n9708), .A2(n9176), .ZN(n6054) );
  NAND2_X1 U7521 ( .A1(n5852), .A2(n9212), .ZN(n5853) );
  NAND2_X1 U7522 ( .A1(n5854), .A2(n5853), .ZN(n9211) );
  AOI22_X1 U7523 ( .A1(n5664), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n4338), .B2(
        P1_REG0_REG_21__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U7524 ( .A1(n5934), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5855) );
  OAI211_X1 U7525 ( .C1(n9211), .C2(n5898), .A(n5856), .B(n5855), .ZN(n9302)
         );
  INV_X1 U7526 ( .A(n9302), .ZN(n8286) );
  NAND2_X1 U7527 ( .A1(n9558), .A2(n8286), .ZN(n5866) );
  NAND2_X1 U7528 ( .A1(n5866), .A2(n9550), .ZN(n5984) );
  OR2_X1 U7529 ( .A1(n9558), .A2(n8286), .ZN(n5983) );
  INV_X1 U7530 ( .A(n5983), .ZN(n5858) );
  INV_X1 U7531 ( .A(n6052), .ZN(n5860) );
  AND2_X1 U7532 ( .A1(n6054), .A2(n5860), .ZN(n6018) );
  NAND2_X1 U7533 ( .A1(n5942), .A2(n5943), .ZN(n6016) );
  AOI21_X1 U7534 ( .B1(n5861), .B2(n6018), .A(n6016), .ZN(n5864) );
  NAND2_X1 U7535 ( .A1(n5983), .A2(n5862), .ZN(n8306) );
  INV_X1 U7536 ( .A(n8306), .ZN(n5863) );
  OAI21_X1 U7537 ( .B1(n5865), .B2(n5864), .A(n5863), .ZN(n5867) );
  NAND2_X1 U7538 ( .A1(n5872), .A2(n8309), .ZN(n5870) );
  NAND2_X1 U7539 ( .A1(n5870), .A2(n8310), .ZN(n5980) );
  AND2_X1 U7540 ( .A1(n8310), .A2(n5871), .ZN(n5985) );
  INV_X1 U7541 ( .A(n5985), .ZN(n5873) );
  NAND2_X1 U7542 ( .A1(n5873), .A2(n5872), .ZN(n5874) );
  MUX2_X1 U7543 ( .A(n5980), .B(n5874), .S(n6075), .Z(n5882) );
  INV_X1 U7544 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9166) );
  INV_X1 U7545 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n9256) );
  OAI21_X1 U7546 ( .B1(n5875), .B2(n9166), .A(n9256), .ZN(n5876) );
  NAND2_X1 U7547 ( .A1(n5876), .A2(n5888), .ZN(n9504) );
  OR2_X1 U7548 ( .A1(n9504), .A2(n5898), .ZN(n5881) );
  INV_X1 U7549 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9503) );
  NAND2_X1 U7550 ( .A1(n5664), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U7551 ( .A1(n4339), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5877) );
  OAI211_X1 U7552 ( .C1(n9503), .C2(n4340), .A(n5878), .B(n5877), .ZN(n5879)
         );
  INV_X1 U7553 ( .A(n5879), .ZN(n5880) );
  NAND2_X1 U7554 ( .A1(n5881), .A2(n5880), .ZN(n9299) );
  INV_X1 U7555 ( .A(n9299), .ZN(n8290) );
  NAND2_X1 U7556 ( .A1(n9502), .A2(n8290), .ZN(n5986) );
  AOI21_X1 U7557 ( .B1(n5883), .B2(n5882), .A(n9507), .ZN(n5887) );
  INV_X1 U7558 ( .A(n8311), .ZN(n5885) );
  INV_X1 U7559 ( .A(n5986), .ZN(n5884) );
  MUX2_X1 U7560 ( .A(n5885), .B(n5884), .S(n6075), .Z(n5886) );
  NAND2_X1 U7561 ( .A1(n5888), .A2(n9221), .ZN(n5889) );
  NAND2_X1 U7562 ( .A1(n5890), .A2(n5889), .ZN(n9222) );
  INV_X1 U7563 ( .A(n9222), .ZN(n9494) );
  INV_X1 U7564 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9673) );
  NAND2_X1 U7565 ( .A1(n4338), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5892) );
  NAND2_X1 U7566 ( .A1(n5934), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5891) );
  OAI211_X1 U7567 ( .C1(n4327), .C2(n9673), .A(n5892), .B(n5891), .ZN(n5893)
         );
  NAND2_X1 U7568 ( .A1(n9493), .A2(n9252), .ZN(n5987) );
  INV_X1 U7569 ( .A(n5987), .ZN(n5894) );
  OR2_X1 U7570 ( .A1(n9478), .A2(n8293), .ZN(n5978) );
  AND2_X1 U7571 ( .A1(n5978), .A2(n8312), .ZN(n5906) );
  OAI21_X1 U7572 ( .B1(n5908), .B2(n5894), .A(n5906), .ZN(n5905) );
  INV_X1 U7573 ( .A(n5896), .ZN(n5895) );
  NAND2_X1 U7574 ( .A1(n5895), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8301) );
  INV_X1 U7575 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U7576 ( .A1(n5896), .A2(n8270), .ZN(n5897) );
  NAND2_X1 U7577 ( .A1(n8301), .A2(n5897), .ZN(n9462) );
  OR2_X1 U7578 ( .A1(n9462), .A2(n5898), .ZN(n5903) );
  INV_X1 U7579 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U7580 ( .A1(n4339), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7581 ( .A1(n5934), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5899) );
  OAI211_X1 U7582 ( .C1(n4327), .C2(n9663), .A(n5900), .B(n5899), .ZN(n5901)
         );
  INV_X1 U7583 ( .A(n5901), .ZN(n5902) );
  NAND2_X1 U7584 ( .A1(n9461), .A2(n9197), .ZN(n8314) );
  INV_X1 U7585 ( .A(n9453), .ZN(n5904) );
  AOI211_X1 U7586 ( .C1(n8313), .C2(n5905), .A(n6075), .B(n5904), .ZN(n5929)
         );
  INV_X1 U7587 ( .A(n5906), .ZN(n5907) );
  AOI21_X1 U7588 ( .B1(n5908), .B2(n5987), .A(n5907), .ZN(n5918) );
  NAND3_X1 U7589 ( .A1(n9453), .A2(n8313), .A3(n6075), .ZN(n5917) );
  OAI21_X1 U7590 ( .B1(n9296), .B2(n6075), .A(n9461), .ZN(n5915) );
  OAI21_X1 U7591 ( .B1(n9197), .B2(n5932), .A(n9741), .ZN(n5914) );
  XNOR2_X1 U7592 ( .A(n8301), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n9440) );
  INV_X1 U7593 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n5912) );
  NAND2_X1 U7594 ( .A1(n5664), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5911) );
  INV_X1 U7595 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7032) );
  OR2_X1 U7596 ( .A1(n5909), .A2(n7032), .ZN(n5910) );
  OAI211_X1 U7597 ( .C1(n5912), .C2(n4341), .A(n5911), .B(n5910), .ZN(n5913)
         );
  AOI21_X1 U7598 ( .B1(n9440), .B2(n5919), .A(n5913), .ZN(n9189) );
  INV_X1 U7599 ( .A(n5941), .ZN(n8315) );
  AOI21_X1 U7600 ( .B1(n5915), .B2(n5914), .A(n8315), .ZN(n5916) );
  OAI211_X1 U7601 ( .C1(n5918), .C2(n5917), .A(n5916), .B(n6023), .ZN(n5928)
         );
  NAND2_X1 U7602 ( .A1(n5919), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7603 ( .A1(n8301), .A2(n5920), .ZN(n5926) );
  INV_X1 U7604 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5923) );
  NAND2_X1 U7605 ( .A1(n5934), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5922) );
  NAND2_X1 U7606 ( .A1(n4338), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5921) );
  OAI211_X1 U7607 ( .C1(n4327), .C2(n5923), .A(n5922), .B(n5921), .ZN(n5924)
         );
  INV_X1 U7608 ( .A(n5924), .ZN(n5925) );
  NAND2_X1 U7609 ( .A1(n9650), .A2(n9196), .ZN(n5976) );
  MUX2_X1 U7610 ( .A(n6023), .B(n5941), .S(n6075), .Z(n5927) );
  MUX2_X1 U7611 ( .A(n5976), .B(n6029), .S(n6075), .Z(n5930) );
  NAND2_X1 U7612 ( .A1(n5931), .A2(n5930), .ZN(n5939) );
  INV_X1 U7613 ( .A(n6891), .ZN(n5933) );
  INV_X1 U7614 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5937) );
  NAND2_X1 U7615 ( .A1(n5934), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5936) );
  NAND2_X1 U7616 ( .A1(n4339), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5935) );
  OAI211_X1 U7617 ( .C1(n4327), .C2(n5937), .A(n5936), .B(n5935), .ZN(n9294)
         );
  OAI21_X1 U7618 ( .B1(n9646), .B2(n9294), .A(n6891), .ZN(n5938) );
  NAND2_X1 U7619 ( .A1(n9646), .A2(n6891), .ZN(n6064) );
  NAND2_X1 U7620 ( .A1(n6023), .A2(n5941), .ZN(n9437) );
  INV_X1 U7621 ( .A(n9470), .ZN(n5966) );
  XNOR2_X1 U7622 ( .A(n9558), .B(n9302), .ZN(n9551) );
  INV_X1 U7623 ( .A(n9565), .ZN(n9567) );
  NAND2_X1 U7624 ( .A1(n5943), .A2(n6054), .ZN(n9594) );
  NAND2_X1 U7625 ( .A1(n5944), .A2(n6051), .ZN(n8278) );
  INV_X1 U7626 ( .A(n8278), .ZN(n9634) );
  NAND2_X1 U7627 ( .A1(n5945), .A2(n6049), .ZN(n6047) );
  INV_X1 U7628 ( .A(n6047), .ZN(n8204) );
  NAND2_X1 U7629 ( .A1(n6042), .A2(n5946), .ZN(n6040) );
  INV_X1 U7630 ( .A(n6040), .ZN(n8225) );
  NAND2_X1 U7631 ( .A1(n5947), .A2(n7787), .ZN(n7797) );
  NAND2_X1 U7632 ( .A1(n7797), .A2(n7790), .ZN(n5948) );
  NAND2_X1 U7633 ( .A1(n5948), .A2(n7791), .ZN(n5999) );
  AND2_X1 U7634 ( .A1(n5999), .A2(n7633), .ZN(n6037) );
  NAND3_X1 U7635 ( .A1(n7791), .A2(n5949), .A3(n7605), .ZN(n5998) );
  INV_X1 U7636 ( .A(n5998), .ZN(n5956) );
  AND2_X1 U7637 ( .A1(n9324), .A2(n7264), .ZN(n5991) );
  NOR2_X1 U7638 ( .A1(n7258), .A2(n5991), .ZN(n7565) );
  NAND2_X1 U7639 ( .A1(n5950), .A2(n5992), .ZN(n7461) );
  INV_X1 U7640 ( .A(n7461), .ZN(n7466) );
  NAND2_X1 U7641 ( .A1(n5951), .A2(n7464), .ZN(n7306) );
  INV_X1 U7642 ( .A(n7306), .ZN(n7308) );
  NAND4_X1 U7643 ( .A1(n7565), .A2(n7466), .A3(n7308), .A4(n7726), .ZN(n5952)
         );
  NAND2_X1 U7644 ( .A1(n5994), .A2(n6036), .ZN(n7504) );
  NOR2_X1 U7645 ( .A1(n5952), .A2(n7504), .ZN(n5955) );
  NAND4_X1 U7646 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(n5957)
         );
  NOR2_X1 U7647 ( .A1(n5957), .A2(n7869), .ZN(n5958) );
  NAND4_X1 U7648 ( .A1(n7991), .A2(n8225), .A3(n6037), .A4(n5958), .ZN(n5959)
         );
  NOR2_X1 U7649 ( .A1(n8127), .A2(n5959), .ZN(n5960) );
  NAND4_X1 U7650 ( .A1(n9634), .A2(n8204), .A3(n8129), .A4(n5960), .ZN(n5961)
         );
  NOR3_X1 U7651 ( .A1(n9594), .A2(n9607), .A3(n5961), .ZN(n5962) );
  NAND4_X1 U7652 ( .A1(n9551), .A2(n9567), .A3(n9581), .A4(n5962), .ZN(n5963)
         );
  NOR3_X1 U7653 ( .A1(n5964), .A2(n9507), .A3(n5963), .ZN(n5965) );
  NAND4_X1 U7654 ( .A1(n9453), .A2(n5966), .A3(n9487), .A4(n5965), .ZN(n5967)
         );
  NOR2_X1 U7655 ( .A1(n9437), .A2(n5967), .ZN(n5971) );
  INV_X1 U7656 ( .A(n9294), .ZN(n5968) );
  NOR2_X1 U7657 ( .A1(n9432), .A2(n5968), .ZN(n6063) );
  INV_X1 U7658 ( .A(n6063), .ZN(n5969) );
  NAND2_X1 U7659 ( .A1(n9432), .A2(n5968), .ZN(n5977) );
  AND2_X1 U7660 ( .A1(n5969), .A2(n5977), .ZN(n5970) );
  NAND4_X1 U7661 ( .A1(n6064), .A2(n8297), .A3(n5971), .A4(n5970), .ZN(n6068)
         );
  INV_X1 U7662 ( .A(n6068), .ZN(n5972) );
  NAND2_X1 U7663 ( .A1(n5972), .A2(n6074), .ZN(n5973) );
  AND2_X1 U7664 ( .A1(n5979), .A2(n5978), .ZN(n6022) );
  NAND2_X1 U7665 ( .A1(n8311), .A2(n5980), .ZN(n5981) );
  NAND2_X1 U7666 ( .A1(n5981), .A2(n5986), .ZN(n5982) );
  NAND2_X1 U7667 ( .A1(n8312), .A2(n5982), .ZN(n6019) );
  NAND2_X1 U7668 ( .A1(n5984), .A2(n5983), .ZN(n8307) );
  AND3_X1 U7669 ( .A1(n5986), .A2(n5985), .A3(n8307), .ZN(n5988) );
  OAI21_X1 U7670 ( .B1(n6019), .B2(n5988), .A(n5987), .ZN(n5990) );
  INV_X1 U7671 ( .A(n8314), .ZN(n5989) );
  AOI211_X1 U7672 ( .C1(n6022), .C2(n5990), .A(n5989), .B(n8315), .ZN(n6026)
         );
  NAND3_X1 U7673 ( .A1(n6027), .A2(n6026), .A3(n8313), .ZN(n6058) );
  INV_X1 U7674 ( .A(n6058), .ZN(n6032) );
  INV_X1 U7675 ( .A(n6056), .ZN(n6021) );
  OAI211_X1 U7676 ( .C1(n7304), .C2(n7650), .A(n6083), .B(n7464), .ZN(n5996)
         );
  INV_X1 U7677 ( .A(n5991), .ZN(n5993) );
  OAI211_X1 U7678 ( .C1(n4461), .C2(n10034), .A(n5993), .B(n5992), .ZN(n5995)
         );
  OAI21_X1 U7679 ( .B1(n5996), .B2(n5995), .A(n5994), .ZN(n5997) );
  OAI21_X1 U7680 ( .B1(n7505), .B2(n5997), .A(n6036), .ZN(n6003) );
  NAND2_X1 U7681 ( .A1(n5999), .A2(n5998), .ZN(n7877) );
  INV_X1 U7682 ( .A(n7877), .ZN(n6002) );
  INV_X1 U7683 ( .A(n6000), .ZN(n6001) );
  AOI211_X1 U7684 ( .C1(n6003), .C2(n6037), .A(n6002), .B(n6001), .ZN(n6005)
         );
  NOR2_X1 U7685 ( .A1(n6005), .A2(n6004), .ZN(n6008) );
  OAI211_X1 U7686 ( .C1(n6008), .C2(n6007), .A(n6045), .B(n6006), .ZN(n6010)
         );
  NAND3_X1 U7687 ( .A1(n6010), .A2(n8202), .A3(n6009), .ZN(n6012) );
  AOI21_X1 U7688 ( .B1(n6013), .B2(n6012), .A(n6011), .ZN(n6014) );
  OAI21_X1 U7689 ( .B1(n6015), .B2(n6014), .A(n6053), .ZN(n6017) );
  AOI21_X1 U7690 ( .B1(n6018), .B2(n6017), .A(n6016), .ZN(n6020) );
  NOR2_X1 U7691 ( .A1(n6019), .A2(n8306), .ZN(n6060) );
  OAI21_X1 U7692 ( .B1(n6021), .B2(n6020), .A(n6060), .ZN(n6031) );
  INV_X1 U7693 ( .A(n6022), .ZN(n6025) );
  INV_X1 U7694 ( .A(n6023), .ZN(n6024) );
  AOI21_X1 U7695 ( .B1(n6026), .B2(n6025), .A(n6024), .ZN(n6030) );
  INV_X1 U7696 ( .A(n6027), .ZN(n6028) );
  AOI21_X1 U7697 ( .B1(n6030), .B2(n6029), .A(n6028), .ZN(n6062) );
  INV_X1 U7698 ( .A(n6064), .ZN(n6076) );
  OAI21_X1 U7699 ( .B1(n6033), .B2(n6076), .A(n6074), .ZN(n6072) );
  NAND2_X1 U7700 ( .A1(n6035), .A2(n6034), .ZN(n6071) );
  NAND2_X1 U7701 ( .A1(n7632), .A2(n6036), .ZN(n7613) );
  NAND2_X1 U7702 ( .A1(n7613), .A2(n6037), .ZN(n7878) );
  INV_X1 U7703 ( .A(n8226), .ZN(n6039) );
  NOR2_X1 U7704 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NAND2_X1 U7705 ( .A1(n8227), .A2(n6041), .ZN(n8224) );
  NAND2_X1 U7706 ( .A1(n8224), .A2(n6042), .ZN(n7990) );
  NAND2_X1 U7707 ( .A1(n7990), .A2(n7991), .ZN(n8095) );
  INV_X1 U7708 ( .A(n8094), .ZN(n6043) );
  NOR2_X1 U7709 ( .A1(n8127), .A2(n6043), .ZN(n6044) );
  NOR2_X1 U7710 ( .A1(n6047), .A2(n6046), .ZN(n6048) );
  NAND2_X1 U7711 ( .A1(n6050), .A2(n6049), .ZN(n9635) );
  NAND2_X1 U7712 ( .A1(n6055), .A2(n6054), .ZN(n9578) );
  NAND2_X1 U7713 ( .A1(n9578), .A2(n9581), .ZN(n6057) );
  INV_X1 U7714 ( .A(n9568), .ZN(n6059) );
  AOI21_X1 U7715 ( .B1(n6060), .B2(n6059), .A(n6058), .ZN(n6061) );
  AOI211_X1 U7716 ( .C1(n6063), .C2(n6891), .A(n6062), .B(n6061), .ZN(n6066)
         );
  OAI21_X1 U7717 ( .B1(n4472), .B2(n6891), .A(n6064), .ZN(n6065) );
  OAI21_X1 U7718 ( .B1(n6066), .B2(n6065), .A(n6810), .ZN(n6069) );
  AOI211_X1 U7719 ( .C1(n6069), .C2(n6068), .A(n6067), .B(n7624), .ZN(n6070)
         );
  OAI21_X1 U7720 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(n6078) );
  NAND2_X1 U7721 ( .A1(n6083), .A2(n6758), .ZN(n6970) );
  AOI211_X1 U7722 ( .C1(n6076), .C2(n7570), .A(n6969), .B(n6970), .ZN(n6077)
         );
  OR2_X1 U7723 ( .A1(n6809), .A2(P1_U3086), .ZN(n6771) );
  NAND2_X1 U7724 ( .A1(n6083), .A2(n7624), .ZN(n6525) );
  OR2_X1 U7725 ( .A1(n6967), .A2(n6525), .ZN(n7562) );
  INV_X1 U7726 ( .A(n6813), .ZN(n9783) );
  INV_X1 U7727 ( .A(n8217), .ZN(n6805) );
  NAND2_X1 U7728 ( .A1(n6805), .A2(n6084), .ZN(n6827) );
  NOR3_X1 U7729 ( .A1(n7562), .A2(n9783), .A3(n6827), .ZN(n6086) );
  OAI21_X1 U7730 ( .B1(n6771), .B2(n6969), .A(P1_B_REG_SCAN_IN), .ZN(n6085) );
  INV_X1 U7731 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6090) );
  XNOR2_X2 U7732 ( .A(n6089), .B(P2_IR_REG_30__SCAN_IN), .ZN(n6093) );
  NAND2_X1 U7733 ( .A1(n6093), .A2(n8219), .ZN(n6131) );
  INV_X1 U7734 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7296) );
  OR2_X1 U7735 ( .A1(n6131), .A2(n7296), .ZN(n6098) );
  NAND2_X2 U7736 ( .A1(n6094), .A2(n8219), .ZN(n6145) );
  OR2_X1 U7737 ( .A1(n6145), .A2(n10225), .ZN(n6097) );
  NAND2_X1 U7738 ( .A1(n6094), .A2(n6092), .ZN(n6133) );
  INV_X1 U7739 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n6095) );
  OR2_X1 U7740 ( .A1(n6133), .A2(n6095), .ZN(n6096) );
  INV_X1 U7741 ( .A(n10154), .ZN(n6107) );
  NAND2_X1 U7742 ( .A1(n6139), .A2(n6848), .ZN(n6105) );
  INV_X1 U7743 ( .A(n7425), .ZN(n6101) );
  OR2_X1 U7744 ( .A1(n6102), .A2(n6101), .ZN(n6103) );
  NAND2_X1 U7745 ( .A1(n6107), .A2(n6106), .ZN(n8330) );
  INV_X1 U7746 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6109) );
  OR2_X1 U7747 ( .A1(n6133), .A2(n6109), .ZN(n6114) );
  NAND2_X1 U7748 ( .A1(n6110), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6113) );
  INV_X1 U7749 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6111) );
  NAND4_X1 U7750 ( .A1(n6115), .A2(n6114), .A3(n6113), .A4(n6112), .ZN(n8708)
         );
  INV_X1 U7751 ( .A(SI_0_), .ZN(n6117) );
  INV_X1 U7752 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7753 ( .B1(n6846), .B2(n6117), .A(n6116), .ZN(n6119) );
  NAND2_X1 U7754 ( .A1(n6119), .A2(n6118), .ZN(n6841) );
  MUX2_X1 U7755 ( .A(n10089), .B(n6841), .S(n6445), .Z(n7214) );
  NAND2_X1 U7756 ( .A1(n8708), .A2(n6451), .ZN(n7350) );
  NAND2_X1 U7757 ( .A1(n7345), .A2(n7350), .ZN(n6121) );
  NAND2_X1 U7758 ( .A1(n10154), .A2(n6106), .ZN(n6120) );
  NAND2_X1 U7759 ( .A1(n6121), .A2(n6120), .ZN(n10151) );
  NAND2_X1 U7760 ( .A1(n6139), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6122) );
  INV_X1 U7761 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n6124) );
  OR2_X1 U7762 ( .A1(n6133), .A2(n6124), .ZN(n6128) );
  INV_X2 U7763 ( .A(n6145), .ZN(n8452) );
  INV_X1 U7764 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10148) );
  OR2_X1 U7765 ( .A1(n6131), .A2(n10148), .ZN(n6125) );
  NAND2_X1 U7766 ( .A1(n6129), .A2(n7225), .ZN(n6130) );
  NAND2_X1 U7767 ( .A1(n8452), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6138) );
  OR2_X1 U7768 ( .A1(n6310), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n6137) );
  INV_X1 U7769 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6132) );
  OR2_X1 U7770 ( .A1(n6149), .A2(n6132), .ZN(n6136) );
  INV_X1 U7771 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6134) );
  OR2_X1 U7772 ( .A1(n6442), .A2(n6134), .ZN(n6135) );
  NAND2_X1 U7773 ( .A1(n6139), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7774 ( .A1(n6318), .A2(n6140), .ZN(n6141) );
  NAND2_X1 U7775 ( .A1(n8453), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n6153) );
  OR2_X1 U7776 ( .A1(n6145), .A2(n6146), .ZN(n6152) );
  NAND2_X1 U7777 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6148) );
  AND2_X1 U7778 ( .A1(n6159), .A2(n6148), .ZN(n7341) );
  OR2_X1 U7779 ( .A1(n6310), .A2(n7341), .ZN(n6151) );
  OR2_X1 U7780 ( .A1(n6149), .A2(n7494), .ZN(n6150) );
  NAND2_X1 U7781 ( .A1(n8450), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6155) );
  NAND2_X1 U7782 ( .A1(n6318), .A2(n7400), .ZN(n6154) );
  OAI211_X1 U7783 ( .C1(n6215), .C2(n6853), .A(n6155), .B(n6154), .ZN(n10177)
         );
  NAND2_X1 U7784 ( .A1(n8453), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n6164) );
  OR2_X1 U7785 ( .A1(n6145), .A2(n6156), .ZN(n6163) );
  NAND2_X1 U7786 ( .A1(n6159), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6160) );
  AND2_X1 U7787 ( .A1(n6169), .A2(n6160), .ZN(n7486) );
  OR2_X1 U7788 ( .A1(n6310), .A2(n7486), .ZN(n6162) );
  OR2_X1 U7789 ( .A1(n6149), .A2(n5479), .ZN(n6161) );
  NAND4_X1 U7790 ( .A1(n6164), .A2(n6163), .A3(n6162), .A4(n6161), .ZN(n8707)
         );
  NAND2_X1 U7791 ( .A1(n8450), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U7792 ( .A1(n6318), .A2(n6165), .ZN(n6166) );
  OAI211_X1 U7793 ( .C1(n6215), .C2(n6855), .A(n6167), .B(n6166), .ZN(n7451)
         );
  OR2_X1 U7794 ( .A1(n8707), .A2(n7451), .ZN(n7478) );
  NAND2_X1 U7795 ( .A1(n8707), .A2(n7451), .ZN(n7477) );
  NAND2_X1 U7796 ( .A1(n8452), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6175) );
  INV_X1 U7797 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n6168) );
  OR2_X1 U7798 ( .A1(n6442), .A2(n6168), .ZN(n6174) );
  NAND2_X1 U7799 ( .A1(n6169), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6170) );
  AND2_X1 U7800 ( .A1(n6184), .A2(n6170), .ZN(n7703) );
  OR2_X1 U7801 ( .A1(n6310), .A2(n7703), .ZN(n6173) );
  INV_X1 U7802 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6171) );
  OR2_X1 U7803 ( .A1(n6149), .A2(n6171), .ZN(n6172) );
  NAND2_X1 U7804 ( .A1(n8450), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n6178) );
  NAND2_X1 U7805 ( .A1(n6318), .A2(n6176), .ZN(n6177) );
  OAI211_X1 U7806 ( .C1(n6215), .C2(n6862), .A(n6178), .B(n6177), .ZN(n7526)
         );
  AND2_X1 U7807 ( .A1(n8706), .A2(n7526), .ZN(n6180) );
  INV_X1 U7808 ( .A(n8706), .ZN(n7676) );
  INV_X1 U7809 ( .A(n7526), .ZN(n10184) );
  NAND2_X1 U7810 ( .A1(n7676), .A2(n10184), .ZN(n6179) );
  NAND2_X1 U7811 ( .A1(n8452), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6189) );
  INV_X1 U7812 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6181) );
  OR2_X1 U7813 ( .A1(n6442), .A2(n6181), .ZN(n6188) );
  NAND2_X1 U7814 ( .A1(n6184), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n6185) );
  AND2_X1 U7815 ( .A1(n6198), .A2(n6185), .ZN(n7735) );
  OR2_X1 U7816 ( .A1(n6310), .A2(n7735), .ZN(n6187) );
  OR2_X1 U7817 ( .A1(n6149), .A2(n7546), .ZN(n6186) );
  NAND4_X1 U7818 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(n8704)
         );
  NAND2_X1 U7819 ( .A1(n6864), .A2(n8451), .ZN(n6191) );
  NAND2_X1 U7820 ( .A1(n8450), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n6190) );
  OAI211_X1 U7821 ( .C1(n6445), .C2(n6866), .A(n6191), .B(n6190), .ZN(n7737)
         );
  INV_X1 U7822 ( .A(n7737), .ZN(n10188) );
  OR2_X1 U7823 ( .A1(n8704), .A2(n10188), .ZN(n8350) );
  NAND2_X1 U7824 ( .A1(n8704), .A2(n10188), .ZN(n7685) );
  NAND2_X1 U7825 ( .A1(n7730), .A2(n8483), .ZN(n6193) );
  INV_X1 U7826 ( .A(n8704), .ZN(n7769) );
  NAND2_X1 U7827 ( .A1(n7769), .A2(n10188), .ZN(n6192) );
  NAND2_X1 U7828 ( .A1(n6868), .A2(n8451), .ZN(n6196) );
  AOI22_X1 U7829 ( .A1(n8450), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6318), .B2(
        n6194), .ZN(n6195) );
  NAND2_X1 U7830 ( .A1(n8453), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7831 ( .A1(n6145), .A2(n6197), .ZN(n6202) );
  NAND2_X1 U7832 ( .A1(n6198), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6199) );
  AND2_X1 U7833 ( .A1(n6207), .A2(n6199), .ZN(n7775) );
  OR2_X1 U7834 ( .A1(n6310), .A2(n7775), .ZN(n6201) );
  OR2_X1 U7835 ( .A1(n6149), .A2(n7687), .ZN(n6200) );
  NAND2_X1 U7836 ( .A1(n7776), .A2(n7774), .ZN(n8353) );
  NAND2_X1 U7837 ( .A1(n8352), .A2(n8353), .ZN(n8481) );
  INV_X1 U7838 ( .A(n8481), .ZN(n7681) );
  OR2_X1 U7839 ( .A1(n7774), .A2(n10193), .ZN(n6204) );
  NAND2_X1 U7840 ( .A1(n8453), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6212) );
  OR2_X1 U7841 ( .A1(n6145), .A2(n10237), .ZN(n6211) );
  INV_X1 U7842 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n6205) );
  NAND2_X1 U7843 ( .A1(n6207), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6208) );
  AND2_X1 U7844 ( .A1(n6220), .A2(n6208), .ZN(n7857) );
  OR2_X1 U7845 ( .A1(n6310), .A2(n7857), .ZN(n6210) );
  OR2_X1 U7846 ( .A1(n6149), .A2(n7825), .ZN(n6209) );
  INV_X2 U7847 ( .A(n6215), .ZN(n8451) );
  NAND2_X1 U7848 ( .A1(n6872), .A2(n8451), .ZN(n6214) );
  AOI22_X1 U7849 ( .A1(n8450), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6318), .B2(
        n7828), .ZN(n6213) );
  NAND2_X1 U7850 ( .A1(n6883), .A2(n8451), .ZN(n6218) );
  AOI22_X1 U7851 ( .A1(n8450), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6318), .B2(
        n6216), .ZN(n6217) );
  NAND2_X1 U7852 ( .A1(n8453), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6225) );
  OR2_X1 U7853 ( .A1(n6145), .A2(n6219), .ZN(n6224) );
  NAND2_X1 U7854 ( .A1(n6220), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6221) );
  AND2_X1 U7855 ( .A1(n6232), .A2(n6221), .ZN(n8032) );
  OR2_X1 U7856 ( .A1(n6310), .A2(n8032), .ZN(n6223) );
  OR2_X1 U7857 ( .A1(n6149), .A2(n5489), .ZN(n6222) );
  NAND2_X1 U7858 ( .A1(n8076), .A2(n8068), .ZN(n6226) );
  NAND2_X1 U7859 ( .A1(n7962), .A2(n6226), .ZN(n6228) );
  OR2_X1 U7860 ( .A1(n8076), .A2(n8068), .ZN(n6227) );
  NAND2_X1 U7861 ( .A1(n6887), .A2(n8451), .ZN(n6230) );
  AOI22_X1 U7862 ( .A1(n8450), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6318), .B2(
        n8714), .ZN(n6229) );
  NAND2_X1 U7863 ( .A1(n6230), .A2(n6229), .ZN(n8057) );
  NAND2_X1 U7864 ( .A1(n8452), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6237) );
  INV_X1 U7865 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n6231) );
  OR2_X1 U7866 ( .A1(n6442), .A2(n6231), .ZN(n6236) );
  NAND2_X1 U7867 ( .A1(n6232), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6233) );
  AND2_X1 U7868 ( .A1(n6244), .A2(n6233), .ZN(n8054) );
  OR2_X1 U7869 ( .A1(n6310), .A2(n8054), .ZN(n6235) );
  OR2_X1 U7870 ( .A1(n6149), .A2(n8711), .ZN(n6234) );
  NAND2_X1 U7871 ( .A1(n8057), .A2(n8174), .ZN(n8382) );
  NAND2_X1 U7872 ( .A1(n8381), .A2(n8382), .ZN(n8074) );
  INV_X1 U7873 ( .A(n8174), .ZN(n8701) );
  NAND2_X1 U7874 ( .A1(n8057), .A2(n8701), .ZN(n6238) );
  NAND2_X1 U7875 ( .A1(n6889), .A2(n8451), .ZN(n6241) );
  OAI22_X1 U7876 ( .A1(n6265), .A2(n6893), .B1(n8015), .B2(n6445), .ZN(n6239)
         );
  INV_X1 U7877 ( .A(n6239), .ZN(n6240) );
  NAND2_X1 U7878 ( .A1(n8453), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6249) );
  OR2_X1 U7879 ( .A1(n6145), .A2(n6242), .ZN(n6248) );
  OR2_X1 U7880 ( .A1(n6149), .A2(n8042), .ZN(n6247) );
  INV_X1 U7881 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8014) );
  NAND2_X1 U7882 ( .A1(n6244), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6245) );
  AND2_X1 U7883 ( .A1(n6257), .A2(n6245), .ZN(n8179) );
  OR2_X1 U7884 ( .A1(n6310), .A2(n8179), .ZN(n6246) );
  NAND4_X1 U7885 ( .A1(n6249), .A2(n6248), .A3(n6247), .A4(n6246), .ZN(n8700)
         );
  OR2_X1 U7886 ( .A1(n10220), .A2(n8700), .ZN(n6250) );
  NAND2_X1 U7887 ( .A1(n10220), .A2(n8700), .ZN(n6251) );
  NAND2_X1 U7888 ( .A1(n6252), .A2(n6251), .ZN(n8118) );
  NAND2_X1 U7889 ( .A1(n6954), .A2(n8451), .ZN(n6254) );
  AOI22_X1 U7890 ( .A1(n8450), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6318), .B2(
        n10091), .ZN(n6253) );
  NAND2_X1 U7891 ( .A1(n8453), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6262) );
  OR2_X1 U7892 ( .A1(n6145), .A2(n10101), .ZN(n6261) );
  INV_X1 U7893 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7894 ( .A1(n6257), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6258) );
  AND2_X1 U7895 ( .A1(n6267), .A2(n6258), .ZN(n8122) );
  OR2_X1 U7896 ( .A1(n6310), .A2(n8122), .ZN(n6260) );
  OR2_X1 U7897 ( .A1(n6149), .A2(n10094), .ZN(n6259) );
  NAND4_X1 U7898 ( .A1(n6262), .A2(n6261), .A3(n6260), .A4(n6259), .ZN(n8977)
         );
  NAND2_X1 U7899 ( .A1(n9143), .A2(n8182), .ZN(n8391) );
  NAND2_X1 U7900 ( .A1(n8118), .A2(n8489), .ZN(n6264) );
  NAND2_X1 U7901 ( .A1(n9143), .A2(n8977), .ZN(n6263) );
  INV_X1 U7902 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6963) );
  OAI22_X1 U7903 ( .A1(n10127), .A2(n6445), .B1(n6265), .B2(n6963), .ZN(n6266)
         );
  NAND2_X1 U7904 ( .A1(n8453), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6272) );
  OR2_X1 U7905 ( .A1(n6145), .A2(n9045), .ZN(n6271) );
  NAND2_X1 U7906 ( .A1(n6267), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6268) );
  AND2_X1 U7907 ( .A1(n6279), .A2(n6268), .ZN(n8980) );
  OR2_X1 U7908 ( .A1(n6310), .A2(n8980), .ZN(n6270) );
  OR2_X1 U7909 ( .A1(n6149), .A2(n8991), .ZN(n6269) );
  NAND4_X1 U7910 ( .A1(n6272), .A2(n6271), .A3(n6270), .A4(n6269), .ZN(n8518)
         );
  OR2_X1 U7911 ( .A1(n8982), .A2(n8518), .ZN(n8398) );
  NAND2_X1 U7912 ( .A1(n8982), .A2(n8518), .ZN(n8397) );
  NAND2_X1 U7913 ( .A1(n8398), .A2(n8397), .ZN(n8986) );
  NAND2_X1 U7914 ( .A1(n8976), .A2(n8986), .ZN(n6274) );
  INV_X1 U7915 ( .A(n8518), .ZN(n8680) );
  OR2_X1 U7916 ( .A1(n8982), .A2(n8680), .ZN(n6273) );
  NAND2_X1 U7917 ( .A1(n6976), .A2(n8451), .ZN(n6276) );
  AOI22_X1 U7918 ( .A1(n6977), .A2(n6318), .B1(n8450), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U7919 ( .A1(n8453), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6284) );
  OR2_X1 U7920 ( .A1(n6145), .A2(n8249), .ZN(n6283) );
  INV_X1 U7921 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7922 ( .A1(n6279), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6280) );
  AND2_X1 U7923 ( .A1(n6288), .A2(n6280), .ZN(n8686) );
  OR2_X1 U7924 ( .A1(n6310), .A2(n8686), .ZN(n6282) );
  OR2_X1 U7925 ( .A1(n6149), .A2(n8728), .ZN(n6281) );
  NAND4_X1 U7926 ( .A1(n6284), .A2(n6283), .A3(n6282), .A4(n6281), .ZN(n8978)
         );
  INV_X1 U7927 ( .A(n8978), .ZN(n8616) );
  OR2_X1 U7928 ( .A1(n8694), .A2(n8616), .ZN(n8401) );
  NAND2_X1 U7929 ( .A1(n8694), .A2(n8616), .ZN(n6458) );
  NAND2_X1 U7930 ( .A1(n8244), .A2(n8242), .ZN(n6286) );
  NAND2_X1 U7931 ( .A1(n8694), .A2(n8978), .ZN(n6285) );
  NAND2_X1 U7932 ( .A1(n6286), .A2(n6285), .ZN(n8967) );
  AOI22_X1 U7933 ( .A1(n8450), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6318), .B2(
        n7198), .ZN(n6287) );
  NAND2_X1 U7934 ( .A1(n8452), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6293) );
  INV_X1 U7935 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9129) );
  OR2_X1 U7936 ( .A1(n6442), .A2(n9129), .ZN(n6292) );
  NAND2_X1 U7937 ( .A1(n6288), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6289) );
  AND2_X1 U7938 ( .A1(n6301), .A2(n6289), .ZN(n8972) );
  OR2_X1 U7939 ( .A1(n6310), .A2(n8972), .ZN(n6291) );
  INV_X1 U7940 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8971) );
  OR2_X1 U7941 ( .A1(n6149), .A2(n8971), .ZN(n6290) );
  NAND4_X1 U7942 ( .A1(n6293), .A2(n6292), .A3(n6291), .A4(n6290), .ZN(n8699)
         );
  NAND2_X1 U7943 ( .A1(n9130), .A2(n8960), .ZN(n8406) );
  INV_X1 U7944 ( .A(n8968), .ZN(n6294) );
  NAND2_X1 U7945 ( .A1(n8967), .A2(n6294), .ZN(n6296) );
  NAND2_X1 U7946 ( .A1(n9130), .A2(n8699), .ZN(n6295) );
  NAND2_X1 U7947 ( .A1(n6296), .A2(n6295), .ZN(n8957) );
  NAND2_X1 U7948 ( .A1(n7326), .A2(n8451), .ZN(n6298) );
  AOI22_X1 U7949 ( .A1(n8450), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6318), .B2(
        n8768), .ZN(n6297) );
  INV_X1 U7950 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7951 ( .A1(n6301), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6302) );
  AND2_X1 U7952 ( .A1(n6311), .A2(n6302), .ZN(n8961) );
  OR2_X1 U7953 ( .A1(n6310), .A2(n8961), .ZN(n6306) );
  INV_X1 U7954 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9125) );
  OR2_X1 U7955 ( .A1(n6442), .A2(n9125), .ZN(n6305) );
  OR2_X1 U7956 ( .A1(n6145), .A2(n9040), .ZN(n6304) );
  OR2_X1 U7957 ( .A1(n6149), .A2(n8962), .ZN(n6303) );
  NAND4_X1 U7958 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n8969)
         );
  INV_X1 U7959 ( .A(n8969), .ZN(n8942) );
  OR2_X1 U7960 ( .A1(n9039), .A2(n8942), .ZN(n8407) );
  NAND2_X1 U7961 ( .A1(n9039), .A2(n8942), .ZN(n8410) );
  NAND2_X1 U7962 ( .A1(n9039), .A2(n8969), .ZN(n6307) );
  NAND2_X1 U7963 ( .A1(n7454), .A2(n8451), .ZN(n6309) );
  AOI22_X1 U7964 ( .A1(n6318), .A2(n8798), .B1(n8450), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U7965 ( .A1(n6311), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7966 ( .A1(n6325), .A2(n6312), .ZN(n8947) );
  NAND2_X1 U7967 ( .A1(n6110), .A2(n8947), .ZN(n6317) );
  INV_X1 U7968 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9035) );
  OR2_X1 U7969 ( .A1(n6145), .A2(n9035), .ZN(n6316) );
  INV_X1 U7970 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9120) );
  OR2_X1 U7971 ( .A1(n6442), .A2(n9120), .ZN(n6315) );
  OR2_X1 U7972 ( .A1(n6149), .A2(n6313), .ZN(n6314) );
  NAND4_X1 U7973 ( .A1(n6317), .A2(n6316), .A3(n6315), .A4(n6314), .ZN(n8926)
         );
  NAND2_X1 U7974 ( .A1(n8657), .A2(n8959), .ZN(n8411) );
  NAND2_X1 U7975 ( .A1(n8924), .A2(n8411), .ZN(n8944) );
  INV_X1 U7976 ( .A(n8944), .ZN(n8940) );
  NAND2_X1 U7977 ( .A1(n7516), .A2(n8451), .ZN(n6320) );
  AOI22_X1 U7978 ( .A1(n8509), .A2(n6318), .B1(n8450), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7979 ( .A1(n8453), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6322) );
  NAND2_X1 U7980 ( .A1(n8452), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6321) );
  AND2_X1 U7981 ( .A1(n6322), .A2(n6321), .ZN(n6329) );
  INV_X1 U7982 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7983 ( .A1(n6325), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6326) );
  NAND2_X1 U7984 ( .A1(n6333), .A2(n6326), .ZN(n8934) );
  NAND2_X1 U7985 ( .A1(n8934), .A2(n6110), .ZN(n6328) );
  OR2_X1 U7986 ( .A1(n6149), .A2(n5530), .ZN(n6327) );
  OR2_X1 U7987 ( .A1(n9115), .A2(n8943), .ZN(n8409) );
  NAND2_X1 U7988 ( .A1(n9115), .A2(n8943), .ZN(n8415) );
  NAND2_X1 U7989 ( .A1(n8409), .A2(n8415), .ZN(n8927) );
  OR2_X1 U7990 ( .A1(n8657), .A2(n8926), .ZN(n8928) );
  AND2_X1 U7991 ( .A1(n8927), .A2(n8928), .ZN(n6330) );
  NAND2_X1 U7992 ( .A1(n7600), .A2(n8451), .ZN(n6332) );
  NAND2_X1 U7993 ( .A1(n8450), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6331) );
  INV_X1 U7994 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8920) );
  NAND2_X1 U7995 ( .A1(n6333), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U7996 ( .A1(n6342), .A2(n6334), .ZN(n8921) );
  NAND2_X1 U7997 ( .A1(n8921), .A2(n6110), .ZN(n6336) );
  AOI22_X1 U7998 ( .A1(n8453), .A2(P2_REG0_REG_20__SCAN_IN), .B1(n8452), .B2(
        P2_REG1_REG_20__SCAN_IN), .ZN(n6335) );
  OAI211_X1 U7999 ( .C1(n6149), .C2(n8920), .A(n6336), .B(n6335), .ZN(n8933)
         );
  INV_X1 U8000 ( .A(n8933), .ZN(n8601) );
  OR2_X1 U8001 ( .A1(n9109), .A2(n8601), .ZN(n8896) );
  NAND2_X1 U8002 ( .A1(n9109), .A2(n8601), .ZN(n8897) );
  INV_X1 U8003 ( .A(n8943), .ZN(n8918) );
  AND2_X1 U8004 ( .A1(n9115), .A2(n8918), .ZN(n8915) );
  NOR2_X1 U8005 ( .A1(n8914), .A2(n8915), .ZN(n6337) );
  OR2_X1 U8006 ( .A1(n9109), .A2(n8933), .ZN(n8902) );
  NAND2_X1 U8007 ( .A1(n8900), .A2(n8902), .ZN(n6347) );
  NAND2_X1 U8008 ( .A1(n7710), .A2(n8451), .ZN(n6339) );
  NAND2_X1 U8009 ( .A1(n8450), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6338) );
  INV_X1 U8010 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8907) );
  INV_X1 U8011 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n6340) );
  NAND2_X1 U8012 ( .A1(n6342), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6343) );
  NAND2_X1 U8013 ( .A1(n6350), .A2(n6343), .ZN(n8908) );
  NAND2_X1 U8014 ( .A1(n8908), .A2(n6110), .ZN(n6345) );
  AOI22_X1 U8015 ( .A1(n8453), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n8452), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6344) );
  OAI211_X1 U8016 ( .C1(n6149), .C2(n8907), .A(n6345), .B(n6344), .ZN(n8917)
         );
  INV_X1 U8017 ( .A(n8917), .ZN(n6346) );
  NAND2_X1 U8018 ( .A1(n9103), .A2(n6346), .ZN(n8421) );
  NAND2_X1 U8019 ( .A1(n8420), .A2(n8421), .ZN(n8901) );
  NAND2_X1 U8020 ( .A1(n6347), .A2(n8901), .ZN(n8883) );
  OR2_X1 U8021 ( .A1(n9103), .A2(n8917), .ZN(n8884) );
  NAND2_X1 U8022 ( .A1(n8883), .A2(n8884), .ZN(n6358) );
  NAND2_X1 U8023 ( .A1(n7809), .A2(n8451), .ZN(n6349) );
  NAND2_X1 U8024 ( .A1(n8450), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U8025 ( .A1(n6350), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U8026 ( .A1(n6362), .A2(n6351), .ZN(n8890) );
  NAND2_X1 U8027 ( .A1(n8890), .A2(n6110), .ZN(n6356) );
  INV_X1 U8028 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U8029 ( .A1(n8453), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6353) );
  NAND2_X1 U8030 ( .A1(n8452), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6352) );
  OAI211_X1 U8031 ( .C1(n8892), .C2(n6149), .A(n6353), .B(n6352), .ZN(n6354)
         );
  INV_X1 U8032 ( .A(n6354), .ZN(n6355) );
  INV_X1 U8033 ( .A(n8905), .ZN(n6357) );
  NOR2_X1 U8034 ( .A1(n9019), .A2(n6357), .ZN(n8323) );
  INV_X1 U8035 ( .A(n8323), .ZN(n6460) );
  NAND2_X1 U8036 ( .A1(n9019), .A2(n6357), .ZN(n8322) );
  OR2_X1 U8037 ( .A1(n9019), .A2(n8905), .ZN(n6359) );
  NAND2_X1 U8038 ( .A1(n7956), .A2(n8451), .ZN(n6361) );
  NAND2_X1 U8039 ( .A1(n8450), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6360) );
  NAND2_X1 U8040 ( .A1(n6362), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6363) );
  NAND2_X1 U8041 ( .A1(n6375), .A2(n6363), .ZN(n8879) );
  NAND2_X1 U8042 ( .A1(n8879), .A2(n6110), .ZN(n6368) );
  INV_X1 U8043 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U8044 ( .A1(n8452), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6365) );
  OAI211_X1 U8045 ( .C1(n6442), .C2(n9095), .A(n6365), .B(n6364), .ZN(n6366)
         );
  INV_X1 U8046 ( .A(n6366), .ZN(n6367) );
  NAND2_X1 U8047 ( .A1(n9096), .A2(n8888), .ZN(n6369) );
  OR2_X1 U8048 ( .A1(n9096), .A2(n8888), .ZN(n6370) );
  INV_X1 U8049 ( .A(n8862), .ZN(n6382) );
  NAND2_X1 U8050 ( .A1(n7979), .A2(n8451), .ZN(n6372) );
  NAND2_X1 U8051 ( .A1(n8450), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6371) );
  INV_X1 U8052 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U8053 ( .A1(n6375), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U8054 ( .A1(n6387), .A2(n6376), .ZN(n8867) );
  NAND2_X1 U8055 ( .A1(n8867), .A2(n6110), .ZN(n6381) );
  INV_X1 U8056 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9089) );
  NAND2_X1 U8057 ( .A1(n8452), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6377) );
  OAI211_X1 U8058 ( .C1(n6442), .C2(n9089), .A(n6378), .B(n6377), .ZN(n6379)
         );
  INV_X1 U8059 ( .A(n6379), .ZN(n6380) );
  NAND2_X1 U8060 ( .A1(n9090), .A2(n8877), .ZN(n8850) );
  NAND2_X1 U8061 ( .A1(n7999), .A2(n8451), .ZN(n6384) );
  NAND2_X1 U8062 ( .A1(n8450), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6383) );
  INV_X1 U8063 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6385) );
  NAND2_X1 U8064 ( .A1(n6387), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6388) );
  NAND2_X1 U8065 ( .A1(n6397), .A2(n6388), .ZN(n8857) );
  NAND2_X1 U8066 ( .A1(n8857), .A2(n6110), .ZN(n6393) );
  INV_X1 U8067 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n9082) );
  NAND2_X1 U8068 ( .A1(n8452), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6390) );
  OAI211_X1 U8069 ( .C1(n9082), .C2(n6442), .A(n6390), .B(n6389), .ZN(n6391)
         );
  INV_X1 U8070 ( .A(n6391), .ZN(n6392) );
  NAND2_X1 U8071 ( .A1(n9083), .A2(n8844), .ZN(n8429) );
  AND2_X1 U8072 ( .A1(n8850), .A2(n8429), .ZN(n6394) );
  OR2_X1 U8073 ( .A1(n9083), .A2(n8844), .ZN(n8430) );
  NAND2_X1 U8074 ( .A1(n8064), .A2(n8451), .ZN(n6396) );
  NAND2_X1 U8075 ( .A1(n8450), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U8076 ( .A1(n6397), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8077 ( .A1(n6409), .A2(n6398), .ZN(n8847) );
  NAND2_X1 U8078 ( .A1(n8847), .A2(n6110), .ZN(n6403) );
  INV_X1 U8079 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9005) );
  NAND2_X1 U8080 ( .A1(n8453), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6400) );
  OAI211_X1 U8081 ( .C1(n6145), .C2(n9005), .A(n6400), .B(n6399), .ZN(n6401)
         );
  INV_X1 U8082 ( .A(n6401), .ZN(n6402) );
  NAND2_X1 U8083 ( .A1(n8145), .A2(n8451), .ZN(n6406) );
  NAND2_X1 U8084 ( .A1(n8450), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6405) );
  INV_X1 U8085 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6407) );
  NAND2_X1 U8086 ( .A1(n6409), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6410) );
  NAND2_X1 U8087 ( .A1(n6418), .A2(n6410), .ZN(n8838) );
  NAND2_X1 U8088 ( .A1(n8838), .A2(n6110), .ZN(n6415) );
  INV_X1 U8089 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n9069) );
  NAND2_X1 U8090 ( .A1(n8452), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6412) );
  OAI211_X1 U8091 ( .C1(n9069), .C2(n6442), .A(n6412), .B(n6411), .ZN(n6413)
         );
  INV_X1 U8092 ( .A(n6413), .ZN(n6414) );
  NAND2_X2 U8093 ( .A1(n6415), .A2(n6414), .ZN(n8845) );
  NAND2_X1 U8094 ( .A1(n9076), .A2(n8698), .ZN(n8832) );
  NAND2_X1 U8095 ( .A1(n8450), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6416) );
  NAND2_X1 U8096 ( .A1(n6418), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6419) );
  NAND2_X1 U8097 ( .A1(n8807), .A2(n6419), .ZN(n8827) );
  NAND2_X1 U8098 ( .A1(n8827), .A2(n6110), .ZN(n6424) );
  INV_X1 U8099 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n9063) );
  NAND2_X1 U8100 ( .A1(n8452), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6420) );
  OAI211_X1 U8101 ( .C1(n6442), .C2(n9063), .A(n6421), .B(n6420), .ZN(n6422)
         );
  INV_X1 U8102 ( .A(n6422), .ZN(n6423) );
  NOR2_X1 U8103 ( .A1(n9064), .A2(n8697), .ZN(n6425) );
  INV_X1 U8104 ( .A(n9064), .ZN(n8998) );
  OAI22_X1 U8105 ( .A1(n8823), .A2(n6425), .B1(n8837), .B2(n8998), .ZN(n6433)
         );
  NAND2_X1 U8106 ( .A1(n8218), .A2(n8451), .ZN(n6427) );
  NAND2_X1 U8107 ( .A1(n8450), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6426) );
  NAND2_X1 U8108 ( .A1(n6427), .A2(n6426), .ZN(n6504) );
  INV_X1 U8109 ( .A(n8807), .ZN(n6428) );
  NAND2_X1 U8110 ( .A1(n6428), .A2(n6110), .ZN(n8455) );
  INV_X1 U8111 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6518) );
  NAND2_X1 U8112 ( .A1(n8452), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6430) );
  OAI211_X1 U8113 ( .C1(n6518), .C2(n6442), .A(n6430), .B(n6429), .ZN(n6431)
         );
  INV_X1 U8114 ( .A(n6431), .ZN(n6432) );
  NAND2_X1 U8115 ( .A1(n6504), .A2(n8825), .ZN(n8446) );
  XNOR2_X1 U8116 ( .A(n6433), .B(n8441), .ZN(n6450) );
  NAND2_X1 U8117 ( .A1(n8509), .A2(n8513), .ZN(n6510) );
  NAND2_X1 U8118 ( .A1(n4376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6435) );
  XNOR2_X1 U8119 ( .A(n6435), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8462) );
  NAND2_X1 U8120 ( .A1(n8326), .A2(n8462), .ZN(n8471) );
  NAND2_X1 U8121 ( .A1(n6436), .A2(n8511), .ZN(n6437) );
  AND2_X1 U8122 ( .A1(n6445), .A2(n6437), .ZN(n7203) );
  NAND2_X1 U8123 ( .A1(n8697), .A2(n10130), .ZN(n6448) );
  INV_X1 U8124 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n6441) );
  INV_X1 U8125 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6438) );
  OR2_X1 U8126 ( .A1(n6145), .A2(n6438), .ZN(n6439) );
  OAI211_X1 U8127 ( .C1(n6442), .C2(n6441), .A(n6440), .B(n6439), .ZN(n6443)
         );
  INV_X1 U8128 ( .A(n6443), .ZN(n6444) );
  NAND2_X1 U8129 ( .A1(n8455), .A2(n6444), .ZN(n8696) );
  NOR2_X2 U8130 ( .A1(n7203), .A2(n8457), .ZN(n10132) );
  NAND2_X1 U8131 ( .A1(n6445), .A2(P2_B_REG_SCAN_IN), .ZN(n6446) );
  AND2_X1 U8132 ( .A1(n10132), .A2(n6446), .ZN(n8805) );
  NAND2_X1 U8133 ( .A1(n8696), .A2(n8805), .ZN(n6447) );
  NAND2_X1 U8134 ( .A1(n6448), .A2(n6447), .ZN(n6449) );
  INV_X1 U8135 ( .A(n7345), .ZN(n6453) );
  INV_X1 U8136 ( .A(n8708), .ZN(n6452) );
  INV_X1 U8137 ( .A(n7214), .ZN(n6451) );
  NAND2_X1 U8138 ( .A1(n6452), .A2(n6451), .ZN(n7216) );
  NAND2_X1 U8139 ( .A1(n6453), .A2(n8329), .ZN(n7346) );
  NAND2_X1 U8140 ( .A1(n7346), .A2(n8333), .ZN(n10144) );
  NAND2_X1 U8141 ( .A1(n10144), .A2(n10150), .ZN(n6454) );
  NAND2_X1 U8142 ( .A1(n6454), .A2(n8338), .ZN(n10136) );
  NAND2_X1 U8143 ( .A1(n7482), .A2(n10177), .ZN(n8361) );
  OR2_X1 U8144 ( .A1(n7482), .A2(n10177), .ZN(n7491) );
  INV_X1 U8145 ( .A(n7451), .ZN(n10179) );
  NAND2_X1 U8146 ( .A1(n8707), .A2(n10179), .ZN(n8366) );
  AND2_X1 U8147 ( .A1(n7491), .A2(n8366), .ZN(n8347) );
  NAND2_X1 U8148 ( .A1(n7476), .A2(n8347), .ZN(n6455) );
  OR2_X1 U8149 ( .A1(n8707), .A2(n10179), .ZN(n8362) );
  NAND2_X1 U8150 ( .A1(n6455), .A2(n8362), .ZN(n7702) );
  NAND2_X1 U8151 ( .A1(n8706), .A2(n10184), .ZN(n8365) );
  NAND2_X1 U8152 ( .A1(n8368), .A2(n8365), .ZN(n8482) );
  INV_X1 U8153 ( .A(n8482), .ZN(n7701) );
  AND2_X1 U8154 ( .A1(n8352), .A2(n7685), .ZN(n8371) );
  NAND2_X1 U8155 ( .A1(n7861), .A2(n7963), .ZN(n8357) );
  NAND2_X1 U8156 ( .A1(n7760), .A2(n8487), .ZN(n7759) );
  NAND2_X1 U8157 ( .A1(n7759), .A2(n8373), .ZN(n7961) );
  OR2_X1 U8158 ( .A1(n8076), .A2(n8075), .ZN(n8378) );
  NAND2_X1 U8159 ( .A1(n8076), .A2(n8075), .ZN(n8377) );
  XNOR2_X1 U8160 ( .A(n10220), .B(n8700), .ZN(n8384) );
  NAND2_X1 U8161 ( .A1(n8043), .A2(n8384), .ZN(n8044) );
  INV_X1 U8162 ( .A(n8700), .ZN(n8386) );
  OR2_X1 U8163 ( .A1(n10220), .A2(n8386), .ZN(n8388) );
  NAND2_X1 U8164 ( .A1(n8044), .A2(n8388), .ZN(n8121) );
  INV_X1 U8165 ( .A(n8397), .ZN(n6457) );
  INV_X1 U8166 ( .A(n6458), .ZN(n8403) );
  INV_X1 U8167 ( .A(n8402), .ZN(n8405) );
  AOI21_X1 U8168 ( .B1(n8966), .B2(n8406), .A(n8405), .ZN(n8955) );
  NAND2_X1 U8169 ( .A1(n8955), .A2(n8954), .ZN(n8953) );
  AND2_X1 U8170 ( .A1(n8409), .A2(n8924), .ZN(n8412) );
  AND2_X1 U8171 ( .A1(n8896), .A2(n8420), .ZN(n8417) );
  INV_X1 U8172 ( .A(n8420), .ZN(n6459) );
  AND2_X1 U8173 ( .A1(n8421), .A2(n8897), .ZN(n8418) );
  NOR2_X1 U8174 ( .A1(n9096), .A2(n8865), .ZN(n8425) );
  AND2_X1 U8175 ( .A1(n9090), .A2(n8854), .ZN(n8474) );
  INV_X1 U8176 ( .A(n8474), .ZN(n6461) );
  NAND2_X1 U8177 ( .A1(n9096), .A2(n8865), .ZN(n8869) );
  AND2_X1 U8178 ( .A1(n6461), .A2(n8869), .ZN(n8428) );
  NAND2_X1 U8179 ( .A1(n8868), .A2(n8428), .ZN(n6462) );
  INV_X1 U8180 ( .A(n8844), .ZN(n8864) );
  OR2_X1 U8181 ( .A1(n9083), .A2(n8864), .ZN(n8432) );
  INV_X1 U8182 ( .A(n8432), .ZN(n6463) );
  NAND2_X1 U8183 ( .A1(n9083), .A2(n8864), .ZN(n8431) );
  NAND2_X1 U8184 ( .A1(n9076), .A2(n8855), .ZN(n8435) );
  INV_X1 U8185 ( .A(n8435), .ZN(n6464) );
  NAND2_X1 U8186 ( .A1(n9070), .A2(n8826), .ZN(n8438) );
  NAND2_X1 U8187 ( .A1(n9064), .A2(n8837), .ZN(n6466) );
  NOR2_X1 U8188 ( .A1(n9064), .A2(n8837), .ZN(n6465) );
  INV_X1 U8189 ( .A(n8462), .ZN(n7207) );
  NAND2_X1 U8190 ( .A1(n5529), .A2(n8513), .ZN(n6500) );
  INV_X1 U8191 ( .A(n8513), .ZN(n6468) );
  NAND2_X1 U8192 ( .A1(n6468), .A2(n7348), .ZN(n10210) );
  AOI21_X1 U8193 ( .B1(n7209), .B2(n6500), .A(n10221), .ZN(n6469) );
  OR2_X1 U8194 ( .A1(n7209), .A2(n8457), .ZN(n7012) );
  AND2_X1 U8195 ( .A1(n6469), .A2(n7012), .ZN(n7965) );
  NAND2_X1 U8196 ( .A1(n8812), .A2(n7965), .ZN(n6470) );
  NAND2_X1 U8197 ( .A1(n8509), .A2(n7207), .ZN(n7349) );
  NOR2_X1 U8198 ( .A1(n7349), .A2(n8513), .ZN(n10207) );
  NOR2_X1 U8199 ( .A1(n8813), .A2(n6472), .ZN(n6517) );
  INV_X1 U8200 ( .A(P2_B_REG_SCAN_IN), .ZN(n6473) );
  XNOR2_X1 U8201 ( .A(n6474), .B(n6473), .ZN(n6475) );
  NAND2_X1 U8202 ( .A1(n6475), .A2(n8065), .ZN(n6477) );
  INV_X1 U8203 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6478) );
  NAND2_X1 U8204 ( .A1(n6483), .A2(n6478), .ZN(n6482) );
  INV_X1 U8205 ( .A(n4333), .ZN(n6480) );
  NAND2_X1 U8206 ( .A1(n6480), .A2(n6484), .ZN(n6481) );
  NAND2_X1 U8207 ( .A1(n6482), .A2(n6481), .ZN(n6513) );
  INV_X1 U8208 ( .A(n6513), .ZN(n9150) );
  INV_X1 U8209 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6899) );
  NAND2_X1 U8210 ( .A1(n6483), .A2(n6899), .ZN(n6485) );
  NAND2_X1 U8211 ( .A1(n6484), .A2(n6474), .ZN(n6897) );
  INV_X1 U8212 ( .A(n7210), .ZN(n7316) );
  AND2_X1 U8213 ( .A1(n9150), .A2(n7316), .ZN(n6508) );
  INV_X1 U8214 ( .A(n6508), .ZN(n6499) );
  NAND2_X1 U8215 ( .A1(n6995), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9149) );
  NOR2_X1 U8216 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .ZN(
        n6490) );
  NOR4_X1 U8217 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6489) );
  NOR4_X1 U8218 ( .A1(P2_D_REG_28__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6488) );
  NOR4_X1 U8219 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6487) );
  NAND4_X1 U8220 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n6496)
         );
  NOR4_X1 U8221 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6494) );
  NOR4_X1 U8222 ( .A1(P2_D_REG_9__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n6493) );
  NOR4_X1 U8223 ( .A1(P2_D_REG_19__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6492) );
  NOR4_X1 U8224 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_10__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6491) );
  NAND4_X1 U8225 ( .A1(n6494), .A2(n6493), .A3(n6492), .A4(n6491), .ZN(n6495)
         );
  OAI21_X1 U8226 ( .B1(n6496), .B2(n6495), .A(n6483), .ZN(n6512) );
  NAND2_X1 U8227 ( .A1(n7209), .A2(n8458), .ZN(n6994) );
  NAND2_X1 U8228 ( .A1(n6512), .A2(n6994), .ZN(n6497) );
  NOR2_X1 U8229 ( .A1(n9149), .A2(n6497), .ZN(n6498) );
  AND2_X1 U8230 ( .A1(n6499), .A2(n6498), .ZN(n7318) );
  INV_X1 U8231 ( .A(n7349), .ZN(n10147) );
  NOR2_X1 U8232 ( .A1(n7009), .A2(n7210), .ZN(n6502) );
  OR2_X1 U8233 ( .A1(n6500), .A2(n7207), .ZN(n6501) );
  NAND2_X1 U8234 ( .A1(n6501), .A2(n8457), .ZN(n7315) );
  MUX2_X1 U8235 ( .A(n6502), .B(n9150), .S(n7315), .Z(n6503) );
  AND2_X2 U8236 ( .A1(n7318), .A2(n6503), .ZN(n10243) );
  OR2_X1 U8237 ( .A1(n6517), .A2(n6505), .ZN(n6507) );
  INV_X1 U8238 ( .A(n6504), .ZN(n8814) );
  NAND2_X1 U8239 ( .A1(n10243), .A2(n10221), .ZN(n9037) );
  NAND2_X1 U8240 ( .A1(n6505), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8241 ( .A1(n6507), .A2(n4962), .ZN(P2_U3488) );
  NAND2_X1 U8242 ( .A1(n6508), .A2(n6512), .ZN(n6992) );
  INV_X1 U8243 ( .A(n6992), .ZN(n6509) );
  NAND2_X1 U8244 ( .A1(n6509), .A2(n7010), .ZN(n7008) );
  NAND2_X1 U8245 ( .A1(n7348), .A2(n8462), .ZN(n8504) );
  OR2_X1 U8246 ( .A1(n6510), .A2(n8504), .ZN(n6993) );
  AND2_X1 U8247 ( .A1(n7012), .A2(n6993), .ZN(n6511) );
  OR2_X1 U8248 ( .A1(n7008), .A2(n6511), .ZN(n6516) );
  NAND3_X1 U8249 ( .A1(n6513), .A2(n7210), .A3(n6512), .ZN(n6999) );
  OR2_X1 U8250 ( .A1(n9149), .A2(n6999), .ZN(n7013) );
  INV_X1 U8251 ( .A(n7013), .ZN(n7005) );
  AND2_X1 U8252 ( .A1(n8457), .A2(n10210), .ZN(n6514) );
  NAND2_X1 U8253 ( .A1(n6993), .A2(n6514), .ZN(n7003) );
  NAND2_X1 U8254 ( .A1(n7349), .A2(n10221), .ZN(n8981) );
  NAND2_X1 U8255 ( .A1(n7003), .A2(n8981), .ZN(n6991) );
  NAND2_X1 U8256 ( .A1(n7005), .A2(n6991), .ZN(n6515) );
  NAND2_X1 U8257 ( .A1(n10222), .A2(n10221), .ZN(n9122) );
  NAND2_X1 U8258 ( .A1(n6519), .A2(n4960), .ZN(P2_U3456) );
  INV_X1 U8259 ( .A(n6525), .ZN(n6520) );
  NAND2_X1 U8260 ( .A1(n9322), .A2(n6549), .ZN(n6527) );
  OR2_X1 U8261 ( .A1(n6521), .A2(n6525), .ZN(n7644) );
  AND2_X1 U8262 ( .A1(n6768), .A2(n6525), .ZN(n6526) );
  INV_X2 U8263 ( .A(n8258), .ZN(n9186) );
  INV_X1 U8264 ( .A(n6533), .ZN(n6531) );
  NAND2_X1 U8265 ( .A1(n9322), .A2(n6746), .ZN(n6529) );
  OR2_X1 U8266 ( .A1(n7436), .A2(n6545), .ZN(n6528) );
  AND2_X1 U8267 ( .A1(n6529), .A2(n6528), .ZN(n6532) );
  INV_X1 U8268 ( .A(n6532), .ZN(n6530) );
  NAND2_X1 U8269 ( .A1(n6531), .A2(n6530), .ZN(n6534) );
  NAND2_X1 U8270 ( .A1(n6533), .A2(n6532), .ZN(n7236) );
  NAND2_X1 U8271 ( .A1(n9324), .A2(n6549), .ZN(n6537) );
  INV_X1 U8272 ( .A(n6557), .ZN(n6535) );
  NAND2_X1 U8273 ( .A1(n6535), .A2(n7572), .ZN(n6536) );
  NAND2_X1 U8274 ( .A1(n6537), .A2(n6536), .ZN(n6541) );
  NOR2_X1 U8275 ( .A1(n6768), .A2(n6875), .ZN(n6538) );
  OR2_X1 U8276 ( .A1(n6541), .A2(n6538), .ZN(n6803) );
  NAND2_X1 U8277 ( .A1(n9324), .A2(n6746), .ZN(n6540) );
  INV_X1 U8278 ( .A(n6768), .ZN(n6785) );
  AOI22_X1 U8279 ( .A1(n7572), .A2(n4330), .B1(n6785), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6539) );
  NAND2_X1 U8280 ( .A1(n6540), .A2(n6539), .ZN(n6802) );
  NAND2_X1 U8281 ( .A1(n6803), .A2(n6802), .ZN(n6544) );
  INV_X1 U8282 ( .A(n6541), .ZN(n6542) );
  NAND2_X1 U8283 ( .A1(n6542), .A2(n9186), .ZN(n6543) );
  NAND2_X1 U8284 ( .A1(n9321), .A2(n4330), .ZN(n6547) );
  NAND2_X1 U8285 ( .A1(n6547), .A2(n6546), .ZN(n6548) );
  XNOR2_X1 U8286 ( .A(n6548), .B(n9186), .ZN(n6553) );
  NAND2_X1 U8287 ( .A1(n9321), .A2(n6746), .ZN(n6551) );
  OR2_X1 U8288 ( .A1(n10050), .A2(n6545), .ZN(n6550) );
  AND2_X1 U8289 ( .A1(n6551), .A2(n6550), .ZN(n6552) );
  NAND2_X1 U8290 ( .A1(n6553), .A2(n6552), .ZN(n6556) );
  OR2_X1 U8291 ( .A1(n6553), .A2(n6552), .ZN(n6554) );
  AND2_X1 U8292 ( .A1(n6556), .A2(n6554), .ZN(n7235) );
  NAND2_X1 U8293 ( .A1(n6555), .A2(n7235), .ZN(n7239) );
  NAND2_X1 U8294 ( .A1(n7239), .A2(n6556), .ZN(n7270) );
  NAND2_X1 U8295 ( .A1(n9320), .A2(n4330), .ZN(n6559) );
  OR2_X1 U8296 ( .A1(n6557), .A2(n7431), .ZN(n6558) );
  NAND2_X1 U8297 ( .A1(n6559), .A2(n6558), .ZN(n6560) );
  NAND2_X1 U8298 ( .A1(n9320), .A2(n6746), .ZN(n6562) );
  OR2_X1 U8299 ( .A1(n7431), .A2(n6545), .ZN(n6561) );
  NAND2_X1 U8300 ( .A1(n6562), .A2(n6561), .ZN(n6568) );
  XNOR2_X1 U8301 ( .A(n6570), .B(n6568), .ZN(n7271) );
  NAND2_X1 U8302 ( .A1(n7270), .A2(n7271), .ZN(n7269) );
  NAND2_X1 U8303 ( .A1(n9319), .A2(n4330), .ZN(n6564) );
  OR2_X1 U8304 ( .A1(n6557), .A2(n7593), .ZN(n6563) );
  NAND2_X1 U8305 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  XNOR2_X1 U8306 ( .A(n6565), .B(n9186), .ZN(n6572) );
  NAND2_X1 U8307 ( .A1(n9319), .A2(n6746), .ZN(n6567) );
  OR2_X1 U8308 ( .A1(n7593), .A2(n6545), .ZN(n6566) );
  NAND2_X1 U8309 ( .A1(n6567), .A2(n6566), .ZN(n6573) );
  XNOR2_X1 U8310 ( .A(n6572), .B(n6573), .ZN(n7280) );
  INV_X1 U8311 ( .A(n6568), .ZN(n6569) );
  NAND2_X1 U8312 ( .A1(n6570), .A2(n6569), .ZN(n7281) );
  AND2_X1 U8313 ( .A1(n7280), .A2(n7281), .ZN(n6571) );
  NAND2_X1 U8314 ( .A1(n7269), .A2(n6571), .ZN(n7279) );
  INV_X1 U8315 ( .A(n6572), .ZN(n6574) );
  NAND2_X1 U8316 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  NAND2_X1 U8317 ( .A1(n7279), .A2(n6575), .ZN(n6583) );
  NAND2_X1 U8318 ( .A1(n9318), .A2(n4330), .ZN(n6577) );
  OR2_X1 U8319 ( .A1(n6557), .A2(n7582), .ZN(n6576) );
  NAND2_X1 U8320 ( .A1(n6577), .A2(n6576), .ZN(n6578) );
  XNOR2_X1 U8321 ( .A(n6578), .B(n8258), .ZN(n6582) );
  INV_X1 U8322 ( .A(n6582), .ZN(n6579) );
  NAND2_X1 U8323 ( .A1(n9318), .A2(n6746), .ZN(n6581) );
  OR2_X1 U8324 ( .A1(n7582), .A2(n6545), .ZN(n6580) );
  AND2_X1 U8325 ( .A1(n6581), .A2(n6580), .ZN(n7533) );
  NAND2_X1 U8326 ( .A1(n9317), .A2(n4330), .ZN(n6585) );
  INV_X2 U8327 ( .A(n6557), .ZN(n9183) );
  NAND2_X1 U8328 ( .A1(n10056), .A2(n9183), .ZN(n6584) );
  NAND2_X1 U8329 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  XNOR2_X1 U8330 ( .A(n6586), .B(n8258), .ZN(n6589) );
  NAND2_X1 U8331 ( .A1(n9317), .A2(n6746), .ZN(n6588) );
  NAND2_X1 U8332 ( .A1(n10056), .A2(n4330), .ZN(n6587) );
  NAND2_X1 U8333 ( .A1(n6588), .A2(n6587), .ZN(n6590) );
  NAND2_X1 U8334 ( .A1(n6589), .A2(n6590), .ZN(n7716) );
  NAND2_X1 U8335 ( .A1(n7715), .A2(n7716), .ZN(n7660) );
  INV_X1 U8336 ( .A(n6589), .ZN(n6592) );
  INV_X1 U8337 ( .A(n6590), .ZN(n6591) );
  NAND2_X1 U8338 ( .A1(n6592), .A2(n6591), .ZN(n7718) );
  NAND2_X1 U8339 ( .A1(n9316), .A2(n4330), .ZN(n6593) );
  OAI21_X1 U8340 ( .B1(n7697), .B2(n6557), .A(n6593), .ZN(n6594) );
  XNOR2_X1 U8341 ( .A(n6594), .B(n9186), .ZN(n6613) );
  OR2_X1 U8342 ( .A1(n7697), .A2(n6545), .ZN(n6596) );
  NAND2_X1 U8343 ( .A1(n9316), .A2(n6746), .ZN(n6595) );
  NAND2_X1 U8344 ( .A1(n6596), .A2(n6595), .ZN(n6612) );
  INV_X1 U8345 ( .A(n6612), .ZN(n6597) );
  NAND2_X1 U8346 ( .A1(n6613), .A2(n6597), .ZN(n6611) );
  AND2_X1 U8347 ( .A1(n7718), .A2(n6611), .ZN(n7811) );
  NAND2_X1 U8348 ( .A1(n7952), .A2(n9183), .ZN(n6599) );
  OR2_X1 U8349 ( .A1(n7881), .A2(n6545), .ZN(n6598) );
  NAND2_X1 U8350 ( .A1(n6599), .A2(n6598), .ZN(n6600) );
  XNOR2_X1 U8351 ( .A(n6600), .B(n8258), .ZN(n7944) );
  NAND2_X1 U8352 ( .A1(n7952), .A2(n4330), .ZN(n6603) );
  OR2_X1 U8353 ( .A1(n7881), .A2(n6601), .ZN(n6602) );
  NAND2_X1 U8354 ( .A1(n6603), .A2(n6602), .ZN(n6617) );
  NAND2_X1 U8355 ( .A1(n10012), .A2(n4330), .ZN(n6605) );
  OR2_X1 U8356 ( .A1(n7788), .A2(n6601), .ZN(n6604) );
  NAND2_X1 U8357 ( .A1(n6605), .A2(n6604), .ZN(n7814) );
  NAND2_X1 U8358 ( .A1(n10012), .A2(n9183), .ZN(n6607) );
  OR2_X1 U8359 ( .A1(n7788), .A2(n6545), .ZN(n6606) );
  NAND2_X1 U8360 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  XNOR2_X1 U8361 ( .A(n6608), .B(n8258), .ZN(n7939) );
  OAI22_X1 U8362 ( .A1(n7944), .A2(n6617), .B1(n7814), .B2(n7939), .ZN(n6615)
         );
  INV_X1 U8363 ( .A(n6615), .ZN(n6609) );
  AND2_X1 U8364 ( .A1(n7811), .A2(n6609), .ZN(n6610) );
  NAND2_X1 U8365 ( .A1(n7660), .A2(n6610), .ZN(n6623) );
  INV_X1 U8366 ( .A(n6611), .ZN(n6614) );
  XNOR2_X1 U8367 ( .A(n6613), .B(n6612), .ZN(n7662) );
  NAND2_X1 U8368 ( .A1(n7939), .A2(n7814), .ZN(n6616) );
  INV_X1 U8369 ( .A(n6617), .ZN(n7943) );
  NAND2_X1 U8370 ( .A1(n6616), .A2(n7943), .ZN(n6619) );
  INV_X1 U8371 ( .A(n6616), .ZN(n6618) );
  AOI22_X1 U8372 ( .A1(n7944), .A2(n6619), .B1(n6618), .B2(n6617), .ZN(n6620)
         );
  NAND2_X1 U8373 ( .A1(n9862), .A2(n9183), .ZN(n6625) );
  OR2_X1 U8374 ( .A1(n8230), .A2(n6545), .ZN(n6624) );
  NAND2_X1 U8375 ( .A1(n6625), .A2(n6624), .ZN(n6626) );
  NOR2_X1 U8376 ( .A1(n8230), .A2(n6601), .ZN(n6627) );
  AOI21_X1 U8377 ( .B1(n9862), .B2(n4330), .A(n6627), .ZN(n9859) );
  NAND2_X1 U8378 ( .A1(n9886), .A2(n9183), .ZN(n6629) );
  NAND2_X1 U8379 ( .A1(n9312), .A2(n4330), .ZN(n6628) );
  NAND2_X1 U8380 ( .A1(n6629), .A2(n6628), .ZN(n6630) );
  XNOR2_X1 U8381 ( .A(n6630), .B(n8258), .ZN(n9876) );
  NAND2_X1 U8382 ( .A1(n9886), .A2(n4330), .ZN(n6632) );
  NAND2_X1 U8383 ( .A1(n9312), .A2(n6746), .ZN(n6631) );
  NAND2_X1 U8384 ( .A1(n6632), .A2(n6631), .ZN(n9877) );
  NAND2_X1 U8385 ( .A1(n9876), .A2(n9877), .ZN(n9875) );
  OAI21_X1 U8386 ( .B1(n9857), .B2(n9859), .A(n9875), .ZN(n6638) );
  INV_X1 U8387 ( .A(n9876), .ZN(n6636) );
  INV_X1 U8388 ( .A(n9857), .ZN(n9879) );
  INV_X1 U8389 ( .A(n9859), .ZN(n6633) );
  OAI21_X1 U8390 ( .B1(n9879), .B2(n6633), .A(n9877), .ZN(n6635) );
  NOR2_X1 U8391 ( .A1(n9877), .A2(n6633), .ZN(n6634) );
  NAND2_X1 U8392 ( .A1(n9872), .A2(n9183), .ZN(n6640) );
  NAND2_X1 U8393 ( .A1(n9311), .A2(n4330), .ZN(n6639) );
  NAND2_X1 U8394 ( .A1(n6640), .A2(n6639), .ZN(n6641) );
  XNOR2_X1 U8395 ( .A(n6641), .B(n9186), .ZN(n6643) );
  AND2_X1 U8396 ( .A1(n9311), .A2(n6746), .ZN(n6642) );
  AOI21_X1 U8397 ( .B1(n9872), .B2(n4330), .A(n6642), .ZN(n6644) );
  NAND2_X1 U8398 ( .A1(n6643), .A2(n6644), .ZN(n6648) );
  INV_X1 U8399 ( .A(n6643), .ZN(n6646) );
  INV_X1 U8400 ( .A(n6644), .ZN(n6645) );
  NAND2_X1 U8401 ( .A1(n6646), .A2(n6645), .ZN(n6647) );
  NAND2_X1 U8402 ( .A1(n8163), .A2(n9183), .ZN(n6650) );
  OR2_X1 U8403 ( .A1(n8105), .A2(n6545), .ZN(n6649) );
  NAND2_X1 U8404 ( .A1(n6650), .A2(n6649), .ZN(n6651) );
  XNOR2_X1 U8405 ( .A(n6651), .B(n8258), .ZN(n6653) );
  NOR2_X1 U8406 ( .A1(n8105), .A2(n6601), .ZN(n6652) );
  AOI21_X1 U8407 ( .B1(n8163), .B2(n4330), .A(n6652), .ZN(n6654) );
  XNOR2_X1 U8408 ( .A(n6653), .B(n6654), .ZN(n7925) );
  INV_X1 U8409 ( .A(n6653), .ZN(n6655) );
  NAND2_X1 U8410 ( .A1(n6655), .A2(n6654), .ZN(n6656) );
  NAND2_X1 U8411 ( .A1(n9728), .A2(n9183), .ZN(n6658) );
  NAND2_X1 U8412 ( .A1(n9309), .A2(n4330), .ZN(n6657) );
  NAND2_X1 U8413 ( .A1(n6658), .A2(n6657), .ZN(n6659) );
  XNOR2_X1 U8414 ( .A(n6659), .B(n9186), .ZN(n6663) );
  NAND2_X1 U8415 ( .A1(n6662), .A2(n6663), .ZN(n8111) );
  NAND2_X1 U8416 ( .A1(n9728), .A2(n4330), .ZN(n6661) );
  NAND2_X1 U8417 ( .A1(n9309), .A2(n6746), .ZN(n6660) );
  NAND2_X1 U8418 ( .A1(n6661), .A2(n6660), .ZN(n8110) );
  NAND2_X1 U8419 ( .A1(n8111), .A2(n8110), .ZN(n8109) );
  NAND2_X1 U8420 ( .A1(n8109), .A2(n8113), .ZN(n6671) );
  INV_X1 U8421 ( .A(n6671), .ZN(n6669) );
  NAND2_X1 U8422 ( .A1(n8274), .A2(n9183), .ZN(n6667) );
  NAND2_X1 U8423 ( .A1(n9308), .A2(n4330), .ZN(n6666) );
  NAND2_X1 U8424 ( .A1(n6667), .A2(n6666), .ZN(n6668) );
  XNOR2_X1 U8425 ( .A(n6668), .B(n9186), .ZN(n6670) );
  INV_X1 U8426 ( .A(n6670), .ZN(n6672) );
  OAI22_X1 U8427 ( .A1(n9781), .A2(n6545), .B1(n8277), .B2(n6601), .ZN(n8166)
         );
  INV_X1 U8428 ( .A(n9240), .ZN(n9307) );
  AOI22_X1 U8429 ( .A1(n9628), .A2(n4330), .B1(n6746), .B2(n9307), .ZN(n6677)
         );
  NAND2_X1 U8430 ( .A1(n9628), .A2(n9183), .ZN(n6675) );
  OR2_X1 U8431 ( .A1(n9240), .A2(n6545), .ZN(n6674) );
  NAND2_X1 U8432 ( .A1(n6675), .A2(n6674), .ZN(n6676) );
  XNOR2_X1 U8433 ( .A(n6676), .B(n8258), .ZN(n6679) );
  XOR2_X1 U8434 ( .A(n6677), .B(n6679), .Z(n9226) );
  INV_X1 U8435 ( .A(n6677), .ZN(n6678) );
  NOR2_X1 U8436 ( .A1(n6679), .A2(n6678), .ZN(n9236) );
  NAND2_X1 U8437 ( .A1(n9610), .A2(n9183), .ZN(n6681) );
  NAND2_X1 U8438 ( .A1(n9306), .A2(n4330), .ZN(n6680) );
  NAND2_X1 U8439 ( .A1(n6681), .A2(n6680), .ZN(n6682) );
  XNOR2_X1 U8440 ( .A(n6682), .B(n9186), .ZN(n6684) );
  AND2_X1 U8441 ( .A1(n9306), .A2(n6746), .ZN(n6683) );
  AOI21_X1 U8442 ( .B1(n9610), .B2(n4330), .A(n6683), .ZN(n6685) );
  XNOR2_X1 U8443 ( .A(n6684), .B(n6685), .ZN(n9235) );
  INV_X1 U8444 ( .A(n6684), .ZN(n6687) );
  INV_X1 U8445 ( .A(n6685), .ZN(n6686) );
  AOI22_X1 U8446 ( .A1(n9708), .A2(n4330), .B1(n6746), .B2(n9305), .ZN(n9173)
         );
  AOI22_X1 U8447 ( .A1(n9708), .A2(n9183), .B1(n4330), .B2(n9305), .ZN(n6688)
         );
  XNOR2_X1 U8448 ( .A(n6688), .B(n8258), .ZN(n9172) );
  NAND2_X1 U8449 ( .A1(n9587), .A2(n9183), .ZN(n6690) );
  NAND2_X1 U8450 ( .A1(n9304), .A2(n4330), .ZN(n6689) );
  NAND2_X1 U8451 ( .A1(n6690), .A2(n6689), .ZN(n6691) );
  XNOR2_X1 U8452 ( .A(n6691), .B(n9186), .ZN(n6701) );
  AND2_X1 U8453 ( .A1(n9304), .A2(n6746), .ZN(n6692) );
  AOI21_X1 U8454 ( .B1(n9587), .B2(n4330), .A(n6692), .ZN(n6702) );
  NAND2_X1 U8455 ( .A1(n6701), .A2(n6702), .ZN(n9170) );
  NAND2_X1 U8456 ( .A1(n9697), .A2(n9183), .ZN(n6694) );
  INV_X1 U8457 ( .A(n9177), .ZN(n9303) );
  NAND2_X1 U8458 ( .A1(n9303), .A2(n4330), .ZN(n6693) );
  NAND2_X1 U8459 ( .A1(n6694), .A2(n6693), .ZN(n6695) );
  XNOR2_X1 U8460 ( .A(n6695), .B(n9186), .ZN(n6698) );
  INV_X1 U8461 ( .A(n6698), .ZN(n6700) );
  NOR2_X1 U8462 ( .A1(n9177), .A2(n6601), .ZN(n6696) );
  AOI21_X1 U8463 ( .B1(n9697), .B2(n4330), .A(n6696), .ZN(n6697) );
  INV_X1 U8464 ( .A(n6697), .ZN(n6699) );
  AOI21_X1 U8465 ( .B1(n6700), .B2(n6699), .A(n6706), .ZN(n9261) );
  INV_X1 U8466 ( .A(n6701), .ZN(n6704) );
  INV_X1 U8467 ( .A(n6702), .ZN(n6703) );
  NAND2_X1 U8468 ( .A1(n6704), .A2(n6703), .ZN(n9262) );
  INV_X1 U8469 ( .A(n6706), .ZN(n6707) );
  NAND2_X1 U8470 ( .A1(n9260), .A2(n6707), .ZN(n9208) );
  OAI22_X1 U8471 ( .A1(n9762), .A2(n6545), .B1(n8286), .B2(n6601), .ZN(n6711)
         );
  NAND2_X1 U8472 ( .A1(n9558), .A2(n9183), .ZN(n6709) );
  NAND2_X1 U8473 ( .A1(n9302), .A2(n4330), .ZN(n6708) );
  NAND2_X1 U8474 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  XNOR2_X1 U8475 ( .A(n6710), .B(n8258), .ZN(n6712) );
  XOR2_X1 U8476 ( .A(n6711), .B(n6712), .Z(n9209) );
  NAND2_X1 U8477 ( .A1(n9208), .A2(n9209), .ZN(n9207) );
  OR2_X1 U8478 ( .A1(n6712), .A2(n6711), .ZN(n6713) );
  NAND2_X1 U8479 ( .A1(n9207), .A2(n6713), .ZN(n6716) );
  AOI22_X1 U8480 ( .A1(n9685), .A2(n9183), .B1(n4330), .B2(n9301), .ZN(n6714)
         );
  XNOR2_X1 U8481 ( .A(n6714), .B(n8258), .ZN(n6715) );
  NAND2_X1 U8482 ( .A1(n6716), .A2(n6715), .ZN(n6718) );
  NAND2_X1 U8483 ( .A1(n6717), .A2(n6718), .ZN(n9273) );
  OAI22_X1 U8484 ( .A1(n9539), .A2(n6545), .B1(n8287), .B2(n6601), .ZN(n9274)
         );
  NOR2_X2 U8485 ( .A1(n9273), .A2(n9274), .ZN(n9161) );
  OAI22_X1 U8486 ( .A1(n9757), .A2(n6557), .B1(n9276), .B2(n6545), .ZN(n6719)
         );
  XNOR2_X1 U8487 ( .A(n6719), .B(n9186), .ZN(n6721) );
  NOR2_X1 U8488 ( .A1(n9276), .A2(n6601), .ZN(n6720) );
  AOI21_X1 U8489 ( .B1(n9527), .B2(n4330), .A(n6720), .ZN(n6722) );
  NAND2_X1 U8490 ( .A1(n6721), .A2(n6722), .ZN(n9249) );
  INV_X1 U8491 ( .A(n6721), .ZN(n6724) );
  INV_X1 U8492 ( .A(n6722), .ZN(n6723) );
  NAND2_X1 U8493 ( .A1(n6724), .A2(n6723), .ZN(n6725) );
  OAI21_X2 U8494 ( .B1(n9161), .B2(n9163), .A(n9162), .ZN(n9160) );
  NAND2_X1 U8495 ( .A1(n9160), .A2(n9249), .ZN(n6736) );
  NAND2_X1 U8496 ( .A1(n9502), .A2(n9183), .ZN(n6727) );
  NAND2_X1 U8497 ( .A1(n9299), .A2(n4330), .ZN(n6726) );
  NAND2_X1 U8498 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  XNOR2_X1 U8499 ( .A(n6728), .B(n9186), .ZN(n6730) );
  AND2_X1 U8500 ( .A1(n9299), .A2(n6746), .ZN(n6729) );
  AOI21_X1 U8501 ( .B1(n9502), .B2(n4330), .A(n6729), .ZN(n6731) );
  NAND2_X1 U8502 ( .A1(n6730), .A2(n6731), .ZN(n6737) );
  INV_X1 U8503 ( .A(n6730), .ZN(n6733) );
  INV_X1 U8504 ( .A(n6731), .ZN(n6732) );
  NAND2_X1 U8505 ( .A1(n6733), .A2(n6732), .ZN(n6734) );
  NAND2_X1 U8506 ( .A1(n6737), .A2(n6734), .ZN(n9248) );
  NAND2_X1 U8507 ( .A1(n9247), .A2(n6737), .ZN(n9216) );
  OAI22_X1 U8508 ( .A1(n9749), .A2(n6545), .B1(n9252), .B2(n6601), .ZN(n6740)
         );
  OAI22_X1 U8509 ( .A1(n9749), .A2(n6557), .B1(n9252), .B2(n6545), .ZN(n6738)
         );
  XNOR2_X1 U8510 ( .A(n6738), .B(n8258), .ZN(n6739) );
  XOR2_X1 U8511 ( .A(n6740), .B(n6739), .Z(n9217) );
  INV_X1 U8512 ( .A(n6739), .ZN(n6742) );
  INV_X1 U8513 ( .A(n6740), .ZN(n6741) );
  NAND2_X1 U8514 ( .A1(n6742), .A2(n6741), .ZN(n6749) );
  AND2_X1 U8515 ( .A1(n6752), .A2(n6749), .ZN(n6748) );
  NAND2_X1 U8516 ( .A1(n9478), .A2(n9183), .ZN(n6744) );
  NAND2_X1 U8517 ( .A1(n9297), .A2(n4330), .ZN(n6743) );
  NAND2_X1 U8518 ( .A1(n6744), .A2(n6743), .ZN(n6745) );
  XNOR2_X1 U8519 ( .A(n6745), .B(n8258), .ZN(n8263) );
  AND2_X1 U8520 ( .A1(n9297), .A2(n6746), .ZN(n6747) );
  AOI21_X1 U8521 ( .B1(n9478), .B2(n4330), .A(n6747), .ZN(n8261) );
  XNOR2_X1 U8522 ( .A(n8263), .B(n8261), .ZN(n6750) );
  OR2_X1 U8523 ( .A1(n10057), .A2(n6810), .ZN(n6765) );
  NOR2_X1 U8524 ( .A1(n6765), .A2(n9783), .ZN(n6757) );
  INV_X1 U8525 ( .A(n6753), .ZN(n6755) );
  AND2_X1 U8526 ( .A1(n6755), .A2(n6754), .ZN(n7559) );
  NAND2_X1 U8527 ( .A1(n7559), .A2(n6756), .ZN(n6773) );
  INV_X1 U8528 ( .A(n6773), .ZN(n6764) );
  NAND2_X1 U8529 ( .A1(n8266), .A2(n9885), .ZN(n6782) );
  NAND2_X1 U8530 ( .A1(n7563), .A2(n6758), .ZN(n7571) );
  INV_X1 U8531 ( .A(n7571), .ZN(n6759) );
  AND2_X1 U8532 ( .A1(n6813), .A2(n6759), .ZN(n6760) );
  NAND2_X1 U8533 ( .A1(n6764), .A2(n6760), .ZN(n6762) );
  NAND2_X1 U8534 ( .A1(n6813), .A2(n7726), .ZN(n6761) );
  INV_X1 U8535 ( .A(n9286), .ZN(n9253) );
  OAI22_X1 U8536 ( .A1(n9197), .A2(n9275), .B1(n9252), .B2(n9253), .ZN(n9473)
         );
  NOR2_X1 U8537 ( .A1(n6522), .A2(n9783), .ZN(n6763) );
  INV_X1 U8538 ( .A(n9479), .ZN(n6777) );
  NAND2_X1 U8539 ( .A1(n6765), .A2(n7571), .ZN(n6766) );
  NAND2_X1 U8540 ( .A1(n6766), .A2(n6773), .ZN(n6769) );
  NAND3_X1 U8541 ( .A1(n6769), .A2(n6768), .A3(n6767), .ZN(n6770) );
  NAND2_X1 U8542 ( .A1(n6770), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6775) );
  NOR2_X1 U8543 ( .A1(n7562), .A2(n9783), .ZN(n6772) );
  AOI21_X1 U8544 ( .B1(n6773), .B2(n6772), .A(n6080), .ZN(n6774) );
  OAI22_X1 U8545 ( .A1(n6777), .A2(n9890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6776), .ZN(n6778) );
  AOI21_X1 U8546 ( .B1(n9473), .B2(n9882), .A(n6778), .ZN(n6779) );
  INV_X1 U8547 ( .A(n6780), .ZN(n6781) );
  OAI21_X1 U8548 ( .B1(n6783), .B2(n6782), .A(n6781), .ZN(P1_U3240) );
  INV_X1 U8549 ( .A(n8705), .ZN(P2_U3893) );
  INV_X1 U8550 ( .A(n10109), .ZN(n8803) );
  INV_X1 U8551 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n6786) );
  NOR2_X1 U8552 ( .A1(n8803), .A2(n6786), .ZN(n6801) );
  OAI22_X1 U8553 ( .A1(n10128), .A2(n4329), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10148), .ZN(n6800) );
  AOI21_X1 U8554 ( .B1(n6789), .B2(n6788), .A(n6787), .ZN(n6794) );
  INV_X1 U8555 ( .A(n8777), .ZN(n10118) );
  AOI21_X1 U8556 ( .B1(n6792), .B2(n6791), .A(n6790), .ZN(n6793) );
  OAI22_X1 U8557 ( .A1(n6794), .A2(n10122), .B1(n10118), .B2(n6793), .ZN(n6799) );
  AOI211_X1 U8558 ( .C1(n6797), .C2(n6796), .A(n6795), .B(n7406), .ZN(n6798)
         );
  OR4_X1 U8559 ( .A1(n6801), .A2(n6800), .A3(n6799), .A4(n6798), .ZN(P2_U3184)
         );
  NAND2_X1 U8560 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6831) );
  XNOR2_X1 U8561 ( .A(n6803), .B(n6802), .ZN(n6958) );
  NAND3_X1 U8562 ( .A1(n6958), .A2(n6805), .A3(n8191), .ZN(n6808) );
  INV_X1 U8563 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6806) );
  OR2_X1 U8564 ( .A1(n8191), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U8565 ( .A1(n6805), .A2(n6804), .ZN(n6874) );
  INV_X1 U8566 ( .A(P1_U3973), .ZN(n9323) );
  AOI21_X1 U8567 ( .B1(n6806), .B2(n6874), .A(n9323), .ZN(n6807) );
  OAI211_X1 U8568 ( .C1(n6831), .C2(n6827), .A(n6808), .B(n6807), .ZN(n9351)
         );
  INV_X1 U8569 ( .A(n9351), .ZN(n6840) );
  NAND2_X1 U8570 ( .A1(n6810), .A2(n6809), .ZN(n6811) );
  NAND2_X1 U8571 ( .A1(n6812), .A2(n6811), .ZN(n6824) );
  INV_X1 U8572 ( .A(n6824), .ZN(n6814) );
  OR2_X1 U8573 ( .A1(n6813), .A2(n6080), .ZN(n6823) );
  AND2_X1 U8574 ( .A1(n6814), .A2(n6823), .ZN(n6877) );
  NAND2_X1 U8575 ( .A1(n6877), .A2(n8191), .ZN(n9993) );
  XNOR2_X1 U8576 ( .A(n6911), .B(n6815), .ZN(n6822) );
  INV_X1 U8577 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6816) );
  XNOR2_X1 U8578 ( .A(n9328), .B(n6816), .ZN(n9334) );
  AND2_X1 U8579 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9333) );
  NAND2_X1 U8580 ( .A1(n9334), .A2(n9333), .ZN(n9332) );
  NAND2_X1 U8581 ( .A1(n4336), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8582 ( .A1(n9332), .A2(n6817), .ZN(n9343) );
  MUX2_X1 U8583 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n5677), .S(n9341), .Z(n9344)
         );
  NAND2_X1 U8584 ( .A1(n9343), .A2(n9344), .ZN(n9342) );
  NAND2_X1 U8585 ( .A1(n9341), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6818) );
  NAND2_X1 U8586 ( .A1(n9342), .A2(n6818), .ZN(n9356) );
  XNOR2_X1 U8587 ( .A(n9354), .B(n6819), .ZN(n9357) );
  NAND2_X1 U8588 ( .A1(n9356), .A2(n9357), .ZN(n9355) );
  NAND2_X1 U8589 ( .A1(n9354), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6820) );
  NAND2_X1 U8590 ( .A1(n9355), .A2(n6820), .ZN(n6821) );
  NAND2_X1 U8591 ( .A1(n6821), .A2(n6822), .ZN(n6909) );
  OAI21_X1 U8592 ( .B1(n6822), .B2(n6821), .A(n6909), .ZN(n6826) );
  NAND2_X1 U8593 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n7284) );
  NAND2_X1 U8594 ( .A1(n6824), .A2(n6823), .ZN(n10008) );
  INV_X1 U8595 ( .A(n10008), .ZN(n9422) );
  NAND2_X1 U8596 ( .A1(n9422), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6825) );
  OAI211_X1 U8597 ( .C1(n9993), .C2(n6826), .A(n7284), .B(n6825), .ZN(n6839)
         );
  INV_X1 U8598 ( .A(n6911), .ZN(n6854) );
  NAND2_X1 U8599 ( .A1(n6877), .A2(n8217), .ZN(n9974) );
  INV_X1 U8600 ( .A(n6827), .ZN(n6828) );
  NAND2_X1 U8601 ( .A1(n6877), .A2(n6828), .ZN(n9999) );
  XNOR2_X1 U8602 ( .A(n6911), .B(n6829), .ZN(n6836) );
  XNOR2_X1 U8603 ( .A(n4336), .B(n6830), .ZN(n9331) );
  INV_X1 U8604 ( .A(n6831), .ZN(n9330) );
  NAND2_X1 U8605 ( .A1(n9331), .A2(n9330), .ZN(n9329) );
  NAND2_X1 U8606 ( .A1(n4336), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6832) );
  NAND2_X1 U8607 ( .A1(n9329), .A2(n6832), .ZN(n9346) );
  MUX2_X1 U8608 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n5676), .S(n9341), .Z(n9347)
         );
  NAND2_X1 U8609 ( .A1(n9346), .A2(n9347), .ZN(n9345) );
  NAND2_X1 U8610 ( .A1(n9341), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6833) );
  NAND2_X1 U8611 ( .A1(n9345), .A2(n6833), .ZN(n9359) );
  XNOR2_X1 U8612 ( .A(n9354), .B(n10022), .ZN(n9360) );
  NAND2_X1 U8613 ( .A1(n9359), .A2(n9360), .ZN(n9358) );
  NAND2_X1 U8614 ( .A1(n9354), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U8615 ( .A1(n9358), .A2(n6834), .ZN(n6835) );
  OAI21_X1 U8616 ( .B1(n6836), .B2(n6835), .A(n6905), .ZN(n6837) );
  OAI22_X1 U8617 ( .A1(n6854), .A2(n9974), .B1(n9999), .B2(n6837), .ZN(n6838)
         );
  OR3_X1 U8618 ( .A1(n6840), .A2(n6839), .A3(n6838), .ZN(P1_U3247) );
  XNOR2_X1 U8619 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  MUX2_X1 U8620 ( .A(n6841), .B(n10089), .S(P2_STATE_REG_SCAN_IN), .Z(n6842)
         );
  INV_X1 U8621 ( .A(n6842), .ZN(P2_U3295) );
  OR2_X1 U8622 ( .A1(n6846), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8565) );
  INV_X1 U8623 ( .A(n8565), .ZN(n9790) );
  AOI22_X1 U8624 ( .A1(n9790), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(n4336), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6843) );
  OAI21_X1 U8625 ( .B1(n6847), .B2(n9792), .A(n6843), .ZN(P1_U3354) );
  AOI22_X1 U8626 ( .A1(n9790), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(n9341), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6844) );
  OAI21_X1 U8627 ( .B1(n6857), .B2(n9792), .A(n6844), .ZN(P1_U3353) );
  AOI22_X1 U8628 ( .A1(n9354), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n9790), .ZN(n6845) );
  OAI21_X1 U8629 ( .B1(n6859), .B2(n9792), .A(n6845), .ZN(P1_U3352) );
  AND2_X1 U8630 ( .A1(n6846), .A2(P2_U3151), .ZN(n9156) );
  INV_X1 U8631 ( .A(n9156), .ZN(n6964) );
  OAI222_X1 U8632 ( .A1(n6964), .A2(n6848), .B1(n9158), .B2(n6847), .C1(
        P2_U3151), .C2(n7425), .ZN(P2_U3294) );
  INV_X1 U8633 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6850) );
  OAI222_X1 U8634 ( .A1(n6964), .A2(n6850), .B1(n9158), .B2(n6853), .C1(
        P2_U3151), .C2(n6849), .ZN(P2_U3291) );
  AOI22_X1 U8635 ( .A1(n6949), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9790), .ZN(n6851) );
  OAI21_X1 U8636 ( .B1(n6855), .B2(n9792), .A(n6851), .ZN(P1_U3350) );
  INV_X1 U8637 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6852) );
  OAI222_X1 U8638 ( .A1(n6854), .A2(P1_U3086), .B1(n9792), .B2(n6853), .C1(
        n6852), .C2(n8565), .ZN(P1_U3351) );
  OAI222_X1 U8639 ( .A1(n6964), .A2(n6856), .B1(n9158), .B2(n6855), .C1(
        P2_U3151), .C2(n5478), .ZN(P2_U3290) );
  OAI222_X1 U8640 ( .A1(n6964), .A2(n6858), .B1(n9158), .B2(n6857), .C1(
        P2_U3151), .C2(n4329), .ZN(P2_U3293) );
  OAI222_X1 U8641 ( .A1(n6964), .A2(n6860), .B1(n9158), .B2(n6859), .C1(
        P2_U3151), .C2(n4742), .ZN(P2_U3292) );
  AOI22_X1 U8642 ( .A1(n6924), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9790), .ZN(n6861) );
  OAI21_X1 U8643 ( .B1(n6862), .B2(n9792), .A(n6861), .ZN(P1_U3349) );
  OAI222_X1 U8644 ( .A1(n6964), .A2(n6863), .B1(n9158), .B2(n6862), .C1(
        P2_U3151), .C2(n7364), .ZN(P2_U3289) );
  INV_X1 U8645 ( .A(n6864), .ZN(n6867) );
  AOI22_X1 U8646 ( .A1(n6937), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9790), .ZN(n6865) );
  OAI21_X1 U8647 ( .B1(n6867), .B2(n9792), .A(n6865), .ZN(P1_U3348) );
  INV_X1 U8648 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n7019) );
  OAI222_X1 U8649 ( .A1(n6964), .A2(n7019), .B1(n9158), .B2(n6867), .C1(
        P2_U3151), .C2(n6866), .ZN(P2_U3288) );
  INV_X1 U8650 ( .A(n6868), .ZN(n6870) );
  OAI222_X1 U8651 ( .A1(n6964), .A2(n6869), .B1(n9158), .B2(n6870), .C1(
        P2_U3151), .C2(n7750), .ZN(P2_U3287) );
  INV_X1 U8652 ( .A(n9370), .ZN(n6871) );
  OAI222_X1 U8653 ( .A1(n6871), .A2(P1_U3086), .B1(n9792), .B2(n6870), .C1(
        n7166), .C2(n8565), .ZN(P1_U3347) );
  NOR2_X1 U8654 ( .A1(n9422), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8655 ( .A(n6872), .ZN(n6881) );
  AOI22_X1 U8656 ( .A1(n7828), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9156), .ZN(n6873) );
  OAI21_X1 U8657 ( .B1(n6881), .B2(n9158), .A(n6873), .ZN(P2_U3286) );
  AOI21_X1 U8658 ( .B1(n8191), .B2(n6875), .A(n6874), .ZN(n6876) );
  XNOR2_X1 U8659 ( .A(n6876), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6880) );
  INV_X1 U8660 ( .A(n6877), .ZN(n6879) );
  AOI22_X1 U8661 ( .A1(n9422), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n6878) );
  OAI21_X1 U8662 ( .B1(n6880), .B2(n6879), .A(n6878), .ZN(P1_U3243) );
  INV_X1 U8663 ( .A(n9400), .ZN(n6882) );
  OAI222_X1 U8664 ( .A1(P1_U3086), .A2(n6882), .B1(n9792), .B2(n6881), .C1(
        n7152), .C2(n8565), .ZN(P1_U3346) );
  INV_X1 U8665 ( .A(n6883), .ZN(n6886) );
  AOI22_X1 U8666 ( .A1(n9853), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n9790), .ZN(n6884) );
  OAI21_X1 U8667 ( .B1(n6886), .B2(n9792), .A(n6884), .ZN(P1_U3345) );
  INV_X1 U8668 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6885) );
  OAI222_X1 U8669 ( .A1(n9158), .A2(n6886), .B1(n7898), .B2(P2_U3151), .C1(
        n6885), .C2(n6964), .ZN(P2_U3285) );
  INV_X1 U8670 ( .A(n6887), .ZN(n6901) );
  AOI22_X1 U8671 ( .A1(n9899), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9790), .ZN(n6888) );
  OAI21_X1 U8672 ( .B1(n6901), .B2(n9792), .A(n6888), .ZN(P1_U3344) );
  INV_X1 U8673 ( .A(n6889), .ZN(n6894) );
  AOI22_X1 U8674 ( .A1(n9903), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9790), .ZN(n6890) );
  OAI21_X1 U8675 ( .B1(n6894), .B2(n9792), .A(n6890), .ZN(P1_U3343) );
  NAND2_X1 U8676 ( .A1(n6891), .A2(P1_U3973), .ZN(n6892) );
  OAI21_X1 U8677 ( .B1(P1_U3973), .B2(n5120), .A(n6892), .ZN(P1_U3585) );
  OAI222_X1 U8678 ( .A1(n9158), .A2(n6894), .B1(n8015), .B2(P2_U3151), .C1(
        n6893), .C2(n6964), .ZN(P2_U3283) );
  INV_X1 U8679 ( .A(n6483), .ZN(n6895) );
  NAND2_X1 U8680 ( .A1(n7010), .A2(n6895), .ZN(n6903) );
  INV_X1 U8681 ( .A(n6896), .ZN(n7958) );
  NOR3_X1 U8682 ( .A1(n6897), .A2(n7958), .A3(P2_U3151), .ZN(n6898) );
  AOI21_X1 U8683 ( .B1(n6903), .B2(n6899), .A(n6898), .ZN(P2_U3376) );
  OAI222_X1 U8684 ( .A1(n6964), .A2(n6902), .B1(n9158), .B2(n6901), .C1(
        P2_U3151), .C2(n6900), .ZN(P2_U3284) );
  AND2_X1 U8685 ( .A1(n6903), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8686 ( .A1(n6903), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8687 ( .A1(n6903), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8688 ( .A1(n6903), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8689 ( .A1(n6903), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8690 ( .A1(n6903), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8691 ( .A1(n6903), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8692 ( .A1(n6903), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8693 ( .A1(n6903), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8694 ( .A1(n6903), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U8695 ( .A1(n6903), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8696 ( .A1(n6903), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8697 ( .A1(n6903), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8698 ( .A1(n6903), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8699 ( .A1(n6903), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8700 ( .A1(n6903), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8701 ( .A1(n6903), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8702 ( .A1(n6903), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8703 ( .A1(n6903), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8704 ( .A1(n6903), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8705 ( .A1(n6903), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8706 ( .A1(n6903), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8707 ( .A1(n6903), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8708 ( .A1(n6903), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8709 ( .A1(n6903), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8710 ( .A1(n6903), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  INV_X1 U8711 ( .A(n6903), .ZN(n6904) );
  INV_X1 U8712 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n7048) );
  NOR2_X1 U8713 ( .A1(n6904), .A2(n7048), .ZN(P2_U3234) );
  INV_X1 U8714 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n7142) );
  NOR2_X1 U8715 ( .A1(n6904), .A2(n7142), .ZN(P2_U3242) );
  INV_X1 U8716 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n7035) );
  NOR2_X1 U8717 ( .A1(n6904), .A2(n7035), .ZN(P2_U3251) );
  INV_X1 U8718 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n7153) );
  NOR2_X1 U8719 ( .A1(n6904), .A2(n7153), .ZN(P2_U3259) );
  XNOR2_X1 U8720 ( .A(n6949), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6947) );
  NOR2_X1 U8721 ( .A1(n6948), .A2(n6947), .ZN(n6946) );
  MUX2_X1 U8722 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7617), .S(n6924), .Z(n6906)
         );
  INV_X1 U8723 ( .A(n6906), .ZN(n6907) );
  NOR2_X1 U8724 ( .A1(n6908), .A2(n6907), .ZN(n6920) );
  AOI211_X1 U8725 ( .C1(n6908), .C2(n6907), .A(n9999), .B(n6920), .ZN(n6919)
         );
  INV_X1 U8726 ( .A(n6909), .ZN(n6910) );
  XNOR2_X1 U8727 ( .A(n6949), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6944) );
  NOR2_X1 U8728 ( .A1(n6945), .A2(n6944), .ZN(n6943) );
  INV_X1 U8729 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6912) );
  MUX2_X1 U8730 ( .A(n6912), .B(P1_REG1_REG_6__SCAN_IN), .S(n6924), .Z(n6913)
         );
  NOR2_X1 U8731 ( .A1(n6914), .A2(n6913), .ZN(n6923) );
  AOI211_X1 U8732 ( .C1(n6914), .C2(n6913), .A(n9993), .B(n6923), .ZN(n6918)
         );
  INV_X1 U8733 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9808) );
  INV_X1 U8734 ( .A(n9974), .ZN(n10005) );
  NAND2_X1 U8735 ( .A1(n10005), .A2(n6924), .ZN(n6916) );
  NAND2_X1 U8736 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n6915) );
  OAI211_X1 U8737 ( .C1(n9808), .C2(n10008), .A(n6916), .B(n6915), .ZN(n6917)
         );
  OR3_X1 U8738 ( .A1(n6919), .A2(n6918), .A3(n6917), .ZN(P1_U3249) );
  XNOR2_X1 U8739 ( .A(n6937), .B(P1_REG2_REG_7__SCAN_IN), .ZN(n6932) );
  NOR2_X1 U8740 ( .A1(n6933), .A2(n6932), .ZN(n6931) );
  XNOR2_X1 U8741 ( .A(n9370), .B(P1_REG2_REG_8__SCAN_IN), .ZN(n6921) );
  NOR2_X1 U8742 ( .A1(n6922), .A2(n6921), .ZN(n9365) );
  AOI211_X1 U8743 ( .C1(n6922), .C2(n6921), .A(n9999), .B(n9365), .ZN(n6930)
         );
  AOI21_X1 U8744 ( .B1(n6924), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6923), .ZN(
        n6936) );
  XNOR2_X1 U8745 ( .A(n6937), .B(P1_REG1_REG_7__SCAN_IN), .ZN(n6935) );
  NOR2_X1 U8746 ( .A1(n6936), .A2(n6935), .ZN(n6934) );
  XNOR2_X1 U8747 ( .A(n9370), .B(P1_REG1_REG_8__SCAN_IN), .ZN(n6925) );
  NOR2_X1 U8748 ( .A1(n6926), .A2(n6925), .ZN(n9369) );
  AOI211_X1 U8749 ( .C1(n6926), .C2(n6925), .A(n9993), .B(n9369), .ZN(n6929)
         );
  INV_X1 U8750 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U8751 ( .A1(n10005), .A2(n9370), .ZN(n6927) );
  NAND2_X1 U8752 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7818) );
  OAI211_X1 U8753 ( .C1(n9817), .C2(n10008), .A(n6927), .B(n7818), .ZN(n6928)
         );
  OR3_X1 U8754 ( .A1(n6930), .A2(n6929), .A3(n6928), .ZN(P1_U3251) );
  AOI211_X1 U8755 ( .C1(n6933), .C2(n6932), .A(n9999), .B(n6931), .ZN(n6942)
         );
  AOI211_X1 U8756 ( .C1(n6936), .C2(n6935), .A(n9993), .B(n6934), .ZN(n6941)
         );
  INV_X1 U8757 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9813) );
  NAND2_X1 U8758 ( .A1(n10005), .A2(n6937), .ZN(n6939) );
  NAND2_X1 U8759 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n6938) );
  OAI211_X1 U8760 ( .C1(n9813), .C2(n10008), .A(n6939), .B(n6938), .ZN(n6940)
         );
  OR3_X1 U8761 ( .A1(n6942), .A2(n6941), .A3(n6940), .ZN(P1_U3250) );
  AOI211_X1 U8762 ( .C1(n6945), .C2(n6944), .A(n6943), .B(n9993), .ZN(n6953)
         );
  AOI211_X1 U8763 ( .C1(n6948), .C2(n6947), .A(n6946), .B(n9999), .ZN(n6952)
         );
  INV_X1 U8764 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n7174) );
  NAND2_X1 U8765 ( .A1(n10005), .A2(n6949), .ZN(n6950) );
  NAND2_X1 U8766 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n7535) );
  OAI211_X1 U8767 ( .C1(n7174), .C2(n10008), .A(n6950), .B(n7535), .ZN(n6951)
         );
  OR3_X1 U8768 ( .A1(n6953), .A2(n6952), .A3(n6951), .ZN(P1_U3248) );
  INV_X1 U8769 ( .A(n6954), .ZN(n6960) );
  AOI22_X1 U8770 ( .A1(n9919), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9790), .ZN(n6955) );
  OAI21_X1 U8771 ( .B1(n6960), .B2(n9792), .A(n6955), .ZN(P1_U3342) );
  INV_X1 U8772 ( .A(n9885), .ZN(n9292) );
  NAND2_X1 U8773 ( .A1(n9890), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7242) );
  INV_X1 U8774 ( .A(n9882), .ZN(n9288) );
  NAND2_X1 U8775 ( .A1(n9322), .A2(n9287), .ZN(n7566) );
  OAI22_X1 U8776 ( .A1(n9288), .A2(n7566), .B1(n9280), .B2(n7264), .ZN(n6956)
         );
  AOI21_X1 U8777 ( .B1(P1_REG3_REG_0__SCAN_IN), .B2(n7242), .A(n6956), .ZN(
        n6957) );
  OAI21_X1 U8778 ( .B1(n6958), .B2(n9292), .A(n6957), .ZN(P1_U3232) );
  INV_X1 U8779 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6961) );
  OAI222_X1 U8780 ( .A1(n6964), .A2(n6961), .B1(n9158), .B2(n6960), .C1(
        P2_U3151), .C2(n6959), .ZN(P2_U3282) );
  INV_X1 U8781 ( .A(n6962), .ZN(n6965) );
  OAI222_X1 U8782 ( .A1(n6964), .A2(n6963), .B1(n9158), .B2(n6965), .C1(
        P2_U3151), .C2(n10127), .ZN(P2_U3281) );
  INV_X1 U8783 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6966) );
  INV_X1 U8784 ( .A(n9407), .ZN(n9948) );
  OAI222_X1 U8785 ( .A1(n8565), .A2(n6966), .B1(n9792), .B2(n6965), .C1(n9948), 
        .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U8786 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7164) );
  INV_X1 U8787 ( .A(n7563), .ZN(n6974) );
  NAND2_X1 U8788 ( .A1(n6522), .A2(n6967), .ZN(n6968) );
  NAND3_X1 U8789 ( .A1(n7562), .A2(n6974), .A3(n6968), .ZN(n7577) );
  NAND2_X1 U8790 ( .A1(n7570), .A2(n6969), .ZN(n6971) );
  INV_X1 U8791 ( .A(n7565), .ZN(n6972) );
  OAI21_X1 U8792 ( .B1(n9723), .B2(n9636), .A(n6972), .ZN(n6973) );
  OAI211_X1 U8793 ( .C1(n6974), .C2(n7264), .A(n6973), .B(n7566), .ZN(n9732)
         );
  NAND2_X1 U8794 ( .A1(n9732), .A2(n10077), .ZN(n6975) );
  OAI21_X1 U8795 ( .B1(n10077), .B2(n7164), .A(n6975), .ZN(P1_U3453) );
  INV_X1 U8796 ( .A(n6976), .ZN(n7196) );
  AOI22_X1 U8797 ( .A1(n6977), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n9156), .ZN(n6978) );
  OAI21_X1 U8798 ( .B1(n7196), .B2(n9158), .A(n6978), .ZN(P2_U3280) );
  INV_X1 U8799 ( .A(n6981), .ZN(n6982) );
  AOI21_X1 U8800 ( .B1(n6979), .B2(n6980), .A(n6982), .ZN(n6986) );
  INV_X1 U8801 ( .A(n9324), .ZN(n6983) );
  OAI22_X1 U8802 ( .A1(n6983), .A2(n9253), .B1(n7304), .B2(n9275), .ZN(n7262)
         );
  AOI22_X1 U8803 ( .A1(n7262), .A2(n9882), .B1(n10034), .B2(n9887), .ZN(n6985)
         );
  NAND2_X1 U8804 ( .A1(n7242), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6984) );
  OAI211_X1 U8805 ( .C1(n6986), .C2(n9292), .A(n6985), .B(n6984), .ZN(P1_U3222) );
  OR2_X1 U8806 ( .A1(n7965), .A2(n10207), .ZN(n10196) );
  NAND2_X1 U8807 ( .A1(n8708), .A2(n7214), .ZN(n8327) );
  INV_X1 U8808 ( .A(n8327), .ZN(n8334) );
  OR2_X1 U8809 ( .A1(n8334), .A2(n8329), .ZN(n8478) );
  OAI21_X1 U8810 ( .B1(n10196), .B2(n10135), .A(n8478), .ZN(n6989) );
  NOR2_X1 U8811 ( .A1(n10154), .A2(n10157), .ZN(n7322) );
  NOR2_X1 U8812 ( .A1(n7214), .A2(n10210), .ZN(n6987) );
  NOR2_X1 U8813 ( .A1(n7322), .A2(n6987), .ZN(n6988) );
  NAND2_X1 U8814 ( .A1(n6989), .A2(n6988), .ZN(n9054) );
  NAND2_X1 U8815 ( .A1(n10222), .A2(n9054), .ZN(n6990) );
  OAI21_X1 U8816 ( .B1(n10222), .B2(n6109), .A(n6990), .ZN(P2_U3390) );
  NAND2_X1 U8817 ( .A1(n6992), .A2(n6991), .ZN(n6998) );
  INV_X1 U8818 ( .A(n6993), .ZN(n7004) );
  NAND2_X1 U8819 ( .A1(n6995), .A2(n6994), .ZN(n6996) );
  AOI21_X1 U8820 ( .B1(n6999), .B2(n7004), .A(n6996), .ZN(n6997) );
  AOI21_X1 U8821 ( .B1(n6998), .B2(n6997), .A(P2_U3151), .ZN(n7002) );
  INV_X1 U8822 ( .A(n7012), .ZN(n7320) );
  NAND2_X1 U8823 ( .A1(n7010), .A2(n7320), .ZN(n8512) );
  INV_X1 U8824 ( .A(n6999), .ZN(n7000) );
  NOR2_X1 U8825 ( .A1(n8512), .A2(n7000), .ZN(n7001) );
  NOR2_X1 U8826 ( .A1(n8673), .A2(P2_U3151), .ZN(n7297) );
  INV_X1 U8827 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7017) );
  OR2_X1 U8828 ( .A1(n7008), .A2(n7003), .ZN(n7007) );
  NAND2_X1 U8829 ( .A1(n7005), .A2(n7004), .ZN(n7006) );
  OR2_X1 U8830 ( .A1(n7008), .A2(n10210), .ZN(n7011) );
  NAND2_X1 U8831 ( .A1(n7011), .A2(n10149), .ZN(n8693) );
  AOI22_X1 U8832 ( .A1(n8664), .A2(n8478), .B1(n6451), .B2(n8693), .ZN(n7016)
         );
  NOR2_X1 U8833 ( .A1(n7013), .A2(n7012), .ZN(n7204) );
  INV_X1 U8834 ( .A(n7203), .ZN(n7014) );
  NAND2_X1 U8835 ( .A1(n7204), .A2(n7014), .ZN(n8676) );
  INV_X1 U8836 ( .A(n8676), .ZN(n8683) );
  NAND2_X1 U8837 ( .A1(n8683), .A2(n6107), .ZN(n7015) );
  OAI211_X1 U8838 ( .C1(n7297), .C2(n7017), .A(n7016), .B(n7015), .ZN(P2_U3172) );
  MUX2_X1 U8839 ( .A(n8518), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8705), .Z(n7194) );
  INV_X1 U8840 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10009) );
  AOI22_X1 U8841 ( .A1(n7019), .A2(keyinput119), .B1(keyinput110), .B2(n10009), 
        .ZN(n7018) );
  OAI221_X1 U8842 ( .B1(n7019), .B2(keyinput119), .C1(n10009), .C2(keyinput110), .A(n7018), .ZN(n7023) );
  XNOR2_X1 U8843 ( .A(n7020), .B(keyinput122), .ZN(n7022) );
  XNOR2_X1 U8844 ( .A(n7142), .B(keyinput115), .ZN(n7021) );
  OR3_X1 U8845 ( .A1(n7023), .A2(n7022), .A3(n7021), .ZN(n7029) );
  INV_X1 U8846 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U8847 ( .A1(n7025), .A2(keyinput116), .B1(keyinput79), .B2(n10249), 
        .ZN(n7024) );
  OAI221_X1 U8848 ( .B1(n7025), .B2(keyinput116), .C1(n10249), .C2(keyinput79), 
        .A(n7024), .ZN(n7028) );
  AOI22_X1 U8849 ( .A1(n5363), .A2(keyinput76), .B1(n5120), .B2(keyinput84), 
        .ZN(n7026) );
  OAI221_X1 U8850 ( .B1(n5363), .B2(keyinput76), .C1(n5120), .C2(keyinput84), 
        .A(n7026), .ZN(n7027) );
  NOR3_X1 U8851 ( .A1(n7029), .A2(n7028), .A3(n7027), .ZN(n7066) );
  AOI22_X1 U8852 ( .A1(n6231), .A2(keyinput65), .B1(n5178), .B2(keyinput126), 
        .ZN(n7030) );
  OAI221_X1 U8853 ( .B1(n6231), .B2(keyinput65), .C1(n5178), .C2(keyinput126), 
        .A(n7030), .ZN(n7039) );
  AOI22_X1 U8854 ( .A1(n7032), .A2(keyinput127), .B1(n7152), .B2(keyinput113), 
        .ZN(n7031) );
  OAI221_X1 U8855 ( .B1(n7032), .B2(keyinput127), .C1(n7152), .C2(keyinput113), 
        .A(n7031), .ZN(n7038) );
  AOI22_X1 U8856 ( .A1(n9770), .A2(keyinput74), .B1(keyinput69), .B2(n7164), 
        .ZN(n7033) );
  OAI221_X1 U8857 ( .B1(n9770), .B2(keyinput74), .C1(n7164), .C2(keyinput69), 
        .A(n7033), .ZN(n7037) );
  AOI22_X1 U8858 ( .A1(n9503), .A2(keyinput64), .B1(keyinput89), .B2(n7035), 
        .ZN(n7034) );
  OAI221_X1 U8859 ( .B1(n9503), .B2(keyinput64), .C1(n7035), .C2(keyinput89), 
        .A(n7034), .ZN(n7036) );
  NOR4_X1 U8860 ( .A1(n7039), .A2(n7038), .A3(n7037), .A4(n7036), .ZN(n7065)
         );
  XOR2_X1 U8861 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput100), .Z(n7043) );
  XNOR2_X1 U8862 ( .A(n9005), .B(keyinput120), .ZN(n7042) );
  XNOR2_X1 U8863 ( .A(n7040), .B(keyinput107), .ZN(n7041) );
  NOR3_X1 U8864 ( .A1(n7043), .A2(n7042), .A3(n7041), .ZN(n7046) );
  XNOR2_X1 U8865 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput97), .ZN(n7045) );
  XNOR2_X1 U8866 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput72), .ZN(n7044) );
  NAND3_X1 U8867 ( .A1(n7046), .A2(n7045), .A3(n7044), .ZN(n7051) );
  AOI22_X1 U8868 ( .A1(n7153), .A2(keyinput121), .B1(keyinput108), .B2(n6205), 
        .ZN(n7047) );
  OAI221_X1 U8869 ( .B1(n7153), .B2(keyinput121), .C1(n6205), .C2(keyinput108), 
        .A(n7047), .ZN(n7050) );
  XNOR2_X1 U8870 ( .A(n7048), .B(keyinput86), .ZN(n7049) );
  NOR3_X1 U8871 ( .A1(n7051), .A2(n7050), .A3(n7049), .ZN(n7064) );
  AOI22_X1 U8872 ( .A1(n9095), .A2(keyinput99), .B1(keyinput70), .B2(n7053), 
        .ZN(n7052) );
  OAI221_X1 U8873 ( .B1(n9095), .B2(keyinput99), .C1(n7053), .C2(keyinput70), 
        .A(n7052), .ZN(n7062) );
  XNOR2_X1 U8874 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput95), .ZN(n7057) );
  XNOR2_X1 U8875 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput103), .ZN(n7056) );
  XNOR2_X1 U8876 ( .A(P2_REG2_REG_17__SCAN_IN), .B(keyinput105), .ZN(n7055) );
  XNOR2_X1 U8877 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput117), .ZN(n7054) );
  NAND4_X1 U8878 ( .A1(n7057), .A2(n7056), .A3(n7055), .A4(n7054), .ZN(n7061)
         );
  INV_X1 U8879 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n9760) );
  XNOR2_X1 U8880 ( .A(n9760), .B(keyinput81), .ZN(n7060) );
  XNOR2_X1 U8881 ( .A(n7058), .B(keyinput66), .ZN(n7059) );
  NOR4_X1 U8882 ( .A1(n7062), .A2(n7061), .A3(n7060), .A4(n7059), .ZN(n7063)
         );
  NAND4_X1 U8883 ( .A1(n7066), .A2(n7065), .A3(n7064), .A4(n7063), .ZN(n7192)
         );
  AOI22_X1 U8884 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(keyinput77), .B1(
        P1_IR_REG_1__SCAN_IN), .B2(keyinput87), .ZN(n7067) );
  OAI221_X1 U8885 ( .B1(P1_DATAO_REG_27__SCAN_IN), .B2(keyinput77), .C1(
        P1_IR_REG_1__SCAN_IN), .C2(keyinput87), .A(n7067), .ZN(n7074) );
  AOI22_X1 U8886 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(keyinput112), .B1(
        P2_IR_REG_7__SCAN_IN), .B2(keyinput124), .ZN(n7068) );
  OAI221_X1 U8887 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(keyinput112), .C1(
        P2_IR_REG_7__SCAN_IN), .C2(keyinput124), .A(n7068), .ZN(n7073) );
  AOI22_X1 U8888 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(keyinput114), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(keyinput85), .ZN(n7069) );
  OAI221_X1 U8889 ( .B1(P2_IR_REG_2__SCAN_IN), .B2(keyinput114), .C1(
        P1_REG3_REG_0__SCAN_IN), .C2(keyinput85), .A(n7069), .ZN(n7072) );
  AOI22_X1 U8890 ( .A1(P1_RD_REG_SCAN_IN), .A2(keyinput68), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput104), .ZN(n7070) );
  OAI221_X1 U8891 ( .B1(P1_RD_REG_SCAN_IN), .B2(keyinput68), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput104), .A(n7070), .ZN(n7071) );
  NOR4_X1 U8892 ( .A1(n7074), .A2(n7073), .A3(n7072), .A4(n7071), .ZN(n7103)
         );
  AOI22_X1 U8893 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(keyinput91), .B1(
        P1_REG2_REG_10__SCAN_IN), .B2(keyinput102), .ZN(n7075) );
  OAI221_X1 U8894 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(keyinput91), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(keyinput102), .A(n7075), .ZN(n7082) );
  AOI22_X1 U8895 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(keyinput83), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput67), .ZN(n7076) );
  OAI221_X1 U8896 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(keyinput83), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput67), .A(n7076), .ZN(n7081) );
  AOI22_X1 U8897 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput101), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput109), .ZN(n7077) );
  OAI221_X1 U8898 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput101), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput109), .A(n7077), .ZN(n7080) );
  AOI22_X1 U8899 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(keyinput123), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(keyinput93), .ZN(n7078) );
  OAI221_X1 U8900 ( .B1(P2_REG0_REG_27__SCAN_IN), .B2(keyinput123), .C1(
        P2_DATAO_REG_8__SCAN_IN), .C2(keyinput93), .A(n7078), .ZN(n7079) );
  NOR4_X1 U8901 ( .A1(n7082), .A2(n7081), .A3(n7080), .A4(n7079), .ZN(n7102)
         );
  AOI22_X1 U8902 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput78), .B1(
        P1_REG3_REG_25__SCAN_IN), .B2(keyinput106), .ZN(n7083) );
  OAI221_X1 U8903 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput78), .C1(
        P1_REG3_REG_25__SCAN_IN), .C2(keyinput106), .A(n7083), .ZN(n7091) );
  AOI22_X1 U8904 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(keyinput111), .B1(
        P2_REG2_REG_22__SCAN_IN), .B2(keyinput96), .ZN(n7084) );
  OAI221_X1 U8905 ( .B1(P2_REG0_REG_3__SCAN_IN), .B2(keyinput111), .C1(
        P2_REG2_REG_22__SCAN_IN), .C2(keyinput96), .A(n7084), .ZN(n7090) );
  INV_X1 U8906 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n9058) );
  AOI22_X1 U8907 ( .A1(n9058), .A2(keyinput94), .B1(n7086), .B2(keyinput75), 
        .ZN(n7085) );
  OAI221_X1 U8908 ( .B1(n9058), .B2(keyinput94), .C1(n7086), .C2(keyinput75), 
        .A(n7085), .ZN(n7089) );
  INV_X1 U8909 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n10046) );
  AOI22_X1 U8910 ( .A1(n7155), .A2(keyinput125), .B1(n10046), .B2(keyinput88), 
        .ZN(n7087) );
  OAI221_X1 U8911 ( .B1(n7155), .B2(keyinput125), .C1(n10046), .C2(keyinput88), 
        .A(n7087), .ZN(n7088) );
  NOR4_X1 U8912 ( .A1(n7091), .A2(n7090), .A3(n7089), .A4(n7088), .ZN(n7101)
         );
  AOI22_X1 U8913 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(keyinput118), .B1(
        P2_REG0_REG_0__SCAN_IN), .B2(keyinput82), .ZN(n7092) );
  OAI221_X1 U8914 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(keyinput118), .C1(
        P2_REG0_REG_0__SCAN_IN), .C2(keyinput82), .A(n7092), .ZN(n7099) );
  AOI22_X1 U8915 ( .A1(P2_REG0_REG_24__SCAN_IN), .A2(keyinput80), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput73), .ZN(n7093) );
  OAI221_X1 U8916 ( .B1(P2_REG0_REG_24__SCAN_IN), .B2(keyinput80), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput73), .A(n7093), .ZN(n7098) );
  AOI22_X1 U8917 ( .A1(P2_REG0_REG_7__SCAN_IN), .A2(keyinput98), .B1(
        P2_IR_REG_17__SCAN_IN), .B2(keyinput92), .ZN(n7094) );
  OAI221_X1 U8918 ( .B1(P2_REG0_REG_7__SCAN_IN), .B2(keyinput98), .C1(
        P2_IR_REG_17__SCAN_IN), .C2(keyinput92), .A(n7094), .ZN(n7097) );
  AOI22_X1 U8919 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput71), .B1(
        P1_REG1_REG_16__SCAN_IN), .B2(keyinput90), .ZN(n7095) );
  OAI221_X1 U8920 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput71), .C1(
        P1_REG1_REG_16__SCAN_IN), .C2(keyinput90), .A(n7095), .ZN(n7096) );
  NOR4_X1 U8921 ( .A1(n7099), .A2(n7098), .A3(n7097), .A4(n7096), .ZN(n7100)
         );
  NAND4_X1 U8922 ( .A1(n7103), .A2(n7102), .A3(n7101), .A4(n7100), .ZN(n7191)
         );
  OAI22_X1 U8923 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput43), .B1(keyinput21), .B2(P1_REG3_REG_0__SCAN_IN), .ZN(n7104) );
  AOI221_X1 U8924 ( .B1(P1_IR_REG_23__SCAN_IN), .B2(keyinput43), .C1(
        P1_REG3_REG_0__SCAN_IN), .C2(keyinput21), .A(n7104), .ZN(n7111) );
  OAI22_X1 U8925 ( .A1(P1_REG0_REG_28__SCAN_IN), .A2(keyinput63), .B1(
        P2_D_REG_31__SCAN_IN), .B2(keyinput22), .ZN(n7105) );
  AOI221_X1 U8926 ( .B1(P1_REG0_REG_28__SCAN_IN), .B2(keyinput63), .C1(
        keyinput22), .C2(P2_D_REG_31__SCAN_IN), .A(n7105), .ZN(n7110) );
  OAI22_X1 U8927 ( .A1(P2_D_REG_14__SCAN_IN), .A2(keyinput25), .B1(keyinput1), 
        .B2(P2_REG0_REG_11__SCAN_IN), .ZN(n7106) );
  AOI221_X1 U8928 ( .B1(P2_D_REG_14__SCAN_IN), .B2(keyinput25), .C1(
        P2_REG0_REG_11__SCAN_IN), .C2(keyinput1), .A(n7106), .ZN(n7109) );
  OAI22_X1 U8929 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(keyinput23), .B1(
        P2_REG3_REG_27__SCAN_IN), .B2(keyinput9), .ZN(n7107) );
  AOI221_X1 U8930 ( .B1(P1_IR_REG_1__SCAN_IN), .B2(keyinput23), .C1(keyinput9), 
        .C2(P2_REG3_REG_27__SCAN_IN), .A(n7107), .ZN(n7108) );
  NAND4_X1 U8931 ( .A1(n7111), .A2(n7110), .A3(n7109), .A4(n7108), .ZN(n7139)
         );
  OAI22_X1 U8932 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(keyinput52), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput14), .ZN(n7112) );
  AOI221_X1 U8933 ( .B1(P2_IR_REG_18__SCAN_IN), .B2(keyinput52), .C1(
        keyinput14), .C2(P2_REG3_REG_3__SCAN_IN), .A(n7112), .ZN(n7119) );
  OAI22_X1 U8934 ( .A1(P2_REG0_REG_27__SCAN_IN), .A2(keyinput59), .B1(
        P2_REG0_REG_24__SCAN_IN), .B2(keyinput16), .ZN(n7113) );
  AOI221_X1 U8935 ( .B1(P2_REG0_REG_27__SCAN_IN), .B2(keyinput59), .C1(
        keyinput16), .C2(P2_REG0_REG_24__SCAN_IN), .A(n7113), .ZN(n7118) );
  OAI22_X1 U8936 ( .A1(SI_24_), .A2(keyinput11), .B1(keyinput35), .B2(
        P2_REG0_REG_23__SCAN_IN), .ZN(n7114) );
  AOI221_X1 U8937 ( .B1(SI_24_), .B2(keyinput11), .C1(P2_REG0_REG_23__SCAN_IN), 
        .C2(keyinput35), .A(n7114), .ZN(n7117) );
  OAI22_X1 U8938 ( .A1(P1_REG2_REG_28__SCAN_IN), .A2(keyinput19), .B1(
        keyinput34), .B2(P2_REG0_REG_7__SCAN_IN), .ZN(n7115) );
  AOI221_X1 U8939 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(keyinput19), .C1(
        P2_REG0_REG_7__SCAN_IN), .C2(keyinput34), .A(n7115), .ZN(n7116) );
  NAND4_X1 U8940 ( .A1(n7119), .A2(n7118), .A3(n7117), .A4(n7116), .ZN(n7138)
         );
  OAI22_X1 U8941 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(keyinput44), .B1(SI_30_), 
        .B2(keyinput6), .ZN(n7120) );
  AOI221_X1 U8942 ( .B1(P2_REG3_REG_9__SCAN_IN), .B2(keyinput44), .C1(
        keyinput6), .C2(SI_30_), .A(n7120), .ZN(n7127) );
  OAI22_X1 U8943 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(keyinput33), .B1(
        P1_ADDR_REG_18__SCAN_IN), .B2(keyinput46), .ZN(n7121) );
  AOI221_X1 U8944 ( .B1(P2_IR_REG_6__SCAN_IN), .B2(keyinput33), .C1(keyinput46), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n7121), .ZN(n7126) );
  OAI22_X1 U8945 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(keyinput55), .B1(
        keyinput12), .B2(P1_REG1_REG_31__SCAN_IN), .ZN(n7122) );
  AOI221_X1 U8946 ( .B1(P1_DATAO_REG_7__SCAN_IN), .B2(keyinput55), .C1(
        P1_REG1_REG_31__SCAN_IN), .C2(keyinput12), .A(n7122), .ZN(n7125) );
  OAI22_X1 U8947 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(keyinput8), .B1(keyinput0), 
        .B2(P1_REG2_REG_24__SCAN_IN), .ZN(n7123) );
  AOI221_X1 U8948 ( .B1(P1_IR_REG_26__SCAN_IN), .B2(keyinput8), .C1(
        P1_REG2_REG_24__SCAN_IN), .C2(keyinput0), .A(n7123), .ZN(n7124) );
  NAND4_X1 U8949 ( .A1(n7127), .A2(n7126), .A3(n7125), .A4(n7124), .ZN(n7137)
         );
  OAI22_X1 U8950 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(keyinput39), .B1(
        P2_REG1_REG_26__SCAN_IN), .B2(keyinput56), .ZN(n7128) );
  AOI221_X1 U8951 ( .B1(P1_IR_REG_28__SCAN_IN), .B2(keyinput39), .C1(
        keyinput56), .C2(P2_REG1_REG_26__SCAN_IN), .A(n7128), .ZN(n7135) );
  OAI22_X1 U8952 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(keyinput58), .B1(keyinput13), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n7129) );
  AOI221_X1 U8953 ( .B1(P1_IR_REG_9__SCAN_IN), .B2(keyinput58), .C1(
        P1_DATAO_REG_27__SCAN_IN), .C2(keyinput13), .A(n7129), .ZN(n7134) );
  OAI22_X1 U8954 ( .A1(P2_REG0_REG_3__SCAN_IN), .A2(keyinput47), .B1(
        P1_ADDR_REG_0__SCAN_IN), .B2(keyinput15), .ZN(n7130) );
  AOI221_X1 U8955 ( .B1(P2_REG0_REG_3__SCAN_IN), .B2(keyinput47), .C1(
        keyinput15), .C2(P1_ADDR_REG_0__SCAN_IN), .A(n7130), .ZN(n7133) );
  OAI22_X1 U8956 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(keyinput38), .B1(
        P2_IR_REG_2__SCAN_IN), .B2(keyinput50), .ZN(n7131) );
  AOI221_X1 U8957 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(keyinput38), .C1(
        keyinput50), .C2(P2_IR_REG_2__SCAN_IN), .A(n7131), .ZN(n7132) );
  NAND4_X1 U8958 ( .A1(n7135), .A2(n7134), .A3(n7133), .A4(n7132), .ZN(n7136)
         );
  NOR4_X1 U8959 ( .A1(n7139), .A2(n7138), .A3(n7137), .A4(n7136), .ZN(n7190)
         );
  AOI22_X1 U8960 ( .A1(n9719), .A2(keyinput26), .B1(keyinput7), .B2(n10022), 
        .ZN(n7140) );
  OAI221_X1 U8961 ( .B1(n9719), .B2(keyinput26), .C1(n10022), .C2(keyinput7), 
        .A(n7140), .ZN(n7149) );
  AOI22_X1 U8962 ( .A1(n5120), .A2(keyinput20), .B1(n7142), .B2(keyinput51), 
        .ZN(n7141) );
  OAI221_X1 U8963 ( .B1(n5120), .B2(keyinput20), .C1(n7142), .C2(keyinput51), 
        .A(n7141), .ZN(n7148) );
  AOI22_X1 U8964 ( .A1(n9770), .A2(keyinput10), .B1(keyinput60), .B2(n5402), 
        .ZN(n7143) );
  OAI221_X1 U8965 ( .B1(n9770), .B2(keyinput10), .C1(n5402), .C2(keyinput60), 
        .A(n7143), .ZN(n7147) );
  XOR2_X1 U8966 ( .A(n6109), .B(keyinput18), .Z(n7145) );
  XNOR2_X1 U8967 ( .A(SI_4_), .B(keyinput2), .ZN(n7144) );
  NAND2_X1 U8968 ( .A1(n7145), .A2(n7144), .ZN(n7146) );
  NOR4_X1 U8969 ( .A1(n7149), .A2(n7148), .A3(n7147), .A4(n7146), .ZN(n7188)
         );
  AOI22_X1 U8970 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(keyinput27), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(keyinput45), .ZN(n7150) );
  OAI221_X1 U8971 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(keyinput27), .C1(
        P1_DATAO_REG_10__SCAN_IN), .C2(keyinput45), .A(n7150), .ZN(n7161) );
  AOI22_X1 U8972 ( .A1(n7153), .A2(keyinput57), .B1(n7152), .B2(keyinput49), 
        .ZN(n7151) );
  OAI221_X1 U8973 ( .B1(n7153), .B2(keyinput57), .C1(n7152), .C2(keyinput49), 
        .A(n7151), .ZN(n7160) );
  AOI22_X1 U8974 ( .A1(n7155), .A2(keyinput61), .B1(n9760), .B2(keyinput17), 
        .ZN(n7154) );
  OAI221_X1 U8975 ( .B1(n7155), .B2(keyinput61), .C1(n9760), .C2(keyinput17), 
        .A(n7154), .ZN(n7159) );
  XNOR2_X1 U8976 ( .A(P1_REG3_REG_1__SCAN_IN), .B(keyinput36), .ZN(n7157) );
  XNOR2_X1 U8977 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput40), .ZN(n7156) );
  NAND2_X1 U8978 ( .A1(n7157), .A2(n7156), .ZN(n7158) );
  NOR4_X1 U8979 ( .A1(n7161), .A2(n7160), .A3(n7159), .A4(n7158), .ZN(n7187)
         );
  AOI22_X1 U8980 ( .A1(n9221), .A2(keyinput42), .B1(keyinput30), .B2(n9058), 
        .ZN(n7162) );
  OAI221_X1 U8981 ( .B1(n9221), .B2(keyinput42), .C1(n9058), .C2(keyinput30), 
        .A(n7162), .ZN(n7172) );
  AOI22_X1 U8982 ( .A1(n7164), .A2(keyinput5), .B1(keyinput37), .B2(n10148), 
        .ZN(n7163) );
  OAI221_X1 U8983 ( .B1(n7164), .B2(keyinput5), .C1(n10148), .C2(keyinput37), 
        .A(n7163), .ZN(n7171) );
  AOI22_X1 U8984 ( .A1(n8892), .A2(keyinput32), .B1(n7166), .B2(keyinput29), 
        .ZN(n7165) );
  OAI221_X1 U8985 ( .B1(n8892), .B2(keyinput32), .C1(n7166), .C2(keyinput29), 
        .A(n7165), .ZN(n7170) );
  XNOR2_X1 U8986 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput28), .ZN(n7168) );
  XNOR2_X1 U8987 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput31), .ZN(n7167) );
  NAND2_X1 U8988 ( .A1(n7168), .A2(n7167), .ZN(n7169) );
  NOR4_X1 U8989 ( .A1(n7172), .A2(n7171), .A3(n7170), .A4(n7169), .ZN(n7186)
         );
  AOI22_X1 U8990 ( .A1(n8962), .A2(keyinput41), .B1(keyinput54), .B2(n7174), 
        .ZN(n7173) );
  OAI221_X1 U8991 ( .B1(n8962), .B2(keyinput41), .C1(n7174), .C2(keyinput54), 
        .A(n7173), .ZN(n7184) );
  AOI22_X1 U8992 ( .A1(n5178), .A2(keyinput62), .B1(n10046), .B2(keyinput24), 
        .ZN(n7175) );
  OAI221_X1 U8993 ( .B1(n5178), .B2(keyinput62), .C1(n10046), .C2(keyinput24), 
        .A(n7175), .ZN(n7183) );
  INV_X1 U8994 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7178) );
  AOI22_X1 U8995 ( .A1(n7178), .A2(keyinput48), .B1(n7177), .B2(keyinput3), 
        .ZN(n7176) );
  OAI221_X1 U8996 ( .B1(n7178), .B2(keyinput48), .C1(n7177), .C2(keyinput3), 
        .A(n7176), .ZN(n7182) );
  XNOR2_X1 U8997 ( .A(P1_RD_REG_SCAN_IN), .B(keyinput4), .ZN(n7180) );
  XNOR2_X1 U8998 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput53), .ZN(n7179) );
  NAND2_X1 U8999 ( .A1(n7180), .A2(n7179), .ZN(n7181) );
  NOR4_X1 U9000 ( .A1(n7184), .A2(n7183), .A3(n7182), .A4(n7181), .ZN(n7185)
         );
  AND4_X1 U9001 ( .A1(n7188), .A2(n7187), .A3(n7186), .A4(n7185), .ZN(n7189)
         );
  OAI211_X1 U9002 ( .C1(n7192), .C2(n7191), .A(n7190), .B(n7189), .ZN(n7193)
         );
  XNOR2_X1 U9003 ( .A(n7194), .B(n7193), .ZN(P2_U3505) );
  INV_X1 U9004 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7195) );
  OAI222_X1 U9005 ( .A1(n9409), .A2(P1_U3086), .B1(n9792), .B2(n7196), .C1(
        n7195), .C2(n8565), .ZN(P1_U3340) );
  INV_X1 U9006 ( .A(n7197), .ZN(n7201) );
  AOI22_X1 U9007 ( .A1(n7198), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9156), .ZN(n7199) );
  OAI21_X1 U9008 ( .B1(n7201), .B2(n9158), .A(n7199), .ZN(P2_U3279) );
  NAND2_X1 U9009 ( .A1(n9323), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7200) );
  OAI21_X1 U9010 ( .B1(n9196), .B2(n9323), .A(n7200), .ZN(P1_U3583) );
  OAI222_X1 U9011 ( .A1(n8565), .A2(n7202), .B1(n9792), .B2(n7201), .C1(
        P1_U3086), .C2(n9973), .ZN(P1_U3339) );
  INV_X1 U9012 ( .A(n8673), .ZN(n8685) );
  NAND2_X1 U9013 ( .A1(P2_U3151), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n7248) );
  INV_X1 U9014 ( .A(n7248), .ZN(n7206) );
  OAI22_X1 U9015 ( .A1(n8681), .A2(n6129), .B1(n7482), .B2(n8676), .ZN(n7205)
         );
  AOI211_X1 U9016 ( .C1(n10139), .C2(n8693), .A(n7206), .B(n7205), .ZN(n7224)
         );
  NAND2_X1 U9017 ( .A1(n8326), .A2(n7207), .ZN(n7208) );
  NAND2_X1 U9018 ( .A1(n7211), .A2(n10154), .ZN(n7218) );
  NAND2_X1 U9019 ( .A1(n7212), .A2(n7218), .ZN(n7291) );
  INV_X1 U9020 ( .A(n7291), .ZN(n7217) );
  NAND2_X1 U9021 ( .A1(n8558), .A2(n7214), .ZN(n7215) );
  NAND2_X1 U9022 ( .A1(n7216), .A2(n7215), .ZN(n7290) );
  NAND2_X1 U9023 ( .A1(n7217), .A2(n7290), .ZN(n7293) );
  XNOR2_X1 U9024 ( .A(n7219), .B(n10131), .ZN(n7229) );
  NAND2_X1 U9025 ( .A1(n7228), .A2(n7229), .ZN(n7227) );
  NAND2_X1 U9026 ( .A1(n7219), .A2(n6129), .ZN(n7220) );
  AND2_X2 U9027 ( .A1(n7227), .A2(n7220), .ZN(n7222) );
  XNOR2_X1 U9028 ( .A(n7213), .B(n10139), .ZN(n7330) );
  OAI211_X1 U9029 ( .C1(n7222), .C2(n7221), .A(n7333), .B(n8664), .ZN(n7223)
         );
  OAI211_X1 U9030 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8685), .A(n7224), .B(
        n7223), .ZN(P2_U3158) );
  INV_X1 U9031 ( .A(n8693), .ZN(n8670) );
  OAI22_X1 U9032 ( .A1(n10154), .A2(n8681), .B1(n8670), .B2(n7225), .ZN(n7226)
         );
  OAI21_X1 U9033 ( .B1(n7229), .B2(n7228), .A(n4331), .ZN(n7230) );
  NAND2_X1 U9034 ( .A1(n7230), .A2(n8664), .ZN(n7231) );
  OAI211_X1 U9035 ( .C1(n7297), .C2(n10148), .A(n7232), .B(n7231), .ZN(
        P2_U3177) );
  NAND2_X1 U9036 ( .A1(n9322), .A2(n9286), .ZN(n7234) );
  NAND2_X1 U9037 ( .A1(n9320), .A2(n9287), .ZN(n7233) );
  AND2_X1 U9038 ( .A1(n7234), .A2(n7233), .ZN(n7654) );
  OAI22_X1 U9039 ( .A1(n7654), .A2(n9288), .B1(n10050), .B2(n9280), .ZN(n7241)
         );
  INV_X1 U9040 ( .A(n7235), .ZN(n7237) );
  NAND3_X1 U9041 ( .A1(n7237), .A2(n6981), .A3(n7236), .ZN(n7238) );
  AOI21_X1 U9042 ( .B1(n7239), .B2(n7238), .A(n9292), .ZN(n7240) );
  AOI211_X1 U9043 ( .C1(P1_REG3_REG_2__SCAN_IN), .C2(n7242), .A(n7241), .B(
        n7240), .ZN(n7243) );
  INV_X1 U9044 ( .A(n7243), .ZN(P1_U3237) );
  OAI21_X1 U9045 ( .B1(n7244), .B2(P2_REG2_REG_3__SCAN_IN), .A(n7392), .ZN(
        n7247) );
  OAI21_X1 U9046 ( .B1(n7245), .B2(P2_REG1_REG_3__SCAN_IN), .A(n7397), .ZN(
        n7246) );
  AOI22_X1 U9047 ( .A1(n8764), .A2(n7247), .B1(n8777), .B2(n7246), .ZN(n7249)
         );
  OAI211_X1 U9048 ( .C1(n10128), .C2(n4742), .A(n7249), .B(n7248), .ZN(n7250)
         );
  AOI21_X1 U9049 ( .B1(n10109), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n7250), .ZN(
        n7256) );
  OAI21_X1 U9050 ( .B1(n7253), .B2(n7252), .A(n7251), .ZN(n7254) );
  NAND2_X1 U9051 ( .A1(n7254), .A2(n5610), .ZN(n7255) );
  NAND2_X1 U9052 ( .A1(n7256), .A2(n7255), .ZN(P2_U3185) );
  NAND2_X1 U9053 ( .A1(n9324), .A2(n7572), .ZN(n7257) );
  OAI21_X1 U9054 ( .B1(n7259), .B2(n7257), .A(n7303), .ZN(n10042) );
  INV_X1 U9055 ( .A(n10042), .ZN(n7265) );
  INV_X1 U9056 ( .A(n7577), .ZN(n10074) );
  XNOR2_X1 U9057 ( .A(n7259), .B(n7258), .ZN(n7260) );
  NOR2_X1 U9058 ( .A1(n7260), .A2(n9596), .ZN(n7261) );
  AOI211_X1 U9059 ( .C1(n10074), .C2(n10042), .A(n7262), .B(n7261), .ZN(n10044) );
  INV_X1 U9060 ( .A(n7649), .ZN(n7263) );
  OAI211_X1 U9061 ( .C1(n7436), .C2(n7264), .A(n7263), .B(n10058), .ZN(n10039)
         );
  OAI211_X1 U9062 ( .C1(n7265), .C2(n10069), .A(n10044), .B(n10039), .ZN(n7438) );
  INV_X2 U9063 ( .A(n10080), .ZN(n10082) );
  NAND2_X1 U9064 ( .A1(n10082), .A2(n10057), .ZN(n9726) );
  OAI22_X1 U9065 ( .A1(n9726), .A2(n7436), .B1(n10082), .B2(n6816), .ZN(n7267)
         );
  AOI21_X1 U9066 ( .B1(n7438), .B2(n10082), .A(n7267), .ZN(n7268) );
  INV_X1 U9067 ( .A(n7268), .ZN(P1_U3523) );
  OAI21_X1 U9068 ( .B1(n7271), .B2(n7270), .A(n7269), .ZN(n7277) );
  NAND2_X1 U9069 ( .A1(n9321), .A2(n9286), .ZN(n7273) );
  NAND2_X1 U9070 ( .A1(n9319), .A2(n9287), .ZN(n7272) );
  NAND2_X1 U9071 ( .A1(n7273), .A2(n7272), .ZN(n7310) );
  AOI22_X1 U9072 ( .A1(n7310), .A2(n9882), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        P1_U3086), .ZN(n7275) );
  INV_X1 U9073 ( .A(n7431), .ZN(n10025) );
  NAND2_X1 U9074 ( .A1(n9887), .A2(n10025), .ZN(n7274) );
  OAI211_X1 U9075 ( .C1(n9890), .C2(P1_REG3_REG_3__SCAN_IN), .A(n7275), .B(
        n7274), .ZN(n7276) );
  AOI21_X1 U9076 ( .B1(n7277), .B2(n9885), .A(n7276), .ZN(n7278) );
  INV_X1 U9077 ( .A(n7278), .ZN(P1_U3218) );
  NAND2_X1 U9078 ( .A1(n7279), .A2(n9885), .ZN(n7289) );
  AOI21_X1 U9079 ( .B1(n7269), .B2(n7281), .A(n7280), .ZN(n7288) );
  NAND2_X1 U9080 ( .A1(n9320), .A2(n9286), .ZN(n7283) );
  NAND2_X1 U9081 ( .A1(n9318), .A2(n9287), .ZN(n7282) );
  AND2_X1 U9082 ( .A1(n7283), .A2(n7282), .ZN(n7468) );
  OAI21_X1 U9083 ( .B1(n7468), .B2(n9288), .A(n7284), .ZN(n7286) );
  NOR2_X1 U9084 ( .A1(n9890), .A2(n7590), .ZN(n7285) );
  AOI211_X1 U9085 ( .C1(n7498), .C2(n9887), .A(n7286), .B(n7285), .ZN(n7287)
         );
  OAI21_X1 U9086 ( .B1(n7289), .B2(n7288), .A(n7287), .ZN(P1_U3230) );
  INV_X1 U9087 ( .A(n7290), .ZN(n7295) );
  INV_X1 U9088 ( .A(n7293), .ZN(n7294) );
  AOI21_X1 U9089 ( .B1(n7295), .B2(n7292), .A(n7294), .ZN(n7301) );
  OAI22_X1 U9090 ( .A1(n6452), .A2(n8681), .B1(n8670), .B2(n6106), .ZN(n7299)
         );
  NOR2_X1 U9091 ( .A1(n7297), .A2(n7296), .ZN(n7298) );
  AOI211_X1 U9092 ( .C1(n8683), .C2(n10131), .A(n7299), .B(n7298), .ZN(n7300)
         );
  OAI21_X1 U9093 ( .B1(n8688), .B2(n7301), .A(n7300), .ZN(P2_U3162) );
  NAND2_X1 U9094 ( .A1(n4461), .A2(n7436), .ZN(n7302) );
  NAND2_X1 U9095 ( .A1(n7303), .A2(n7302), .ZN(n7645) );
  NAND2_X1 U9096 ( .A1(n7645), .A2(n7652), .ZN(n7647) );
  NAND2_X1 U9097 ( .A1(n7647), .A2(n7305), .ZN(n7307) );
  NAND2_X1 U9098 ( .A1(n7307), .A2(n7306), .ZN(n7460) );
  OAI21_X1 U9099 ( .B1(n7307), .B2(n7306), .A(n7460), .ZN(n10029) );
  INV_X1 U9100 ( .A(n10029), .ZN(n7312) );
  XNOR2_X1 U9101 ( .A(n7309), .B(n7308), .ZN(n7311) );
  AOI21_X1 U9102 ( .B1(n7311), .B2(n9636), .A(n7310), .ZN(n10031) );
  OAI211_X1 U9103 ( .C1(n7648), .C2(n7431), .A(n10058), .B(n7463), .ZN(n10027)
         );
  OAI211_X1 U9104 ( .C1(n7312), .C2(n10062), .A(n10031), .B(n10027), .ZN(n7433) );
  OAI22_X1 U9105 ( .A1(n9726), .A2(n7431), .B1(n10082), .B2(n6819), .ZN(n7313)
         );
  AOI21_X1 U9106 ( .B1(n7433), .B2(n10082), .A(n7313), .ZN(n7314) );
  INV_X1 U9107 ( .A(n7314), .ZN(P1_U3525) );
  MUX2_X1 U9108 ( .A(n9150), .B(n7316), .S(n7315), .Z(n7317) );
  NAND2_X1 U9109 ( .A1(n7318), .A2(n7317), .ZN(n7319) );
  INV_X2 U9110 ( .A(n10162), .ZN(n10160) );
  OR2_X1 U9111 ( .A1(n7319), .A2(n8981), .ZN(n8949) );
  INV_X1 U9112 ( .A(n10149), .ZN(n10140) );
  AOI22_X1 U9113 ( .A1(n10138), .A2(n6451), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n10140), .ZN(n7325) );
  INV_X1 U9114 ( .A(n8478), .ZN(n7321) );
  NOR3_X1 U9115 ( .A1(n7321), .A2(n10221), .A3(n7320), .ZN(n7323) );
  OAI21_X1 U9116 ( .B1(n7323), .B2(n7322), .A(n10160), .ZN(n7324) );
  OAI211_X1 U9117 ( .C1(n6108), .C2(n10160), .A(n7325), .B(n7324), .ZN(
        P2_U3233) );
  INV_X1 U9118 ( .A(n7326), .ZN(n7329) );
  AOI22_X1 U9119 ( .A1(n8768), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9156), .ZN(n7327) );
  OAI21_X1 U9120 ( .B1(n7329), .B2(n9158), .A(n7327), .ZN(P2_U3278) );
  AOI22_X1 U9121 ( .A1(n9984), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9790), .ZN(n7328) );
  OAI21_X1 U9122 ( .B1(n7329), .B2(n9792), .A(n7328), .ZN(P1_U3338) );
  INV_X1 U9123 ( .A(n7330), .ZN(n7331) );
  XNOR2_X1 U9124 ( .A(n7213), .B(n10177), .ZN(n7334) );
  INV_X1 U9125 ( .A(n7334), .ZN(n7335) );
  INV_X1 U9126 ( .A(n7337), .ZN(n7441) );
  AOI21_X1 U9127 ( .B1(n7336), .B2(n7338), .A(n7441), .ZN(n7344) );
  NAND2_X1 U9128 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n7402) );
  INV_X1 U9129 ( .A(n7402), .ZN(n7340) );
  INV_X1 U9130 ( .A(n8707), .ZN(n7706) );
  OAI22_X1 U9131 ( .A1(n8681), .A2(n10156), .B1(n7706), .B2(n8676), .ZN(n7339)
         );
  AOI211_X1 U9132 ( .C1(n10177), .C2(n8693), .A(n7340), .B(n7339), .ZN(n7343)
         );
  INV_X1 U9133 ( .A(n7341), .ZN(n7495) );
  NAND2_X1 U9134 ( .A1(n8673), .A2(n7495), .ZN(n7342) );
  OAI211_X1 U9135 ( .C1(n7344), .C2(n8688), .A(n7343), .B(n7342), .ZN(P2_U3170) );
  INV_X1 U9136 ( .A(n7346), .ZN(n7347) );
  AOI21_X1 U9137 ( .B1(n7216), .B2(n7345), .A(n7347), .ZN(n10164) );
  NOR2_X1 U9138 ( .A1(n7349), .A2(n7348), .ZN(n7480) );
  OR2_X1 U9139 ( .A1(n7965), .A2(n7480), .ZN(n10159) );
  NAND2_X1 U9140 ( .A1(n10160), .A2(n10159), .ZN(n8988) );
  XNOR2_X1 U9141 ( .A(n7345), .B(n7350), .ZN(n7351) );
  AOI222_X1 U9142 ( .A1(n10135), .A2(n7351), .B1(n10131), .B2(n10132), .C1(
        n8708), .C2(n10130), .ZN(n10163) );
  MUX2_X1 U9143 ( .A(n7424), .B(n10163), .S(n10160), .Z(n7354) );
  AOI22_X1 U9144 ( .A1(n10138), .A2(n7352), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10140), .ZN(n7353) );
  OAI211_X1 U9145 ( .C1(n10164), .C2(n8988), .A(n7354), .B(n7353), .ZN(
        P2_U3232) );
  INV_X1 U9146 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7374) );
  OAI21_X1 U9147 ( .B1(n7357), .B2(n7356), .A(n7355), .ZN(n7358) );
  NAND2_X1 U9148 ( .A1(n7358), .A2(n5610), .ZN(n7373) );
  INV_X1 U9149 ( .A(n7359), .ZN(n7360) );
  NAND2_X1 U9150 ( .A1(n7361), .A2(n7360), .ZN(n7363) );
  OAI21_X1 U9151 ( .B1(n7378), .B2(n7363), .A(n7362), .ZN(n7371) );
  NAND2_X1 U9152 ( .A1(P2_U3151), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7523) );
  OAI21_X1 U9153 ( .B1(n10128), .B2(n7364), .A(n7523), .ZN(n7370) );
  NAND3_X1 U9154 ( .A1(n7375), .A2(n7366), .A3(n5540), .ZN(n7368) );
  AOI21_X1 U9155 ( .B1(n7368), .B2(n7367), .A(n10118), .ZN(n7369) );
  AOI211_X1 U9156 ( .C1(n8764), .C2(n7371), .A(n7370), .B(n7369), .ZN(n7372)
         );
  OAI211_X1 U9157 ( .C1(n8803), .C2(n7374), .A(n7373), .B(n7372), .ZN(P2_U3188) );
  OAI21_X1 U9158 ( .B1(n7376), .B2(P2_REG1_REG_5__SCAN_IN), .A(n7375), .ZN(
        n7382) );
  INV_X1 U9159 ( .A(n7377), .ZN(n7380) );
  INV_X1 U9160 ( .A(n7378), .ZN(n7379) );
  OAI21_X1 U9161 ( .B1(n7380), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7379), .ZN(
        n7381) );
  AOI22_X1 U9162 ( .A1(n7382), .A2(n8777), .B1(n8764), .B2(n7381), .ZN(n7383)
         );
  NAND2_X1 U9163 ( .A1(P2_U3151), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7448) );
  OAI211_X1 U9164 ( .C1(n10128), .C2(n5478), .A(n7383), .B(n7448), .ZN(n7388)
         );
  AOI211_X1 U9165 ( .C1(n7386), .C2(n7385), .A(n7406), .B(n7384), .ZN(n7387)
         );
  AOI211_X1 U9166 ( .C1(n10109), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n7388), .B(
        n7387), .ZN(n7389) );
  INV_X1 U9167 ( .A(n7389), .ZN(P2_U3187) );
  AND3_X1 U9168 ( .A1(n7392), .A2(n7391), .A3(n7390), .ZN(n7393) );
  OAI21_X1 U9169 ( .B1(n7394), .B2(n7393), .A(n8764), .ZN(n7404) );
  AND3_X1 U9170 ( .A1(n7397), .A2(n7396), .A3(n7395), .ZN(n7398) );
  OAI21_X1 U9171 ( .B1(n7399), .B2(n7398), .A(n8777), .ZN(n7403) );
  NAND2_X1 U9172 ( .A1(n10090), .A2(n7400), .ZN(n7401) );
  NAND4_X1 U9173 ( .A1(n7404), .A2(n7403), .A3(n7402), .A4(n7401), .ZN(n7410)
         );
  AOI211_X1 U9174 ( .C1(n7408), .C2(n7407), .A(n7406), .B(n7405), .ZN(n7409)
         );
  AOI211_X1 U9175 ( .C1(n10109), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7410), .B(
        n7409), .ZN(n7411) );
  INV_X1 U9176 ( .A(n7411), .ZN(P2_U3186) );
  AND2_X1 U9177 ( .A1(n7412), .A2(n10225), .ZN(n7413) );
  OAI21_X1 U9178 ( .B1(n7414), .B2(n7413), .A(n8777), .ZN(n7421) );
  INV_X1 U9179 ( .A(n7415), .ZN(n7419) );
  NAND2_X1 U9180 ( .A1(n7417), .A2(n7416), .ZN(n7418) );
  NAND3_X1 U9181 ( .A1(n5610), .A2(n7419), .A3(n7418), .ZN(n7420) );
  OAI211_X1 U9182 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n7296), .A(n7421), .B(n7420), .ZN(n7428) );
  AOI21_X1 U9183 ( .B1(n7424), .B2(n7423), .A(n7422), .ZN(n7426) );
  OAI22_X1 U9184 ( .A1(n10122), .A2(n7426), .B1(n10128), .B2(n7425), .ZN(n7427) );
  AOI211_X1 U9185 ( .C1(n10109), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n7428), .B(
        n7427), .ZN(n7429) );
  INV_X1 U9186 ( .A(n7429), .ZN(P2_U3183) );
  INV_X1 U9187 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n7430) );
  OAI22_X1 U9188 ( .A1(n9780), .A2(n7431), .B1(n10077), .B2(n7430), .ZN(n7432)
         );
  AOI21_X1 U9189 ( .B1(n7433), .B2(n10077), .A(n7432), .ZN(n7434) );
  INV_X1 U9190 ( .A(n7434), .ZN(P1_U3462) );
  INV_X1 U9191 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7435) );
  OAI22_X1 U9192 ( .A1(n9780), .A2(n7436), .B1(n10077), .B2(n7435), .ZN(n7437)
         );
  AOI21_X1 U9193 ( .B1(n7438), .B2(n10077), .A(n7437), .ZN(n7439) );
  INV_X1 U9194 ( .A(n7439), .ZN(P1_U3456) );
  INV_X1 U9195 ( .A(n7442), .ZN(n7440) );
  XNOR2_X1 U9196 ( .A(n8552), .B(n7451), .ZN(n7518) );
  XNOR2_X1 U9197 ( .A(n7518), .B(n8707), .ZN(n7444) );
  NOR3_X1 U9198 ( .A1(n7441), .A2(n7440), .A3(n7444), .ZN(n7447) );
  NAND2_X1 U9199 ( .A1(n7443), .A2(n7442), .ZN(n7445) );
  INV_X1 U9200 ( .A(n7520), .ZN(n7446) );
  OAI21_X1 U9201 ( .B1(n7447), .B2(n7446), .A(n8664), .ZN(n7453) );
  INV_X1 U9202 ( .A(n7448), .ZN(n7450) );
  OAI22_X1 U9203 ( .A1(n8681), .A2(n7482), .B1(n7676), .B2(n8676), .ZN(n7449)
         );
  AOI211_X1 U9204 ( .C1(n7451), .C2(n8693), .A(n7450), .B(n7449), .ZN(n7452)
         );
  OAI211_X1 U9205 ( .C1(n7486), .C2(n8685), .A(n7453), .B(n7452), .ZN(P2_U3167) );
  INV_X1 U9206 ( .A(n7454), .ZN(n7457) );
  AOI22_X1 U9207 ( .A1(n8798), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9156), .ZN(n7455) );
  OAI21_X1 U9208 ( .B1(n7457), .B2(n9158), .A(n7455), .ZN(P2_U3277) );
  AOI22_X1 U9209 ( .A1(n10004), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n9790), .ZN(n7456) );
  OAI21_X1 U9210 ( .B1(n7457), .B2(n9792), .A(n7456), .ZN(P1_U3337) );
  NAND2_X1 U9211 ( .A1(n7460), .A2(n7459), .ZN(n7462) );
  NAND2_X1 U9212 ( .A1(n7462), .A2(n7461), .ZN(n7501) );
  OAI21_X1 U9213 ( .B1(n7462), .B2(n7461), .A(n7501), .ZN(n7589) );
  AOI211_X1 U9214 ( .C1(n7498), .C2(n7463), .A(n9627), .B(n4590), .ZN(n7595)
         );
  NAND2_X1 U9215 ( .A1(n7465), .A2(n7464), .ZN(n7467) );
  XNOR2_X1 U9216 ( .A(n7467), .B(n7466), .ZN(n7469) );
  OAI21_X1 U9217 ( .B1(n7469), .B2(n9596), .A(n7468), .ZN(n7596) );
  AOI211_X1 U9218 ( .C1(n9723), .C2(n7589), .A(n7595), .B(n7596), .ZN(n7475)
         );
  OAI22_X1 U9219 ( .A1(n9726), .A2(n7593), .B1(n10082), .B2(n6815), .ZN(n7470)
         );
  INV_X1 U9220 ( .A(n7470), .ZN(n7471) );
  OAI21_X1 U9221 ( .B1(n7475), .B2(n10080), .A(n7471), .ZN(P1_U3526) );
  INV_X1 U9222 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7472) );
  OAI22_X1 U9223 ( .A1(n9780), .A2(n7593), .B1(n10077), .B2(n7472), .ZN(n7473)
         );
  INV_X1 U9224 ( .A(n7473), .ZN(n7474) );
  OAI21_X1 U9225 ( .B1(n7475), .B2(n10075), .A(n7474), .ZN(P1_U3465) );
  NAND2_X1 U9226 ( .A1(n7476), .A2(n7491), .ZN(n7479) );
  NAND2_X1 U9227 ( .A1(n7478), .A2(n7477), .ZN(n8479) );
  XNOR2_X1 U9228 ( .A(n7479), .B(n8479), .ZN(n10180) );
  NAND2_X1 U9229 ( .A1(n10160), .A2(n7480), .ZN(n8819) );
  INV_X1 U9230 ( .A(n7965), .ZN(n7765) );
  XNOR2_X1 U9231 ( .A(n7481), .B(n8479), .ZN(n7484) );
  OAI22_X1 U9232 ( .A1(n7676), .A2(n10157), .B1(n7482), .B2(n10155), .ZN(n7483) );
  AOI21_X1 U9233 ( .B1(n7484), .B2(n10135), .A(n7483), .ZN(n7485) );
  OAI21_X1 U9234 ( .B1(n10180), .B2(n7765), .A(n7485), .ZN(n10182) );
  NAND2_X1 U9235 ( .A1(n10182), .A2(n10160), .ZN(n7489) );
  OAI22_X1 U9236 ( .A1(n8949), .A2(n10179), .B1(n7486), .B2(n10149), .ZN(n7487) );
  AOI21_X1 U9237 ( .B1(n10162), .B2(P2_REG2_REG_5__SCAN_IN), .A(n7487), .ZN(
        n7488) );
  OAI211_X1 U9238 ( .C1(n10180), .C2(n8819), .A(n7489), .B(n7488), .ZN(
        P2_U3228) );
  NAND2_X1 U9239 ( .A1(n7491), .A2(n8361), .ZN(n8477) );
  XNOR2_X1 U9240 ( .A(n7490), .B(n8477), .ZN(n10173) );
  XOR2_X1 U9241 ( .A(n8477), .B(n7492), .Z(n7493) );
  MUX2_X1 U9242 ( .A(n7494), .B(n10174), .S(n10160), .Z(n7497) );
  AOI22_X1 U9243 ( .A1(n10138), .A2(n10177), .B1(n10140), .B2(n7495), .ZN(
        n7496) );
  OAI211_X1 U9244 ( .C1(n8988), .C2(n10173), .A(n7497), .B(n7496), .ZN(
        P2_U3229) );
  INV_X1 U9245 ( .A(n9319), .ZN(n7499) );
  NAND2_X1 U9246 ( .A1(n7501), .A2(n7500), .ZN(n7502) );
  NAND2_X1 U9247 ( .A1(n7502), .A2(n7504), .ZN(n7604) );
  OAI21_X1 U9248 ( .B1(n7502), .B2(n7504), .A(n7604), .ZN(n7576) );
  AOI211_X1 U9249 ( .C1(n7602), .C2(n7503), .A(n9627), .B(n7608), .ZN(n7584)
         );
  XNOR2_X1 U9250 ( .A(n7505), .B(n7504), .ZN(n7509) );
  NAND2_X1 U9251 ( .A1(n9319), .A2(n9286), .ZN(n7507) );
  NAND2_X1 U9252 ( .A1(n9317), .A2(n9287), .ZN(n7506) );
  NAND2_X1 U9253 ( .A1(n7507), .A2(n7506), .ZN(n7534) );
  INV_X1 U9254 ( .A(n7534), .ZN(n7508) );
  OAI21_X1 U9255 ( .B1(n7509), .B2(n9596), .A(n7508), .ZN(n7585) );
  AOI211_X1 U9256 ( .C1(n9723), .C2(n7576), .A(n7584), .B(n7585), .ZN(n7515)
         );
  OAI22_X1 U9257 ( .A1(n9780), .A2(n7582), .B1(n10077), .B2(n5699), .ZN(n7510)
         );
  INV_X1 U9258 ( .A(n7510), .ZN(n7511) );
  OAI21_X1 U9259 ( .B1(n7515), .B2(n10075), .A(n7511), .ZN(P1_U3468) );
  INV_X1 U9260 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7512) );
  OAI22_X1 U9261 ( .A1(n9726), .A2(n7582), .B1(n10082), .B2(n7512), .ZN(n7513)
         );
  INV_X1 U9262 ( .A(n7513), .ZN(n7514) );
  OAI21_X1 U9263 ( .B1(n7515), .B2(n10080), .A(n7514), .ZN(P1_U3527) );
  INV_X1 U9264 ( .A(n7516), .ZN(n7621) );
  AOI22_X1 U9265 ( .A1(n8509), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n9156), .ZN(n7517) );
  OAI21_X1 U9266 ( .B1(n7621), .B2(n9158), .A(n7517), .ZN(P2_U3276) );
  NAND2_X1 U9267 ( .A1(n7518), .A2(n7706), .ZN(n7519) );
  XNOR2_X1 U9268 ( .A(n7213), .B(n7526), .ZN(n7669) );
  XNOR2_X1 U9269 ( .A(n7669), .B(n8706), .ZN(n7521) );
  OAI211_X1 U9270 ( .C1(n7522), .C2(n7521), .A(n7672), .B(n8664), .ZN(n7528)
         );
  INV_X1 U9271 ( .A(n7523), .ZN(n7525) );
  OAI22_X1 U9272 ( .A1(n8681), .A2(n7706), .B1(n7769), .B2(n8676), .ZN(n7524)
         );
  AOI211_X1 U9273 ( .C1(n7526), .C2(n8693), .A(n7525), .B(n7524), .ZN(n7527)
         );
  OAI211_X1 U9274 ( .C1(n7703), .C2(n8685), .A(n7528), .B(n7527), .ZN(P2_U3179) );
  AND2_X1 U9275 ( .A1(n7530), .A2(n7529), .ZN(n7532) );
  OAI21_X1 U9276 ( .B1(n7533), .B2(n7532), .A(n7531), .ZN(n7539) );
  NOR2_X1 U9277 ( .A1(n9890), .A2(n7579), .ZN(n7538) );
  NAND2_X1 U9278 ( .A1(n7534), .A2(n9882), .ZN(n7536) );
  OAI211_X1 U9279 ( .C1(n7582), .C2(n9280), .A(n7536), .B(n7535), .ZN(n7537)
         );
  AOI211_X1 U9280 ( .C1(n7539), .C2(n9885), .A(n7538), .B(n7537), .ZN(n7540)
         );
  INV_X1 U9281 ( .A(n7540), .ZN(P1_U3227) );
  OAI21_X1 U9282 ( .B1(n7543), .B2(n7542), .A(n7541), .ZN(n7556) );
  AOI21_X1 U9283 ( .B1(n7546), .B2(n7545), .A(n7544), .ZN(n7547) );
  NOR2_X1 U9284 ( .A1(n7547), .A2(n10122), .ZN(n7555) );
  AOI21_X1 U9285 ( .B1(n10234), .B2(n7549), .A(n7548), .ZN(n7553) );
  AND2_X1 U9286 ( .A1(P2_U3151), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7678) );
  AOI21_X1 U9287 ( .B1(n10090), .B2(n7550), .A(n7678), .ZN(n7552) );
  NAND2_X1 U9288 ( .A1(n10109), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7551) );
  OAI211_X1 U9289 ( .C1(n7553), .C2(n10118), .A(n7552), .B(n7551), .ZN(n7554)
         );
  AOI211_X1 U9290 ( .C1(n7556), .C2(n5610), .A(n7555), .B(n7554), .ZN(n7557)
         );
  INV_X1 U9291 ( .A(n7557), .ZN(P2_U3189) );
  NAND3_X1 U9292 ( .A1(n7560), .A2(n7559), .A3(n7558), .ZN(n7561) );
  INV_X1 U9293 ( .A(n7562), .ZN(n7564) );
  NOR3_X1 U9294 ( .A1(n7565), .A2(n7564), .A3(n7563), .ZN(n7569) );
  OAI21_X1 U9295 ( .B1(n10021), .B2(n7567), .A(n7566), .ZN(n7568) );
  OAI21_X1 U9296 ( .B1(n7569), .B2(n7568), .A(n10023), .ZN(n7574) );
  OR2_X1 U9297 ( .A1(n10045), .A2(n7570), .ZN(n10038) );
  NOR2_X1 U9298 ( .A1(n10038), .A2(n9627), .ZN(n9547) );
  INV_X1 U9299 ( .A(n9629), .ZN(n10035) );
  OAI21_X1 U9300 ( .B1(n9547), .B2(n10035), .A(n7572), .ZN(n7573) );
  OAI211_X1 U9301 ( .C1(n5669), .C2(n10023), .A(n7574), .B(n7573), .ZN(
        P1_U3293) );
  NAND2_X1 U9302 ( .A1(n8705), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7575) );
  OAI21_X1 U9303 ( .B1(n8825), .B2(n8705), .A(n7575), .ZN(P2_U3520) );
  INV_X1 U9304 ( .A(n7576), .ZN(n7588) );
  AND2_X1 U9305 ( .A1(n7577), .A2(n7644), .ZN(n7578) );
  INV_X1 U9306 ( .A(n7579), .ZN(n7580) );
  INV_X1 U9307 ( .A(n10021), .ZN(n10032) );
  AOI22_X1 U9308 ( .A1(n10033), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n7580), .B2(
        n10032), .ZN(n7581) );
  OAI21_X1 U9309 ( .B1(n9629), .B2(n7582), .A(n7581), .ZN(n7583) );
  AOI21_X1 U9310 ( .B1(n7584), .B2(n10015), .A(n7583), .ZN(n7587) );
  NAND2_X1 U9311 ( .A1(n7585), .A2(n10023), .ZN(n7586) );
  OAI211_X1 U9312 ( .C1(n7588), .C2(n10020), .A(n7587), .B(n7586), .ZN(
        P1_U3288) );
  INV_X1 U9313 ( .A(n7589), .ZN(n7599) );
  INV_X1 U9314 ( .A(n7590), .ZN(n7591) );
  AOI22_X1 U9315 ( .A1(n10033), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7591), .B2(
        n10032), .ZN(n7592) );
  OAI21_X1 U9316 ( .B1(n9629), .B2(n7593), .A(n7592), .ZN(n7594) );
  AOI21_X1 U9317 ( .B1(n7595), .B2(n10015), .A(n7594), .ZN(n7598) );
  NAND2_X1 U9318 ( .A1(n7596), .A2(n10023), .ZN(n7597) );
  OAI211_X1 U9319 ( .C1(n7599), .C2(n10020), .A(n7598), .B(n7597), .ZN(
        P1_U3289) );
  INV_X1 U9320 ( .A(n7600), .ZN(n7623) );
  AOI22_X1 U9321 ( .A1(n8462), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n9156), .ZN(n7601) );
  OAI21_X1 U9322 ( .B1(n7623), .B2(n9158), .A(n7601), .ZN(P2_U3275) );
  NAND2_X1 U9323 ( .A1(n7604), .A2(n7603), .ZN(n7606) );
  NAND2_X1 U9324 ( .A1(n7633), .A2(n7605), .ZN(n7612) );
  OAI21_X1 U9325 ( .B1(n7606), .B2(n7612), .A(n7625), .ZN(n7607) );
  INV_X1 U9326 ( .A(n7607), .ZN(n10063) );
  INV_X1 U9327 ( .A(n7608), .ZN(n7609) );
  AOI21_X1 U9328 ( .B1(n10056), .B2(n7609), .A(n7627), .ZN(n10059) );
  OAI22_X1 U9329 ( .A1(n9629), .A2(n7610), .B1(n7714), .B2(n10021), .ZN(n7611)
         );
  AOI21_X1 U9330 ( .B1(n10059), .B2(n9547), .A(n7611), .ZN(n7619) );
  XNOR2_X1 U9331 ( .A(n7613), .B(n7612), .ZN(n7616) );
  NAND2_X1 U9332 ( .A1(n9318), .A2(n9286), .ZN(n7615) );
  NAND2_X1 U9333 ( .A1(n9316), .A2(n9287), .ZN(n7614) );
  NAND2_X1 U9334 ( .A1(n7615), .A2(n7614), .ZN(n7712) );
  AOI21_X1 U9335 ( .B1(n7616), .B2(n9636), .A(n7712), .ZN(n10061) );
  MUX2_X1 U9336 ( .A(n10061), .B(n7617), .S(n10033), .Z(n7618) );
  OAI211_X1 U9337 ( .C1(n10063), .C2(n10020), .A(n7619), .B(n7618), .ZN(
        P1_U3287) );
  OAI222_X1 U9338 ( .A1(P1_U3086), .A2(n9418), .B1(n9792), .B2(n7621), .C1(
        n7620), .C2(n8565), .ZN(P1_U3336) );
  INV_X1 U9339 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7622) );
  OAI222_X1 U9340 ( .A1(n7624), .A2(P1_U3086), .B1(n9792), .B2(n7623), .C1(
        n7622), .C2(n8565), .ZN(P1_U3335) );
  OAI21_X1 U9341 ( .B1(n7626), .B2(n7636), .A(n7785), .ZN(n7693) );
  INV_X1 U9342 ( .A(n7693), .ZN(n7643) );
  INV_X1 U9343 ( .A(n7627), .ZN(n7628) );
  AOI211_X1 U9344 ( .C1(n7784), .C2(n7628), .A(n9627), .B(n4351), .ZN(n7692)
         );
  INV_X1 U9345 ( .A(n7665), .ZN(n7629) );
  AOI22_X1 U9346 ( .A1(n10033), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7629), .B2(
        n10032), .ZN(n7630) );
  OAI21_X1 U9347 ( .B1(n9629), .B2(n7697), .A(n7630), .ZN(n7631) );
  AOI21_X1 U9348 ( .B1(n7692), .B2(n10015), .A(n7631), .ZN(n7642) );
  INV_X1 U9349 ( .A(n7632), .ZN(n7635) );
  OAI21_X1 U9350 ( .B1(n7635), .B2(n7634), .A(n7633), .ZN(n7796) );
  XNOR2_X1 U9351 ( .A(n7796), .B(n7636), .ZN(n7640) );
  OR2_X1 U9352 ( .A1(n7788), .A2(n9275), .ZN(n7638) );
  NAND2_X1 U9353 ( .A1(n9317), .A2(n9286), .ZN(n7637) );
  NAND2_X1 U9354 ( .A1(n7638), .A2(n7637), .ZN(n7663) );
  INV_X1 U9355 ( .A(n7663), .ZN(n7639) );
  OAI21_X1 U9356 ( .B1(n7640), .B2(n9596), .A(n7639), .ZN(n7691) );
  NAND2_X1 U9357 ( .A1(n7691), .A2(n10023), .ZN(n7641) );
  OAI211_X1 U9358 ( .C1(n7643), .C2(n10020), .A(n7642), .B(n7641), .ZN(
        P1_U3286) );
  NOR2_X1 U9359 ( .A1(n10045), .A2(n7644), .ZN(n10041) );
  OR2_X1 U9360 ( .A1(n7645), .A2(n7652), .ZN(n7646) );
  NAND2_X1 U9361 ( .A1(n7647), .A2(n7646), .ZN(n10053) );
  OAI211_X1 U9362 ( .C1(n10050), .C2(n7649), .A(n4579), .B(n10058), .ZN(n10049) );
  AOI22_X1 U9363 ( .A1(n10035), .A2(n7650), .B1(n10032), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n7651) );
  OAI21_X1 U9364 ( .B1(n10049), .B2(n10038), .A(n7651), .ZN(n7658) );
  XNOR2_X1 U9365 ( .A(n7652), .B(n7653), .ZN(n7656) );
  NAND2_X1 U9366 ( .A1(n10053), .A2(n10074), .ZN(n7655) );
  OAI211_X1 U9367 ( .C1(n7656), .C2(n9596), .A(n7655), .B(n7654), .ZN(n10051)
         );
  MUX2_X1 U9368 ( .A(n10051), .B(P1_REG2_REG_2__SCAN_IN), .S(n10045), .Z(n7657) );
  AOI211_X1 U9369 ( .C1(n10041), .C2(n10053), .A(n7658), .B(n7657), .ZN(n7659)
         );
  INV_X1 U9370 ( .A(n7659), .ZN(P1_U3291) );
  NAND2_X1 U9371 ( .A1(n7660), .A2(n7718), .ZN(n7661) );
  XOR2_X1 U9372 ( .A(n7662), .B(n7661), .Z(n7668) );
  AOI22_X1 U9373 ( .A1(n7663), .A2(n9882), .B1(P1_REG3_REG_7__SCAN_IN), .B2(
        P1_U3086), .ZN(n7664) );
  OAI21_X1 U9374 ( .B1(n9890), .B2(n7665), .A(n7664), .ZN(n7666) );
  AOI21_X1 U9375 ( .B1(n7784), .B2(n9887), .A(n7666), .ZN(n7667) );
  OAI21_X1 U9376 ( .B1(n7668), .B2(n9292), .A(n7667), .ZN(P1_U3213) );
  INV_X1 U9377 ( .A(n7669), .ZN(n7670) );
  NAND2_X1 U9378 ( .A1(n7670), .A2(n8706), .ZN(n7671) );
  XNOR2_X1 U9379 ( .A(n8552), .B(n7737), .ZN(n7770) );
  XNOR2_X1 U9380 ( .A(n7770), .B(n8704), .ZN(n7673) );
  OAI21_X1 U9381 ( .B1(n7674), .B2(n7673), .A(n7772), .ZN(n7675) );
  NAND2_X1 U9382 ( .A1(n7675), .A2(n8664), .ZN(n7680) );
  OAI22_X1 U9383 ( .A1(n8681), .A2(n7676), .B1(n7774), .B2(n8676), .ZN(n7677)
         );
  AOI211_X1 U9384 ( .C1(n7737), .C2(n8693), .A(n7678), .B(n7677), .ZN(n7679)
         );
  OAI211_X1 U9385 ( .C1(n7735), .C2(n8685), .A(n7680), .B(n7679), .ZN(P2_U3153) );
  AOI21_X1 U9386 ( .B1(n7682), .B2(n7681), .A(n10153), .ZN(n7684) );
  OAI22_X1 U9387 ( .A1(n7769), .A2(n10155), .B1(n7963), .B2(n10157), .ZN(n7683) );
  AOI21_X1 U9388 ( .B1(n7684), .B2(n4966), .A(n7683), .ZN(n10192) );
  NAND2_X1 U9389 ( .A1(n7729), .A2(n7685), .ZN(n7686) );
  XNOR2_X1 U9390 ( .A(n7686), .B(n8481), .ZN(n10195) );
  INV_X1 U9391 ( .A(n8988), .ZN(n10142) );
  NOR2_X1 U9392 ( .A1(n8949), .A2(n10193), .ZN(n7689) );
  OAI22_X1 U9393 ( .A1(n10160), .A2(n7687), .B1(n7775), .B2(n10149), .ZN(n7688) );
  AOI211_X1 U9394 ( .C1(n10195), .C2(n10142), .A(n7689), .B(n7688), .ZN(n7690)
         );
  OAI21_X1 U9395 ( .B1(n10192), .B2(n10162), .A(n7690), .ZN(P2_U3225) );
  AOI211_X1 U9396 ( .C1(n9723), .C2(n7693), .A(n7692), .B(n7691), .ZN(n7700)
         );
  INV_X1 U9397 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7694) );
  OAI22_X1 U9398 ( .A1(n9726), .A2(n7697), .B1(n10082), .B2(n7694), .ZN(n7695)
         );
  INV_X1 U9399 ( .A(n7695), .ZN(n7696) );
  OAI21_X1 U9400 ( .B1(n7700), .B2(n10080), .A(n7696), .ZN(P1_U3529) );
  OAI22_X1 U9401 ( .A1(n9780), .A2(n7697), .B1(n10077), .B2(n5725), .ZN(n7698)
         );
  INV_X1 U9402 ( .A(n7698), .ZN(n7699) );
  OAI21_X1 U9403 ( .B1(n7700), .B2(n10075), .A(n7699), .ZN(P1_U3474) );
  XNOR2_X1 U9404 ( .A(n7702), .B(n7701), .ZN(n10187) );
  OAI22_X1 U9405 ( .A1(n8949), .A2(n10184), .B1(n7703), .B2(n10149), .ZN(n7708) );
  XNOR2_X1 U9406 ( .A(n7704), .B(n8482), .ZN(n7705) );
  OAI222_X1 U9407 ( .A1(n10157), .A2(n7769), .B1(n10155), .B2(n7706), .C1(
        n7705), .C2(n10153), .ZN(n10185) );
  MUX2_X1 U9408 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n10185), .S(n10160), .Z(n7707) );
  AOI211_X1 U9409 ( .C1(n10142), .C2(n10187), .A(n7708), .B(n7707), .ZN(n7709)
         );
  INV_X1 U9410 ( .A(n7709), .ZN(P2_U3227) );
  INV_X1 U9411 ( .A(n7710), .ZN(n7725) );
  AOI22_X1 U9412 ( .A1(n8326), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9156), .ZN(n7711) );
  OAI21_X1 U9413 ( .B1(n7725), .B2(n9158), .A(n7711), .ZN(P2_U3274) );
  AOI22_X1 U9414 ( .A1(n7712), .A2(n9882), .B1(P1_REG3_REG_6__SCAN_IN), .B2(
        P1_U3086), .ZN(n7713) );
  OAI21_X1 U9415 ( .B1(n9890), .B2(n7714), .A(n7713), .ZN(n7722) );
  INV_X1 U9416 ( .A(n7660), .ZN(n7719) );
  AOI21_X1 U9417 ( .B1(n7716), .B2(n7718), .A(n7715), .ZN(n7717) );
  AOI21_X1 U9418 ( .B1(n7719), .B2(n7718), .A(n7717), .ZN(n7720) );
  NOR2_X1 U9419 ( .A1(n7720), .A2(n9292), .ZN(n7721) );
  AOI211_X1 U9420 ( .C1(n10056), .C2(n9887), .A(n7722), .B(n7721), .ZN(n7723)
         );
  INV_X1 U9421 ( .A(n7723), .ZN(P1_U3239) );
  OAI222_X1 U9422 ( .A1(n7726), .A2(P1_U3086), .B1(n9792), .B2(n7725), .C1(
        n7724), .C2(n8565), .ZN(P1_U3334) );
  NAND2_X1 U9423 ( .A1(n7727), .A2(n8483), .ZN(n7728) );
  NAND2_X1 U9424 ( .A1(n7729), .A2(n7728), .ZN(n10189) );
  XNOR2_X1 U9425 ( .A(n7730), .B(n8483), .ZN(n7731) );
  NAND2_X1 U9426 ( .A1(n7731), .A2(n10135), .ZN(n7733) );
  INV_X1 U9427 ( .A(n7774), .ZN(n8703) );
  AOI22_X1 U9428 ( .A1(n8703), .A2(n10132), .B1(n10130), .B2(n8706), .ZN(n7732) );
  OAI211_X1 U9429 ( .C1(n7765), .C2(n10189), .A(n7733), .B(n7732), .ZN(n10191)
         );
  MUX2_X1 U9430 ( .A(n10191), .B(P2_REG2_REG_7__SCAN_IN), .S(n10162), .Z(n7734) );
  INV_X1 U9431 ( .A(n7734), .ZN(n7739) );
  INV_X1 U9432 ( .A(n7735), .ZN(n7736) );
  AOI22_X1 U9433 ( .A1(n10138), .A2(n7737), .B1(n10140), .B2(n7736), .ZN(n7738) );
  OAI211_X1 U9434 ( .C1(n10189), .C2(n8819), .A(n7739), .B(n7738), .ZN(
        P2_U3226) );
  AOI21_X1 U9435 ( .B1(n7742), .B2(n7741), .A(n7740), .ZN(n7758) );
  INV_X1 U9436 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7743) );
  NOR2_X1 U9437 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7743), .ZN(n7778) );
  INV_X1 U9438 ( .A(n7778), .ZN(n7749) );
  OAI21_X1 U9439 ( .B1(n7746), .B2(n7745), .A(n7744), .ZN(n7747) );
  NAND2_X1 U9440 ( .A1(n5610), .A2(n7747), .ZN(n7748) );
  OAI211_X1 U9441 ( .C1(n10128), .C2(n7750), .A(n7749), .B(n7748), .ZN(n7756)
         );
  AOI21_X1 U9442 ( .B1(n7753), .B2(n7752), .A(n7751), .ZN(n7754) );
  NOR2_X1 U9443 ( .A1(n7754), .A2(n10118), .ZN(n7755) );
  AOI211_X1 U9444 ( .C1(n10109), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7756), .B(
        n7755), .ZN(n7757) );
  OAI21_X1 U9445 ( .B1(n7758), .B2(n10122), .A(n7757), .ZN(P2_U3190) );
  OAI21_X1 U9446 ( .B1(n7760), .B2(n8487), .A(n7759), .ZN(n10200) );
  XNOR2_X1 U9447 ( .A(n7761), .B(n8487), .ZN(n7762) );
  NAND2_X1 U9448 ( .A1(n7762), .A2(n10135), .ZN(n7764) );
  AOI22_X1 U9449 ( .A1(n10132), .A2(n8068), .B1(n8703), .B2(n10130), .ZN(n7763) );
  OAI211_X1 U9450 ( .C1(n7765), .C2(n10200), .A(n7764), .B(n7763), .ZN(n10202)
         );
  NAND2_X1 U9451 ( .A1(n10202), .A2(n10160), .ZN(n7768) );
  OAI22_X1 U9452 ( .A1(n10160), .A2(n7825), .B1(n7857), .B2(n10149), .ZN(n7766) );
  AOI21_X1 U9453 ( .B1(n10138), .B2(n7861), .A(n7766), .ZN(n7767) );
  OAI211_X1 U9454 ( .C1(n10200), .C2(n8819), .A(n7768), .B(n7767), .ZN(
        P2_U3224) );
  NAND2_X1 U9455 ( .A1(n7770), .A2(n7769), .ZN(n7771) );
  XNOR2_X1 U9456 ( .A(n4342), .B(n10193), .ZN(n7849) );
  OAI21_X1 U9457 ( .B1(n7774), .B2(n4332), .A(n7852), .ZN(n7782) );
  INV_X1 U9458 ( .A(n7775), .ZN(n7777) );
  AOI22_X1 U9459 ( .A1(n7777), .A2(n8673), .B1(n8693), .B2(n7776), .ZN(n7780)
         );
  AOI21_X1 U9460 ( .B1(n8672), .B2(n8704), .A(n7778), .ZN(n7779) );
  OAI211_X1 U9461 ( .C1(n7963), .C2(n8676), .A(n7780), .B(n7779), .ZN(n7781)
         );
  AOI21_X1 U9462 ( .B1(n7782), .B2(n8664), .A(n7781), .ZN(n7783) );
  INV_X1 U9463 ( .A(n7783), .ZN(P2_U3161) );
  NAND2_X1 U9464 ( .A1(n7787), .A2(n7786), .ZN(n7911) );
  NAND2_X1 U9465 ( .A1(n7909), .A2(n7911), .ZN(n7908) );
  INV_X1 U9466 ( .A(n7788), .ZN(n9315) );
  NAND2_X1 U9467 ( .A1(n7788), .A2(n4589), .ZN(n7789) );
  NAND2_X1 U9468 ( .A1(n7908), .A2(n7789), .ZN(n7792) );
  NAND2_X1 U9469 ( .A1(n7791), .A2(n7790), .ZN(n7798) );
  OAI21_X1 U9470 ( .B1(n7792), .B2(n7798), .A(n7868), .ZN(n7841) );
  INV_X1 U9471 ( .A(n7841), .ZN(n7808) );
  INV_X1 U9472 ( .A(n7793), .ZN(n7794) );
  AOI21_X1 U9473 ( .B1(n7796), .B2(n7795), .A(n7794), .ZN(n7910) );
  OAI21_X1 U9474 ( .B1(n7910), .B2(n7911), .A(n7797), .ZN(n7799) );
  XNOR2_X1 U9475 ( .A(n7799), .B(n7798), .ZN(n7800) );
  NAND2_X1 U9476 ( .A1(n9315), .A2(n9286), .ZN(n7948) );
  OAI21_X1 U9477 ( .B1(n7800), .B2(n9596), .A(n7948), .ZN(n7839) );
  INV_X1 U9478 ( .A(n7952), .ZN(n7844) );
  INV_X1 U9479 ( .A(n7915), .ZN(n7801) );
  OAI211_X1 U9480 ( .C1(n7801), .C2(n7844), .A(n10058), .B(n7871), .ZN(n7802)
         );
  INV_X1 U9481 ( .A(n8230), .ZN(n9313) );
  NAND2_X1 U9482 ( .A1(n9313), .A2(n9287), .ZN(n7949) );
  NAND2_X1 U9483 ( .A1(n7802), .A2(n7949), .ZN(n7840) );
  NAND2_X1 U9484 ( .A1(n7840), .A2(n10015), .ZN(n7805) );
  INV_X1 U9485 ( .A(n7803), .ZN(n7951) );
  AOI22_X1 U9486 ( .A1(n10033), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7951), .B2(
        n10032), .ZN(n7804) );
  OAI211_X1 U9487 ( .C1(n7844), .C2(n9629), .A(n7805), .B(n7804), .ZN(n7806)
         );
  AOI21_X1 U9488 ( .B1(n7839), .B2(n10023), .A(n7806), .ZN(n7807) );
  OAI21_X1 U9489 ( .B1(n7808), .B2(n10020), .A(n7807), .ZN(P1_U3284) );
  INV_X1 U9490 ( .A(n7809), .ZN(n7890) );
  AOI22_X1 U9491 ( .A1(n8513), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n9156), .ZN(n7810) );
  OAI21_X1 U9492 ( .B1(n7890), .B2(n9158), .A(n7810), .ZN(P2_U3273) );
  NAND2_X1 U9493 ( .A1(n7660), .A2(n7811), .ZN(n7813) );
  AND2_X1 U9494 ( .A1(n7813), .A2(n7812), .ZN(n7941) );
  XOR2_X1 U9495 ( .A(n7939), .B(n7941), .Z(n7815) );
  NOR2_X1 U9496 ( .A1(n7815), .A2(n7814), .ZN(n7940) );
  AOI21_X1 U9497 ( .B1(n7815), .B2(n7814), .A(n7940), .ZN(n7822) );
  OR2_X1 U9498 ( .A1(n7881), .A2(n9275), .ZN(n7817) );
  NAND2_X1 U9499 ( .A1(n9316), .A2(n9286), .ZN(n7816) );
  NAND2_X1 U9500 ( .A1(n7817), .A2(n7816), .ZN(n7914) );
  NAND2_X1 U9501 ( .A1(n7914), .A2(n9882), .ZN(n7819) );
  OAI211_X1 U9502 ( .C1(n9890), .C2(n10010), .A(n7819), .B(n7818), .ZN(n7820)
         );
  AOI21_X1 U9503 ( .B1(n10012), .B2(n9887), .A(n7820), .ZN(n7821) );
  OAI21_X1 U9504 ( .B1(n7822), .B2(n9292), .A(n7821), .ZN(P1_U3221) );
  AOI21_X1 U9505 ( .B1(n7825), .B2(n7824), .A(n7823), .ZN(n7838) );
  AOI21_X1 U9506 ( .B1(n7827), .B2(n10237), .A(n7826), .ZN(n7835) );
  NOR2_X1 U9507 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6205), .ZN(n7858) );
  AOI21_X1 U9508 ( .B1(n10090), .B2(n7828), .A(n7858), .ZN(n7834) );
  OAI21_X1 U9509 ( .B1(n7831), .B2(n7830), .A(n7829), .ZN(n7832) );
  NAND2_X1 U9510 ( .A1(n5610), .A2(n7832), .ZN(n7833) );
  OAI211_X1 U9511 ( .C1(n10118), .C2(n7835), .A(n7834), .B(n7833), .ZN(n7836)
         );
  AOI21_X1 U9512 ( .B1(n10109), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7836), .ZN(
        n7837) );
  OAI21_X1 U9513 ( .B1(n7838), .B2(n10122), .A(n7837), .ZN(P2_U3191) );
  AOI211_X1 U9514 ( .C1(n9723), .C2(n7841), .A(n7840), .B(n7839), .ZN(n7847)
         );
  INV_X1 U9515 ( .A(n9726), .ZN(n8162) );
  AOI22_X1 U9516 ( .A1(n8162), .A2(n7952), .B1(n10080), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n7842) );
  OAI21_X1 U9517 ( .B1(n7847), .B2(n10080), .A(n7842), .ZN(P1_U3531) );
  INV_X1 U9518 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7843) );
  OAI22_X1 U9519 ( .A1(n7844), .A2(n9780), .B1(n10077), .B2(n7843), .ZN(n7845)
         );
  INV_X1 U9520 ( .A(n7845), .ZN(n7846) );
  OAI21_X1 U9521 ( .B1(n7847), .B2(n10075), .A(n7846), .ZN(P1_U3480) );
  INV_X1 U9522 ( .A(n7849), .ZN(n7850) );
  NAND2_X1 U9523 ( .A1(n7848), .A2(n7850), .ZN(n7851) );
  XNOR2_X1 U9524 ( .A(n4342), .B(n7861), .ZN(n8026) );
  XNOR2_X1 U9525 ( .A(n8026), .B(n7963), .ZN(n7854) );
  AOI21_X1 U9526 ( .B1(n7853), .B2(n7854), .A(n8688), .ZN(n7856) );
  INV_X1 U9527 ( .A(n7854), .ZN(n7855) );
  NAND2_X1 U9528 ( .A1(n7856), .A2(n8029), .ZN(n7866) );
  INV_X1 U9529 ( .A(n7857), .ZN(n7864) );
  NAND2_X1 U9530 ( .A1(n8672), .A2(n8703), .ZN(n7860) );
  INV_X1 U9531 ( .A(n7858), .ZN(n7859) );
  OAI211_X1 U9532 ( .C1(n8075), .C2(n8676), .A(n7860), .B(n7859), .ZN(n7863)
         );
  INV_X1 U9533 ( .A(n7861), .ZN(n10198) );
  NOR2_X1 U9534 ( .A1(n8670), .A2(n10198), .ZN(n7862) );
  AOI211_X1 U9535 ( .C1(n7864), .C2(n8673), .A(n7863), .B(n7862), .ZN(n7865)
         );
  NAND2_X1 U9536 ( .A1(n7866), .A2(n7865), .ZN(P2_U3171) );
  INV_X1 U9537 ( .A(n7881), .ZN(n9314) );
  NAND2_X1 U9538 ( .A1(n7881), .A2(n7844), .ZN(n7867) );
  OAI21_X1 U9539 ( .B1(n7870), .B2(n7869), .A(n7982), .ZN(n7933) );
  INV_X1 U9540 ( .A(n7933), .ZN(n7888) );
  INV_X1 U9541 ( .A(n9862), .ZN(n7872) );
  NOR2_X1 U9542 ( .A1(n7872), .A2(n9629), .ZN(n7875) );
  OAI22_X1 U9543 ( .A1(n10023), .A2(n7873), .B1(n9865), .B2(n10021), .ZN(n7874) );
  AOI211_X1 U9544 ( .C1(n7932), .C2(n10015), .A(n7875), .B(n7874), .ZN(n7887)
         );
  INV_X1 U9545 ( .A(n8227), .ZN(n7880) );
  AOI21_X1 U9546 ( .B1(n7878), .B2(n7877), .A(n7876), .ZN(n7879) );
  OAI21_X1 U9547 ( .B1(n7880), .B2(n7879), .A(n9636), .ZN(n7885) );
  OR2_X1 U9548 ( .A1(n7881), .A2(n9253), .ZN(n7883) );
  NAND2_X1 U9549 ( .A1(n9312), .A2(n9287), .ZN(n7882) );
  NAND2_X1 U9550 ( .A1(n7883), .A2(n7882), .ZN(n9861) );
  INV_X1 U9551 ( .A(n9861), .ZN(n7884) );
  NAND2_X1 U9552 ( .A1(n7885), .A2(n7884), .ZN(n7931) );
  NAND2_X1 U9553 ( .A1(n7931), .A2(n10023), .ZN(n7886) );
  OAI211_X1 U9554 ( .C1(n7888), .C2(n10020), .A(n7887), .B(n7886), .ZN(
        P1_U3283) );
  OAI222_X1 U9555 ( .A1(P1_U3086), .A2(n7891), .B1(n9792), .B2(n7890), .C1(
        n7889), .C2(n8565), .ZN(P1_U3333) );
  AOI21_X1 U9556 ( .B1(n4423), .B2(n7893), .A(n7892), .ZN(n7907) );
  OAI21_X1 U9557 ( .B1(n7896), .B2(n7895), .A(n7894), .ZN(n7901) );
  INV_X1 U9558 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n7897) );
  OR2_X1 U9559 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7897), .ZN(n8033) );
  OAI21_X1 U9560 ( .B1(n10128), .B2(n7898), .A(n8033), .ZN(n7900) );
  INV_X1 U9561 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n9822) );
  NOR2_X1 U9562 ( .A1(n8803), .A2(n9822), .ZN(n7899) );
  AOI211_X1 U9563 ( .C1(n5610), .C2(n7901), .A(n7900), .B(n7899), .ZN(n7906)
         );
  AOI21_X1 U9564 ( .B1(n4422), .B2(n7903), .A(n7902), .ZN(n7904) );
  OR2_X1 U9565 ( .A1(n7904), .A2(n10122), .ZN(n7905) );
  OAI211_X1 U9566 ( .C1(n7907), .C2(n10118), .A(n7906), .B(n7905), .ZN(
        P2_U3192) );
  OAI21_X1 U9567 ( .B1(n7909), .B2(n7911), .A(n7908), .ZN(n10016) );
  INV_X1 U9568 ( .A(n10016), .ZN(n7916) );
  XOR2_X1 U9569 ( .A(n7911), .B(n7910), .Z(n7912) );
  NOR2_X1 U9570 ( .A1(n7912), .A2(n9596), .ZN(n7913) );
  AOI211_X1 U9571 ( .C1(n10074), .C2(n10016), .A(n7914), .B(n7913), .ZN(n10019) );
  OAI211_X1 U9572 ( .C1(n4351), .C2(n4589), .A(n10058), .B(n7915), .ZN(n10013)
         );
  OAI211_X1 U9573 ( .C1(n7916), .C2(n10069), .A(n10019), .B(n10013), .ZN(n7921) );
  NAND2_X1 U9574 ( .A1(n7921), .A2(n10082), .ZN(n7918) );
  NAND2_X1 U9575 ( .A1(n8162), .A2(n10012), .ZN(n7917) );
  OAI211_X1 U9576 ( .C1(n10082), .C2(n5734), .A(n7918), .B(n7917), .ZN(
        P1_U3530) );
  INV_X1 U9577 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7919) );
  OAI22_X1 U9578 ( .A1(n9780), .A2(n4589), .B1(n10077), .B2(n7919), .ZN(n7920)
         );
  AOI21_X1 U9579 ( .B1(n7921), .B2(n10077), .A(n7920), .ZN(n7922) );
  INV_X1 U9580 ( .A(n7922), .ZN(P1_U3477) );
  OAI21_X1 U9581 ( .B1(n7925), .B2(n7924), .A(n7923), .ZN(n7926) );
  NAND2_X1 U9582 ( .A1(n7926), .A2(n9885), .ZN(n7930) );
  INV_X1 U9583 ( .A(n7927), .ZN(n8099) );
  INV_X1 U9584 ( .A(n9890), .ZN(n9270) );
  AOI22_X1 U9585 ( .A1(n9286), .A2(n9311), .B1(n9309), .B2(n9287), .ZN(n8097)
         );
  NAND2_X1 U9586 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n9934) );
  OAI21_X1 U9587 ( .B1(n8097), .B2(n9288), .A(n9934), .ZN(n7928) );
  AOI21_X1 U9588 ( .B1(n8099), .B2(n9270), .A(n7928), .ZN(n7929) );
  OAI211_X1 U9589 ( .C1(n4593), .C2(n9280), .A(n7930), .B(n7929), .ZN(P1_U3234) );
  AOI211_X1 U9590 ( .C1(n7933), .C2(n9723), .A(n7932), .B(n7931), .ZN(n7938)
         );
  INV_X1 U9591 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7934) );
  NOR2_X1 U9592 ( .A1(n10077), .A2(n7934), .ZN(n7935) );
  AOI21_X1 U9593 ( .B1(n9862), .B2(n5396), .A(n7935), .ZN(n7936) );
  OAI21_X1 U9594 ( .B1(n7938), .B2(n10075), .A(n7936), .ZN(P1_U3483) );
  AOI22_X1 U9595 ( .A1(n9862), .A2(n8162), .B1(n10080), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n7937) );
  OAI21_X1 U9596 ( .B1(n7938), .B2(n10080), .A(n7937), .ZN(P1_U3532) );
  INV_X1 U9597 ( .A(n7939), .ZN(n7942) );
  AOI21_X1 U9598 ( .B1(n7942), .B2(n7941), .A(n7940), .ZN(n7946) );
  XNOR2_X1 U9599 ( .A(n7944), .B(n7943), .ZN(n7945) );
  XNOR2_X1 U9600 ( .A(n7946), .B(n7945), .ZN(n7955) );
  INV_X1 U9601 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7947) );
  NOR2_X1 U9602 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7947), .ZN(n9375) );
  AOI21_X1 U9603 ( .B1(n7949), .B2(n7948), .A(n9288), .ZN(n7950) );
  AOI211_X1 U9604 ( .C1(n7951), .C2(n9270), .A(n9375), .B(n7950), .ZN(n7954)
         );
  NAND2_X1 U9605 ( .A1(n7952), .A2(n9887), .ZN(n7953) );
  OAI211_X1 U9606 ( .C1(n7955), .C2(n9292), .A(n7954), .B(n7953), .ZN(P1_U3231) );
  INV_X1 U9607 ( .A(n7956), .ZN(n7960) );
  AOI21_X1 U9608 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9790), .A(n6080), .ZN(
        n7957) );
  OAI21_X1 U9609 ( .B1(n7960), .B2(n9792), .A(n7957), .ZN(P1_U3332) );
  NAND2_X1 U9610 ( .A1(n7958), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8516) );
  NAND2_X1 U9611 ( .A1(n9156), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n7959) );
  OAI211_X1 U9612 ( .C1(n7960), .C2(n9158), .A(n8516), .B(n7959), .ZN(P2_U3272) );
  XNOR2_X1 U9613 ( .A(n8076), .B(n8068), .ZN(n8485) );
  XOR2_X1 U9614 ( .A(n7961), .B(n8485), .Z(n10208) );
  INV_X1 U9615 ( .A(n10208), .ZN(n7971) );
  XNOR2_X1 U9616 ( .A(n7962), .B(n8485), .ZN(n7967) );
  OAI22_X1 U9617 ( .A1(n8174), .A2(n10157), .B1(n7963), .B2(n10155), .ZN(n7964) );
  AOI21_X1 U9618 ( .B1(n10208), .B2(n7965), .A(n7964), .ZN(n7966) );
  OAI21_X1 U9619 ( .B1(n10153), .B2(n7967), .A(n7966), .ZN(n10205) );
  NAND2_X1 U9620 ( .A1(n10205), .A2(n10160), .ZN(n7970) );
  OAI22_X1 U9621 ( .A1(n10160), .A2(n5489), .B1(n8032), .B2(n10149), .ZN(n7968) );
  AOI21_X1 U9622 ( .B1(n10138), .B2(n8076), .A(n7968), .ZN(n7969) );
  OAI211_X1 U9623 ( .C1(n7971), .C2(n8819), .A(n7970), .B(n7969), .ZN(P2_U3223) );
  XNOR2_X1 U9624 ( .A(n7972), .B(n8486), .ZN(n10212) );
  OAI211_X1 U9625 ( .C1(n4425), .C2(n8074), .A(n10135), .B(n7973), .ZN(n7975)
         );
  AOI22_X1 U9626 ( .A1(n8068), .A2(n10130), .B1(n10132), .B2(n8700), .ZN(n7974) );
  NAND2_X1 U9627 ( .A1(n7975), .A2(n7974), .ZN(n10214) );
  NAND2_X1 U9628 ( .A1(n10214), .A2(n10160), .ZN(n7978) );
  OAI22_X1 U9629 ( .A1(n10160), .A2(n8711), .B1(n8054), .B2(n10149), .ZN(n7976) );
  AOI21_X1 U9630 ( .B1(n10138), .B2(n8057), .A(n7976), .ZN(n7977) );
  OAI211_X1 U9631 ( .C1(n8988), .C2(n10212), .A(n7978), .B(n7977), .ZN(
        P2_U3222) );
  INV_X1 U9632 ( .A(n7979), .ZN(n7997) );
  AOI22_X1 U9633 ( .A1(n7980), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9156), .ZN(n7981) );
  OAI21_X1 U9634 ( .B1(n7997), .B2(n9158), .A(n7981), .ZN(P2_U3271) );
  NAND2_X1 U9635 ( .A1(n9886), .A2(n9312), .ZN(n7985) );
  XNOR2_X1 U9636 ( .A(n8090), .B(n7991), .ZN(n8003) );
  INV_X1 U9637 ( .A(n8003), .ZN(n7995) );
  INV_X1 U9638 ( .A(n4968), .ZN(n7986) );
  AOI211_X1 U9639 ( .C1(n9872), .C2(n8234), .A(n9627), .B(n7986), .ZN(n8002)
         );
  INV_X1 U9640 ( .A(n9872), .ZN(n8092) );
  NOR2_X1 U9641 ( .A1(n8092), .A2(n9629), .ZN(n7989) );
  OAI22_X1 U9642 ( .A1(n10023), .A2(n7987), .B1(n9874), .B2(n10021), .ZN(n7988) );
  AOI211_X1 U9643 ( .C1(n8002), .C2(n10015), .A(n7989), .B(n7988), .ZN(n7994)
         );
  OAI211_X1 U9644 ( .C1(n7991), .C2(n7990), .A(n8095), .B(n9636), .ZN(n7992)
         );
  INV_X1 U9645 ( .A(n8105), .ZN(n9310) );
  AOI22_X1 U9646 ( .A1(n9310), .A2(n9287), .B1(n9286), .B2(n9312), .ZN(n9866)
         );
  NAND2_X1 U9647 ( .A1(n7992), .A2(n9866), .ZN(n8001) );
  NAND2_X1 U9648 ( .A1(n8001), .A2(n10023), .ZN(n7993) );
  OAI211_X1 U9649 ( .C1(n7995), .C2(n10020), .A(n7994), .B(n7993), .ZN(
        P1_U3281) );
  OAI222_X1 U9650 ( .A1(n7998), .A2(P1_U3086), .B1(n9792), .B2(n7997), .C1(
        n7996), .C2(n8565), .ZN(P1_U3331) );
  INV_X1 U9651 ( .A(n7999), .ZN(n8050) );
  AOI22_X1 U9652 ( .A1(n4333), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9156), .ZN(n8000) );
  OAI21_X1 U9653 ( .B1(n8050), .B2(n9158), .A(n8000), .ZN(P2_U3270) );
  AOI211_X1 U9654 ( .C1(n8003), .C2(n9723), .A(n8002), .B(n8001), .ZN(n8008)
         );
  AOI22_X1 U9655 ( .A1(n9872), .A2(n8162), .B1(n10080), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n8004) );
  OAI21_X1 U9656 ( .B1(n8008), .B2(n10080), .A(n8004), .ZN(P1_U3534) );
  INV_X1 U9657 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n8005) );
  OAI22_X1 U9658 ( .A1(n8092), .A2(n9780), .B1(n10077), .B2(n8005), .ZN(n8006)
         );
  INV_X1 U9659 ( .A(n8006), .ZN(n8007) );
  OAI21_X1 U9660 ( .B1(n8008), .B2(n10075), .A(n8007), .ZN(P1_U3489) );
  AOI21_X1 U9661 ( .B1(n4409), .B2(n8010), .A(n8009), .ZN(n8025) );
  OAI21_X1 U9662 ( .B1(n8013), .B2(n8012), .A(n8011), .ZN(n8018) );
  OR2_X1 U9663 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8014), .ZN(n8180) );
  OAI21_X1 U9664 ( .B1(n10128), .B2(n8015), .A(n8180), .ZN(n8017) );
  INV_X1 U9665 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n9797) );
  NOR2_X1 U9666 ( .A1(n8803), .A2(n9797), .ZN(n8016) );
  AOI211_X1 U9667 ( .C1(n5610), .C2(n8018), .A(n8017), .B(n8016), .ZN(n8024)
         );
  AOI21_X1 U9668 ( .B1(n8021), .B2(n8020), .A(n8019), .ZN(n8022) );
  OR2_X1 U9669 ( .A1(n8022), .A2(n10122), .ZN(n8023) );
  OAI211_X1 U9670 ( .C1(n8025), .C2(n10118), .A(n8024), .B(n8023), .ZN(
        P2_U3194) );
  INV_X1 U9671 ( .A(n8026), .ZN(n8027) );
  NAND2_X1 U9672 ( .A1(n8027), .A2(n8702), .ZN(n8028) );
  AND2_X2 U9673 ( .A1(n8029), .A2(n8028), .ZN(n8072) );
  XNOR2_X1 U9674 ( .A(n8072), .B(n8068), .ZN(n8030) );
  XNOR2_X1 U9675 ( .A(n8076), .B(n4342), .ZN(n8067) );
  NAND2_X1 U9676 ( .A1(n8030), .A2(n8067), .ZN(n8053) );
  OAI21_X1 U9677 ( .B1(n8030), .B2(n8067), .A(n8053), .ZN(n8031) );
  NAND2_X1 U9678 ( .A1(n8031), .A2(n8664), .ZN(n8039) );
  INV_X1 U9679 ( .A(n8032), .ZN(n8037) );
  NAND2_X1 U9680 ( .A1(n8672), .A2(n8702), .ZN(n8034) );
  OAI211_X1 U9681 ( .C1(n8174), .C2(n8676), .A(n8034), .B(n8033), .ZN(n8036)
         );
  INV_X1 U9682 ( .A(n8076), .ZN(n10204) );
  NOR2_X1 U9683 ( .A1(n8670), .A2(n10204), .ZN(n8035) );
  AOI211_X1 U9684 ( .C1(n8037), .C2(n8673), .A(n8036), .B(n8035), .ZN(n8038)
         );
  NAND2_X1 U9685 ( .A1(n8039), .A2(n8038), .ZN(P2_U3157) );
  INV_X1 U9686 ( .A(n8384), .ZN(n8490) );
  XNOR2_X1 U9687 ( .A(n8040), .B(n8490), .ZN(n8041) );
  OAI222_X1 U9688 ( .A1(n10157), .A2(n8182), .B1(n10155), .B2(n8174), .C1(
        n10153), .C2(n8041), .ZN(n10218) );
  INV_X1 U9689 ( .A(n10218), .ZN(n8048) );
  OAI22_X1 U9690 ( .A1(n10160), .A2(n8042), .B1(n8179), .B2(n10149), .ZN(n8046) );
  NOR2_X1 U9691 ( .A1(n8043), .A2(n8384), .ZN(n10217) );
  INV_X1 U9692 ( .A(n8044), .ZN(n10216) );
  NOR3_X1 U9693 ( .A1(n10217), .A2(n10216), .A3(n8988), .ZN(n8045) );
  AOI211_X1 U9694 ( .C1(n10138), .C2(n10220), .A(n8046), .B(n8045), .ZN(n8047)
         );
  OAI21_X1 U9695 ( .B1(n8048), .B2(n10162), .A(n8047), .ZN(P2_U3221) );
  OAI222_X1 U9696 ( .A1(n8051), .A2(P1_U3086), .B1(n9792), .B2(n8050), .C1(
        n8049), .C2(n8565), .ZN(P1_U3330) );
  XNOR2_X1 U9697 ( .A(n8074), .B(n8558), .ZN(n8173) );
  NAND2_X1 U9698 ( .A1(n8072), .A2(n8075), .ZN(n8052) );
  NAND3_X1 U9699 ( .A1(n8053), .A2(n8173), .A3(n8052), .ZN(n8172) );
  NAND2_X1 U9700 ( .A1(n8172), .A2(n8664), .ZN(n8063) );
  AOI21_X1 U9701 ( .B1(n8053), .B2(n8052), .A(n8173), .ZN(n8062) );
  INV_X1 U9702 ( .A(n8054), .ZN(n8060) );
  NAND2_X1 U9703 ( .A1(n8672), .A2(n8068), .ZN(n8056) );
  AND2_X1 U9704 ( .A1(P2_U3151), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n8713) );
  INV_X1 U9705 ( .A(n8713), .ZN(n8055) );
  OAI211_X1 U9706 ( .C1(n8386), .C2(n8676), .A(n8056), .B(n8055), .ZN(n8059)
         );
  INV_X1 U9707 ( .A(n8057), .ZN(n10211) );
  NOR2_X1 U9708 ( .A1(n8670), .A2(n10211), .ZN(n8058) );
  AOI211_X1 U9709 ( .C1(n8060), .C2(n8673), .A(n8059), .B(n8058), .ZN(n8061)
         );
  OAI21_X1 U9710 ( .B1(n8063), .B2(n8062), .A(n8061), .ZN(P2_U3176) );
  INV_X1 U9711 ( .A(n8064), .ZN(n8143) );
  AOI22_X1 U9712 ( .A1(n8065), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9156), .ZN(n8066) );
  OAI21_X1 U9713 ( .B1(n8143), .B2(n9158), .A(n8066), .ZN(P2_U3269) );
  INV_X1 U9714 ( .A(n8067), .ZN(n8069) );
  NAND2_X1 U9715 ( .A1(n8069), .A2(n8068), .ZN(n8070) );
  NAND3_X1 U9716 ( .A1(n10204), .A2(n8558), .A3(n8075), .ZN(n8073) );
  OAI211_X1 U9717 ( .C1(n8558), .C2(n8701), .A(n8074), .B(n8073), .ZN(n8079)
         );
  NAND3_X1 U9718 ( .A1(n8076), .A2(n8075), .A3(n4342), .ZN(n8077) );
  OAI211_X1 U9719 ( .C1(n8701), .C2(n4342), .A(n8486), .B(n8077), .ZN(n8078)
         );
  XNOR2_X1 U9720 ( .A(n10220), .B(n8558), .ZN(n8080) );
  NOR2_X1 U9721 ( .A1(n8080), .A2(n8700), .ZN(n8175) );
  AOI21_X1 U9722 ( .B1(n8079), .B2(n8078), .A(n8175), .ZN(n8082) );
  INV_X1 U9723 ( .A(n8080), .ZN(n8081) );
  NOR2_X1 U9724 ( .A1(n8081), .A2(n8386), .ZN(n8176) );
  XNOR2_X1 U9725 ( .A(n9143), .B(n4342), .ZN(n8148) );
  XNOR2_X1 U9726 ( .A(n8148), .B(n8977), .ZN(n8149) );
  XOR2_X1 U9727 ( .A(n8150), .B(n8149), .Z(n8088) );
  AOI22_X1 U9728 ( .A1(n8672), .A2(n8700), .B1(P2_REG3_REG_13__SCAN_IN), .B2(
        P2_U3151), .ZN(n8085) );
  NAND2_X1 U9729 ( .A1(n8683), .A2(n8518), .ZN(n8084) );
  OAI211_X1 U9730 ( .C1(n8685), .C2(n8122), .A(n8085), .B(n8084), .ZN(n8086)
         );
  AOI21_X1 U9731 ( .B1(n9143), .B2(n8693), .A(n8086), .ZN(n8087) );
  OAI21_X1 U9732 ( .B1(n8088), .B2(n8688), .A(n8087), .ZN(P2_U3174) );
  XOR2_X1 U9733 ( .A(n8127), .B(n8128), .Z(n8158) );
  INV_X1 U9734 ( .A(n8158), .ZN(n8104) );
  NAND2_X1 U9735 ( .A1(n8095), .A2(n8094), .ZN(n8096) );
  XOR2_X1 U9736 ( .A(n8127), .B(n8096), .Z(n8098) );
  OAI21_X1 U9737 ( .B1(n8098), .B2(n9596), .A(n8097), .ZN(n8156) );
  AOI211_X1 U9738 ( .C1(n8163), .C2(n4968), .A(n9627), .B(n4420), .ZN(n8157)
         );
  NAND2_X1 U9739 ( .A1(n8157), .A2(n10015), .ZN(n8101) );
  AOI22_X1 U9740 ( .A1(n10033), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8099), .B2(
        n10032), .ZN(n8100) );
  OAI211_X1 U9741 ( .C1(n4593), .C2(n9629), .A(n8101), .B(n8100), .ZN(n8102)
         );
  AOI21_X1 U9742 ( .B1(n10023), .B2(n8156), .A(n8102), .ZN(n8103) );
  OAI21_X1 U9743 ( .B1(n8104), .B2(n10020), .A(n8103), .ZN(P1_U3280) );
  OR2_X1 U9744 ( .A1(n8105), .A2(n9253), .ZN(n8107) );
  NAND2_X1 U9745 ( .A1(n9308), .A2(n9287), .ZN(n8106) );
  NAND2_X1 U9746 ( .A1(n8107), .A2(n8106), .ZN(n8132) );
  AOI22_X1 U9747 ( .A1(n8132), .A2(n9882), .B1(P1_REG3_REG_14__SCAN_IN), .B2(
        P1_U3086), .ZN(n8108) );
  OAI21_X1 U9748 ( .B1(n9890), .B2(n8135), .A(n8108), .ZN(n8116) );
  INV_X1 U9749 ( .A(n8109), .ZN(n8114) );
  AOI21_X1 U9750 ( .B1(n8113), .B2(n8111), .A(n8110), .ZN(n8112) );
  AOI211_X1 U9751 ( .C1(n8114), .C2(n8113), .A(n9292), .B(n8112), .ZN(n8115)
         );
  AOI211_X1 U9752 ( .C1(n9728), .C2(n9887), .A(n8116), .B(n8115), .ZN(n8117)
         );
  INV_X1 U9753 ( .A(n8117), .ZN(P1_U3215) );
  INV_X1 U9754 ( .A(n8981), .ZN(n8120) );
  XNOR2_X1 U9755 ( .A(n8118), .B(n8489), .ZN(n8119) );
  OAI222_X1 U9756 ( .A1(n10155), .A2(n8386), .B1(n10157), .B2(n8680), .C1(
        n8119), .C2(n10153), .ZN(n9048) );
  AOI21_X1 U9757 ( .B1(n8120), .B2(n9143), .A(n9048), .ZN(n8125) );
  XNOR2_X1 U9758 ( .A(n8121), .B(n8489), .ZN(n9146) );
  OAI22_X1 U9759 ( .A1(n10160), .A2(n10094), .B1(n8122), .B2(n10149), .ZN(
        n8123) );
  AOI21_X1 U9760 ( .B1(n9146), .B2(n10142), .A(n8123), .ZN(n8124) );
  OAI21_X1 U9761 ( .B1(n8125), .B2(n10162), .A(n8124), .ZN(P2_U3220) );
  XNOR2_X1 U9762 ( .A(n4418), .B(n8129), .ZN(n9731) );
  AOI21_X1 U9763 ( .B1(n8131), .B2(n8130), .A(n9596), .ZN(n8133) );
  AOI21_X1 U9764 ( .B1(n8133), .B2(n8203), .A(n8132), .ZN(n9730) );
  NAND2_X1 U9765 ( .A1(n10033), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n8134) );
  OAI21_X1 U9766 ( .B1(n10021), .B2(n8135), .A(n8134), .ZN(n8136) );
  AOI21_X1 U9767 ( .B1(n9728), .B2(n10035), .A(n8136), .ZN(n8139) );
  OAI21_X1 U9768 ( .B1(n4420), .B2(n8192), .A(n10058), .ZN(n8137) );
  NOR2_X1 U9769 ( .A1(n8137), .A2(n8194), .ZN(n9727) );
  NAND2_X1 U9770 ( .A1(n9727), .A2(n10015), .ZN(n8138) );
  OAI211_X1 U9771 ( .C1(n9730), .C2(n10045), .A(n8139), .B(n8138), .ZN(n8140)
         );
  INV_X1 U9772 ( .A(n8140), .ZN(n8141) );
  OAI21_X1 U9773 ( .B1(n9731), .B2(n10020), .A(n8141), .ZN(P1_U3279) );
  OAI222_X1 U9774 ( .A1(n8144), .A2(P1_U3086), .B1(n9792), .B2(n8143), .C1(
        n8142), .C2(n8565), .ZN(P1_U3329) );
  INV_X1 U9775 ( .A(n8145), .ZN(n8190) );
  AOI21_X1 U9776 ( .B1(n9156), .B2(P1_DATAO_REG_27__SCAN_IN), .A(n8146), .ZN(
        n8147) );
  OAI21_X1 U9777 ( .B1(n8190), .B2(n9158), .A(n8147), .ZN(P2_U3268) );
  XNOR2_X1 U9778 ( .A(n8982), .B(n4342), .ZN(n8519) );
  XNOR2_X1 U9779 ( .A(n8519), .B(n8518), .ZN(n8520) );
  XOR2_X1 U9780 ( .A(n8521), .B(n8520), .Z(n8155) );
  INV_X1 U9781 ( .A(n8982), .ZN(n9136) );
  AOI22_X1 U9782 ( .A1(n8683), .A2(n8978), .B1(P2_REG3_REG_14__SCAN_IN), .B2(
        P2_U3151), .ZN(n8152) );
  NAND2_X1 U9783 ( .A1(n8672), .A2(n8977), .ZN(n8151) );
  OAI211_X1 U9784 ( .C1(n8980), .C2(n8685), .A(n8152), .B(n8151), .ZN(n8153)
         );
  AOI21_X1 U9785 ( .B1(n9136), .B2(n8693), .A(n8153), .ZN(n8154) );
  OAI21_X1 U9786 ( .B1(n8155), .B2(n8688), .A(n8154), .ZN(P2_U3155) );
  AOI211_X1 U9787 ( .C1(n8158), .C2(n9723), .A(n8157), .B(n8156), .ZN(n8165)
         );
  INV_X1 U9788 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n8159) );
  NOR2_X1 U9789 ( .A1(n10077), .A2(n8159), .ZN(n8160) );
  AOI21_X1 U9790 ( .B1(n8163), .B2(n5396), .A(n8160), .ZN(n8161) );
  OAI21_X1 U9791 ( .B1(n8165), .B2(n10075), .A(n8161), .ZN(P1_U3492) );
  AOI22_X1 U9792 ( .A1(n8163), .A2(n8162), .B1(n10080), .B2(
        P1_REG1_REG_13__SCAN_IN), .ZN(n8164) );
  OAI21_X1 U9793 ( .B1(n8165), .B2(n10080), .A(n8164), .ZN(P1_U3535) );
  AOI21_X1 U9794 ( .B1(n8167), .B2(n8166), .A(n4412), .ZN(n8171) );
  OAI22_X1 U9795 ( .A1(n8193), .A2(n9253), .B1(n9240), .B2(n9275), .ZN(n8206)
         );
  NAND2_X1 U9796 ( .A1(n8206), .A2(n9882), .ZN(n8168) );
  NAND2_X1 U9797 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9961) );
  OAI211_X1 U9798 ( .C1(n9890), .C2(n8198), .A(n8168), .B(n9961), .ZN(n8169)
         );
  AOI21_X1 U9799 ( .B1(n8274), .B2(n9887), .A(n8169), .ZN(n8170) );
  OAI21_X1 U9800 ( .B1(n8171), .B2(n9292), .A(n8170), .ZN(P1_U3241) );
  OAI21_X1 U9801 ( .B1(n8174), .B2(n8173), .A(n8172), .ZN(n8178) );
  NOR2_X1 U9802 ( .A1(n8176), .A2(n8175), .ZN(n8177) );
  XNOR2_X1 U9803 ( .A(n8178), .B(n8177), .ZN(n8188) );
  INV_X1 U9804 ( .A(n8179), .ZN(n8186) );
  NAND2_X1 U9805 ( .A1(n8672), .A2(n8701), .ZN(n8181) );
  OAI211_X1 U9806 ( .C1(n8182), .C2(n8676), .A(n8181), .B(n8180), .ZN(n8185)
         );
  INV_X1 U9807 ( .A(n10220), .ZN(n8183) );
  NOR2_X1 U9808 ( .A1(n8183), .A2(n8670), .ZN(n8184) );
  AOI211_X1 U9809 ( .C1(n8186), .C2(n8673), .A(n8185), .B(n8184), .ZN(n8187)
         );
  OAI21_X1 U9810 ( .B1(n8188), .B2(n8688), .A(n8187), .ZN(P2_U3164) );
  OAI222_X1 U9811 ( .A1(P1_U3086), .A2(n8191), .B1(n9792), .B2(n8190), .C1(
        n8189), .C2(n8565), .ZN(P1_U3328) );
  XNOR2_X1 U9812 ( .A(n8276), .B(n8204), .ZN(n9724) );
  INV_X1 U9813 ( .A(n9724), .ZN(n8211) );
  INV_X1 U9814 ( .A(n8194), .ZN(n8197) );
  INV_X1 U9815 ( .A(n8195), .ZN(n8196) );
  AOI211_X1 U9816 ( .C1(n8274), .C2(n8197), .A(n9627), .B(n8196), .ZN(n9722)
         );
  NOR2_X1 U9817 ( .A1(n9781), .A2(n9629), .ZN(n8201) );
  OAI22_X1 U9818 ( .A1(n10023), .A2(n8199), .B1(n8198), .B2(n10021), .ZN(n8200) );
  AOI211_X1 U9819 ( .C1(n9722), .C2(n10015), .A(n8201), .B(n8200), .ZN(n8210)
         );
  NAND2_X1 U9820 ( .A1(n8203), .A2(n8202), .ZN(n8205) );
  XNOR2_X1 U9821 ( .A(n8205), .B(n8204), .ZN(n8208) );
  INV_X1 U9822 ( .A(n8206), .ZN(n8207) );
  OAI21_X1 U9823 ( .B1(n8208), .B2(n9596), .A(n8207), .ZN(n9721) );
  NAND2_X1 U9824 ( .A1(n9721), .A2(n10023), .ZN(n8209) );
  OAI211_X1 U9825 ( .C1(n8211), .C2(n10020), .A(n8210), .B(n8209), .ZN(
        P1_U3278) );
  INV_X1 U9826 ( .A(n8212), .ZN(n8216) );
  NAND2_X1 U9827 ( .A1(n9156), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8213) );
  OAI211_X1 U9828 ( .C1(n8216), .C2(n9158), .A(n8214), .B(n8213), .ZN(P2_U3267) );
  OAI222_X1 U9829 ( .A1(P1_U3086), .A2(n8217), .B1(n9792), .B2(n8216), .C1(
        n8215), .C2(n8565), .ZN(P1_U3327) );
  INV_X1 U9830 ( .A(n8218), .ZN(n8568) );
  AOI22_X1 U9831 ( .A1(n8219), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9156), .ZN(n8220) );
  OAI21_X1 U9832 ( .B1(n8568), .B2(n9158), .A(n8220), .ZN(P2_U3266) );
  INV_X1 U9833 ( .A(n8442), .ZN(n9159) );
  OAI222_X1 U9834 ( .A1(n8565), .A2(n8222), .B1(n9792), .B2(n9159), .C1(
        P1_U3086), .C2(n5359), .ZN(P1_U3325) );
  XNOR2_X1 U9835 ( .A(n8223), .B(n8225), .ZN(n10070) );
  INV_X1 U9836 ( .A(n8224), .ZN(n8229) );
  AOI21_X1 U9837 ( .B1(n8227), .B2(n8226), .A(n8225), .ZN(n8228) );
  NOR3_X1 U9838 ( .A1(n8229), .A2(n8228), .A3(n9596), .ZN(n8233) );
  OR2_X1 U9839 ( .A1(n8230), .A2(n9253), .ZN(n8232) );
  NAND2_X1 U9840 ( .A1(n9311), .A2(n9287), .ZN(n8231) );
  NAND2_X1 U9841 ( .A1(n8232), .A2(n8231), .ZN(n9883) );
  NOR2_X1 U9842 ( .A1(n8233), .A2(n9883), .ZN(n10066) );
  INV_X1 U9843 ( .A(n10066), .ZN(n8240) );
  OAI211_X1 U9844 ( .C1(n8235), .C2(n10068), .A(n10058), .B(n8234), .ZN(n10065) );
  NAND2_X1 U9845 ( .A1(n10033), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n8236) );
  OAI21_X1 U9846 ( .B1(n10021), .B2(n9889), .A(n8236), .ZN(n8237) );
  AOI21_X1 U9847 ( .B1(n4595), .B2(n10035), .A(n8237), .ZN(n8238) );
  OAI21_X1 U9848 ( .B1(n10065), .B2(n10038), .A(n8238), .ZN(n8239) );
  AOI21_X1 U9849 ( .B1(n8240), .B2(n10023), .A(n8239), .ZN(n8241) );
  OAI21_X1 U9850 ( .B1(n10070), .B2(n10020), .A(n8241), .ZN(P1_U3282) );
  XNOR2_X1 U9851 ( .A(n8243), .B(n8242), .ZN(n8256) );
  NAND2_X1 U9852 ( .A1(n10222), .A2(n10196), .ZN(n9142) );
  INV_X1 U9853 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8246) );
  XNOR2_X1 U9854 ( .A(n8244), .B(n8493), .ZN(n8245) );
  AOI222_X1 U9855 ( .A1(n10135), .A2(n8245), .B1(n8699), .B2(n10132), .C1(
        n8518), .C2(n10130), .ZN(n8252) );
  MUX2_X1 U9856 ( .A(n8246), .B(n8252), .S(n10222), .Z(n8248) );
  NAND2_X1 U9857 ( .A1(n8694), .A2(n9144), .ZN(n8247) );
  OAI211_X1 U9858 ( .C1(n8256), .C2(n9142), .A(n8248), .B(n8247), .ZN(P2_U3435) );
  NAND2_X1 U9859 ( .A1(n10243), .A2(n10196), .ZN(n9049) );
  MUX2_X1 U9860 ( .A(n8249), .B(n8252), .S(n10243), .Z(n8251) );
  INV_X1 U9861 ( .A(n9037), .ZN(n9050) );
  NAND2_X1 U9862 ( .A1(n8694), .A2(n9050), .ZN(n8250) );
  OAI211_X1 U9863 ( .C1(n9049), .C2(n8256), .A(n8251), .B(n8250), .ZN(P2_U3474) );
  MUX2_X1 U9864 ( .A(n8728), .B(n8252), .S(n10160), .Z(n8255) );
  INV_X1 U9865 ( .A(n8686), .ZN(n8253) );
  AOI22_X1 U9866 ( .A1(n8694), .A2(n10138), .B1(n10140), .B2(n8253), .ZN(n8254) );
  OAI211_X1 U9867 ( .C1(n8256), .C2(n8988), .A(n8255), .B(n8254), .ZN(P2_U3218) );
  AOI22_X1 U9868 ( .A1(n9461), .A2(n9183), .B1(n4330), .B2(n9296), .ZN(n8257)
         );
  XOR2_X1 U9869 ( .A(n8258), .B(n8257), .Z(n8260) );
  OAI22_X1 U9870 ( .A1(n9741), .A2(n6545), .B1(n9197), .B2(n6601), .ZN(n8259)
         );
  NOR2_X1 U9871 ( .A1(n8260), .A2(n8259), .ZN(n9202) );
  AOI21_X1 U9872 ( .B1(n8260), .B2(n8259), .A(n9202), .ZN(n8264) );
  INV_X1 U9873 ( .A(n8261), .ZN(n8262) );
  NAND2_X1 U9874 ( .A1(n8263), .A2(n8262), .ZN(n8265) );
  AOI21_X1 U9875 ( .B1(n8266), .B2(n8265), .A(n8264), .ZN(n8267) );
  OAI21_X1 U9876 ( .B1(n9195), .B2(n8267), .A(n9885), .ZN(n8273) );
  OR2_X1 U9877 ( .A1(n9189), .A2(n9275), .ZN(n8269) );
  NAND2_X1 U9878 ( .A1(n9297), .A2(n9286), .ZN(n8268) );
  NAND2_X1 U9879 ( .A1(n8269), .A2(n8268), .ZN(n9455) );
  OAI22_X1 U9880 ( .A1(n9462), .A2(n9890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8270), .ZN(n8271) );
  AOI21_X1 U9881 ( .B1(n9455), .B2(n9882), .A(n8271), .ZN(n8272) );
  NAND2_X1 U9882 ( .A1(n9610), .A2(n9306), .ZN(n8280) );
  NAND2_X1 U9883 ( .A1(n9590), .A2(n8281), .ZN(n8282) );
  OAI21_X1 U9884 ( .B1(n9604), .B2(n9176), .A(n8282), .ZN(n9582) );
  INV_X1 U9885 ( .A(n9582), .ZN(n8284) );
  NAND2_X1 U9886 ( .A1(n8288), .A2(n4955), .ZN(n9518) );
  INV_X1 U9887 ( .A(n9276), .ZN(n9300) );
  INV_X1 U9888 ( .A(n9252), .ZN(n9298) );
  NOR2_X1 U9889 ( .A1(n9478), .A2(n9297), .ZN(n8294) );
  OAI22_X1 U9890 ( .A1(n9450), .A2(n9453), .B1(n9461), .B2(n9296), .ZN(n9438)
         );
  NAND2_X1 U9891 ( .A1(n9438), .A2(n9437), .ZN(n9436) );
  INV_X1 U9892 ( .A(n9189), .ZN(n9295) );
  NAND2_X1 U9893 ( .A1(n9436), .A2(n8295), .ZN(n8298) );
  INV_X1 U9894 ( .A(n8298), .ZN(n8296) );
  NAND2_X1 U9895 ( .A1(n8296), .A2(n8316), .ZN(n8300) );
  NAND2_X1 U9896 ( .A1(n8298), .A2(n8297), .ZN(n8299) );
  NAND2_X1 U9897 ( .A1(n8300), .A2(n8299), .ZN(n9654) );
  AOI21_X1 U9898 ( .B1(n9650), .B2(n9439), .A(n9428), .ZN(n9651) );
  INV_X1 U9899 ( .A(n9650), .ZN(n8305) );
  INV_X1 U9900 ( .A(n8301), .ZN(n8302) );
  NAND3_X1 U9901 ( .A1(n8302), .A2(P1_REG3_REG_28__SCAN_IN), .A3(n10032), .ZN(
        n8304) );
  NAND2_X1 U9902 ( .A1(n10033), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8303) );
  OAI211_X1 U9903 ( .C1(n8305), .C2(n9629), .A(n8304), .B(n8303), .ZN(n8320)
         );
  NAND2_X1 U9904 ( .A1(n9452), .A2(n9453), .ZN(n9451) );
  INV_X1 U9905 ( .A(n9437), .ZN(n9443) );
  AOI22_X1 U9906 ( .A1(n9295), .A2(n9286), .B1(n8317), .B2(n9294), .ZN(n8318)
         );
  NOR2_X1 U9907 ( .A1(n4345), .A2(n10033), .ZN(n8319) );
  AOI211_X1 U9908 ( .C1(n9651), .C2(n9547), .A(n8320), .B(n8319), .ZN(n8321)
         );
  NAND2_X1 U9909 ( .A1(n8869), .A2(n8322), .ZN(n8324) );
  MUX2_X1 U9910 ( .A(n8324), .B(n8323), .S(n8458), .Z(n8325) );
  NOR2_X1 U9911 ( .A1(n8325), .A2(n8425), .ZN(n8424) );
  AND2_X1 U9912 ( .A1(n8327), .A2(n8326), .ZN(n8328) );
  OAI21_X1 U9913 ( .B1(n8329), .B2(n8328), .A(n8457), .ZN(n8337) );
  OAI21_X1 U9914 ( .B1(n8337), .B2(n8331), .A(n8333), .ZN(n8332) );
  MUX2_X1 U9915 ( .A(n8333), .B(n8332), .S(n8457), .Z(n8344) );
  NOR2_X1 U9916 ( .A1(n7345), .A2(n8334), .ZN(n8336) );
  AOI21_X1 U9917 ( .B1(n8337), .B2(n8336), .A(n8335), .ZN(n8343) );
  NAND2_X1 U9918 ( .A1(n8338), .A2(n8346), .ZN(n8341) );
  NAND2_X1 U9919 ( .A1(n8360), .A2(n8339), .ZN(n8340) );
  MUX2_X1 U9920 ( .A(n8341), .B(n8340), .S(n8458), .Z(n8342) );
  AOI21_X1 U9921 ( .B1(n8344), .B2(n8343), .A(n8342), .ZN(n8345) );
  OR2_X1 U9922 ( .A1(n8345), .A2(n8477), .ZN(n8364) );
  OAI21_X1 U9923 ( .B1(n8364), .B2(n4643), .A(n8347), .ZN(n8348) );
  NAND3_X1 U9924 ( .A1(n8348), .A2(n8362), .A3(n8368), .ZN(n8349) );
  INV_X1 U9925 ( .A(n8483), .ZN(n8369) );
  NAND3_X1 U9926 ( .A1(n8349), .A2(n8369), .A3(n8365), .ZN(n8351) );
  NAND3_X1 U9927 ( .A1(n8351), .A2(n8353), .A3(n8350), .ZN(n8359) );
  NAND2_X1 U9928 ( .A1(n8373), .A2(n8352), .ZN(n8355) );
  NAND2_X1 U9929 ( .A1(n8357), .A2(n8353), .ZN(n8354) );
  MUX2_X1 U9930 ( .A(n8355), .B(n8354), .S(n8457), .Z(n8356) );
  INV_X1 U9931 ( .A(n8356), .ZN(n8375) );
  NAND2_X1 U9932 ( .A1(n8377), .A2(n8357), .ZN(n8358) );
  INV_X1 U9933 ( .A(n8360), .ZN(n8363) );
  OAI211_X1 U9934 ( .C1(n8364), .C2(n8363), .A(n8362), .B(n8361), .ZN(n8367)
         );
  NAND3_X1 U9935 ( .A1(n8367), .A2(n8366), .A3(n8365), .ZN(n8370) );
  NAND3_X1 U9936 ( .A1(n8370), .A2(n8369), .A3(n8368), .ZN(n8372) );
  NAND2_X1 U9937 ( .A1(n8372), .A2(n8371), .ZN(n8376) );
  NAND2_X1 U9938 ( .A1(n8378), .A2(n8373), .ZN(n8374) );
  NAND2_X1 U9939 ( .A1(n8382), .A2(n8377), .ZN(n8380) );
  NAND2_X1 U9940 ( .A1(n8381), .A2(n8378), .ZN(n8379) );
  MUX2_X1 U9941 ( .A(n8380), .B(n8379), .S(n8458), .Z(n8385) );
  MUX2_X1 U9942 ( .A(n8382), .B(n8381), .S(n8457), .Z(n8383) );
  NAND2_X1 U9943 ( .A1(n10220), .A2(n8386), .ZN(n8387) );
  MUX2_X1 U9944 ( .A(n8388), .B(n8387), .S(n8457), .Z(n8389) );
  INV_X1 U9945 ( .A(n8391), .ZN(n8393) );
  MUX2_X1 U9946 ( .A(n8393), .B(n4655), .S(n8457), .Z(n8394) );
  NOR2_X1 U9947 ( .A1(n8986), .A2(n8394), .ZN(n8395) );
  NAND2_X1 U9948 ( .A1(n8396), .A2(n8395), .ZN(n8400) );
  MUX2_X1 U9949 ( .A(n8398), .B(n8397), .S(n8458), .Z(n8399) );
  INV_X1 U9950 ( .A(n8406), .ZN(n8408) );
  NAND2_X1 U9951 ( .A1(n8411), .A2(n8410), .ZN(n8413) );
  OAI21_X1 U9952 ( .B1(n8414), .B2(n8413), .A(n8412), .ZN(n8416) );
  MUX2_X1 U9953 ( .A(n8418), .B(n8417), .S(n8458), .Z(n8419) );
  MUX2_X1 U9954 ( .A(n8421), .B(n8420), .S(n8457), .Z(n8422) );
  INV_X1 U9955 ( .A(n8425), .ZN(n8476) );
  AND2_X1 U9956 ( .A1(n8427), .A2(n8476), .ZN(n8426) );
  INV_X1 U9957 ( .A(n8427), .ZN(n8475) );
  NAND2_X1 U9958 ( .A1(n8430), .A2(n8429), .ZN(n8859) );
  AND2_X1 U9959 ( .A1(n8434), .A2(n8435), .ZN(n8842) );
  MUX2_X1 U9960 ( .A(n8432), .B(n8431), .S(n8458), .Z(n8433) );
  MUX2_X1 U9961 ( .A(n8435), .B(n8434), .S(n8458), .Z(n8436) );
  MUX2_X1 U9962 ( .A(n8438), .B(n8437), .S(n8457), .Z(n8439) );
  MUX2_X1 U9963 ( .A(n8697), .B(n9064), .S(n8457), .Z(n8448) );
  NAND2_X1 U9964 ( .A1(n8442), .A2(n8451), .ZN(n8444) );
  NAND2_X1 U9965 ( .A1(n8450), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8443) );
  INV_X1 U9966 ( .A(n8696), .ZN(n8445) );
  NAND2_X1 U9967 ( .A1(n9059), .A2(n8445), .ZN(n8502) );
  NAND2_X1 U9968 ( .A1(n8996), .A2(n8696), .ZN(n8501) );
  INV_X1 U9969 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8456) );
  AOI22_X1 U9970 ( .A1(n8453), .A2(P2_REG0_REG_31__SCAN_IN), .B1(n8452), .B2(
        P2_REG1_REG_31__SCAN_IN), .ZN(n8454) );
  OAI211_X1 U9971 ( .C1(n6149), .C2(n8456), .A(n8455), .B(n8454), .ZN(n8806)
         );
  NAND2_X1 U9972 ( .A1(n8502), .A2(n8458), .ZN(n8460) );
  INV_X1 U9973 ( .A(n8806), .ZN(n8468) );
  INV_X1 U9974 ( .A(n8464), .ZN(n8465) );
  NAND3_X1 U9975 ( .A1(n8470), .A2(n8996), .A3(n8468), .ZN(n8473) );
  INV_X1 U9976 ( .A(n8501), .ZN(n8469) );
  OAI21_X1 U9977 ( .B1(n8470), .B2(n8469), .A(n9055), .ZN(n8472) );
  AOI21_X1 U9978 ( .B1(n8473), .B2(n8472), .A(n8471), .ZN(n8508) );
  INV_X1 U9979 ( .A(n8822), .ZN(n8499) );
  NOR2_X1 U9980 ( .A1(n8475), .A2(n8474), .ZN(n8870) );
  NAND2_X1 U9981 ( .A1(n8476), .A2(n8869), .ZN(n8875) );
  INV_X1 U9982 ( .A(n8914), .ZN(n8911) );
  NOR4_X1 U9983 ( .A1(n7345), .A2(n8478), .A3(n8477), .A4(n8335), .ZN(n8480)
         );
  NAND3_X1 U9984 ( .A1(n8480), .A2(n10137), .A3(n8479), .ZN(n8484) );
  NOR4_X1 U9985 ( .A1(n8484), .A2(n8483), .A3(n8482), .A4(n8481), .ZN(n8488)
         );
  NAND4_X1 U9986 ( .A1(n8488), .A2(n8487), .A3(n8486), .A4(n8485), .ZN(n8491)
         );
  NOR4_X1 U9987 ( .A1(n8986), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n8492)
         );
  NAND4_X1 U9988 ( .A1(n8954), .A2(n8493), .A3(n8968), .A4(n8492), .ZN(n8494)
         );
  OR4_X1 U9989 ( .A1(n8911), .A2(n8944), .A3(n8927), .A4(n8494), .ZN(n8495) );
  NOR4_X1 U9990 ( .A1(n8875), .A2(n8496), .A3(n8901), .A4(n8495), .ZN(n8497)
         );
  NAND4_X1 U9991 ( .A1(n8842), .A2(n8870), .A3(n8497), .A4(n8859), .ZN(n8498)
         );
  NOR4_X1 U9992 ( .A1(n8500), .A2(n8499), .A3(n8834), .A4(n8498), .ZN(n8503)
         );
  NAND4_X1 U9993 ( .A1(n4964), .A2(n8503), .A3(n8502), .A4(n8501), .ZN(n8506)
         );
  INV_X1 U9994 ( .A(n8504), .ZN(n8505) );
  NOR3_X1 U9995 ( .A1(n8512), .A2(n8511), .A3(n8510), .ZN(n8515) );
  OAI21_X1 U9996 ( .B1(n8516), .B2(n8513), .A(P2_B_REG_SCAN_IN), .ZN(n8514) );
  OAI22_X1 U9997 ( .A1(n8517), .A2(n8516), .B1(n8515), .B2(n8514), .ZN(
        P2_U3296) );
  XNOR2_X1 U9998 ( .A(n8694), .B(n4342), .ZN(n8522) );
  XOR2_X1 U9999 ( .A(n8978), .B(n8522), .Z(n8690) );
  INV_X1 U10000 ( .A(n8522), .ZN(n8523) );
  NOR2_X2 U10001 ( .A1(n8687), .A2(n4949), .ZN(n8613) );
  XNOR2_X1 U10002 ( .A(n9130), .B(n4342), .ZN(n8614) );
  NAND2_X1 U10003 ( .A1(n8613), .A2(n8614), .ZN(n8526) );
  INV_X1 U10004 ( .A(n8613), .ZN(n8525) );
  INV_X1 U10005 ( .A(n8614), .ZN(n8524) );
  XNOR2_X1 U10006 ( .A(n9039), .B(n8558), .ZN(n8527) );
  NOR2_X1 U10007 ( .A1(n8527), .A2(n8969), .ZN(n8660) );
  AOI21_X1 U10008 ( .B1(n8527), .B2(n8969), .A(n8660), .ZN(n8624) );
  XNOR2_X1 U10009 ( .A(n8657), .B(n4342), .ZN(n8531) );
  XNOR2_X1 U10010 ( .A(n8531), .B(n8926), .ZN(n8659) );
  AND2_X1 U10011 ( .A1(n8624), .A2(n8659), .ZN(n8528) );
  NAND2_X1 U10012 ( .A1(n8622), .A2(n8528), .ZN(n8663) );
  INV_X1 U10013 ( .A(n8659), .ZN(n8530) );
  INV_X1 U10014 ( .A(n8660), .ZN(n8529) );
  NAND2_X1 U10015 ( .A1(n8531), .A2(n8959), .ZN(n8532) );
  XNOR2_X1 U10016 ( .A(n9115), .B(n4342), .ZN(n8584) );
  INV_X1 U10017 ( .A(n8584), .ZN(n8534) );
  XNOR2_X1 U10018 ( .A(n9109), .B(n8558), .ZN(n8536) );
  AOI21_X1 U10019 ( .B1(n8536), .B2(n8933), .A(n8595), .ZN(n8642) );
  XNOR2_X1 U10020 ( .A(n9103), .B(n4342), .ZN(n8538) );
  XNOR2_X1 U10021 ( .A(n8538), .B(n8917), .ZN(n8594) );
  NAND2_X1 U10022 ( .A1(n8537), .A2(n8594), .ZN(n8597) );
  INV_X1 U10023 ( .A(n8538), .ZN(n8539) );
  NAND2_X1 U10024 ( .A1(n8650), .A2(n8905), .ZN(n8541) );
  NOR2_X1 U10025 ( .A1(n8650), .A2(n8905), .ZN(n8540) );
  XNOR2_X1 U10026 ( .A(n9096), .B(n4342), .ZN(n8543) );
  INV_X1 U10027 ( .A(n8542), .ZN(n8544) );
  NAND2_X1 U10028 ( .A1(n8544), .A2(n8543), .ZN(n8633) );
  XNOR2_X1 U10029 ( .A(n9090), .B(n4342), .ZN(n8546) );
  NAND2_X1 U10030 ( .A1(n8546), .A2(n8854), .ZN(n8545) );
  INV_X1 U10031 ( .A(n8545), .ZN(n8547) );
  XNOR2_X1 U10032 ( .A(n8546), .B(n8877), .ZN(n8635) );
  XOR2_X1 U10033 ( .A(n4342), .B(n9083), .Z(n8550) );
  INV_X1 U10034 ( .A(n8550), .ZN(n8549) );
  NOR2_X1 U10035 ( .A1(n8550), .A2(n8844), .ZN(n8551) );
  XNOR2_X1 U10036 ( .A(n9076), .B(n8552), .ZN(n8553) );
  XNOR2_X1 U10037 ( .A(n8555), .B(n8553), .ZN(n8671) );
  NAND2_X1 U10038 ( .A1(n8671), .A2(n8855), .ZN(n8557) );
  INV_X1 U10039 ( .A(n8553), .ZN(n8554) );
  OR2_X1 U10040 ( .A1(n8555), .A2(n8554), .ZN(n8556) );
  NAND2_X1 U10041 ( .A1(n8557), .A2(n8556), .ZN(n8569) );
  XNOR2_X1 U10042 ( .A(n9070), .B(n8558), .ZN(n8559) );
  NAND2_X1 U10043 ( .A1(n8559), .A2(n8845), .ZN(n8560) );
  OAI21_X1 U10044 ( .B1(n8559), .B2(n8845), .A(n8560), .ZN(n8570) );
  AOI22_X1 U10045 ( .A1(n8845), .A2(n8672), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8562) );
  NAND2_X1 U10046 ( .A1(n8827), .A2(n8673), .ZN(n8561) );
  OAI211_X1 U10047 ( .C1(n8825), .C2(n8676), .A(n8562), .B(n8561), .ZN(n8563)
         );
  AOI21_X1 U10048 ( .B1(n9064), .B2(n8693), .A(n8563), .ZN(n8564) );
  OAI222_X1 U10049 ( .A1(n9792), .A2(n8568), .B1(n8567), .B2(P1_U3086), .C1(
        n8566), .C2(n8565), .ZN(P1_U3326) );
  INV_X1 U10050 ( .A(n9070), .ZN(n9002) );
  AOI21_X1 U10051 ( .B1(n8569), .B2(n8570), .A(n8688), .ZN(n8572) );
  NAND2_X1 U10052 ( .A1(n8572), .A2(n8571), .ZN(n8576) );
  AOI22_X1 U10053 ( .A1(n8698), .A2(n8672), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8573) );
  OAI21_X1 U10054 ( .B1(n8837), .B2(n8676), .A(n8573), .ZN(n8574) );
  AOI21_X1 U10055 ( .B1(n8838), .B2(n8673), .A(n8574), .ZN(n8575) );
  OAI211_X1 U10056 ( .C1(n9002), .C2(n8670), .A(n8576), .B(n8575), .ZN(
        P2_U3154) );
  XNOR2_X1 U10057 ( .A(n8577), .B(n8888), .ZN(n8582) );
  AOI22_X1 U10058 ( .A1(n8672), .A2(n8905), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8579) );
  NAND2_X1 U10059 ( .A1(n8673), .A2(n8879), .ZN(n8578) );
  OAI211_X1 U10060 ( .C1(n8854), .C2(n8676), .A(n8579), .B(n8578), .ZN(n8580)
         );
  AOI21_X1 U10061 ( .B1(n9096), .B2(n8693), .A(n8580), .ZN(n8581) );
  OAI21_X1 U10062 ( .B1(n8582), .B2(n8688), .A(n8581), .ZN(P2_U3156) );
  INV_X1 U10063 ( .A(n8583), .ZN(n8586) );
  XNOR2_X1 U10064 ( .A(n8584), .B(n8918), .ZN(n8585) );
  XNOR2_X1 U10065 ( .A(n8586), .B(n8585), .ZN(n8592) );
  NAND2_X1 U10066 ( .A1(n8672), .A2(n8926), .ZN(n8588) );
  OAI211_X1 U10067 ( .C1(n8601), .C2(n8676), .A(n8588), .B(n8587), .ZN(n8589)
         );
  AOI21_X1 U10068 ( .B1(n8934), .B2(n8673), .A(n8589), .ZN(n8591) );
  NAND2_X1 U10069 ( .A1(n9115), .A2(n8693), .ZN(n8590) );
  OAI211_X1 U10070 ( .C1(n8592), .C2(n8688), .A(n8591), .B(n8590), .ZN(
        P2_U3159) );
  INV_X1 U10071 ( .A(n9103), .ZN(n8605) );
  INV_X1 U10072 ( .A(n8593), .ZN(n8596) );
  NOR3_X1 U10073 ( .A1(n8596), .A2(n8595), .A3(n8594), .ZN(n8599) );
  INV_X1 U10074 ( .A(n8597), .ZN(n8598) );
  OAI21_X1 U10075 ( .B1(n8599), .B2(n8598), .A(n8664), .ZN(n8604) );
  AOI22_X1 U10076 ( .A1(n8683), .A2(n8905), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8600) );
  OAI21_X1 U10077 ( .B1(n8601), .B2(n8681), .A(n8600), .ZN(n8602) );
  AOI21_X1 U10078 ( .B1(n8908), .B2(n8673), .A(n8602), .ZN(n8603) );
  OAI211_X1 U10079 ( .C1(n8605), .C2(n8670), .A(n8604), .B(n8603), .ZN(
        P2_U3163) );
  XOR2_X1 U10080 ( .A(n8607), .B(n8606), .Z(n8612) );
  AOI22_X1 U10081 ( .A1(n8698), .A2(n8683), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8609) );
  NAND2_X1 U10082 ( .A1(n8673), .A2(n8857), .ZN(n8608) );
  OAI211_X1 U10083 ( .C1(n8854), .C2(n8681), .A(n8609), .B(n8608), .ZN(n8610)
         );
  AOI21_X1 U10084 ( .B1(n9083), .B2(n8693), .A(n8610), .ZN(n8611) );
  OAI21_X1 U10085 ( .B1(n8612), .B2(n8688), .A(n8611), .ZN(P2_U3165) );
  XNOR2_X1 U10086 ( .A(n8614), .B(n8960), .ZN(n8615) );
  XNOR2_X1 U10087 ( .A(n8613), .B(n8615), .ZN(n8621) );
  NAND2_X1 U10088 ( .A1(P2_U3151), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8754) );
  OAI21_X1 U10089 ( .B1(n8681), .B2(n8616), .A(n8754), .ZN(n8617) );
  AOI21_X1 U10090 ( .B1(n8683), .B2(n8969), .A(n8617), .ZN(n8618) );
  OAI21_X1 U10091 ( .B1(n8972), .B2(n8685), .A(n8618), .ZN(n8619) );
  AOI21_X1 U10092 ( .B1(n9130), .B2(n8693), .A(n8619), .ZN(n8620) );
  OAI21_X1 U10093 ( .B1(n8621), .B2(n8688), .A(n8620), .ZN(P2_U3166) );
  INV_X1 U10094 ( .A(n9039), .ZN(n8631) );
  NAND2_X1 U10095 ( .A1(n8623), .A2(n8624), .ZN(n8658) );
  OAI21_X1 U10096 ( .B1(n8624), .B2(n8623), .A(n8658), .ZN(n8625) );
  NAND2_X1 U10097 ( .A1(n8625), .A2(n8664), .ZN(n8630) );
  INV_X1 U10098 ( .A(n8961), .ZN(n8628) );
  AND2_X1 U10099 ( .A1(P2_U3151), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8767) );
  AOI21_X1 U10100 ( .B1(n8683), .B2(n8926), .A(n8767), .ZN(n8626) );
  OAI21_X1 U10101 ( .B1(n8960), .B2(n8681), .A(n8626), .ZN(n8627) );
  AOI21_X1 U10102 ( .B1(n8628), .B2(n8673), .A(n8627), .ZN(n8629) );
  OAI211_X1 U10103 ( .C1(n8631), .C2(n8670), .A(n8630), .B(n8629), .ZN(
        P2_U3168) );
  NAND2_X1 U10104 ( .A1(n8632), .A2(n8633), .ZN(n8634) );
  XOR2_X1 U10105 ( .A(n8635), .B(n8634), .Z(n8640) );
  AOI22_X1 U10106 ( .A1(n8844), .A2(n8683), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8637) );
  NAND2_X1 U10107 ( .A1(n8673), .A2(n8867), .ZN(n8636) );
  OAI211_X1 U10108 ( .C1(n8865), .C2(n8681), .A(n8637), .B(n8636), .ZN(n8638)
         );
  AOI21_X1 U10109 ( .B1(n9090), .B2(n8693), .A(n8638), .ZN(n8639) );
  OAI21_X1 U10110 ( .B1(n8640), .B2(n8688), .A(n8639), .ZN(P2_U3169) );
  INV_X1 U10111 ( .A(n9109), .ZN(n8648) );
  OAI21_X1 U10112 ( .B1(n8642), .B2(n8641), .A(n8593), .ZN(n8643) );
  NAND2_X1 U10113 ( .A1(n8643), .A2(n8664), .ZN(n8647) );
  AOI22_X1 U10114 ( .A1(n8683), .A2(n8917), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8644) );
  OAI21_X1 U10115 ( .B1(n8943), .B2(n8681), .A(n8644), .ZN(n8645) );
  AOI21_X1 U10116 ( .B1(n8921), .B2(n8673), .A(n8645), .ZN(n8646) );
  OAI211_X1 U10117 ( .C1(n8648), .C2(n8670), .A(n8647), .B(n8646), .ZN(
        P2_U3173) );
  XNOR2_X1 U10118 ( .A(n8650), .B(n8905), .ZN(n8651) );
  XNOR2_X1 U10119 ( .A(n8649), .B(n8651), .ZN(n8656) );
  AOI22_X1 U10120 ( .A1(n8672), .A2(n8917), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8653) );
  NAND2_X1 U10121 ( .A1(n8673), .A2(n8890), .ZN(n8652) );
  OAI211_X1 U10122 ( .C1(n8865), .C2(n8676), .A(n8653), .B(n8652), .ZN(n8654)
         );
  AOI21_X1 U10123 ( .B1(n9019), .B2(n8693), .A(n8654), .ZN(n8655) );
  OAI21_X1 U10124 ( .B1(n8656), .B2(n8688), .A(n8655), .ZN(P2_U3175) );
  INV_X1 U10125 ( .A(n8657), .ZN(n9123) );
  INV_X1 U10126 ( .A(n8658), .ZN(n8661) );
  NOR3_X1 U10127 ( .A1(n8661), .A2(n8660), .A3(n8659), .ZN(n8665) );
  OAI21_X1 U10128 ( .B1(n8665), .B2(n4414), .A(n8664), .ZN(n8669) );
  NAND2_X1 U10129 ( .A1(n8672), .A2(n8969), .ZN(n8666) );
  NAND2_X1 U10130 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8790) );
  OAI211_X1 U10131 ( .C1(n8943), .C2(n8676), .A(n8666), .B(n8790), .ZN(n8667)
         );
  AOI21_X1 U10132 ( .B1(n8947), .B2(n8673), .A(n8667), .ZN(n8668) );
  OAI211_X1 U10133 ( .C1(n9123), .C2(n8670), .A(n8669), .B(n8668), .ZN(
        P2_U3178) );
  XNOR2_X1 U10134 ( .A(n4335), .B(n8698), .ZN(n8679) );
  AOI22_X1 U10135 ( .A1(n8844), .A2(n8672), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8675) );
  NAND2_X1 U10136 ( .A1(n8847), .A2(n8673), .ZN(n8674) );
  OAI211_X1 U10137 ( .C1(n8826), .C2(n8676), .A(n8675), .B(n8674), .ZN(n8677)
         );
  AOI21_X1 U10138 ( .B1(n9076), .B2(n8693), .A(n8677), .ZN(n8678) );
  OAI21_X1 U10139 ( .B1(n8679), .B2(n8688), .A(n8678), .ZN(P2_U3180) );
  NAND2_X1 U10140 ( .A1(P2_U3151), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n8736) );
  OAI21_X1 U10141 ( .B1(n8681), .B2(n8680), .A(n8736), .ZN(n8682) );
  AOI21_X1 U10142 ( .B1(n8683), .B2(n8699), .A(n8682), .ZN(n8684) );
  OAI21_X1 U10143 ( .B1(n8686), .B2(n8685), .A(n8684), .ZN(n8692) );
  AOI211_X1 U10144 ( .C1(n8690), .C2(n8689), .A(n8688), .B(n8687), .ZN(n8691)
         );
  AOI211_X1 U10145 ( .C1(n8694), .C2(n8693), .A(n8692), .B(n8691), .ZN(n8695)
         );
  INV_X1 U10146 ( .A(n8695), .ZN(P2_U3181) );
  MUX2_X1 U10147 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8806), .S(P2_U3893), .Z(
        P2_U3522) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8696), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10149 ( .A(n8697), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8705), .Z(
        P2_U3519) );
  MUX2_X1 U10150 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8845), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10151 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8698), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U10152 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8844), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10153 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8877), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10154 ( .A(n8888), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8705), .Z(
        P2_U3514) );
  MUX2_X1 U10155 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8905), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10156 ( .A(n8917), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8705), .Z(
        P2_U3512) );
  MUX2_X1 U10157 ( .A(n8933), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8705), .Z(
        P2_U3511) );
  MUX2_X1 U10158 ( .A(n8918), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8705), .Z(
        P2_U3510) );
  MUX2_X1 U10159 ( .A(n8926), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8705), .Z(
        P2_U3509) );
  MUX2_X1 U10160 ( .A(n8969), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8705), .Z(
        P2_U3508) );
  MUX2_X1 U10161 ( .A(n8699), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8705), .Z(
        P2_U3507) );
  MUX2_X1 U10162 ( .A(n8978), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8705), .Z(
        P2_U3506) );
  MUX2_X1 U10163 ( .A(n8977), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8705), .Z(
        P2_U3504) );
  MUX2_X1 U10164 ( .A(n8700), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8705), .Z(
        P2_U3503) );
  MUX2_X1 U10165 ( .A(n8701), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8705), .Z(
        P2_U3502) );
  MUX2_X1 U10166 ( .A(n8068), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8705), .Z(
        P2_U3501) );
  MUX2_X1 U10167 ( .A(n8702), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8705), .Z(
        P2_U3500) );
  MUX2_X1 U10168 ( .A(n8703), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8705), .Z(
        P2_U3499) );
  MUX2_X1 U10169 ( .A(n8704), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8705), .Z(
        P2_U3498) );
  MUX2_X1 U10170 ( .A(n8706), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8705), .Z(
        P2_U3497) );
  MUX2_X1 U10171 ( .A(n8707), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8705), .Z(
        P2_U3496) );
  MUX2_X1 U10172 ( .A(n10133), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8705), .Z(
        P2_U3495) );
  MUX2_X1 U10173 ( .A(n10131), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8705), .Z(
        P2_U3493) );
  MUX2_X1 U10174 ( .A(n6107), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8705), .Z(
        P2_U3492) );
  MUX2_X1 U10175 ( .A(n8708), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8705), .Z(
        P2_U3491) );
  AOI21_X1 U10176 ( .B1(n8711), .B2(n8710), .A(n8709), .ZN(n8712) );
  OR2_X1 U10177 ( .A1(n8712), .A2(n10122), .ZN(n8725) );
  AOI21_X1 U10178 ( .B1(n10090), .B2(n8714), .A(n8713), .ZN(n8724) );
  NAND2_X1 U10179 ( .A1(n8715), .A2(n10240), .ZN(n8716) );
  NAND2_X1 U10180 ( .A1(n8716), .A2(n4838), .ZN(n8721) );
  OAI21_X1 U10181 ( .B1(n8719), .B2(n8718), .A(n8717), .ZN(n8720) );
  AOI22_X1 U10182 ( .A1(n8777), .A2(n8721), .B1(n5610), .B2(n8720), .ZN(n8723)
         );
  NAND2_X1 U10183 ( .A1(n10109), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n8722) );
  NAND4_X1 U10184 ( .A1(n8725), .A2(n8724), .A3(n8723), .A4(n8722), .ZN(
        P2_U3193) );
  AOI21_X1 U10185 ( .B1(n8728), .B2(n8727), .A(n8726), .ZN(n8743) );
  INV_X1 U10186 ( .A(n8729), .ZN(n8730) );
  NOR2_X1 U10187 ( .A1(n8730), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8732) );
  OAI21_X1 U10188 ( .B1(n8732), .B2(n8731), .A(n8777), .ZN(n8742) );
  OAI21_X1 U10189 ( .B1(n8735), .B2(n8734), .A(n8733), .ZN(n8740) );
  OAI21_X1 U10190 ( .B1(n10128), .B2(n8737), .A(n8736), .ZN(n8739) );
  INV_X1 U10191 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n9832) );
  NOR2_X1 U10192 ( .A1(n8803), .A2(n9832), .ZN(n8738) );
  AOI211_X1 U10193 ( .C1(n5610), .C2(n8740), .A(n8739), .B(n8738), .ZN(n8741)
         );
  OAI211_X1 U10194 ( .C1(n8743), .C2(n10122), .A(n8742), .B(n8741), .ZN(
        P2_U3197) );
  AOI21_X1 U10195 ( .B1(n4401), .B2(n8745), .A(n8744), .ZN(n8761) );
  AND2_X1 U10196 ( .A1(n8747), .A2(n8746), .ZN(n8750) );
  INV_X1 U10197 ( .A(n8748), .ZN(n8749) );
  OAI21_X1 U10198 ( .B1(n8750), .B2(n8749), .A(n8777), .ZN(n8760) );
  OAI21_X1 U10199 ( .B1(n8753), .B2(n8752), .A(n8751), .ZN(n8758) );
  OAI21_X1 U10200 ( .B1(n10128), .B2(n8755), .A(n8754), .ZN(n8757) );
  INV_X1 U10201 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n9835) );
  NOR2_X1 U10202 ( .A1(n8803), .A2(n9835), .ZN(n8756) );
  AOI211_X1 U10203 ( .C1(n5610), .C2(n8758), .A(n8757), .B(n8756), .ZN(n8759)
         );
  OAI211_X1 U10204 ( .C1(n8761), .C2(n10122), .A(n8760), .B(n8759), .ZN(
        P2_U3198) );
  INV_X1 U10205 ( .A(n8762), .ZN(n8763) );
  NOR2_X1 U10206 ( .A1(n8763), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8766) );
  OAI21_X1 U10207 ( .B1(n8766), .B2(n8765), .A(n8764), .ZN(n8781) );
  AOI21_X1 U10208 ( .B1(n10090), .B2(n8768), .A(n8767), .ZN(n8780) );
  AND2_X1 U10209 ( .A1(n8769), .A2(n9040), .ZN(n8770) );
  OAI21_X1 U10210 ( .B1(n8774), .B2(n8773), .A(n8772), .ZN(n8775) );
  NAND2_X1 U10211 ( .A1(n10109), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n8778) );
  NAND4_X1 U10212 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), .ZN(
        P2_U3199) );
  INV_X1 U10213 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n8804) );
  INV_X1 U10214 ( .A(n8782), .ZN(n8785) );
  INV_X1 U10215 ( .A(n8783), .ZN(n8784) );
  NAND2_X1 U10216 ( .A1(n8785), .A2(n8784), .ZN(n8786) );
  AOI21_X1 U10217 ( .B1(n8787), .B2(n8786), .A(n10122), .ZN(n8793) );
  AOI21_X1 U10218 ( .B1(n4366), .B2(n8789), .A(n8788), .ZN(n8791) );
  OAI21_X1 U10219 ( .B1(n10118), .B2(n8791), .A(n8790), .ZN(n8792) );
  NOR2_X1 U10220 ( .A1(n8793), .A2(n8792), .ZN(n8802) );
  NOR2_X1 U10221 ( .A1(n8795), .A2(n8794), .ZN(n8797) );
  INV_X1 U10222 ( .A(n8797), .ZN(n8796) );
  NAND2_X1 U10223 ( .A1(n5610), .A2(n8796), .ZN(n8800) );
  AOI21_X1 U10224 ( .B1(P2_U3893), .B2(n8797), .A(n10090), .ZN(n8799) );
  MUX2_X1 U10225 ( .A(n8800), .B(n8799), .S(n8798), .Z(n8801) );
  OAI211_X1 U10226 ( .C1(n8804), .C2(n8803), .A(n8802), .B(n8801), .ZN(
        P2_U3200) );
  AND2_X1 U10227 ( .A1(n8806), .A2(n8805), .ZN(n9056) );
  NOR2_X1 U10228 ( .A1(n8807), .A2(n10149), .ZN(n8816) );
  AOI21_X1 U10229 ( .B1(n9056), .B2(n10160), .A(n8816), .ZN(n8811) );
  NAND2_X1 U10230 ( .A1(n10162), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8808) );
  OAI211_X1 U10231 ( .C1(n8809), .C2(n8949), .A(n8811), .B(n8808), .ZN(
        P2_U3202) );
  NAND2_X1 U10232 ( .A1(n10162), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8810) );
  OAI211_X1 U10233 ( .C1(n8996), .C2(n8949), .A(n8811), .B(n8810), .ZN(
        P2_U3203) );
  INV_X1 U10234 ( .A(n8812), .ZN(n8820) );
  NAND2_X1 U10235 ( .A1(n8813), .A2(n10160), .ZN(n8818) );
  NOR2_X1 U10236 ( .A1(n8814), .A2(n8949), .ZN(n8815) );
  AOI211_X1 U10237 ( .C1(n10162), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8816), .B(
        n8815), .ZN(n8817) );
  OAI211_X1 U10238 ( .C1(n8820), .C2(n8819), .A(n8818), .B(n8817), .ZN(
        P2_U3204) );
  XNOR2_X1 U10239 ( .A(n8823), .B(n8822), .ZN(n8824) );
  OAI222_X1 U10240 ( .A1(n10155), .A2(n8826), .B1(n10157), .B2(n8825), .C1(
        n8824), .C2(n10153), .ZN(n8997) );
  INV_X1 U10241 ( .A(n8997), .ZN(n9062) );
  MUX2_X1 U10242 ( .A(n4543), .B(n9062), .S(n10160), .Z(n8829) );
  AOI22_X1 U10243 ( .A1(n9064), .A2(n10138), .B1(n10140), .B2(n8827), .ZN(
        n8828) );
  OAI211_X1 U10244 ( .C1(n9067), .C2(n8988), .A(n8829), .B(n8828), .ZN(
        P2_U3205) );
  NAND2_X1 U10245 ( .A1(n8833), .A2(n8832), .ZN(n8835) );
  XNOR2_X1 U10246 ( .A(n8835), .B(n8834), .ZN(n8836) );
  OAI222_X1 U10247 ( .A1(n10155), .A2(n8855), .B1(n10157), .B2(n8837), .C1(
        n8836), .C2(n10153), .ZN(n9001) );
  INV_X1 U10248 ( .A(n9001), .ZN(n9068) );
  MUX2_X1 U10249 ( .A(n4541), .B(n9068), .S(n10160), .Z(n8840) );
  AOI22_X1 U10250 ( .A1(n9070), .A2(n10138), .B1(n10140), .B2(n8838), .ZN(
        n8839) );
  OAI211_X1 U10251 ( .C1(n9073), .C2(n8988), .A(n8840), .B(n8839), .ZN(
        P2_U3206) );
  XOR2_X1 U10252 ( .A(n8842), .B(n8841), .Z(n9079) );
  XNOR2_X1 U10253 ( .A(n8843), .B(n8842), .ZN(n8846) );
  AOI222_X1 U10254 ( .A1(n10135), .A2(n8846), .B1(n8845), .B2(n10132), .C1(
        n8844), .C2(n10130), .ZN(n9074) );
  MUX2_X1 U10255 ( .A(n4540), .B(n9074), .S(n10160), .Z(n8849) );
  AOI22_X1 U10256 ( .A1(n9076), .A2(n10138), .B1(n10140), .B2(n8847), .ZN(
        n8848) );
  OAI211_X1 U10257 ( .C1(n9079), .C2(n8988), .A(n8849), .B(n8848), .ZN(
        P2_U3207) );
  INV_X1 U10258 ( .A(n9083), .ZN(n9009) );
  NOR2_X1 U10259 ( .A1(n9009), .A2(n8981), .ZN(n8856) );
  NAND2_X1 U10260 ( .A1(n8851), .A2(n8850), .ZN(n8852) );
  XOR2_X1 U10261 ( .A(n8859), .B(n8852), .Z(n8853) );
  OAI222_X1 U10262 ( .A1(n10157), .A2(n8855), .B1(n10155), .B2(n8854), .C1(
        n10153), .C2(n8853), .ZN(n9080) );
  AOI211_X1 U10263 ( .C1(n10140), .C2(n8857), .A(n8856), .B(n9080), .ZN(n8861)
         );
  XOR2_X1 U10264 ( .A(n8859), .B(n8858), .Z(n9008) );
  AOI22_X1 U10265 ( .A1(n9008), .A2(n10142), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10162), .ZN(n8860) );
  OAI21_X1 U10266 ( .B1(n8861), .B2(n10162), .A(n8860), .ZN(P2_U3208) );
  INV_X1 U10267 ( .A(n9090), .ZN(n9013) );
  NOR2_X1 U10268 ( .A1(n9013), .A2(n8981), .ZN(n8866) );
  XNOR2_X1 U10269 ( .A(n8862), .B(n8870), .ZN(n8863) );
  OAI222_X1 U10270 ( .A1(n10155), .A2(n8865), .B1(n10157), .B2(n8864), .C1(
        n10153), .C2(n8863), .ZN(n9087) );
  AOI211_X1 U10271 ( .C1(n10140), .C2(n8867), .A(n8866), .B(n9087), .ZN(n8873)
         );
  NAND2_X1 U10272 ( .A1(n8868), .A2(n8869), .ZN(n8871) );
  XNOR2_X1 U10273 ( .A(n8871), .B(n8870), .ZN(n9012) );
  AOI22_X1 U10274 ( .A1(n9012), .A2(n10142), .B1(P2_REG2_REG_24__SCAN_IN), 
        .B2(n10162), .ZN(n8872) );
  OAI21_X1 U10275 ( .B1(n8873), .B2(n10162), .A(n8872), .ZN(P2_U3209) );
  XOR2_X1 U10276 ( .A(n8874), .B(n8875), .Z(n9099) );
  XNOR2_X1 U10277 ( .A(n8876), .B(n8875), .ZN(n8878) );
  AOI222_X1 U10278 ( .A1(n10135), .A2(n8878), .B1(n8905), .B2(n10130), .C1(
        n8877), .C2(n10132), .ZN(n9094) );
  MUX2_X1 U10279 ( .A(n4537), .B(n9094), .S(n10160), .Z(n8881) );
  AOI22_X1 U10280 ( .A1(n9096), .A2(n10138), .B1(n10140), .B2(n8879), .ZN(
        n8880) );
  OAI211_X1 U10281 ( .C1(n9099), .C2(n8988), .A(n8881), .B(n8880), .ZN(
        P2_U3210) );
  XNOR2_X1 U10282 ( .A(n8882), .B(n8885), .ZN(n9022) );
  NAND3_X1 U10283 ( .A1(n8883), .A2(n8885), .A3(n8884), .ZN(n8886) );
  NAND2_X1 U10284 ( .A1(n8887), .A2(n8886), .ZN(n8889) );
  AOI222_X1 U10285 ( .A1(n10135), .A2(n8889), .B1(n8888), .B2(n10132), .C1(
        n8917), .C2(n10130), .ZN(n9021) );
  OR2_X1 U10286 ( .A1(n9021), .A2(n10162), .ZN(n8895) );
  INV_X1 U10287 ( .A(n8890), .ZN(n8891) );
  OAI22_X1 U10288 ( .A1(n10160), .A2(n8892), .B1(n8891), .B2(n10149), .ZN(
        n8893) );
  AOI21_X1 U10289 ( .B1(n9019), .B2(n10138), .A(n8893), .ZN(n8894) );
  OAI211_X1 U10290 ( .C1(n9022), .C2(n8988), .A(n8895), .B(n8894), .ZN(
        P2_U3211) );
  NAND2_X1 U10291 ( .A1(n8912), .A2(n8896), .ZN(n8898) );
  NAND2_X1 U10292 ( .A1(n8898), .A2(n8897), .ZN(n8899) );
  XNOR2_X1 U10293 ( .A(n8899), .B(n8901), .ZN(n9106) );
  INV_X1 U10294 ( .A(n8901), .ZN(n8903) );
  NAND3_X1 U10295 ( .A1(n8900), .A2(n8903), .A3(n8902), .ZN(n8904) );
  NAND2_X1 U10296 ( .A1(n8883), .A2(n8904), .ZN(n8906) );
  AOI222_X1 U10297 ( .A1(n10135), .A2(n8906), .B1(n8933), .B2(n10130), .C1(
        n8905), .C2(n10132), .ZN(n9101) );
  MUX2_X1 U10298 ( .A(n8907), .B(n9101), .S(n10160), .Z(n8910) );
  AOI22_X1 U10299 ( .A1(n9103), .A2(n10138), .B1(n10140), .B2(n8908), .ZN(
        n8909) );
  OAI211_X1 U10300 ( .C1(n9106), .C2(n8988), .A(n8910), .B(n8909), .ZN(
        P2_U3212) );
  XNOR2_X1 U10301 ( .A(n8912), .B(n8911), .ZN(n9112) );
  INV_X1 U10302 ( .A(n8913), .ZN(n8930) );
  OAI21_X1 U10303 ( .B1(n8930), .B2(n8915), .A(n8914), .ZN(n8916) );
  NAND2_X1 U10304 ( .A1(n8916), .A2(n8900), .ZN(n8919) );
  AOI222_X1 U10305 ( .A1(n10135), .A2(n8919), .B1(n8918), .B2(n10130), .C1(
        n8917), .C2(n10132), .ZN(n9107) );
  MUX2_X1 U10306 ( .A(n8920), .B(n9107), .S(n10160), .Z(n8923) );
  AOI22_X1 U10307 ( .A1(n9109), .A2(n10138), .B1(n10140), .B2(n8921), .ZN(
        n8922) );
  OAI211_X1 U10308 ( .C1(n9112), .C2(n8988), .A(n8923), .B(n8922), .ZN(
        P2_U3213) );
  NAND2_X1 U10309 ( .A1(n4971), .A2(n8924), .ZN(n8925) );
  XOR2_X1 U10310 ( .A(n8927), .B(n8925), .Z(n9118) );
  AND2_X1 U10311 ( .A1(n8926), .A2(n10130), .ZN(n8932) );
  AOI21_X1 U10312 ( .B1(n8937), .B2(n8928), .A(n8927), .ZN(n8929) );
  NOR3_X1 U10313 ( .A1(n8930), .A2(n8929), .A3(n10153), .ZN(n8931) );
  AOI211_X1 U10314 ( .C1(n10132), .C2(n8933), .A(n8932), .B(n8931), .ZN(n9113)
         );
  MUX2_X1 U10315 ( .A(n5530), .B(n9113), .S(n10160), .Z(n8936) );
  AOI22_X1 U10316 ( .A1(n9115), .A2(n10138), .B1(n10140), .B2(n8934), .ZN(
        n8935) );
  OAI211_X1 U10317 ( .C1(n9118), .C2(n8988), .A(n8936), .B(n8935), .ZN(
        P2_U3214) );
  INV_X1 U10318 ( .A(n8937), .ZN(n8938) );
  AOI21_X1 U10319 ( .B1(n8940), .B2(n8939), .A(n8938), .ZN(n8941) );
  OAI222_X1 U10320 ( .A1(n10157), .A2(n8943), .B1(n10155), .B2(n8942), .C1(
        n10153), .C2(n8941), .ZN(n9033) );
  INV_X1 U10321 ( .A(n4971), .ZN(n8946) );
  AND2_X1 U10322 ( .A1(n8945), .A2(n8944), .ZN(n9032) );
  NOR3_X1 U10323 ( .A1(n8946), .A2(n9032), .A3(n8988), .ZN(n8951) );
  AOI22_X1 U10324 ( .A1(n10162), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n10140), 
        .B2(n8947), .ZN(n8948) );
  OAI21_X1 U10325 ( .B1(n9123), .B2(n8949), .A(n8948), .ZN(n8950) );
  AOI211_X1 U10326 ( .C1(n9033), .C2(n10160), .A(n8951), .B(n8950), .ZN(n8952)
         );
  INV_X1 U10327 ( .A(n8952), .ZN(P2_U3215) );
  OAI21_X1 U10328 ( .B1(n8955), .B2(n8954), .A(n8953), .ZN(n8956) );
  INV_X1 U10329 ( .A(n8956), .ZN(n9127) );
  XNOR2_X1 U10330 ( .A(n8957), .B(n4575), .ZN(n8958) );
  OAI222_X1 U10331 ( .A1(n10155), .A2(n8960), .B1(n10157), .B2(n8959), .C1(
        n8958), .C2(n10153), .ZN(n9038) );
  NAND2_X1 U10332 ( .A1(n9038), .A2(n10160), .ZN(n8965) );
  OAI22_X1 U10333 ( .A1(n10160), .A2(n8962), .B1(n8961), .B2(n10149), .ZN(
        n8963) );
  AOI21_X1 U10334 ( .B1(n9039), .B2(n10138), .A(n8963), .ZN(n8964) );
  OAI211_X1 U10335 ( .C1(n9127), .C2(n8988), .A(n8965), .B(n8964), .ZN(
        P2_U3216) );
  XNOR2_X1 U10336 ( .A(n8966), .B(n8968), .ZN(n9133) );
  XNOR2_X1 U10337 ( .A(n8967), .B(n8968), .ZN(n8970) );
  AOI222_X1 U10338 ( .A1(n10135), .A2(n8970), .B1(n8969), .B2(n10132), .C1(
        n8978), .C2(n10130), .ZN(n9128) );
  MUX2_X1 U10339 ( .A(n8971), .B(n9128), .S(n10160), .Z(n8975) );
  INV_X1 U10340 ( .A(n8972), .ZN(n8973) );
  AOI22_X1 U10341 ( .A1(n9130), .A2(n10138), .B1(n10140), .B2(n8973), .ZN(
        n8974) );
  OAI211_X1 U10342 ( .C1(n9133), .C2(n8988), .A(n8975), .B(n8974), .ZN(
        P2_U3217) );
  XOR2_X1 U10343 ( .A(n8976), .B(n8986), .Z(n8979) );
  AOI222_X1 U10344 ( .A1(n10135), .A2(n8979), .B1(n8978), .B2(n10132), .C1(
        n8977), .C2(n10130), .ZN(n9134) );
  INV_X1 U10345 ( .A(n9134), .ZN(n8984) );
  OAI22_X1 U10346 ( .A1(n8982), .A2(n8981), .B1(n8980), .B2(n10149), .ZN(n8983) );
  OAI21_X1 U10347 ( .B1(n8984), .B2(n8983), .A(n10160), .ZN(n8990) );
  INV_X1 U10348 ( .A(n8986), .ZN(n8987) );
  XNOR2_X1 U10349 ( .A(n8985), .B(n8987), .ZN(n9139) );
  OR2_X1 U10350 ( .A1(n9139), .A2(n8988), .ZN(n8989) );
  OAI211_X1 U10351 ( .C1(n10160), .C2(n8991), .A(n8990), .B(n8989), .ZN(
        P2_U3219) );
  INV_X1 U10352 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U10353 ( .A1(n9055), .A2(n9050), .ZN(n8992) );
  NAND2_X1 U10354 ( .A1(n9056), .A2(n10243), .ZN(n8994) );
  OAI211_X1 U10355 ( .C1(n10243), .C2(n8993), .A(n8992), .B(n8994), .ZN(
        P2_U3490) );
  NAND2_X1 U10356 ( .A1(n6505), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8995) );
  OAI211_X1 U10357 ( .C1(n8996), .C2(n9037), .A(n8995), .B(n8994), .ZN(
        P2_U3489) );
  MUX2_X1 U10358 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8997), .S(n10243), .Z(
        n9000) );
  OAI22_X1 U10359 ( .A1(n9067), .A2(n9049), .B1(n8998), .B2(n9037), .ZN(n8999)
         );
  OR2_X1 U10360 ( .A1(n9000), .A2(n8999), .ZN(P2_U3487) );
  MUX2_X1 U10361 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9001), .S(n10243), .Z(
        n9004) );
  OAI22_X1 U10362 ( .A1(n9073), .A2(n9049), .B1(n9002), .B2(n9037), .ZN(n9003)
         );
  OR2_X1 U10363 ( .A1(n9004), .A2(n9003), .ZN(P2_U3486) );
  MUX2_X1 U10364 ( .A(n9005), .B(n9074), .S(n10243), .Z(n9007) );
  NAND2_X1 U10365 ( .A1(n9076), .A2(n9050), .ZN(n9006) );
  OAI211_X1 U10366 ( .C1(n9049), .C2(n9079), .A(n9007), .B(n9006), .ZN(
        P2_U3485) );
  MUX2_X1 U10367 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9080), .S(n10243), .Z(
        n9011) );
  INV_X1 U10368 ( .A(n9008), .ZN(n9086) );
  OAI22_X1 U10369 ( .A1(n9086), .A2(n9049), .B1(n9009), .B2(n9037), .ZN(n9010)
         );
  OR2_X1 U10370 ( .A1(n9011), .A2(n9010), .ZN(P2_U3484) );
  MUX2_X1 U10371 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9087), .S(n10243), .Z(
        n9015) );
  INV_X1 U10372 ( .A(n9012), .ZN(n9093) );
  OAI22_X1 U10373 ( .A1(n9093), .A2(n9049), .B1(n9013), .B2(n9037), .ZN(n9014)
         );
  OR2_X1 U10374 ( .A1(n9015), .A2(n9014), .ZN(P2_U3483) );
  INV_X1 U10375 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9016) );
  MUX2_X1 U10376 ( .A(n9016), .B(n9094), .S(n10243), .Z(n9018) );
  NAND2_X1 U10377 ( .A1(n9096), .A2(n9050), .ZN(n9017) );
  OAI211_X1 U10378 ( .C1(n9099), .C2(n9049), .A(n9018), .B(n9017), .ZN(
        P2_U3482) );
  INV_X1 U10379 ( .A(n10196), .ZN(n10215) );
  NAND2_X1 U10380 ( .A1(n9019), .A2(n10221), .ZN(n9020) );
  OAI211_X1 U10381 ( .C1(n10215), .C2(n9022), .A(n9021), .B(n9020), .ZN(n9100)
         );
  MUX2_X1 U10382 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9100), .S(n10243), .Z(
        P2_U3481) );
  INV_X1 U10383 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9023) );
  MUX2_X1 U10384 ( .A(n9023), .B(n9101), .S(n10243), .Z(n9025) );
  NAND2_X1 U10385 ( .A1(n9103), .A2(n9050), .ZN(n9024) );
  OAI211_X1 U10386 ( .C1(n9049), .C2(n9106), .A(n9025), .B(n9024), .ZN(
        P2_U3480) );
  INV_X1 U10387 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9026) );
  MUX2_X1 U10388 ( .A(n9026), .B(n9107), .S(n10243), .Z(n9028) );
  NAND2_X1 U10389 ( .A1(n9109), .A2(n9050), .ZN(n9027) );
  OAI211_X1 U10390 ( .C1(n9049), .C2(n9112), .A(n9028), .B(n9027), .ZN(
        P2_U3479) );
  INV_X1 U10391 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9029) );
  MUX2_X1 U10392 ( .A(n9029), .B(n9113), .S(n10243), .Z(n9031) );
  NAND2_X1 U10393 ( .A1(n9115), .A2(n9050), .ZN(n9030) );
  OAI211_X1 U10394 ( .C1(n9118), .C2(n9049), .A(n9031), .B(n9030), .ZN(
        P2_U3478) );
  NOR2_X1 U10395 ( .A1(n9032), .A2(n10215), .ZN(n9034) );
  AOI21_X1 U10396 ( .B1(n9034), .B2(n4971), .A(n9033), .ZN(n9119) );
  MUX2_X1 U10397 ( .A(n9035), .B(n9119), .S(n10243), .Z(n9036) );
  OAI21_X1 U10398 ( .B1(n9123), .B2(n9037), .A(n9036), .ZN(P2_U3477) );
  AOI21_X1 U10399 ( .B1(n10221), .B2(n9039), .A(n9038), .ZN(n9124) );
  MUX2_X1 U10400 ( .A(n9040), .B(n9124), .S(n10243), .Z(n9041) );
  OAI21_X1 U10401 ( .B1(n9127), .B2(n9049), .A(n9041), .ZN(P2_U3476) );
  INV_X1 U10402 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9042) );
  MUX2_X1 U10403 ( .A(n9042), .B(n9128), .S(n10243), .Z(n9044) );
  NAND2_X1 U10404 ( .A1(n9130), .A2(n9050), .ZN(n9043) );
  OAI211_X1 U10405 ( .C1(n9133), .C2(n9049), .A(n9044), .B(n9043), .ZN(
        P2_U3475) );
  MUX2_X1 U10406 ( .A(n9045), .B(n9134), .S(n10243), .Z(n9047) );
  NAND2_X1 U10407 ( .A1(n9136), .A2(n9050), .ZN(n9046) );
  OAI211_X1 U10408 ( .C1(n9139), .C2(n9049), .A(n9047), .B(n9046), .ZN(
        P2_U3473) );
  INV_X1 U10409 ( .A(n9048), .ZN(n9140) );
  MUX2_X1 U10410 ( .A(n10101), .B(n9140), .S(n10243), .Z(n9053) );
  INV_X1 U10411 ( .A(n9049), .ZN(n9051) );
  AOI22_X1 U10412 ( .A1(n9146), .A2(n9051), .B1(n9050), .B2(n9143), .ZN(n9052)
         );
  NAND2_X1 U10413 ( .A1(n9053), .A2(n9052), .ZN(P2_U3472) );
  MUX2_X1 U10414 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n9054), .S(n10243), .Z(
        P2_U3459) );
  NAND2_X1 U10415 ( .A1(n9055), .A2(n9144), .ZN(n9057) );
  NAND2_X1 U10416 ( .A1(n9056), .A2(n10222), .ZN(n9060) );
  OAI211_X1 U10417 ( .C1(n9058), .C2(n10222), .A(n9057), .B(n9060), .ZN(
        P2_U3458) );
  NAND2_X1 U10418 ( .A1(n9059), .A2(n9144), .ZN(n9061) );
  OAI211_X1 U10419 ( .C1(n6441), .C2(n10222), .A(n9061), .B(n9060), .ZN(
        P2_U3457) );
  MUX2_X1 U10420 ( .A(n9063), .B(n9062), .S(n10222), .Z(n9066) );
  NAND2_X1 U10421 ( .A1(n9064), .A2(n9144), .ZN(n9065) );
  OAI211_X1 U10422 ( .C1(n9067), .C2(n9142), .A(n9066), .B(n9065), .ZN(
        P2_U3455) );
  MUX2_X1 U10423 ( .A(n9069), .B(n9068), .S(n10222), .Z(n9072) );
  NAND2_X1 U10424 ( .A1(n9070), .A2(n9144), .ZN(n9071) );
  OAI211_X1 U10425 ( .C1(n9073), .C2(n9142), .A(n9072), .B(n9071), .ZN(
        P2_U3454) );
  INV_X1 U10426 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9075) );
  MUX2_X1 U10427 ( .A(n9075), .B(n9074), .S(n10222), .Z(n9078) );
  NAND2_X1 U10428 ( .A1(n9076), .A2(n9144), .ZN(n9077) );
  OAI211_X1 U10429 ( .C1(n9079), .C2(n9142), .A(n9078), .B(n9077), .ZN(
        P2_U3453) );
  INV_X1 U10430 ( .A(n9080), .ZN(n9081) );
  MUX2_X1 U10431 ( .A(n9082), .B(n9081), .S(n10222), .Z(n9085) );
  NAND2_X1 U10432 ( .A1(n9083), .A2(n9144), .ZN(n9084) );
  OAI211_X1 U10433 ( .C1(n9086), .C2(n9142), .A(n9085), .B(n9084), .ZN(
        P2_U3452) );
  INV_X1 U10434 ( .A(n9087), .ZN(n9088) );
  MUX2_X1 U10435 ( .A(n9089), .B(n9088), .S(n10222), .Z(n9092) );
  NAND2_X1 U10436 ( .A1(n9090), .A2(n9144), .ZN(n9091) );
  OAI211_X1 U10437 ( .C1(n9093), .C2(n9142), .A(n9092), .B(n9091), .ZN(
        P2_U3451) );
  MUX2_X1 U10438 ( .A(n9095), .B(n9094), .S(n10222), .Z(n9098) );
  NAND2_X1 U10439 ( .A1(n9096), .A2(n9144), .ZN(n9097) );
  OAI211_X1 U10440 ( .C1(n9099), .C2(n9142), .A(n9098), .B(n9097), .ZN(
        P2_U3450) );
  MUX2_X1 U10441 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9100), .S(n10222), .Z(
        P2_U3449) );
  INV_X1 U10442 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n9102) );
  MUX2_X1 U10443 ( .A(n9102), .B(n9101), .S(n10222), .Z(n9105) );
  NAND2_X1 U10444 ( .A1(n9103), .A2(n9144), .ZN(n9104) );
  OAI211_X1 U10445 ( .C1(n9106), .C2(n9142), .A(n9105), .B(n9104), .ZN(
        P2_U3448) );
  INV_X1 U10446 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9108) );
  MUX2_X1 U10447 ( .A(n9108), .B(n9107), .S(n10222), .Z(n9111) );
  NAND2_X1 U10448 ( .A1(n9109), .A2(n9144), .ZN(n9110) );
  OAI211_X1 U10449 ( .C1(n9112), .C2(n9142), .A(n9111), .B(n9110), .ZN(
        P2_U3447) );
  INV_X1 U10450 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9114) );
  MUX2_X1 U10451 ( .A(n9114), .B(n9113), .S(n10222), .Z(n9117) );
  NAND2_X1 U10452 ( .A1(n9115), .A2(n9144), .ZN(n9116) );
  OAI211_X1 U10453 ( .C1(n9118), .C2(n9142), .A(n9117), .B(n9116), .ZN(
        P2_U3446) );
  MUX2_X1 U10454 ( .A(n9120), .B(n9119), .S(n10222), .Z(n9121) );
  OAI21_X1 U10455 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(P2_U3444) );
  MUX2_X1 U10456 ( .A(n9125), .B(n9124), .S(n10222), .Z(n9126) );
  OAI21_X1 U10457 ( .B1(n9127), .B2(n9142), .A(n9126), .ZN(P2_U3441) );
  MUX2_X1 U10458 ( .A(n9129), .B(n9128), .S(n10222), .Z(n9132) );
  NAND2_X1 U10459 ( .A1(n9130), .A2(n9144), .ZN(n9131) );
  OAI211_X1 U10460 ( .C1(n9133), .C2(n9142), .A(n9132), .B(n9131), .ZN(
        P2_U3438) );
  INV_X1 U10461 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9135) );
  MUX2_X1 U10462 ( .A(n9135), .B(n9134), .S(n10222), .Z(n9138) );
  NAND2_X1 U10463 ( .A1(n9136), .A2(n9144), .ZN(n9137) );
  OAI211_X1 U10464 ( .C1(n9139), .C2(n9142), .A(n9138), .B(n9137), .ZN(
        P2_U3432) );
  INV_X1 U10465 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9141) );
  MUX2_X1 U10466 ( .A(n9141), .B(n9140), .S(n10222), .Z(n9148) );
  INV_X1 U10467 ( .A(n9142), .ZN(n9145) );
  AOI22_X1 U10468 ( .A1(n9146), .A2(n9145), .B1(n9144), .B2(n9143), .ZN(n9147)
         );
  NAND2_X1 U10469 ( .A1(n9148), .A2(n9147), .ZN(P2_U3429) );
  MUX2_X1 U10470 ( .A(n9150), .B(P2_D_REG_1__SCAN_IN), .S(n9149), .Z(P2_U3377)
         );
  INV_X1 U10471 ( .A(n9151), .ZN(n9793) );
  NOR4_X1 U10472 ( .A1(n9153), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3151), .A4(
        n9152), .ZN(n9154) );
  AOI21_X1 U10473 ( .B1(n9156), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9154), .ZN(
        n9155) );
  OAI21_X1 U10474 ( .B1(n9793), .B2(n9158), .A(n9155), .ZN(P2_U3264) );
  AOI22_X1 U10475 ( .A1(n6093), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9156), .ZN(n9157) );
  OAI21_X1 U10476 ( .B1(n9159), .B2(n9158), .A(n9157), .ZN(P2_U3265) );
  INV_X1 U10477 ( .A(n9160), .ZN(n9165) );
  NOR3_X1 U10478 ( .A1(n9161), .A2(n9163), .A3(n9162), .ZN(n9164) );
  OAI21_X1 U10479 ( .B1(n9165), .B2(n9164), .A(n9885), .ZN(n9169) );
  AOI22_X1 U10480 ( .A1(n9299), .A2(n9287), .B1(n9286), .B2(n9301), .ZN(n9522)
         );
  OAI22_X1 U10481 ( .A1(n9522), .A2(n9288), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9166), .ZN(n9167) );
  AOI21_X1 U10482 ( .B1(n9528), .B2(n9270), .A(n9167), .ZN(n9168) );
  OAI211_X1 U10483 ( .C1(n9757), .C2(n9280), .A(n9169), .B(n9168), .ZN(
        P1_U3216) );
  NAND2_X1 U10484 ( .A1(n9262), .A2(n9170), .ZN(n9175) );
  XNOR2_X1 U10485 ( .A(n4819), .B(n9172), .ZN(n9285) );
  AOI22_X1 U10486 ( .A1(n9285), .A2(n9173), .B1(n9172), .B2(n9171), .ZN(n9174)
         );
  XOR2_X1 U10487 ( .A(n9175), .B(n9174), .Z(n9182) );
  OAI22_X1 U10488 ( .A1(n9177), .A2(n9275), .B1(n9176), .B2(n9253), .ZN(n9579)
         );
  NOR2_X1 U10489 ( .A1(n9178), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9421) );
  AOI21_X1 U10490 ( .B1(n9579), .B2(n9882), .A(n9421), .ZN(n9179) );
  OAI21_X1 U10491 ( .B1(n9890), .B2(n9583), .A(n9179), .ZN(n9180) );
  AOI21_X1 U10492 ( .B1(n9587), .B2(n9887), .A(n9180), .ZN(n9181) );
  OAI21_X1 U10493 ( .B1(n9182), .B2(n9292), .A(n9181), .ZN(P1_U3219) );
  INV_X1 U10494 ( .A(n9202), .ZN(n9193) );
  NAND2_X1 U10495 ( .A1(n9655), .A2(n9183), .ZN(n9185) );
  OR2_X1 U10496 ( .A1(n9189), .A2(n6545), .ZN(n9184) );
  NAND2_X1 U10497 ( .A1(n9185), .A2(n9184), .ZN(n9187) );
  XNOR2_X1 U10498 ( .A(n9187), .B(n9186), .ZN(n9191) );
  NAND2_X1 U10499 ( .A1(n9655), .A2(n4330), .ZN(n9188) );
  OAI21_X1 U10500 ( .B1(n9189), .B2(n6601), .A(n9188), .ZN(n9190) );
  XNOR2_X1 U10501 ( .A(n9191), .B(n9190), .ZN(n9201) );
  INV_X1 U10502 ( .A(n9201), .ZN(n9192) );
  NAND4_X1 U10503 ( .A1(n9194), .A2(n9193), .A3(n9192), .A4(n9885), .ZN(n9206)
         );
  NAND3_X1 U10504 ( .A1(n9195), .A2(n9885), .A3(n9201), .ZN(n9205) );
  OAI22_X1 U10505 ( .A1(n9197), .A2(n9253), .B1(n9196), .B2(n9275), .ZN(n9445)
         );
  INV_X1 U10506 ( .A(n9445), .ZN(n9199) );
  AOI22_X1 U10507 ( .A1(n9440), .A2(n9270), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n9198) );
  OAI21_X1 U10508 ( .B1(n9199), .B2(n9288), .A(n9198), .ZN(n9200) );
  AOI21_X1 U10509 ( .B1(n9655), .B2(n9887), .A(n9200), .ZN(n9204) );
  NAND3_X1 U10510 ( .A1(n9202), .A2(n9885), .A3(n9201), .ZN(n9203) );
  NAND4_X1 U10511 ( .A1(n9206), .A2(n9205), .A3(n9204), .A4(n9203), .ZN(
        P1_U3220) );
  OAI21_X1 U10512 ( .B1(n9209), .B2(n9208), .A(n9207), .ZN(n9210) );
  NAND2_X1 U10513 ( .A1(n9210), .A2(n9885), .ZN(n9215) );
  INV_X1 U10514 ( .A(n9211), .ZN(n9559) );
  AOI22_X1 U10515 ( .A1(n9301), .A2(n9287), .B1(n9303), .B2(n9286), .ZN(n9554)
         );
  OAI22_X1 U10516 ( .A1(n9554), .A2(n9288), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9212), .ZN(n9213) );
  AOI21_X1 U10517 ( .B1(n9559), .B2(n9270), .A(n9213), .ZN(n9214) );
  OAI211_X1 U10518 ( .C1(n9762), .C2(n9280), .A(n9215), .B(n9214), .ZN(
        P1_U3223) );
  OAI21_X1 U10519 ( .B1(n9217), .B2(n9216), .A(n6752), .ZN(n9218) );
  NAND2_X1 U10520 ( .A1(n9218), .A2(n9885), .ZN(n9225) );
  NAND2_X1 U10521 ( .A1(n9297), .A2(n9287), .ZN(n9220) );
  NAND2_X1 U10522 ( .A1(n9299), .A2(n9286), .ZN(n9219) );
  NAND2_X1 U10523 ( .A1(n9220), .A2(n9219), .ZN(n9489) );
  OAI22_X1 U10524 ( .A1(n9222), .A2(n9890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9221), .ZN(n9223) );
  AOI21_X1 U10525 ( .B1(n9489), .B2(n9882), .A(n9223), .ZN(n9224) );
  OAI211_X1 U10526 ( .C1(n9749), .C2(n9280), .A(n9225), .B(n9224), .ZN(
        P1_U3225) );
  AOI21_X1 U10527 ( .B1(n9227), .B2(n9226), .A(n9237), .ZN(n9233) );
  NAND2_X1 U10528 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9976) );
  NAND2_X1 U10529 ( .A1(n9308), .A2(n9286), .ZN(n9229) );
  NAND2_X1 U10530 ( .A1(n9306), .A2(n9287), .ZN(n9228) );
  NAND2_X1 U10531 ( .A1(n9229), .A2(n9228), .ZN(n9638) );
  NAND2_X1 U10532 ( .A1(n9638), .A2(n9882), .ZN(n9230) );
  OAI211_X1 U10533 ( .C1(n9890), .C2(n9630), .A(n9976), .B(n9230), .ZN(n9231)
         );
  AOI21_X1 U10534 ( .B1(n9628), .B2(n9887), .A(n9231), .ZN(n9232) );
  OAI21_X1 U10535 ( .B1(n9233), .B2(n9292), .A(n9232), .ZN(P1_U3226) );
  INV_X1 U10536 ( .A(n9234), .ZN(n9239) );
  OAI21_X1 U10537 ( .B1(n9237), .B2(n9236), .A(n9235), .ZN(n9238) );
  NAND3_X1 U10538 ( .A1(n9239), .A2(n9885), .A3(n9238), .ZN(n9246) );
  OR2_X1 U10539 ( .A1(n9240), .A2(n9253), .ZN(n9242) );
  NAND2_X1 U10540 ( .A1(n9305), .A2(n9287), .ZN(n9241) );
  NAND2_X1 U10541 ( .A1(n9242), .A2(n9241), .ZN(n9618) );
  NAND2_X1 U10542 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9989) );
  INV_X1 U10543 ( .A(n9989), .ZN(n9244) );
  NOR2_X1 U10544 ( .A1(n9890), .A2(n9611), .ZN(n9243) );
  AOI211_X1 U10545 ( .C1(n9882), .C2(n9618), .A(n9244), .B(n9243), .ZN(n9245)
         );
  OAI211_X1 U10546 ( .C1(n9772), .C2(n9280), .A(n9246), .B(n9245), .ZN(
        P1_U3228) );
  INV_X1 U10547 ( .A(n9247), .ZN(n9251) );
  AND3_X1 U10548 ( .A1(n9160), .A2(n9249), .A3(n9248), .ZN(n9250) );
  OAI21_X1 U10549 ( .B1(n9251), .B2(n9250), .A(n9885), .ZN(n9259) );
  OR2_X1 U10550 ( .A1(n9252), .A2(n9275), .ZN(n9255) );
  OR2_X1 U10551 ( .A1(n9276), .A2(n9253), .ZN(n9254) );
  NAND2_X1 U10552 ( .A1(n9255), .A2(n9254), .ZN(n9511) );
  OAI22_X1 U10553 ( .A1(n9504), .A2(n9890), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9256), .ZN(n9257) );
  AOI21_X1 U10554 ( .B1(n9511), .B2(n9882), .A(n9257), .ZN(n9258) );
  OAI211_X1 U10555 ( .C1(n9753), .C2(n9280), .A(n9259), .B(n9258), .ZN(
        P1_U3229) );
  INV_X1 U10556 ( .A(n9697), .ZN(n9575) );
  INV_X1 U10557 ( .A(n9260), .ZN(n9265) );
  AOI21_X1 U10558 ( .B1(n9263), .B2(n9262), .A(n9261), .ZN(n9264) );
  OAI21_X1 U10559 ( .B1(n9265), .B2(n9264), .A(n9885), .ZN(n9272) );
  INV_X1 U10560 ( .A(n9266), .ZN(n9572) );
  AND2_X1 U10561 ( .A1(n9304), .A2(n9286), .ZN(n9267) );
  AOI21_X1 U10562 ( .B1(n9302), .B2(n9287), .A(n9267), .ZN(n9569) );
  OAI22_X1 U10563 ( .A1(n9569), .A2(n9288), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9268), .ZN(n9269) );
  AOI21_X1 U10564 ( .B1(n9572), .B2(n9270), .A(n9269), .ZN(n9271) );
  OAI211_X1 U10565 ( .C1(n9575), .C2(n9280), .A(n9272), .B(n9271), .ZN(
        P1_U3233) );
  AOI21_X1 U10566 ( .B1(n9274), .B2(n9273), .A(n9161), .ZN(n9284) );
  OR2_X1 U10567 ( .A1(n9276), .A2(n9275), .ZN(n9278) );
  NAND2_X1 U10568 ( .A1(n9302), .A2(n9286), .ZN(n9277) );
  NAND2_X1 U10569 ( .A1(n9278), .A2(n9277), .ZN(n9542) );
  OAI22_X1 U10570 ( .A1(n9890), .A2(n9536), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9279), .ZN(n9282) );
  NOR2_X1 U10571 ( .A1(n9539), .A2(n9280), .ZN(n9281) );
  AOI211_X1 U10572 ( .C1(n9882), .C2(n9542), .A(n9282), .B(n9281), .ZN(n9283)
         );
  OAI21_X1 U10573 ( .B1(n9284), .B2(n9292), .A(n9283), .ZN(P1_U3235) );
  XNOR2_X1 U10574 ( .A(n9285), .B(n4818), .ZN(n9293) );
  NOR2_X1 U10575 ( .A1(n9890), .A2(n9600), .ZN(n9290) );
  AOI22_X1 U10576 ( .A1(n9304), .A2(n9287), .B1(n9306), .B2(n9286), .ZN(n9595)
         );
  NAND2_X1 U10577 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10006)
         );
  OAI21_X1 U10578 ( .B1(n9595), .B2(n9288), .A(n10006), .ZN(n9289) );
  AOI211_X1 U10579 ( .C1(n9708), .C2(n9887), .A(n9290), .B(n9289), .ZN(n9291)
         );
  OAI21_X1 U10580 ( .B1(n9293), .B2(n9292), .A(n9291), .ZN(P1_U3238) );
  MUX2_X1 U10581 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9294), .S(P1_U3973), .Z(
        P1_U3584) );
  MUX2_X1 U10582 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9295), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10583 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9296), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10584 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9297), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10585 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9298), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10586 ( .A(n9299), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9323), .Z(
        P1_U3578) );
  MUX2_X1 U10587 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9300), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10588 ( .A(n9301), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9323), .Z(
        P1_U3576) );
  MUX2_X1 U10589 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9302), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10590 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9303), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10591 ( .A(n9304), .B(P1_DATAO_REG_19__SCAN_IN), .S(n9323), .Z(
        P1_U3573) );
  MUX2_X1 U10592 ( .A(n9305), .B(P1_DATAO_REG_18__SCAN_IN), .S(n9323), .Z(
        P1_U3572) );
  MUX2_X1 U10593 ( .A(n9306), .B(P1_DATAO_REG_17__SCAN_IN), .S(n9323), .Z(
        P1_U3571) );
  MUX2_X1 U10594 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9307), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10595 ( .A(n9308), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9323), .Z(
        P1_U3569) );
  MUX2_X1 U10596 ( .A(n9309), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9323), .Z(
        P1_U3568) );
  MUX2_X1 U10597 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9310), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10598 ( .A(n9311), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9323), .Z(
        P1_U3566) );
  MUX2_X1 U10599 ( .A(n9312), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9323), .Z(
        P1_U3565) );
  MUX2_X1 U10600 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9313), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10601 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9314), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10602 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9315), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10603 ( .A(n9316), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9323), .Z(
        P1_U3561) );
  MUX2_X1 U10604 ( .A(n9317), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9323), .Z(
        P1_U3560) );
  MUX2_X1 U10605 ( .A(n9318), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9323), .Z(
        P1_U3559) );
  MUX2_X1 U10606 ( .A(n9319), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9323), .Z(
        P1_U3558) );
  MUX2_X1 U10607 ( .A(n9320), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9323), .Z(
        P1_U3557) );
  MUX2_X1 U10608 ( .A(n9321), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9323), .Z(
        P1_U3556) );
  MUX2_X1 U10609 ( .A(n9322), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9323), .Z(
        P1_U3555) );
  MUX2_X1 U10610 ( .A(n9324), .B(P1_DATAO_REG_0__SCAN_IN), .S(n9323), .Z(
        P1_U3554) );
  INV_X1 U10611 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9326) );
  OAI22_X1 U10612 ( .A1(n10008), .A2(n9326), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9325), .ZN(n9327) );
  AOI21_X1 U10613 ( .B1(n10005), .B2(n4336), .A(n9327), .ZN(n9337) );
  INV_X1 U10614 ( .A(n9999), .ZN(n9987) );
  OAI211_X1 U10615 ( .C1(n9331), .C2(n9330), .A(n9987), .B(n9329), .ZN(n9336)
         );
  INV_X1 U10616 ( .A(n9993), .ZN(n9986) );
  OAI211_X1 U10617 ( .C1(n9334), .C2(n9333), .A(n9986), .B(n9332), .ZN(n9335)
         );
  NAND3_X1 U10618 ( .A1(n9337), .A2(n9336), .A3(n9335), .ZN(P1_U3244) );
  INV_X1 U10619 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9339) );
  OAI22_X1 U10620 ( .A1(n10008), .A2(n9339), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9338), .ZN(n9340) );
  AOI21_X1 U10621 ( .B1(n10005), .B2(n9341), .A(n9340), .ZN(n9350) );
  OAI211_X1 U10622 ( .C1(n9344), .C2(n9343), .A(n9986), .B(n9342), .ZN(n9349)
         );
  OAI211_X1 U10623 ( .C1(n9347), .C2(n9346), .A(n9987), .B(n9345), .ZN(n9348)
         );
  NAND4_X1 U10624 ( .A1(n9351), .A2(n9350), .A3(n9349), .A4(n9348), .ZN(
        P1_U3245) );
  INV_X1 U10625 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U10626 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_U3086), .ZN(n9352) );
  OAI21_X1 U10627 ( .B1(n10008), .B2(n9798), .A(n9352), .ZN(n9353) );
  AOI21_X1 U10628 ( .B1(n10005), .B2(n9354), .A(n9353), .ZN(n9363) );
  OAI211_X1 U10629 ( .C1(n9357), .C2(n9356), .A(n9986), .B(n9355), .ZN(n9362)
         );
  OAI211_X1 U10630 ( .C1(n9360), .C2(n9359), .A(n9987), .B(n9358), .ZN(n9361)
         );
  NAND3_X1 U10631 ( .A1(n9363), .A2(n9362), .A3(n9361), .ZN(P1_U3246) );
  XNOR2_X1 U10632 ( .A(n9400), .B(n9364), .ZN(n9367) );
  NAND2_X1 U10633 ( .A1(n9366), .A2(n9367), .ZN(n9382) );
  OAI21_X1 U10634 ( .B1(n9367), .B2(n9366), .A(n9382), .ZN(n9368) );
  NAND2_X1 U10635 ( .A1(n9368), .A2(n9987), .ZN(n9379) );
  MUX2_X1 U10636 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n9371), .S(n9400), .Z(n9372)
         );
  NAND2_X1 U10637 ( .A1(n9373), .A2(n9372), .ZN(n9399) );
  OAI21_X1 U10638 ( .B1(n9373), .B2(n9372), .A(n9399), .ZN(n9374) );
  NAND2_X1 U10639 ( .A1(n9374), .A2(n9986), .ZN(n9378) );
  AOI21_X1 U10640 ( .B1(n9422), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9375), .ZN(
        n9377) );
  NAND2_X1 U10641 ( .A1(n10005), .A2(n9400), .ZN(n9376) );
  NAND4_X1 U10642 ( .A1(n9379), .A2(n9378), .A3(n9377), .A4(n9376), .ZN(
        P1_U3252) );
  XNOR2_X1 U10643 ( .A(n9919), .B(n9380), .ZN(n9920) );
  NOR2_X1 U10644 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n9903), .ZN(n9381) );
  AOI21_X1 U10645 ( .B1(n9903), .B2(P1_REG2_REG_12__SCAN_IN), .A(n9381), .ZN(
        n9910) );
  OAI21_X1 U10646 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9400), .A(n9382), .ZN(
        n9850) );
  NAND2_X1 U10647 ( .A1(n9853), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n9383) );
  OAI21_X1 U10648 ( .B1(n9853), .B2(P1_REG2_REG_10__SCAN_IN), .A(n9383), .ZN(
        n9849) );
  NOR2_X1 U10649 ( .A1(n9850), .A2(n9849), .ZN(n9848) );
  NAND2_X1 U10650 ( .A1(n9899), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9384) );
  OAI21_X1 U10651 ( .B1(n9899), .B2(P1_REG2_REG_11__SCAN_IN), .A(n9384), .ZN(
        n9892) );
  NOR2_X1 U10652 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  AOI21_X1 U10653 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n9899), .A(n9891), .ZN(
        n9909) );
  NAND2_X1 U10654 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  OAI21_X1 U10655 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9903), .A(n9908), .ZN(
        n9921) );
  INV_X1 U10656 ( .A(n9921), .ZN(n9385) );
  NAND2_X1 U10657 ( .A1(n9920), .A2(n9385), .ZN(n9924) );
  NAND2_X1 U10658 ( .A1(n9919), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n9386) );
  NAND2_X1 U10659 ( .A1(P1_REG2_REG_14__SCAN_IN), .A2(n9407), .ZN(n9387) );
  OAI21_X1 U10660 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n9407), .A(n9387), .ZN(
        n9938) );
  NOR2_X1 U10661 ( .A1(n9388), .A2(n9409), .ZN(n9389) );
  XNOR2_X1 U10662 ( .A(n9973), .B(n9631), .ZN(n9967) );
  NAND2_X1 U10663 ( .A1(n9390), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n9391) );
  XNOR2_X1 U10664 ( .A(n9984), .B(n9612), .ZN(n9981) );
  NAND2_X1 U10665 ( .A1(n9980), .A2(n9981), .ZN(n9979) );
  OR2_X1 U10666 ( .A1(n9984), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U10667 ( .A1(n10004), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n9394) );
  OAI21_X1 U10668 ( .B1(n10004), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9394), .ZN(
        n10001) );
  INV_X1 U10669 ( .A(n10001), .ZN(n9393) );
  NAND2_X1 U10670 ( .A1(n9997), .A2(n9394), .ZN(n9395) );
  XNOR2_X1 U10671 ( .A(n9395), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9416) );
  INV_X1 U10672 ( .A(n9416), .ZN(n9415) );
  OR2_X1 U10673 ( .A1(n9919), .A2(n9396), .ZN(n9398) );
  NAND2_X1 U10674 ( .A1(n9919), .A2(n9396), .ZN(n9397) );
  NAND2_X1 U10675 ( .A1(n9398), .A2(n9397), .ZN(n9927) );
  OR2_X1 U10676 ( .A1(n9903), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n9404) );
  OAI21_X1 U10677 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9400), .A(n9399), .ZN(
        n9846) );
  MUX2_X1 U10678 ( .A(n9401), .B(P1_REG1_REG_10__SCAN_IN), .S(n9853), .Z(n9847) );
  NOR2_X1 U10679 ( .A1(n9846), .A2(n9847), .ZN(n9845) );
  MUX2_X1 U10680 ( .A(n9402), .B(P1_REG1_REG_11__SCAN_IN), .S(n9899), .Z(n9895) );
  NOR2_X1 U10681 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  MUX2_X1 U10682 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9403), .S(n9903), .Z(n9905) );
  NAND2_X1 U10683 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  NAND2_X1 U10684 ( .A1(n9927), .A2(n9928), .ZN(n9926) );
  NAND2_X1 U10685 ( .A1(n9919), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n9405) );
  NAND2_X1 U10686 ( .A1(n9926), .A2(n9405), .ZN(n9943) );
  XNOR2_X1 U10687 ( .A(n9407), .B(n9406), .ZN(n9944) );
  NOR2_X1 U10688 ( .A1(n9408), .A2(n9409), .ZN(n9410) );
  XNOR2_X1 U10689 ( .A(n9409), .B(n9408), .ZN(n9955) );
  NOR2_X1 U10690 ( .A1(n9410), .A2(n9953), .ZN(n9965) );
  XNOR2_X1 U10691 ( .A(n9973), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9964) );
  AOI22_X1 U10692 ( .A1(n9965), .A2(n9964), .B1(n9719), .B2(n9973), .ZN(n9983)
         );
  XNOR2_X1 U10693 ( .A(n9984), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9982) );
  OAI22_X1 U10694 ( .A1(n9983), .A2(n9982), .B1(n9984), .B2(
        P1_REG1_REG_17__SCAN_IN), .ZN(n9995) );
  NAND2_X1 U10695 ( .A1(n10004), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n9411) );
  OAI21_X1 U10696 ( .B1(n10004), .B2(P1_REG1_REG_18__SCAN_IN), .A(n9411), .ZN(
        n9994) );
  NOR2_X1 U10697 ( .A1(n9995), .A2(n9994), .ZN(n9992) );
  INV_X1 U10698 ( .A(n9411), .ZN(n9412) );
  NOR2_X1 U10699 ( .A1(n9992), .A2(n9412), .ZN(n9413) );
  XNOR2_X1 U10700 ( .A(n9413), .B(n9704), .ZN(n9417) );
  NAND2_X1 U10701 ( .A1(n9417), .A2(n9986), .ZN(n9414) );
  OAI22_X1 U10702 ( .A1(n9417), .A2(n9993), .B1(n9416), .B2(n9999), .ZN(n9419)
         );
  AOI211_X1 U10703 ( .C1(P1_ADDR_REG_19__SCAN_IN), .C2(n9422), .A(n9421), .B(
        n9420), .ZN(n9423) );
  INV_X1 U10704 ( .A(n9423), .ZN(P1_U3262) );
  NAND2_X1 U10705 ( .A1(n9424), .A2(n10015), .ZN(n9427) );
  INV_X1 U10706 ( .A(n9647), .ZN(n9425) );
  NOR2_X1 U10707 ( .A1(n9425), .A2(n10033), .ZN(n9433) );
  AOI21_X1 U10708 ( .B1(n10033), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9433), .ZN(
        n9426) );
  OAI211_X1 U10709 ( .C1(n9646), .C2(n9629), .A(n9427), .B(n9426), .ZN(
        P1_U3263) );
  INV_X1 U10710 ( .A(n9428), .ZN(n9431) );
  INV_X1 U10711 ( .A(n9429), .ZN(n9430) );
  NAND2_X1 U10712 ( .A1(n9648), .A2(n10015), .ZN(n9435) );
  AOI21_X1 U10713 ( .B1(n10033), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9433), .ZN(
        n9434) );
  OAI211_X1 U10714 ( .C1(n4472), .C2(n9629), .A(n9435), .B(n9434), .ZN(
        P1_U3264) );
  AOI21_X1 U10715 ( .B1(n9655), .B2(n9458), .A(n4600), .ZN(n9656) );
  INV_X1 U10716 ( .A(n9655), .ZN(n9442) );
  AOI22_X1 U10717 ( .A1(n9440), .A2(n10032), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n10033), .ZN(n9441) );
  OAI21_X1 U10718 ( .B1(n9442), .B2(n9629), .A(n9441), .ZN(n9448) );
  XNOR2_X1 U10719 ( .A(n9444), .B(n9443), .ZN(n9446) );
  NOR2_X1 U10720 ( .A1(n9658), .A2(n10045), .ZN(n9447) );
  AOI211_X1 U10721 ( .C1(n9656), .C2(n9547), .A(n9448), .B(n9447), .ZN(n9449)
         );
  OAI21_X1 U10722 ( .B1(n9659), .B2(n10020), .A(n9449), .ZN(P1_U3265) );
  XNOR2_X1 U10723 ( .A(n9450), .B(n9453), .ZN(n9662) );
  INV_X1 U10724 ( .A(n9662), .ZN(n9468) );
  OAI21_X1 U10725 ( .B1(n9453), .B2(n9452), .A(n9451), .ZN(n9454) );
  NAND2_X1 U10726 ( .A1(n9454), .A2(n9636), .ZN(n9457) );
  INV_X1 U10727 ( .A(n9455), .ZN(n9456) );
  NAND2_X1 U10728 ( .A1(n9457), .A2(n9456), .ZN(n9660) );
  INV_X1 U10729 ( .A(n9476), .ZN(n9460) );
  INV_X1 U10730 ( .A(n9458), .ZN(n9459) );
  AOI211_X1 U10731 ( .C1(n9461), .C2(n9460), .A(n9627), .B(n9459), .ZN(n9661)
         );
  NAND2_X1 U10732 ( .A1(n9661), .A2(n10015), .ZN(n9465) );
  INV_X1 U10733 ( .A(n9462), .ZN(n9463) );
  AOI22_X1 U10734 ( .A1(n9463), .A2(n10032), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n10033), .ZN(n9464) );
  OAI211_X1 U10735 ( .C1(n9741), .C2(n9629), .A(n9465), .B(n9464), .ZN(n9466)
         );
  AOI21_X1 U10736 ( .B1(n9660), .B2(n10023), .A(n9466), .ZN(n9467) );
  OAI21_X1 U10737 ( .B1(n9468), .B2(n10020), .A(n9467), .ZN(P1_U3266) );
  XNOR2_X1 U10738 ( .A(n9469), .B(n9470), .ZN(n9667) );
  INV_X1 U10739 ( .A(n9667), .ZN(n9484) );
  XNOR2_X1 U10740 ( .A(n9471), .B(n9470), .ZN(n9472) );
  NAND2_X1 U10741 ( .A1(n9472), .A2(n9636), .ZN(n9475) );
  INV_X1 U10742 ( .A(n9473), .ZN(n9474) );
  NAND2_X1 U10743 ( .A1(n9475), .A2(n9474), .ZN(n9665) );
  INV_X1 U10744 ( .A(n9492), .ZN(n9477) );
  AOI211_X1 U10745 ( .C1(n9478), .C2(n9477), .A(n9627), .B(n9476), .ZN(n9666)
         );
  NAND2_X1 U10746 ( .A1(n9666), .A2(n10015), .ZN(n9481) );
  AOI22_X1 U10747 ( .A1(n9479), .A2(n10032), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n10033), .ZN(n9480) );
  OAI211_X1 U10748 ( .C1(n9745), .C2(n9629), .A(n9481), .B(n9480), .ZN(n9482)
         );
  AOI21_X1 U10749 ( .B1(n10023), .B2(n9665), .A(n9482), .ZN(n9483) );
  OAI21_X1 U10750 ( .B1(n9484), .B2(n10020), .A(n9483), .ZN(P1_U3267) );
  XNOR2_X1 U10751 ( .A(n9485), .B(n9487), .ZN(n9672) );
  INV_X1 U10752 ( .A(n9672), .ZN(n9499) );
  OAI211_X1 U10753 ( .C1(n9488), .C2(n9487), .A(n9486), .B(n9636), .ZN(n9491)
         );
  INV_X1 U10754 ( .A(n9489), .ZN(n9490) );
  NAND2_X1 U10755 ( .A1(n9491), .A2(n9490), .ZN(n9670) );
  AOI211_X1 U10756 ( .C1(n9493), .C2(n9501), .A(n9627), .B(n9492), .ZN(n9671)
         );
  NAND2_X1 U10757 ( .A1(n9671), .A2(n10015), .ZN(n9496) );
  AOI22_X1 U10758 ( .A1(n9494), .A2(n10032), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n10033), .ZN(n9495) );
  OAI211_X1 U10759 ( .C1(n9749), .C2(n9629), .A(n9496), .B(n9495), .ZN(n9497)
         );
  AOI21_X1 U10760 ( .B1(n10023), .B2(n9670), .A(n9497), .ZN(n9498) );
  OAI21_X1 U10761 ( .B1(n9499), .B2(n10020), .A(n9498), .ZN(P1_U3268) );
  XNOR2_X1 U10762 ( .A(n9500), .B(n9507), .ZN(n9677) );
  INV_X1 U10763 ( .A(n9677), .ZN(n9516) );
  AOI211_X1 U10764 ( .C1(n9502), .C2(n9524), .A(n9627), .B(n4578), .ZN(n9676)
         );
  NOR2_X1 U10765 ( .A1(n9753), .A2(n9629), .ZN(n9506) );
  OAI22_X1 U10766 ( .A1(n9504), .A2(n10021), .B1(n9503), .B2(n10023), .ZN(
        n9505) );
  AOI211_X1 U10767 ( .C1(n9676), .C2(n10015), .A(n9506), .B(n9505), .ZN(n9515)
         );
  NAND2_X1 U10768 ( .A1(n9508), .A2(n9507), .ZN(n9509) );
  NAND3_X1 U10769 ( .A1(n9510), .A2(n9636), .A3(n9509), .ZN(n9513) );
  INV_X1 U10770 ( .A(n9511), .ZN(n9512) );
  NAND2_X1 U10771 ( .A1(n9513), .A2(n9512), .ZN(n9675) );
  NAND2_X1 U10772 ( .A1(n9675), .A2(n10023), .ZN(n9514) );
  OAI211_X1 U10773 ( .C1(n9516), .C2(n10020), .A(n9515), .B(n9514), .ZN(
        P1_U3269) );
  XNOR2_X1 U10774 ( .A(n9518), .B(n9517), .ZN(n9682) );
  INV_X1 U10775 ( .A(n9682), .ZN(n9533) );
  XNOR2_X1 U10776 ( .A(n9520), .B(n9519), .ZN(n9521) );
  NAND2_X1 U10777 ( .A1(n9521), .A2(n9636), .ZN(n9523) );
  NAND2_X1 U10778 ( .A1(n9523), .A2(n9522), .ZN(n9680) );
  INV_X1 U10779 ( .A(n9535), .ZN(n9526) );
  INV_X1 U10780 ( .A(n9524), .ZN(n9525) );
  AOI211_X1 U10781 ( .C1(n9527), .C2(n9526), .A(n9627), .B(n9525), .ZN(n9681)
         );
  NAND2_X1 U10782 ( .A1(n9681), .A2(n10015), .ZN(n9530) );
  AOI22_X1 U10783 ( .A1(n9528), .A2(n10032), .B1(P1_REG2_REG_23__SCAN_IN), 
        .B2(n10033), .ZN(n9529) );
  OAI211_X1 U10784 ( .C1(n9757), .C2(n9629), .A(n9530), .B(n9529), .ZN(n9531)
         );
  AOI21_X1 U10785 ( .B1(n10023), .B2(n9680), .A(n9531), .ZN(n9532) );
  OAI21_X1 U10786 ( .B1(n9533), .B2(n10020), .A(n9532), .ZN(P1_U3270) );
  XOR2_X1 U10787 ( .A(n9534), .B(n9540), .Z(n9689) );
  AOI21_X1 U10788 ( .B1(n9685), .B2(n9556), .A(n9535), .ZN(n9686) );
  INV_X1 U10789 ( .A(n9536), .ZN(n9537) );
  AOI22_X1 U10790 ( .A1(n9537), .A2(n10032), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n10033), .ZN(n9538) );
  OAI21_X1 U10791 ( .B1(n9539), .B2(n9629), .A(n9538), .ZN(n9546) );
  INV_X1 U10792 ( .A(n9540), .ZN(n9541) );
  AOI21_X1 U10793 ( .B1(n9541), .B2(n4408), .A(n9596), .ZN(n9544) );
  AOI21_X1 U10794 ( .B1(n9544), .B2(n9543), .A(n9542), .ZN(n9688) );
  NOR2_X1 U10795 ( .A1(n9688), .A2(n10045), .ZN(n9545) );
  AOI211_X1 U10796 ( .C1(n9686), .C2(n9547), .A(n9546), .B(n9545), .ZN(n9548)
         );
  OAI21_X1 U10797 ( .B1(n9689), .B2(n10020), .A(n9548), .ZN(P1_U3271) );
  XOR2_X1 U10798 ( .A(n9551), .B(n9549), .Z(n9692) );
  INV_X1 U10799 ( .A(n9692), .ZN(n9564) );
  OAI21_X1 U10800 ( .B1(n9568), .B2(n9565), .A(n9550), .ZN(n9552) );
  XNOR2_X1 U10801 ( .A(n9552), .B(n9551), .ZN(n9553) );
  NAND2_X1 U10802 ( .A1(n9553), .A2(n9636), .ZN(n9555) );
  NAND2_X1 U10803 ( .A1(n9555), .A2(n9554), .ZN(n9690) );
  INV_X1 U10804 ( .A(n9556), .ZN(n9557) );
  AOI211_X1 U10805 ( .C1(n9558), .C2(n9571), .A(n9627), .B(n9557), .ZN(n9691)
         );
  NAND2_X1 U10806 ( .A1(n9691), .A2(n10015), .ZN(n9561) );
  AOI22_X1 U10807 ( .A1(n9559), .A2(n10032), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n10033), .ZN(n9560) );
  OAI211_X1 U10808 ( .C1(n9762), .C2(n9629), .A(n9561), .B(n9560), .ZN(n9562)
         );
  AOI21_X1 U10809 ( .B1(n10023), .B2(n9690), .A(n9562), .ZN(n9563) );
  OAI21_X1 U10810 ( .B1(n9564), .B2(n10020), .A(n9563), .ZN(P1_U3272) );
  XNOR2_X1 U10811 ( .A(n9566), .B(n9565), .ZN(n9699) );
  XNOR2_X1 U10812 ( .A(n9568), .B(n9567), .ZN(n9570) );
  OAI21_X1 U10813 ( .B1(n9570), .B2(n9596), .A(n9569), .ZN(n9696) );
  AOI211_X1 U10814 ( .C1(n9697), .C2(n4350), .A(n9627), .B(n4585), .ZN(n9695)
         );
  NAND2_X1 U10815 ( .A1(n9695), .A2(n10015), .ZN(n9574) );
  AOI22_X1 U10816 ( .A1(n9572), .A2(n10032), .B1(n10033), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9573) );
  OAI211_X1 U10817 ( .C1(n9575), .C2(n9629), .A(n9574), .B(n9573), .ZN(n9576)
         );
  AOI21_X1 U10818 ( .B1(n10023), .B2(n9696), .A(n9576), .ZN(n9577) );
  OAI21_X1 U10819 ( .B1(n9699), .B2(n10020), .A(n9577), .ZN(P1_U3273) );
  XNOR2_X1 U10820 ( .A(n9578), .B(n9581), .ZN(n9580) );
  AOI21_X1 U10821 ( .B1(n9580), .B2(n9636), .A(n9579), .ZN(n9701) );
  XOR2_X1 U10822 ( .A(n9582), .B(n9581), .Z(n9702) );
  OR2_X1 U10823 ( .A1(n9702), .A2(n10020), .ZN(n9589) );
  OAI22_X1 U10824 ( .A1(n10023), .A2(n9584), .B1(n9583), .B2(n10021), .ZN(
        n9586) );
  OAI211_X1 U10825 ( .C1(n9598), .C2(n9767), .A(n10058), .B(n4350), .ZN(n9700)
         );
  NOR2_X1 U10826 ( .A1(n9700), .A2(n10038), .ZN(n9585) );
  AOI211_X1 U10827 ( .C1(n10035), .C2(n9587), .A(n9586), .B(n9585), .ZN(n9588)
         );
  OAI211_X1 U10828 ( .C1(n10033), .C2(n9701), .A(n9589), .B(n9588), .ZN(
        P1_U3274) );
  XNOR2_X1 U10829 ( .A(n9590), .B(n9594), .ZN(n9710) );
  NAND2_X1 U10830 ( .A1(n9592), .A2(n9591), .ZN(n9593) );
  XOR2_X1 U10831 ( .A(n9594), .B(n9593), .Z(n9597) );
  OAI21_X1 U10832 ( .B1(n9597), .B2(n9596), .A(n9595), .ZN(n9707) );
  INV_X1 U10833 ( .A(n9609), .ZN(n9599) );
  AOI211_X1 U10834 ( .C1(n9708), .C2(n9599), .A(n9627), .B(n9598), .ZN(n9706)
         );
  NAND2_X1 U10835 ( .A1(n9706), .A2(n10015), .ZN(n9603) );
  INV_X1 U10836 ( .A(n9600), .ZN(n9601) );
  AOI22_X1 U10837 ( .A1(n10033), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9601), 
        .B2(n10032), .ZN(n9602) );
  OAI211_X1 U10838 ( .C1(n9604), .C2(n9629), .A(n9603), .B(n9602), .ZN(n9605)
         );
  AOI21_X1 U10839 ( .B1(n10023), .B2(n9707), .A(n9605), .ZN(n9606) );
  OAI21_X1 U10840 ( .B1(n9710), .B2(n10020), .A(n9606), .ZN(P1_U3275) );
  XNOR2_X1 U10841 ( .A(n9608), .B(n9607), .ZN(n9713) );
  INV_X1 U10842 ( .A(n9713), .ZN(n9623) );
  AOI211_X1 U10843 ( .C1(n9610), .C2(n9625), .A(n9627), .B(n9609), .ZN(n9712)
         );
  NOR2_X1 U10844 ( .A1(n9772), .A2(n9629), .ZN(n9614) );
  OAI22_X1 U10845 ( .A1(n10023), .A2(n9612), .B1(n9611), .B2(n10021), .ZN(
        n9613) );
  AOI211_X1 U10846 ( .C1(n9712), .C2(n10015), .A(n9614), .B(n9613), .ZN(n9622)
         );
  XNOR2_X1 U10847 ( .A(n9616), .B(n9615), .ZN(n9617) );
  NAND2_X1 U10848 ( .A1(n9617), .A2(n9636), .ZN(n9620) );
  INV_X1 U10849 ( .A(n9618), .ZN(n9619) );
  NAND2_X1 U10850 ( .A1(n9620), .A2(n9619), .ZN(n9711) );
  NAND2_X1 U10851 ( .A1(n9711), .A2(n10023), .ZN(n9621) );
  OAI211_X1 U10852 ( .C1(n9623), .C2(n10020), .A(n9622), .B(n9621), .ZN(
        P1_U3276) );
  XNOR2_X1 U10853 ( .A(n9624), .B(n9634), .ZN(n9718) );
  INV_X1 U10854 ( .A(n9718), .ZN(n9643) );
  INV_X1 U10855 ( .A(n9625), .ZN(n9626) );
  AOI211_X1 U10856 ( .C1(n9628), .C2(n8195), .A(n9627), .B(n9626), .ZN(n9717)
         );
  INV_X1 U10857 ( .A(n9628), .ZN(n9776) );
  NOR2_X1 U10858 ( .A1(n9776), .A2(n9629), .ZN(n9633) );
  OAI22_X1 U10859 ( .A1(n10023), .A2(n9631), .B1(n9630), .B2(n10021), .ZN(
        n9632) );
  AOI211_X1 U10860 ( .C1(n9717), .C2(n10015), .A(n9633), .B(n9632), .ZN(n9642)
         );
  XNOR2_X1 U10861 ( .A(n9635), .B(n9634), .ZN(n9637) );
  NAND2_X1 U10862 ( .A1(n9637), .A2(n9636), .ZN(n9640) );
  INV_X1 U10863 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U10864 ( .A1(n9640), .A2(n9639), .ZN(n9716) );
  NAND2_X1 U10865 ( .A1(n9716), .A2(n10023), .ZN(n9641) );
  OAI211_X1 U10866 ( .C1(n9643), .C2(n10020), .A(n9642), .B(n9641), .ZN(
        P1_U3277) );
  OAI21_X1 U10867 ( .B1(n9646), .B2(n9726), .A(n9645), .ZN(P1_U3553) );
  NOR2_X1 U10868 ( .A1(n9648), .A2(n9647), .ZN(n9733) );
  MUX2_X1 U10869 ( .A(n5937), .B(n9733), .S(n10082), .Z(n9649) );
  OAI21_X1 U10870 ( .B1(n4472), .B2(n9726), .A(n9649), .ZN(P1_U3552) );
  AOI22_X1 U10871 ( .A1(n9651), .A2(n10058), .B1(n10057), .B2(n9650), .ZN(
        n9652) );
  OAI21_X1 U10872 ( .B1(n9654), .B2(n10062), .A(n9653), .ZN(n9736) );
  MUX2_X1 U10873 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9736), .S(n10082), .Z(
        P1_U3551) );
  AOI22_X1 U10874 ( .A1(n9656), .A2(n10058), .B1(n10057), .B2(n9655), .ZN(
        n9657) );
  OAI211_X1 U10875 ( .C1(n9659), .C2(n10062), .A(n9658), .B(n9657), .ZN(n9737)
         );
  MUX2_X1 U10876 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9737), .S(n10082), .Z(
        P1_U3550) );
  MUX2_X1 U10877 ( .A(n9663), .B(n9738), .S(n10082), .Z(n9664) );
  OAI21_X1 U10878 ( .B1(n9741), .B2(n9726), .A(n9664), .ZN(P1_U3549) );
  MUX2_X1 U10879 ( .A(n9668), .B(n9742), .S(n10082), .Z(n9669) );
  OAI21_X1 U10880 ( .B1(n9745), .B2(n9726), .A(n9669), .ZN(P1_U3548) );
  MUX2_X1 U10881 ( .A(n9673), .B(n9746), .S(n10082), .Z(n9674) );
  OAI21_X1 U10882 ( .B1(n9749), .B2(n9726), .A(n9674), .ZN(P1_U3547) );
  INV_X1 U10883 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9678) );
  AOI211_X1 U10884 ( .C1(n9677), .C2(n9723), .A(n9676), .B(n9675), .ZN(n9750)
         );
  MUX2_X1 U10885 ( .A(n9678), .B(n9750), .S(n10082), .Z(n9679) );
  OAI21_X1 U10886 ( .B1(n9753), .B2(n9726), .A(n9679), .ZN(P1_U3546) );
  AOI211_X1 U10887 ( .C1(n9682), .C2(n9723), .A(n9681), .B(n9680), .ZN(n9754)
         );
  MUX2_X1 U10888 ( .A(n9683), .B(n9754), .S(n10082), .Z(n9684) );
  OAI21_X1 U10889 ( .B1(n9757), .B2(n9726), .A(n9684), .ZN(P1_U3545) );
  AOI22_X1 U10890 ( .A1(n9686), .A2(n10058), .B1(n10057), .B2(n9685), .ZN(
        n9687) );
  OAI211_X1 U10891 ( .C1(n9689), .C2(n10062), .A(n9688), .B(n9687), .ZN(n9758)
         );
  MUX2_X1 U10892 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9758), .S(n10082), .Z(
        P1_U3544) );
  INV_X1 U10893 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n9693) );
  AOI211_X1 U10894 ( .C1(n9692), .C2(n9723), .A(n9691), .B(n9690), .ZN(n9759)
         );
  MUX2_X1 U10895 ( .A(n9693), .B(n9759), .S(n10082), .Z(n9694) );
  OAI21_X1 U10896 ( .B1(n9762), .B2(n9726), .A(n9694), .ZN(P1_U3543) );
  AOI211_X1 U10897 ( .C1(n10057), .C2(n9697), .A(n9696), .B(n9695), .ZN(n9698)
         );
  OAI21_X1 U10898 ( .B1(n9699), .B2(n10062), .A(n9698), .ZN(n9763) );
  MUX2_X1 U10899 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9763), .S(n10082), .Z(
        P1_U3542) );
  OAI211_X1 U10900 ( .C1(n9702), .C2(n10062), .A(n9701), .B(n9700), .ZN(n9703)
         );
  INV_X1 U10901 ( .A(n9703), .ZN(n9764) );
  MUX2_X1 U10902 ( .A(n9704), .B(n9764), .S(n10082), .Z(n9705) );
  OAI21_X1 U10903 ( .B1(n9767), .B2(n9726), .A(n9705), .ZN(P1_U3541) );
  AOI211_X1 U10904 ( .C1(n10057), .C2(n9708), .A(n9707), .B(n9706), .ZN(n9709)
         );
  OAI21_X1 U10905 ( .B1(n9710), .B2(n10062), .A(n9709), .ZN(n9768) );
  MUX2_X1 U10906 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9768), .S(n10082), .Z(
        P1_U3540) );
  AOI211_X1 U10907 ( .C1(n9713), .C2(n9723), .A(n9712), .B(n9711), .ZN(n9769)
         );
  MUX2_X1 U10908 ( .A(n9714), .B(n9769), .S(n10082), .Z(n9715) );
  OAI21_X1 U10909 ( .B1(n9772), .B2(n9726), .A(n9715), .ZN(P1_U3539) );
  AOI211_X1 U10910 ( .C1(n9718), .C2(n9723), .A(n9717), .B(n9716), .ZN(n9773)
         );
  MUX2_X1 U10911 ( .A(n9719), .B(n9773), .S(n10082), .Z(n9720) );
  OAI21_X1 U10912 ( .B1(n9776), .B2(n9726), .A(n9720), .ZN(P1_U3538) );
  AOI211_X1 U10913 ( .C1(n9724), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9777)
         );
  MUX2_X1 U10914 ( .A(n9954), .B(n9777), .S(n10082), .Z(n9725) );
  OAI21_X1 U10915 ( .B1(n9781), .B2(n9726), .A(n9725), .ZN(P1_U3537) );
  AOI21_X1 U10916 ( .B1(n10057), .B2(n9728), .A(n9727), .ZN(n9729) );
  OAI211_X1 U10917 ( .C1(n9731), .C2(n10062), .A(n9730), .B(n9729), .ZN(n9782)
         );
  MUX2_X1 U10918 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9782), .S(n10082), .Z(
        P1_U3536) );
  MUX2_X1 U10919 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9732), .S(n10082), .Z(
        P1_U3522) );
  INV_X1 U10920 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9734) );
  MUX2_X1 U10921 ( .A(n9734), .B(n9733), .S(n10077), .Z(n9735) );
  OAI21_X1 U10922 ( .B1(n4472), .B2(n9780), .A(n9735), .ZN(P1_U3520) );
  MUX2_X1 U10923 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9736), .S(n10077), .Z(
        P1_U3519) );
  MUX2_X1 U10924 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9737), .S(n10077), .Z(
        P1_U3518) );
  INV_X1 U10925 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n9739) );
  MUX2_X1 U10926 ( .A(n9739), .B(n9738), .S(n10077), .Z(n9740) );
  OAI21_X1 U10927 ( .B1(n9741), .B2(n9780), .A(n9740), .ZN(P1_U3517) );
  INV_X1 U10928 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9743) );
  MUX2_X1 U10929 ( .A(n9743), .B(n9742), .S(n10077), .Z(n9744) );
  OAI21_X1 U10930 ( .B1(n9745), .B2(n9780), .A(n9744), .ZN(P1_U3516) );
  INV_X1 U10931 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9747) );
  MUX2_X1 U10932 ( .A(n9747), .B(n9746), .S(n10077), .Z(n9748) );
  OAI21_X1 U10933 ( .B1(n9749), .B2(n9780), .A(n9748), .ZN(P1_U3515) );
  INV_X1 U10934 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9751) );
  MUX2_X1 U10935 ( .A(n9751), .B(n9750), .S(n10077), .Z(n9752) );
  OAI21_X1 U10936 ( .B1(n9753), .B2(n9780), .A(n9752), .ZN(P1_U3514) );
  INV_X1 U10937 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9755) );
  MUX2_X1 U10938 ( .A(n9755), .B(n9754), .S(n10077), .Z(n9756) );
  OAI21_X1 U10939 ( .B1(n9757), .B2(n9780), .A(n9756), .ZN(P1_U3513) );
  MUX2_X1 U10940 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9758), .S(n10077), .Z(
        P1_U3512) );
  MUX2_X1 U10941 ( .A(n9760), .B(n9759), .S(n10077), .Z(n9761) );
  OAI21_X1 U10942 ( .B1(n9762), .B2(n9780), .A(n9761), .ZN(P1_U3511) );
  MUX2_X1 U10943 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9763), .S(n10077), .Z(
        P1_U3510) );
  INV_X1 U10944 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n9765) );
  MUX2_X1 U10945 ( .A(n9765), .B(n9764), .S(n10077), .Z(n9766) );
  OAI21_X1 U10946 ( .B1(n9767), .B2(n9780), .A(n9766), .ZN(P1_U3509) );
  MUX2_X1 U10947 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9768), .S(n10077), .Z(
        P1_U3507) );
  MUX2_X1 U10948 ( .A(n9770), .B(n9769), .S(n10077), .Z(n9771) );
  OAI21_X1 U10949 ( .B1(n9772), .B2(n9780), .A(n9771), .ZN(P1_U3504) );
  INV_X1 U10950 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9774) );
  MUX2_X1 U10951 ( .A(n9774), .B(n9773), .S(n10077), .Z(n9775) );
  OAI21_X1 U10952 ( .B1(n9776), .B2(n9780), .A(n9775), .ZN(P1_U3501) );
  INV_X1 U10953 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9778) );
  MUX2_X1 U10954 ( .A(n9778), .B(n9777), .S(n10077), .Z(n9779) );
  OAI21_X1 U10955 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(P1_U3498) );
  MUX2_X1 U10956 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9782), .S(n10077), .Z(
        P1_U3495) );
  NOR2_X1 U10957 ( .A1(n9784), .A2(n9783), .ZN(n10047) );
  MUX2_X1 U10958 ( .A(P1_D_REG_1__SCAN_IN), .B(n9785), .S(n10047), .Z(P1_U3440) );
  MUX2_X1 U10959 ( .A(P1_D_REG_0__SCAN_IN), .B(n9786), .S(n10047), .Z(P1_U3439) );
  NOR4_X1 U10960 ( .A1(n9787), .A2(P1_IR_REG_30__SCAN_IN), .A3(P1_U3086), .A4(
        n9788), .ZN(n9789) );
  AOI21_X1 U10961 ( .B1(n9790), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9789), .ZN(
        n9791) );
  OAI21_X1 U10962 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(P1_U3324) );
  MUX2_X1 U10963 ( .A(n9794), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U10964 ( .A1(n9796), .A2(n9795), .ZN(n9844) );
  NOR2_X1 U10965 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9840) );
  NOR2_X1 U10966 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9837) );
  NOR2_X1 U10967 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9834) );
  NOR2_X1 U10968 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9831) );
  NOR2_X1 U10969 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9829) );
  NOR2_X1 U10970 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9827) );
  INV_X1 U10971 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9918) );
  AOI22_X1 U10972 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(n9918), .B1(
        P1_ADDR_REG_12__SCAN_IN), .B2(n9797), .ZN(n10264) );
  NAND2_X1 U10973 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9825) );
  INV_X1 U10974 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9902) );
  XNOR2_X1 U10975 ( .A(n9902), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(n10266) );
  NOR2_X1 U10976 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n10267) );
  NOR2_X1 U10977 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9805) );
  XNOR2_X1 U10978 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10285) );
  NAND2_X1 U10979 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9803) );
  XNOR2_X1 U10980 ( .A(n9798), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U10981 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n9801) );
  AOI21_X1 U10982 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10245) );
  NOR2_X1 U10983 ( .A1(n10249), .A2(n10248), .ZN(n10247) );
  NOR2_X1 U10984 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n10244), .ZN(n9799) );
  NOR2_X1 U10985 ( .A1(n10245), .A2(n9799), .ZN(n10281) );
  XOR2_X1 U10986 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10280) );
  NAND2_X1 U10987 ( .A1(n10281), .A2(n10280), .ZN(n9800) );
  NAND2_X1 U10988 ( .A1(n9801), .A2(n9800), .ZN(n10282) );
  NAND2_X1 U10989 ( .A1(n10283), .A2(n10282), .ZN(n9802) );
  NAND2_X1 U10990 ( .A1(n9803), .A2(n9802), .ZN(n10284) );
  NOR2_X1 U10991 ( .A1(n10285), .A2(n10284), .ZN(n9804) );
  NOR2_X1 U10992 ( .A1(n9805), .A2(n9804), .ZN(n9806) );
  NOR2_X1 U10993 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9806), .ZN(n10273) );
  AND2_X1 U10994 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n9806), .ZN(n10272) );
  NOR2_X1 U10995 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10272), .ZN(n9807) );
  NOR2_X1 U10996 ( .A1(n10273), .A2(n9807), .ZN(n9809) );
  NAND2_X1 U10997 ( .A1(n9809), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9811) );
  XNOR2_X1 U10998 ( .A(n9809), .B(n9808), .ZN(n10271) );
  NAND2_X1 U10999 ( .A1(n10271), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9810) );
  NAND2_X1 U11000 ( .A1(n9811), .A2(n9810), .ZN(n9812) );
  NAND2_X1 U11001 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9812), .ZN(n9815) );
  XNOR2_X1 U11002 ( .A(n9813), .B(n9812), .ZN(n10278) );
  NAND2_X1 U11003 ( .A1(n10278), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9814) );
  NAND2_X1 U11004 ( .A1(n9815), .A2(n9814), .ZN(n9816) );
  NAND2_X1 U11005 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9816), .ZN(n9819) );
  XNOR2_X1 U11006 ( .A(n9817), .B(n9816), .ZN(n10279) );
  NAND2_X1 U11007 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10279), .ZN(n9818) );
  NAND2_X1 U11008 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  AND2_X1 U11009 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n9820), .ZN(n9821) );
  INV_X1 U11010 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n10277) );
  XNOR2_X1 U11011 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n9820), .ZN(n10276) );
  NOR2_X1 U11012 ( .A1(n10277), .A2(n10276), .ZN(n10275) );
  NOR2_X1 U11013 ( .A1(n9821), .A2(n10275), .ZN(n10270) );
  INV_X1 U11014 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9855) );
  NOR2_X1 U11015 ( .A1(n9855), .A2(n9822), .ZN(n10268) );
  INV_X1 U11016 ( .A(n10268), .ZN(n9823) );
  OAI21_X1 U11017 ( .B1(n10267), .B2(n10270), .A(n9823), .ZN(n10265) );
  NAND2_X1 U11018 ( .A1(n10266), .A2(n10265), .ZN(n9824) );
  NAND2_X1 U11019 ( .A1(n9825), .A2(n9824), .ZN(n10263) );
  NOR2_X1 U11020 ( .A1(n10264), .A2(n10263), .ZN(n9826) );
  NOR2_X1 U11021 ( .A1(n9827), .A2(n9826), .ZN(n10262) );
  INV_X1 U11022 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9936) );
  XOR2_X1 U11023 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n9936), .Z(n10261) );
  NOR2_X1 U11024 ( .A1(n10262), .A2(n10261), .ZN(n9828) );
  NOR2_X1 U11025 ( .A1(n9829), .A2(n9828), .ZN(n10260) );
  INV_X1 U11026 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9952) );
  XOR2_X1 U11027 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(n9952), .Z(n10259) );
  NOR2_X1 U11028 ( .A1(n10260), .A2(n10259), .ZN(n9830) );
  NOR2_X1 U11029 ( .A1(n9831), .A2(n9830), .ZN(n10258) );
  INV_X1 U11030 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9963) );
  AOI22_X1 U11031 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(n9963), .B1(
        P1_ADDR_REG_15__SCAN_IN), .B2(n9832), .ZN(n10257) );
  NOR2_X1 U11032 ( .A1(n10258), .A2(n10257), .ZN(n9833) );
  NOR2_X1 U11033 ( .A1(n9834), .A2(n9833), .ZN(n10256) );
  INV_X1 U11034 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9978) );
  AOI22_X1 U11035 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(n9978), .B1(
        P1_ADDR_REG_16__SCAN_IN), .B2(n9835), .ZN(n10255) );
  NOR2_X1 U11036 ( .A1(n10256), .A2(n10255), .ZN(n9836) );
  NOR2_X1 U11037 ( .A1(n9837), .A2(n9836), .ZN(n10254) );
  INV_X1 U11038 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n9991) );
  INV_X1 U11039 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9838) );
  AOI22_X1 U11040 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n9991), .B1(
        P1_ADDR_REG_17__SCAN_IN), .B2(n9838), .ZN(n10253) );
  NOR2_X1 U11041 ( .A1(n10254), .A2(n10253), .ZN(n9839) );
  NOR2_X1 U11042 ( .A1(n9840), .A2(n9839), .ZN(n9841) );
  NOR2_X1 U11043 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9841), .ZN(n10250) );
  AND2_X1 U11044 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n9841), .ZN(n10251) );
  NOR2_X1 U11045 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10251), .ZN(n9842) );
  NOR2_X1 U11046 ( .A1(n10250), .A2(n9842), .ZN(n9843) );
  XOR2_X1 U11047 ( .A(n9844), .B(n9843), .Z(ADD_1068_U4) );
  AOI211_X1 U11048 ( .C1(n9847), .C2(n9846), .A(n9993), .B(n9845), .ZN(n9852)
         );
  AOI211_X1 U11049 ( .C1(n9850), .C2(n9849), .A(n9999), .B(n9848), .ZN(n9851)
         );
  AOI211_X1 U11050 ( .C1(n10005), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9854)
         );
  NAND2_X1 U11051 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n9863) );
  OAI211_X1 U11052 ( .C1(n9855), .C2(n10008), .A(n9854), .B(n9863), .ZN(
        P1_U3253) );
  XNOR2_X1 U11053 ( .A(n9856), .B(n9857), .ZN(n9858) );
  NAND2_X1 U11054 ( .A1(n9858), .A2(n9859), .ZN(n9878) );
  OAI21_X1 U11055 ( .B1(n9859), .B2(n9858), .A(n9878), .ZN(n9860) );
  AOI222_X1 U11056 ( .A1(n9887), .A2(n9862), .B1(n9861), .B2(n9882), .C1(n9860), .C2(n9885), .ZN(n9864) );
  OAI211_X1 U11057 ( .C1(n9890), .C2(n9865), .A(n9864), .B(n9863), .ZN(
        P1_U3217) );
  INV_X1 U11058 ( .A(n9866), .ZN(n9871) );
  OAI21_X1 U11059 ( .B1(n9869), .B2(n9868), .A(n9867), .ZN(n9870) );
  AOI222_X1 U11060 ( .A1(n9887), .A2(n9872), .B1(n9871), .B2(n9882), .C1(n9870), .C2(n9885), .ZN(n9873) );
  NAND2_X1 U11061 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n9916) );
  OAI211_X1 U11062 ( .C1(n9890), .C2(n9874), .A(n9873), .B(n9916), .ZN(
        P1_U3224) );
  OAI21_X1 U11063 ( .B1(n9877), .B2(n9876), .A(n9875), .ZN(n9881) );
  OAI21_X1 U11064 ( .B1(n9879), .B2(n9856), .A(n9878), .ZN(n9880) );
  XOR2_X1 U11065 ( .A(n9881), .B(n9880), .Z(n9884) );
  AOI222_X1 U11066 ( .A1(n9887), .A2(n4595), .B1(n9885), .B2(n9884), .C1(n9883), .C2(n9882), .ZN(n9888) );
  NAND2_X1 U11067 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n9900) );
  OAI211_X1 U11068 ( .C1(n9890), .C2(n9889), .A(n9888), .B(n9900), .ZN(
        P1_U3236) );
  XNOR2_X1 U11069 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  AOI211_X1 U11070 ( .C1(n9893), .C2(n9892), .A(n9891), .B(n9999), .ZN(n9898)
         );
  AOI211_X1 U11071 ( .C1(n9896), .C2(n9895), .A(n9894), .B(n9993), .ZN(n9897)
         );
  AOI211_X1 U11072 ( .C1(n10005), .C2(n9899), .A(n9898), .B(n9897), .ZN(n9901)
         );
  OAI211_X1 U11073 ( .C1(n9902), .C2(n10008), .A(n9901), .B(n9900), .ZN(
        P1_U3254) );
  INV_X1 U11074 ( .A(n9903), .ZN(n9914) );
  OAI21_X1 U11075 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9907) );
  NAND2_X1 U11076 ( .A1(n9986), .A2(n9907), .ZN(n9913) );
  OAI21_X1 U11077 ( .B1(n9910), .B2(n9909), .A(n9908), .ZN(n9911) );
  NAND2_X1 U11078 ( .A1(n9987), .A2(n9911), .ZN(n9912) );
  OAI211_X1 U11079 ( .C1(n9974), .C2(n9914), .A(n9913), .B(n9912), .ZN(n9915)
         );
  INV_X1 U11080 ( .A(n9915), .ZN(n9917) );
  OAI211_X1 U11081 ( .C1(n9918), .C2(n10008), .A(n9917), .B(n9916), .ZN(
        P1_U3255) );
  INV_X1 U11082 ( .A(n9919), .ZN(n9932) );
  INV_X1 U11083 ( .A(n9920), .ZN(n9922) );
  NAND2_X1 U11084 ( .A1(n9922), .A2(n9921), .ZN(n9923) );
  NAND2_X1 U11085 ( .A1(n9924), .A2(n9923), .ZN(n9925) );
  OR2_X1 U11086 ( .A1(n9999), .A2(n9925), .ZN(n9931) );
  OAI21_X1 U11087 ( .B1(n9928), .B2(n9927), .A(n9926), .ZN(n9929) );
  OR2_X1 U11088 ( .A1(n9993), .A2(n9929), .ZN(n9930) );
  OAI211_X1 U11089 ( .C1(n9974), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9933)
         );
  INV_X1 U11090 ( .A(n9933), .ZN(n9935) );
  OAI211_X1 U11091 ( .C1(n9936), .C2(n10008), .A(n9935), .B(n9934), .ZN(
        P1_U3256) );
  AOI21_X1 U11092 ( .B1(n9939), .B2(n9938), .A(n9937), .ZN(n9940) );
  NAND2_X1 U11093 ( .A1(n9987), .A2(n9940), .ZN(n9947) );
  INV_X1 U11094 ( .A(n9941), .ZN(n9942) );
  OAI21_X1 U11095 ( .B1(n9944), .B2(n9943), .A(n9942), .ZN(n9945) );
  OR2_X1 U11096 ( .A1(n9993), .A2(n9945), .ZN(n9946) );
  OAI211_X1 U11097 ( .C1(n9974), .C2(n9948), .A(n9947), .B(n9946), .ZN(n9949)
         );
  INV_X1 U11098 ( .A(n9949), .ZN(n9951) );
  NAND2_X1 U11099 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n9950) );
  OAI211_X1 U11100 ( .C1(n9952), .C2(n10008), .A(n9951), .B(n9950), .ZN(
        P1_U3257) );
  AOI211_X1 U11101 ( .C1(n9955), .C2(n9954), .A(n9953), .B(n9993), .ZN(n9959)
         );
  AOI211_X1 U11102 ( .C1(n9957), .C2(n8199), .A(n9956), .B(n9999), .ZN(n9958)
         );
  AOI211_X1 U11103 ( .C1(n10005), .C2(n9960), .A(n9959), .B(n9958), .ZN(n9962)
         );
  OAI211_X1 U11104 ( .C1(n9963), .C2(n10008), .A(n9962), .B(n9961), .ZN(
        P1_U3258) );
  XNOR2_X1 U11105 ( .A(n9965), .B(n9964), .ZN(n9966) );
  NAND2_X1 U11106 ( .A1(n9966), .A2(n9986), .ZN(n9972) );
  NAND2_X1 U11107 ( .A1(n9968), .A2(n9967), .ZN(n9969) );
  NAND3_X1 U11108 ( .A1(n9970), .A2(n9987), .A3(n9969), .ZN(n9971) );
  OAI211_X1 U11109 ( .C1(n9974), .C2(n9973), .A(n9972), .B(n9971), .ZN(n9975)
         );
  INV_X1 U11110 ( .A(n9975), .ZN(n9977) );
  OAI211_X1 U11111 ( .C1(n9978), .C2(n10008), .A(n9977), .B(n9976), .ZN(
        P1_U3259) );
  OAI21_X1 U11112 ( .B1(n9981), .B2(n9980), .A(n9979), .ZN(n9988) );
  XNOR2_X1 U11113 ( .A(n9983), .B(n9982), .ZN(n9985) );
  AOI222_X1 U11114 ( .A1(n9988), .A2(n9987), .B1(n9986), .B2(n9985), .C1(n9984), .C2(n10005), .ZN(n9990) );
  OAI211_X1 U11115 ( .C1(n9991), .C2(n10008), .A(n9990), .B(n9989), .ZN(
        P1_U3260) );
  AOI211_X1 U11116 ( .C1(n9995), .C2(n9994), .A(n9993), .B(n9992), .ZN(n10003)
         );
  INV_X1 U11117 ( .A(n9996), .ZN(n10000) );
  INV_X1 U11118 ( .A(n9997), .ZN(n9998) );
  AOI211_X1 U11119 ( .C1(n10001), .C2(n10000), .A(n9999), .B(n9998), .ZN(
        n10002) );
  AOI211_X1 U11120 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n10007) );
  OAI211_X1 U11121 ( .C1(n10009), .C2(n10008), .A(n10007), .B(n10006), .ZN(
        P1_U3261) );
  INV_X1 U11122 ( .A(n10010), .ZN(n10011) );
  AOI222_X1 U11123 ( .A1(n10012), .A2(n10035), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n10045), .C1(n10011), .C2(n10032), .ZN(n10018) );
  INV_X1 U11124 ( .A(n10013), .ZN(n10014) );
  AOI22_X1 U11125 ( .A1(n10016), .A2(n10041), .B1(n10015), .B2(n10014), .ZN(
        n10017) );
  OAI211_X1 U11126 ( .C1(n10045), .C2(n10019), .A(n10018), .B(n10017), .ZN(
        P1_U3285) );
  OAI22_X1 U11127 ( .A1(n10023), .A2(n10022), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n10021), .ZN(n10024) );
  AOI21_X1 U11128 ( .B1(n10035), .B2(n10025), .A(n10024), .ZN(n10026) );
  OAI21_X1 U11129 ( .B1(n10038), .B2(n10027), .A(n10026), .ZN(n10028) );
  AOI21_X1 U11130 ( .B1(n10029), .B2(n4616), .A(n10028), .ZN(n10030) );
  OAI21_X1 U11131 ( .B1(n10045), .B2(n10031), .A(n10030), .ZN(P1_U3290) );
  AOI22_X1 U11132 ( .A1(n10033), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n10032), .ZN(n10037) );
  NAND2_X1 U11133 ( .A1(n10035), .A2(n10034), .ZN(n10036) );
  OAI211_X1 U11134 ( .C1(n10039), .C2(n10038), .A(n10037), .B(n10036), .ZN(
        n10040) );
  AOI21_X1 U11135 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  OAI21_X1 U11136 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(P1_U3292) );
  AND2_X1 U11137 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10048), .ZN(P1_U3294) );
  AND2_X1 U11138 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10048), .ZN(P1_U3295) );
  AND2_X1 U11139 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10048), .ZN(P1_U3296) );
  NOR2_X1 U11140 ( .A1(n10047), .A2(n10046), .ZN(P1_U3297) );
  AND2_X1 U11141 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10048), .ZN(P1_U3298) );
  AND2_X1 U11142 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10048), .ZN(P1_U3299) );
  AND2_X1 U11143 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10048), .ZN(P1_U3300) );
  AND2_X1 U11144 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10048), .ZN(P1_U3301) );
  AND2_X1 U11145 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10048), .ZN(P1_U3302) );
  AND2_X1 U11146 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10048), .ZN(P1_U3303) );
  AND2_X1 U11147 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10048), .ZN(P1_U3304) );
  AND2_X1 U11148 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10048), .ZN(P1_U3305) );
  AND2_X1 U11149 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10048), .ZN(P1_U3306) );
  AND2_X1 U11150 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10048), .ZN(P1_U3307) );
  AND2_X1 U11151 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10048), .ZN(P1_U3308) );
  AND2_X1 U11152 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10048), .ZN(P1_U3309) );
  AND2_X1 U11153 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10048), .ZN(P1_U3310) );
  AND2_X1 U11154 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10048), .ZN(P1_U3311) );
  AND2_X1 U11155 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10048), .ZN(P1_U3312) );
  AND2_X1 U11156 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10048), .ZN(P1_U3313) );
  AND2_X1 U11157 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10048), .ZN(P1_U3314) );
  AND2_X1 U11158 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10048), .ZN(P1_U3315) );
  AND2_X1 U11159 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10048), .ZN(P1_U3316) );
  AND2_X1 U11160 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10048), .ZN(P1_U3317) );
  AND2_X1 U11161 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10048), .ZN(P1_U3318) );
  AND2_X1 U11162 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10048), .ZN(P1_U3319) );
  AND2_X1 U11163 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10048), .ZN(P1_U3320) );
  AND2_X1 U11164 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10048), .ZN(P1_U3321) );
  AND2_X1 U11165 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10048), .ZN(P1_U3322) );
  AND2_X1 U11166 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10048), .ZN(P1_U3323) );
  INV_X1 U11167 ( .A(n10069), .ZN(n10054) );
  INV_X1 U11168 ( .A(n10057), .ZN(n10067) );
  OAI21_X1 U11169 ( .B1(n10050), .B2(n10067), .A(n10049), .ZN(n10052) );
  AOI211_X1 U11170 ( .C1(n10054), .C2(n10053), .A(n10052), .B(n10051), .ZN(
        n10078) );
  INV_X1 U11171 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10055) );
  AOI22_X1 U11172 ( .A1(n10077), .A2(n10078), .B1(n10055), .B2(n10075), .ZN(
        P1_U3459) );
  AOI22_X1 U11173 ( .A1(n10059), .A2(n10058), .B1(n10057), .B2(n10056), .ZN(
        n10060) );
  OAI211_X1 U11174 ( .C1(n10063), .C2(n10062), .A(n10061), .B(n10060), .ZN(
        n10064) );
  INV_X1 U11175 ( .A(n10064), .ZN(n10079) );
  AOI22_X1 U11176 ( .A1(n10077), .A2(n10079), .B1(n5709), .B2(n10075), .ZN(
        P1_U3471) );
  INV_X1 U11177 ( .A(n10070), .ZN(n10073) );
  OAI211_X1 U11178 ( .C1(n10068), .C2(n10067), .A(n10066), .B(n10065), .ZN(
        n10072) );
  NOR2_X1 U11179 ( .A1(n10070), .A2(n10069), .ZN(n10071) );
  AOI211_X1 U11180 ( .C1(n10074), .C2(n10073), .A(n10072), .B(n10071), .ZN(
        n10081) );
  INV_X1 U11181 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U11182 ( .A1(n10077), .A2(n10081), .B1(n10076), .B2(n10075), .ZN(
        P1_U3486) );
  AOI22_X1 U11183 ( .A1(n10082), .A2(n10078), .B1(n5677), .B2(n10080), .ZN(
        P1_U3524) );
  AOI22_X1 U11184 ( .A1(n10082), .A2(n10079), .B1(n6912), .B2(n10080), .ZN(
        P1_U3528) );
  AOI22_X1 U11185 ( .A1(n10082), .A2(n10081), .B1(n9402), .B2(n10080), .ZN(
        P1_U3533) );
  AOI22_X1 U11186 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n10109), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3151), .ZN(n10088) );
  INV_X1 U11187 ( .A(n10083), .ZN(n10086) );
  XNOR2_X1 U11188 ( .A(n10084), .B(n10089), .ZN(n10085) );
  OAI21_X1 U11189 ( .B1(n5610), .B2(n10086), .A(n10085), .ZN(n10087) );
  OAI211_X1 U11190 ( .C1(n10128), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        P2_U3182) );
  AOI22_X1 U11191 ( .A1(n10091), .A2(n10090), .B1(n10109), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10108) );
  AOI21_X1 U11192 ( .B1(n10094), .B2(n10093), .A(n10092), .ZN(n10105) );
  OAI21_X1 U11193 ( .B1(n10097), .B2(n10096), .A(n10095), .ZN(n10098) );
  NAND2_X1 U11194 ( .A1(n5610), .A2(n10098), .ZN(n10104) );
  AOI21_X1 U11195 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10102) );
  OR2_X1 U11196 ( .A1(n10102), .A2(n10118), .ZN(n10103) );
  OAI211_X1 U11197 ( .C1(n10105), .C2(n10122), .A(n10104), .B(n10103), .ZN(
        n10106) );
  INV_X1 U11198 ( .A(n10106), .ZN(n10107) );
  OAI211_X1 U11199 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n6255), .A(n10108), .B(
        n10107), .ZN(P2_U3195) );
  AOI22_X1 U11200 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(n10109), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3151), .ZN(n10126) );
  AOI21_X1 U11201 ( .B1(n4407), .B2(n10111), .A(n10110), .ZN(n10123) );
  OAI21_X1 U11202 ( .B1(n10114), .B2(n10113), .A(n10112), .ZN(n10115) );
  NAND2_X1 U11203 ( .A1(n5610), .A2(n10115), .ZN(n10121) );
  AOI21_X1 U11204 ( .B1(n10117), .B2(n10116), .A(n4364), .ZN(n10119) );
  OR2_X1 U11205 ( .A1(n10119), .A2(n10118), .ZN(n10120) );
  OAI211_X1 U11206 ( .C1(n10123), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        n10124) );
  INV_X1 U11207 ( .A(n10124), .ZN(n10125) );
  OAI211_X1 U11208 ( .C1(n10128), .C2(n10127), .A(n10126), .B(n10125), .ZN(
        P2_U3196) );
  XOR2_X1 U11209 ( .A(n10137), .B(n10129), .Z(n10134) );
  AOI222_X1 U11210 ( .A1(n10135), .A2(n10134), .B1(n10133), .B2(n10132), .C1(
        n10131), .C2(n10130), .ZN(n10170) );
  XNOR2_X1 U11211 ( .A(n10136), .B(n10137), .ZN(n10172) );
  AOI222_X1 U11212 ( .A1(n10172), .A2(n10142), .B1(n10141), .B2(n10140), .C1(
        n10139), .C2(n10138), .ZN(n10143) );
  OAI221_X1 U11213 ( .B1(n10162), .B2(n10170), .C1(n10160), .C2(n6132), .A(
        n10143), .ZN(P2_U3230) );
  XNOR2_X1 U11214 ( .A(n10144), .B(n10150), .ZN(n10169) );
  AND2_X1 U11215 ( .A1(n10145), .A2(n10221), .ZN(n10168) );
  INV_X1 U11216 ( .A(n10168), .ZN(n10146) );
  OAI22_X1 U11217 ( .A1(n10149), .A2(n10148), .B1(n10147), .B2(n10146), .ZN(
        n10158) );
  XNOR2_X1 U11218 ( .A(n10151), .B(n10150), .ZN(n10152) );
  OAI222_X1 U11219 ( .A1(n10157), .A2(n10156), .B1(n10155), .B2(n10154), .C1(
        n10153), .C2(n10152), .ZN(n10167) );
  AOI211_X1 U11220 ( .C1(n10169), .C2(n10159), .A(n10158), .B(n10167), .ZN(
        n10161) );
  AOI22_X1 U11221 ( .A1(n10162), .A2(n4536), .B1(n10161), .B2(n10160), .ZN(
        P2_U3231) );
  INV_X1 U11222 ( .A(n10163), .ZN(n10166) );
  OAI22_X1 U11223 ( .A1(n10164), .A2(n10215), .B1(n10210), .B2(n6106), .ZN(
        n10165) );
  NOR2_X1 U11224 ( .A1(n10166), .A2(n10165), .ZN(n10226) );
  AOI22_X1 U11225 ( .A1(n10224), .A2(n6095), .B1(n10226), .B2(n10222), .ZN(
        P2_U3393) );
  AOI211_X1 U11226 ( .C1(n10169), .C2(n10196), .A(n10168), .B(n10167), .ZN(
        n10228) );
  AOI22_X1 U11227 ( .A1(n10224), .A2(n6124), .B1(n10228), .B2(n10222), .ZN(
        P2_U3396) );
  OAI21_X1 U11228 ( .B1(n4525), .B2(n10210), .A(n10170), .ZN(n10171) );
  AOI21_X1 U11229 ( .B1(n10196), .B2(n10172), .A(n10171), .ZN(n10230) );
  AOI22_X1 U11230 ( .A1(n10224), .A2(n6134), .B1(n10230), .B2(n10222), .ZN(
        P2_U3399) );
  INV_X1 U11231 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10178) );
  NOR2_X1 U11232 ( .A1(n10173), .A2(n10215), .ZN(n10176) );
  INV_X1 U11233 ( .A(n10174), .ZN(n10175) );
  AOI211_X1 U11234 ( .C1(n10221), .C2(n10177), .A(n10176), .B(n10175), .ZN(
        n10231) );
  AOI22_X1 U11235 ( .A1(n10224), .A2(n10178), .B1(n10231), .B2(n10222), .ZN(
        P2_U3402) );
  INV_X1 U11236 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10183) );
  INV_X1 U11237 ( .A(n10207), .ZN(n10199) );
  OAI22_X1 U11238 ( .A1(n10180), .A2(n10199), .B1(n10179), .B2(n10210), .ZN(
        n10181) );
  NOR2_X1 U11239 ( .A1(n10182), .A2(n10181), .ZN(n10232) );
  AOI22_X1 U11240 ( .A1(n10224), .A2(n10183), .B1(n10232), .B2(n10222), .ZN(
        P2_U3405) );
  NOR2_X1 U11241 ( .A1(n10184), .A2(n10210), .ZN(n10186) );
  AOI211_X1 U11242 ( .C1(n10187), .C2(n10196), .A(n10186), .B(n10185), .ZN(
        n10233) );
  AOI22_X1 U11243 ( .A1(n10224), .A2(n6168), .B1(n10233), .B2(n10222), .ZN(
        P2_U3408) );
  OAI22_X1 U11244 ( .A1(n10189), .A2(n10199), .B1(n10188), .B2(n10210), .ZN(
        n10190) );
  NOR2_X1 U11245 ( .A1(n10191), .A2(n10190), .ZN(n10235) );
  AOI22_X1 U11246 ( .A1(n10224), .A2(n6181), .B1(n10235), .B2(n10222), .ZN(
        P2_U3411) );
  INV_X1 U11247 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10197) );
  OAI21_X1 U11248 ( .B1(n10193), .B2(n10210), .A(n10192), .ZN(n10194) );
  AOI21_X1 U11249 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(n10236) );
  AOI22_X1 U11250 ( .A1(n10224), .A2(n10197), .B1(n10236), .B2(n10222), .ZN(
        P2_U3414) );
  INV_X1 U11251 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10203) );
  OAI22_X1 U11252 ( .A1(n10200), .A2(n10199), .B1(n10198), .B2(n10210), .ZN(
        n10201) );
  NOR2_X1 U11253 ( .A1(n10202), .A2(n10201), .ZN(n10238) );
  AOI22_X1 U11254 ( .A1(n10224), .A2(n10203), .B1(n10238), .B2(n10222), .ZN(
        P2_U3417) );
  INV_X1 U11255 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10209) );
  NOR2_X1 U11256 ( .A1(n10204), .A2(n10210), .ZN(n10206) );
  AOI211_X1 U11257 ( .C1(n10208), .C2(n10207), .A(n10206), .B(n10205), .ZN(
        n10239) );
  AOI22_X1 U11258 ( .A1(n10224), .A2(n10209), .B1(n10239), .B2(n10222), .ZN(
        P2_U3420) );
  OAI22_X1 U11259 ( .A1(n10212), .A2(n10215), .B1(n10211), .B2(n10210), .ZN(
        n10213) );
  NOR2_X1 U11260 ( .A1(n10214), .A2(n10213), .ZN(n10241) );
  AOI22_X1 U11261 ( .A1(n10224), .A2(n6231), .B1(n10241), .B2(n10222), .ZN(
        P2_U3423) );
  INV_X1 U11262 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10223) );
  NOR3_X1 U11263 ( .A1(n10217), .A2(n10216), .A3(n10215), .ZN(n10219) );
  AOI211_X1 U11264 ( .C1(n10221), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10242) );
  AOI22_X1 U11265 ( .A1(n10224), .A2(n10223), .B1(n10242), .B2(n10222), .ZN(
        P2_U3426) );
  AOI22_X1 U11266 ( .A1(n10243), .A2(n10226), .B1(n10225), .B2(n6505), .ZN(
        P2_U3460) );
  INV_X1 U11267 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U11268 ( .A1(n10243), .A2(n10228), .B1(n10227), .B2(n6505), .ZN(
        P2_U3461) );
  INV_X1 U11269 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U11270 ( .A1(n10243), .A2(n10230), .B1(n10229), .B2(n6505), .ZN(
        P2_U3462) );
  AOI22_X1 U11271 ( .A1(n10243), .A2(n10231), .B1(n6146), .B2(n6505), .ZN(
        P2_U3463) );
  AOI22_X1 U11272 ( .A1(n10243), .A2(n10232), .B1(n6156), .B2(n6505), .ZN(
        P2_U3464) );
  AOI22_X1 U11273 ( .A1(n10243), .A2(n10233), .B1(n5541), .B2(n6505), .ZN(
        P2_U3465) );
  AOI22_X1 U11274 ( .A1(n10243), .A2(n10235), .B1(n10234), .B2(n6505), .ZN(
        P2_U3466) );
  AOI22_X1 U11275 ( .A1(n10243), .A2(n10236), .B1(n6197), .B2(n6505), .ZN(
        P2_U3467) );
  AOI22_X1 U11276 ( .A1(n10243), .A2(n10238), .B1(n10237), .B2(n6505), .ZN(
        P2_U3468) );
  AOI22_X1 U11277 ( .A1(n10243), .A2(n10239), .B1(n6219), .B2(n6505), .ZN(
        P2_U3469) );
  AOI22_X1 U11278 ( .A1(n10243), .A2(n10241), .B1(n10240), .B2(n6505), .ZN(
        P2_U3470) );
  AOI22_X1 U11279 ( .A1(n10243), .A2(n10242), .B1(n6242), .B2(n6505), .ZN(
        P2_U3471) );
  NOR2_X1 U11280 ( .A1(n10245), .A2(n10244), .ZN(n10246) );
  XOR2_X1 U11281 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10246), .Z(ADD_1068_U5) );
  AOI21_X1 U11282 ( .B1(n10249), .B2(n10248), .A(n10247), .ZN(ADD_1068_U46) );
  NOR2_X1 U11283 ( .A1(n10251), .A2(n10250), .ZN(n10252) );
  XOR2_X1 U11284 ( .A(n10252), .B(P2_ADDR_REG_18__SCAN_IN), .Z(ADD_1068_U55)
         );
  XNOR2_X1 U11285 ( .A(n10254), .B(n10253), .ZN(ADD_1068_U56) );
  XNOR2_X1 U11286 ( .A(n10256), .B(n10255), .ZN(ADD_1068_U57) );
  XNOR2_X1 U11287 ( .A(n10258), .B(n10257), .ZN(ADD_1068_U58) );
  XNOR2_X1 U11288 ( .A(n10260), .B(n10259), .ZN(ADD_1068_U59) );
  XNOR2_X1 U11289 ( .A(n10262), .B(n10261), .ZN(ADD_1068_U60) );
  XNOR2_X1 U11290 ( .A(n10264), .B(n10263), .ZN(ADD_1068_U61) );
  XOR2_X1 U11291 ( .A(n10266), .B(n10265), .Z(ADD_1068_U62) );
  NOR2_X1 U11292 ( .A1(n10268), .A2(n10267), .ZN(n10269) );
  XNOR2_X1 U11293 ( .A(n10270), .B(n10269), .ZN(ADD_1068_U63) );
  XOR2_X1 U11294 ( .A(n10271), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1068_U50) );
  NOR2_X1 U11295 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  XOR2_X1 U11296 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10274), .Z(ADD_1068_U51) );
  AOI21_X1 U11297 ( .B1(n10277), .B2(n10276), .A(n10275), .ZN(ADD_1068_U47) );
  XOR2_X1 U11298 ( .A(n10278), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1068_U49) );
  XOR2_X1 U11299 ( .A(n10279), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1068_U48) );
  XOR2_X1 U11300 ( .A(n10281), .B(n10280), .Z(ADD_1068_U54) );
  XOR2_X1 U11301 ( .A(n10283), .B(n10282), .Z(ADD_1068_U53) );
  XNOR2_X1 U11302 ( .A(n10285), .B(n10284), .ZN(ADD_1068_U52) );
  OR2_X1 U6822 ( .A1(n5356), .A2(n9788), .ZN(n5358) );
  NAND2_X1 U4877 ( .A1(n9787), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5355) );
  NAND3_X1 U4872 ( .A1(n4790), .A2(n4787), .A3(n6969), .ZN(n6967) );
  CLKBUF_X1 U4985 ( .A(n8671), .Z(n4335) );
endmodule

