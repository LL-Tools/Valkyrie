

module b22_C_SARLock_k_64_8 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput0,
         keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, keyinput6,
         keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, keyinput12,
         keyinput13, keyinput14, keyinput15, keyinput16, keyinput17,
         keyinput18, keyinput19, keyinput20, keyinput21, keyinput22,
         keyinput23, keyinput24, keyinput25, keyinput26, keyinput27,
         keyinput28, keyinput29, keyinput30, keyinput31, keyinput32,
         keyinput33, keyinput34, keyinput35, keyinput36, keyinput37,
         keyinput38, keyinput39, keyinput40, keyinput41, keyinput42,
         keyinput43, keyinput44, keyinput45, keyinput46, keyinput47,
         keyinput48, keyinput49, keyinput50, keyinput51, keyinput52,
         keyinput53, keyinput54, keyinput55, keyinput56, keyinput57,
         keyinput58, keyinput59, keyinput60, keyinput61, keyinput62,
         keyinput63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164;

  INV_X4 U7171 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  AOI21_X1 U7172 ( .B1(n6669), .B2(n6473), .A(n6668), .ZN(n11647) );
  INV_X1 U7173 ( .A(n12441), .ZN(n12471) );
  CLKBUF_X1 U7174 ( .A(n8269), .Z(n11653) );
  CLKBUF_X2 U7175 ( .A(n7448), .Z(n11979) );
  NAND2_X1 U7176 ( .A1(n6635), .A2(n10208), .ZN(n11686) );
  BUF_X2 U7177 ( .A(n9970), .Z(n6425) );
  INV_X1 U7178 ( .A(n14831), .ZN(n14855) );
  CLKBUF_X1 U7179 ( .A(n7503), .Z(n6464) );
  CLKBUF_X2 U7180 ( .A(n7551), .Z(n8110) );
  INV_X1 U7181 ( .A(n13436), .ZN(n13461) );
  INV_X1 U7182 ( .A(n13464), .ZN(n11515) );
  CLKBUF_X2 U7183 ( .A(n7524), .Z(n9379) );
  NOR2_X1 U7184 ( .A1(n9208), .A2(n9207), .ZN(n13767) );
  OR2_X1 U7185 ( .A1(n12402), .A2(n12403), .ZN(n12400) );
  INV_X2 U7186 ( .A(n11804), .ZN(n11808) );
  AND2_X1 U7187 ( .A1(n12400), .A2(n8702), .ZN(n12387) );
  INV_X1 U7188 ( .A(n8263), .ZN(n9975) );
  AOI21_X1 U7189 ( .B1(n11395), .B2(n8731), .A(n6498), .ZN(n8733) );
  OR2_X1 U7190 ( .A1(n7943), .A2(n9204), .ZN(n7238) );
  OR2_X2 U7191 ( .A1(n7575), .A2(n6896), .ZN(n9932) );
  INV_X1 U7192 ( .A(n6466), .ZN(n7235) );
  INV_X1 U7193 ( .A(n9363), .ZN(n9475) );
  NAND2_X1 U7194 ( .A1(n7942), .A2(n7941), .ZN(n7964) );
  INV_X1 U7195 ( .A(n8839), .ZN(n12029) );
  XNOR2_X1 U7196 ( .A(n8883), .B(n8881), .ZN(n12096) );
  AND2_X1 U7197 ( .A1(n8220), .A2(n12736), .ZN(n8269) );
  INV_X1 U7198 ( .A(n12388), .ZN(n12420) );
  INV_X1 U7200 ( .A(n9379), .ZN(n7923) );
  AND2_X1 U7201 ( .A1(n7646), .A2(n7645), .ZN(n10247) );
  INV_X1 U7202 ( .A(n13028), .ZN(n13202) );
  OAI21_X1 U7203 ( .B1(n11904), .B2(n11903), .A(n13357), .ZN(n13367) );
  NAND2_X1 U7204 ( .A1(n13535), .A2(n13536), .ZN(n9740) );
  XNOR2_X1 U7205 ( .A(n14266), .B(n14267), .ZN(n14308) );
  NAND2_X1 U7206 ( .A1(n8206), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8207) );
  NOR2_X1 U7207 ( .A1(n8758), .A2(n8757), .ZN(n8759) );
  NOR2_X1 U7208 ( .A1(n8333), .A2(n8332), .ZN(n10108) );
  CLKBUF_X3 U7210 ( .A(n7842), .Z(n14833) );
  INV_X1 U7211 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n7563) );
  INV_X1 U7212 ( .A(n9744), .ZN(n6434) );
  NAND2_X1 U7213 ( .A1(n8891), .A2(n8890), .ZN(n12115) );
  INV_X1 U7214 ( .A(n9474), .ZN(n11852) );
  XNOR2_X1 U7215 ( .A(n14311), .B(n7142), .ZN(n14373) );
  XNOR2_X1 U7216 ( .A(n8207), .B(n8215), .ZN(n8211) );
  NAND2_X1 U7217 ( .A1(n9363), .A2(n11852), .ZN(n13453) );
  AND2_X1 U7218 ( .A1(n8220), .A2(n8223), .ZN(n6422) );
  AND2_X1 U7219 ( .A1(n13970), .A2(n6448), .ZN(n6423) );
  NAND2_X1 U7220 ( .A1(n8211), .A2(n8210), .ZN(n9970) );
  OAI21_X1 U7221 ( .B1(n10022), .B2(n10023), .A(n6554), .ZN(n7033) );
  XNOR2_X1 U7222 ( .A(n9984), .B(n6695), .ZN(n10022) );
  CLKBUF_X1 U7223 ( .A(n11644), .Z(n6424) );
  NAND2_X2 U7224 ( .A1(n9205), .A2(n9184), .ZN(n9274) );
  NOR2_X4 U7225 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n9205) );
  NAND2_X2 U7226 ( .A1(n7573), .A2(n7572), .ZN(n7639) );
  NAND2_X2 U7227 ( .A1(n7568), .A2(n7567), .ZN(n7573) );
  OR2_X2 U7228 ( .A1(n12067), .A2(n12066), .ZN(n12068) );
  NOR2_X2 U7229 ( .A1(n9273), .A2(n9186), .ZN(n7365) );
  NOR2_X1 U7230 ( .A1(n10825), .A2(n14559), .ZN(n10919) );
  OR2_X1 U7231 ( .A1(n7593), .A2(n7594), .ZN(n7595) );
  XNOR2_X2 U7232 ( .A(n14323), .B(n7133), .ZN(n14380) );
  AND2_X2 U7233 ( .A1(n6851), .A2(n6571), .ZN(n14323) );
  NOR2_X2 U7234 ( .A1(n15027), .A2(n12319), .ZN(n12320) );
  OAI21_X2 U7235 ( .B1(n11245), .B2(n7431), .A(n7429), .ZN(n14073) );
  XNOR2_X2 U7236 ( .A(n13039), .B(n12980), .ZN(n13037) );
  BUF_X4 U7237 ( .A(n11608), .Z(n6426) );
  NOR2_X2 U7238 ( .A1(n8630), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8642) );
  OAI22_X2 U7239 ( .A1(n13437), .A2(n9066), .B1(n7943), .B2(n9065), .ZN(n9107)
         );
  INV_X1 U7240 ( .A(n8852), .ZN(n6427) );
  CLKBUF_X3 U7241 ( .A(n13453), .Z(n6428) );
  XOR2_X2 U7242 ( .A(n10769), .B(n10763), .Z(n10674) );
  AND2_X2 U7243 ( .A1(n10672), .A2(n10671), .ZN(n10769) );
  AOI21_X2 U7244 ( .B1(n7138), .B2(n7137), .A(n7136), .ZN(n14298) );
  INV_X1 U7245 ( .A(n6422), .ZN(n6429) );
  INV_X4 U7246 ( .A(n6422), .ZN(n6430) );
  AOI21_X1 U7247 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n9975), .A(n10042), .ZN(
        n10057) );
  XNOR2_X1 U7248 ( .A(n8297), .B(P3_IR_REG_2__SCAN_IN), .ZN(n10067) );
  NOR2_X2 U7249 ( .A1(n14600), .A2(n14599), .ZN(n14598) );
  NOR2_X2 U7250 ( .A1(n14596), .A2(n14336), .ZN(n14600) );
  NOR2_X1 U7251 ( .A1(n6453), .A2(n11589), .ZN(n14118) );
  OR2_X1 U7252 ( .A1(n13898), .A2(n13897), .ZN(n14108) );
  AND2_X1 U7253 ( .A1(n13923), .A2(n7424), .ZN(n6453) );
  OAI21_X1 U7254 ( .B1(n13980), .B2(n6907), .A(n6906), .ZN(n6910) );
  INV_X1 U7255 ( .A(n13054), .ZN(n13214) );
  INV_X1 U7256 ( .A(n12116), .ZN(n6432) );
  NAND2_X1 U7257 ( .A1(n7969), .A2(n7968), .ZN(n13230) );
  AND2_X1 U7258 ( .A1(n7024), .A2(n7018), .ZN(n15008) );
  NAND2_X1 U7259 ( .A1(n7023), .A2(n7022), .ZN(n14987) );
  NAND2_X1 U7260 ( .A1(n11066), .A2(n8847), .ZN(n11022) );
  OAI21_X1 U7261 ( .B1(n7412), .B2(n6435), .A(n11243), .ZN(n6452) );
  INV_X1 U7262 ( .A(n13484), .ZN(n6435) );
  INV_X1 U7263 ( .A(n9740), .ZN(n13533) );
  NAND2_X1 U7264 ( .A1(n13544), .A2(n13543), .ZN(n13539) );
  INV_X1 U7265 ( .A(n13548), .ZN(n10604) );
  AND3_X1 U7266 ( .A1(n8371), .A2(n8370), .A3(n8369), .ZN(n11062) );
  NAND2_X2 U7267 ( .A1(n14855), .A2(n11624), .ZN(n9927) );
  NOR2_X1 U7268 ( .A1(n8357), .A2(n8270), .ZN(n8271) );
  CLKBUF_X2 U7269 ( .A(n9623), .Z(n11978) );
  INV_X1 U7270 ( .A(n9883), .ZN(n9835) );
  INV_X2 U7271 ( .A(n8119), .ZN(n7692) );
  NAND2_X1 U7272 ( .A1(n11966), .A2(n14075), .ZN(n9623) );
  NAND2_X4 U7273 ( .A1(n9970), .A2(n11553), .ZN(n8310) );
  INV_X1 U7274 ( .A(n13749), .ZN(n7348) );
  INV_X1 U7275 ( .A(n13748), .ZN(n10338) );
  INV_X4 U7276 ( .A(n11966), .ZN(n10324) );
  INV_X2 U7277 ( .A(n9091), .ZN(n6433) );
  BUF_X1 U7278 ( .A(n7584), .Z(n9066) );
  NAND2_X4 U7279 ( .A1(n9508), .A2(n10954), .ZN(n9533) );
  CLKBUF_X2 U7280 ( .A(n9500), .Z(n13440) );
  NAND2_X1 U7281 ( .A1(n9475), .A2(n11852), .ZN(n11557) );
  CLKBUF_X1 U7283 ( .A(n7485), .Z(n7486) );
  AND2_X1 U7284 ( .A1(n8470), .A2(n8198), .ZN(n6634) );
  INV_X1 U7285 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n14401) );
  NAND2_X1 U7286 ( .A1(n6440), .A2(n6438), .ZN(P1_U3523) );
  NAND2_X1 U7287 ( .A1(n14209), .A2(n14729), .ZN(n6440) );
  NAND2_X1 U7288 ( .A1(n14121), .A2(n14120), .ZN(n14209) );
  INV_X1 U7289 ( .A(n6437), .ZN(n14121) );
  AOI21_X1 U7290 ( .B1(n14105), .B2(n14183), .A(n6508), .ZN(n6664) );
  OAI21_X1 U7291 ( .B1(n14118), .B2(n13957), .A(n11615), .ZN(n6437) );
  AOI21_X1 U7292 ( .B1(n11614), .B2(n14183), .A(n11613), .ZN(n11615) );
  AOI21_X1 U7293 ( .B1(n11673), .B2(n11672), .A(n11671), .ZN(n11674) );
  NAND2_X1 U7294 ( .A1(n12049), .A2(n8888), .ZN(n8891) );
  OR2_X1 U7295 ( .A1(n12397), .A2(n12403), .ZN(n12398) );
  NAND2_X1 U7296 ( .A1(n12993), .A2(n12986), .ZN(n12996) );
  AND2_X1 U7297 ( .A1(n7256), .A2(n12984), .ZN(n13017) );
  NAND2_X1 U7298 ( .A1(n8748), .A2(n11792), .ZN(n12416) );
  INV_X1 U7299 ( .A(n9107), .ZN(n13180) );
  OR2_X1 U7300 ( .A1(n13029), .A2(n12982), .ZN(n7256) );
  OAI21_X1 U7301 ( .B1(n8664), .B2(n6992), .A(n6990), .ZN(n8690) );
  OR2_X1 U7302 ( .A1(n7079), .A2(n13016), .ZN(n7076) );
  NAND2_X1 U7303 ( .A1(n6892), .A2(n12981), .ZN(n13029) );
  NAND2_X1 U7304 ( .A1(n12987), .A2(n9131), .ZN(n12986) );
  NAND2_X1 U7305 ( .A1(n14128), .A2(n6577), .ZN(n13925) );
  OR2_X1 U7306 ( .A1(n12440), .A2(n8662), .ZN(n8664) );
  XNOR2_X1 U7307 ( .A(n7215), .B(n9064), .ZN(n13437) );
  NAND2_X1 U7308 ( .A1(n13939), .A2(n13938), .ZN(n14128) );
  NAND2_X1 U7309 ( .A1(n13038), .A2(n12979), .ZN(n6892) );
  INV_X1 U7310 ( .A(n12955), .ZN(n13185) );
  NAND2_X1 U7311 ( .A1(n12457), .A2(n8746), .ZN(n12444) );
  INV_X1 U7312 ( .A(n13495), .ZN(n6447) );
  NAND2_X1 U7313 ( .A1(n9060), .A2(n9059), .ZN(n9068) );
  NAND2_X1 U7314 ( .A1(n11579), .A2(n11578), .ZN(n14115) );
  NAND2_X1 U7315 ( .A1(n13970), .A2(n7439), .ZN(n13948) );
  NOR2_X1 U7316 ( .A1(n11838), .A2(n11668), .ZN(n11672) );
  OR2_X1 U7317 ( .A1(n7003), .A2(n7002), .ZN(n7000) );
  NAND2_X1 U7318 ( .A1(n8091), .A2(n8090), .ZN(n13196) );
  XNOR2_X1 U7319 ( .A(n9055), .B(n9054), .ZN(n11975) );
  NAND2_X1 U7320 ( .A1(n8624), .A2(n8623), .ZN(n12468) );
  NAND2_X1 U7321 ( .A1(n11565), .A2(n7432), .ZN(n13970) );
  NOR2_X1 U7323 ( .A1(n13949), .A2(n6449), .ZN(n6448) );
  NAND2_X1 U7324 ( .A1(n11476), .A2(n11475), .ZN(n13928) );
  AND2_X1 U7325 ( .A1(n7123), .A2(n7121), .ZN(n14392) );
  OAI21_X1 U7326 ( .B1(n6460), .B2(n7421), .A(n7419), .ZN(n13995) );
  AND2_X1 U7327 ( .A1(n11525), .A2(n11524), .ZN(n6460) );
  INV_X1 U7328 ( .A(n7439), .ZN(n6449) );
  XNOR2_X1 U7329 ( .A(n8892), .B(n12404), .ZN(n12116) );
  AND2_X1 U7330 ( .A1(n8028), .A2(n8027), .ZN(n13054) );
  AND2_X1 U7331 ( .A1(n8548), .A2(n8547), .ZN(n8550) );
  AND2_X1 U7332 ( .A1(n11791), .A2(n11792), .ZN(n12431) );
  NAND2_X1 U7333 ( .A1(n6446), .A2(n11510), .ZN(n14041) );
  CLKBUF_X1 U7334 ( .A(n8738), .Z(n6683) );
  NAND2_X1 U7335 ( .A1(n14349), .A2(n14348), .ZN(n14354) );
  OAI21_X1 U7336 ( .B1(n12963), .B2(n6878), .A(n6877), .ZN(n6876) );
  NAND2_X1 U7337 ( .A1(n11569), .A2(n11568), .ZN(n13978) );
  NAND2_X1 U7338 ( .A1(n6443), .A2(n11506), .ZN(n14055) );
  NAND2_X1 U7339 ( .A1(n6443), .A2(n6441), .ZN(n6446) );
  NAND2_X1 U7340 ( .A1(n7990), .A2(n7989), .ZN(n13226) );
  NAND2_X1 U7341 ( .A1(n11423), .A2(n6444), .ZN(n6443) );
  NAND2_X1 U7342 ( .A1(n13427), .A2(n13426), .ZN(n13425) );
  NAND2_X1 U7343 ( .A1(n7351), .A2(n7350), .ZN(n11224) );
  INV_X1 U7344 ( .A(n11331), .ZN(n11245) );
  NAND2_X1 U7345 ( .A1(n11541), .A2(n11540), .ZN(n14010) );
  NAND2_X1 U7346 ( .A1(n7413), .A2(n7412), .ZN(n11242) );
  NAND2_X1 U7347 ( .A1(n11022), .A2(n8849), .ZN(n11164) );
  NAND2_X1 U7348 ( .A1(n11171), .A2(n11714), .ZN(n11395) );
  NOR2_X1 U7349 ( .A1(n11504), .A2(n6445), .ZN(n6444) );
  AOI21_X1 U7350 ( .B1(n14987), .B2(n12317), .A(n15024), .ZN(n12318) );
  NAND2_X1 U7351 ( .A1(n10918), .A2(n10917), .ZN(n10928) );
  NOR2_X1 U7352 ( .A1(n6442), .A2(n11511), .ZN(n6441) );
  INV_X1 U7353 ( .A(n6452), .ZN(n6451) );
  NAND2_X1 U7354 ( .A1(n11172), .A2(n11821), .ZN(n11171) );
  INV_X1 U7355 ( .A(n11506), .ZN(n6442) );
  XNOR2_X1 U7356 ( .A(n7964), .B(SI_20_), .ZN(n7963) );
  INV_X1 U7357 ( .A(n11422), .ZN(n6445) );
  NAND2_X1 U7358 ( .A1(n6782), .A2(n6780), .ZN(n11859) );
  NAND2_X1 U7359 ( .A1(n7006), .A2(n6494), .ZN(n11066) );
  NAND2_X1 U7360 ( .A1(n10845), .A2(n10844), .ZN(n10847) );
  NAND2_X1 U7361 ( .A1(n10956), .A2(n6542), .ZN(n7006) );
  NAND2_X1 U7362 ( .A1(n10503), .A2(n10511), .ZN(n10845) );
  NAND2_X1 U7363 ( .A1(n10564), .A2(n10491), .ZN(n10503) );
  NAND2_X1 U7364 ( .A1(n7859), .A2(n7858), .ZN(n13258) );
  NAND2_X1 U7365 ( .A1(n10800), .A2(n10801), .ZN(n10956) );
  NAND2_X1 U7366 ( .A1(n11227), .A2(n11226), .ZN(n13612) );
  AND4_X1 U7367 ( .A1(n8687), .A2(n8686), .A3(n8685), .A4(n8684), .ZN(n12433)
         );
  NAND2_X1 U7368 ( .A1(n6450), .A2(n7407), .ZN(n10278) );
  NAND2_X1 U7369 ( .A1(n7795), .A2(n7794), .ZN(n11152) );
  NAND2_X1 U7370 ( .A1(n7734), .A2(n7733), .ZN(n10875) );
  NAND2_X1 U7371 ( .A1(n10915), .A2(n10914), .ZN(n14575) );
  NAND2_X1 U7372 ( .A1(n10218), .A2(n7406), .ZN(n6450) );
  NAND2_X1 U7373 ( .A1(n10212), .A2(n10211), .ZN(n10218) );
  NAND2_X1 U7374 ( .A1(n9851), .A2(n13471), .ZN(n10212) );
  AND2_X2 U7375 ( .A1(n7707), .A2(n7706), .ZN(n14923) );
  AND2_X2 U7376 ( .A1(n10187), .A2(n15114), .ZN(n14462) );
  OAI21_X1 U7377 ( .B1(n10397), .B2(n15060), .A(n6541), .ZN(n7035) );
  NOR2_X1 U7378 ( .A1(n10443), .A2(n12864), .ZN(n10245) );
  XNOR2_X1 U7379 ( .A(n14316), .B(n7140), .ZN(n15157) );
  AND2_X1 U7380 ( .A1(n15107), .A2(n8726), .ZN(n15101) );
  NAND2_X1 U7381 ( .A1(n7141), .A2(n14314), .ZN(n14316) );
  NAND2_X1 U7382 ( .A1(n10490), .A2(n10489), .ZN(n13572) );
  AND4_X1 U7383 ( .A1(n8348), .A2(n8347), .A3(n8346), .A4(n8345), .ZN(n10747)
         );
  NAND3_X1 U7384 ( .A1(n6636), .A2(n8272), .A3(n8273), .ZN(n10087) );
  NAND4_X2 U7385 ( .A1(n8309), .A2(n8308), .A3(n8307), .A4(n8306), .ZN(n12149)
         );
  CLKBUF_X1 U7386 ( .A(n15105), .Z(n6670) );
  NAND2_X1 U7387 ( .A1(n7348), .A2(n7349), .ZN(n13536) );
  OR2_X1 U7388 ( .A1(n14729), .A2(n6439), .ZN(n6438) );
  AND4_X1 U7389 ( .A1(n8292), .A2(n8291), .A3(n8290), .A4(n8289), .ZN(n15105)
         );
  NAND2_X1 U7390 ( .A1(n7033), .A2(n7032), .ZN(n10353) );
  NAND2_X1 U7391 ( .A1(n10265), .A2(n10264), .ZN(n13556) );
  INV_X1 U7392 ( .A(n10597), .ZN(n7349) );
  NAND2_X1 U7393 ( .A1(n9739), .A2(n9738), .ZN(n9741) );
  OR2_X1 U7394 ( .A1(n9282), .A2(n11841), .ZN(n7015) );
  AND2_X1 U7395 ( .A1(n9676), .A2(n9675), .ZN(n10597) );
  NAND2_X1 U7396 ( .A1(n13529), .A2(n13530), .ZN(n9712) );
  BUF_X2 U7397 ( .A(n8293), .Z(n11663) );
  AND2_X1 U7398 ( .A1(n10095), .A2(n9983), .ZN(n9984) );
  BUF_X2 U7399 ( .A(n8293), .Z(n8430) );
  NAND2_X1 U7400 ( .A1(n6649), .A2(n6650), .ZN(n9330) );
  CLKBUF_X1 U7401 ( .A(n12304), .Z(n6717) );
  OR2_X1 U7402 ( .A1(n9433), .A2(n9432), .ZN(n6845) );
  INV_X2 U7403 ( .A(n6591), .ZN(n13703) );
  OR2_X1 U7404 ( .A1(n9710), .A2(n13523), .ZN(n13529) );
  NAND4_X2 U7405 ( .A1(n9524), .A2(n9523), .A3(n9522), .A4(n9521), .ZN(n9710)
         );
  NAND2_X2 U7406 ( .A1(n9501), .A2(n13440), .ZN(n14075) );
  NAND4_X1 U7407 ( .A1(n7520), .A2(n7519), .A3(n7518), .A4(n7517), .ZN(n12870)
         );
  OR2_X1 U7408 ( .A1(n10072), .A2(n9979), .ZN(n10094) );
  CLKBUF_X1 U7409 ( .A(n9632), .Z(n6688) );
  INV_X1 U7410 ( .A(n10616), .ZN(n11682) );
  NAND2_X1 U7411 ( .A1(n12729), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8217) );
  INV_X1 U7412 ( .A(n13957), .ZN(n6436) );
  OR2_X1 U7413 ( .A1(n8762), .A2(n8783), .ZN(n6650) );
  NAND2_X1 U7414 ( .A1(n9916), .A2(n13001), .ZN(n14936) );
  AND2_X2 U7415 ( .A1(n9533), .A2(n9544), .ZN(n11966) );
  AND2_X1 U7416 ( .A1(n9978), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10072) );
  XNOR2_X1 U7417 ( .A(n6796), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10616) );
  AND2_X1 U7418 ( .A1(n6526), .A2(n6854), .ZN(n14266) );
  NOR2_X1 U7419 ( .A1(n8761), .A2(n8763), .ZN(n8783) );
  CLKBUF_X3 U7420 ( .A(n11557), .Z(n6467) );
  NAND2_X1 U7421 ( .A1(n8218), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8219) );
  MUX2_X1 U7422 ( .A(n8765), .B(n8760), .S(P3_IR_REG_25__SCAN_IN), .Z(n8761)
         );
  XNOR2_X1 U7423 ( .A(n8209), .B(n8208), .ZN(n8210) );
  OR2_X1 U7424 ( .A1(n8507), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8534) );
  MUX2_X1 U7425 ( .A(n8765), .B(n8764), .S(P3_IR_REG_26__SCAN_IN), .Z(n8766)
         );
  INV_X1 U7426 ( .A(n6426), .ZN(n13450) );
  NOR2_X1 U7427 ( .A1(n8715), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n6797) );
  OR2_X1 U7428 ( .A1(n7608), .A2(n7607), .ZN(n7636) );
  INV_X1 U7429 ( .A(n13286), .ZN(n7516) );
  NAND2_X2 U7430 ( .A1(n9475), .A2(n9474), .ZN(n11606) );
  NAND2_X1 U7431 ( .A1(n7514), .A2(n13282), .ZN(n13286) );
  XNOR2_X1 U7432 ( .A(n9493), .B(P1_IR_REG_20__SCAN_IN), .ZN(n13442) );
  OR2_X1 U7433 ( .A1(n6860), .A2(n14262), .ZN(n6855) );
  NOR2_X1 U7434 ( .A1(n10056), .A2(n7016), .ZN(n9977) );
  CLKBUF_X1 U7435 ( .A(n11202), .Z(n6700) );
  AND2_X1 U7436 ( .A1(n8756), .A2(n7209), .ZN(n8763) );
  OR2_X1 U7437 ( .A1(n8440), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8462) );
  OAI21_X1 U7438 ( .B1(n9495), .B2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9283) );
  NAND2_X2 U7439 ( .A1(n9496), .A2(n9495), .ZN(n13920) );
  XNOR2_X1 U7440 ( .A(n7510), .B(P2_IR_REG_30__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U7441 ( .A1(n13282), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7510) );
  INV_X2 U7442 ( .A(n14238), .ZN(n10724) );
  XNOR2_X1 U7443 ( .A(n9287), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U7444 ( .A1(n14236), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9359) );
  NOR2_X1 U7445 ( .A1(n10043), .A2(n15119), .ZN(n10042) );
  AND2_X1 U7446 ( .A1(n7436), .A2(n9195), .ZN(n9360) );
  NAND2_X2 U7447 ( .A1(n9617), .A2(P2_U3088), .ZN(n13303) );
  NAND2_X1 U7448 ( .A1(n6634), .A2(n8331), .ZN(n6799) );
  NOR2_X1 U7449 ( .A1(n9193), .A2(n9192), .ZN(n9194) );
  AND2_X2 U7450 ( .A1(n6937), .A2(n6936), .ZN(n9212) );
  AND3_X1 U7451 ( .A1(n8195), .A2(n8194), .A3(n8193), .ZN(n8470) );
  NAND2_X1 U7452 ( .A1(n6638), .A2(n6637), .ZN(n8263) );
  AND3_X1 U7453 ( .A1(n7463), .A2(n7462), .A3(n7461), .ZN(n6474) );
  NOR2_X1 U7454 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n7461) );
  NOR2_X1 U7455 ( .A1(P3_IR_REG_10__SCAN_IN), .A2(P3_IR_REG_6__SCAN_IN), .ZN(
        n8195) );
  NOR2_X1 U7456 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_7__SCAN_IN), .ZN(
        n8194) );
  NOR2_X1 U7457 ( .A1(P3_IR_REG_8__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n8193) );
  NOR2_X1 U7458 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7463) );
  NOR2_X1 U7459 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n7462) );
  INV_X1 U7460 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n12257) );
  NOR2_X1 U7461 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n9178) );
  NOR2_X1 U7462 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n9179) );
  INV_X4 U7463 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  INV_X1 U7464 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n9874) );
  NOR2_X1 U7465 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n7458) );
  NOR2_X1 U7466 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n9188) );
  INV_X1 U7467 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9286) );
  INV_X1 U7468 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n9284) );
  INV_X1 U7469 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n6439) );
  NOR2_X1 U7470 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n7457) );
  NOR2_X1 U7471 ( .A1(P3_IR_REG_17__SCAN_IN), .A2(P3_IR_REG_18__SCAN_IN), .ZN(
        n8212) );
  INV_X1 U7472 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n9997) );
  INV_X1 U7473 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n6638) );
  INV_X1 U7474 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6637) );
  INV_X4 U7475 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7476 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7199) );
  INV_X1 U7477 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n9276) );
  NOR2_X1 U7478 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n9183) );
  INV_X1 U7479 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n9223) );
  NAND2_X1 U7480 ( .A1(n11423), .A2(n11422), .ZN(n11505) );
  NAND2_X1 U7481 ( .A1(n14041), .A2(n14040), .ZN(n11525) );
  AOI21_X1 U7482 ( .B1(n13923), .B2(n7427), .A(n6447), .ZN(n11589) );
  NAND2_X2 U7483 ( .A1(n13925), .A2(n13924), .ZN(n13923) );
  NAND2_X1 U7484 ( .A1(n13995), .A2(n13996), .ZN(n11565) );
  NAND2_X1 U7485 ( .A1(n10565), .A2(n13478), .ZN(n10564) );
  OAI21_X2 U7486 ( .B1(n7413), .B2(n6435), .A(n6451), .ZN(n11331) );
  NAND2_X1 U7487 ( .A1(n12285), .A2(n8726), .ZN(n15103) );
  XNOR2_X1 U7488 ( .A(n14260), .B(n14261), .ZN(n14305) );
  XNOR2_X1 U7489 ( .A(n6682), .B(P1_ADDR_REG_1__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U7490 ( .A1(n13923), .A2(n7424), .ZN(n7426) );
  AND2_X2 U7491 ( .A1(n8785), .A2(n8203), .ZN(n8756) );
  OAI21_X1 U7492 ( .B1(n8950), .B2(n8949), .A(n8948), .ZN(n8952) );
  NOR2_X2 U7493 ( .A1(n7832), .A2(P2_IR_REG_15__SCAN_IN), .ZN(n7853) );
  CLKBUF_X1 U7494 ( .A(n12059), .Z(n6454) );
  AND2_X1 U7495 ( .A1(n10528), .A2(n7010), .ZN(n6455) );
  NAND2_X1 U7496 ( .A1(n12116), .A2(n6456), .ZN(n6457) );
  NAND2_X1 U7497 ( .A1(n6432), .A2(n12115), .ZN(n6458) );
  NAND2_X1 U7498 ( .A1(n6457), .A2(n6458), .ZN(n12122) );
  INV_X1 U7499 ( .A(n12115), .ZN(n6456) );
  INV_X1 U7501 ( .A(n6460), .ZN(n14032) );
  OR2_X2 U7502 ( .A1(n8173), .A2(n8174), .ZN(n9170) );
  OAI21_X1 U7503 ( .B1(n8969), .B2(n7332), .A(n7328), .ZN(n8977) );
  CLKBUF_X1 U7504 ( .A(n7226), .Z(n6461) );
  NAND2_X1 U7505 ( .A1(n12088), .A2(n8877), .ZN(n12043) );
  OAI222_X1 U7506 ( .A1(n10724), .A2(n11646), .B1(P1_U3086), .B2(n9363), .C1(
        n13446), .C2(n14252), .ZN(P1_U3325) );
  NOR2_X2 U7507 ( .A1(n13900), .A2(n13883), .ZN(n13882) );
  OR2_X1 U7508 ( .A1(n9360), .A2(n10377), .ZN(n9361) );
  NOR2_X2 U7509 ( .A1(n14344), .A2(n14604), .ZN(n14607) );
  AOI21_X2 U7510 ( .B1(n14057), .B2(n14056), .A(n11593), .ZN(n14038) );
  AND2_X2 U7511 ( .A1(n6463), .A2(n7504), .ZN(n6485) );
  NAND2_X2 U7512 ( .A1(n9711), .A2(n9517), .ZN(n13524) );
  NAND2_X1 U7513 ( .A1(n7426), .A2(n6527), .ZN(n14107) );
  OAI222_X1 U7515 ( .A1(n12744), .A2(n12739), .B1(P3_U3151), .B2(n8211), .C1(
        n12747), .C2(n12738), .ZN(P3_U3267) );
  AOI21_X1 U7516 ( .B1(n7274), .B2(n7272), .A(n13667), .ZN(n6720) );
  NOR2_X2 U7517 ( .A1(n8374), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8388) );
  NOR2_X2 U7518 ( .A1(n12316), .A2(n14971), .ZN(n14990) );
  AND2_X1 U7519 ( .A1(n14856), .A2(n7504), .ZN(n6462) );
  AND2_X1 U7520 ( .A1(n14856), .A2(n7504), .ZN(n14816) );
  CLKBUF_X1 U7521 ( .A(n7503), .Z(n6463) );
  XNOR2_X1 U7522 ( .A(n7315), .B(n7314), .ZN(n7503) );
  XNOR2_X1 U7523 ( .A(n12325), .B(n6698), .ZN(n14442) );
  NOR2_X2 U7524 ( .A1(n10567), .A2(n13572), .ZN(n10566) );
  BUF_X8 U7525 ( .A(n11606), .Z(n6465) );
  BUF_X8 U7526 ( .A(n13703), .Z(n6466) );
  NOR2_X2 U7527 ( .A1(n8534), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8536) );
  NOR2_X2 U7528 ( .A1(n10120), .A2(n13548), .ZN(n10234) );
  XNOR2_X1 U7529 ( .A(n9290), .B(n9289), .ZN(n9299) );
  NAND2_X1 U7530 ( .A1(n8953), .A2(n7345), .ZN(n7344) );
  NOR2_X1 U7531 ( .A1(n12479), .A2(n11775), .ZN(n6823) );
  NAND2_X1 U7532 ( .A1(n6662), .A2(n6661), .ZN(n7326) );
  INV_X1 U7533 ( .A(n9034), .ZN(n6661) );
  OR2_X1 U7534 ( .A1(n8173), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n7472) );
  INV_X1 U7535 ( .A(n10283), .ZN(n7359) );
  AND2_X1 U7536 ( .A1(n7358), .A2(n13476), .ZN(n7357) );
  OR2_X1 U7537 ( .A1(n10282), .A2(n7359), .ZN(n7358) );
  NAND2_X1 U7538 ( .A1(n6926), .A2(n6924), .ZN(n7875) );
  AOI21_X1 U7539 ( .B1(n6928), .B2(n6930), .A(n6925), .ZN(n6924) );
  INV_X1 U7540 ( .A(n7871), .ZN(n6925) );
  AND2_X1 U7541 ( .A1(n13220), .A2(n13094), .ZN(n13077) );
  NAND2_X1 U7542 ( .A1(n13156), .A2(n13157), .ZN(n12963) );
  AND2_X1 U7543 ( .A1(n14081), .A2(n13616), .ZN(n6912) );
  NOR2_X1 U7544 ( .A1(n8958), .A2(n8957), .ZN(n8960) );
  INV_X1 U7545 ( .A(n8972), .ZN(n7336) );
  OR2_X1 U7546 ( .A1(n8974), .A2(n8973), .ZN(n7337) );
  AOI21_X1 U7547 ( .B1(n13606), .B2(n13605), .A(n6466), .ZN(n13625) );
  AND2_X1 U7548 ( .A1(n7311), .A2(n7313), .ZN(n7310) );
  NAND2_X1 U7549 ( .A1(n6469), .A2(n7312), .ZN(n7311) );
  AOI21_X1 U7550 ( .B1(n6824), .B2(n6823), .A(n6821), .ZN(n11784) );
  OAI21_X1 U7551 ( .B1(n6993), .B2(n6992), .A(n8688), .ZN(n6991) );
  INV_X1 U7552 ( .A(n7827), .ZN(n7830) );
  NOR2_X1 U7553 ( .A1(n7768), .A2(n7222), .ZN(n7221) );
  INV_X1 U7554 ( .A(n7749), .ZN(n7222) );
  INV_X1 U7555 ( .A(n12736), .ZN(n8223) );
  INV_X1 U7556 ( .A(n11998), .ZN(n8220) );
  INV_X1 U7557 ( .A(n7208), .ZN(n7207) );
  AOI21_X1 U7558 ( .B1(n12494), .B2(n8743), .A(n6550), .ZN(n7208) );
  OR2_X1 U7559 ( .A1(n12472), .A2(n12482), .ZN(n11779) );
  NOR2_X1 U7560 ( .A1(n6477), .A2(n6553), .ZN(n6963) );
  INV_X1 U7561 ( .A(n11755), .ZN(n8739) );
  NAND2_X1 U7562 ( .A1(n11209), .A2(n8403), .ZN(n11308) );
  NAND2_X1 U7563 ( .A1(n8767), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8209) );
  NOR2_X2 U7564 ( .A1(n6799), .A2(n7194), .ZN(n8785) );
  NAND2_X1 U7565 ( .A1(n7195), .A2(n6505), .ZN(n7194) );
  INV_X1 U7566 ( .A(n7196), .ZN(n7195) );
  INV_X1 U7567 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n8213) );
  OAI21_X1 U7568 ( .B1(P2_DATAO_REG_12__SCAN_IN), .B2(n9645), .A(n8241), .ZN(
        n8242) );
  NAND2_X1 U7569 ( .A1(n6735), .A2(n6734), .ZN(n8241) );
  AOI21_X1 U7570 ( .B1(n6736), .B2(n7044), .A(n6609), .ZN(n6734) );
  INV_X1 U7571 ( .A(n8240), .ZN(n7045) );
  INV_X1 U7572 ( .A(n6700), .ZN(n9129) );
  NOR2_X1 U7573 ( .A1(n9147), .A2(n6712), .ZN(n6711) );
  NAND2_X1 U7574 ( .A1(n13208), .A2(n12980), .ZN(n7089) );
  AOI21_X1 U7575 ( .B1(n7088), .B2(n13037), .A(n7086), .ZN(n7085) );
  NAND2_X1 U7576 ( .A1(n13053), .A2(n7090), .ZN(n7088) );
  INV_X1 U7577 ( .A(n7089), .ZN(n7086) );
  NOR2_X1 U7578 ( .A1(n13092), .A2(n7107), .ZN(n7106) );
  INV_X1 U7579 ( .A(n12936), .ZN(n7107) );
  AND2_X1 U7580 ( .A1(n10879), .A2(n8970), .ZN(n10578) );
  INV_X1 U7581 ( .A(n7814), .ZN(n7464) );
  AND2_X1 U7582 ( .A1(n7484), .A2(n7314), .ZN(n8136) );
  INV_X1 U7583 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8135) );
  INV_X1 U7584 ( .A(n13943), .ZN(n11953) );
  NOR2_X2 U7585 ( .A1(n10948), .A2(n13601), .ZN(n11096) );
  NAND2_X1 U7586 ( .A1(n14042), .A2(n14028), .ZN(n14025) );
  INV_X1 U7587 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n9293) );
  INV_X1 U7588 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n9292) );
  INV_X1 U7589 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n9291) );
  NAND2_X1 U7590 ( .A1(n7227), .A2(n8046), .ZN(n8065) );
  NAND2_X1 U7591 ( .A1(n8044), .A2(n8043), .ZN(n7227) );
  INV_X1 U7592 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n9191) );
  INV_X1 U7593 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n9190) );
  INV_X1 U7594 ( .A(n6929), .ZN(n6928) );
  OAI21_X1 U7595 ( .B1(n6932), .B2(n6930), .A(n7850), .ZN(n6929) );
  INV_X1 U7596 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U7597 ( .A1(n14263), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6859) );
  OR2_X1 U7598 ( .A1(n14263), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6860) );
  INV_X1 U7599 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14270) );
  OAI21_X1 U7600 ( .B1(n14287), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n14286), .ZN(
        n14340) );
  OR2_X1 U7601 ( .A1(n14338), .A2(n14337), .ZN(n14286) );
  OAI22_X1 U7602 ( .A1(n6792), .A2(n6789), .B1(n6795), .B2(n6791), .ZN(n6788)
         );
  NOR2_X1 U7603 ( .A1(n6795), .A2(n12116), .ZN(n6789) );
  INV_X1 U7604 ( .A(n8894), .ZN(n7002) );
  INV_X1 U7605 ( .A(n7004), .ZN(n7003) );
  OAI22_X1 U7606 ( .A1(n11999), .A2(n7005), .B1(n12388), .B2(n8893), .ZN(n7004) );
  INV_X1 U7607 ( .A(n8837), .ZN(n12031) );
  NAND2_X1 U7608 ( .A1(n11685), .A2(n15101), .ZN(n8817) );
  INV_X1 U7609 ( .A(n10087), .ZN(n6635) );
  NAND2_X1 U7610 ( .A1(n7008), .A2(n6594), .ZN(n7007) );
  NAND2_X1 U7611 ( .A1(n10008), .A2(n10007), .ZN(n10355) );
  NAND2_X1 U7612 ( .A1(n7035), .A2(n7034), .ZN(n10672) );
  INV_X1 U7613 ( .A(n10399), .ZN(n7034) );
  INV_X1 U7614 ( .A(n7200), .ZN(n6668) );
  INV_X1 U7615 ( .A(n12416), .ZN(n6669) );
  INV_X1 U7616 ( .A(n7203), .ZN(n7202) );
  NAND2_X1 U7617 ( .A1(n6967), .A2(n6966), .ZN(n12480) );
  AOI21_X1 U7618 ( .B1(n6968), .B2(n6971), .A(n6552), .ZN(n6966) );
  AOI21_X1 U7619 ( .B1(n7183), .B2(n7186), .A(n11732), .ZN(n7182) );
  AND2_X1 U7620 ( .A1(n9970), .A2(n9617), .ZN(n8293) );
  OR2_X1 U7621 ( .A1(n11848), .A2(n11682), .ZN(n15138) );
  OAI21_X1 U7622 ( .B1(n8626), .B2(n8625), .A(n6613), .ZN(n7050) );
  NAND2_X1 U7623 ( .A1(n8584), .A2(n8213), .ZN(n8715) );
  NAND2_X1 U7624 ( .A1(n6721), .A2(n7039), .ZN(n8569) );
  NAND2_X1 U7625 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n7040), .ZN(n7039) );
  NAND2_X1 U7626 ( .A1(n8551), .A2(n8552), .ZN(n6721) );
  AOI21_X1 U7627 ( .B1(n8382), .B2(n6728), .A(n6725), .ZN(n6724) );
  NAND2_X1 U7628 ( .A1(n6726), .A2(n8237), .ZN(n6725) );
  NAND2_X1 U7629 ( .A1(n6737), .A2(n6740), .ZN(n8366) );
  AOI21_X1 U7630 ( .B1(n6741), .B2(n8349), .A(n6561), .ZN(n6740) );
  NAND2_X1 U7631 ( .A1(n11459), .A2(n7870), .ZN(n7889) );
  NAND2_X1 U7632 ( .A1(n7156), .A2(n6515), .ZN(n10645) );
  INV_X1 U7633 ( .A(n10646), .ZN(n7155) );
  AND2_X1 U7634 ( .A1(n7747), .A2(n7724), .ZN(n7174) );
  INV_X1 U7635 ( .A(n12870), .ZN(n11471) );
  OR2_X1 U7636 ( .A1(n7882), .A2(n7881), .ZN(n7905) );
  AND2_X1 U7637 ( .A1(n8078), .A2(n8077), .ZN(n12983) );
  AND2_X1 U7638 ( .A1(n7911), .A2(n7910), .ZN(n12961) );
  AND3_X1 U7639 ( .A1(n7841), .A2(n7840), .A3(n7839), .ZN(n11364) );
  AND4_X1 U7640 ( .A1(n7781), .A2(n7780), .A3(n7779), .A4(n7778), .ZN(n11122)
         );
  AND2_X1 U7641 ( .A1(n11470), .A2(n13286), .ZN(n7552) );
  XNOR2_X1 U7642 ( .A(n12896), .B(n12895), .ZN(n12883) );
  NOR2_X1 U7643 ( .A1(n13190), .A2(n6952), .ZN(n6950) );
  AND2_X1 U7644 ( .A1(n9087), .A2(n9086), .ZN(n12955) );
  NOR2_X1 U7645 ( .A1(n13069), .A2(n12939), .ZN(n13049) );
  NAND2_X1 U7646 ( .A1(n6884), .A2(n6484), .ZN(n6883) );
  INV_X1 U7647 ( .A(n6887), .ZN(n6884) );
  OAI22_X1 U7648 ( .A1(n13161), .A2(n12960), .B1(n13255), .B2(n12959), .ZN(
        n13156) );
  OR2_X1 U7649 ( .A1(n10875), .A2(n10736), .ZN(n10879) );
  OAI21_X1 U7650 ( .B1(n9925), .B2(n6869), .A(n10153), .ZN(n6868) );
  NAND2_X1 U7651 ( .A1(n7524), .A2(n11553), .ZN(n7584) );
  AND2_X1 U7652 ( .A1(n8005), .A2(n8004), .ZN(n13220) );
  AND2_X1 U7653 ( .A1(n7835), .A2(n7834), .ZN(n11375) );
  AND2_X1 U7654 ( .A1(n14856), .A2(n9171), .ZN(n14943) );
  AND2_X1 U7655 ( .A1(n11202), .A2(n11050), .ZN(n14856) );
  OR2_X1 U7656 ( .A1(n11447), .A2(n8150), .ZN(n9176) );
  INV_X1 U7657 ( .A(n10812), .ZN(n7404) );
  AOI21_X1 U7658 ( .B1(n7373), .B2(n7376), .A(n6547), .ZN(n7371) );
  NAND2_X1 U7659 ( .A1(n6774), .A2(n6496), .ZN(n6773) );
  INV_X1 U7660 ( .A(n13378), .ZN(n6774) );
  NAND2_X1 U7661 ( .A1(n13466), .A2(n13465), .ZN(n13883) );
  NOR2_X1 U7662 ( .A1(n13495), .A2(n7428), .ZN(n7424) );
  AOI21_X1 U7663 ( .B1(n6899), .B2(n6901), .A(n6564), .ZN(n6897) );
  NOR2_X1 U7664 ( .A1(n7434), .A2(n7433), .ZN(n7432) );
  INV_X1 U7665 ( .A(n11564), .ZN(n7433) );
  AND2_X1 U7666 ( .A1(n7352), .A2(n13604), .ZN(n7350) );
  NAND2_X1 U7667 ( .A1(n7354), .A2(n6514), .ZN(n10510) );
  INV_X1 U7668 ( .A(n13478), .ZN(n6902) );
  INV_X1 U7669 ( .A(n14183), .ZN(n14166) );
  XNOR2_X1 U7670 ( .A(n9201), .B(P1_IR_REG_23__SCAN_IN), .ZN(n9288) );
  OR2_X1 U7671 ( .A1(n14248), .A2(n13864), .ZN(n9237) );
  NAND2_X1 U7672 ( .A1(n9194), .A2(n9195), .ZN(n9294) );
  NAND2_X1 U7673 ( .A1(n6708), .A2(n7812), .ZN(n7829) );
  NAND2_X1 U7674 ( .A1(n7730), .A2(n7729), .ZN(n7750) );
  INV_X1 U7675 ( .A(n6472), .ZN(n7147) );
  NAND2_X1 U7676 ( .A1(n6539), .A2(n6820), .ZN(n6755) );
  INV_X1 U7677 ( .A(n6754), .ZN(n6753) );
  NAND2_X1 U7678 ( .A1(n7437), .A2(n11845), .ZN(n6819) );
  INV_X1 U7679 ( .A(n14520), .ZN(n14498) );
  AND2_X1 U7680 ( .A1(n14492), .A2(n7808), .ZN(n7172) );
  OAI21_X1 U7681 ( .B1(n12901), .B2(n14786), .A(n6691), .ZN(n6690) );
  AOI21_X1 U7682 ( .B1(n12902), .B2(n14765), .A(n14805), .ZN(n6691) );
  NOR2_X1 U7683 ( .A1(n7500), .A2(n7440), .ZN(n7501) );
  NAND2_X1 U7684 ( .A1(n7855), .A2(n7495), .ZN(n7502) );
  XNOR2_X1 U7685 ( .A(n7259), .B(n12944), .ZN(n13188) );
  AOI21_X1 U7686 ( .B1(n6922), .B2(n14814), .A(n12951), .ZN(n13187) );
  NAND2_X1 U7687 ( .A1(n11448), .A2(n9199), .ZN(n9544) );
  AND2_X1 U7688 ( .A1(n14244), .A2(n14248), .ZN(n9199) );
  NAND2_X1 U7689 ( .A1(n6862), .A2(n6861), .ZN(n14348) );
  NOR2_X1 U7690 ( .A1(n14347), .A2(n6472), .ZN(n6861) );
  AOI22_X1 U7691 ( .A1(n6424), .A2(n6433), .B1(n12870), .B2(n9091), .ZN(n8931)
         );
  INV_X1 U7692 ( .A(n13555), .ZN(n7291) );
  NAND2_X1 U7693 ( .A1(n8939), .A2(n8938), .ZN(n8943) );
  AOI22_X1 U7694 ( .A1(n10177), .A2(n9080), .B1(n9091), .B2(n12867), .ZN(n8949) );
  INV_X1 U7695 ( .A(n13574), .ZN(n7288) );
  OR2_X1 U7696 ( .A1(n7335), .A2(n7331), .ZN(n7330) );
  NOR2_X1 U7697 ( .A1(n8967), .A2(n8968), .ZN(n7331) );
  NOR2_X1 U7698 ( .A1(n7338), .A2(n7336), .ZN(n7335) );
  AND2_X1 U7699 ( .A1(n10578), .A2(n7334), .ZN(n7333) );
  NAND2_X1 U7700 ( .A1(n7338), .A2(n7336), .ZN(n7334) );
  INV_X1 U7701 ( .A(n13602), .ZN(n7280) );
  AOI21_X1 U7702 ( .B1(n6653), .B2(n8987), .A(n8986), .ZN(n8990) );
  NAND2_X1 U7703 ( .A1(n6833), .A2(n11695), .ZN(n6832) );
  NAND2_X1 U7704 ( .A1(n11692), .A2(n11691), .ZN(n6833) );
  INV_X1 U7705 ( .A(n11694), .ZN(n6831) );
  NOR2_X1 U7706 ( .A1(n13663), .A2(n13664), .ZN(n7275) );
  OAI21_X1 U7707 ( .B1(n11701), .B2(n11709), .A(n11808), .ZN(n6838) );
  NAND2_X1 U7708 ( .A1(n6837), .A2(n11804), .ZN(n6836) );
  INV_X1 U7709 ( .A(n11702), .ZN(n6837) );
  NOR2_X1 U7710 ( .A1(n7322), .A2(n9016), .ZN(n7319) );
  INV_X1 U7711 ( .A(n9018), .ZN(n7322) );
  INV_X1 U7712 ( .A(n9021), .ZN(n7318) );
  NOR2_X1 U7713 ( .A1(n9018), .A2(n9017), .ZN(n7323) );
  INV_X1 U7714 ( .A(n7319), .ZN(n7316) );
  NAND2_X1 U7715 ( .A1(n7321), .A2(n9020), .ZN(n7320) );
  INV_X1 U7716 ( .A(n7323), .ZN(n7321) );
  NAND2_X1 U7717 ( .A1(n7281), .A2(n7282), .ZN(n13680) );
  NAND2_X1 U7718 ( .A1(n7285), .A2(n13675), .ZN(n7282) );
  INV_X1 U7719 ( .A(n13676), .ZN(n7285) );
  NOR2_X1 U7720 ( .A1(n7307), .A2(n7313), .ZN(n7309) );
  AOI21_X1 U7721 ( .B1(n7310), .B2(n7307), .A(n7306), .ZN(n7305) );
  INV_X1 U7722 ( .A(n9031), .ZN(n7306) );
  INV_X1 U7723 ( .A(n7310), .ZN(n7308) );
  OAI21_X1 U7724 ( .B1(n9025), .B2(n9023), .A(n9022), .ZN(n9027) );
  OR2_X1 U7725 ( .A1(n7309), .A2(n7305), .ZN(n7304) );
  NAND2_X1 U7726 ( .A1(n11768), .A2(n12525), .ZN(n6828) );
  NAND2_X1 U7727 ( .A1(n11767), .A2(n11766), .ZN(n6827) );
  INV_X1 U7728 ( .A(n11801), .ZN(n6813) );
  NAND2_X1 U7729 ( .A1(n6809), .A2(n6810), .ZN(n6814) );
  INV_X1 U7730 ( .A(n11795), .ZN(n6810) );
  NOR2_X1 U7731 ( .A1(n6815), .A2(n11789), .ZN(n6811) );
  INV_X1 U7732 ( .A(n12431), .ZN(n6815) );
  INV_X1 U7733 ( .A(n6814), .ZN(n6804) );
  AND2_X1 U7734 ( .A1(n7269), .A2(n13692), .ZN(n7268) );
  INV_X1 U7735 ( .A(n13691), .ZN(n7269) );
  NAND2_X1 U7736 ( .A1(n6808), .A2(n11835), .ZN(n6801) );
  INV_X1 U7737 ( .A(n8676), .ZN(n6992) );
  NOR2_X1 U7738 ( .A1(n8611), .A2(n6973), .ZN(n6972) );
  INV_X1 U7739 ( .A(n8566), .ZN(n6973) );
  INV_X1 U7740 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n7455) );
  INV_X1 U7741 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n7454) );
  INV_X1 U7742 ( .A(n8161), .ZN(n7233) );
  NAND2_X1 U7743 ( .A1(n7920), .A2(n9809), .ZN(n7941) );
  NAND2_X1 U7744 ( .A1(n11839), .A2(n6747), .ZN(n6746) );
  AND2_X1 U7745 ( .A1(n11835), .A2(n6748), .ZN(n6747) );
  NOR2_X1 U7746 ( .A1(n11836), .A2(n6749), .ZN(n6748) );
  NAND2_X1 U7747 ( .A1(n6809), .A2(n6522), .ZN(n6749) );
  NAND2_X1 U7748 ( .A1(n11667), .A2(n11666), .ZN(n11838) );
  NOR2_X1 U7749 ( .A1(n6431), .A2(n7017), .ZN(n7016) );
  OR2_X1 U7750 ( .A1(n10060), .A2(n6643), .ZN(n10000) );
  NOR2_X1 U7751 ( .A1(n6431), .A2(n9998), .ZN(n6643) );
  NOR2_X1 U7752 ( .A1(n12343), .A2(n12342), .ZN(n12345) );
  NOR2_X1 U7753 ( .A1(n12431), .A2(n6994), .ZN(n6993) );
  INV_X1 U7754 ( .A(n8663), .ZN(n6994) );
  OR2_X1 U7755 ( .A1(n12713), .A2(n12498), .ZN(n11769) );
  OR2_X1 U7756 ( .A1(n12539), .A2(n12511), .ZN(n11760) );
  NAND2_X1 U7757 ( .A1(n8737), .A2(n11743), .ZN(n8738) );
  INV_X1 U7758 ( .A(n6965), .ZN(n6964) );
  OAI21_X1 U7759 ( .B1(n8482), .B2(n6486), .A(n8499), .ZN(n6965) );
  INV_X1 U7760 ( .A(n11736), .ZN(n7192) );
  INV_X1 U7761 ( .A(n11741), .ZN(n7188) );
  NOR2_X1 U7762 ( .A1(n7066), .A2(n7065), .ZN(n7064) );
  NAND2_X1 U7763 ( .A1(n6616), .A2(n7071), .ZN(n7065) );
  NAND2_X1 U7764 ( .A1(n8677), .A2(n7072), .ZN(n7069) );
  NAND2_X1 U7765 ( .A1(n8247), .A2(n8246), .ZN(n8248) );
  NAND2_X1 U7766 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n10725), .ZN(n8246) );
  NOR2_X1 U7767 ( .A1(n7054), .A2(n12205), .ZN(n6732) );
  INV_X1 U7768 ( .A(n8244), .ZN(n7055) );
  NOR2_X1 U7769 ( .A1(P3_IR_REG_13__SCAN_IN), .A2(P3_IR_REG_4__SCAN_IN), .ZN(
        n8197) );
  XNOR2_X1 U7770 ( .A(n10177), .B(n7692), .ZN(n7594) );
  INV_X1 U7771 ( .A(n7080), .ZN(n7078) );
  INV_X1 U7772 ( .A(n6885), .ZN(n6879) );
  INV_X1 U7773 ( .A(n12927), .ZN(n7098) );
  NAND2_X1 U7774 ( .A1(n13174), .A2(n6948), .ZN(n6947) );
  INV_X1 U7775 ( .A(n13258), .ZN(n6948) );
  INV_X1 U7776 ( .A(n11123), .ZN(n7249) );
  NAND2_X1 U7777 ( .A1(n7113), .A2(n10157), .ZN(n7112) );
  NOR2_X1 U7778 ( .A1(n10240), .A2(n7114), .ZN(n7113) );
  INV_X1 U7779 ( .A(n10159), .ZN(n7114) );
  NAND2_X1 U7780 ( .A1(n7468), .A2(n6894), .ZN(n6893) );
  INV_X1 U7781 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n6894) );
  INV_X1 U7782 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n7493) );
  OR2_X1 U7783 ( .A1(n7562), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n7615) );
  NAND2_X2 U7784 ( .A1(n13449), .A2(n13444), .ZN(n6591) );
  AND2_X1 U7785 ( .A1(n6900), .A2(n13495), .ZN(n6899) );
  NAND2_X1 U7786 ( .A1(n13924), .A2(n11598), .ZN(n6900) );
  INV_X1 U7787 ( .A(n11598), .ZN(n6901) );
  NOR2_X1 U7788 ( .A1(n13961), .A2(n13352), .ZN(n7360) );
  NOR2_X1 U7789 ( .A1(n13952), .A2(n6909), .ZN(n6908) );
  INV_X1 U7790 ( .A(n7441), .ZN(n6909) );
  NOR2_X1 U7791 ( .A1(n13612), .A2(n6940), .ZN(n6939) );
  INV_X1 U7792 ( .A(n6941), .ZN(n6940) );
  INV_X1 U7793 ( .A(n7416), .ZN(n7415) );
  OAI21_X1 U7794 ( .B1(n7417), .B2(n6470), .A(n13485), .ZN(n7416) );
  INV_X1 U7795 ( .A(n7418), .ZN(n7417) );
  NAND2_X1 U7796 ( .A1(n10904), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10938) );
  XNOR2_X1 U7797 ( .A(n14115), .B(n13903), .ZN(n13495) );
  NAND2_X1 U7798 ( .A1(n11596), .A2(n11595), .ZN(n13988) );
  AOI21_X1 U7799 ( .B1(n6435), .B2(n7353), .A(n6545), .ZN(n7352) );
  INV_X1 U7800 ( .A(n11089), .ZN(n7353) );
  INV_X1 U7801 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9285) );
  NAND2_X1 U7802 ( .A1(n7875), .A2(n6481), .ZN(n7229) );
  NAND2_X1 U7803 ( .A1(n6931), .A2(n7831), .ZN(n6930) );
  INV_X1 U7804 ( .A(n7851), .ZN(n6931) );
  NOR2_X1 U7805 ( .A1(n7828), .A2(n6933), .ZN(n6932) );
  INV_X1 U7806 ( .A(n7812), .ZN(n6933) );
  BUF_X1 U7807 ( .A(n7228), .Z(n6708) );
  AOI21_X1 U7808 ( .B1(n7219), .B2(n7220), .A(n7217), .ZN(n7216) );
  INV_X1 U7809 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n9182) );
  INV_X1 U7810 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n9181) );
  OR2_X1 U7811 ( .A1(n7605), .A2(n7610), .ZN(n7604) );
  OR2_X1 U7812 ( .A1(n9232), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n9245) );
  NAND4_X1 U7813 ( .A1(n14401), .A2(n7475), .A3(P1_ADDR_REG_19__SCAN_IN), .A4(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n6936) );
  NAND4_X1 U7814 ( .A1(n7474), .A2(n12908), .A3(n7210), .A4(
        P3_ADDR_REG_19__SCAN_IN), .ZN(n6937) );
  INV_X1 U7815 ( .A(P2_RD_REG_SCAN_IN), .ZN(n7475) );
  INV_X1 U7816 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n6682) );
  INV_X1 U7817 ( .A(n7134), .ZN(n14260) );
  NAND2_X1 U7818 ( .A1(n14259), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n7135) );
  NOR2_X1 U7819 ( .A1(n6857), .A2(P1_ADDR_REG_4__SCAN_IN), .ZN(n6856) );
  INV_X1 U7820 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n14267) );
  NOR2_X1 U7821 ( .A1(n14275), .A2(n14274), .ZN(n14294) );
  NOR2_X1 U7822 ( .A1(n14315), .A2(n14273), .ZN(n14274) );
  NOR2_X1 U7823 ( .A1(n8883), .A2(n8882), .ZN(n7009) );
  NAND2_X1 U7824 ( .A1(n10528), .A2(n7010), .ZN(n10744) );
  AND2_X1 U7825 ( .A1(n8831), .A2(n8826), .ZN(n7010) );
  AOI22_X1 U7826 ( .A1(n8841), .A2(n8842), .B1(n8840), .B2(n12145), .ZN(n8843)
         );
  NAND2_X1 U7827 ( .A1(n8889), .A2(n12421), .ZN(n8890) );
  INV_X1 U7828 ( .A(n8210), .ZN(n11846) );
  OR2_X1 U7829 ( .A1(n12749), .A2(n8784), .ZN(n9203) );
  XNOR2_X1 U7830 ( .A(n10067), .B(n7017), .ZN(n10058) );
  NOR2_X1 U7831 ( .A1(n10061), .A2(n10062), .ZN(n10060) );
  INV_X1 U7832 ( .A(n9987), .ZN(n7032) );
  NAND2_X1 U7833 ( .A1(n10355), .A2(n10356), .ZN(n10387) );
  OR2_X1 U7834 ( .A1(n10771), .A2(n10772), .ZN(n7030) );
  AND2_X1 U7835 ( .A1(n7030), .A2(n7029), .ZN(n12313) );
  INV_X1 U7836 ( .A(n10773), .ZN(n7029) );
  NOR2_X1 U7837 ( .A1(n12313), .A2(n7028), .ZN(n12315) );
  AND2_X1 U7838 ( .A1(n12314), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7028) );
  OR2_X1 U7839 ( .A1(n15019), .A2(n15018), .ZN(n15021) );
  NAND2_X1 U7840 ( .A1(n8664), .A2(n6993), .ZN(n12435) );
  NAND2_X1 U7841 ( .A1(n6958), .A2(n8637), .ZN(n12454) );
  INV_X1 U7842 ( .A(n12137), .ZN(n12456) );
  NAND2_X1 U7843 ( .A1(n8745), .A2(n11779), .ZN(n12457) );
  AND4_X1 U7844 ( .A1(n8621), .A2(n8620), .A3(n8619), .A4(n8618), .ZN(n12470)
         );
  OAI21_X1 U7845 ( .B1(n12520), .B2(n11770), .A(n11769), .ZN(n12488) );
  OR2_X1 U7846 ( .A1(n12488), .A2(n12494), .ZN(n12490) );
  AOI21_X1 U7847 ( .B1(n12576), .B2(n7180), .A(n7179), .ZN(n7178) );
  AND2_X1 U7848 ( .A1(n8525), .A2(n8739), .ZN(n12559) );
  AND4_X1 U7849 ( .A1(n8512), .A2(n8511), .A3(n8510), .A4(n8509), .ZN(n12597)
         );
  NAND2_X1 U7850 ( .A1(n6959), .A2(n6538), .ZN(n11382) );
  NAND2_X1 U7851 ( .A1(n11308), .A2(n8456), .ZN(n6959) );
  NAND2_X1 U7852 ( .A1(n11388), .A2(n11827), .ZN(n11387) );
  NOR2_X1 U7853 ( .A1(n7185), .A2(n7184), .ZN(n7183) );
  INV_X1 U7854 ( .A(n11731), .ZN(n7184) );
  NOR2_X1 U7855 ( .A1(n8732), .A2(n7186), .ZN(n7185) );
  INV_X1 U7856 ( .A(n11729), .ZN(n7186) );
  CLKBUF_X1 U7857 ( .A(n8733), .Z(n6684) );
  AND4_X1 U7858 ( .A1(n8410), .A2(n8409), .A3(n8408), .A4(n8407), .ZN(n11398)
         );
  INV_X1 U7859 ( .A(n6980), .ZN(n11057) );
  AOI21_X1 U7860 ( .B1(n6978), .B2(n11817), .A(n6551), .ZN(n6976) );
  INV_X1 U7861 ( .A(n6978), .ZN(n6977) );
  NOR2_X1 U7862 ( .A1(n11822), .A2(n6979), .ZN(n6978) );
  INV_X1 U7863 ( .A(n8338), .ZN(n6979) );
  INV_X1 U7864 ( .A(n11698), .ZN(n11822) );
  NAND2_X1 U7865 ( .A1(n10729), .A2(n11696), .ZN(n10728) );
  AND4_X1 U7866 ( .A1(n8326), .A2(n8325), .A3(n8324), .A4(n8323), .ZN(n10685)
         );
  NAND2_X1 U7867 ( .A1(n8287), .A2(n8286), .ZN(n15083) );
  INV_X1 U7868 ( .A(n12571), .ZN(n15104) );
  INV_X1 U7869 ( .A(n12569), .ZN(n15106) );
  NAND2_X1 U7870 ( .A1(n12387), .A2(n12386), .ZN(n12385) );
  AND2_X1 U7871 ( .A1(n11848), .A2(n11682), .ZN(n11804) );
  AOI21_X1 U7872 ( .B1(n12731), .B2(n11663), .A(n11652), .ZN(n14465) );
  NOR2_X1 U7873 ( .A1(n8310), .A2(n12727), .ZN(n11652) );
  AND2_X1 U7874 ( .A1(n14458), .A2(n14457), .ZN(n14469) );
  NAND2_X1 U7875 ( .A1(n8260), .A2(n8259), .ZN(n8703) );
  NAND2_X1 U7876 ( .A1(n8615), .A2(n8614), .ZN(n11776) );
  INV_X1 U7877 ( .A(n14482), .ZN(n15139) );
  NAND2_X1 U7878 ( .A1(n8285), .A2(n6537), .ZN(n8726) );
  NOR2_X1 U7879 ( .A1(n7069), .A2(n8256), .ZN(n7066) );
  NAND2_X1 U7880 ( .A1(n8756), .A2(n6497), .ZN(n8767) );
  NAND2_X1 U7881 ( .A1(n14251), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n7072) );
  NAND2_X1 U7882 ( .A1(n8255), .A2(n8254), .ZN(n8666) );
  NAND2_X1 U7883 ( .A1(n8765), .A2(n7013), .ZN(n7012) );
  XNOR2_X1 U7884 ( .A(n8253), .B(n7046), .ZN(n8651) );
  NAND2_X1 U7885 ( .A1(n8251), .A2(n6751), .ZN(n8626) );
  NAND2_X1 U7886 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n6752), .ZN(n6751) );
  INV_X1 U7887 ( .A(n6797), .ZN(n8717) );
  NAND2_X1 U7888 ( .A1(n7038), .A2(n7036), .ZN(n8583) );
  NAND2_X1 U7889 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n7037), .ZN(n7036) );
  NAND2_X1 U7890 ( .A1(n8569), .A2(n8567), .ZN(n7038) );
  NAND2_X1 U7891 ( .A1(n8245), .A2(n6722), .ZN(n8551) );
  NAND2_X1 U7892 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n6723), .ZN(n6722) );
  NAND2_X1 U7893 ( .A1(n6733), .A2(n8243), .ZN(n8502) );
  NAND2_X1 U7894 ( .A1(n8483), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6733) );
  XNOR2_X1 U7895 ( .A(n8242), .B(P2_DATAO_REG_13__SCAN_IN), .ZN(n8483) );
  AOI21_X1 U7896 ( .B1(n7043), .B2(n6476), .A(n6560), .ZN(n6736) );
  XNOR2_X1 U7897 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n8411) );
  NAND2_X1 U7898 ( .A1(n8239), .A2(n8238), .ZN(n8412) );
  XNOR2_X1 U7899 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n8428) );
  INV_X1 U7900 ( .A(n8236), .ZN(n6729) );
  INV_X1 U7901 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n8396) );
  OAI21_X1 U7902 ( .B1(n8366), .B2(n8234), .A(n8235), .ZN(n8382) );
  AND2_X1 U7903 ( .A1(n9230), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8234) );
  OR2_X1 U7904 ( .A1(n8352), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n8472) );
  AOI21_X1 U7905 ( .B1(n8311), .B2(n7057), .A(n6557), .ZN(n7056) );
  INV_X1 U7906 ( .A(n9769), .ZN(n7161) );
  OR2_X1 U7907 ( .A1(n7819), .A2(n7818), .ZN(n7837) );
  INV_X1 U7908 ( .A(n7948), .ZN(n7946) );
  AND2_X1 U7909 ( .A1(n7935), .A2(n7151), .ZN(n7150) );
  NAND2_X1 U7910 ( .A1(n7153), .A2(n7152), .ZN(n7151) );
  NAND2_X1 U7911 ( .A1(n12817), .A2(n6533), .ZN(n12784) );
  INV_X1 U7912 ( .A(n12861), .ZN(n10736) );
  NAND2_X1 U7913 ( .A1(n12794), .A2(n8080), .ZN(n12841) );
  AOI211_X1 U7914 ( .C1(n9152), .C2(n9151), .A(n13001), .B(n9158), .ZN(n9153)
         );
  AND2_X1 U7915 ( .A1(n8015), .A2(n8014), .ZN(n12974) );
  AND2_X1 U7916 ( .A1(n7888), .A2(n7887), .ZN(n12958) );
  AND4_X1 U7917 ( .A1(n7653), .A2(n7652), .A3(n7651), .A4(n7650), .ZN(n10242)
         );
  NOR2_X2 U7918 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n7544) );
  NAND2_X1 U7919 ( .A1(n14752), .A2(n14753), .ZN(n14751) );
  NOR2_X1 U7920 ( .A1(n9420), .A2(n6846), .ZN(n9433) );
  AND2_X1 U7921 ( .A1(n9390), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6846) );
  OR2_X1 U7922 ( .A1(n7085), .A2(n6511), .ZN(n7080) );
  OR2_X1 U7923 ( .A1(n7082), .A2(n6511), .ZN(n7079) );
  AOI21_X1 U7924 ( .B1(n7084), .B2(n7083), .A(n6555), .ZN(n7082) );
  INV_X1 U7925 ( .A(n6493), .ZN(n7083) );
  NAND2_X1 U7926 ( .A1(n13052), .A2(n12978), .ZN(n13038) );
  AND2_X1 U7927 ( .A1(n13055), .A2(n13039), .ZN(n13040) );
  NAND2_X1 U7928 ( .A1(n13214), .A2(n12977), .ZN(n7090) );
  NAND2_X1 U7929 ( .A1(n6488), .A2(n12976), .ZN(n13052) );
  AND2_X1 U7930 ( .A1(n13054), .A2(n13077), .ZN(n13055) );
  NAND2_X1 U7931 ( .A1(n6621), .A2(n13066), .ZN(n13075) );
  INV_X1 U7932 ( .A(n7109), .ZN(n13069) );
  INV_X1 U7933 ( .A(n7106), .ZN(n7105) );
  NAND2_X1 U7934 ( .A1(n13110), .A2(n12934), .ZN(n7108) );
  NAND2_X1 U7935 ( .A1(n7108), .A2(n7106), .ZN(n13089) );
  AND2_X1 U7936 ( .A1(n12932), .A2(n12931), .ZN(n13124) );
  OR2_X1 U7937 ( .A1(n13131), .A2(n12929), .ZN(n12932) );
  NOR2_X1 U7938 ( .A1(n12965), .A2(n6888), .ZN(n6887) );
  INV_X1 U7939 ( .A(n12962), .ZN(n6888) );
  AND2_X1 U7940 ( .A1(n12933), .A2(n9133), .ZN(n13125) );
  NOR2_X1 U7941 ( .A1(n11368), .A2(n13258), .ZN(n13168) );
  NOR2_X1 U7942 ( .A1(n11368), .A2(n6947), .ZN(n13171) );
  NAND2_X1 U7943 ( .A1(n7102), .A2(n7101), .ZN(n13162) );
  INV_X1 U7944 ( .A(n13165), .ZN(n7101) );
  INV_X1 U7945 ( .A(n13164), .ZN(n7102) );
  INV_X1 U7946 ( .A(n11355), .ZN(n7242) );
  NAND2_X1 U7947 ( .A1(n7245), .A2(n7244), .ZN(n7243) );
  INV_X1 U7948 ( .A(n11354), .ZN(n7245) );
  INV_X1 U7949 ( .A(n7248), .ZN(n6875) );
  AOI21_X1 U7950 ( .B1(n7248), .B2(n6874), .A(n6873), .ZN(n6872) );
  INV_X1 U7951 ( .A(n11120), .ZN(n6874) );
  INV_X1 U7952 ( .A(n7246), .ZN(n6873) );
  AOI21_X1 U7953 ( .B1(n7248), .B2(n7247), .A(n6531), .ZN(n7246) );
  NAND2_X1 U7954 ( .A1(n11114), .A2(n11113), .ZN(n11133) );
  NAND2_X1 U7955 ( .A1(n11121), .A2(n11120), .ZN(n14504) );
  AND2_X1 U7956 ( .A1(n10878), .A2(n10879), .ZN(n7120) );
  OR2_X1 U7957 ( .A1(n10579), .A2(n10585), .ZN(n10880) );
  NAND2_X1 U7958 ( .A1(n10472), .A2(n10471), .ZN(n10577) );
  AND2_X1 U7959 ( .A1(n10252), .A2(n10470), .ZN(n10479) );
  NAND2_X1 U7960 ( .A1(n9920), .A2(n9919), .ZN(n10540) );
  XNOR2_X1 U7961 ( .A(n8937), .B(n11625), .ZN(n10539) );
  XNOR2_X1 U7962 ( .A(n11202), .B(n6485), .ZN(n9916) );
  NAND2_X1 U7963 ( .A1(n9938), .A2(n9937), .ZN(n14814) );
  XNOR2_X1 U7964 ( .A(n11644), .B(n12870), .ZN(n11637) );
  INV_X1 U7965 ( .A(n13155), .ZN(n13248) );
  NAND2_X1 U7966 ( .A1(n7754), .A2(n7753), .ZN(n14942) );
  INV_X1 U7967 ( .A(n14943), .ZN(n14933) );
  AND2_X1 U7968 ( .A1(n8141), .A2(n8149), .ZN(n14845) );
  AND2_X1 U7969 ( .A1(n8134), .A2(n6483), .ZN(n8148) );
  XNOR2_X1 U7970 ( .A(n8153), .B(n8152), .ZN(n9377) );
  INV_X1 U7971 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8152) );
  INV_X1 U7972 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n7488) );
  INV_X1 U7973 ( .A(n9288), .ZN(n9543) );
  INV_X1 U7974 ( .A(n13934), .ZN(n13310) );
  NAND2_X1 U7975 ( .A1(n11859), .A2(n11858), .ZN(n14555) );
  OR2_X1 U7976 ( .A1(n10287), .A2(n10286), .ZN(n10496) );
  NOR2_X1 U7977 ( .A1(n11229), .A2(n11228), .ZN(n11237) );
  INV_X1 U7978 ( .A(n10715), .ZN(n7402) );
  NAND2_X1 U7979 ( .A1(n10711), .A2(n6783), .ZN(n6782) );
  AND2_X1 U7980 ( .A1(n7403), .A2(n10710), .ZN(n6783) );
  NOR2_X1 U7981 ( .A1(n11518), .A2(n13325), .ZN(n11530) );
  OAI21_X1 U7982 ( .B1(n13386), .B2(n7395), .A(n7393), .ZN(n13399) );
  AOI21_X1 U7983 ( .B1(n7396), .B2(n7394), .A(n6519), .ZN(n7393) );
  INV_X1 U7984 ( .A(n7396), .ZN(n7395) );
  AND2_X1 U7985 ( .A1(n11432), .A2(n11431), .ZN(n13628) );
  NAND2_X1 U7986 ( .A1(n13861), .A2(n13860), .ZN(n13900) );
  NAND2_X1 U7987 ( .A1(n13931), .A2(n7443), .ZN(n13916) );
  NAND2_X1 U7988 ( .A1(n13933), .A2(n13932), .ZN(n13931) );
  AND2_X1 U7989 ( .A1(n7423), .A2(n11538), .ZN(n7422) );
  OR2_X1 U7990 ( .A1(n13612), .A2(n14537), .ZN(n13616) );
  AND2_X1 U7991 ( .A1(n11236), .A2(n13610), .ZN(n6913) );
  AND4_X1 U7992 ( .A1(n11086), .A2(n11085), .A3(n11084), .A4(n11083), .ZN(
        n11885) );
  NAND2_X1 U7993 ( .A1(n14588), .A2(n13343), .ZN(n7418) );
  NAND2_X1 U7994 ( .A1(n10911), .A2(n10910), .ZN(n10934) );
  NAND2_X1 U7995 ( .A1(n10840), .A2(n7367), .ZN(n10911) );
  NOR2_X1 U7996 ( .A1(n10846), .A2(n7368), .ZN(n7367) );
  INV_X1 U7997 ( .A(n10839), .ZN(n7368) );
  NAND2_X1 U7998 ( .A1(n10510), .A2(n7369), .ZN(n10840) );
  AND2_X1 U7999 ( .A1(n13479), .A2(n10509), .ZN(n7369) );
  AOI21_X1 U8000 ( .B1(n7357), .B2(n7359), .A(n6509), .ZN(n7355) );
  NAND2_X1 U8001 ( .A1(n10550), .A2(n10723), .ZN(n10567) );
  OAI21_X1 U8002 ( .B1(n10260), .B2(n13474), .A(n10266), .ZN(n7408) );
  NAND2_X1 U8003 ( .A1(n10281), .A2(n10280), .ZN(n10555) );
  INV_X1 U8004 ( .A(n13474), .ZN(n10554) );
  NAND2_X1 U8005 ( .A1(n10218), .A2(n10217), .ZN(n10261) );
  AOI21_X1 U8006 ( .B1(n7411), .B2(n13539), .A(n6534), .ZN(n7409) );
  OR2_X1 U8007 ( .A1(n13457), .A2(n6468), .ZN(n14020) );
  OR2_X1 U8008 ( .A1(n13457), .A2(n9525), .ZN(n14060) );
  INV_X1 U8009 ( .A(n14060), .ZN(n14083) );
  NAND2_X1 U8010 ( .A1(n9741), .A2(n9740), .ZN(n9831) );
  OR2_X1 U8011 ( .A1(n6426), .A2(n14618), .ZN(n9512) );
  INV_X1 U8012 ( .A(n13978), .ZN(n14142) );
  INV_X1 U8013 ( .A(n14028), .ZN(n14157) );
  NAND2_X1 U8014 ( .A1(n11517), .A2(n11516), .ZN(n14043) );
  NAND2_X1 U8015 ( .A1(n11509), .A2(n11508), .ZN(n14175) );
  AND2_X1 U8016 ( .A1(n13957), .A2(n14716), .ZN(n14192) );
  AND2_X1 U8017 ( .A1(n9786), .A2(n9536), .ZN(n14587) );
  NAND2_X1 U8018 ( .A1(n13441), .A2(n9509), .ZN(n14183) );
  AND3_X1 U8019 ( .A1(n9194), .A2(n6566), .A3(n9289), .ZN(n7436) );
  XNOR2_X1 U8020 ( .A(n9068), .B(n9070), .ZN(n13445) );
  NAND2_X1 U8021 ( .A1(n8088), .A2(n8087), .ZN(n8159) );
  INV_X1 U8022 ( .A(n9357), .ZN(n6630) );
  INV_X1 U8023 ( .A(n8001), .ZN(n7225) );
  AND2_X1 U8024 ( .A1(n12257), .A2(n7294), .ZN(n7293) );
  INV_X1 U8025 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U8026 ( .A1(n7875), .A2(n7874), .ZN(n7894) );
  NOR2_X1 U8027 ( .A1(n7612), .A2(n6707), .ZN(n6706) );
  INV_X1 U8028 ( .A(n7610), .ZN(n6707) );
  AND2_X1 U8029 ( .A1(n7611), .A2(n7583), .ZN(n9836) );
  OR2_X1 U8030 ( .A1(n7582), .A2(n7606), .ZN(n7583) );
  NAND2_X1 U8031 ( .A1(n6631), .A2(n14307), .ZN(n14310) );
  NAND2_X1 U8032 ( .A1(n14318), .A2(n14317), .ZN(n14319) );
  OAI22_X1 U8033 ( .A1(P1_ADDR_REG_13__SCAN_IN), .A2(n15017), .B1(n14289), 
        .B2(n14288), .ZN(n14345) );
  NOR2_X1 U8034 ( .A1(n6475), .A2(n12134), .ZN(n6785) );
  NAND2_X1 U8035 ( .A1(n6788), .A2(n6790), .ZN(n6787) );
  NAND2_X1 U8036 ( .A1(n6795), .A2(n12116), .ZN(n6790) );
  INV_X1 U8037 ( .A(n7450), .ZN(n7011) );
  INV_X1 U8038 ( .A(n6999), .ZN(n6998) );
  OAI21_X1 U8039 ( .B1(n7001), .B2(n6502), .A(n7000), .ZN(n6999) );
  NAND2_X1 U8040 ( .A1(n7003), .A2(n7002), .ZN(n7001) );
  INV_X1 U8041 ( .A(n12141), .ZN(n12596) );
  AND3_X1 U8042 ( .A1(n8454), .A2(n8453), .A3(n8452), .ZN(n11316) );
  AND3_X1 U8043 ( .A1(n8300), .A2(n8299), .A3(n8298), .ZN(n10434) );
  OR2_X1 U8044 ( .A1(n8310), .A2(SI_2_), .ZN(n8299) );
  NAND2_X1 U8045 ( .A1(n8680), .A2(n8679), .ZN(n12422) );
  NAND2_X1 U8046 ( .A1(n8919), .A2(n15114), .ZN(n12132) );
  INV_X1 U8047 ( .A(n12510), .ZN(n12139) );
  INV_X1 U8048 ( .A(n10685), .ZN(n11704) );
  XNOR2_X1 U8049 ( .A(n12315), .B(n12333), .ZN(n14972) );
  NAND2_X1 U8050 ( .A1(n9991), .A2(n9990), .ZN(n15050) );
  INV_X1 U8051 ( .A(n12373), .ZN(n6703) );
  NOR2_X1 U8052 ( .A1(n12370), .A2(n6705), .ZN(n6704) );
  OAI22_X1 U8053 ( .A1(n12362), .A2(n12361), .B1(n12371), .B2(n12664), .ZN(
        n12364) );
  AOI211_X1 U8054 ( .C1(n15035), .C2(n12375), .A(n6642), .B(n6608), .ZN(n6641)
         );
  INV_X1 U8055 ( .A(n12365), .ZN(n6642) );
  NOR2_X1 U8056 ( .A1(n6989), .A2(n6988), .ZN(n6987) );
  NOR2_X1 U8057 ( .A1(n11665), .A2(n14456), .ZN(n6988) );
  NOR2_X1 U8058 ( .A1(n12000), .A2(n15106), .ZN(n6989) );
  NAND2_X1 U8059 ( .A1(n12406), .A2(n6646), .ZN(n12623) );
  INV_X1 U8060 ( .A(n6647), .ZN(n6646) );
  OAI21_X1 U8061 ( .B1(n12408), .B2(n15093), .A(n12407), .ZN(n6647) );
  NAND2_X1 U8062 ( .A1(n6750), .A2(n8693), .ZN(n12412) );
  NAND2_X1 U8063 ( .A1(n12740), .A2(n11663), .ZN(n6750) );
  NAND2_X1 U8064 ( .A1(n8599), .A2(n8598), .ZN(n12505) );
  AND3_X1 U8065 ( .A1(n8480), .A2(n8479), .A3(n8478), .ZN(n14477) );
  AND3_X1 U8066 ( .A1(n8356), .A2(n8355), .A3(n8354), .ZN(n15072) );
  OR2_X1 U8067 ( .A1(n8310), .A2(SI_5_), .ZN(n8355) );
  INV_X1 U8068 ( .A(n8703), .ZN(n12686) );
  OAI21_X1 U8069 ( .B1(n12619), .B2(n15139), .A(n12620), .ZN(n12683) );
  AND2_X1 U8070 ( .A1(n8641), .A2(n8640), .ZN(n12700) );
  OR2_X1 U8071 ( .A1(n15144), .A2(n15138), .ZN(n12724) );
  XNOR2_X1 U8072 ( .A(n8214), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11848) );
  OAI21_X1 U8073 ( .B1(n8717), .B2(P3_IR_REG_21__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8214) );
  NAND2_X1 U8074 ( .A1(n8587), .A2(n8715), .ZN(n12363) );
  NAND2_X1 U8075 ( .A1(n6663), .A2(n9085), .ZN(n7734) );
  INV_X1 U8076 ( .A(n10821), .ZN(n6663) );
  INV_X1 U8077 ( .A(n10470), .ZN(n14916) );
  AND2_X1 U8078 ( .A1(n11015), .A2(n7782), .ZN(n6689) );
  NAND2_X1 U8079 ( .A1(n11282), .A2(n7847), .ZN(n11461) );
  NAND2_X1 U8080 ( .A1(n7720), .A2(n7719), .ZN(n10655) );
  INV_X1 U8081 ( .A(n10648), .ZN(n6715) );
  INV_X1 U8082 ( .A(n13122), .ZN(n13237) );
  AND2_X1 U8083 ( .A1(n8180), .A2(n8155), .ZN(n14494) );
  INV_X1 U8084 ( .A(n12983), .ZN(n12941) );
  INV_X1 U8085 ( .A(n11122), .ZN(n12859) );
  AND3_X1 U8086 ( .A1(n7528), .A2(n7529), .A3(n7527), .ZN(n7531) );
  OAI21_X1 U8087 ( .B1(n10314), .B2(n10313), .A(n10312), .ZN(n10695) );
  INV_X1 U8088 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n12908) );
  NOR2_X1 U8089 ( .A1(n12898), .A2(n12897), .ZN(n12899) );
  NOR2_X1 U8090 ( .A1(n12893), .A2(n12892), .ZN(n12894) );
  NAND2_X2 U8091 ( .A1(n8163), .A2(n8162), .ZN(n13190) );
  OR3_X1 U8092 ( .A1(n13077), .A2(n13076), .A3(n13169), .ZN(n13219) );
  OAI21_X1 U8093 ( .B1(n12963), .B2(n6885), .A(n6881), .ZN(n13101) );
  AND2_X1 U8094 ( .A1(n7817), .A2(n7816), .ZN(n14520) );
  AND2_X1 U8095 ( .A1(n7620), .A2(n7619), .ZN(n14895) );
  NAND2_X1 U8096 ( .A1(n8164), .A2(n14854), .ZN(n14819) );
  AND2_X2 U8097 ( .A1(n11158), .A2(n11149), .ZN(n14970) );
  AND2_X1 U8098 ( .A1(n13186), .A2(n6895), .ZN(n6672) );
  OR2_X1 U8099 ( .A1(n13188), .A2(n13261), .ZN(n6895) );
  INV_X1 U8100 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7509) );
  NAND2_X1 U8101 ( .A1(n7379), .A2(n7377), .ZN(n13322) );
  AOI21_X1 U8102 ( .B1(n7380), .B2(n7381), .A(n7378), .ZN(n7377) );
  INV_X1 U8103 ( .A(n13323), .ZN(n7378) );
  INV_X1 U8104 ( .A(n7386), .ZN(n11984) );
  OAI21_X1 U8105 ( .B1(n13349), .B2(n6563), .A(n7387), .ZN(n7386) );
  AOI21_X1 U8106 ( .B1(n7388), .B2(n13307), .A(n6565), .ZN(n7387) );
  NAND2_X1 U8107 ( .A1(n6487), .A2(n9630), .ZN(n9679) );
  INV_X1 U8108 ( .A(n13338), .ZN(n6778) );
  NAND2_X1 U8109 ( .A1(n7372), .A2(n7371), .ZN(n13339) );
  NAND2_X1 U8110 ( .A1(n6500), .A2(n6764), .ZN(n10327) );
  NAND2_X1 U8111 ( .A1(n13392), .A2(n13391), .ZN(n14540) );
  NAND2_X1 U8112 ( .A1(n10628), .A2(n10627), .ZN(n10711) );
  NAND2_X1 U8113 ( .A1(n6489), .A2(n7212), .ZN(n7211) );
  INV_X1 U8114 ( .A(n13722), .ZN(n7212) );
  INV_X1 U8115 ( .A(n7214), .ZN(n7213) );
  OAI21_X1 U8116 ( .B1(n13729), .B2(n13728), .A(n13726), .ZN(n7214) );
  AND2_X1 U8117 ( .A1(n13513), .A2(n13514), .ZN(n13727) );
  OR2_X1 U8118 ( .A1(n6426), .A2(n9633), .ZN(n9636) );
  INV_X1 U8119 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n7474) );
  NAND2_X1 U8120 ( .A1(n6680), .A2(n6678), .ZN(n6677) );
  NAND2_X1 U8121 ( .A1(n13853), .A2(n14640), .ZN(n6680) );
  NOR2_X1 U8122 ( .A1(n13852), .A2(n6679), .ZN(n6678) );
  XNOR2_X1 U8123 ( .A(n13875), .B(n13880), .ZN(n14106) );
  NAND2_X1 U8124 ( .A1(n11565), .A2(n11564), .ZN(n13968) );
  NAND2_X1 U8125 ( .A1(n10932), .A2(n10931), .ZN(n13601) );
  NAND2_X1 U8126 ( .A1(n10495), .A2(n10494), .ZN(n13576) );
  AND2_X1 U8127 ( .A1(n9196), .A2(n9294), .ZN(n11448) );
  INV_X1 U8128 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14300) );
  AOI21_X1 U8129 ( .B1(n14370), .B2(n14304), .A(n14367), .ZN(n15160) );
  AOI21_X1 U8130 ( .B1(n14344), .B2(n7147), .A(n7144), .ZN(n14611) );
  NOR2_X1 U8131 ( .A1(n7149), .A2(n7146), .ZN(n7145) );
  OR2_X1 U8132 ( .A1(n14614), .A2(P2_ADDR_REG_16__SCAN_IN), .ZN(n7123) );
  INV_X1 U8133 ( .A(n14359), .ZN(n7122) );
  OR2_X1 U8134 ( .A1(n14353), .A2(n6865), .ZN(n6864) );
  AND2_X1 U8135 ( .A1(n14393), .A2(n7129), .ZN(n7127) );
  NAND2_X1 U8136 ( .A1(n11644), .A2(n9091), .ZN(n8924) );
  NAND2_X1 U8137 ( .A1(n7291), .A2(n13554), .ZN(n7290) );
  NAND2_X1 U8138 ( .A1(n8947), .A2(n8946), .ZN(n7296) );
  INV_X1 U8139 ( .A(n13573), .ZN(n7286) );
  NOR2_X1 U8140 ( .A1(n7288), .A2(n13573), .ZN(n7287) );
  NAND2_X1 U8141 ( .A1(n7333), .A2(n6536), .ZN(n7332) );
  AND2_X1 U8142 ( .A1(n7329), .A2(n7337), .ZN(n7328) );
  NAND2_X1 U8143 ( .A1(n7279), .A2(n13602), .ZN(n7278) );
  INV_X1 U8144 ( .A(n13603), .ZN(n7279) );
  NAND2_X1 U8145 ( .A1(n6651), .A2(n6652), .ZN(n8993) );
  NAND2_X1 U8146 ( .A1(n8989), .A2(n8988), .ZN(n6652) );
  AND2_X1 U8147 ( .A1(n13651), .A2(n6572), .ZN(n6718) );
  NAND2_X1 U8148 ( .A1(n13663), .A2(n13664), .ZN(n7276) );
  AOI21_X1 U8149 ( .B1(n6830), .B2(n6829), .A(n11698), .ZN(n11706) );
  NOR2_X1 U8150 ( .A1(n6521), .A2(n11696), .ZN(n6829) );
  NAND2_X1 U8151 ( .A1(n6832), .A2(n6831), .ZN(n6830) );
  OAI21_X1 U8152 ( .B1(n9002), .B2(n9001), .A(n6562), .ZN(n7341) );
  INV_X1 U8153 ( .A(n7275), .ZN(n7272) );
  INV_X1 U8154 ( .A(n13667), .ZN(n7273) );
  AOI21_X1 U8155 ( .B1(n6835), .B2(n6834), .A(n6504), .ZN(n11726) );
  NOR2_X1 U8156 ( .A1(n11719), .A2(n11718), .ZN(n6834) );
  OR2_X1 U8157 ( .A1(n13671), .A2(n13672), .ZN(n13673) );
  NAND2_X1 U8158 ( .A1(n7284), .A2(n13676), .ZN(n7283) );
  INV_X1 U8159 ( .A(n13675), .ZN(n7284) );
  AOI21_X1 U8160 ( .B1(n9020), .B2(n7319), .A(n7318), .ZN(n7317) );
  AOI21_X1 U8161 ( .B1(n6469), .B2(n7309), .A(n7303), .ZN(n7302) );
  AND2_X1 U8162 ( .A1(n7305), .A2(n7308), .ZN(n7303) );
  NAND2_X1 U8163 ( .A1(n6619), .A2(n6618), .ZN(n13681) );
  INV_X1 U8164 ( .A(n13679), .ZN(n6618) );
  NAND2_X1 U8165 ( .A1(n6826), .A2(n6825), .ZN(n6824) );
  NOR2_X1 U8166 ( .A1(n12494), .A2(n11772), .ZN(n6825) );
  NAND2_X1 U8167 ( .A1(n6828), .A2(n6827), .ZN(n6826) );
  NAND2_X1 U8168 ( .A1(n6556), .A2(n6822), .ZN(n6821) );
  INV_X1 U8169 ( .A(n12467), .ZN(n6822) );
  INV_X1 U8170 ( .A(n9037), .ZN(n7327) );
  NAND2_X1 U8171 ( .A1(n7268), .A2(n7266), .ZN(n7264) );
  NAND2_X1 U8172 ( .A1(n7267), .A2(n13691), .ZN(n7266) );
  INV_X1 U8173 ( .A(n13692), .ZN(n7267) );
  NAND2_X1 U8174 ( .A1(n6803), .A2(n6802), .ZN(n6808) );
  OAI21_X1 U8175 ( .B1(n6814), .B2(n6811), .A(n6813), .ZN(n6800) );
  AND2_X1 U8176 ( .A1(n11835), .A2(n11804), .ZN(n6807) );
  NOR2_X1 U8177 ( .A1(n12386), .A2(n11800), .ZN(n11835) );
  AND2_X1 U8178 ( .A1(n12670), .A2(n12070), .ZN(n11755) );
  NOR2_X1 U8179 ( .A1(P3_IR_REG_22__SCAN_IN), .A2(P3_IR_REG_21__SCAN_IN), .ZN(
        n8202) );
  NAND2_X1 U8180 ( .A1(n7197), .A2(n8200), .ZN(n7196) );
  INV_X1 U8181 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n8200) );
  INV_X1 U8182 ( .A(n7198), .ZN(n7197) );
  NOR2_X1 U8183 ( .A1(P3_IR_REG_12__SCAN_IN), .A2(P3_IR_REG_5__SCAN_IN), .ZN(
        n8196) );
  NAND2_X1 U8184 ( .A1(n13183), .A2(n12948), .ZN(n6713) );
  INV_X1 U8185 ( .A(n7916), .ZN(n7918) );
  INV_X1 U8186 ( .A(n7787), .ZN(n7217) );
  OAI21_X1 U8187 ( .B1(n9212), .B2(n6710), .A(n6709), .ZN(n7602) );
  NAND2_X1 U8188 ( .A1(n9212), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n6709) );
  OAI21_X1 U8189 ( .B1(n9212), .B2(n6693), .A(n6692), .ZN(n7580) );
  NAND2_X1 U8190 ( .A1(n9212), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n6692) );
  INV_X1 U8191 ( .A(P1_RD_REG_SCAN_IN), .ZN(n7210) );
  INV_X1 U8192 ( .A(n6859), .ZN(n6857) );
  INV_X1 U8193 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14277) );
  OAI21_X1 U8194 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14279), .A(n14278), .ZN(
        n14280) );
  OR2_X1 U8195 ( .A1(n8616), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U8196 ( .A1(n12078), .A2(n12137), .ZN(n7008) );
  NAND2_X1 U8197 ( .A1(n11837), .A2(n14460), .ZN(n11670) );
  NAND2_X1 U8198 ( .A1(n10099), .A2(n10002), .ZN(n10004) );
  NAND2_X1 U8199 ( .A1(n10667), .A2(n10668), .ZN(n10762) );
  NAND2_X1 U8200 ( .A1(n12331), .A2(n6595), .ZN(n12334) );
  NAND2_X1 U8201 ( .A1(n14425), .A2(n6639), .ZN(n12348) );
  NAND2_X1 U8202 ( .A1(n12322), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6639) );
  AOI21_X1 U8203 ( .B1(n7203), .B2(n11803), .A(n11802), .ZN(n7200) );
  INV_X1 U8204 ( .A(n6991), .ZN(n6990) );
  NAND2_X1 U8205 ( .A1(n12403), .A2(n7204), .ZN(n7203) );
  NAND2_X1 U8206 ( .A1(n11798), .A2(n11796), .ZN(n7204) );
  AND2_X1 U8207 ( .A1(n6975), .A2(n6969), .ZN(n6968) );
  NAND2_X1 U8208 ( .A1(n6972), .A2(n6970), .ZN(n6969) );
  AND2_X1 U8209 ( .A1(n8610), .A2(n12494), .ZN(n6975) );
  INV_X1 U8210 ( .A(n6972), .ZN(n6971) );
  NAND2_X1 U8211 ( .A1(n7178), .A2(n11829), .ZN(n7177) );
  NAND2_X1 U8212 ( .A1(n12146), .A2(n11180), .ZN(n11715) );
  NAND2_X1 U8213 ( .A1(n9203), .A2(n9329), .ZN(n9971) );
  NAND2_X1 U8214 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13297), .ZN(n7071) );
  INV_X1 U8215 ( .A(P3_IR_REG_26__SCAN_IN), .ZN(n8205) );
  AND2_X1 U8216 ( .A1(n7013), .A2(n8204), .ZN(n7209) );
  INV_X1 U8217 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n8204) );
  AND2_X1 U8218 ( .A1(n7048), .A2(n7047), .ZN(n8253) );
  NAND2_X1 U8219 ( .A1(n11297), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7047) );
  NAND2_X1 U8220 ( .A1(n7050), .A2(n7049), .ZN(n7048) );
  INV_X1 U8221 ( .A(n8638), .ZN(n7049) );
  NOR2_X1 U8222 ( .A1(n6716), .A2(n7196), .ZN(n7193) );
  NAND2_X1 U8223 ( .A1(n8199), .A2(n7199), .ZN(n7198) );
  INV_X1 U8224 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n8199) );
  INV_X1 U8225 ( .A(n8238), .ZN(n7041) );
  AOI21_X1 U8226 ( .B1(n6730), .B2(n8236), .A(n6593), .ZN(n6728) );
  NAND2_X1 U8227 ( .A1(n6728), .A2(n6729), .ZN(n6726) );
  NOR2_X1 U8228 ( .A1(n6742), .A2(n6739), .ZN(n6738) );
  INV_X1 U8229 ( .A(n8233), .ZN(n6741) );
  INV_X1 U8230 ( .A(n8232), .ZN(n7057) );
  INV_X1 U8231 ( .A(n7167), .ZN(n7166) );
  AOI21_X1 U8232 ( .B1(n7167), .B2(n7165), .A(n7164), .ZN(n7163) );
  INV_X1 U8233 ( .A(n8103), .ZN(n7164) );
  INV_X1 U8234 ( .A(n8080), .ZN(n7165) );
  NOR2_X1 U8235 ( .A1(n6506), .A2(n7170), .ZN(n7169) );
  INV_X1 U8236 ( .A(n7982), .ZN(n7170) );
  OR2_X1 U8237 ( .A1(n13190), .A2(n12946), .ZN(n9131) );
  NOR2_X1 U8238 ( .A1(n13202), .A2(n13208), .ZN(n6954) );
  NAND2_X1 U8239 ( .A1(n7106), .A2(n7104), .ZN(n7103) );
  INV_X1 U8240 ( .A(n12934), .ZN(n7104) );
  NAND2_X1 U8241 ( .A1(n6946), .A2(n13155), .ZN(n6945) );
  INV_X1 U8242 ( .A(n6947), .ZN(n6946) );
  NAND2_X1 U8243 ( .A1(n6872), .A2(n6875), .ZN(n6871) );
  INV_X1 U8244 ( .A(n6492), .ZN(n7247) );
  NOR2_X1 U8245 ( .A1(n10875), .A2(n10653), .ZN(n6957) );
  AND2_X1 U8246 ( .A1(n10441), .A2(n14909), .ZN(n10252) );
  INV_X1 U8247 ( .A(n9926), .ZN(n6869) );
  NOR2_X1 U8248 ( .A1(n7096), .A2(n7094), .ZN(n7093) );
  INV_X1 U8249 ( .A(n9929), .ZN(n7094) );
  INV_X1 U8250 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8174) );
  OR3_X1 U8251 ( .A1(n7688), .A2(P2_IR_REG_6__SCAN_IN), .A3(
        P2_IR_REG_7__SCAN_IN), .ZN(n7700) );
  OR2_X1 U8252 ( .A1(n7770), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n7688) );
  INV_X1 U8253 ( .A(n13385), .ZN(n7394) );
  NAND2_X1 U8254 ( .A1(n6779), .A2(n9544), .ZN(n7448) );
  NAND2_X1 U8255 ( .A1(n7236), .A2(n7235), .ZN(n13508) );
  NOR2_X1 U8256 ( .A1(n13508), .A2(n13503), .ZN(n13506) );
  NAND2_X1 U8257 ( .A1(n13700), .A2(n13702), .ZN(n7270) );
  INV_X1 U8258 ( .A(n11557), .ZN(n9632) );
  AOI21_X1 U8259 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n13833), .A(n13832), .ZN(
        n13842) );
  NOR2_X1 U8260 ( .A1(n13998), .A2(n13978), .ZN(n13958) );
  NOR2_X1 U8261 ( .A1(n14025), .A2(n14010), .ZN(n6942) );
  INV_X1 U8262 ( .A(n11543), .ZN(n11559) );
  NAND2_X1 U8263 ( .A1(n11559), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11558) );
  NAND2_X1 U8264 ( .A1(n11542), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11543) );
  INV_X1 U8265 ( .A(n13642), .ZN(n13659) );
  OR2_X1 U8266 ( .A1(n13638), .A2(n14084), .ZN(n11503) );
  NOR2_X1 U8267 ( .A1(n13474), .A2(n13473), .ZN(n7406) );
  NAND2_X1 U8268 ( .A1(n10555), .A2(n10282), .ZN(n7356) );
  AND2_X1 U8269 ( .A1(n13523), .A2(n9744), .ZN(n9742) );
  NAND2_X1 U8270 ( .A1(n7230), .A2(n7231), .ZN(n9084) );
  AOI21_X1 U8271 ( .B1(n7232), .B2(n8158), .A(n6614), .ZN(n7231) );
  NAND4_X1 U8272 ( .A1(n9188), .A2(n9284), .A3(n9286), .A4(n9187), .ZN(n9193)
         );
  INV_X1 U8273 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9187) );
  AOI21_X1 U8274 ( .B1(n8003), .B2(n7225), .A(n8021), .ZN(n7223) );
  NAND2_X1 U8275 ( .A1(n7967), .A2(n7966), .ZN(n7985) );
  NAND2_X1 U8276 ( .A1(n7965), .A2(SI_20_), .ZN(n7966) );
  AND2_X1 U8277 ( .A1(n7941), .A2(n7922), .ZN(n7939) );
  INV_X1 U8278 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n9185) );
  AOI21_X1 U8279 ( .B1(n7221), .B2(n7728), .A(n6559), .ZN(n7219) );
  INV_X1 U8280 ( .A(n7221), .ZN(n7220) );
  INV_X1 U8281 ( .A(n7681), .ZN(n6916) );
  NAND2_X1 U8282 ( .A1(n9212), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6934) );
  INV_X1 U8283 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14261) );
  AOI21_X1 U8284 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14277), .A(n14276), .ZN(
        n14322) );
  NOR2_X1 U8285 ( .A1(n14294), .A2(n14293), .ZN(n14276) );
  OR2_X1 U8286 ( .A1(n14281), .A2(n14280), .ZN(n14328) );
  NAND2_X1 U8287 ( .A1(n12116), .A2(n6794), .ZN(n6793) );
  INV_X1 U8288 ( .A(n8890), .ZN(n6794) );
  INV_X1 U8289 ( .A(n11999), .ZN(n6795) );
  INV_X1 U8290 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n12217) );
  OAI21_X1 U8291 ( .B1(n12059), .B2(n8865), .A(n8867), .ZN(n12067) );
  AND2_X1 U8292 ( .A1(n8642), .A2(n12014), .ZN(n8655) );
  INV_X1 U8293 ( .A(n8884), .ZN(n12075) );
  NAND2_X1 U8294 ( .A1(n8435), .A2(n6960), .ZN(n11403) );
  INV_X1 U8295 ( .A(n6961), .ZN(n6960) );
  OAI21_X1 U8296 ( .B1(n8310), .B2(SI_9_), .A(n8434), .ZN(n6961) );
  INV_X1 U8297 ( .A(n15101), .ZN(n11681) );
  XNOR2_X1 U8298 ( .A(n10434), .B(n8852), .ZN(n8822) );
  OAI22_X1 U8299 ( .A1(n11842), .A2(n15113), .B1(n11844), .B2(n11843), .ZN(
        n6754) );
  NAND2_X1 U8300 ( .A1(n11840), .A2(n6745), .ZN(n6744) );
  NOR2_X1 U8301 ( .A1(n11837), .A2(n6746), .ZN(n6745) );
  INV_X1 U8302 ( .A(n11841), .ZN(n6820) );
  OR2_X1 U8303 ( .A1(n8357), .A2(n9998), .ZN(n8289) );
  AOI21_X1 U8304 ( .B1(n10051), .B2(n10196), .A(n9995), .ZN(n10044) );
  AND2_X1 U8305 ( .A1(n10044), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10046) );
  NAND2_X1 U8306 ( .A1(n10074), .A2(n10001), .ZN(n10101) );
  NAND2_X1 U8307 ( .A1(n10101), .A2(n10100), .ZN(n10099) );
  XNOR2_X1 U8308 ( .A(n10004), .B(n6695), .ZN(n10026) );
  XNOR2_X1 U8309 ( .A(n10762), .B(n10770), .ZN(n10669) );
  XNOR2_X1 U8310 ( .A(n12334), .B(n12333), .ZN(n14977) );
  INV_X1 U8311 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n15017) );
  NAND2_X1 U8312 ( .A1(n15021), .A2(n12301), .ZN(n15043) );
  OR2_X1 U8313 ( .A1(n15043), .A2(n15044), .ZN(n15040) );
  AND2_X1 U8314 ( .A1(n14410), .A2(n14409), .ZN(n14411) );
  NAND2_X1 U8315 ( .A1(n14407), .A2(n12346), .ZN(n14427) );
  NOR2_X1 U8316 ( .A1(n14411), .A2(n6701), .ZN(n14433) );
  NOR2_X1 U8317 ( .A1(n6702), .A2(n14413), .ZN(n6701) );
  INV_X1 U8318 ( .A(n12308), .ZN(n6702) );
  NOR2_X1 U8319 ( .A1(n14422), .A2(n12323), .ZN(n12325) );
  XNOR2_X1 U8320 ( .A(n12348), .B(n6698), .ZN(n14444) );
  AOI21_X1 U8321 ( .B1(n14444), .B2(P3_REG1_REG_17__SCAN_IN), .A(n6697), .ZN(
        n12362) );
  AND2_X1 U8322 ( .A1(n12348), .A2(n12349), .ZN(n6697) );
  OR2_X1 U8323 ( .A1(n14459), .A2(n8221), .ZN(n12392) );
  OR2_X1 U8324 ( .A1(n8669), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8681) );
  INV_X1 U8325 ( .A(n7206), .ZN(n7205) );
  OAI21_X1 U8326 ( .B1(n7207), .B2(n8743), .A(n8744), .ZN(n7206) );
  NOR2_X1 U8327 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n8591), .ZN(n8600) );
  AND4_X1 U8328 ( .A1(n8607), .A2(n8606), .A3(n8605), .A4(n8604), .ZN(n12510)
         );
  OR2_X1 U8329 ( .A1(n12509), .A2(n12508), .ZN(n12513) );
  NAND2_X1 U8330 ( .A1(n12106), .A2(n8576), .ZN(n8591) );
  AND2_X1 U8331 ( .A1(n11760), .A2(n11765), .ZN(n12525) );
  NAND2_X1 U8332 ( .A1(n6974), .A2(n8566), .ZN(n12491) );
  NAND2_X1 U8333 ( .A1(n12542), .A2(n11830), .ZN(n6974) );
  OR2_X1 U8334 ( .A1(n12491), .A2(n12525), .ZN(n12523) );
  AND2_X1 U8335 ( .A1(n8558), .A2(n8557), .ZN(n8576) );
  AND4_X1 U8336 ( .A1(n8498), .A2(n8497), .A3(n8496), .A4(n8495), .ZN(n12581)
         );
  INV_X1 U8337 ( .A(n7191), .ZN(n7190) );
  AOI21_X1 U8338 ( .B1(n7189), .B2(n7191), .A(n7188), .ZN(n7187) );
  NOR2_X1 U8339 ( .A1(n8736), .A2(n7192), .ZN(n7191) );
  NOR2_X1 U8340 ( .A1(n8462), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8492) );
  INV_X1 U8341 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8491) );
  AND4_X1 U8342 ( .A1(n8446), .A2(n8445), .A3(n8444), .A4(n8443), .ZN(n12611)
         );
  AND2_X1 U8343 ( .A1(n8388), .A2(n12217), .ZN(n8420) );
  AND4_X1 U8344 ( .A1(n8394), .A2(n8393), .A3(n8392), .A4(n8391), .ZN(n11399)
         );
  NAND2_X1 U8345 ( .A1(n11714), .A2(n11715), .ZN(n11711) );
  OR2_X1 U8346 ( .A1(n8358), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8374) );
  NAND2_X1 U8347 ( .A1(n11057), .A2(n11056), .ZN(n11055) );
  AND2_X1 U8348 ( .A1(n8728), .A2(n11702), .ZN(n11814) );
  NAND2_X1 U8349 ( .A1(n11053), .A2(n11814), .ZN(n11052) );
  NAND2_X1 U8350 ( .A1(n10978), .A2(n11822), .ZN(n10977) );
  NAND2_X1 U8351 ( .A1(n8319), .A2(n8318), .ZN(n10687) );
  NAND2_X1 U8352 ( .A1(n10682), .A2(n11815), .ZN(n10681) );
  AND2_X2 U8353 ( .A1(n11689), .A2(n11693), .ZN(n15085) );
  NAND2_X1 U8354 ( .A1(n8755), .A2(n8789), .ZN(n15090) );
  AND4_X2 U8355 ( .A1(n8276), .A2(n8277), .A3(n8275), .A4(n8278), .ZN(n15107)
         );
  OR2_X1 U8356 ( .A1(n6429), .A2(n9907), .ZN(n8278) );
  AND3_X1 U8357 ( .A1(n8336), .A2(n8335), .A3(n8334), .ZN(n8827) );
  OR2_X1 U8358 ( .A1(n8310), .A2(SI_4_), .ZN(n8335) );
  INV_X1 U8359 ( .A(n9971), .ZN(n8918) );
  INV_X1 U8360 ( .A(n11661), .ZN(n7075) );
  NAND2_X1 U8361 ( .A1(n7061), .A2(n7060), .ZN(n8704) );
  AOI21_X1 U8362 ( .B1(n7064), .B2(n7069), .A(n6617), .ZN(n7060) );
  INV_X1 U8363 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n8215) );
  INV_X1 U8364 ( .A(n7071), .ZN(n7063) );
  XNOR2_X1 U8365 ( .A(n8787), .B(n8203), .ZN(n9968) );
  NAND2_X1 U8366 ( .A1(n8250), .A2(n8249), .ZN(n8613) );
  AND2_X1 U8367 ( .A1(n8718), .A2(n8717), .ZN(n8800) );
  XNOR2_X1 U8368 ( .A(n8248), .B(n10976), .ZN(n8597) );
  AND2_X1 U8369 ( .A1(n7193), .A2(n8212), .ZN(n8584) );
  INV_X1 U8370 ( .A(n7193), .ZN(n8570) );
  OAI211_X1 U8371 ( .C1(n8243), .C2(n7054), .A(n6731), .B(n7051), .ZN(n8515)
         );
  AOI21_X1 U8372 ( .B1(n7053), .B2(n7055), .A(n6601), .ZN(n7051) );
  OR2_X1 U8373 ( .A1(n8431), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n8449) );
  OR2_X1 U8374 ( .A1(n8399), .A2(P3_IR_REG_8__SCAN_IN), .ZN(n8431) );
  INV_X1 U8375 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n8330) );
  AND2_X2 U8376 ( .A1(n9975), .A2(n8192), .ZN(n8331) );
  NOR2_X1 U8377 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n8192) );
  XNOR2_X1 U8378 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8261) );
  AND2_X1 U8379 ( .A1(n8229), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8279) );
  NOR2_X1 U8380 ( .A1(n7648), .A2(n7647), .ZN(n7672) );
  NOR2_X1 U8381 ( .A1(n12750), .A2(n7168), .ZN(n7167) );
  INV_X1 U8382 ( .A(n8084), .ZN(n7168) );
  AOI21_X1 U8383 ( .B1(n9896), .B2(n7159), .A(n6520), .ZN(n7158) );
  INV_X1 U8384 ( .A(n7658), .ZN(n7159) );
  AND2_X1 U8385 ( .A1(n9896), .A2(n7161), .ZN(n7157) );
  NAND2_X1 U8386 ( .A1(n7776), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7796) );
  OR2_X1 U8387 ( .A1(n7796), .A2(n10970), .ZN(n7819) );
  XNOR2_X1 U8388 ( .A(n8119), .B(n11644), .ZN(n7533) );
  NAND2_X1 U8389 ( .A1(n7903), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n7927) );
  OR2_X1 U8390 ( .A1(n8176), .A2(n9397), .ZN(n12913) );
  CLKBUF_X1 U8391 ( .A(n7162), .Z(n6625) );
  INV_X1 U8392 ( .A(n14833), .ZN(n8118) );
  AND2_X1 U8393 ( .A1(n7955), .A2(n7954), .ZN(n12967) );
  AND4_X1 U8394 ( .A1(n7711), .A2(n7710), .A3(n7709), .A4(n7708), .ZN(n10582)
         );
  AND4_X1 U8395 ( .A1(n7718), .A2(n7717), .A3(n7716), .A4(n7715), .ZN(n10475)
         );
  AND4_X1 U8396 ( .A1(n7626), .A2(n7625), .A3(n7624), .A4(n7623), .ZN(n10155)
         );
  XNOR2_X1 U8397 ( .A(n14742), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n14746) );
  NAND2_X1 U8398 ( .A1(n14751), .A2(n9375), .ZN(n14766) );
  AND2_X1 U8399 ( .A1(n14766), .A2(n14767), .ZN(n14763) );
  NOR2_X1 U8400 ( .A1(n14763), .A2(n6839), .ZN(n9422) );
  NOR2_X1 U8401 ( .A1(n9388), .A2(n6840), .ZN(n6839) );
  OR2_X1 U8402 ( .A1(n9559), .A2(n9558), .ZN(n6843) );
  AND2_X1 U8403 ( .A1(n6843), .A2(n6842), .ZN(n9587) );
  NAND2_X1 U8404 ( .A1(n9590), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6842) );
  NAND2_X1 U8405 ( .A1(n9587), .A2(n9586), .ZN(n9795) );
  NOR2_X1 U8406 ( .A1(n10136), .A2(n6850), .ZN(n10140) );
  AND2_X1 U8407 ( .A1(n10137), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6850) );
  NOR2_X1 U8408 ( .A1(n10140), .A2(n10139), .ZN(n10305) );
  AND2_X1 U8409 ( .A1(n10132), .A2(n10131), .ZN(n10314) );
  NOR2_X1 U8410 ( .A1(n10305), .A2(n6849), .ZN(n10306) );
  AND2_X1 U8411 ( .A1(n10308), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8412 ( .A1(n10306), .A2(n10307), .ZN(n10692) );
  NOR2_X1 U8413 ( .A1(n10867), .A2(n6848), .ZN(n10869) );
  AND2_X1 U8414 ( .A1(n10868), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6848) );
  NOR2_X1 U8415 ( .A1(n10869), .A2(n10870), .ZN(n11184) );
  NOR2_X1 U8416 ( .A1(n11184), .A2(n6847), .ZN(n11336) );
  AND2_X1 U8417 ( .A1(n11185), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U8418 ( .A1(n14794), .A2(n6615), .ZN(n12896) );
  NOR2_X1 U8419 ( .A1(n12883), .A2(n12884), .ZN(n12898) );
  OAI21_X1 U8420 ( .B1(n12875), .B2(n12876), .A(n14801), .ZN(n12890) );
  INV_X1 U8421 ( .A(n7486), .ZN(n7500) );
  NAND2_X1 U8422 ( .A1(n9072), .A2(n9071), .ZN(n9151) );
  NAND2_X1 U8423 ( .A1(n12996), .A2(n6671), .ZN(n12945) );
  OR2_X1 U8424 ( .A1(n13190), .A2(n12943), .ZN(n6671) );
  NAND2_X1 U8425 ( .A1(n7078), .A2(n13006), .ZN(n7077) );
  AOI21_X1 U8426 ( .B1(n7255), .B2(n12982), .A(n6516), .ZN(n7253) );
  INV_X1 U8427 ( .A(n12986), .ZN(n12994) );
  AND2_X1 U8428 ( .A1(n13016), .A2(n12984), .ZN(n7255) );
  AND2_X1 U8429 ( .A1(n8106), .A2(n8072), .ZN(n13026) );
  NAND2_X1 U8430 ( .A1(n13055), .A2(n6954), .ZN(n13023) );
  NAND2_X1 U8431 ( .A1(n12971), .A2(n6879), .ZN(n6878) );
  AOI21_X1 U8432 ( .B1(n12971), .B2(n6882), .A(n12970), .ZN(n6877) );
  NAND2_X1 U8433 ( .A1(n6886), .A2(n6484), .ZN(n6885) );
  INV_X1 U8434 ( .A(n12966), .ZN(n6886) );
  NOR3_X1 U8435 ( .A1(n11368), .A2(n6945), .A3(n6949), .ZN(n13139) );
  INV_X1 U8436 ( .A(n7100), .ZN(n7099) );
  AOI21_X1 U8437 ( .B1(n7100), .B2(n7098), .A(n6546), .ZN(n7097) );
  AOI21_X1 U8438 ( .B1(n13165), .B2(n12927), .A(n6518), .ZN(n7100) );
  NOR2_X1 U8439 ( .A1(n11368), .A2(n6945), .ZN(n13150) );
  AOI21_X1 U8440 ( .B1(n7241), .B2(n11358), .A(n6512), .ZN(n7240) );
  NAND2_X1 U8441 ( .A1(n7836), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7862) );
  INV_X1 U8442 ( .A(n7837), .ZN(n7836) );
  AND2_X1 U8443 ( .A1(n14520), .A2(n11132), .ZN(n11276) );
  NAND2_X1 U8444 ( .A1(n11265), .A2(n11264), .ZN(n11267) );
  OAI21_X1 U8445 ( .B1(n11133), .B2(n11138), .A(n11115), .ZN(n11265) );
  NAND2_X1 U8446 ( .A1(n7119), .A2(n7118), .ZN(n14509) );
  AOI21_X1 U8447 ( .B1(n7120), .B2(n10585), .A(n6529), .ZN(n7118) );
  NAND2_X1 U8448 ( .A1(n10479), .A2(n6957), .ZN(n10885) );
  NAND2_X1 U8449 ( .A1(n10479), .A2(n14923), .ZN(n10587) );
  AOI21_X1 U8450 ( .B1(n10448), .B2(n6891), .A(n10245), .ZN(n6890) );
  INV_X1 U8451 ( .A(n10243), .ZN(n6891) );
  NAND2_X1 U8452 ( .A1(n6674), .A2(n10448), .ZN(n6889) );
  INV_X1 U8453 ( .A(n10244), .ZN(n6674) );
  NAND2_X1 U8454 ( .A1(n7111), .A2(n7110), .ZN(n10450) );
  AND2_X1 U8455 ( .A1(n10248), .A2(n7112), .ZN(n7111) );
  AND2_X1 U8456 ( .A1(n10163), .A2(n10247), .ZN(n10441) );
  NAND2_X1 U8457 ( .A1(n7117), .A2(n7116), .ZN(n7115) );
  NAND2_X1 U8458 ( .A1(n7115), .A2(n7113), .ZN(n10447) );
  NOR2_X1 U8459 ( .A1(n10174), .A2(n9942), .ZN(n10163) );
  AND2_X1 U8460 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7621) );
  XNOR2_X1 U8461 ( .A(n9942), .B(n12866), .ZN(n10152) );
  NAND2_X1 U8462 ( .A1(n6944), .A2(n14887), .ZN(n10174) );
  NAND2_X1 U8463 ( .A1(n9930), .A2(n9929), .ZN(n14811) );
  NAND2_X1 U8464 ( .A1(n11636), .A2(n9928), .ZN(n10536) );
  NAND2_X1 U8465 ( .A1(n11637), .A2(n11638), .ZN(n11636) );
  NAND2_X1 U8466 ( .A1(n7250), .A2(n11123), .ZN(n11137) );
  NAND2_X1 U8467 ( .A1(n7251), .A2(n6492), .ZN(n7250) );
  INV_X1 U8468 ( .A(n14504), .ZN(n7251) );
  CLKBUF_X1 U8469 ( .A(n14936), .Z(n6660) );
  OR2_X1 U8470 ( .A1(n7584), .A2(n9674), .ZN(n7549) );
  XNOR2_X1 U8471 ( .A(n8140), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8149) );
  AND2_X1 U8472 ( .A1(n7507), .A2(n6474), .ZN(n7252) );
  OR2_X1 U8473 ( .A1(n8136), .A2(n13281), .ZN(n7483) );
  INV_X1 U8474 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n7494) );
  NOR2_X1 U8475 ( .A1(n7700), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n7704) );
  INV_X1 U8476 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n7453) );
  INV_X1 U8477 ( .A(n6773), .ZN(n6771) );
  OR2_X1 U8478 ( .A1(n7382), .A2(n7442), .ZN(n7380) );
  AND2_X1 U8479 ( .A1(n13407), .A2(n7383), .ZN(n7382) );
  NAND2_X1 U8480 ( .A1(n7384), .A2(n11908), .ZN(n7383) );
  INV_X1 U8481 ( .A(n13368), .ZN(n7384) );
  NAND2_X1 U8482 ( .A1(n7385), .A2(n11908), .ZN(n7381) );
  OR2_X1 U8483 ( .A1(n9538), .A2(n13716), .ZN(n9780) );
  INV_X1 U8484 ( .A(n13307), .ZN(n7389) );
  INV_X1 U8485 ( .A(n13416), .ZN(n7392) );
  INV_X1 U8486 ( .A(n11958), .ZN(n7391) );
  INV_X1 U8487 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10286) );
  NOR2_X1 U8488 ( .A1(n13330), .A2(n7397), .ZN(n7396) );
  INV_X1 U8489 ( .A(n11925), .ZN(n7397) );
  NAND2_X1 U8490 ( .A1(n13425), .A2(n7398), .ZN(n13357) );
  AND2_X1 U8491 ( .A1(n11900), .A2(n7399), .ZN(n7398) );
  INV_X1 U8492 ( .A(n13360), .ZN(n7399) );
  INV_X1 U8493 ( .A(n10408), .ZN(n6760) );
  NAND2_X1 U8494 ( .A1(n6766), .A2(n6764), .ZN(n6763) );
  OR2_X1 U8495 ( .A1(n10321), .A2(n6765), .ZN(n6762) );
  NAND2_X1 U8496 ( .A1(n6767), .A2(n10326), .ZN(n6765) );
  AND2_X1 U8497 ( .A1(n11530), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11542) );
  NAND2_X1 U8498 ( .A1(n13399), .A2(n13400), .ZN(n13398) );
  AND2_X1 U8499 ( .A1(n10828), .A2(n10827), .ZN(n10904) );
  NOR2_X1 U8500 ( .A1(n10496), .A2(n11044), .ZN(n10828) );
  NAND2_X1 U8501 ( .A1(n14555), .A2(n14554), .ZN(n14568) );
  INV_X1 U8502 ( .A(n14554), .ZN(n7376) );
  AND2_X1 U8503 ( .A1(n11870), .A2(n7374), .ZN(n7373) );
  NAND2_X1 U8504 ( .A1(n14554), .A2(n7375), .ZN(n7374) );
  INV_X1 U8505 ( .A(n11858), .ZN(n7375) );
  NAND2_X1 U8506 ( .A1(n13367), .A2(n13368), .ZN(n13366) );
  OR2_X1 U8507 ( .A1(n11437), .A2(n11436), .ZN(n11518) );
  NAND2_X1 U8508 ( .A1(n11237), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11437) );
  NAND2_X1 U8509 ( .A1(n14542), .A2(n11893), .ZN(n11899) );
  NAND2_X1 U8510 ( .A1(n13506), .A2(n13711), .ZN(n13510) );
  INV_X2 U8511 ( .A(n6428), .ZN(n11600) );
  NAND2_X1 U8512 ( .A1(n9632), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9638) );
  AOI22_X1 U8513 ( .A1(n9661), .A2(n9662), .B1(P1_REG1_REG_4__SCAN_IN), .B2(
        n9837), .ZN(n9304) );
  NAND2_X1 U8514 ( .A1(n9411), .A2(n6676), .ZN(n9412) );
  OR2_X1 U8515 ( .A1(n10488), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8516 ( .A1(n9412), .A2(n9413), .ZN(n9601) );
  AOI21_X1 U8517 ( .B1(n10822), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9728), .ZN(
        n9730) );
  NAND2_X1 U8518 ( .A1(n9821), .A2(n6675), .ZN(n9822) );
  OR2_X1 U8519 ( .A1(n10913), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8520 ( .A1(n9822), .A2(n9823), .ZN(n10415) );
  AOI21_X1 U8521 ( .B1(n13818), .B2(P1_REG1_REG_16__SCAN_IN), .A(n13817), .ZN(
        n13821) );
  NAND2_X1 U8522 ( .A1(n9298), .A2(n7361), .ZN(n9320) );
  NAND2_X1 U8523 ( .A1(n9195), .A2(n12257), .ZN(n10458) );
  NAND2_X1 U8524 ( .A1(n13807), .A2(n11513), .ZN(n6679) );
  INV_X1 U8525 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n13325) );
  NAND2_X1 U8526 ( .A1(n13877), .A2(n13913), .ZN(n7425) );
  INV_X1 U8527 ( .A(n14115), .ZN(n13877) );
  OAI21_X1 U8528 ( .B1(n13916), .B2(n6901), .A(n6899), .ZN(n13876) );
  NAND2_X1 U8529 ( .A1(n13915), .A2(n11598), .ZN(n11599) );
  INV_X1 U8530 ( .A(n6943), .ZN(n13936) );
  INV_X1 U8531 ( .A(n6908), .ZN(n6907) );
  AOI21_X1 U8532 ( .B1(n6908), .B2(n13493), .A(n7360), .ZN(n6906) );
  OR2_X1 U8533 ( .A1(n14142), .A2(n13990), .ZN(n7439) );
  INV_X1 U8534 ( .A(n11570), .ZN(n11494) );
  AND2_X1 U8535 ( .A1(n13979), .A2(n6908), .ZN(n13950) );
  NAND2_X1 U8536 ( .A1(n13979), .A2(n7441), .ZN(n13951) );
  INV_X1 U8537 ( .A(n13732), .ZN(n13990) );
  NAND2_X1 U8538 ( .A1(n11571), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11570) );
  NAND2_X1 U8539 ( .A1(n13980), .A2(n7434), .ZN(n13979) );
  AOI21_X1 U8540 ( .B1(n7422), .B2(n14033), .A(n7420), .ZN(n7419) );
  INV_X1 U8541 ( .A(n7422), .ZN(n7421) );
  INV_X1 U8542 ( .A(n11552), .ZN(n7420) );
  NAND2_X1 U8543 ( .A1(n6942), .A2(n7363), .ZN(n13998) );
  INV_X1 U8544 ( .A(n6942), .ZN(n14012) );
  NOR2_X1 U8545 ( .A1(n14063), .A2(n14043), .ZN(n14042) );
  OR2_X1 U8546 ( .A1(n14175), .A2(n14065), .ZN(n14063) );
  AND2_X1 U8547 ( .A1(n11096), .A2(n6479), .ZN(n14074) );
  NAND2_X1 U8548 ( .A1(n11096), .A2(n6939), .ZN(n14076) );
  AOI21_X1 U8549 ( .B1(n7430), .B2(n13617), .A(n6543), .ZN(n7429) );
  NAND2_X1 U8550 ( .A1(n11096), .A2(n14582), .ZN(n11324) );
  AOI21_X1 U8551 ( .B1(n7415), .B2(n7417), .A(n6544), .ZN(n7412) );
  INV_X1 U8552 ( .A(n10919), .ZN(n10920) );
  AND2_X1 U8553 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9856) );
  NAND2_X1 U8554 ( .A1(n10221), .A2(n13473), .ZN(n10281) );
  NAND2_X1 U8555 ( .A1(n9544), .A2(n9235), .ZN(n13715) );
  INV_X1 U8556 ( .A(n13539), .ZN(n13470) );
  NAND2_X1 U8557 ( .A1(n7351), .A2(n7352), .ZN(n11327) );
  NAND2_X1 U8558 ( .A1(n9834), .A2(n6914), .ZN(n14706) );
  AOI22_X1 U8559 ( .A1(n11514), .A2(n9833), .B1(n7361), .B2(n6523), .ZN(n6914)
         );
  INV_X1 U8560 ( .A(n14587), .ZN(n14712) );
  OAI21_X1 U8561 ( .B1(n9068), .B2(n9069), .A(n9062), .ZN(n7215) );
  XNOR2_X1 U8562 ( .A(n9084), .B(n9083), .ZN(n13462) );
  XNOR2_X1 U8563 ( .A(n8159), .B(n8089), .ZN(n13293) );
  OR2_X1 U8564 ( .A1(n10458), .A2(n9193), .ZN(n9200) );
  NAND2_X1 U8565 ( .A1(n9495), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9493) );
  NAND2_X1 U8566 ( .A1(n7229), .A2(n7897), .ZN(n7917) );
  NAND2_X1 U8567 ( .A1(n6923), .A2(n6928), .ZN(n7872) );
  OR2_X1 U8568 ( .A1(n6708), .A2(n6930), .ZN(n6923) );
  NAND2_X1 U8569 ( .A1(n6927), .A2(n7831), .ZN(n7852) );
  NAND2_X1 U8570 ( .A1(n6708), .A2(n6932), .ZN(n6927) );
  NAND2_X1 U8571 ( .A1(n7750), .A2(n7749), .ZN(n7769) );
  OR2_X1 U8572 ( .A1(n10035), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n9354) );
  OR2_X1 U8573 ( .A1(n9354), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n9876) );
  AND2_X1 U8574 ( .A1(n9234), .A2(n9245), .ZN(n10214) );
  OAI21_X1 U8575 ( .B1(n9212), .B2(P2_DATAO_REG_0__SCAN_IN), .A(n6673), .ZN(
        n7477) );
  NAND2_X1 U8576 ( .A1(n9212), .A2(n8229), .ZN(n6673) );
  AND2_X1 U8577 ( .A1(n14258), .A2(P3_ADDR_REG_1__SCAN_IN), .ZN(n7136) );
  INV_X1 U8578 ( .A(n14299), .ZN(n7138) );
  INV_X1 U8579 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n14258) );
  XNOR2_X1 U8580 ( .A(n14295), .B(P1_ADDR_REG_4__SCAN_IN), .ZN(n14296) );
  NOR2_X1 U8581 ( .A1(n14269), .A2(n14268), .ZN(n14312) );
  OR2_X1 U8582 ( .A1(n14374), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n6851) );
  OAI21_X1 U8583 ( .B1(n14381), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n7447), .ZN(
        n14335) );
  AOI22_X1 U8584 ( .A1(P3_ADDR_REG_11__SCAN_IN), .A2(n14285), .B1(n14332), 
        .B2(n14284), .ZN(n14338) );
  INV_X1 U8585 ( .A(n7148), .ZN(n7146) );
  OR2_X1 U8586 ( .A1(n14608), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7148) );
  INV_X1 U8587 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n6865) );
  OR2_X1 U8588 ( .A1(n14611), .A2(P2_ADDR_REG_15__SCAN_IN), .ZN(n14349) );
  AND4_X1 U8589 ( .A1(n8541), .A2(n8540), .A3(n8539), .A4(n8538), .ZN(n12582)
         );
  INV_X1 U8590 ( .A(n12700), .ZN(n12019) );
  AND4_X1 U8591 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n12511)
         );
  AOI21_X1 U8592 ( .B1(n8817), .B2(n10202), .A(n8816), .ZN(n8819) );
  NAND2_X1 U8593 ( .A1(n12043), .A2(n12042), .ZN(n12041) );
  INV_X1 U8594 ( .A(n12572), .ZN(n12070) );
  NAND2_X1 U8595 ( .A1(n10528), .A2(n8826), .ZN(n10746) );
  NAND2_X1 U8596 ( .A1(n7006), .A2(n8843), .ZN(n11068) );
  NAND2_X1 U8597 ( .A1(n8629), .A2(n8628), .ZN(n12472) );
  NAND2_X1 U8598 ( .A1(n10430), .A2(n10431), .ZN(n10527) );
  NAND2_X1 U8599 ( .A1(n8906), .A2(n8905), .ZN(n12117) );
  AND4_X1 U8600 ( .A1(n8380), .A2(n8379), .A3(n8378), .A4(n8377), .ZN(n11210)
         );
  OR2_X1 U8601 ( .A1(n8910), .A2(n11847), .ZN(n12126) );
  NAND2_X1 U8602 ( .A1(n12006), .A2(n8861), .ZN(n12125) );
  INV_X1 U8603 ( .A(n12511), .ZN(n12543) );
  INV_X1 U8604 ( .A(n12582), .ZN(n12556) );
  INV_X1 U8605 ( .A(n12581), .ZN(n12140) );
  INV_X1 U8606 ( .A(n12611), .ZN(n12142) );
  INV_X1 U8607 ( .A(n11398), .ZN(n12143) );
  INV_X1 U8608 ( .A(n11399), .ZN(n12145) );
  INV_X1 U8609 ( .A(n11210), .ZN(n12146) );
  INV_X1 U8610 ( .A(n10747), .ZN(n12148) );
  OR2_X1 U8611 ( .A1(n11655), .A2(n8304), .ZN(n8307) );
  NOR2_X1 U8612 ( .A1(n6491), .A2(n8271), .ZN(n6636) );
  INV_X1 U8613 ( .A(n15107), .ZN(n12285) );
  NOR2_X1 U8614 ( .A1(n9203), .A2(n9325), .ZN(n12284) );
  INV_X1 U8615 ( .A(n9999), .ZN(n10082) );
  NAND2_X1 U8616 ( .A1(n9963), .A2(n9962), .ZN(n10020) );
  INV_X1 U8617 ( .A(n7033), .ZN(n9988) );
  NAND2_X1 U8618 ( .A1(n10389), .A2(n10390), .ZN(n10393) );
  NAND2_X1 U8619 ( .A1(n10393), .A2(n10392), .ZN(n10667) );
  INV_X1 U8620 ( .A(n7035), .ZN(n10400) );
  NAND2_X1 U8621 ( .A1(n10761), .A2(n10760), .ZN(n12287) );
  INV_X1 U8622 ( .A(n7030), .ZN(n10774) );
  NAND2_X1 U8623 ( .A1(n7023), .A2(n7021), .ZN(n7024) );
  AND2_X1 U8624 ( .A1(n7022), .A2(n12339), .ZN(n7021) );
  NAND2_X1 U8625 ( .A1(n14987), .A2(n7019), .ZN(n7025) );
  OR2_X1 U8626 ( .A1(n12317), .A2(n15024), .ZN(n7027) );
  INV_X1 U8627 ( .A(n7031), .ZN(n14404) );
  INV_X1 U8628 ( .A(n12324), .ZN(n14441) );
  NAND2_X1 U8629 ( .A1(n12416), .A2(n11797), .ZN(n7201) );
  NAND2_X1 U8630 ( .A1(n12435), .A2(n8676), .ZN(n12418) );
  NAND2_X1 U8631 ( .A1(n8664), .A2(n8663), .ZN(n12432) );
  NAND2_X1 U8632 ( .A1(n8668), .A2(n8667), .ZN(n12631) );
  AND2_X1 U8633 ( .A1(n8653), .A2(n8652), .ZN(n12638) );
  NAND2_X1 U8634 ( .A1(n12490), .A2(n8743), .ZN(n12478) );
  NAND2_X1 U8635 ( .A1(n8575), .A2(n8574), .ZN(n12539) );
  OAI21_X1 U8636 ( .B1(n6683), .B2(n11829), .A(n7178), .ZN(n12560) );
  NAND2_X1 U8637 ( .A1(n6683), .A2(n11745), .ZN(n12577) );
  NAND2_X1 U8638 ( .A1(n11387), .A2(n11736), .ZN(n12592) );
  NAND2_X1 U8639 ( .A1(n8488), .A2(n8487), .ZN(n14475) );
  NAND2_X1 U8640 ( .A1(n11383), .A2(n8482), .ZN(n12593) );
  OAI21_X1 U8641 ( .B1(n6684), .B2(n7186), .A(n7183), .ZN(n11321) );
  NAND2_X1 U8642 ( .A1(n6684), .A2(n8732), .ZN(n12602) );
  AND3_X1 U8643 ( .A1(n8417), .A2(n8416), .A3(n8415), .ZN(n12615) );
  AND3_X1 U8644 ( .A1(n8386), .A2(n8385), .A3(n8384), .ZN(n15057) );
  NAND2_X1 U8645 ( .A1(n10728), .A2(n6978), .ZN(n10980) );
  INV_X1 U8646 ( .A(n12587), .ZN(n15081) );
  NAND2_X1 U8647 ( .A1(n10368), .A2(n12375), .ZN(n15113) );
  NAND2_X1 U8648 ( .A1(n15120), .A2(n15095), .ZN(n15116) );
  INV_X1 U8649 ( .A(n15114), .ZN(n15098) );
  INV_X1 U8650 ( .A(n6987), .ZN(n6983) );
  NAND2_X1 U8651 ( .A1(n6981), .A2(n15109), .ZN(n6984) );
  NAND2_X1 U8652 ( .A1(n15149), .A2(n14476), .ZN(n12682) );
  AND2_X1 U8653 ( .A1(n14467), .A2(n14466), .ZN(n14486) );
  NAND2_X1 U8654 ( .A1(n15144), .A2(n8811), .ZN(n6985) );
  INV_X1 U8655 ( .A(n12412), .ZN(n12690) );
  NOR2_X1 U8656 ( .A1(n6648), .A2(n12623), .ZN(n12687) );
  AND2_X1 U8657 ( .A1(n12624), .A2(n6605), .ZN(n6648) );
  INV_X1 U8658 ( .A(n11776), .ZN(n12708) );
  OR2_X1 U8659 ( .A1(n12654), .A2(n12653), .ZN(n12709) );
  NAND2_X1 U8660 ( .A1(n8590), .A2(n8589), .ZN(n12713) );
  INV_X1 U8661 ( .A(n15057), .ZN(n11180) );
  INV_X1 U8662 ( .A(n8827), .ZN(n11703) );
  INV_X1 U8663 ( .A(n8726), .ZN(n10785) );
  NAND2_X1 U8664 ( .A1(n8771), .A2(n8770), .ZN(n10183) );
  XNOR2_X1 U8665 ( .A(n7074), .B(n7073), .ZN(n12731) );
  INV_X1 U8666 ( .A(n11651), .ZN(n7073) );
  OAI22_X1 U8667 ( .A1(n11660), .A2(n7075), .B1(n13446), .B2(
        P1_DATAO_REG_30__SCAN_IN), .ZN(n7074) );
  NAND2_X1 U8668 ( .A1(n6623), .A2(n6622), .ZN(n12729) );
  INV_X1 U8669 ( .A(n8218), .ZN(n6623) );
  XNOR2_X1 U8670 ( .A(n8692), .B(n8691), .ZN(n12740) );
  NAND2_X1 U8671 ( .A1(n7067), .A2(n7062), .ZN(n8692) );
  NOR2_X1 U8672 ( .A1(n7066), .A2(n7063), .ZN(n7062) );
  INV_X1 U8673 ( .A(SI_26_), .ZN(n12745) );
  INV_X1 U8674 ( .A(n7072), .ZN(n7068) );
  OAI21_X1 U8675 ( .B1(n8756), .B2(n7014), .A(n7012), .ZN(n8758) );
  NAND2_X1 U8676 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_24__SCAN_IN), 
        .ZN(n7014) );
  INV_X1 U8677 ( .A(n7050), .ZN(n8639) );
  NOR2_X1 U8678 ( .A1(n6797), .A2(n8765), .ZN(n6796) );
  INV_X1 U8679 ( .A(SI_19_), .ZN(n9809) );
  INV_X1 U8680 ( .A(SI_17_), .ZN(n9653) );
  INV_X1 U8681 ( .A(SI_15_), .ZN(n9532) );
  NAND2_X1 U8682 ( .A1(n7052), .A2(n8244), .ZN(n8528) );
  NAND2_X1 U8683 ( .A1(n8502), .A2(n8500), .ZN(n7052) );
  INV_X1 U8684 ( .A(SI_13_), .ZN(n9333) );
  INV_X1 U8685 ( .A(SI_12_), .ZN(n9244) );
  OAI21_X1 U8686 ( .B1(n8239), .B2(n7044), .A(n6736), .ZN(n8469) );
  INV_X1 U8687 ( .A(SI_11_), .ZN(n9260) );
  NAND2_X1 U8688 ( .A1(n7042), .A2(n8240), .ZN(n8448) );
  NAND2_X1 U8689 ( .A1(n8412), .A2(n8411), .ZN(n7042) );
  INV_X1 U8690 ( .A(n6727), .ZN(n8395) );
  AOI21_X1 U8691 ( .B1(n8382), .B2(n8381), .A(n6729), .ZN(n6727) );
  NAND2_X1 U8692 ( .A1(n6743), .A2(n8233), .ZN(n8350) );
  NAND2_X1 U8693 ( .A1(n8328), .A2(n8327), .ZN(n6743) );
  NAND2_X1 U8694 ( .A1(n7059), .A2(n8232), .ZN(n8313) );
  NAND2_X1 U8695 ( .A1(n8263), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U8696 ( .A1(n7160), .A2(n7658), .ZN(n9897) );
  NAND2_X1 U8697 ( .A1(n6625), .A2(n7161), .ZN(n7160) );
  NAND2_X1 U8698 ( .A1(n12841), .A2(n8084), .ZN(n12751) );
  NAND2_X1 U8699 ( .A1(n12841), .A2(n7167), .ZN(n12753) );
  INV_X1 U8700 ( .A(n13220), .ZN(n13081) );
  NAND2_X1 U8701 ( .A1(n10655), .A2(n7724), .ZN(n10792) );
  OR2_X1 U8702 ( .A1(n7532), .A2(n11472), .ZN(n11628) );
  INV_X1 U8703 ( .A(n6424), .ZN(n14865) );
  NAND2_X1 U8704 ( .A1(n12817), .A2(n7960), .ZN(n12786) );
  NAND2_X1 U8705 ( .A1(n7889), .A2(n11453), .ZN(n11458) );
  INV_X1 U8706 ( .A(n11462), .ZN(n6626) );
  NOR2_X1 U8707 ( .A1(n9695), .A2(n9692), .ZN(n7599) );
  AND2_X1 U8708 ( .A1(n9693), .A2(n9646), .ZN(n6699) );
  AND2_X1 U8709 ( .A1(n12784), .A2(n7982), .ZN(n12819) );
  NAND2_X1 U8710 ( .A1(n7765), .A2(n10734), .ZN(n11011) );
  AND2_X1 U8711 ( .A1(n11458), .A2(n7893), .ZN(n12833) );
  INV_X1 U8712 ( .A(n6625), .ZN(n9770) );
  INV_X1 U8713 ( .A(n10247), .ZN(n14901) );
  INV_X1 U8714 ( .A(n14494), .ZN(n12816) );
  INV_X1 U8715 ( .A(n11375), .ZN(n11287) );
  INV_X1 U8716 ( .A(n10155), .ZN(n12866) );
  INV_X1 U8717 ( .A(n11625), .ZN(n12869) );
  OAI22_X1 U8718 ( .A1(n14757), .A2(n14758), .B1(n7546), .B2(n9387), .ZN(
        n14775) );
  AOI21_X1 U8719 ( .B1(n14773), .B2(n9424), .A(n9423), .ZN(n9437) );
  INV_X1 U8720 ( .A(n6845), .ZN(n9431) );
  NOR2_X1 U8721 ( .A1(n9386), .A2(n9385), .ZN(n9555) );
  AND2_X1 U8722 ( .A1(n6845), .A2(n6844), .ZN(n9386) );
  NAND2_X1 U8723 ( .A1(n9391), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6844) );
  INV_X1 U8724 ( .A(n6843), .ZN(n9584) );
  AOI21_X1 U8725 ( .B1(n14789), .B2(n9565), .A(n9564), .ZN(n9589) );
  NAND2_X1 U8726 ( .A1(n9795), .A2(n6841), .ZN(n9796) );
  OR2_X1 U8727 ( .A1(n9799), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6841) );
  NOR2_X1 U8728 ( .A1(n9802), .A2(n9801), .ZN(n10128) );
  AOI211_X1 U8729 ( .C1(n10698), .C2(n10703), .A(n10697), .B(n10699), .ZN(
        n10863) );
  XNOR2_X1 U8730 ( .A(n11336), .B(n11335), .ZN(n11187) );
  INV_X1 U8731 ( .A(n9151), .ZN(n13183) );
  NAND2_X1 U8732 ( .A1(n7256), .A2(n7255), .ZN(n13194) );
  OAI21_X1 U8733 ( .B1(n13049), .B2(n7080), .A(n7079), .ZN(n13007) );
  NAND2_X1 U8734 ( .A1(n7084), .A2(n7081), .ZN(n13020) );
  NAND2_X1 U8735 ( .A1(n13049), .A2(n6493), .ZN(n7081) );
  OR3_X1 U8736 ( .A1(n13041), .A2(n13040), .A3(n13169), .ZN(n13206) );
  NAND2_X1 U8737 ( .A1(n7087), .A2(n7090), .ZN(n13034) );
  OR2_X1 U8738 ( .A1(n13049), .A2(n13053), .ZN(n7087) );
  OR3_X1 U8739 ( .A1(n13056), .A2(n13055), .A3(n13169), .ZN(n13212) );
  NAND2_X1 U8740 ( .A1(n7108), .A2(n12936), .ZN(n13086) );
  AND2_X1 U8741 ( .A1(n7945), .A2(n7944), .ZN(n13122) );
  NAND2_X1 U8742 ( .A1(n6880), .A2(n6484), .ZN(n13116) );
  NAND2_X1 U8743 ( .A1(n12963), .A2(n6887), .ZN(n6880) );
  NAND2_X1 U8744 ( .A1(n12963), .A2(n12962), .ZN(n13137) );
  NAND2_X1 U8745 ( .A1(n13162), .A2(n12927), .ZN(n13147) );
  OR3_X1 U8746 ( .A1(n13171), .A2(n13170), .A3(n13169), .ZN(n13252) );
  NAND2_X1 U8747 ( .A1(n7243), .A2(n7241), .ZN(n12957) );
  NAND2_X1 U8748 ( .A1(n7243), .A2(n11355), .ZN(n11356) );
  OAI21_X1 U8749 ( .B1(n11121), .B2(n6875), .A(n6872), .ZN(n11272) );
  NAND2_X1 U8750 ( .A1(n10880), .A2(n10879), .ZN(n10881) );
  AND2_X1 U8751 ( .A1(n7691), .A2(n7690), .ZN(n10470) );
  NAND2_X1 U8752 ( .A1(n10244), .A2(n10243), .ZN(n10439) );
  NAND2_X1 U8753 ( .A1(n9836), .A2(n9085), .ZN(n6620) );
  INV_X1 U8754 ( .A(n9932), .ZN(n14879) );
  OR2_X1 U8755 ( .A1(n14844), .A2(n14832), .ZN(n14824) );
  INV_X1 U8756 ( .A(n13178), .ZN(n14828) );
  INV_X1 U8757 ( .A(n14824), .ZN(n13141) );
  INV_X1 U8758 ( .A(n14819), .ZN(n14839) );
  INV_X2 U8759 ( .A(n14515), .ZN(n14844) );
  OR3_X1 U8760 ( .A1(n13223), .A2(n13222), .A3(n13221), .ZN(n13273) );
  OR2_X1 U8761 ( .A1(n13235), .A2(n13234), .ZN(n13275) );
  AND2_X2 U8762 ( .A1(n11158), .A2(n14850), .ZN(n14952) );
  AND2_X1 U8763 ( .A1(n9176), .A2(n8154), .ZN(n14854) );
  INV_X1 U8764 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n13285) );
  MUX2_X1 U8765 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7513), .S(
        P2_IR_REG_29__SCAN_IN), .Z(n7514) );
  INV_X1 U8766 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11297) );
  INV_X1 U8767 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11204) );
  INV_X1 U8768 ( .A(n6464), .ZN(n11050) );
  INV_X1 U8769 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U8770 ( .A1(n7490), .A2(n7489), .ZN(n7492) );
  NAND2_X1 U8771 ( .A1(n7488), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7489) );
  INV_X1 U8772 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n12226) );
  INV_X1 U8773 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n9645) );
  INV_X1 U8774 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n9230) );
  INV_X1 U8775 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n9231) );
  INV_X1 U8776 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n9227) );
  NAND2_X1 U8777 ( .A1(n10716), .A2(n10715), .ZN(n10813) );
  NAND2_X1 U8778 ( .A1(n10711), .A2(n10710), .ZN(n10716) );
  OAI21_X1 U8779 ( .B1(n6777), .B2(n6769), .A(n6768), .ZN(n13306) );
  AOI21_X1 U8780 ( .B1(n6770), .B2(n6776), .A(n7388), .ZN(n6768) );
  INV_X1 U8781 ( .A(n6770), .ZN(n6769) );
  NOR2_X1 U8782 ( .A1(n6490), .A2(n6771), .ZN(n6770) );
  NAND2_X1 U8783 ( .A1(n14540), .A2(n7370), .ZN(n14542) );
  AND2_X1 U8784 ( .A1(n14538), .A2(n14539), .ZN(n7370) );
  NAND2_X1 U8785 ( .A1(n9884), .A2(n9886), .ZN(n9887) );
  INV_X1 U8786 ( .A(n9885), .ZN(n9886) );
  OAI21_X1 U8787 ( .B1(n13367), .B2(n7381), .A(n7380), .ZN(n13324) );
  AND2_X1 U8788 ( .A1(n10813), .A2(n7403), .ZN(n11036) );
  NAND2_X1 U8789 ( .A1(n10813), .A2(n10812), .ZN(n10814) );
  NAND2_X1 U8790 ( .A1(n9629), .A2(n6756), .ZN(n9630) );
  NAND2_X1 U8791 ( .A1(n9628), .A2(n11853), .ZN(n9629) );
  INV_X1 U8792 ( .A(n9627), .ZN(n9628) );
  NAND2_X1 U8793 ( .A1(n13384), .A2(n11925), .ZN(n13329) );
  NAND2_X1 U8794 ( .A1(n6772), .A2(n6773), .ZN(n13349) );
  NAND2_X1 U8795 ( .A1(n13425), .A2(n11900), .ZN(n13359) );
  AND2_X1 U8796 ( .A1(n11426), .A2(n11425), .ZN(n14181) );
  NAND2_X1 U8797 ( .A1(n6777), .A2(n11944), .ZN(n13377) );
  NOR2_X1 U8798 ( .A1(n7400), .A2(n6781), .ZN(n6780) );
  INV_X1 U8799 ( .A(n11041), .ZN(n6781) );
  AND2_X1 U8800 ( .A1(n6782), .A2(n7401), .ZN(n11042) );
  NAND2_X1 U8801 ( .A1(n13322), .A2(n11921), .ZN(n13386) );
  NAND2_X1 U8802 ( .A1(n13386), .A2(n13385), .ZN(n13384) );
  NAND2_X1 U8803 ( .A1(n13340), .A2(n11879), .ZN(n13392) );
  NAND2_X1 U8804 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  AND2_X1 U8805 ( .A1(n13332), .A2(n14083), .ZN(n13418) );
  OAI21_X1 U8806 ( .B1(n11859), .B2(n7376), .A(n7373), .ZN(n14571) );
  AND2_X1 U8807 ( .A1(n13422), .A2(n14712), .ZN(n14576) );
  NAND2_X1 U8808 ( .A1(n13366), .A2(n11908), .ZN(n13408) );
  NAND2_X1 U8809 ( .A1(n10623), .A2(n10622), .ZN(n10628) );
  OR3_X1 U8810 ( .A1(n9548), .A2(n9538), .A3(n9537), .ZN(n14570) );
  XNOR2_X1 U8811 ( .A(n11899), .B(n11897), .ZN(n13427) );
  INV_X1 U8812 ( .A(n14570), .ZN(n14553) );
  INV_X1 U8813 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n12233) );
  OR2_X1 U8814 ( .A1(n6428), .A2(n9518), .ZN(n9524) );
  OR2_X1 U8815 ( .A1(n6426), .A2(n9520), .ZN(n9522) );
  OR2_X1 U8816 ( .A1(n11557), .A2(n9307), .ZN(n9521) );
  CLKBUF_X1 U8817 ( .A(n9745), .Z(n13752) );
  AOI21_X1 U8818 ( .B1(n10263), .B2(P1_REG1_REG_6__SCAN_IN), .A(n9460), .ZN(
        n9449) );
  AND2_X1 U8819 ( .A1(n9763), .A2(n9705), .ZN(n13802) );
  AOI21_X1 U8820 ( .B1(n13802), .B2(P1_REG1_REG_13__SCAN_IN), .A(n13793), .ZN(
        n10416) );
  NOR2_X1 U8821 ( .A1(n13863), .A2(n14075), .ZN(n14093) );
  AOI21_X1 U8822 ( .B1(n13895), .B2(n13879), .A(n7347), .ZN(n13881) );
  AND2_X1 U8823 ( .A1(n14111), .A2(n13878), .ZN(n7347) );
  AND2_X1 U8824 ( .A1(n13901), .A2(n13900), .ZN(n14109) );
  NAND2_X1 U8825 ( .A1(n11492), .A2(n11491), .ZN(n13943) );
  NAND2_X1 U8826 ( .A1(n14031), .A2(n7422), .ZN(n14009) );
  AND2_X1 U8827 ( .A1(n11529), .A2(n11528), .ZN(n14028) );
  INV_X1 U8828 ( .A(n14181), .ZN(n13638) );
  AND2_X1 U8829 ( .A1(n11433), .A2(n13616), .ZN(n14082) );
  NAND2_X1 U8830 ( .A1(n14195), .A2(n7430), .ZN(n11417) );
  NAND2_X1 U8831 ( .A1(n11245), .A2(n11244), .ZN(n14195) );
  NAND2_X1 U8832 ( .A1(n11223), .A2(n11222), .ZN(n14546) );
  NAND2_X1 U8833 ( .A1(n11090), .A2(n11089), .ZN(n11219) );
  NAND2_X1 U8834 ( .A1(n7414), .A2(n7418), .ZN(n11095) );
  NAND2_X1 U8835 ( .A1(n10928), .A2(n6470), .ZN(n7414) );
  NAND2_X1 U8836 ( .A1(n10840), .A2(n10839), .ZN(n10842) );
  NAND2_X1 U8837 ( .A1(n10510), .A2(n10509), .ZN(n10512) );
  NAND2_X1 U8838 ( .A1(n7354), .A2(n7355), .ZN(n10568) );
  INV_X1 U8839 ( .A(n10550), .ZN(n10298) );
  OR2_X1 U8840 ( .A1(n14673), .A2(n10258), .ZN(n14091) );
  NAND2_X1 U8841 ( .A1(n10549), .A2(n10554), .ZN(n10548) );
  NAND2_X1 U8842 ( .A1(n10261), .A2(n10260), .ZN(n10549) );
  NAND2_X1 U8843 ( .A1(n10112), .A2(n13539), .ZN(n10111) );
  NAND2_X1 U8844 ( .A1(n9831), .A2(n9830), .ZN(n10112) );
  OR2_X1 U8845 ( .A1(n14650), .A2(n9786), .ZN(n14666) );
  INV_X1 U8846 ( .A(n14091), .ZN(n14655) );
  INV_X1 U8847 ( .A(n14666), .ZN(n13994) );
  OR2_X1 U8848 ( .A1(n9745), .A2(n6434), .ZN(n9517) );
  OR2_X1 U8849 ( .A1(n10262), .A2(n13436), .ZN(n10265) );
  AND2_X2 U8850 ( .A1(n9573), .A2(n9782), .ZN(n14734) );
  AND2_X1 U8851 ( .A1(n13448), .A2(n13447), .ZN(n14206) );
  OR3_X1 U8852 ( .A1(n14145), .A2(n14144), .A3(n14143), .ZN(n14215) );
  INV_X1 U8853 ( .A(n14043), .ZN(n14228) );
  NAND2_X1 U8854 ( .A1(n10824), .A2(n10823), .ZN(n14559) );
  AOI22_X1 U8855 ( .A1(n11514), .A2(n13767), .B1(n7361), .B2(n6524), .ZN(n9675) );
  INV_X1 U8856 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n9358) );
  OR2_X1 U8857 ( .A1(n8159), .A2(n8158), .ZN(n7234) );
  NOR2_X1 U8858 ( .A1(n9296), .A2(n9297), .ZN(n6629) );
  XNOR2_X1 U8859 ( .A(n9197), .B(P1_IR_REG_26__SCAN_IN), .ZN(n14244) );
  INV_X1 U8860 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14251) );
  XNOR2_X1 U8861 ( .A(n9198), .B(P1_IR_REG_25__SCAN_IN), .ZN(n14248) );
  OAI21_X1 U8862 ( .B1(n11554), .B2(n7225), .A(n8003), .ZN(n8022) );
  NAND2_X1 U8863 ( .A1(n7295), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9287) );
  AND2_X1 U8864 ( .A1(n7293), .A2(n6573), .ZN(n7292) );
  INV_X1 U8865 ( .A(n13442), .ZN(n10954) );
  INV_X1 U8866 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n9878) );
  INV_X1 U8867 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n9766) );
  INV_X1 U8868 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n9707) );
  INV_X1 U8869 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n9552) );
  INV_X1 U8870 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n9356) );
  NAND2_X1 U8871 ( .A1(n7731), .A2(n7750), .ZN(n10821) );
  OR2_X1 U8872 ( .A1(n7730), .A2(n7729), .ZN(n7731) );
  OR2_X1 U8873 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  INV_X1 U8874 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n12253) );
  INV_X1 U8875 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n9280) );
  OR2_X1 U8876 ( .A1(n9279), .A2(n9278), .ZN(n9406) );
  INV_X1 U8877 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n9247) );
  INV_X1 U8878 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n9229) );
  NAND2_X1 U8879 ( .A1(n7611), .A2(n6706), .ZN(n7613) );
  NAND2_X1 U8880 ( .A1(n14303), .A2(n14302), .ZN(n14369) );
  XNOR2_X1 U8881 ( .A(n14296), .B(n7139), .ZN(n15153) );
  INV_X1 U8882 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7139) );
  OAI21_X1 U8883 ( .B1(n14306), .B2(n14778), .A(n15159), .ZN(n15152) );
  INV_X1 U8884 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7142) );
  INV_X1 U8885 ( .A(n14324), .ZN(n7133) );
  XNOR2_X1 U8886 ( .A(n14331), .B(n14330), .ZN(n14381) );
  NOR2_X1 U8887 ( .A1(n14335), .A2(n14334), .ZN(n6853) );
  AND2_X1 U8888 ( .A1(n14335), .A2(n14334), .ZN(n14596) );
  AND2_X1 U8889 ( .A1(n14343), .A2(n14342), .ZN(n14603) );
  NOR2_X1 U8890 ( .A1(n14354), .A2(n14353), .ZN(n14614) );
  NAND2_X1 U8891 ( .A1(n6499), .A2(n7129), .ZN(n7132) );
  CLKBUF_X2 U8892 ( .A(n12284), .Z(P3_U3897) );
  NAND2_X1 U8893 ( .A1(n6787), .A2(n6997), .ZN(n6786) );
  NAND2_X1 U8894 ( .A1(n6471), .A2(n7001), .ZN(n6996) );
  NAND2_X1 U8895 ( .A1(n6817), .A2(n6816), .ZN(P3_U3296) );
  OR2_X1 U8896 ( .A1(n11850), .A2(n11849), .ZN(n6816) );
  NAND2_X1 U8897 ( .A1(n6818), .A2(n8903), .ZN(n6817) );
  INV_X1 U8898 ( .A(n6640), .ZN(n12376) );
  OAI211_X1 U8899 ( .C1(n12366), .C2(n12367), .A(n6501), .B(n6641), .ZN(n6640)
         );
  OAI21_X1 U8900 ( .B1(n8810), .B2(n15150), .A(n6658), .ZN(P3_U3488) );
  NOR2_X1 U8901 ( .A1(n6480), .A2(n6659), .ZN(n6658) );
  AND2_X1 U8902 ( .A1(n6984), .A2(n6982), .ZN(n8810) );
  NOR2_X1 U8903 ( .A1(n15149), .A2(n8795), .ZN(n6659) );
  OAI21_X1 U8904 ( .B1(n12685), .B2(n15144), .A(n6685), .ZN(P3_U3455) );
  INV_X1 U8905 ( .A(n6686), .ZN(n6685) );
  OAI22_X1 U8906 ( .A1(n12686), .A2(n12724), .B1(n12684), .B2(n15143), .ZN(
        n6686) );
  AND2_X1 U8907 ( .A1(n10966), .A2(n7808), .ZN(n14493) );
  INV_X1 U8908 ( .A(n6690), .ZN(n12904) );
  INV_X1 U8909 ( .A(n7257), .ZN(n12990) );
  OAI21_X1 U8910 ( .B1(n13188), .B2(n13178), .A(n7258), .ZN(n7257) );
  AOI21_X1 U8911 ( .B1(n13184), .B2(n14507), .A(n12989), .ZN(n7258) );
  OR2_X1 U8912 ( .A1(n14970), .A2(n6920), .ZN(n6919) );
  NAND2_X1 U8913 ( .A1(n13267), .A2(n14970), .ZN(n6921) );
  INV_X1 U8914 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6920) );
  INV_X1 U8915 ( .A(n9235), .ZN(n9202) );
  AOI21_X1 U8916 ( .B1(n13727), .B2(n7213), .A(n7211), .ZN(n7260) );
  NAND2_X1 U8917 ( .A1(n6681), .A2(n6677), .ZN(n13859) );
  NAND2_X1 U8918 ( .A1(n13856), .A2(n13920), .ZN(n6681) );
  OR2_X1 U8919 ( .A1(n14734), .A2(n6904), .ZN(n6903) );
  NAND2_X1 U8920 ( .A1(n14207), .A2(n14734), .ZN(n6905) );
  INV_X1 U8921 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6904) );
  MUX2_X1 U8922 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14207), .S(n14729), .Z(
        P1_U3525) );
  NOR2_X1 U8923 ( .A1(n14607), .A2(n14608), .ZN(n14606) );
  INV_X1 U8924 ( .A(n14348), .ZN(n14612) );
  INV_X1 U8925 ( .A(n7127), .ZN(n7124) );
  AOI21_X1 U8926 ( .B1(n7402), .B2(n7403), .A(n11035), .ZN(n7401) );
  NAND2_X2 U8927 ( .A1(n9533), .A2(n9506), .ZN(n11853) );
  NOR2_X1 U8928 ( .A1(n9030), .A2(n9029), .ZN(n6469) );
  INV_X1 U8929 ( .A(n13493), .ZN(n7434) );
  NAND2_X1 U8930 ( .A1(n6460), .A2(n11537), .ZN(n14031) );
  INV_X1 U8931 ( .A(n7044), .ZN(n7043) );
  OAI21_X1 U8932 ( .B1(n8411), .B2(n7045), .A(n8447), .ZN(n7044) );
  OR2_X1 U8933 ( .A1(n14588), .A2(n13343), .ZN(n6470) );
  INV_X1 U8934 ( .A(n7401), .ZN(n7400) );
  AND2_X1 U8935 ( .A1(n6998), .A2(n6997), .ZN(n6471) );
  AND2_X1 U8936 ( .A1(n14608), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6472) );
  INV_X1 U8937 ( .A(n11358), .ZN(n7244) );
  NAND2_X1 U8938 ( .A1(n11502), .A2(n11501), .ZN(n13961) );
  AOI21_X1 U8939 ( .B1(n13416), .B2(n7391), .A(n6558), .ZN(n7390) );
  INV_X1 U8940 ( .A(n7390), .ZN(n7388) );
  NAND2_X1 U8941 ( .A1(n9030), .A2(n9029), .ZN(n7312) );
  INV_X1 U8942 ( .A(n7312), .ZN(n7307) );
  AND2_X1 U8943 ( .A1(n11803), .A2(n11796), .ZN(n6473) );
  INV_X1 U8944 ( .A(n13039), .ZN(n13208) );
  NAND2_X2 U8945 ( .A1(n6620), .A2(n7586), .ZN(n10177) );
  AND2_X1 U8946 ( .A1(n6788), .A2(n6535), .ZN(n6475) );
  INV_X1 U8947 ( .A(n13617), .ZN(n11244) );
  AND2_X1 U8948 ( .A1(n13604), .A2(n13610), .ZN(n13617) );
  OR2_X1 U8949 ( .A1(n7045), .A2(n7041), .ZN(n6476) );
  NAND2_X1 U8950 ( .A1(n12583), .A2(n8544), .ZN(n6477) );
  INV_X1 U8951 ( .A(n7431), .ZN(n7430) );
  NAND2_X1 U8952 ( .A1(n13487), .A2(n11246), .ZN(n7431) );
  AND2_X1 U8953 ( .A1(n6957), .A2(n6956), .ZN(n6478) );
  AND2_X1 U8954 ( .A1(n6939), .A2(n6938), .ZN(n6479) );
  XNOR2_X1 U8955 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n8349) );
  INV_X1 U8956 ( .A(n8349), .ZN(n6742) );
  INV_X1 U8957 ( .A(n11750), .ZN(n7179) );
  AND2_X1 U8958 ( .A1(n8796), .A2(n8797), .ZN(n6480) );
  AND2_X1 U8959 ( .A1(n6602), .A2(n7874), .ZN(n6481) );
  AND2_X1 U8960 ( .A1(n7027), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n6482) );
  OR2_X1 U8961 ( .A1(n8132), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n6483) );
  INV_X1 U8962 ( .A(n7026), .ZN(n7019) );
  NAND2_X1 U8963 ( .A1(n7492), .A2(n7491), .ZN(n7504) );
  INV_X1 U8964 ( .A(n7448), .ZN(n11932) );
  INV_X1 U8965 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n14265) );
  INV_X1 U8966 ( .A(n8937), .ZN(n10545) );
  NAND2_X1 U8967 ( .A1(n7549), .A2(n7548), .ZN(n8937) );
  INV_X1 U8968 ( .A(n13754), .ZN(n7362) );
  OR2_X1 U8969 ( .A1(n13244), .A2(n12964), .ZN(n6484) );
  NOR2_X1 U8970 ( .A1(n14475), .A2(n12140), .ZN(n6486) );
  NAND2_X2 U8971 ( .A1(n11998), .A2(n8223), .ZN(n8357) );
  AND2_X1 U8972 ( .A1(n6758), .A2(n6757), .ZN(n6487) );
  AND2_X1 U8973 ( .A1(n13075), .A2(n12975), .ZN(n6488) );
  OR4_X1 U8974 ( .A1(n13714), .A2(n13713), .A3(n13712), .A4(n13717), .ZN(n6489) );
  NAND2_X1 U8975 ( .A1(n11977), .A2(n11976), .ZN(n14111) );
  OR2_X1 U8976 ( .A1(n7392), .A2(n13350), .ZN(n6490) );
  AND2_X1 U8977 ( .A1(n8269), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n6491) );
  OR2_X1 U8978 ( .A1(n14527), .A2(n11122), .ZN(n6492) );
  AND2_X1 U8979 ( .A1(n7089), .A2(n7090), .ZN(n6493) );
  AND2_X1 U8980 ( .A1(n8843), .A2(n8844), .ZN(n6494) );
  INV_X1 U8981 ( .A(n6792), .ZN(n6791) );
  NAND2_X1 U8982 ( .A1(n7005), .A2(n6793), .ZN(n6792) );
  OR2_X1 U8983 ( .A1(n14360), .A2(n7130), .ZN(n6495) );
  INV_X1 U8984 ( .A(n8954), .ZN(n7345) );
  OR2_X1 U8985 ( .A1(n11949), .A2(n11948), .ZN(n6496) );
  AND2_X1 U8986 ( .A1(n7209), .A2(n8205), .ZN(n6497) );
  NOR2_X1 U8987 ( .A1(n11124), .A2(n7249), .ZN(n7248) );
  NOR2_X1 U8988 ( .A1(n8730), .A2(n11722), .ZN(n6498) );
  OR2_X1 U8989 ( .A1(n14360), .A2(n14393), .ZN(n6499) );
  OR2_X1 U8990 ( .A1(n10321), .A2(n6766), .ZN(n6500) );
  AND2_X1 U8991 ( .A1(n11751), .A2(n11750), .ZN(n12576) );
  OR2_X1 U8992 ( .A1(n12374), .A2(n15042), .ZN(n6501) );
  INV_X1 U8993 ( .A(n10003), .ZN(n6695) );
  INV_X1 U8994 ( .A(n11830), .ZN(n6970) );
  NOR2_X1 U8995 ( .A1(n11999), .A2(n6432), .ZN(n6502) );
  AND2_X1 U8996 ( .A1(n6982), .A2(n15143), .ZN(n6503) );
  INV_X1 U8997 ( .A(n14942), .ZN(n6956) );
  INV_X1 U8998 ( .A(n12980), .ZN(n12853) );
  AND2_X1 U8999 ( .A1(n8058), .A2(n8057), .ZN(n12980) );
  OR2_X1 U9000 ( .A1(n11725), .A2(n12603), .ZN(n6504) );
  AND4_X1 U9001 ( .A1(n8212), .A2(n8202), .A3(n8201), .A4(n8213), .ZN(n6505)
         );
  BUF_X2 U9002 ( .A(n6433), .Z(n9080) );
  AND2_X1 U9003 ( .A1(n12818), .A2(n7997), .ZN(n6506) );
  AND2_X1 U9004 ( .A1(n8311), .A2(n8294), .ZN(n6507) );
  OR2_X1 U9005 ( .A1(n14104), .A2(n14103), .ZN(n6508) );
  AND2_X1 U9006 ( .A1(n13563), .A2(n10712), .ZN(n6509) );
  INV_X1 U9007 ( .A(n12749), .ZN(n6649) );
  NOR2_X1 U9008 ( .A1(n10815), .A2(n7404), .ZN(n7403) );
  OR3_X1 U9009 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6510) );
  AND2_X1 U9010 ( .A1(n13028), .A2(n12941), .ZN(n6511) );
  INV_X1 U9011 ( .A(n14742), .ZN(n9372) );
  AND2_X1 U9012 ( .A1(n8069), .A2(n8068), .ZN(n13028) );
  AND2_X1 U9013 ( .A1(n13258), .A2(n12956), .ZN(n6512) );
  AND2_X1 U9014 ( .A1(n6890), .A2(n10246), .ZN(n6513) );
  AND2_X1 U9015 ( .A1(n7355), .A2(n6902), .ZN(n6514) );
  AND2_X1 U9016 ( .A1(n7158), .A2(n7155), .ZN(n6515) );
  AND2_X1 U9017 ( .A1(n13196), .A2(n12985), .ZN(n6516) );
  AND2_X1 U9018 ( .A1(n12447), .A2(n11834), .ZN(n6517) );
  AND2_X1 U9019 ( .A1(n13155), .A2(n12928), .ZN(n6518) );
  AND2_X1 U9020 ( .A1(n11928), .A2(n11927), .ZN(n6519) );
  AND2_X1 U9021 ( .A1(n7680), .A2(n7679), .ZN(n6520) );
  AND2_X1 U9022 ( .A1(n11697), .A2(n11804), .ZN(n6521) );
  INV_X1 U9023 ( .A(n11836), .ZN(n6667) );
  AND2_X1 U9024 ( .A1(n12431), .A2(n6517), .ZN(n6522) );
  INV_X1 U9025 ( .A(n6882), .ZN(n6881) );
  OAI21_X1 U9026 ( .B1(n12966), .B2(n6883), .A(n12968), .ZN(n6882) );
  INV_X1 U9027 ( .A(n14257), .ZN(n7137) );
  INV_X1 U9028 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n10377) );
  AND2_X1 U9029 ( .A1(n11553), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6523) );
  AND2_X1 U9030 ( .A1(n11553), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n6524) );
  AND2_X1 U9031 ( .A1(n8036), .A2(n8035), .ZN(n12977) );
  AND2_X1 U9032 ( .A1(n6984), .A2(n6987), .ZN(n6525) );
  OR2_X1 U9033 ( .A1(n14264), .A2(n14265), .ZN(n6526) );
  INV_X1 U9034 ( .A(n10157), .ZN(n7116) );
  AND2_X1 U9035 ( .A1(n7775), .A2(n7774), .ZN(n14527) );
  AND2_X1 U9036 ( .A1(n13897), .A2(n7425), .ZN(n6527) );
  AND2_X1 U9037 ( .A1(n7902), .A2(n7901), .ZN(n13155) );
  INV_X1 U9038 ( .A(n13607), .ZN(n14582) );
  NAND2_X1 U9039 ( .A1(n11093), .A2(n11092), .ZN(n13607) );
  AND2_X1 U9040 ( .A1(n14031), .A2(n11538), .ZN(n6528) );
  NAND2_X1 U9041 ( .A1(n13055), .A2(n6951), .ZN(n6955) );
  AND2_X1 U9042 ( .A1(n14942), .A2(n11112), .ZN(n6529) );
  INV_X1 U9043 ( .A(n7363), .ZN(n13997) );
  NAND2_X1 U9044 ( .A1(n14253), .A2(n7361), .ZN(n7363) );
  AND2_X1 U9045 ( .A1(n13384), .A2(n7396), .ZN(n6530) );
  AND2_X1 U9046 ( .A1(n11152), .A2(n12858), .ZN(n6531) );
  AND2_X1 U9047 ( .A1(n14353), .A2(n6865), .ZN(n6532) );
  AND2_X1 U9048 ( .A1(n7171), .A2(n7960), .ZN(n6533) );
  AND2_X1 U9049 ( .A1(n10124), .A2(n9883), .ZN(n6534) );
  OR2_X1 U9050 ( .A1(n6792), .A2(n6795), .ZN(n6535) );
  INV_X1 U9051 ( .A(n6776), .ZN(n6775) );
  NAND2_X1 U9052 ( .A1(n6496), .A2(n11944), .ZN(n6776) );
  OR2_X1 U9053 ( .A1(n7339), .A2(n7340), .ZN(n6536) );
  AND2_X1 U9054 ( .A1(n8284), .A2(n8283), .ZN(n6537) );
  AND2_X1 U9055 ( .A1(n8459), .A2(n8460), .ZN(n6538) );
  XOR2_X1 U9056 ( .A(n6744), .B(n12363), .Z(n6539) );
  NAND2_X1 U9057 ( .A1(n6502), .A2(n8894), .ZN(n6540) );
  INV_X1 U9058 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n8208) );
  OR2_X1 U9059 ( .A1(n10396), .A2(n10395), .ZN(n6541) );
  AND4_X1 U9060 ( .A1(n8839), .A2(n8837), .A3(n10955), .A4(n8836), .ZN(n6542)
         );
  OR2_X1 U9061 ( .A1(n9624), .A2(n9625), .ZN(n6758) );
  NOR2_X1 U9062 ( .A1(n13612), .A2(n14086), .ZN(n6543) );
  NOR2_X1 U9063 ( .A1(n13601), .A2(n13740), .ZN(n6544) );
  NOR2_X1 U9064 ( .A1(n13607), .A2(n14536), .ZN(n6545) );
  NOR2_X1 U9065 ( .A1(n13155), .A2(n12928), .ZN(n6546) );
  NOR2_X1 U9066 ( .A1(n11873), .A2(n11872), .ZN(n6547) );
  OR2_X1 U9067 ( .A1(n14413), .A2(n12320), .ZN(n6548) );
  XOR2_X1 U9068 ( .A(n14403), .B(n14402), .Z(n6549) );
  AND2_X1 U9069 ( .A1(n11776), .A2(n12470), .ZN(n6550) );
  AND2_X1 U9070 ( .A1(n10747), .A2(n10984), .ZN(n6551) );
  NAND2_X1 U9071 ( .A1(n13439), .A2(n13438), .ZN(n13862) );
  INV_X1 U9072 ( .A(n13862), .ZN(n7236) );
  AND2_X1 U9073 ( .A1(n12505), .A2(n12139), .ZN(n6552) );
  AND2_X1 U9074 ( .A1(n6964), .A2(n6486), .ZN(n6553) );
  INV_X1 U9075 ( .A(n7428), .ZN(n7427) );
  NOR2_X1 U9076 ( .A1(n13417), .A2(n13310), .ZN(n7428) );
  OR2_X1 U9077 ( .A1(n6695), .A2(n9984), .ZN(n6554) );
  AND2_X1 U9078 ( .A1(n13202), .A2(n12983), .ZN(n6555) );
  INV_X1 U9079 ( .A(n6952), .ZN(n6951) );
  NAND2_X1 U9080 ( .A1(n6953), .A2(n6954), .ZN(n6952) );
  INV_X1 U9081 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n8765) );
  INV_X1 U9082 ( .A(n7154), .ZN(n7153) );
  NAND2_X1 U9083 ( .A1(n12832), .A2(n7893), .ZN(n7154) );
  NOR2_X1 U9084 ( .A1(n11778), .A2(n11777), .ZN(n6556) );
  AND2_X1 U9085 ( .A1(n12233), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6557) );
  AND2_X1 U9086 ( .A1(n11965), .A2(n11964), .ZN(n6558) );
  AND2_X1 U9087 ( .A1(n7767), .A2(n9260), .ZN(n6559) );
  AND2_X1 U9088 ( .A1(n9552), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n6560) );
  AND2_X1 U9089 ( .A1(n9231), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n6561) );
  OR2_X1 U9090 ( .A1(n7342), .A2(n9006), .ZN(n6562) );
  OR2_X1 U9091 ( .A1(n6490), .A2(n7389), .ZN(n6563) );
  NOR2_X1 U9092 ( .A1(n13877), .A2(n13903), .ZN(n6564) );
  AND2_X1 U9093 ( .A1(n11974), .A2(n11973), .ZN(n6565) );
  AND2_X1 U9094 ( .A1(n7880), .A2(n7879), .ZN(n13174) );
  INV_X1 U9095 ( .A(n13174), .ZN(n13255) );
  INV_X1 U9096 ( .A(n14033), .ZN(n11537) );
  INV_X1 U9097 ( .A(n6767), .ZN(n6766) );
  INV_X1 U9098 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7013) );
  AND3_X1 U9099 ( .A1(n9291), .A2(n9292), .A3(n9293), .ZN(n6566) );
  OR2_X1 U9100 ( .A1(n9037), .A2(n9039), .ZN(n6567) );
  OR2_X1 U9101 ( .A1(n7345), .A2(n8953), .ZN(n6568) );
  OR2_X1 U9102 ( .A1(n12422), .A2(n12433), .ZN(n11797) );
  OR2_X1 U9103 ( .A1(n7327), .A2(n9038), .ZN(n6569) );
  INV_X1 U9104 ( .A(n13479), .ZN(n10511) );
  OR2_X1 U9105 ( .A1(n14310), .A2(n14309), .ZN(n6570) );
  OR2_X1 U9106 ( .A1(n14320), .A2(n14319), .ZN(n6571) );
  AND2_X1 U9107 ( .A1(n13652), .A2(n13650), .ZN(n6572) );
  AND3_X1 U9108 ( .A1(n9286), .A2(n9285), .A3(n9284), .ZN(n6573) );
  NAND2_X1 U9109 ( .A1(n6863), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14257) );
  AND2_X1 U9110 ( .A1(n13617), .A2(n13739), .ZN(n6574) );
  AND2_X1 U9111 ( .A1(n7371), .A2(n6778), .ZN(n6575) );
  INV_X1 U9112 ( .A(n9004), .ZN(n7342) );
  AND2_X1 U9113 ( .A1(n12937), .A2(n7103), .ZN(n6576) );
  AND3_X1 U9114 ( .A1(n7467), .A2(n7466), .A3(n7465), .ZN(n7507) );
  NOR2_X1 U9115 ( .A1(n12922), .A2(n7242), .ZN(n7241) );
  OR2_X1 U9116 ( .A1(n11953), .A2(n13953), .ZN(n6577) );
  NOR2_X1 U9117 ( .A1(n7275), .A2(n7273), .ZN(n6578) );
  INV_X1 U9118 ( .A(n10878), .ZN(n10882) );
  AND2_X1 U9119 ( .A1(n6497), .A2(n8208), .ZN(n6579) );
  OR2_X1 U9120 ( .A1(n7291), .A2(n13554), .ZN(n6580) );
  AND2_X1 U9121 ( .A1(n6871), .A2(n11271), .ZN(n6581) );
  AND2_X1 U9122 ( .A1(n13697), .A2(n7266), .ZN(n6582) );
  AND2_X1 U9123 ( .A1(n7264), .A2(n13696), .ZN(n6583) );
  AND2_X1 U9124 ( .A1(n6471), .A2(n6540), .ZN(n6584) );
  INV_X1 U9125 ( .A(n11800), .ZN(n12403) );
  AND2_X1 U9126 ( .A1(n7276), .A2(n13661), .ZN(n6585) );
  AND2_X1 U9127 ( .A1(n6763), .A2(n6760), .ZN(n6586) );
  INV_X1 U9128 ( .A(n7442), .ZN(n7385) );
  NAND2_X1 U9129 ( .A1(n7280), .A2(n13603), .ZN(n6587) );
  NAND2_X1 U9130 ( .A1(n13701), .A2(n7271), .ZN(n6588) );
  AND2_X1 U9131 ( .A1(n6478), .A2(n14527), .ZN(n6589) );
  INV_X1 U9132 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n7314) );
  NAND2_X1 U9133 ( .A1(n13196), .A2(n12942), .ZN(n6590) );
  INV_X1 U9134 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n9289) );
  NAND2_X1 U9135 ( .A1(n8892), .A2(n12433), .ZN(n7005) );
  INV_X1 U9136 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7037) );
  NOR2_X1 U9137 ( .A1(n13737), .A2(n6466), .ZN(n6592) );
  AND2_X2 U9138 ( .A1(n7502), .A2(n7501), .ZN(n12903) );
  OAI21_X1 U9139 ( .B1(n11383), .B2(n6486), .A(n6964), .ZN(n12551) );
  AND2_X1 U9140 ( .A1(n7925), .A2(n7924), .ZN(n13244) );
  INV_X1 U9141 ( .A(n13244), .ZN(n6949) );
  NAND2_X1 U9142 ( .A1(n11458), .A2(n7153), .ZN(n12769) );
  NAND2_X1 U9143 ( .A1(n12872), .A2(n14831), .ZN(n9136) );
  NAND2_X1 U9144 ( .A1(n11119), .A2(n11118), .ZN(n11121) );
  INV_X1 U9145 ( .A(n7054), .ZN(n7053) );
  OAI21_X1 U9146 ( .B1(n8500), .B2(n7055), .A(n8526), .ZN(n7054) );
  INV_X1 U9147 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6935) );
  XNOR2_X1 U9148 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n8327) );
  INV_X1 U9149 ( .A(n8327), .ZN(n6739) );
  XOR2_X1 U9150 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .Z(n6593) );
  INV_X1 U9151 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7040) );
  INV_X1 U9152 ( .A(n13196), .ZN(n6953) );
  INV_X1 U9153 ( .A(n14008), .ZN(n7423) );
  INV_X1 U9154 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n6622) );
  INV_X1 U9155 ( .A(n11745), .ZN(n7180) );
  OR2_X1 U9156 ( .A1(n8884), .A2(n12471), .ZN(n6594) );
  INV_X1 U9157 ( .A(n8381), .ZN(n6730) );
  XNOR2_X1 U9158 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n8381) );
  OR2_X1 U9159 ( .A1(n12332), .A2(n8404), .ZN(n6595) );
  AND2_X1 U9160 ( .A1(n14195), .A2(n11246), .ZN(n6596) );
  INV_X1 U9161 ( .A(n7550), .ZN(n7587) );
  OR2_X1 U9162 ( .A1(n11907), .A2(n11906), .ZN(n11908) );
  AND2_X1 U9163 ( .A1(n10880), .A2(n7120), .ZN(n6597) );
  AND2_X1 U9164 ( .A1(n8887), .A2(n7452), .ZN(n6598) );
  OR2_X1 U9165 ( .A1(n6716), .A2(P3_IR_REG_14__SCAN_IN), .ZN(n6599) );
  OR2_X1 U9166 ( .A1(n7918), .A2(n12267), .ZN(n6600) );
  AND2_X1 U9167 ( .A1(n9878), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n6601) );
  NAND2_X1 U9168 ( .A1(n7895), .A2(n9653), .ZN(n6602) );
  INV_X1 U9169 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10180) );
  AND2_X1 U9170 ( .A1(n11224), .A2(n13610), .ZN(n6603) );
  INV_X1 U9171 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n6723) );
  AND2_X1 U9172 ( .A1(n6600), .A2(n7897), .ZN(n6604) );
  NOR2_X1 U9173 ( .A1(n15113), .A2(n11848), .ZN(n6605) );
  INV_X1 U9174 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6752) );
  INV_X1 U9175 ( .A(n11453), .ZN(n7152) );
  AND2_X1 U9176 ( .A1(n10479), .A2(n6478), .ZN(n6606) );
  NAND2_X1 U9177 ( .A1(n12317), .A2(n15024), .ZN(n7026) );
  AND2_X1 U9178 ( .A1(n11096), .A2(n6941), .ZN(n6607) );
  AND2_X1 U9179 ( .A1(n14998), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n6608) );
  XOR2_X1 U9180 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .Z(n6609) );
  NAND2_X1 U9181 ( .A1(n10327), .A2(n6759), .ZN(n10621) );
  NAND2_X1 U9182 ( .A1(n11420), .A2(n11419), .ZN(n14188) );
  INV_X1 U9183 ( .A(n14188), .ZN(n6938) );
  INV_X1 U9184 ( .A(n11827), .ZN(n7189) );
  NAND2_X1 U9185 ( .A1(n7356), .A2(n10283), .ZN(n10507) );
  AND2_X1 U9186 ( .A1(n6889), .A2(n6890), .ZN(n6610) );
  AND2_X1 U9187 ( .A1(n10728), .A2(n8338), .ZN(n6611) );
  AND2_X1 U9188 ( .A1(n7115), .A2(n10159), .ZN(n6612) );
  NAND2_X1 U9189 ( .A1(n11204), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6613) );
  AND2_X1 U9190 ( .A1(n9057), .A2(n12739), .ZN(n6614) );
  INV_X1 U9191 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10457) );
  INV_X1 U9192 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10380) );
  INV_X1 U9193 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11051) );
  NOR2_X1 U9194 ( .A1(n9054), .A2(n7233), .ZN(n7232) );
  OAI21_X1 U9195 ( .B1(n7022), .B2(n7026), .A(n6482), .ZN(n7020) );
  INV_X1 U9196 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7070) );
  NAND4_X2 U9197 ( .A1(n9638), .A2(n9637), .A3(n9636), .A4(n9635), .ZN(n13749)
         );
  INV_X1 U9198 ( .A(n12134), .ZN(n6997) );
  INV_X1 U9199 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14245) );
  INV_X1 U9200 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13294) );
  INV_X1 U9201 ( .A(n14817), .ZN(n6944) );
  NAND2_X1 U9202 ( .A1(n8895), .A2(n8918), .ZN(n12134) );
  AND2_X1 U9203 ( .A1(n14804), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6615) );
  AND2_X1 U9204 ( .A1(n8809), .A2(n8808), .ZN(n15144) );
  OR2_X1 U9205 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7070), .ZN(n6616) );
  AND2_X1 U9206 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n7070), .ZN(n6617) );
  AND2_X1 U9207 ( .A1(n12903), .A2(n6485), .ZN(n9913) );
  INV_X1 U9208 ( .A(n12349), .ZN(n6698) );
  INV_X1 U9209 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n7017) );
  INV_X1 U9210 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6693) );
  INV_X1 U9211 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6710) );
  INV_X1 U9212 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7046) );
  INV_X1 U9213 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n6624) );
  INV_X1 U9214 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6840) );
  INV_X1 U9215 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7140) );
  INV_X1 U9216 ( .A(n13680), .ZN(n6619) );
  NAND2_X1 U9217 ( .A1(n9195), .A2(n7435), .ZN(n9357) );
  NOR2_X1 U9218 ( .A1(n6630), .A2(n6629), .ZN(n6628) );
  OAI21_X1 U9219 ( .B1(n13693), .B2(n7268), .A(n6582), .ZN(n13698) );
  OR2_X1 U9220 ( .A1(n15154), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n6852) );
  NAND2_X1 U9221 ( .A1(n14373), .A2(n14372), .ZN(n7141) );
  NAND3_X1 U9222 ( .A1(n6855), .A2(n6858), .A3(n6859), .ZN(n14295) );
  NOR2_X1 U9223 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(n14392), .ZN(n14360) );
  NOR2_X1 U9224 ( .A1(n14343), .A2(n14342), .ZN(n14604) );
  XNOR2_X1 U9225 ( .A(n14299), .B(n14257), .ZN(n14301) );
  NAND2_X1 U9226 ( .A1(n15153), .A2(n15152), .ZN(n6631) );
  NAND2_X1 U9227 ( .A1(n14325), .A2(n14326), .ZN(n14331) );
  AOI21_X1 U9228 ( .B1(n14601), .B2(n14339), .A(n14598), .ZN(n14343) );
  XNOR2_X1 U9229 ( .A(n14319), .B(n14320), .ZN(n14374) );
  XNOR2_X1 U9230 ( .A(n7844), .B(n7845), .ZN(n11281) );
  NAND2_X2 U9231 ( .A1(n7173), .A2(n7807), .ZN(n10966) );
  OAI21_X2 U9232 ( .B1(n11592), .B2(n11591), .A(n11590), .ZN(n14057) );
  OR2_X1 U9233 ( .A1(n10267), .A2(n9066), .ZN(n7671) );
  NAND2_X1 U9234 ( .A1(n9746), .A2(n13529), .ZN(n9747) );
  NAND2_X2 U9235 ( .A1(n7162), .A2(n7157), .ZN(n7156) );
  NAND2_X1 U9236 ( .A1(n11088), .A2(n11087), .ZN(n11090) );
  NAND2_X1 U9237 ( .A1(n9852), .A2(n13536), .ZN(n10115) );
  OAI21_X1 U9238 ( .B1(n14192), .B2(n14106), .A(n6664), .ZN(n14207) );
  NAND2_X1 U9239 ( .A1(n8993), .A2(n8994), .ZN(n8992) );
  NAND2_X1 U9240 ( .A1(n9014), .A2(n9013), .ZN(n9015) );
  NOR2_X1 U9241 ( .A1(n8930), .A2(n8929), .ZN(n8934) );
  NOR2_X1 U9242 ( .A1(n8960), .A2(n8959), .ZN(n8964) );
  INV_X1 U9243 ( .A(n13072), .ZN(n6621) );
  NAND2_X2 U9244 ( .A1(n7524), .A2(n9617), .ZN(n7943) );
  AND2_X4 U9245 ( .A1(n9913), .A2(n11202), .ZN(n9091) );
  NAND2_X1 U9246 ( .A1(n9924), .A2(n9923), .ZN(n10169) );
  NAND2_X1 U9247 ( .A1(n12991), .A2(n12987), .ZN(n7259) );
  INV_X1 U9248 ( .A(n8990), .ZN(n6651) );
  NAND2_X1 U9249 ( .A1(n6921), .A2(n6919), .ZN(P2_U3528) );
  NAND2_X1 U9250 ( .A1(n7253), .A2(n7254), .ZN(n12992) );
  NAND2_X1 U9251 ( .A1(n12090), .A2(n12089), .ZN(n12088) );
  MUX2_X1 U9252 ( .A(n11686), .B(n8818), .S(n8852), .Z(n10205) );
  OAI21_X2 U9253 ( .B1(n11301), .B2(n7011), .A(n11299), .ZN(n12008) );
  NAND2_X2 U9254 ( .A1(n11998), .A2(n12736), .ZN(n11655) );
  XNOR2_X2 U9255 ( .A(n8217), .B(n6624), .ZN(n11998) );
  AOI21_X2 U9256 ( .B1(n11164), .B2(n8851), .A(n8850), .ZN(n11255) );
  NAND2_X1 U9257 ( .A1(n6798), .A2(n8864), .ZN(n12059) );
  NAND2_X1 U9258 ( .A1(n9747), .A2(n13533), .ZN(n9852) );
  NAND2_X1 U9259 ( .A1(n10115), .A2(n13470), .ZN(n10114) );
  NAND2_X1 U9260 ( .A1(n10936), .A2(n10935), .ZN(n11088) );
  NAND2_X1 U9261 ( .A1(n6665), .A2(n13530), .ZN(n9746) );
  NAND2_X1 U9262 ( .A1(n11254), .A2(n8856), .ZN(n11301) );
  NAND2_X1 U9263 ( .A1(n11224), .A2(n6913), .ZN(n11433) );
  AOI21_X1 U9264 ( .B1(n9157), .B2(n9156), .A(n9155), .ZN(n9166) );
  NAND2_X1 U9265 ( .A1(n10114), .A2(n13543), .ZN(n9853) );
  NAND2_X1 U9266 ( .A1(n12125), .A2(n8862), .ZN(n6798) );
  INV_X1 U9267 ( .A(n9745), .ZN(n6666) );
  NAND4_X1 U9268 ( .A1(n9514), .A2(n9512), .A3(n9511), .A4(n9513), .ZN(n9745)
         );
  INV_X1 U9269 ( .A(n13527), .ZN(n6665) );
  NAND2_X1 U9270 ( .A1(n6898), .A2(n6897), .ZN(n13895) );
  OAI21_X2 U9271 ( .B1(n13988), .B2(n13996), .A(n11597), .ZN(n13980) );
  XNOR2_X1 U9272 ( .A(n13881), .B(n13880), .ZN(n14105) );
  OAI21_X1 U9273 ( .B1(n9212), .B2(n6935), .A(n6934), .ZN(n7476) );
  XNOR2_X2 U9274 ( .A(n8019), .B(n8017), .ZN(n12759) );
  NAND2_X1 U9275 ( .A1(n12773), .A2(n7938), .ZN(n7956) );
  NAND2_X2 U9276 ( .A1(n6627), .A2(n6626), .ZN(n11459) );
  INV_X1 U9277 ( .A(n11461), .ZN(n6627) );
  NAND2_X1 U9278 ( .A1(n9696), .A2(n7601), .ZN(n9755) );
  NAND2_X1 U9279 ( .A1(n7698), .A2(n7697), .ZN(n7726) );
  NAND2_X1 U9280 ( .A1(n7226), .A2(n7542), .ZN(n7568) );
  NAND2_X1 U9281 ( .A1(n6632), .A2(n7919), .ZN(n7940) );
  AND2_X4 U9282 ( .A1(n7366), .A2(n7365), .ZN(n9195) );
  OR2_X1 U9283 ( .A1(n9618), .A2(n13436), .ZN(n9621) );
  NAND2_X1 U9284 ( .A1(n10847), .A2(n10846), .ZN(n10918) );
  NAND2_X1 U9285 ( .A1(n10278), .A2(n10284), .ZN(n10486) );
  NAND2_X1 U9286 ( .A1(n6905), .A2(n6903), .ZN(P1_U3557) );
  NAND2_X2 U9287 ( .A1(n9299), .A2(n14619), .ZN(n7364) );
  NAND2_X2 U9288 ( .A1(n9295), .A2(n6628), .ZN(n14619) );
  NAND2_X1 U9289 ( .A1(n7229), .A2(n6604), .ZN(n6632) );
  XNOR2_X1 U9290 ( .A(n6633), .B(n6549), .ZN(SUB_1596_U4) );
  NAND2_X1 U9291 ( .A1(n7125), .A2(n7132), .ZN(n6633) );
  NAND2_X1 U9292 ( .A1(n8819), .A2(n10205), .ZN(n10204) );
  NOR2_X1 U9293 ( .A1(n14603), .A2(P2_ADDR_REG_13__SCAN_IN), .ZN(n14344) );
  NAND2_X4 U9294 ( .A1(n14936), .A2(n9128), .ZN(n8119) );
  NAND2_X1 U9295 ( .A1(n8000), .A2(n7999), .ZN(n8019) );
  NAND3_X1 U9296 ( .A1(n7300), .A2(n8947), .A3(n7299), .ZN(n7298) );
  NAND2_X1 U9297 ( .A1(n8941), .A2(n8940), .ZN(n7300) );
  INV_X4 U9298 ( .A(n7943), .ZN(n8026) );
  NAND2_X1 U9299 ( .A1(n14408), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n14407) );
  NAND2_X1 U9300 ( .A1(n10766), .A2(n10767), .ZN(n12331) );
  OAI211_X1 U9301 ( .C1(n7261), .C2(n13730), .A(n6644), .B(n7260), .ZN(
        P1_U3242) );
  NAND2_X1 U9302 ( .A1(n7261), .A2(n13723), .ZN(n6644) );
  NAND2_X1 U9303 ( .A1(n13668), .A2(n13669), .ZN(n13671) );
  NAND2_X1 U9304 ( .A1(n6645), .A2(n7270), .ZN(n13706) );
  NAND3_X1 U9305 ( .A1(n13698), .A2(n13699), .A3(n6588), .ZN(n6645) );
  INV_X1 U9306 ( .A(n10460), .ZN(n7405) );
  NAND2_X1 U9307 ( .A1(n10726), .A2(n11700), .ZN(n10978) );
  NAND2_X1 U9308 ( .A1(n10527), .A2(n8824), .ZN(n10528) );
  NAND2_X1 U9309 ( .A1(n8740), .A2(n8739), .ZN(n12545) );
  NAND2_X1 U9310 ( .A1(n12283), .A2(n15094), .ZN(n11693) );
  NAND2_X1 U9311 ( .A1(n8983), .A2(n8982), .ZN(n6654) );
  AND2_X1 U9312 ( .A1(n7324), .A2(n7325), .ZN(n9025) );
  NAND2_X1 U9313 ( .A1(n6655), .A2(n6654), .ZN(n6653) );
  OAI22_X1 U9314 ( .A1(n7341), .A2(n9003), .B1(n9005), .B2(n9004), .ZN(n9009)
         );
  NAND2_X1 U9315 ( .A1(n8985), .A2(n8984), .ZN(n6655) );
  INV_X1 U9316 ( .A(n6653), .ZN(n8989) );
  NAND2_X1 U9317 ( .A1(n6656), .A2(n6569), .ZN(n9042) );
  INV_X1 U9318 ( .A(n9036), .ZN(n6657) );
  NAND3_X1 U9319 ( .A1(n6657), .A2(n6567), .A3(n7326), .ZN(n6656) );
  AOI21_X1 U9320 ( .B1(n13352), .B2(n11616), .A(n6423), .ZN(n13939) );
  NAND2_X1 U9321 ( .A1(n12760), .A2(n8020), .ZN(n12802) );
  AND2_X2 U9322 ( .A1(n9754), .A2(n7632), .ZN(n7162) );
  XNOR2_X1 U9323 ( .A(n11647), .B(n6667), .ZN(n12381) );
  NOR2_X1 U9324 ( .A1(n7438), .A2(n6983), .ZN(n6982) );
  AOI21_X1 U9325 ( .B1(n7639), .B2(n7638), .A(n7637), .ZN(n7643) );
  AND3_X1 U9326 ( .A1(n7297), .A2(n7298), .A3(n7296), .ZN(n8950) );
  INV_X1 U9327 ( .A(n9035), .ZN(n6662) );
  INV_X4 U9328 ( .A(n7587), .ZN(n9073) );
  OAI21_X2 U9329 ( .B1(n7660), .B2(n6918), .A(n6915), .ZN(n7686) );
  OAI21_X1 U9330 ( .B1(n8977), .B2(n8976), .A(n8975), .ZN(n8979) );
  NAND2_X1 U9331 ( .A1(n9712), .A2(n9711), .ZN(n9739) );
  OAI21_X1 U9332 ( .B1(n14298), .B2(n14297), .A(n7135), .ZN(n7134) );
  NAND2_X1 U9333 ( .A1(n9854), .A2(n9853), .ZN(n7346) );
  NAND2_X1 U9334 ( .A1(n14023), .A2(n11594), .ZN(n14004) );
  NAND2_X1 U9335 ( .A1(n6666), .A2(n6434), .ZN(n13527) );
  OAI21_X1 U9336 ( .B1(n8933), .B2(n8934), .A(n8932), .ZN(n8936) );
  NAND2_X1 U9337 ( .A1(n9126), .A2(n9125), .ZN(n9162) );
  AOI21_X1 U9338 ( .B1(n9035), .B2(n9034), .A(n9033), .ZN(n9036) );
  OAI21_X1 U9339 ( .B1(n8964), .B2(n8963), .A(n8962), .ZN(n8966) );
  NAND3_X1 U9340 ( .A1(n8952), .A2(n8951), .A3(n6568), .ZN(n7343) );
  NAND2_X1 U9341 ( .A1(n8945), .A2(n8944), .ZN(n7299) );
  INV_X1 U9342 ( .A(n8971), .ZN(n7338) );
  OAI211_X1 U9343 ( .C1(n9015), .C2(n7323), .A(n7316), .B(n9019), .ZN(n7324)
         );
  NAND2_X1 U9344 ( .A1(n13187), .A2(n6672), .ZN(n13267) );
  NAND2_X1 U9345 ( .A1(n7791), .A2(n7790), .ZN(n7810) );
  NAND2_X1 U9346 ( .A1(n7600), .A2(n7599), .ZN(n9696) );
  NAND2_X1 U9347 ( .A1(n6943), .A2(n13417), .ZN(n11617) );
  NAND2_X1 U9348 ( .A1(n14491), .A2(n7826), .ZN(n7844) );
  NAND2_X1 U9349 ( .A1(n7566), .A2(n7565), .ZN(n7575) );
  INV_X1 U9350 ( .A(n8766), .ZN(n8768) );
  OAI211_X1 U9351 ( .C1(n13049), .C2(n7077), .A(n7076), .B(n6590), .ZN(n6696)
         );
  NAND2_X1 U9352 ( .A1(n6911), .A2(n14033), .ZN(n14023) );
  NAND2_X1 U9353 ( .A1(n7538), .A2(n7537), .ZN(n7226) );
  NAND2_X1 U9354 ( .A1(n14036), .A2(n13659), .ZN(n14019) );
  NAND2_X1 U9355 ( .A1(n10555), .A2(n7357), .ZN(n7354) );
  INV_X1 U9356 ( .A(n6910), .ZN(n13933) );
  NAND2_X1 U9357 ( .A1(n9579), .A2(n9580), .ZN(n9647) );
  AOI21_X2 U9358 ( .B1(n10647), .B2(n10646), .A(n6715), .ZN(n7720) );
  NAND2_X1 U9359 ( .A1(n11011), .A2(n6689), .ZN(n11021) );
  NAND2_X1 U9360 ( .A1(n9755), .A2(n9756), .ZN(n9754) );
  NAND2_X2 U9361 ( .A1(n10655), .A2(n7174), .ZN(n10790) );
  NAND2_X1 U9362 ( .A1(n11021), .A2(n7786), .ZN(n10965) );
  NAND2_X1 U9363 ( .A1(n7333), .A2(n7330), .ZN(n7329) );
  NAND2_X2 U9364 ( .A1(n7156), .A2(n7158), .ZN(n10647) );
  NAND2_X1 U9365 ( .A1(n6889), .A2(n6513), .ZN(n10464) );
  NAND2_X1 U9366 ( .A1(n7239), .A2(n7240), .ZN(n13161) );
  NOR2_X2 U9367 ( .A1(n7814), .A2(n7508), .ZN(n7511) );
  INV_X1 U9368 ( .A(n6876), .ZN(n13091) );
  NOR2_X1 U9369 ( .A1(n10169), .A2(n6869), .ZN(n6866) );
  INV_X1 U9370 ( .A(n9830), .ZN(n7411) );
  OR2_X1 U9371 ( .A1(n9674), .A2(n13436), .ZN(n9676) );
  INV_X4 U9372 ( .A(n8852), .ZN(n10202) );
  NAND2_X1 U9373 ( .A1(n14607), .A2(n7148), .ZN(n6862) );
  NOR2_X1 U9374 ( .A1(n6853), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n14336) );
  NOR2_X2 U9375 ( .A1(n10034), .A2(n9274), .ZN(n7366) );
  NAND4_X1 U9376 ( .A1(n9180), .A2(n9178), .A3(n9179), .A4(n9874), .ZN(n10034)
         );
  NAND2_X1 U9377 ( .A1(n6687), .A2(n13670), .ZN(n13674) );
  NAND2_X1 U9378 ( .A1(n13671), .A2(n13672), .ZN(n6687) );
  OR2_X2 U9379 ( .A1(n13560), .A2(n13559), .ZN(n13561) );
  OAI22_X2 U9380 ( .A1(n13575), .A2(n7287), .B1(n13574), .B2(n7286), .ZN(
        n13579) );
  NAND2_X1 U9381 ( .A1(n7265), .A2(n6583), .ZN(n13695) );
  INV_X1 U9382 ( .A(n6720), .ZN(n13668) );
  NAND2_X1 U9383 ( .A1(n11191), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n11192) );
  BUF_X1 U9384 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n14739) );
  XNOR2_X2 U9385 ( .A(n7473), .B(P2_IR_REG_1__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U9386 ( .A1(n7460), .A2(n7771), .ZN(n7814) );
  INV_X1 U9387 ( .A(n6696), .ZN(n12993) );
  NOR2_X1 U9388 ( .A1(n9979), .A2(n6694), .ZN(n9978) );
  AND2_X1 U9389 ( .A1(n9977), .A2(n10082), .ZN(n6694) );
  XNOR2_X2 U9390 ( .A(n10395), .B(n10396), .ZN(n10397) );
  NOR2_X1 U9391 ( .A1(n15029), .A2(n15028), .ZN(n15027) );
  XNOR2_X1 U9392 ( .A(n12320), .B(n14413), .ZN(n14405) );
  NAND2_X1 U9393 ( .A1(n15012), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n15011) );
  XNOR2_X1 U9394 ( .A(n12945), .B(n12944), .ZN(n6922) );
  NAND2_X1 U9395 ( .A1(n7810), .A2(n7809), .ZN(n7228) );
  NAND2_X1 U9396 ( .A1(n9647), .A2(n6699), .ZN(n7600) );
  NAND2_X2 U9397 ( .A1(n8063), .A2(n12791), .ZN(n12794) );
  NAND2_X1 U9398 ( .A1(n10966), .A2(n7172), .ZN(n14491) );
  XNOR2_X1 U9399 ( .A(n6704), .B(n6703), .ZN(n12374) );
  AND2_X1 U9400 ( .A1(n12372), .A2(n12371), .ZN(n6705) );
  NOR2_X1 U9401 ( .A1(n7636), .A2(n7635), .ZN(n7637) );
  NAND2_X1 U9402 ( .A1(n7234), .A2(n8161), .ZN(n9055) );
  INV_X1 U9403 ( .A(n7085), .ZN(n7084) );
  NAND2_X2 U9404 ( .A1(n7726), .A2(n7725), .ZN(n7730) );
  NAND2_X1 U9405 ( .A1(n9148), .A2(n6711), .ZN(n9158) );
  NAND3_X1 U9406 ( .A1(n6713), .A2(n12988), .A3(n13006), .ZN(n6712) );
  NAND2_X1 U9407 ( .A1(n6714), .A2(n12846), .ZN(n8167) );
  NAND2_X1 U9408 ( .A1(n8166), .A2(n14494), .ZN(n6714) );
  XNOR2_X2 U9409 ( .A(n7483), .B(n8135), .ZN(n11202) );
  NAND2_X1 U9410 ( .A1(n7644), .A2(n7660), .ZN(n10262) );
  INV_X1 U9411 ( .A(n7408), .ZN(n7407) );
  NAND2_X1 U9412 ( .A1(n7201), .A2(n11796), .ZN(n12397) );
  NAND2_X1 U9413 ( .A1(n6984), .A2(n6503), .ZN(n6986) );
  NAND2_X1 U9414 ( .A1(n6986), .A2(n6985), .ZN(n8814) );
  OAI21_X2 U9415 ( .B1(n12488), .B2(n7207), .A(n7205), .ZN(n12466) );
  NOR2_X2 U9416 ( .A1(n12149), .A2(n10892), .ZN(n11697) );
  INV_X8 U9417 ( .A(n9617), .ZN(n11553) );
  NAND2_X1 U9418 ( .A1(n7263), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U9419 ( .A1(n13609), .A2(n6574), .ZN(n13606) );
  NAND2_X1 U9420 ( .A1(n13614), .A2(n13615), .ZN(n13609) );
  NAND2_X1 U9421 ( .A1(n6719), .A2(n6718), .ZN(n13662) );
  NAND2_X1 U9422 ( .A1(n13634), .A2(n13633), .ZN(n6719) );
  INV_X4 U9423 ( .A(n7364), .ZN(n11514) );
  XNOR2_X1 U9424 ( .A(n12340), .B(n15024), .ZN(n15012) );
  INV_X1 U9425 ( .A(n6724), .ZN(n8429) );
  NAND2_X1 U9426 ( .A1(n8483), .A2(n6732), .ZN(n6731) );
  NAND2_X1 U9427 ( .A1(n8239), .A2(n6736), .ZN(n6735) );
  NAND2_X1 U9428 ( .A1(n8328), .A2(n6738), .ZN(n6737) );
  NAND3_X1 U9429 ( .A1(n6755), .A2(n6819), .A3(n6753), .ZN(n6818) );
  NAND2_X1 U9430 ( .A1(n9679), .A2(n6758), .ZN(n9680) );
  NAND2_X1 U9431 ( .A1(n9626), .A2(n9627), .ZN(n6756) );
  NAND2_X1 U9432 ( .A1(n9625), .A2(n9624), .ZN(n6757) );
  NAND3_X1 U9433 ( .A1(n6762), .A2(n6586), .A3(n6761), .ZN(n6759) );
  NAND2_X1 U9434 ( .A1(n10321), .A2(n6764), .ZN(n6761) );
  NAND3_X1 U9435 ( .A1(n6762), .A2(n6763), .A3(n6761), .ZN(n10407) );
  INV_X1 U9436 ( .A(n10326), .ZN(n6764) );
  NAND2_X1 U9437 ( .A1(n10621), .A2(n10620), .ZN(n10623) );
  NAND2_X1 U9438 ( .A1(n10322), .A2(n10323), .ZN(n6767) );
  NAND2_X1 U9439 ( .A1(n13315), .A2(n13316), .ZN(n6777) );
  NAND2_X1 U9440 ( .A1(n6777), .A2(n6775), .ZN(n6772) );
  NAND2_X1 U9441 ( .A1(n7372), .A2(n6575), .ZN(n13340) );
  INV_X1 U9442 ( .A(n9544), .ZN(n9534) );
  INV_X2 U9443 ( .A(n7448), .ZN(n11967) );
  INV_X1 U9444 ( .A(n9533), .ZN(n6779) );
  INV_X1 U9445 ( .A(n9195), .ZN(n10037) );
  NAND2_X1 U9446 ( .A1(n9195), .A2(n7293), .ZN(n10460) );
  NAND2_X1 U9447 ( .A1(n9195), .A2(n7292), .ZN(n7295) );
  OR2_X1 U9448 ( .A1(n9195), .A2(n10377), .ZN(n10378) );
  NAND2_X1 U9449 ( .A1(n8891), .A2(n6785), .ZN(n6784) );
  OAI211_X1 U9450 ( .C1(n8891), .C2(n6786), .A(n6784), .B(n12004), .ZN(
        P3_U3154) );
  AND2_X4 U9451 ( .A1(n7015), .A2(n8815), .ZN(n8852) );
  NOR2_X1 U9452 ( .A1(n6716), .A2(n7198), .ZN(n8516) );
  NAND2_X1 U9453 ( .A1(n6716), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8503) );
  INV_X1 U9454 ( .A(n6800), .ZN(n6802) );
  NAND2_X1 U9455 ( .A1(n11806), .A2(n6801), .ZN(n6805) );
  NAND3_X1 U9456 ( .A1(n11790), .A2(n12447), .A3(n6804), .ZN(n6803) );
  INV_X1 U9457 ( .A(n12417), .ZN(n6809) );
  NAND2_X1 U9458 ( .A1(n6806), .A2(n6805), .ZN(n11811) );
  AOI21_X1 U9459 ( .B1(n6808), .B2(n6807), .A(n6812), .ZN(n6806) );
  INV_X1 U9460 ( .A(n11807), .ZN(n6812) );
  NAND3_X1 U9461 ( .A1(n6838), .A2(n11720), .A3(n6836), .ZN(n6835) );
  AND2_X2 U9462 ( .A1(n6852), .A2(n6570), .ZN(n14311) );
  NOR2_X1 U9463 ( .A1(n14596), .A2(n6853), .ZN(n14597) );
  NAND3_X1 U9464 ( .A1(n6858), .A2(n6856), .A3(n6855), .ZN(n6854) );
  NOR2_X1 U9465 ( .A1(n14262), .A2(n14263), .ZN(n14264) );
  NAND2_X1 U9466 ( .A1(n14262), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n6858) );
  AND2_X1 U9467 ( .A1(n14354), .A2(n14353), .ZN(n14615) );
  OAI21_X1 U9468 ( .B1(n14354), .B2(n6532), .A(n6864), .ZN(n14358) );
  NOR2_X2 U9469 ( .A1(n7562), .A2(n7456), .ZN(n7460) );
  NAND2_X1 U9470 ( .A1(n7544), .A2(n7453), .ZN(n7562) );
  OAI21_X1 U9471 ( .B1(n6868), .B2(n6866), .A(n10156), .ZN(n10241) );
  NAND2_X1 U9472 ( .A1(n6867), .A2(n9926), .ZN(n10154) );
  NAND2_X1 U9473 ( .A1(n10169), .A2(n9925), .ZN(n6867) );
  NAND2_X1 U9474 ( .A1(n11121), .A2(n6872), .ZN(n6870) );
  NAND2_X1 U9475 ( .A1(n6870), .A2(n6581), .ZN(n11275) );
  OAI21_X2 U9476 ( .B1(n8132), .B2(n6893), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n8173) );
  NOR2_X1 U9477 ( .A1(n7584), .A2(n9832), .ZN(n6896) );
  OR2_X2 U9478 ( .A1(n11090), .A2(n13484), .ZN(n7351) );
  NAND2_X1 U9479 ( .A1(n13916), .A2(n6899), .ZN(n6898) );
  NAND2_X1 U9480 ( .A1(n13916), .A2(n13917), .ZN(n13915) );
  INV_X1 U9481 ( .A(n14019), .ZN(n6911) );
  NAND2_X1 U9482 ( .A1(n14038), .A2(n14037), .ZN(n14036) );
  NAND2_X1 U9483 ( .A1(n11433), .A2(n6912), .ZN(n14080) );
  NAND2_X2 U9484 ( .A1(n7364), .A2(n11553), .ZN(n13464) );
  AOI21_X1 U9485 ( .B1(n7663), .B2(n6917), .A(n6916), .ZN(n6915) );
  INV_X1 U9486 ( .A(n7659), .ZN(n6917) );
  INV_X1 U9487 ( .A(n7663), .ZN(n6918) );
  NAND2_X1 U9488 ( .A1(n7664), .A2(n7663), .ZN(n7682) );
  NAND2_X1 U9489 ( .A1(n7660), .A2(n7659), .ZN(n7664) );
  NAND2_X1 U9490 ( .A1(n7643), .A2(n7642), .ZN(n7660) );
  NAND2_X1 U9491 ( .A1(n7228), .A2(n6928), .ZN(n6926) );
  NOR2_X1 U9492 ( .A1(n14546), .A2(n13607), .ZN(n6941) );
  NOR2_X2 U9493 ( .A1(n10551), .A2(n13556), .ZN(n10550) );
  NOR2_X2 U9494 ( .A1(n14115), .A2(n11617), .ZN(n13861) );
  NOR2_X2 U9495 ( .A1(n13959), .A2(n13943), .ZN(n6943) );
  OAI211_X2 U9496 ( .C1(n7584), .C2(n9618), .A(n7238), .B(n7237), .ZN(n11644)
         );
  NAND2_X1 U9497 ( .A1(n13055), .A2(n6950), .ZN(n12998) );
  INV_X1 U9498 ( .A(n6955), .ZN(n13011) );
  NAND2_X1 U9499 ( .A1(n6589), .A2(n10479), .ZN(n14505) );
  NAND2_X1 U9500 ( .A1(n12454), .A2(n12459), .ZN(n8650) );
  NAND2_X1 U9501 ( .A1(n12468), .A2(n8636), .ZN(n6958) );
  NAND2_X1 U9502 ( .A1(n11383), .A2(n6964), .ZN(n6962) );
  NAND2_X1 U9503 ( .A1(n6962), .A2(n6963), .ZN(n8548) );
  NAND2_X1 U9504 ( .A1(n12542), .A2(n6968), .ZN(n6967) );
  OAI21_X1 U9505 ( .B1(n10729), .B2(n6977), .A(n6976), .ZN(n6980) );
  XNOR2_X1 U9506 ( .A(n8714), .B(n6667), .ZN(n6981) );
  NAND2_X1 U9507 ( .A1(n12115), .A2(n6584), .ZN(n6995) );
  OAI211_X1 U9508 ( .C1(n12115), .C2(n6996), .A(n8921), .B(n6995), .ZN(
        P3_U3160) );
  OAI21_X2 U9509 ( .B1(n12076), .B2(n7007), .A(n6598), .ZN(n12049) );
  AOI21_X2 U9510 ( .B1(n12096), .B2(n12482), .A(n7009), .ZN(n12076) );
  NAND2_X1 U9511 ( .A1(n10744), .A2(n8832), .ZN(n10800) );
  NOR2_X2 U9512 ( .A1(n10057), .A2(n10058), .ZN(n10056) );
  INV_X1 U9513 ( .A(n14990), .ZN(n7023) );
  AOI21_X1 U9514 ( .B1(n14990), .B2(n7019), .A(n7020), .ZN(n7018) );
  INV_X1 U9515 ( .A(n14989), .ZN(n7022) );
  NAND3_X1 U9516 ( .A1(n7025), .A2(n7027), .A3(n7024), .ZN(n15009) );
  INV_X1 U9517 ( .A(n9978), .ZN(n10073) );
  NAND2_X1 U9518 ( .A1(n10094), .A2(n9982), .ZN(n10095) );
  AND2_X2 U9519 ( .A1(n7031), .A2(n6548), .ZN(n14424) );
  OR2_X2 U9520 ( .A1(n14405), .A2(n14406), .ZN(n7031) );
  AND2_X2 U9521 ( .A1(n10353), .A2(n10352), .ZN(n10395) );
  OR2_X2 U9522 ( .A1(n14442), .A2(n14443), .ZN(n12324) );
  NAND2_X1 U9523 ( .A1(n8296), .A2(n6507), .ZN(n7058) );
  NAND2_X1 U9524 ( .A1(n7058), .A2(n7056), .ZN(n8328) );
  NAND2_X1 U9525 ( .A1(n8296), .A2(n8294), .ZN(n7059) );
  OR2_X1 U9526 ( .A1(n8666), .A2(n7069), .ZN(n7067) );
  NAND2_X1 U9527 ( .A1(n8666), .A2(n7064), .ZN(n7061) );
  AOI21_X1 U9528 ( .B1(n8666), .B2(n8256), .A(n7068), .ZN(n8678) );
  NOR2_X1 U9529 ( .A1(n12318), .A2(n15008), .ZN(n15029) );
  NOR2_X2 U9530 ( .A1(n14424), .A2(n14423), .ZN(n14422) );
  NAND2_X1 U9531 ( .A1(n9930), .A2(n7093), .ZN(n7092) );
  NAND2_X1 U9532 ( .A1(n14826), .A2(n9933), .ZN(n7091) );
  NAND3_X1 U9533 ( .A1(n7092), .A2(n7091), .A3(n10170), .ZN(n9936) );
  NAND2_X1 U9534 ( .A1(n7095), .A2(n9933), .ZN(n10171) );
  NAND2_X1 U9535 ( .A1(n14811), .A2(n14810), .ZN(n7095) );
  INV_X1 U9536 ( .A(n9933), .ZN(n7096) );
  OAI21_X1 U9537 ( .B1(n13164), .B2(n7099), .A(n7097), .ZN(n13131) );
  OAI21_X1 U9538 ( .B1(n13110), .B2(n7105), .A(n6576), .ZN(n7109) );
  NAND2_X1 U9539 ( .A1(n10158), .A2(n7113), .ZN(n7110) );
  INV_X1 U9540 ( .A(n10158), .ZN(n7117) );
  NAND2_X1 U9541 ( .A1(n10579), .A2(n7120), .ZN(n7119) );
  NOR2_X1 U9542 ( .A1(n14615), .A2(n7122), .ZN(n7121) );
  NAND3_X1 U9543 ( .A1(n6495), .A2(n7128), .A3(n7124), .ZN(n14395) );
  NOR2_X1 U9544 ( .A1(n7127), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n7126) );
  NAND3_X1 U9545 ( .A1(n6495), .A2(n7128), .A3(n7126), .ZN(n7125) );
  NAND2_X1 U9546 ( .A1(n14360), .A2(n7129), .ZN(n7128) );
  INV_X1 U9547 ( .A(n14396), .ZN(n7129) );
  NAND2_X1 U9548 ( .A1(n7131), .A2(n14396), .ZN(n7130) );
  INV_X1 U9549 ( .A(n14393), .ZN(n7131) );
  NAND2_X1 U9550 ( .A1(n7143), .A2(n7145), .ZN(n7144) );
  NAND2_X1 U9551 ( .A1(n14604), .A2(n7147), .ZN(n7143) );
  INV_X1 U9552 ( .A(n14347), .ZN(n7149) );
  OAI21_X2 U9553 ( .B1(n7889), .B2(n7154), .A(n7150), .ZN(n12773) );
  OAI21_X2 U9554 ( .B1(n12794), .B2(n7166), .A(n7163), .ZN(n8122) );
  NAND2_X1 U9555 ( .A1(n12784), .A2(n7169), .ZN(n8000) );
  INV_X1 U9556 ( .A(n12787), .ZN(n7171) );
  INV_X1 U9557 ( .A(n10965), .ZN(n7173) );
  NAND2_X1 U9558 ( .A1(n10790), .A2(n7748), .ZN(n7765) );
  NAND3_X1 U9559 ( .A1(n7460), .A2(n7771), .A3(n6474), .ZN(n7485) );
  NOR2_X2 U9560 ( .A1(n7485), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7484) );
  NAND2_X1 U9561 ( .A1(n7175), .A2(n7176), .ZN(n8740) );
  NAND2_X1 U9562 ( .A1(n8738), .A2(n7178), .ZN(n7175) );
  AND2_X1 U9563 ( .A1(n12559), .A2(n7177), .ZN(n7176) );
  NAND2_X1 U9564 ( .A1(n7181), .A2(n7182), .ZN(n8735) );
  NAND2_X1 U9565 ( .A1(n8733), .A2(n7183), .ZN(n7181) );
  OAI21_X2 U9566 ( .B1(n11388), .B2(n7190), .A(n7187), .ZN(n12584) );
  INV_X1 U9567 ( .A(n12584), .ZN(n8737) );
  OAI21_X1 U9568 ( .B1(n12416), .B2(n11799), .A(n7202), .ZN(n12399) );
  AND2_X1 U9569 ( .A1(n8756), .A2(n7013), .ZN(n8757) );
  AND2_X2 U9570 ( .A1(n8756), .A2(n6579), .ZN(n8216) );
  OR2_X1 U9571 ( .A1(n13437), .A2(n13436), .ZN(n13439) );
  OAI21_X1 U9572 ( .B1(n7730), .B2(n7220), .A(n7219), .ZN(n7788) );
  NAND2_X1 U9573 ( .A1(n7218), .A2(n7216), .ZN(n7791) );
  NAND2_X1 U9574 ( .A1(n7730), .A2(n7219), .ZN(n7218) );
  NAND2_X1 U9575 ( .A1(n11554), .A2(n8003), .ZN(n7224) );
  NAND2_X1 U9576 ( .A1(n7224), .A2(n7223), .ZN(n8025) );
  INV_X1 U9577 ( .A(n6461), .ZN(n7540) );
  NAND2_X1 U9578 ( .A1(n7478), .A2(n7479), .ZN(n7538) );
  OAI21_X2 U9579 ( .B1(n8065), .B2(n8064), .A(n8066), .ZN(n8086) );
  NAND2_X1 U9580 ( .A1(n8159), .A2(n7232), .ZN(n7230) );
  NAND2_X1 U9581 ( .A1(n7522), .A2(n14742), .ZN(n7237) );
  NAND2_X2 U9582 ( .A1(n7472), .A2(n7471), .ZN(n7524) );
  NAND2_X1 U9583 ( .A1(n11354), .A2(n7241), .ZN(n7239) );
  NAND2_X1 U9584 ( .A1(n7464), .A2(n7252), .ZN(n8132) );
  NAND2_X1 U9585 ( .A1(n13029), .A2(n7255), .ZN(n7254) );
  NAND2_X1 U9586 ( .A1(n13709), .A2(n13708), .ZN(n7262) );
  NAND2_X1 U9587 ( .A1(n13705), .A2(n13704), .ZN(n7263) );
  NAND2_X1 U9588 ( .A1(n13693), .A2(n7266), .ZN(n7265) );
  INV_X1 U9589 ( .A(n13700), .ZN(n7271) );
  NAND2_X1 U9590 ( .A1(n13662), .A2(n6585), .ZN(n7274) );
  NAND2_X1 U9591 ( .A1(n7274), .A2(n6578), .ZN(n13666) );
  NAND2_X1 U9592 ( .A1(n7277), .A2(n7278), .ZN(n13614) );
  NAND3_X1 U9593 ( .A1(n13600), .A2(n13599), .A3(n6587), .ZN(n7277) );
  NAND3_X1 U9594 ( .A1(n13674), .A2(n13673), .A3(n7283), .ZN(n7281) );
  NAND2_X1 U9595 ( .A1(n13579), .A2(n13580), .ZN(n13578) );
  NAND3_X1 U9596 ( .A1(n13553), .A2(n13552), .A3(n6580), .ZN(n7289) );
  NAND2_X1 U9597 ( .A1(n7289), .A2(n7290), .ZN(n13560) );
  NAND3_X1 U9598 ( .A1(n7300), .A2(n7299), .A3(n8946), .ZN(n7297) );
  NAND2_X1 U9599 ( .A1(n9028), .A2(n7304), .ZN(n7301) );
  NAND2_X1 U9600 ( .A1(n7301), .A2(n7302), .ZN(n9035) );
  INV_X1 U9601 ( .A(n9032), .ZN(n7313) );
  NOR2_X1 U9602 ( .A1(n7484), .A2(n13281), .ZN(n7315) );
  OAI21_X1 U9603 ( .B1(n9015), .B2(n7320), .A(n7317), .ZN(n7325) );
  INV_X1 U9604 ( .A(n8967), .ZN(n7339) );
  INV_X1 U9605 ( .A(n8968), .ZN(n7340) );
  NAND2_X1 U9606 ( .A1(n7343), .A2(n7344), .ZN(n8958) );
  OAI21_X1 U9607 ( .B1(n9853), .B2(n9854), .A(n7346), .ZN(n9855) );
  NAND2_X1 U9608 ( .A1(n7346), .A2(n10220), .ZN(n10221) );
  CLKBUF_X1 U9609 ( .A(n7364), .Z(n7361) );
  NAND2_X2 U9610 ( .A1(n7364), .A2(n9617), .ZN(n13436) );
  NAND2_X1 U9611 ( .A1(n11514), .A2(n7362), .ZN(n9619) );
  MUX2_X1 U9612 ( .A(n14255), .B(n14621), .S(n11514), .Z(n9744) );
  NAND2_X1 U9613 ( .A1(n11859), .A2(n7373), .ZN(n7372) );
  NAND2_X1 U9614 ( .A1(n13367), .A2(n7380), .ZN(n7379) );
  OAI21_X1 U9615 ( .B1(n13349), .B2(n13350), .A(n11958), .ZN(n13415) );
  NAND2_X1 U9616 ( .A1(n7405), .A2(n9285), .ZN(n9495) );
  NAND2_X1 U9617 ( .A1(n7410), .A2(n7409), .ZN(n9851) );
  NAND3_X1 U9618 ( .A1(n9741), .A2(n9740), .A3(n13539), .ZN(n7410) );
  NAND2_X1 U9619 ( .A1(n10928), .A2(n7415), .ZN(n7413) );
  AND2_X1 U9620 ( .A1(n7425), .A2(n7426), .ZN(n13898) );
  AND2_X1 U9621 ( .A1(n9194), .A2(n6566), .ZN(n7435) );
  NAND2_X1 U9622 ( .A1(n11647), .A2(n11810), .ZN(n11673) );
  INV_X1 U9623 ( .A(n10684), .ZN(n8319) );
  NAND2_X1 U9624 ( .A1(n8303), .A2(n8302), .ZN(n10684) );
  INV_X1 U9625 ( .A(n14119), .ZN(n14120) );
  NAND2_X1 U9626 ( .A1(n8650), .A2(n8649), .ZN(n12440) );
  OAI211_X1 U9627 ( .C1(n8191), .C2(n13190), .A(n8190), .B(n8189), .ZN(
        P2_U3192) );
  NAND2_X1 U9628 ( .A1(n8167), .A2(n13190), .ZN(n8190) );
  NAND2_X1 U9629 ( .A1(n9508), .A2(n14254), .ZN(n13457) );
  AND2_X1 U9630 ( .A1(n13440), .A2(n13442), .ZN(n13505) );
  NOR2_X1 U9631 ( .A1(n9379), .A2(n7546), .ZN(n7547) );
  INV_X1 U9632 ( .A(n14075), .ZN(n14163) );
  OAI21_X1 U9633 ( .B1(n14118), .B2(n14716), .A(n14117), .ZN(n14119) );
  NAND2_X1 U9634 ( .A1(n11173), .A2(n8387), .ZN(n11209) );
  AOI22_X1 U9635 ( .A1(n9710), .A2(n11967), .B1(n9737), .B2(n11966), .ZN(n9622) );
  INV_X1 U9636 ( .A(n11637), .ZN(n9918) );
  INV_X1 U9637 ( .A(n8172), .ZN(n8109) );
  INV_X1 U9638 ( .A(n6485), .ZN(n9128) );
  NAND2_X1 U9639 ( .A1(n8768), .A2(n8767), .ZN(n12749) );
  INV_X1 U9640 ( .A(n9379), .ZN(n7522) );
  AOI211_X1 U9641 ( .C1(n13001), .C2(n9158), .A(n9154), .B(n9153), .ZN(n9155)
         );
  NAND2_X1 U9642 ( .A1(n8025), .A2(n8024), .ZN(n8044) );
  NOR2_X1 U9643 ( .A1(n11553), .A2(P3_STATE_REG_SCAN_IN), .ZN(n14376) );
  NAND2_X1 U9644 ( .A1(n7963), .A2(n7962), .ZN(n7967) );
  AOI22_X1 U9645 ( .A1(n9932), .A2(n9091), .B1(n12868), .B2(n6433), .ZN(n8947)
         );
  AND2_X1 U9646 ( .A1(n7515), .A2(n13286), .ZN(n7551) );
  INV_X1 U9647 ( .A(n7515), .ZN(n11470) );
  XNOR2_X1 U9648 ( .A(n12363), .B(n11674), .ZN(n7437) );
  AND2_X1 U9649 ( .A1(n12381), .A2(n14482), .ZN(n7438) );
  AND2_X1 U9650 ( .A1(n7499), .A2(n7498), .ZN(n7440) );
  OR2_X1 U9651 ( .A1(n14142), .A2(n13732), .ZN(n7441) );
  AND2_X1 U9652 ( .A1(n11915), .A2(n11914), .ZN(n7442) );
  OR2_X1 U9653 ( .A1(n11953), .A2(n13731), .ZN(n7443) );
  NOR2_X1 U9654 ( .A1(n7943), .A2(n9218), .ZN(n7444) );
  AND2_X1 U9655 ( .A1(n8703), .A2(n12132), .ZN(n7445) );
  INV_X1 U9656 ( .A(n13301), .ZN(n13289) );
  AND2_X1 U9657 ( .A1(n8117), .A2(n8116), .ZN(n12943) );
  INV_X1 U9658 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n10755) );
  NOR2_X1 U9659 ( .A1(n7776), .A2(n7756), .ZN(n7446) );
  INV_X1 U9660 ( .A(n12988), .ZN(n12944) );
  INV_X1 U9661 ( .A(n11295), .ZN(n9167) );
  INV_X1 U9662 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n10725) );
  INV_X1 U9663 ( .A(n12843), .ZN(n12947) );
  NAND2_X1 U9664 ( .A1(n9397), .A2(n9378), .ZN(n12843) );
  OR2_X1 U9665 ( .A1(n14331), .A2(n14330), .ZN(n7447) );
  INV_X1 U9666 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7818) );
  NAND2_X1 U9667 ( .A1(n9915), .A2(n14819), .ZN(n14515) );
  AND2_X1 U9668 ( .A1(n9114), .A2(n9105), .ZN(n7449) );
  AND2_X1 U9669 ( .A1(n13887), .A2(n14044), .ZN(n14650) );
  INV_X1 U9670 ( .A(n14650), .ZN(n14047) );
  INV_X1 U9671 ( .A(n14254), .ZN(n9526) );
  INV_X1 U9672 ( .A(n13861), .ZN(n13899) );
  INV_X2 U9673 ( .A(n14462), .ZN(n15120) );
  AND2_X2 U9674 ( .A1(n10186), .A2(n8794), .ZN(n15149) );
  NAND2_X1 U9675 ( .A1(n8857), .A2(n12581), .ZN(n7450) );
  NOR2_X1 U9676 ( .A1(n8741), .A2(n12531), .ZN(n7451) );
  OR3_X1 U9677 ( .A1(n12075), .A2(n12441), .A3(n12137), .ZN(n7452) );
  INV_X1 U9678 ( .A(n12421), .ZN(n12442) );
  AND4_X1 U9679 ( .A1(n8675), .A2(n8674), .A3(n8673), .A4(n8672), .ZN(n12421)
         );
  NAND2_X1 U9680 ( .A1(n6433), .A2(n12870), .ZN(n8923) );
  NAND2_X1 U9681 ( .A1(n12869), .A2(n9091), .ZN(n8938) );
  OAI22_X1 U9682 ( .A1(n14895), .A2(n9092), .B1(n10155), .B2(n9043), .ZN(n8954) );
  INV_X1 U9683 ( .A(n8955), .ZN(n8956) );
  INV_X1 U9684 ( .A(n8961), .ZN(n8962) );
  INV_X1 U9685 ( .A(n11686), .ZN(n11677) );
  INV_X1 U9686 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n8201) );
  AOI21_X1 U9687 ( .B1(n9042), .B2(n9041), .A(n9040), .ZN(n9049) );
  NAND2_X1 U9688 ( .A1(n9116), .A2(n9117), .ZN(n9118) );
  INV_X1 U9689 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n8203) );
  AND2_X1 U9690 ( .A1(n9119), .A2(n9118), .ZN(n9120) );
  INV_X1 U9691 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n7881) );
  INV_X1 U9692 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n7465) );
  INV_X1 U9693 ( .A(n11856), .ZN(n11857) );
  NAND2_X1 U9694 ( .A1(n11839), .A2(n11670), .ZN(n11671) );
  AND2_X1 U9695 ( .A1(n8536), .A2(n8519), .ZN(n8558) );
  INV_X1 U9696 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n8419) );
  INV_X1 U9697 ( .A(n11815), .ZN(n8318) );
  INV_X1 U9698 ( .A(n7905), .ZN(n7903) );
  NAND2_X1 U9699 ( .A1(n8007), .A2(n8006), .ZN(n8030) );
  OR2_X1 U9700 ( .A1(n7927), .A2(n7926), .ZN(n7948) );
  OR2_X1 U9701 ( .A1(n7713), .A2(n7712), .ZN(n7737) );
  OR2_X1 U9702 ( .A1(n9379), .A2(n9388), .ZN(n7565) );
  INV_X1 U9703 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n7468) );
  NAND2_X1 U9704 ( .A1(n11855), .A2(n11857), .ZN(n11858) );
  INV_X1 U9705 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n10223) );
  INV_X1 U9706 ( .A(n13487), .ZN(n11236) );
  INV_X1 U9707 ( .A(n13961), .ZN(n11616) );
  INV_X1 U9708 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n9184) );
  NOR2_X1 U9709 ( .A1(n14260), .A2(n14261), .ZN(n14263) );
  INV_X1 U9710 ( .A(n10745), .ZN(n8831) );
  INV_X1 U9711 ( .A(n8798), .ZN(n8799) );
  INV_X1 U9712 ( .A(SI_18_), .ZN(n12267) );
  OR2_X1 U9713 ( .A1(n11655), .A2(n8274), .ZN(n8276) );
  INV_X1 U9714 ( .A(n14982), .ZN(n12333) );
  OR2_X1 U9715 ( .A1(n8681), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U9716 ( .A1(n8690), .A2(n8689), .ZN(n12402) );
  AND2_X1 U9717 ( .A1(n11746), .A2(n11745), .ZN(n11743) );
  OR2_X1 U9718 ( .A1(n8422), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8440) );
  OAI21_X1 U9719 ( .B1(n8782), .B2(n8781), .A(n8780), .ZN(n8802) );
  AND2_X1 U9720 ( .A1(n8197), .A2(n8196), .ZN(n8198) );
  NOR2_X1 U9721 ( .A1(n7737), .A2(n7736), .ZN(n7755) );
  OR2_X1 U9722 ( .A1(n8052), .A2(n12797), .ZN(n8071) );
  NAND2_X1 U9723 ( .A1(n7946), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n7971) );
  AND2_X1 U9724 ( .A1(n7755), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7776) );
  OR2_X1 U9725 ( .A1(n8071), .A2(n8070), .ZN(n8106) );
  OR2_X1 U9726 ( .A1(n7971), .A2(n7970), .ZN(n8009) );
  INV_X1 U9727 ( .A(n13190), .ZN(n12909) );
  NAND2_X1 U9728 ( .A1(n7860), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n7882) );
  AND2_X1 U9729 ( .A1(n9129), .A2(n6464), .ZN(n9378) );
  NAND2_X1 U9730 ( .A1(n7522), .A2(n7521), .ZN(n7526) );
  INV_X1 U9731 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10937) );
  INV_X1 U9732 ( .A(n10810), .ZN(n10811) );
  AND2_X1 U9733 ( .A1(n14566), .A2(n14567), .ZN(n11870) );
  INV_X1 U9734 ( .A(n11493), .ZN(n11485) );
  INV_X1 U9735 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n11228) );
  INV_X1 U9736 ( .A(n14111), .ZN(n13860) );
  INV_X1 U9737 ( .A(n11484), .ZN(n11477) );
  INV_X1 U9738 ( .A(n11558), .ZN(n11571) );
  INV_X1 U9739 ( .A(n11096), .ZN(n11097) );
  NAND2_X1 U9740 ( .A1(n13958), .A2(n11616), .ZN(n13959) );
  OR2_X1 U9741 ( .A1(n8910), .A2(n8907), .ZN(n12109) );
  OR2_X1 U9742 ( .A1(n8804), .A2(n8803), .ZN(n8910) );
  INV_X1 U9743 ( .A(n10388), .ZN(n10396) );
  INV_X1 U9744 ( .A(n10763), .ZN(n10770) );
  NOR2_X1 U9745 ( .A1(n8694), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8696) );
  AND2_X1 U9746 ( .A1(n11786), .A2(n11785), .ZN(n12447) );
  OR2_X1 U9747 ( .A1(n8310), .A2(n10366), .ZN(n8598) );
  AND2_X1 U9748 ( .A1(n12535), .A2(n12534), .ZN(n12660) );
  NAND2_X1 U9749 ( .A1(n8550), .A2(n8549), .ZN(n12542) );
  INV_X1 U9750 ( .A(n11743), .ZN(n12583) );
  INV_X1 U9751 ( .A(n11732), .ZN(n11320) );
  INV_X1 U9752 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8339) );
  OR2_X1 U9753 ( .A1(n9282), .A2(n10183), .ZN(n8798) );
  AND2_X1 U9754 ( .A1(n11736), .A2(n11735), .ZN(n11827) );
  AND2_X1 U9755 ( .A1(n8801), .A2(n11675), .ZN(n15093) );
  INV_X1 U9756 ( .A(n9330), .ZN(n8780) );
  XNOR2_X1 U9757 ( .A(n8122), .B(n8121), .ZN(n8166) );
  INV_X1 U9758 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U9759 ( .A1(n8180), .A2(n8179), .ZN(n12783) );
  NOR2_X1 U9760 ( .A1(n8183), .A2(n14851), .ZN(n8180) );
  OR2_X1 U9761 ( .A1(n8182), .A2(n8109), .ZN(n8117) );
  INV_X1 U9762 ( .A(n12874), .ZN(n12882) );
  INV_X1 U9763 ( .A(n10578), .ZN(n10585) );
  INV_X1 U9764 ( .A(n14816), .ZN(n13169) );
  OR3_X1 U9765 ( .A1(n13139), .A2(n13138), .A3(n13169), .ZN(n13242) );
  INV_X1 U9766 ( .A(n14814), .ZN(n14834) );
  NAND2_X1 U9767 ( .A1(n10707), .A2(n10709), .ZN(n10710) );
  OR2_X1 U9768 ( .A1(n10938), .A2(n10937), .ZN(n11077) );
  INV_X1 U9769 ( .A(n13983), .ZN(n13352) );
  INV_X1 U9770 ( .A(n13418), .ZN(n14565) );
  INV_X1 U9771 ( .A(n13928), .ZN(n13417) );
  INV_X1 U9772 ( .A(n6465), .ZN(n11545) );
  INV_X1 U9773 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n14259) );
  INV_X1 U9774 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n11044) );
  INV_X1 U9775 ( .A(n6468), .ZN(n9525) );
  INV_X1 U9776 ( .A(n13958), .ZN(n13974) );
  OR2_X1 U9777 ( .A1(n14075), .A2(n13920), .ZN(n9785) );
  INV_X1 U9778 ( .A(n9712), .ZN(n13469) );
  NAND2_X1 U9779 ( .A1(n9507), .A2(n11853), .ZN(n13957) );
  INV_X1 U9780 ( .A(n13740), .ZN(n14564) );
  INV_X1 U9781 ( .A(n13480), .ZN(n10846) );
  INV_X1 U9782 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n14233) );
  NOR2_X1 U9783 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n14308), .ZN(n14268) );
  OAI22_X1 U9784 ( .A1(n14312), .A2(n14271), .B1(P1_ADDR_REG_6__SCAN_IN), .B2(
        n14270), .ZN(n14272) );
  INV_X1 U9785 ( .A(n12049), .ZN(n12050) );
  INV_X1 U9786 ( .A(n12109), .ZN(n12128) );
  INV_X1 U9787 ( .A(n12126), .ZN(n12107) );
  OR2_X1 U9788 ( .A1(n6430), .A2(n8709), .ZN(n11659) );
  AND4_X1 U9789 ( .A1(n8635), .A2(n8634), .A3(n8633), .A4(n8632), .ZN(n12482)
         );
  INV_X1 U9790 ( .A(n12367), .ZN(n15048) );
  INV_X1 U9791 ( .A(n12363), .ZN(n12375) );
  AND2_X1 U9792 ( .A1(n8696), .A2(n8911), .ZN(n14459) );
  AND3_X1 U9793 ( .A1(n9989), .A2(n6425), .A3(n11804), .ZN(n12569) );
  AND2_X1 U9794 ( .A1(n8719), .A2(n11804), .ZN(n12571) );
  INV_X1 U9795 ( .A(n15093), .ZN(n15109) );
  NAND2_X1 U9796 ( .A1(n15116), .A2(n10897), .ZN(n12589) );
  INV_X1 U9797 ( .A(n11406), .ZN(n11319) );
  AND3_X1 U9798 ( .A1(n8798), .A2(n8804), .A3(n8788), .ZN(n10186) );
  INV_X1 U9799 ( .A(n15138), .ZN(n14476) );
  OR2_X1 U9800 ( .A1(n15090), .A2(n6605), .ZN(n14482) );
  AND2_X1 U9801 ( .A1(n9968), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9329) );
  NOR2_X1 U9802 ( .A1(n8181), .A2(n12783), .ZN(n8188) );
  INV_X1 U9803 ( .A(n14895), .ZN(n9942) );
  INV_X1 U9804 ( .A(n14502), .ZN(n12842) );
  NAND2_X1 U9805 ( .A1(n8165), .A2(n14819), .ZN(n14499) );
  INV_X1 U9806 ( .A(n8110), .ZN(n9078) );
  AND2_X1 U9807 ( .A1(n7933), .A2(n7932), .ZN(n12964) );
  INV_X1 U9808 ( .A(n14765), .ZN(n14795) );
  AND2_X1 U9809 ( .A1(n9384), .A2(n13295), .ZN(n14765) );
  OAI21_X1 U9810 ( .B1(n12943), .B2(n12843), .A(n12950), .ZN(n12951) );
  INV_X1 U9811 ( .A(n14820), .ZN(n14507) );
  AND2_X1 U9812 ( .A1(n6660), .A2(n14945), .ZN(n13261) );
  INV_X1 U9813 ( .A(n13261), .ZN(n14913) );
  NOR2_X1 U9814 ( .A1(n11148), .A2(n11147), .ZN(n11158) );
  INV_X1 U9815 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n13281) );
  AND2_X1 U9816 ( .A1(n9543), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9235) );
  OR2_X1 U9817 ( .A1(n11077), .A2(n11076), .ZN(n11229) );
  NOR2_X1 U9818 ( .A1(n9548), .A2(n9780), .ZN(n13332) );
  INV_X1 U9819 ( .A(n13503), .ZN(n13866) );
  AND2_X1 U9820 ( .A1(n11536), .A2(n11535), .ZN(n13522) );
  INV_X1 U9821 ( .A(n13873), .ZN(n13897) );
  INV_X1 U9822 ( .A(n14020), .ZN(n14085) );
  OR2_X1 U9823 ( .A1(n9785), .A2(n13715), .ZN(n14044) );
  AND2_X1 U9824 ( .A1(n10123), .A2(n13920), .ZN(n14659) );
  AOI21_X1 U9825 ( .B1(n9505), .B2(n9504), .A(n9503), .ZN(n9782) );
  INV_X1 U9826 ( .A(n14192), .ZN(n14725) );
  NOR2_X1 U9827 ( .A1(n9780), .A2(n9502), .ZN(n9573) );
  OAI211_X1 U9828 ( .C1(n11448), .C2(n9237), .A(n14244), .B(n9236), .ZN(n9499)
         );
  AND2_X1 U9829 ( .A1(n10038), .A2(n10037), .ZN(n13818) );
  AND2_X1 U9830 ( .A1(n9327), .A2(n9354), .ZN(n10493) );
  AND2_X1 U9831 ( .A1(n10012), .A2(n10011), .ZN(n14998) );
  NOR2_X1 U9832 ( .A1(n8920), .A2(n7445), .ZN(n8921) );
  INV_X1 U9833 ( .A(n12505), .ZN(n12651) );
  INV_X1 U9834 ( .A(n12117), .ZN(n12130) );
  INV_X1 U9835 ( .A(n12433), .ZN(n12404) );
  INV_X1 U9836 ( .A(n12470), .ZN(n12499) );
  INV_X1 U9837 ( .A(n12597), .ZN(n12570) );
  NAND2_X1 U9838 ( .A1(P3_U3897), .A2(n8211), .ZN(n15042) );
  INV_X1 U9839 ( .A(n12589), .ZN(n12618) );
  NAND2_X1 U9840 ( .A1(n8918), .A2(n8917), .ZN(n15114) );
  NAND2_X1 U9841 ( .A1(n11319), .A2(n14476), .ZN(n12587) );
  INV_X1 U9842 ( .A(n15149), .ZN(n15150) );
  INV_X2 U9843 ( .A(n15144), .ZN(n15143) );
  NAND2_X1 U9844 ( .A1(n9330), .A2(n9329), .ZN(n9334) );
  INV_X1 U9845 ( .A(n9329), .ZN(n9325) );
  INV_X1 U9846 ( .A(n8800), .ZN(n10368) );
  INV_X1 U9847 ( .A(SI_16_), .ZN(n12244) );
  INV_X1 U9848 ( .A(n14375), .ZN(n12726) );
  NOR2_X1 U9849 ( .A1(n8188), .A2(n8187), .ZN(n8189) );
  INV_X1 U9850 ( .A(n12943), .ZN(n12946) );
  INV_X1 U9851 ( .A(n12964), .ZN(n12930) );
  INV_X1 U9852 ( .A(n11364), .ZN(n12856) );
  INV_X1 U9853 ( .A(n10582), .ZN(n12862) );
  CLKBUF_X2 U9854 ( .A(P2_U3947), .Z(n12871) );
  INV_X1 U9855 ( .A(n14805), .ZN(n12878) );
  OR2_X1 U9856 ( .A1(n9393), .A2(n13295), .ZN(n14786) );
  OR2_X1 U9857 ( .A1(n9915), .A2(n12903), .ZN(n14820) );
  AND2_X1 U9858 ( .A1(n14840), .A2(n9917), .ZN(n13178) );
  INV_X1 U9859 ( .A(n14970), .ZN(n14968) );
  OR2_X1 U9860 ( .A1(n13246), .A2(n13245), .ZN(n13277) );
  INV_X1 U9861 ( .A(n14952), .ZN(n14950) );
  INV_X1 U9862 ( .A(n14848), .ZN(n14846) );
  INV_X1 U9863 ( .A(n14854), .ZN(n14851) );
  INV_X1 U9864 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n13297) );
  INV_X1 U9865 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n12205) );
  NAND2_X1 U9866 ( .A1(n9891), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14580) );
  INV_X1 U9867 ( .A(n14576), .ZN(n13434) );
  INV_X1 U9868 ( .A(n13522), .ZN(n13734) );
  INV_X1 U9869 ( .A(n13628), .ZN(n14084) );
  INV_X1 U9870 ( .A(n14637), .ZN(n13807) );
  INV_X1 U9871 ( .A(n14627), .ZN(n14645) );
  INV_X1 U9872 ( .A(n14047), .ZN(n14673) );
  INV_X1 U9873 ( .A(n14734), .ZN(n14732) );
  INV_X1 U9874 ( .A(n13612), .ZN(n13435) );
  INV_X1 U9875 ( .A(n14729), .ZN(n14727) );
  AND2_X2 U9876 ( .A1(n9573), .A2(n9572), .ZN(n14729) );
  INV_X1 U9877 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n9643) );
  NOR2_X1 U9878 ( .A1(P2_U3088), .A2(n9382), .ZN(P2_U3947) );
  NOR2_X2 U9879 ( .A1(n9544), .A2(n9202), .ZN(P1_U4016) );
  INV_X2 U9880 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n7616) );
  NAND4_X1 U9881 ( .A1(n7563), .A2(n7455), .A3(n7616), .A4(n7454), .ZN(n7456)
         );
  NOR2_X1 U9882 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n7459) );
  INV_X1 U9883 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n7666) );
  AND4_X2 U9884 ( .A1(n7459), .A2(n7458), .A3(n7457), .A4(n7666), .ZN(n7771)
         );
  NOR2_X1 U9885 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n7467) );
  NOR2_X1 U9886 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n7466) );
  INV_X1 U9887 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n7469) );
  NAND2_X1 U9888 ( .A1(n8174), .A2(n7469), .ZN(n7470) );
  NAND2_X1 U9889 ( .A1(n9170), .A2(n7470), .ZN(n7471) );
  NAND2_X1 U9890 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n14739), .ZN(n7473) );
  INV_X2 U9891 ( .A(n9212), .ZN(n9617) );
  NAND2_X1 U9892 ( .A1(n7476), .A2(SI_1_), .ZN(n7537) );
  OAI21_X1 U9893 ( .B1(n7476), .B2(SI_1_), .A(n7537), .ZN(n7481) );
  INV_X1 U9894 ( .A(n7481), .ZN(n7478) );
  INV_X1 U9895 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8280) );
  INV_X1 U9896 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n8229) );
  INV_X1 U9897 ( .A(SI_0_), .ZN(n9515) );
  NOR2_X1 U9898 ( .A1(n7477), .A2(n9515), .ZN(n7479) );
  INV_X1 U9899 ( .A(n7479), .ZN(n7480) );
  NAND2_X1 U9900 ( .A1(n7481), .A2(n7480), .ZN(n7482) );
  NAND2_X1 U9901 ( .A1(n7538), .A2(n7482), .ZN(n9618) );
  INV_X1 U9902 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U9903 ( .A1(n7486), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7487) );
  NAND2_X1 U9904 ( .A1(n7487), .A2(P2_IR_REG_20__SCAN_IN), .ZN(n7490) );
  INV_X1 U9905 ( .A(n7484), .ZN(n7491) );
  NAND2_X1 U9906 ( .A1(n7464), .A2(n7493), .ZN(n7832) );
  NAND2_X1 U9907 ( .A1(n7853), .A2(n7494), .ZN(n7855) );
  AND2_X1 U9908 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n7495) );
  INV_X1 U9909 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n7497) );
  INV_X1 U9910 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n7496) );
  NAND3_X1 U9911 ( .A1(n7497), .A2(n7496), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n7499) );
  XNOR2_X1 U9912 ( .A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_19__SCAN_IN), .ZN(
        n7498) );
  INV_X2 U9913 ( .A(n12903), .ZN(n13001) );
  NAND2_X1 U9914 ( .A1(n6462), .A2(n13001), .ZN(n7842) );
  NOR2_X1 U9915 ( .A1(P2_IR_REG_27__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n7506) );
  NOR2_X1 U9916 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n7505) );
  NAND4_X1 U9917 ( .A1(n6474), .A2(n7507), .A3(n7506), .A4(n7505), .ZN(n7508)
         );
  NAND2_X1 U9918 ( .A1(n7511), .A2(n7509), .ZN(n13282) );
  INV_X1 U9919 ( .A(n7511), .ZN(n7512) );
  NAND2_X1 U9920 ( .A1(n7512), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7513) );
  AND2_X4 U9921 ( .A1(n7515), .A2(n7516), .ZN(n8172) );
  NAND2_X1 U9922 ( .A1(n8172), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n7520) );
  NAND2_X1 U9923 ( .A1(n7552), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n7519) );
  NAND2_X1 U9924 ( .A1(n7551), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n7518) );
  AND2_X2 U9925 ( .A1(n11470), .A2(n7516), .ZN(n7550) );
  NAND2_X1 U9926 ( .A1(n7550), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n7517) );
  NAND2_X1 U9927 ( .A1(n7842), .A2(n12870), .ZN(n7534) );
  XNOR2_X1 U9928 ( .A(n7533), .B(n7534), .ZN(n11629) );
  INV_X1 U9929 ( .A(n14739), .ZN(n7521) );
  NAND2_X1 U9930 ( .A1(n11553), .A2(SI_0_), .ZN(n7523) );
  XNOR2_X1 U9931 ( .A(n7523), .B(n8229), .ZN(n13304) );
  NAND2_X1 U9932 ( .A1(n9379), .A2(n13304), .ZN(n7525) );
  NAND2_X2 U9933 ( .A1(n7526), .A2(n7525), .ZN(n14831) );
  AND2_X1 U9934 ( .A1(n8119), .A2(n14831), .ZN(n7532) );
  NAND2_X1 U9935 ( .A1(n7552), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n7529) );
  NAND2_X1 U9936 ( .A1(n7550), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7528) );
  NAND2_X1 U9937 ( .A1(n7551), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n7527) );
  NAND2_X1 U9938 ( .A1(n8172), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7530) );
  NAND2_X1 U9939 ( .A1(n7531), .A2(n7530), .ZN(n12872) );
  INV_X1 U9940 ( .A(n12872), .ZN(n11624) );
  OAI21_X1 U9941 ( .B1(n14831), .B2(n7842), .A(n9927), .ZN(n11472) );
  NAND2_X1 U9942 ( .A1(n11629), .A2(n11628), .ZN(n11627) );
  INV_X1 U9943 ( .A(n7533), .ZN(n7535) );
  NAND2_X1 U9944 ( .A1(n7535), .A2(n7534), .ZN(n7536) );
  NAND2_X1 U9945 ( .A1(n11627), .A2(n7536), .ZN(n9579) );
  MUX2_X1 U9946 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9212), .Z(n7539) );
  NAND2_X1 U9947 ( .A1(n7539), .A2(SI_2_), .ZN(n7567) );
  OAI21_X1 U9948 ( .B1(n7539), .B2(SI_2_), .A(n7567), .ZN(n7541) );
  NAND2_X1 U9949 ( .A1(n7540), .A2(n7541), .ZN(n7543) );
  INV_X1 U9950 ( .A(n7541), .ZN(n7542) );
  NAND2_X1 U9951 ( .A1(n7543), .A2(n7568), .ZN(n9674) );
  OR2_X1 U9952 ( .A1(n7544), .A2(n13281), .ZN(n7545) );
  XNOR2_X1 U9953 ( .A(n7545), .B(P2_IR_REG_2__SCAN_IN), .ZN(n14755) );
  INV_X1 U9954 ( .A(n14755), .ZN(n7546) );
  INV_X1 U9955 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9218) );
  NOR2_X1 U9956 ( .A1(n7547), .A2(n7444), .ZN(n7548) );
  XNOR2_X1 U9957 ( .A(n10545), .B(n8119), .ZN(n7557) );
  NAND2_X1 U9958 ( .A1(n8172), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n7556) );
  NAND2_X1 U9959 ( .A1(n9073), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U9960 ( .A1(n8110), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n7554) );
  INV_X2 U9961 ( .A(n7552), .ZN(n8114) );
  INV_X2 U9962 ( .A(n8114), .ZN(n9050) );
  NAND2_X1 U9963 ( .A1(n9050), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n7553) );
  AND4_X2 U9964 ( .A1(n7556), .A2(n7555), .A3(n7554), .A4(n7553), .ZN(n11625)
         );
  NAND2_X1 U9965 ( .A1(n12869), .A2(n7842), .ZN(n7558) );
  NAND2_X1 U9966 ( .A1(n7557), .A2(n7558), .ZN(n9646) );
  INV_X1 U9967 ( .A(n7557), .ZN(n7560) );
  INV_X1 U9968 ( .A(n7558), .ZN(n7559) );
  NAND2_X1 U9969 ( .A1(n7560), .A2(n7559), .ZN(n7561) );
  AND2_X1 U9970 ( .A1(n9646), .A2(n7561), .ZN(n9580) );
  NAND2_X1 U9971 ( .A1(n8026), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9972 ( .A1(n7562), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7564) );
  XNOR2_X1 U9973 ( .A(n7564), .B(n7563), .ZN(n9388) );
  INV_X1 U9974 ( .A(n7573), .ZN(n7570) );
  MUX2_X1 U9975 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), 
        .S(n9212), .Z(n7569) );
  NAND2_X1 U9976 ( .A1(n7569), .A2(SI_3_), .ZN(n7603) );
  OAI21_X1 U9977 ( .B1(n7569), .B2(SI_3_), .A(n7603), .ZN(n7571) );
  NAND2_X1 U9978 ( .A1(n7570), .A2(n7571), .ZN(n7574) );
  INV_X1 U9979 ( .A(n7571), .ZN(n7572) );
  NAND2_X1 U9980 ( .A1(n7574), .A2(n7639), .ZN(n9832) );
  XNOR2_X1 U9981 ( .A(n9932), .B(n8119), .ZN(n7598) );
  INV_X1 U9982 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9650) );
  NAND2_X1 U9983 ( .A1(n8172), .A2(n9650), .ZN(n7579) );
  NAND2_X1 U9984 ( .A1(n8110), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n7578) );
  INV_X2 U9985 ( .A(n8114), .ZN(n9074) );
  NAND2_X1 U9986 ( .A1(n9074), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9987 ( .A1(n9073), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n7576) );
  NAND4_X1 U9988 ( .A1(n7579), .A2(n7578), .A3(n7577), .A4(n7576), .ZN(n12868)
         );
  NAND2_X1 U9989 ( .A1(n14833), .A2(n12868), .ZN(n7596) );
  XNOR2_X1 U9990 ( .A(n7598), .B(n7596), .ZN(n9693) );
  NAND2_X1 U9991 ( .A1(n7639), .A2(n7603), .ZN(n7582) );
  NAND2_X1 U9992 ( .A1(n7580), .A2(SI_4_), .ZN(n7610) );
  OAI21_X1 U9993 ( .B1(n7580), .B2(SI_4_), .A(n7610), .ZN(n7581) );
  INV_X1 U9994 ( .A(n7581), .ZN(n7606) );
  NAND2_X1 U9995 ( .A1(n7582), .A2(n7606), .ZN(n7611) );
  INV_X4 U9996 ( .A(n9066), .ZN(n9085) );
  NAND2_X1 U9997 ( .A1(n7615), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7585) );
  XNOR2_X1 U9998 ( .A(n7585), .B(P2_IR_REG_4__SCAN_IN), .ZN(n9390) );
  AOI22_X1 U9999 ( .A1(n8026), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n7923), .B2(
        n9390), .ZN(n7586) );
  NAND2_X1 U10000 ( .A1(n9073), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7592) );
  NAND2_X1 U10001 ( .A1(n8110), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7591) );
  NOR2_X1 U10002 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7588) );
  NOR2_X1 U10003 ( .A1(n7621), .A2(n7588), .ZN(n9689) );
  NAND2_X1 U10004 ( .A1(n8172), .A2(n9689), .ZN(n7590) );
  NAND2_X1 U10005 ( .A1(n9050), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n7589) );
  NAND4_X1 U10006 ( .A1(n7592), .A2(n7591), .A3(n7590), .A4(n7589), .ZN(n12867) );
  NAND2_X1 U10007 ( .A1(n14833), .A2(n12867), .ZN(n7593) );
  NAND2_X1 U10008 ( .A1(n7594), .A2(n7593), .ZN(n7601) );
  NAND2_X1 U10009 ( .A1(n7601), .A2(n7595), .ZN(n9695) );
  INV_X1 U10010 ( .A(n7596), .ZN(n7597) );
  AND2_X1 U10011 ( .A1(n7598), .A2(n7597), .ZN(n9692) );
  NAND2_X1 U10012 ( .A1(n7602), .A2(SI_5_), .ZN(n7634) );
  OAI21_X1 U10013 ( .B1(n7602), .B2(SI_5_), .A(n7634), .ZN(n7605) );
  AND2_X1 U10014 ( .A1(n7603), .A2(n7604), .ZN(n7633) );
  NAND2_X1 U10015 ( .A1(n7639), .A2(n7633), .ZN(n7609) );
  INV_X1 U10016 ( .A(n7604), .ZN(n7608) );
  INV_X1 U10017 ( .A(n7605), .ZN(n7612) );
  AND2_X1 U10018 ( .A1(n7612), .A2(n7606), .ZN(n7607) );
  NAND2_X1 U10019 ( .A1(n7609), .A2(n7636), .ZN(n7614) );
  NAND2_X1 U10020 ( .A1(n7614), .A2(n7613), .ZN(n10213) );
  OR2_X1 U10021 ( .A1(n10213), .A2(n9066), .ZN(n7620) );
  INV_X1 U10022 ( .A(n7615), .ZN(n7617) );
  NAND2_X1 U10023 ( .A1(n7617), .A2(n7616), .ZN(n7770) );
  NAND2_X1 U10024 ( .A1(n7770), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7618) );
  XNOR2_X1 U10025 ( .A(n7618), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9391) );
  AOI22_X1 U10026 ( .A1(n8026), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n7923), .B2(
        n9391), .ZN(n7619) );
  XNOR2_X1 U10027 ( .A(n14895), .B(n8119), .ZN(n7627) );
  NAND2_X1 U10028 ( .A1(n9073), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7626) );
  NAND2_X1 U10029 ( .A1(n9050), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n7625) );
  NAND2_X1 U10030 ( .A1(n7621), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7648) );
  OAI21_X1 U10031 ( .B1(n7621), .B2(P2_REG3_REG_5__SCAN_IN), .A(n7648), .ZN(
        n9944) );
  INV_X1 U10032 ( .A(n9944), .ZN(n7622) );
  NAND2_X1 U10033 ( .A1(n8172), .A2(n7622), .ZN(n7624) );
  NAND2_X1 U10034 ( .A1(n8110), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n7623) );
  NAND2_X1 U10035 ( .A1(n12866), .A2(n14833), .ZN(n7628) );
  NAND2_X1 U10036 ( .A1(n7627), .A2(n7628), .ZN(n7632) );
  INV_X1 U10037 ( .A(n7627), .ZN(n7630) );
  INV_X1 U10038 ( .A(n7628), .ZN(n7629) );
  NAND2_X1 U10039 ( .A1(n7630), .A2(n7629), .ZN(n7631) );
  AND2_X1 U10040 ( .A1(n7632), .A2(n7631), .ZN(n9756) );
  AND2_X1 U10041 ( .A1(n7633), .A2(n7634), .ZN(n7638) );
  INV_X1 U10042 ( .A(n7634), .ZN(n7635) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11553), .Z(n7640) );
  NAND2_X1 U10044 ( .A1(n7640), .A2(SI_6_), .ZN(n7659) );
  OAI21_X1 U10045 ( .B1(n7640), .B2(SI_6_), .A(n7659), .ZN(n7641) );
  INV_X1 U10046 ( .A(n7641), .ZN(n7642) );
  OR2_X1 U10047 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  OR2_X1 U10048 ( .A1(n10262), .A2(n9066), .ZN(n7646) );
  NAND2_X1 U10049 ( .A1(n7688), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7667) );
  XNOR2_X1 U10050 ( .A(n7667), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9561) );
  AOI22_X1 U10051 ( .A1(n8026), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n7923), .B2(
        n9561), .ZN(n7645) );
  XNOR2_X1 U10052 ( .A(n10247), .B(n8119), .ZN(n7654) );
  NAND2_X1 U10053 ( .A1(n9073), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7653) );
  NAND2_X1 U10054 ( .A1(n9050), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n7652) );
  INV_X1 U10055 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7647) );
  AND2_X1 U10056 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  NOR2_X1 U10057 ( .A1(n7672), .A2(n7649), .ZN(n9771) );
  NAND2_X1 U10058 ( .A1(n8172), .A2(n9771), .ZN(n7651) );
  NAND2_X1 U10059 ( .A1(n8110), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7650) );
  INV_X1 U10060 ( .A(n10242), .ZN(n12865) );
  NAND2_X1 U10061 ( .A1(n12865), .A2(n14833), .ZN(n7655) );
  XNOR2_X1 U10062 ( .A(n7654), .B(n7655), .ZN(n9769) );
  INV_X1 U10063 ( .A(n7654), .ZN(n7657) );
  INV_X1 U10064 ( .A(n7655), .ZN(n7656) );
  NAND2_X1 U10065 ( .A1(n7657), .A2(n7656), .ZN(n7658) );
  MUX2_X1 U10066 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11553), .Z(n7661) );
  NAND2_X1 U10067 ( .A1(n7661), .A2(SI_7_), .ZN(n7681) );
  OAI21_X1 U10068 ( .B1(n7661), .B2(SI_7_), .A(n7681), .ZN(n7662) );
  INV_X1 U10069 ( .A(n7662), .ZN(n7663) );
  OR2_X1 U10070 ( .A1(n7664), .A2(n7663), .ZN(n7665) );
  NAND2_X1 U10071 ( .A1(n7682), .A2(n7665), .ZN(n10267) );
  NAND2_X1 U10072 ( .A1(n7667), .A2(n7666), .ZN(n7668) );
  NAND2_X1 U10073 ( .A1(n7668), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7669) );
  XNOR2_X1 U10074 ( .A(n7669), .B(P2_IR_REG_7__SCAN_IN), .ZN(n14785) );
  AOI22_X1 U10075 ( .A1(n8026), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n7923), .B2(
        n14785), .ZN(n7670) );
  NAND2_X1 U10076 ( .A1(n7671), .A2(n7670), .ZN(n10443) );
  XNOR2_X1 U10077 ( .A(n10443), .B(n8119), .ZN(n7680) );
  NAND2_X1 U10078 ( .A1(n9050), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n7677) );
  NAND2_X1 U10079 ( .A1(n9073), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n7676) );
  NAND2_X1 U10080 ( .A1(n7672), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7713) );
  OR2_X1 U10081 ( .A1(n7672), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n7673) );
  AND2_X1 U10082 ( .A1(n7713), .A2(n7673), .ZN(n10442) );
  NAND2_X1 U10083 ( .A1(n8172), .A2(n10442), .ZN(n7675) );
  NAND2_X1 U10084 ( .A1(n8110), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7674) );
  NAND4_X1 U10085 ( .A1(n7677), .A2(n7676), .A3(n7675), .A4(n7674), .ZN(n12864) );
  NAND2_X1 U10086 ( .A1(n14833), .A2(n12864), .ZN(n7678) );
  XNOR2_X1 U10087 ( .A(n7680), .B(n7678), .ZN(n9896) );
  INV_X1 U10088 ( .A(n7678), .ZN(n7679) );
  MUX2_X1 U10089 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11553), .Z(n7683) );
  NAND2_X1 U10090 ( .A1(n7683), .A2(SI_8_), .ZN(n7693) );
  OAI21_X1 U10091 ( .B1(n7683), .B2(SI_8_), .A(n7693), .ZN(n7684) );
  INV_X1 U10092 ( .A(n7684), .ZN(n7685) );
  NAND2_X1 U10093 ( .A1(n7686), .A2(n7685), .ZN(n7694) );
  OR2_X1 U10094 ( .A1(n7686), .A2(n7685), .ZN(n7687) );
  NAND2_X1 U10095 ( .A1(n7694), .A2(n7687), .ZN(n10487) );
  OR2_X1 U10096 ( .A1(n10487), .A2(n9066), .ZN(n7691) );
  NAND2_X1 U10097 ( .A1(n7700), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7689) );
  XNOR2_X1 U10098 ( .A(n7689), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9590) );
  AOI22_X1 U10099 ( .A1(n8026), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n7923), .B2(
        n9590), .ZN(n7690) );
  XNOR2_X1 U10100 ( .A(n10470), .B(n7692), .ZN(n10646) );
  NAND2_X1 U10101 ( .A1(n7694), .A2(n7693), .ZN(n7698) );
  MUX2_X1 U10102 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11553), .Z(n7695) );
  NAND2_X1 U10103 ( .A1(n7695), .A2(SI_9_), .ZN(n7725) );
  OAI21_X1 U10104 ( .B1(n7695), .B2(SI_9_), .A(n7725), .ZN(n7696) );
  INV_X1 U10105 ( .A(n7696), .ZN(n7697) );
  NAND2_X1 U10106 ( .A1(n7726), .A2(n7699), .ZN(n10492) );
  OR2_X1 U10107 ( .A1(n10492), .A2(n9066), .ZN(n7707) );
  INV_X1 U10108 ( .A(n7704), .ZN(n7701) );
  NAND2_X1 U10109 ( .A1(n7701), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7702) );
  MUX2_X1 U10110 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7702), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n7705) );
  INV_X1 U10111 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n7703) );
  NAND2_X1 U10112 ( .A1(n7704), .A2(n7703), .ZN(n7751) );
  NAND2_X1 U10113 ( .A1(n7705), .A2(n7751), .ZN(n9591) );
  INV_X1 U10114 ( .A(n9591), .ZN(n9799) );
  AOI22_X1 U10115 ( .A1(n8026), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n7923), .B2(
        n9799), .ZN(n7706) );
  XNOR2_X1 U10116 ( .A(n14923), .B(n7692), .ZN(n7721) );
  NAND2_X1 U10117 ( .A1(n9050), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U10118 ( .A1(n9073), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7710) );
  INV_X1 U10119 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7712) );
  XNOR2_X1 U10120 ( .A(n7737), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n10641) );
  NAND2_X1 U10121 ( .A1(n8172), .A2(n10641), .ZN(n7709) );
  NAND2_X1 U10122 ( .A1(n8110), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U10123 ( .A1(n12862), .A2(n14833), .ZN(n7722) );
  XNOR2_X1 U10124 ( .A(n7721), .B(n7722), .ZN(n10648) );
  NAND2_X1 U10125 ( .A1(n9050), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n7718) );
  NAND2_X1 U10126 ( .A1(n9073), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7717) );
  NAND2_X1 U10127 ( .A1(n7713), .A2(n7712), .ZN(n7714) );
  AND2_X1 U10128 ( .A1(n7737), .A2(n7714), .ZN(n10253) );
  NAND2_X1 U10129 ( .A1(n8172), .A2(n10253), .ZN(n7716) );
  NAND2_X1 U10130 ( .A1(n8110), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n7715) );
  INV_X1 U10131 ( .A(n10475), .ZN(n12863) );
  AND2_X1 U10132 ( .A1(n12863), .A2(n14833), .ZN(n10145) );
  NAND2_X1 U10133 ( .A1(n10645), .A2(n10145), .ZN(n7719) );
  INV_X1 U10134 ( .A(n7721), .ZN(n7723) );
  NAND2_X1 U10135 ( .A1(n7723), .A2(n7722), .ZN(n7724) );
  MUX2_X1 U10136 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11553), .Z(n7727) );
  NAND2_X1 U10137 ( .A1(n7727), .A2(SI_10_), .ZN(n7749) );
  OAI21_X1 U10138 ( .B1(n7727), .B2(SI_10_), .A(n7749), .ZN(n7728) );
  INV_X1 U10139 ( .A(n7728), .ZN(n7729) );
  NAND2_X1 U10140 ( .A1(n7751), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7732) );
  XNOR2_X1 U10141 ( .A(n7732), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U10142 ( .A1(n8026), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7923), 
        .B2(n10137), .ZN(n7733) );
  XNOR2_X1 U10143 ( .A(n10875), .B(n8119), .ZN(n7743) );
  NAND2_X1 U10144 ( .A1(n9050), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7742) );
  NAND2_X1 U10145 ( .A1(n9073), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7741) );
  INV_X1 U10146 ( .A(n7737), .ZN(n7735) );
  AOI21_X1 U10147 ( .B1(n7735), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n7738) );
  NAND2_X1 U10148 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n7736) );
  OR2_X1 U10149 ( .A1(n7738), .A2(n7755), .ZN(n10789) );
  INV_X1 U10150 ( .A(n10789), .ZN(n10589) );
  NAND2_X1 U10151 ( .A1(n8172), .A2(n10589), .ZN(n7740) );
  NAND2_X1 U10152 ( .A1(n8110), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n7739) );
  NAND4_X1 U10153 ( .A1(n7742), .A2(n7741), .A3(n7740), .A4(n7739), .ZN(n12861) );
  AND2_X1 U10154 ( .A1(n14833), .A2(n12861), .ZN(n7744) );
  NAND2_X1 U10155 ( .A1(n7743), .A2(n7744), .ZN(n7748) );
  INV_X1 U10156 ( .A(n7743), .ZN(n10737) );
  INV_X1 U10157 ( .A(n7744), .ZN(n7745) );
  NAND2_X1 U10158 ( .A1(n10737), .A2(n7745), .ZN(n7746) );
  NAND2_X1 U10159 ( .A1(n7748), .A2(n7746), .ZN(n10793) );
  INV_X1 U10160 ( .A(n10793), .ZN(n7747) );
  MUX2_X1 U10161 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11553), .Z(n7766) );
  XNOR2_X1 U10162 ( .A(n7766), .B(SI_11_), .ZN(n7768) );
  XNOR2_X1 U10163 ( .A(n7769), .B(n7768), .ZN(n10912) );
  NAND2_X1 U10164 ( .A1(n10912), .A2(n9085), .ZN(n7754) );
  OAI21_X1 U10165 ( .B1(n7751), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7752) );
  XNOR2_X1 U10166 ( .A(n7752), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10308) );
  AOI22_X1 U10167 ( .A1(n8026), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10308), 
        .B2(n7923), .ZN(n7753) );
  XNOR2_X1 U10168 ( .A(n14942), .B(n8119), .ZN(n7761) );
  NAND2_X1 U10169 ( .A1(n9050), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n7760) );
  NAND2_X1 U10170 ( .A1(n9073), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7759) );
  NOR2_X1 U10171 ( .A1(n7755), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10172 ( .A1(n8172), .A2(n7446), .ZN(n7758) );
  NAND2_X1 U10173 ( .A1(n8110), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7757) );
  NAND4_X1 U10174 ( .A1(n7760), .A2(n7759), .A3(n7758), .A4(n7757), .ZN(n12860) );
  AND2_X1 U10175 ( .A1(n14833), .A2(n12860), .ZN(n7762) );
  NAND2_X1 U10176 ( .A1(n7761), .A2(n7762), .ZN(n7782) );
  INV_X1 U10177 ( .A(n7761), .ZN(n11012) );
  INV_X1 U10178 ( .A(n7762), .ZN(n7763) );
  NAND2_X1 U10179 ( .A1(n11012), .A2(n7763), .ZN(n7764) );
  AND2_X1 U10180 ( .A1(n7782), .A2(n7764), .ZN(n10734) );
  INV_X1 U10181 ( .A(n7766), .ZN(n7767) );
  MUX2_X1 U10182 ( .A(n9643), .B(n9645), .S(n11553), .Z(n7789) );
  XNOR2_X1 U10183 ( .A(n7789), .B(SI_12_), .ZN(n7787) );
  XNOR2_X1 U10184 ( .A(n7788), .B(n7787), .ZN(n10929) );
  NAND2_X1 U10185 ( .A1(n10929), .A2(n9085), .ZN(n7775) );
  INV_X1 U10186 ( .A(n7770), .ZN(n7772) );
  NAND2_X1 U10187 ( .A1(n7772), .A2(n7771), .ZN(n7792) );
  NAND2_X1 U10188 ( .A1(n7792), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7773) );
  XNOR2_X1 U10189 ( .A(n7773), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10696) );
  AOI22_X1 U10190 ( .A1(n8026), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7923), 
        .B2(n10696), .ZN(n7774) );
  XNOR2_X1 U10191 ( .A(n14527), .B(n7692), .ZN(n7783) );
  NAND2_X1 U10192 ( .A1(n9050), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n7781) );
  NAND2_X1 U10193 ( .A1(n9073), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7780) );
  OR2_X1 U10194 ( .A1(n7776), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7777) );
  AND2_X1 U10195 ( .A1(n7796), .A2(n7777), .ZN(n14512) );
  NAND2_X1 U10196 ( .A1(n8172), .A2(n14512), .ZN(n7779) );
  NAND2_X1 U10197 ( .A1(n8110), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7778) );
  NAND2_X1 U10198 ( .A1(n12859), .A2(n7842), .ZN(n7784) );
  XNOR2_X1 U10199 ( .A(n7783), .B(n7784), .ZN(n11015) );
  INV_X1 U10200 ( .A(n7783), .ZN(n7785) );
  NAND2_X1 U10201 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  NAND2_X1 U10202 ( .A1(n7789), .A2(n9244), .ZN(n7790) );
  MUX2_X1 U10203 ( .A(n9707), .B(n12205), .S(n11553), .Z(n7811) );
  XNOR2_X1 U10204 ( .A(n7811), .B(SI_13_), .ZN(n7809) );
  XNOR2_X1 U10205 ( .A(n7810), .B(n7809), .ZN(n11091) );
  NAND2_X1 U10206 ( .A1(n11091), .A2(n9085), .ZN(n7795) );
  OAI21_X1 U10207 ( .B1(n7792), .B2(P2_IR_REG_12__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n7793) );
  XNOR2_X1 U10208 ( .A(n7793), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10868) );
  AOI22_X1 U10209 ( .A1(n8026), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n7923), 
        .B2(n10868), .ZN(n7794) );
  XNOR2_X1 U10210 ( .A(n11152), .B(n8119), .ZN(n7802) );
  NAND2_X1 U10211 ( .A1(n7796), .A2(n10970), .ZN(n7797) );
  AND2_X1 U10212 ( .A1(n7819), .A2(n7797), .ZN(n11139) );
  NAND2_X1 U10213 ( .A1(n11139), .A2(n8172), .ZN(n7801) );
  NAND2_X1 U10214 ( .A1(n9073), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7800) );
  NAND2_X1 U10215 ( .A1(n8110), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7799) );
  NAND2_X1 U10216 ( .A1(n9074), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n7798) );
  NAND4_X1 U10217 ( .A1(n7801), .A2(n7800), .A3(n7799), .A4(n7798), .ZN(n12858) );
  AND2_X1 U10218 ( .A1(n7842), .A2(n12858), .ZN(n7803) );
  NAND2_X1 U10219 ( .A1(n7802), .A2(n7803), .ZN(n7808) );
  INV_X1 U10220 ( .A(n7802), .ZN(n7805) );
  INV_X1 U10221 ( .A(n7803), .ZN(n7804) );
  NAND2_X1 U10222 ( .A1(n7805), .A2(n7804), .ZN(n7806) );
  NAND2_X1 U10223 ( .A1(n7808), .A2(n7806), .ZN(n10964) );
  INV_X1 U10224 ( .A(n10964), .ZN(n7807) );
  NAND2_X1 U10225 ( .A1(n7811), .A2(n9333), .ZN(n7812) );
  MUX2_X1 U10226 ( .A(n9766), .B(n12226), .S(n11553), .Z(n7827) );
  XNOR2_X1 U10227 ( .A(n7827), .B(SI_14_), .ZN(n7813) );
  XNOR2_X1 U10228 ( .A(n7829), .B(n7813), .ZN(n11220) );
  NAND2_X1 U10229 ( .A1(n11220), .A2(n9085), .ZN(n7817) );
  NAND2_X1 U10230 ( .A1(n7814), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7815) );
  XNOR2_X1 U10231 ( .A(n7815), .B(P2_IR_REG_14__SCAN_IN), .ZN(n11185) );
  AOI22_X1 U10232 ( .A1(n8026), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n7923), 
        .B2(n11185), .ZN(n7816) );
  XNOR2_X1 U10233 ( .A(n14520), .B(n7692), .ZN(n7823) );
  NAND2_X1 U10234 ( .A1(n7819), .A2(n7818), .ZN(n7820) );
  NAND2_X1 U10235 ( .A1(n7837), .A2(n7820), .ZN(n14503) );
  AOI22_X1 U10236 ( .A1(n8110), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n9074), .B2(
        P2_REG0_REG_14__SCAN_IN), .ZN(n7822) );
  NAND2_X1 U10237 ( .A1(n9073), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7821) );
  OAI211_X1 U10238 ( .C1(n14503), .C2(n8109), .A(n7822), .B(n7821), .ZN(n12857) );
  NAND2_X1 U10239 ( .A1(n14833), .A2(n12857), .ZN(n7824) );
  XNOR2_X1 U10240 ( .A(n7823), .B(n7824), .ZN(n14492) );
  INV_X1 U10241 ( .A(n7823), .ZN(n7825) );
  NAND2_X1 U10242 ( .A1(n7825), .A2(n7824), .ZN(n7826) );
  NOR2_X1 U10243 ( .A1(n7830), .A2(SI_14_), .ZN(n7828) );
  NAND2_X1 U10244 ( .A1(n7830), .A2(SI_14_), .ZN(n7831) );
  MUX2_X1 U10245 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(P1_DATAO_REG_15__SCAN_IN), 
        .S(n11553), .Z(n7848) );
  XNOR2_X1 U10246 ( .A(n7848), .B(SI_15_), .ZN(n7851) );
  XNOR2_X1 U10247 ( .A(n7852), .B(n7851), .ZN(n11225) );
  NAND2_X1 U10248 ( .A1(n11225), .A2(n9085), .ZN(n7835) );
  NAND2_X1 U10249 ( .A1(n7832), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7833) );
  XNOR2_X1 U10250 ( .A(n7833), .B(P2_IR_REG_15__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U10251 ( .A1(n8026), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n7923), 
        .B2(n11342), .ZN(n7834) );
  XNOR2_X1 U10252 ( .A(n11375), .B(n7692), .ZN(n7845) );
  INV_X1 U10253 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n11195) );
  NAND2_X1 U10254 ( .A1(n7837), .A2(n11195), .ZN(n7838) );
  NAND2_X1 U10255 ( .A1(n7862), .A2(n7838), .ZN(n11285) );
  OR2_X1 U10256 ( .A1(n11285), .A2(n8109), .ZN(n7841) );
  AOI22_X1 U10257 ( .A1(n9074), .A2(P2_REG0_REG_15__SCAN_IN), .B1(n9073), .B2(
        P2_REG1_REG_15__SCAN_IN), .ZN(n7840) );
  NAND2_X1 U10258 ( .A1(n8110), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n7839) );
  NOR2_X1 U10259 ( .A1(n11364), .A2(n8118), .ZN(n7843) );
  NAND2_X1 U10260 ( .A1(n11281), .A2(n7843), .ZN(n11282) );
  INV_X1 U10261 ( .A(n7844), .ZN(n7846) );
  NAND2_X1 U10262 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  INV_X1 U10263 ( .A(n7848), .ZN(n7849) );
  NAND2_X1 U10264 ( .A1(n7849), .A2(n9532), .ZN(n7850) );
  MUX2_X1 U10265 ( .A(n6723), .B(n10180), .S(n11553), .Z(n7873) );
  XNOR2_X1 U10266 ( .A(n7873), .B(SI_16_), .ZN(n7871) );
  XNOR2_X1 U10267 ( .A(n7872), .B(n7871), .ZN(n11418) );
  NAND2_X1 U10268 ( .A1(n11418), .A2(n9085), .ZN(n7859) );
  NOR2_X1 U10269 ( .A1(n7853), .A2(n13281), .ZN(n7854) );
  MUX2_X1 U10270 ( .A(n13281), .B(n7854), .S(P2_IR_REG_16__SCAN_IN), .Z(n7857)
         );
  INV_X1 U10271 ( .A(n7855), .ZN(n7856) );
  OR2_X1 U10272 ( .A1(n7857), .A2(n7856), .ZN(n12874) );
  AOI22_X1 U10273 ( .A1(n8026), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n7923), 
        .B2(n12882), .ZN(n7858) );
  XNOR2_X1 U10274 ( .A(n13258), .B(n7692), .ZN(n11454) );
  INV_X1 U10275 ( .A(n7862), .ZN(n7860) );
  INV_X1 U10276 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U10277 ( .A1(n7862), .A2(n7861), .ZN(n7863) );
  NAND2_X1 U10278 ( .A1(n7882), .A2(n7863), .ZN(n11463) );
  OR2_X1 U10279 ( .A1(n11463), .A2(n8109), .ZN(n7868) );
  INV_X1 U10280 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n11367) );
  NAND2_X1 U10281 ( .A1(n9050), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n7865) );
  NAND2_X1 U10282 ( .A1(n9073), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7864) );
  OAI211_X1 U10283 ( .C1(n11367), .C2(n9078), .A(n7865), .B(n7864), .ZN(n7866)
         );
  INV_X1 U10284 ( .A(n7866), .ZN(n7867) );
  NAND2_X1 U10285 ( .A1(n7868), .A2(n7867), .ZN(n12956) );
  NAND2_X1 U10286 ( .A1(n12956), .A2(n14833), .ZN(n7869) );
  XNOR2_X1 U10287 ( .A(n11454), .B(n7869), .ZN(n11462) );
  NAND2_X1 U10288 ( .A1(n11454), .A2(n7869), .ZN(n7870) );
  NAND2_X1 U10289 ( .A1(n7873), .A2(n12244), .ZN(n7874) );
  MUX2_X1 U10290 ( .A(n7040), .B(n10380), .S(n11553), .Z(n7895) );
  XNOR2_X1 U10291 ( .A(n7895), .B(SI_17_), .ZN(n7876) );
  XNOR2_X1 U10292 ( .A(n7894), .B(n7876), .ZN(n11424) );
  NAND2_X1 U10293 ( .A1(n11424), .A2(n9085), .ZN(n7880) );
  NAND2_X1 U10294 ( .A1(n7855), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7877) );
  MUX2_X1 U10295 ( .A(P2_IR_REG_31__SCAN_IN), .B(n7877), .S(
        P2_IR_REG_17__SCAN_IN), .Z(n7878) );
  OR2_X1 U10296 ( .A1(n7855), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n7899) );
  AND2_X1 U10297 ( .A1(n7878), .A2(n7899), .ZN(n14804) );
  AOI22_X1 U10298 ( .A1(n8026), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n7923), 
        .B2(n14804), .ZN(n7879) );
  XNOR2_X1 U10299 ( .A(n13174), .B(n8119), .ZN(n7892) );
  NAND2_X1 U10300 ( .A1(n7882), .A2(n7881), .ZN(n7883) );
  AND2_X1 U10301 ( .A1(n7905), .A2(n7883), .ZN(n13172) );
  NAND2_X1 U10302 ( .A1(n13172), .A2(n8172), .ZN(n7888) );
  INV_X1 U10303 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12875) );
  NAND2_X1 U10304 ( .A1(n9050), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n7885) );
  NAND2_X1 U10305 ( .A1(n9073), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n7884) );
  OAI211_X1 U10306 ( .C1(n12875), .C2(n9078), .A(n7885), .B(n7884), .ZN(n7886)
         );
  INV_X1 U10307 ( .A(n7886), .ZN(n7887) );
  NOR2_X1 U10308 ( .A1(n12958), .A2(n8118), .ZN(n7890) );
  XNOR2_X1 U10309 ( .A(n7892), .B(n7890), .ZN(n11453) );
  INV_X1 U10310 ( .A(n7890), .ZN(n7891) );
  NAND2_X1 U10311 ( .A1(n7892), .A2(n7891), .ZN(n7893) );
  INV_X1 U10312 ( .A(n7895), .ZN(n7896) );
  NAND2_X1 U10313 ( .A1(n7896), .A2(SI_17_), .ZN(n7897) );
  MUX2_X1 U10314 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n11553), .Z(n7916) );
  XNOR2_X1 U10315 ( .A(n7916), .B(SI_18_), .ZN(n7898) );
  XNOR2_X1 U10316 ( .A(n7917), .B(n7898), .ZN(n11507) );
  NAND2_X1 U10317 ( .A1(n11507), .A2(n9085), .ZN(n7902) );
  NAND2_X1 U10318 ( .A1(n7899), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7900) );
  XNOR2_X1 U10319 ( .A(n7900), .B(P2_IR_REG_18__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U10320 ( .A1(n8026), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n7923), 
        .B2(n12891), .ZN(n7901) );
  XNOR2_X1 U10321 ( .A(n13155), .B(n7692), .ZN(n7912) );
  INV_X1 U10322 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7904) );
  NAND2_X1 U10323 ( .A1(n7905), .A2(n7904), .ZN(n7906) );
  NAND2_X1 U10324 ( .A1(n7927), .A2(n7906), .ZN(n13152) );
  OR2_X1 U10325 ( .A1(n13152), .A2(n8109), .ZN(n7911) );
  INV_X1 U10326 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n12884) );
  NAND2_X1 U10327 ( .A1(n9074), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n7908) );
  NAND2_X1 U10328 ( .A1(n8110), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n7907) );
  OAI211_X1 U10329 ( .C1(n7587), .C2(n12884), .A(n7908), .B(n7907), .ZN(n7909)
         );
  INV_X1 U10330 ( .A(n7909), .ZN(n7910) );
  NOR2_X1 U10331 ( .A1(n12961), .A2(n8118), .ZN(n7913) );
  NAND2_X1 U10332 ( .A1(n7912), .A2(n7913), .ZN(n7934) );
  INV_X1 U10333 ( .A(n7912), .ZN(n12770) );
  INV_X1 U10334 ( .A(n7913), .ZN(n7914) );
  NAND2_X1 U10335 ( .A1(n12770), .A2(n7914), .ZN(n7915) );
  AND2_X1 U10336 ( .A1(n7934), .A2(n7915), .ZN(n12832) );
  NAND2_X1 U10337 ( .A1(n7918), .A2(n12267), .ZN(n7919) );
  MUX2_X1 U10338 ( .A(n10725), .B(n10755), .S(n11553), .Z(n7920) );
  INV_X1 U10339 ( .A(n7920), .ZN(n7921) );
  NAND2_X1 U10340 ( .A1(n7921), .A2(SI_19_), .ZN(n7922) );
  XNOR2_X1 U10341 ( .A(n7940), .B(n7939), .ZN(n11512) );
  NAND2_X1 U10342 ( .A1(n11512), .A2(n9085), .ZN(n7925) );
  AOI22_X1 U10343 ( .A1(n8026), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n7923), 
        .B2(n12903), .ZN(n7924) );
  XNOR2_X1 U10344 ( .A(n13244), .B(n7692), .ZN(n12809) );
  INV_X1 U10345 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7926) );
  NAND2_X1 U10346 ( .A1(n7927), .A2(n7926), .ZN(n7928) );
  AND2_X1 U10347 ( .A1(n7948), .A2(n7928), .ZN(n13140) );
  NAND2_X1 U10348 ( .A1(n13140), .A2(n8172), .ZN(n7933) );
  INV_X1 U10349 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n12240) );
  NAND2_X1 U10350 ( .A1(n8110), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n7930) );
  NAND2_X1 U10351 ( .A1(n7550), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n7929) );
  OAI211_X1 U10352 ( .C1(n8114), .C2(n12240), .A(n7930), .B(n7929), .ZN(n7931)
         );
  INV_X1 U10353 ( .A(n7931), .ZN(n7932) );
  NAND2_X1 U10354 ( .A1(n12930), .A2(n14833), .ZN(n7936) );
  XNOR2_X1 U10355 ( .A(n12809), .B(n7936), .ZN(n12779) );
  AND2_X1 U10356 ( .A1(n12779), .A2(n7934), .ZN(n7935) );
  INV_X1 U10357 ( .A(n12809), .ZN(n7937) );
  NAND2_X1 U10358 ( .A1(n7937), .A2(n7936), .ZN(n7938) );
  NAND2_X1 U10359 ( .A1(n7940), .A2(n7939), .ZN(n7942) );
  INV_X1 U10360 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n11527) );
  MUX2_X1 U10361 ( .A(n11527), .B(n10976), .S(n11553), .Z(n7961) );
  XNOR2_X1 U10362 ( .A(n7963), .B(n7961), .ZN(n11526) );
  NAND2_X1 U10363 ( .A1(n11526), .A2(n9085), .ZN(n7945) );
  OR2_X1 U10364 ( .A1(n7943), .A2(n10976), .ZN(n7944) );
  XNOR2_X1 U10365 ( .A(n13122), .B(n8119), .ZN(n7959) );
  INV_X1 U10366 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n7947) );
  NAND2_X1 U10367 ( .A1(n7948), .A2(n7947), .ZN(n7949) );
  NAND2_X1 U10368 ( .A1(n7971), .A2(n7949), .ZN(n13119) );
  OR2_X1 U10369 ( .A1(n13119), .A2(n8109), .ZN(n7955) );
  INV_X1 U10370 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n7952) );
  NAND2_X1 U10371 ( .A1(n9074), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n7951) );
  NAND2_X1 U10372 ( .A1(n7550), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n7950) );
  OAI211_X1 U10373 ( .C1(n7952), .C2(n9078), .A(n7951), .B(n7950), .ZN(n7953)
         );
  INV_X1 U10374 ( .A(n7953), .ZN(n7954) );
  NOR2_X1 U10375 ( .A1(n12967), .A2(n8118), .ZN(n7957) );
  XNOR2_X1 U10376 ( .A(n7959), .B(n7957), .ZN(n12810) );
  NAND2_X2 U10377 ( .A1(n7956), .A2(n12810), .ZN(n12817) );
  INV_X1 U10378 ( .A(n7957), .ZN(n7958) );
  NAND2_X1 U10379 ( .A1(n7959), .A2(n7958), .ZN(n7960) );
  INV_X1 U10380 ( .A(n7961), .ZN(n7962) );
  INV_X1 U10381 ( .A(n7964), .ZN(n7965) );
  MUX2_X1 U10382 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11553), .Z(n7986) );
  XNOR2_X1 U10383 ( .A(n7986), .B(SI_21_), .ZN(n7983) );
  XNOR2_X1 U10384 ( .A(n7985), .B(n7983), .ZN(n11539) );
  NAND2_X1 U10385 ( .A1(n11539), .A2(n9085), .ZN(n7969) );
  OR2_X1 U10386 ( .A1(n7943), .A2(n11051), .ZN(n7968) );
  XNOR2_X1 U10387 ( .A(n13230), .B(n7692), .ZN(n7978) );
  INV_X1 U10388 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n7970) );
  NAND2_X1 U10389 ( .A1(n7971), .A2(n7970), .ZN(n7972) );
  AND2_X1 U10390 ( .A1(n8009), .A2(n7972), .ZN(n13102) );
  NAND2_X1 U10391 ( .A1(n13102), .A2(n8172), .ZN(n7977) );
  INV_X1 U10392 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n13104) );
  NAND2_X1 U10393 ( .A1(n9074), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n7974) );
  NAND2_X1 U10394 ( .A1(n9073), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n7973) );
  OAI211_X1 U10395 ( .C1(n13104), .C2(n9078), .A(n7974), .B(n7973), .ZN(n7975)
         );
  INV_X1 U10396 ( .A(n7975), .ZN(n7976) );
  NAND2_X1 U10397 ( .A1(n7977), .A2(n7976), .ZN(n12969) );
  NAND2_X1 U10398 ( .A1(n12969), .A2(n14833), .ZN(n7979) );
  XNOR2_X1 U10399 ( .A(n7978), .B(n7979), .ZN(n12787) );
  INV_X1 U10400 ( .A(n7978), .ZN(n7981) );
  INV_X1 U10401 ( .A(n7979), .ZN(n7980) );
  NAND2_X1 U10402 ( .A1(n7981), .A2(n7980), .ZN(n7982) );
  INV_X1 U10403 ( .A(n7983), .ZN(n7984) );
  NAND2_X1 U10404 ( .A1(n7985), .A2(n7984), .ZN(n7988) );
  NAND2_X1 U10405 ( .A1(n7986), .A2(SI_21_), .ZN(n7987) );
  NAND2_X2 U10406 ( .A1(n7988), .A2(n7987), .ZN(n8002) );
  XNOR2_X2 U10407 ( .A(n8002), .B(SI_22_), .ZN(n11554) );
  MUX2_X1 U10408 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n11553), .Z(n8001) );
  XNOR2_X1 U10409 ( .A(n11554), .B(n8001), .ZN(n11201) );
  NAND2_X1 U10410 ( .A1(n11201), .A2(n9085), .ZN(n7990) );
  OR2_X1 U10411 ( .A1(n7943), .A2(n11204), .ZN(n7989) );
  XNOR2_X1 U10412 ( .A(n13226), .B(n8119), .ZN(n12818) );
  XNOR2_X1 U10413 ( .A(n8009), .B(P2_REG3_REG_22__SCAN_IN), .ZN(n13095) );
  NAND2_X1 U10414 ( .A1(n13095), .A2(n8172), .ZN(n7996) );
  INV_X1 U10415 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10416 ( .A1(n9074), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n7992) );
  NAND2_X1 U10417 ( .A1(n7550), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n7991) );
  OAI211_X1 U10418 ( .C1(n7993), .C2(n9078), .A(n7992), .B(n7991), .ZN(n7994)
         );
  INV_X1 U10419 ( .A(n7994), .ZN(n7995) );
  NAND2_X1 U10420 ( .A1(n7996), .A2(n7995), .ZN(n12972) );
  AND2_X1 U10421 ( .A1(n12972), .A2(n14833), .ZN(n7997) );
  INV_X1 U10422 ( .A(n12818), .ZN(n7998) );
  INV_X1 U10423 ( .A(n7997), .ZN(n12820) );
  NAND2_X1 U10424 ( .A1(n7998), .A2(n12820), .ZN(n7999) );
  NAND2_X1 U10425 ( .A1(n8002), .A2(SI_22_), .ZN(n8003) );
  MUX2_X1 U10426 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11553), .Z(n8023) );
  XNOR2_X1 U10427 ( .A(n8023), .B(SI_23_), .ZN(n8021) );
  XNOR2_X1 U10428 ( .A(n8022), .B(n8021), .ZN(n11566) );
  NAND2_X1 U10429 ( .A1(n11566), .A2(n9085), .ZN(n8005) );
  OR2_X1 U10430 ( .A1(n7943), .A2(n11297), .ZN(n8004) );
  XNOR2_X1 U10431 ( .A(n13220), .B(n7692), .ZN(n8017) );
  INV_X1 U10432 ( .A(n8009), .ZN(n8007) );
  AND2_X1 U10433 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_23__SCAN_IN), 
        .ZN(n8006) );
  INV_X1 U10434 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n12824) );
  INV_X1 U10435 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8008) );
  OAI21_X1 U10436 ( .B1(n8009), .B2(n12824), .A(n8008), .ZN(n8010) );
  NAND2_X1 U10437 ( .A1(n8030), .A2(n8010), .ZN(n13078) );
  OR2_X1 U10438 ( .A1(n13078), .A2(n8109), .ZN(n8015) );
  INV_X1 U10439 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n13079) );
  NAND2_X1 U10440 ( .A1(n9074), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n8012) );
  NAND2_X1 U10441 ( .A1(n7550), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n8011) );
  OAI211_X1 U10442 ( .C1(n13079), .C2(n9078), .A(n8012), .B(n8011), .ZN(n8013)
         );
  INV_X1 U10443 ( .A(n8013), .ZN(n8014) );
  NOR2_X1 U10444 ( .A1(n12974), .A2(n8118), .ZN(n8016) );
  NAND2_X1 U10445 ( .A1(n12759), .A2(n8016), .ZN(n12760) );
  INV_X1 U10446 ( .A(n8017), .ZN(n8018) );
  OR2_X1 U10447 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND2_X1 U10448 ( .A1(n8023), .A2(SI_23_), .ZN(n8024) );
  MUX2_X1 U10449 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n11553), .Z(n8045) );
  XNOR2_X1 U10450 ( .A(n8045), .B(SI_24_), .ZN(n8042) );
  XNOR2_X1 U10451 ( .A(n8044), .B(n8042), .ZN(n11499) );
  NAND2_X1 U10452 ( .A1(n11499), .A2(n9085), .ZN(n8028) );
  NAND2_X1 U10453 ( .A1(n8026), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8027) );
  XNOR2_X1 U10454 ( .A(n13054), .B(n7692), .ZN(n8037) );
  INV_X1 U10455 ( .A(n8030), .ZN(n8029) );
  NAND2_X1 U10456 ( .A1(n8029), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n8052) );
  INV_X1 U10457 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n12804) );
  NAND2_X1 U10458 ( .A1(n8030), .A2(n12804), .ZN(n8031) );
  NAND2_X1 U10459 ( .A1(n8052), .A2(n8031), .ZN(n13058) );
  OR2_X1 U10460 ( .A1(n13058), .A2(n8109), .ZN(n8036) );
  INV_X1 U10461 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n13057) );
  NAND2_X1 U10462 ( .A1(n9074), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n8033) );
  NAND2_X1 U10463 ( .A1(n9073), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n8032) );
  OAI211_X1 U10464 ( .C1(n13057), .C2(n9078), .A(n8033), .B(n8032), .ZN(n8034)
         );
  INV_X1 U10465 ( .A(n8034), .ZN(n8035) );
  NOR2_X1 U10466 ( .A1(n12977), .A2(n8118), .ZN(n8038) );
  NAND2_X1 U10467 ( .A1(n8037), .A2(n8038), .ZN(n8041) );
  INV_X1 U10468 ( .A(n8037), .ZN(n12793) );
  INV_X1 U10469 ( .A(n8038), .ZN(n8039) );
  NAND2_X1 U10470 ( .A1(n12793), .A2(n8039), .ZN(n8040) );
  AND2_X1 U10471 ( .A1(n8041), .A2(n8040), .ZN(n12803) );
  NAND2_X1 U10472 ( .A1(n12802), .A2(n12803), .ZN(n12801) );
  NAND2_X1 U10473 ( .A1(n12801), .A2(n8041), .ZN(n8063) );
  INV_X1 U10474 ( .A(n8042), .ZN(n8043) );
  NAND2_X1 U10475 ( .A1(n8045), .A2(SI_24_), .ZN(n8046) );
  INV_X1 U10476 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13302) );
  MUX2_X1 U10477 ( .A(n14251), .B(n13302), .S(n11553), .Z(n8047) );
  INV_X1 U10478 ( .A(SI_25_), .ZN(n11292) );
  NAND2_X1 U10479 ( .A1(n8047), .A2(n11292), .ZN(n8066) );
  INV_X1 U10480 ( .A(n8047), .ZN(n8048) );
  NAND2_X1 U10481 ( .A1(n8048), .A2(SI_25_), .ZN(n8049) );
  NAND2_X1 U10482 ( .A1(n8066), .A2(n8049), .ZN(n8064) );
  XNOR2_X1 U10483 ( .A(n8065), .B(n8064), .ZN(n13299) );
  NAND2_X1 U10484 ( .A1(n13299), .A2(n9085), .ZN(n8051) );
  OR2_X1 U10485 ( .A1(n7943), .A2(n13302), .ZN(n8050) );
  AND2_X2 U10486 ( .A1(n8051), .A2(n8050), .ZN(n13039) );
  XNOR2_X1 U10487 ( .A(n13039), .B(n7692), .ZN(n8059) );
  INV_X1 U10488 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n12797) );
  NAND2_X1 U10489 ( .A1(n8052), .A2(n12797), .ZN(n8053) );
  NAND2_X1 U10490 ( .A1(n8071), .A2(n8053), .ZN(n13043) );
  OR2_X1 U10491 ( .A1(n13043), .A2(n8109), .ZN(n8058) );
  INV_X1 U10492 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n12228) );
  NAND2_X1 U10493 ( .A1(n8110), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n8055) );
  NAND2_X1 U10494 ( .A1(n9073), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n8054) );
  OAI211_X1 U10495 ( .C1(n8114), .C2(n12228), .A(n8055), .B(n8054), .ZN(n8056)
         );
  INV_X1 U10496 ( .A(n8056), .ZN(n8057) );
  NOR2_X1 U10497 ( .A1(n12980), .A2(n8118), .ZN(n8060) );
  NAND2_X1 U10498 ( .A1(n8059), .A2(n8060), .ZN(n8079) );
  INV_X1 U10499 ( .A(n8059), .ZN(n12838) );
  INV_X1 U10500 ( .A(n8060), .ZN(n8061) );
  NAND2_X1 U10501 ( .A1(n12838), .A2(n8061), .ZN(n8062) );
  AND2_X1 U10502 ( .A1(n8079), .A2(n8062), .ZN(n12791) );
  MUX2_X1 U10503 ( .A(n14245), .B(n13297), .S(n11553), .Z(n8085) );
  XNOR2_X1 U10504 ( .A(n8085), .B(SI_26_), .ZN(n8067) );
  XNOR2_X1 U10505 ( .A(n8086), .B(n8067), .ZN(n13296) );
  NAND2_X1 U10506 ( .A1(n13296), .A2(n9085), .ZN(n8069) );
  OR2_X1 U10507 ( .A1(n7943), .A2(n13297), .ZN(n8068) );
  XNOR2_X1 U10508 ( .A(n13028), .B(n8119), .ZN(n8083) );
  INV_X1 U10509 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8070) );
  NAND2_X1 U10510 ( .A1(n8071), .A2(n8070), .ZN(n8072) );
  NAND2_X1 U10511 ( .A1(n13026), .A2(n8172), .ZN(n8078) );
  INV_X1 U10512 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8075) );
  NAND2_X1 U10513 ( .A1(n9074), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n8074) );
  NAND2_X1 U10514 ( .A1(n7550), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n8073) );
  OAI211_X1 U10515 ( .C1(n8075), .C2(n9078), .A(n8074), .B(n8073), .ZN(n8076)
         );
  INV_X1 U10516 ( .A(n8076), .ZN(n8077) );
  NOR2_X1 U10517 ( .A1(n12983), .A2(n8118), .ZN(n8081) );
  XNOR2_X1 U10518 ( .A(n8083), .B(n8081), .ZN(n12850) );
  AND2_X1 U10519 ( .A1(n12850), .A2(n8079), .ZN(n8080) );
  INV_X1 U10520 ( .A(n8081), .ZN(n8082) );
  NAND2_X1 U10521 ( .A1(n8083), .A2(n8082), .ZN(n8084) );
  OAI21_X1 U10522 ( .B1(n8086), .B2(n12745), .A(n8085), .ZN(n8088) );
  NAND2_X1 U10523 ( .A1(n8086), .A2(n12745), .ZN(n8087) );
  MUX2_X1 U10524 ( .A(n7070), .B(n13294), .S(n11553), .Z(n8157) );
  XNOR2_X1 U10525 ( .A(n8157), .B(SI_27_), .ZN(n8089) );
  NAND2_X1 U10526 ( .A1(n13293), .A2(n9085), .ZN(n8091) );
  OR2_X1 U10527 ( .A1(n7943), .A2(n13294), .ZN(n8090) );
  XNOR2_X1 U10528 ( .A(n13196), .B(n8119), .ZN(n8098) );
  XNOR2_X1 U10529 ( .A(n8106), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n13012) );
  NAND2_X1 U10530 ( .A1(n13012), .A2(n8172), .ZN(n8097) );
  INV_X1 U10531 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n8094) );
  NAND2_X1 U10532 ( .A1(n9074), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n8093) );
  NAND2_X1 U10533 ( .A1(n9073), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n8092) );
  OAI211_X1 U10534 ( .C1(n8094), .C2(n9078), .A(n8093), .B(n8092), .ZN(n8095)
         );
  INV_X1 U10535 ( .A(n8095), .ZN(n8096) );
  NAND2_X1 U10536 ( .A1(n8097), .A2(n8096), .ZN(n12985) );
  AND2_X1 U10537 ( .A1(n12985), .A2(n14833), .ZN(n8099) );
  NAND2_X1 U10538 ( .A1(n8098), .A2(n8099), .ZN(n8103) );
  INV_X1 U10539 ( .A(n8098), .ZN(n8101) );
  INV_X1 U10540 ( .A(n8099), .ZN(n8100) );
  NAND2_X1 U10541 ( .A1(n8101), .A2(n8100), .ZN(n8102) );
  NAND2_X1 U10542 ( .A1(n8103), .A2(n8102), .ZN(n12750) );
  NAND2_X1 U10543 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n8104) );
  NOR2_X1 U10544 ( .A1(n8106), .A2(n8104), .ZN(n12953) );
  INV_X1 U10545 ( .A(n12953), .ZN(n8108) );
  INV_X1 U10546 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n12754) );
  INV_X1 U10547 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8105) );
  OAI21_X1 U10548 ( .B1(n8106), .B2(n12754), .A(n8105), .ZN(n8107) );
  NAND2_X1 U10549 ( .A1(n8108), .A2(n8107), .ZN(n8182) );
  INV_X1 U10550 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8113) );
  NAND2_X1 U10551 ( .A1(n8110), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n8112) );
  NAND2_X1 U10552 ( .A1(n9073), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n8111) );
  OAI211_X1 U10553 ( .C1(n8114), .C2(n8113), .A(n8112), .B(n8111), .ZN(n8115)
         );
  INV_X1 U10554 ( .A(n8115), .ZN(n8116) );
  NOR2_X1 U10555 ( .A1(n12943), .A2(n8118), .ZN(n8120) );
  XNOR2_X1 U10556 ( .A(n8120), .B(n8119), .ZN(n8121) );
  INV_X1 U10557 ( .A(n8166), .ZN(n8156) );
  NOR4_X1 U10558 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8131) );
  OR4_X1 U10559 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8128) );
  NOR4_X1 U10560 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8126) );
  NOR4_X1 U10561 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8125) );
  NOR4_X1 U10562 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8124) );
  NOR4_X1 U10563 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8123) );
  NAND4_X1 U10564 ( .A1(n8126), .A2(n8125), .A3(n8124), .A4(n8123), .ZN(n8127)
         );
  NOR4_X1 U10565 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n8128), .A4(n8127), .ZN(n8130) );
  NOR4_X1 U10566 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8129) );
  NAND3_X1 U10567 ( .A1(n8131), .A2(n8130), .A3(n8129), .ZN(n8142) );
  NAND2_X1 U10568 ( .A1(n8132), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8133) );
  MUX2_X1 U10569 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8133), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8134) );
  INV_X1 U10570 ( .A(n8148), .ZN(n13300) );
  NAND2_X1 U10571 ( .A1(n8136), .A2(n8135), .ZN(n8151) );
  OAI21_X1 U10572 ( .B1(n8151), .B2(P2_IR_REG_23__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8137) );
  MUX2_X1 U10573 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8137), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8138) );
  NAND2_X1 U10574 ( .A1(n8138), .A2(n8132), .ZN(n11447) );
  INV_X1 U10575 ( .A(P2_B_REG_SCAN_IN), .ZN(n12911) );
  XOR2_X1 U10576 ( .A(n11447), .B(n12911), .Z(n8139) );
  NAND2_X1 U10577 ( .A1(n13300), .A2(n8139), .ZN(n8141) );
  NAND2_X1 U10578 ( .A1(n6483), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8140) );
  NAND2_X1 U10579 ( .A1(n8142), .A2(n14845), .ZN(n9909) );
  INV_X1 U10580 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14849) );
  NAND2_X1 U10581 ( .A1(n14845), .A2(n14849), .ZN(n8144) );
  INV_X1 U10582 ( .A(n8149), .ZN(n13298) );
  NAND2_X1 U10583 ( .A1(n11447), .A2(n13298), .ZN(n8143) );
  NAND2_X1 U10584 ( .A1(n8144), .A2(n8143), .ZN(n14850) );
  INV_X1 U10585 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14852) );
  NAND2_X1 U10586 ( .A1(n14845), .A2(n14852), .ZN(n8146) );
  NAND2_X1 U10587 ( .A1(n13298), .A2(n13300), .ZN(n8145) );
  NAND2_X1 U10588 ( .A1(n8146), .A2(n8145), .ZN(n14853) );
  NOR2_X1 U10589 ( .A1(n14850), .A2(n14853), .ZN(n8147) );
  NAND2_X1 U10590 ( .A1(n9909), .A2(n8147), .ZN(n8183) );
  NAND2_X1 U10591 ( .A1(n8149), .A2(n8148), .ZN(n8150) );
  NAND2_X1 U10592 ( .A1(n8151), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8153) );
  AND2_X1 U10593 ( .A1(n9377), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8154) );
  NAND2_X1 U10594 ( .A1(n13001), .A2(n7504), .ZN(n9171) );
  NOR2_X1 U10595 ( .A1(n14943), .A2(n9378), .ZN(n8155) );
  NAND2_X1 U10596 ( .A1(n8156), .A2(n14494), .ZN(n8191) );
  INV_X1 U10597 ( .A(n8157), .ZN(n8160) );
  NOR2_X1 U10598 ( .A1(n8160), .A2(SI_27_), .ZN(n8158) );
  NAND2_X1 U10599 ( .A1(n8160), .A2(SI_27_), .ZN(n8161) );
  MUX2_X1 U10600 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n11553), .Z(n9056) );
  XNOR2_X1 U10601 ( .A(n9056), .B(SI_28_), .ZN(n9054) );
  NAND2_X1 U10602 ( .A1(n11975), .A2(n9085), .ZN(n8163) );
  INV_X1 U10603 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n13292) );
  OR2_X1 U10604 ( .A1(n7943), .A2(n13292), .ZN(n8162) );
  INV_X1 U10605 ( .A(n7504), .ZN(n9160) );
  AND2_X1 U10606 ( .A1(n14856), .A2(n9160), .ZN(n9943) );
  NAND2_X1 U10607 ( .A1(n8180), .A2(n9943), .ZN(n8165) );
  NAND2_X1 U10608 ( .A1(n14816), .A2(n12903), .ZN(n11146) );
  INV_X1 U10609 ( .A(n11146), .ZN(n8164) );
  INV_X1 U10610 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8170) );
  NAND2_X1 U10611 ( .A1(n9074), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n8169) );
  NAND2_X1 U10612 ( .A1(n9073), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n8168) );
  OAI211_X1 U10613 ( .C1(n8170), .C2(n9078), .A(n8169), .B(n8168), .ZN(n8171)
         );
  AOI21_X1 U10614 ( .B1(n12953), .B2(n8172), .A(n8171), .ZN(n9088) );
  INV_X1 U10615 ( .A(n9378), .ZN(n8176) );
  NAND2_X1 U10616 ( .A1(n8173), .A2(n8174), .ZN(n9169) );
  NAND2_X1 U10617 ( .A1(n9169), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8175) );
  XNOR2_X1 U10618 ( .A(n8175), .B(P2_IR_REG_28__SCAN_IN), .ZN(n9397) );
  OR2_X1 U10619 ( .A1(n9088), .A2(n12913), .ZN(n8178) );
  NAND2_X1 U10620 ( .A1(n12985), .A2(n12947), .ZN(n8177) );
  NAND2_X1 U10621 ( .A1(n8178), .A2(n8177), .ZN(n12995) );
  INV_X1 U10622 ( .A(n12995), .ZN(n8181) );
  INV_X1 U10623 ( .A(n9171), .ZN(n8179) );
  INV_X1 U10624 ( .A(n8182), .ZN(n13000) );
  NAND2_X1 U10625 ( .A1(n8183), .A2(n11146), .ZN(n8185) );
  NAND2_X1 U10626 ( .A1(n9378), .A2(n9171), .ZN(n9908) );
  AND3_X1 U10627 ( .A1(n9176), .A2(n9377), .A3(n9908), .ZN(n8184) );
  NAND2_X1 U10628 ( .A1(n8185), .A2(n8184), .ZN(n9578) );
  NAND2_X1 U10629 ( .A1(n9578), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14502) );
  AOI22_X1 U10630 ( .A1(n13000), .A2(n12842), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n8186) );
  INV_X1 U10631 ( .A(n8186), .ZN(n8187) );
  INV_X1 U10632 ( .A(P3_REG1_REG_29__SCAN_IN), .ZN(n8795) );
  INV_X1 U10633 ( .A(n8216), .ZN(n8206) );
  INV_X2 U10634 ( .A(n11846), .ZN(n12304) );
  OR2_X1 U10635 ( .A1(n8211), .A2(n12304), .ZN(n9989) );
  NAND2_X1 U10636 ( .A1(n8216), .A2(n8215), .ZN(n8218) );
  XNOR2_X2 U10637 ( .A(n8219), .B(n6622), .ZN(n12736) );
  NAND2_X1 U10638 ( .A1(n11653), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n8228) );
  INV_X1 U10639 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n12684) );
  OR2_X1 U10640 ( .A1(n11655), .A2(n12684), .ZN(n8227) );
  INV_X1 U10641 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n12106) );
  NOR2_X1 U10642 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8340) );
  NAND2_X1 U10643 ( .A1(n8340), .A2(n8339), .ZN(n8358) );
  NAND2_X1 U10644 ( .A1(n8420), .A2(n8419), .ZN(n8422) );
  NAND2_X1 U10645 ( .A1(n8492), .A2(n8491), .ZN(n8507) );
  INV_X1 U10646 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n8519) );
  INV_X1 U10647 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8557) );
  INV_X1 U10648 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12091) );
  NAND2_X1 U10649 ( .A1(n8600), .A2(n12091), .ZN(n8616) );
  INV_X1 U10650 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n12014) );
  INV_X1 U10651 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n12081) );
  NAND2_X1 U10652 ( .A1(n8655), .A2(n12081), .ZN(n8669) );
  INV_X1 U10653 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8911) );
  NOR2_X1 U10654 ( .A1(n8696), .A2(n8911), .ZN(n8221) );
  INV_X1 U10655 ( .A(n12392), .ZN(n8222) );
  OR2_X1 U10656 ( .A1(n6430), .A2(n8222), .ZN(n8226) );
  INV_X1 U10657 ( .A(n8357), .ZN(n8343) );
  INV_X1 U10658 ( .A(n8343), .ZN(n8490) );
  INV_X1 U10659 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n8224) );
  OR2_X1 U10660 ( .A1(n8490), .A2(n8224), .ZN(n8225) );
  AND4_X2 U10661 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(n12000)
         );
  AOI22_X1 U10662 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n11051), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n6752), .ZN(n8612) );
  AOI22_X1 U10663 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n10755), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n10725), .ZN(n8582) );
  AOI22_X1 U10664 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n10457), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n7037), .ZN(n8567) );
  AOI22_X1 U10665 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n10380), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n7040), .ZN(n8552) );
  XNOR2_X1 U10666 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .ZN(n8513) );
  NAND2_X1 U10667 ( .A1(n8261), .A2(n8279), .ZN(n8231) );
  NAND2_X1 U10668 ( .A1(n9204), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8230) );
  NAND2_X1 U10669 ( .A1(n8231), .A2(n8230), .ZN(n8296) );
  XNOR2_X1 U10670 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n8294) );
  NAND2_X1 U10671 ( .A1(n9218), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8232) );
  XNOR2_X1 U10672 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n8311) );
  NAND2_X1 U10673 ( .A1(n9227), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8233) );
  NAND2_X1 U10674 ( .A1(n9229), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8235) );
  NAND2_X1 U10675 ( .A1(n9247), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8236) );
  NAND2_X1 U10676 ( .A1(n9280), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8237) );
  NAND2_X1 U10677 ( .A1(n8429), .A2(n8428), .ZN(n8239) );
  NAND2_X1 U10678 ( .A1(n12253), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8238) );
  NAND2_X1 U10679 ( .A1(n9356), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8240) );
  XNOR2_X1 U10680 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n8447) );
  NAND2_X1 U10681 ( .A1(n9707), .A2(n8242), .ZN(n8243) );
  XNOR2_X1 U10682 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n8500) );
  NAND2_X1 U10683 ( .A1(n9766), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8244) );
  XNOR2_X1 U10684 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .ZN(n8526) );
  NAND2_X1 U10685 ( .A1(n8513), .A2(n8515), .ZN(n8245) );
  NAND2_X1 U10686 ( .A1(n8582), .A2(n8583), .ZN(n8247) );
  NAND2_X1 U10687 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n8248), .ZN(n8250) );
  NAND2_X1 U10688 ( .A1(n8597), .A2(n11527), .ZN(n8249) );
  NAND2_X1 U10689 ( .A1(n8612), .A2(n8613), .ZN(n8251) );
  INV_X1 U10690 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8252) );
  AOI22_X1 U10691 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(
        P1_DATAO_REG_22__SCAN_IN), .B1(n11204), .B2(n8252), .ZN(n8625) );
  INV_X1 U10692 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U10693 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(
        P1_DATAO_REG_23__SCAN_IN), .B1(n11297), .B2(n11567), .ZN(n8638) );
  INV_X1 U10694 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11500) );
  NAND2_X1 U10695 ( .A1(n8651), .A2(n11500), .ZN(n8255) );
  NAND2_X1 U10696 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n8253), .ZN(n8254) );
  NAND2_X1 U10697 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(n13302), .ZN(n8256) );
  AOI22_X1 U10698 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n13297), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n14245), .ZN(n8677) );
  INV_X1 U10699 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14242) );
  AOI22_X1 U10700 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13292), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n14242), .ZN(n8257) );
  INV_X1 U10701 ( .A(n8257), .ZN(n8258) );
  XNOR2_X1 U10702 ( .A(n8704), .B(n8258), .ZN(n12737) );
  NAND2_X1 U10703 ( .A1(n12737), .A2(n8293), .ZN(n8260) );
  INV_X1 U10704 ( .A(SI_28_), .ZN(n12739) );
  OR2_X1 U10705 ( .A1(n8310), .A2(n12739), .ZN(n8259) );
  XNOR2_X1 U10706 ( .A(n8261), .B(n8279), .ZN(n9252) );
  NAND2_X1 U10707 ( .A1(n8430), .A2(n9252), .ZN(n8267) );
  INV_X1 U10708 ( .A(SI_1_), .ZN(n9253) );
  OR2_X1 U10709 ( .A1(n8310), .A2(n9253), .ZN(n8266) );
  NAND2_X1 U10710 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), 
        .ZN(n8262) );
  MUX2_X1 U10711 ( .A(n8262), .B(P3_IR_REG_31__SCAN_IN), .S(n9997), .Z(n8264)
         );
  NAND2_X1 U10712 ( .A1(n8264), .A2(n8263), .ZN(n9974) );
  OR2_X1 U10713 ( .A1(n6425), .A2(n9974), .ZN(n8265) );
  AND3_X2 U10714 ( .A1(n8267), .A2(n8266), .A3(n8265), .ZN(n15100) );
  INV_X1 U10715 ( .A(n15100), .ZN(n10208) );
  INV_X1 U10716 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n8268) );
  OR2_X1 U10717 ( .A1(n11655), .A2(n8268), .ZN(n8273) );
  INV_X1 U10718 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n15115) );
  OR2_X1 U10719 ( .A1(n6429), .A2(n15115), .ZN(n8272) );
  INV_X1 U10720 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n8270) );
  NAND2_X1 U10721 ( .A1(n10087), .A2(n15100), .ZN(n11685) );
  NAND2_X1 U10722 ( .A1(n11686), .A2(n11685), .ZN(n15102) );
  INV_X1 U10723 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9907) );
  INV_X1 U10724 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n8274) );
  INV_X1 U10725 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10782) );
  OR2_X1 U10726 ( .A1(n8490), .A2(n10782), .ZN(n8275) );
  NAND2_X1 U10727 ( .A1(n8269), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8277) );
  INV_X1 U10728 ( .A(n8279), .ZN(n8282) );
  NAND2_X1 U10729 ( .A1(n8280), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8281) );
  NAND2_X1 U10730 ( .A1(n8282), .A2(n8281), .ZN(n9264) );
  NAND2_X1 U10731 ( .A1(n8430), .A2(n9264), .ZN(n8285) );
  OR2_X1 U10732 ( .A1(n8310), .A2(n9515), .ZN(n8284) );
  INV_X1 U10733 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n9994) );
  OR2_X1 U10734 ( .A1(n6425), .A2(n9994), .ZN(n8283) );
  NAND2_X1 U10735 ( .A1(n15102), .A2(n15103), .ZN(n8287) );
  INV_X1 U10736 ( .A(n10087), .ZN(n15088) );
  NAND2_X1 U10737 ( .A1(n15088), .A2(n15100), .ZN(n8286) );
  NAND2_X1 U10738 ( .A1(n8269), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8292) );
  INV_X1 U10739 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n10437) );
  OR2_X1 U10740 ( .A1(n6429), .A2(n10437), .ZN(n8291) );
  INV_X1 U10741 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n8288) );
  OR2_X1 U10742 ( .A1(n11655), .A2(n8288), .ZN(n8290) );
  INV_X1 U10743 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n9998) );
  INV_X1 U10744 ( .A(n8294), .ZN(n8295) );
  XNOR2_X1 U10745 ( .A(n8296), .B(n8295), .ZN(n9271) );
  NAND2_X1 U10746 ( .A1(n11663), .A2(n9271), .ZN(n8300) );
  OR2_X1 U10747 ( .A1(n6425), .A2(n6431), .ZN(n8298) );
  NAND2_X1 U10748 ( .A1(n15105), .A2(n10434), .ZN(n11689) );
  INV_X1 U10749 ( .A(n15105), .ZN(n12283) );
  INV_X1 U10750 ( .A(n10434), .ZN(n15094) );
  INV_X1 U10751 ( .A(n15085), .ZN(n8301) );
  NAND2_X1 U10752 ( .A1(n15083), .A2(n8301), .ZN(n8303) );
  NAND2_X1 U10753 ( .A1(n6670), .A2(n15094), .ZN(n8302) );
  NAND2_X1 U10754 ( .A1(n8269), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8309) );
  OR2_X1 U10755 ( .A1(n6430), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n8308) );
  INV_X1 U10756 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n8304) );
  INV_X1 U10757 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n8305) );
  OR2_X1 U10758 ( .A1(n8710), .A2(n8305), .ZN(n8306) );
  INV_X1 U10759 ( .A(n8311), .ZN(n8312) );
  XNOR2_X1 U10760 ( .A(n8313), .B(n8312), .ZN(n9269) );
  NAND2_X1 U10761 ( .A1(n11663), .A2(n9269), .ZN(n8317) );
  INV_X1 U10762 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10763 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6510), .ZN(n8314) );
  XNOR2_X1 U10764 ( .A(n8315), .B(n8314), .ZN(n9999) );
  OR2_X1 U10765 ( .A1(n6425), .A2(n10082), .ZN(n8316) );
  OAI211_X1 U10766 ( .C1(n8310), .C2(SI_3_), .A(n8317), .B(n8316), .ZN(n10892)
         );
  INV_X1 U10767 ( .A(n11697), .ZN(n8727) );
  NAND2_X1 U10768 ( .A1(n12149), .A2(n10892), .ZN(n11695) );
  AND2_X2 U10769 ( .A1(n8727), .A2(n11695), .ZN(n11815) );
  INV_X1 U10770 ( .A(n10892), .ZN(n15080) );
  NAND2_X1 U10771 ( .A1(n12149), .A2(n15080), .ZN(n8320) );
  NAND2_X1 U10772 ( .A1(n10687), .A2(n8320), .ZN(n10729) );
  NAND2_X1 U10773 ( .A1(n8269), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8326) );
  INV_X1 U10774 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n9993) );
  OR2_X1 U10775 ( .A1(n8490), .A2(n9993), .ZN(n8325) );
  AND2_X1 U10776 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8321) );
  NOR2_X1 U10777 ( .A1(n8340), .A2(n8321), .ZN(n10898) );
  OR2_X1 U10778 ( .A1(n6430), .A2(n10898), .ZN(n8324) );
  INV_X1 U10779 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n8322) );
  OR2_X1 U10780 ( .A1(n11655), .A2(n8322), .ZN(n8323) );
  XNOR2_X1 U10781 ( .A(n8328), .B(n6739), .ZN(n9220) );
  NAND2_X1 U10782 ( .A1(n8430), .A2(n9220), .ZN(n8336) );
  NOR2_X1 U10783 ( .A1(n8331), .A2(n8765), .ZN(n8329) );
  MUX2_X1 U10784 ( .A(n8765), .B(n8329), .S(P3_IR_REG_4__SCAN_IN), .Z(n8333)
         );
  NAND2_X1 U10785 ( .A1(n8331), .A2(n8330), .ZN(n8352) );
  INV_X1 U10786 ( .A(n8352), .ZN(n8332) );
  OR2_X1 U10787 ( .A1(n6425), .A2(n10108), .ZN(n8334) );
  NAND2_X1 U10788 ( .A1(n10685), .A2(n8827), .ZN(n11700) );
  NAND2_X1 U10789 ( .A1(n11704), .A2(n11703), .ZN(n8337) );
  NAND2_X1 U10790 ( .A1(n11700), .A2(n8337), .ZN(n11696) );
  OR2_X1 U10791 ( .A1(n10685), .A2(n11703), .ZN(n8338) );
  NAND2_X1 U10792 ( .A1(n8269), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8348) );
  OR2_X1 U10793 ( .A1(n8340), .A2(n8339), .ZN(n8341) );
  AND2_X1 U10794 ( .A1(n8358), .A2(n8341), .ZN(n15074) );
  OR2_X1 U10795 ( .A1(n6430), .A2(n15074), .ZN(n8347) );
  INV_X1 U10796 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n8342) );
  OR2_X1 U10797 ( .A1(n11655), .A2(n8342), .ZN(n8346) );
  INV_X1 U10798 ( .A(n8343), .ZN(n8710) );
  INV_X1 U10799 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n8344) );
  OR2_X1 U10800 ( .A1(n8710), .A2(n8344), .ZN(n8345) );
  XNOR2_X1 U10801 ( .A(n8350), .B(n6742), .ZN(n9267) );
  NAND2_X1 U10802 ( .A1(n8430), .A2(n9267), .ZN(n8356) );
  NAND2_X1 U10803 ( .A1(n8352), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8351) );
  MUX2_X1 U10804 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8351), .S(
        P3_IR_REG_5__SCAN_IN), .Z(n8353) );
  NAND2_X1 U10805 ( .A1(n8353), .A2(n8472), .ZN(n10003) );
  OR2_X1 U10806 ( .A1(n6425), .A2(n6695), .ZN(n8354) );
  NAND2_X1 U10807 ( .A1(n10747), .A2(n15072), .ZN(n11707) );
  INV_X1 U10808 ( .A(n15072), .ZN(n10984) );
  NAND2_X1 U10809 ( .A1(n12148), .A2(n10984), .ZN(n11699) );
  NAND2_X1 U10810 ( .A1(n11707), .A2(n11699), .ZN(n11698) );
  NAND2_X1 U10811 ( .A1(n11653), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8364) );
  INV_X1 U10812 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n10006) );
  OR2_X1 U10813 ( .A1(n8710), .A2(n10006), .ZN(n8363) );
  NAND2_X1 U10814 ( .A1(n8358), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8359) );
  AND2_X1 U10815 ( .A1(n8374), .A2(n8359), .ZN(n15067) );
  OR2_X1 U10816 ( .A1(n6430), .A2(n15067), .ZN(n8362) );
  INV_X1 U10817 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n8360) );
  OR2_X1 U10818 ( .A1(n11655), .A2(n8360), .ZN(n8361) );
  NAND4_X1 U10819 ( .A1(n8364), .A2(n8363), .A3(n8362), .A4(n8361), .ZN(n12147) );
  XNOR2_X1 U10820 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n8365) );
  XNOR2_X1 U10821 ( .A(n8366), .B(n8365), .ZN(n9261) );
  NAND2_X1 U10822 ( .A1(n8430), .A2(n9261), .ZN(n8371) );
  INV_X1 U10823 ( .A(SI_6_), .ZN(n9262) );
  OR2_X1 U10824 ( .A1(n8310), .A2(n9262), .ZN(n8370) );
  NAND2_X1 U10825 ( .A1(n8472), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8368) );
  INV_X1 U10826 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n8367) );
  XNOR2_X1 U10827 ( .A(n8368), .B(n8367), .ZN(n10354) );
  OR2_X1 U10828 ( .A1(n6425), .A2(n10354), .ZN(n8369) );
  NOR2_X1 U10829 ( .A1(n12147), .A2(n11062), .ZN(n11709) );
  INV_X1 U10830 ( .A(n11709), .ZN(n8728) );
  NAND2_X1 U10831 ( .A1(n12147), .A2(n11062), .ZN(n11702) );
  INV_X1 U10832 ( .A(n11814), .ZN(n11056) );
  INV_X1 U10833 ( .A(n11062), .ZN(n15065) );
  NAND2_X1 U10834 ( .A1(n12147), .A2(n15065), .ZN(n8372) );
  NAND2_X1 U10835 ( .A1(n11055), .A2(n8372), .ZN(n11174) );
  NAND2_X1 U10836 ( .A1(n8269), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8380) );
  INV_X1 U10837 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n8373) );
  OR2_X1 U10838 ( .A1(n8357), .A2(n8373), .ZN(n8379) );
  AND2_X1 U10839 ( .A1(n8374), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8375) );
  NOR2_X1 U10840 ( .A1(n8388), .A2(n8375), .ZN(n15054) );
  OR2_X1 U10841 ( .A1(n6430), .A2(n15054), .ZN(n8378) );
  INV_X1 U10842 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n8376) );
  OR2_X1 U10843 ( .A1(n11655), .A2(n8376), .ZN(n8377) );
  XNOR2_X1 U10844 ( .A(n8382), .B(n8381), .ZN(n9255) );
  NAND2_X1 U10845 ( .A1(n8430), .A2(n9255), .ZN(n8386) );
  OR2_X1 U10846 ( .A1(n8310), .A2(SI_7_), .ZN(n8385) );
  NOR2_X1 U10847 ( .A1(n8472), .A2(P3_IR_REG_6__SCAN_IN), .ZN(n8397) );
  OR2_X1 U10848 ( .A1(n8397), .A2(n8765), .ZN(n8383) );
  XNOR2_X1 U10849 ( .A(n8383), .B(n8396), .ZN(n10388) );
  OR2_X1 U10850 ( .A1(n6425), .A2(n10396), .ZN(n8384) );
  NAND2_X1 U10851 ( .A1(n11210), .A2(n15057), .ZN(n11714) );
  NAND2_X1 U10852 ( .A1(n11174), .A2(n11711), .ZN(n11173) );
  OR2_X1 U10853 ( .A1(n11210), .A2(n11180), .ZN(n8387) );
  NAND2_X1 U10854 ( .A1(n8269), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8394) );
  INV_X1 U10855 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n10391) );
  OR2_X1 U10856 ( .A1(n8710), .A2(n10391), .ZN(n8393) );
  NOR2_X1 U10857 ( .A1(n8388), .A2(n12217), .ZN(n8389) );
  OR2_X1 U10858 ( .A1(n8420), .A2(n8389), .ZN(n12036) );
  INV_X1 U10859 ( .A(n12036), .ZN(n11214) );
  OR2_X1 U10860 ( .A1(n6430), .A2(n11214), .ZN(n8392) );
  INV_X1 U10861 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n8390) );
  OR2_X1 U10862 ( .A1(n11655), .A2(n8390), .ZN(n8391) );
  INV_X1 U10863 ( .A(SI_8_), .ZN(n9215) );
  XNOR2_X1 U10864 ( .A(n8395), .B(n6593), .ZN(n9213) );
  NAND2_X1 U10865 ( .A1(n8430), .A2(n9213), .ZN(n8402) );
  NAND2_X1 U10866 ( .A1(n8397), .A2(n8396), .ZN(n8399) );
  NAND2_X1 U10867 ( .A1(n8399), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8398) );
  MUX2_X1 U10868 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8398), .S(
        P3_IR_REG_8__SCAN_IN), .Z(n8400) );
  NAND2_X1 U10869 ( .A1(n8400), .A2(n8431), .ZN(n10666) );
  OR2_X1 U10870 ( .A1(n6425), .A2(n10666), .ZN(n8401) );
  OAI211_X1 U10871 ( .C1(n8310), .C2(n9215), .A(n8402), .B(n8401), .ZN(n12035)
         );
  INV_X1 U10872 ( .A(n12035), .ZN(n8833) );
  NAND2_X1 U10873 ( .A1(n11399), .A2(n8833), .ZN(n8403) );
  OR2_X1 U10874 ( .A1(n11399), .A2(n8833), .ZN(n11307) );
  NAND2_X1 U10875 ( .A1(n8269), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8410) );
  INV_X1 U10876 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8404) );
  OR2_X1 U10877 ( .A1(n8710), .A2(n8404), .ZN(n8409) );
  NAND2_X1 U10878 ( .A1(n8422), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8405) );
  AND2_X1 U10879 ( .A1(n8440), .A2(n8405), .ZN(n12612) );
  OR2_X1 U10880 ( .A1(n6430), .A2(n12612), .ZN(n8408) );
  INV_X1 U10881 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n8406) );
  OR2_X1 U10882 ( .A1(n11655), .A2(n8406), .ZN(n8407) );
  XNOR2_X1 U10883 ( .A(n8412), .B(n8411), .ZN(n9257) );
  NAND2_X1 U10884 ( .A1(n11663), .A2(n9257), .ZN(n8417) );
  OR2_X1 U10885 ( .A1(n8310), .A2(SI_10_), .ZN(n8416) );
  NAND2_X1 U10886 ( .A1(n8449), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8414) );
  INV_X1 U10887 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n8413) );
  XNOR2_X1 U10888 ( .A(n8414), .B(n8413), .ZN(n12314) );
  INV_X1 U10889 ( .A(n12314), .ZN(n12332) );
  OR2_X1 U10890 ( .A1(n6425), .A2(n12332), .ZN(n8415) );
  NAND2_X1 U10891 ( .A1(n11398), .A2(n12615), .ZN(n11731) );
  INV_X1 U10892 ( .A(n12615), .ZN(n15137) );
  NAND2_X1 U10893 ( .A1(n12143), .A2(n15137), .ZN(n11729) );
  NAND2_X1 U10894 ( .A1(n11731), .A2(n11729), .ZN(n12607) );
  INV_X1 U10895 ( .A(n12607), .ZN(n8436) );
  NAND2_X1 U10896 ( .A1(n8269), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8427) );
  INV_X1 U10897 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n8418) );
  OR2_X1 U10898 ( .A1(n8710), .A2(n8418), .ZN(n8426) );
  OR2_X1 U10899 ( .A1(n8420), .A2(n8419), .ZN(n8421) );
  AND2_X1 U10900 ( .A1(n8422), .A2(n8421), .ZN(n11404) );
  OR2_X1 U10901 ( .A1(n6430), .A2(n11404), .ZN(n8425) );
  INV_X1 U10902 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10903 ( .A1(n11655), .A2(n8423), .ZN(n8424) );
  NAND4_X1 U10904 ( .A1(n8427), .A2(n8426), .A3(n8425), .A4(n8424), .ZN(n12144) );
  XNOR2_X1 U10905 ( .A(n8429), .B(n8428), .ZN(n9250) );
  NAND2_X1 U10906 ( .A1(n8430), .A2(n9250), .ZN(n8435) );
  NAND2_X1 U10907 ( .A1(n8431), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8432) );
  MUX2_X1 U10908 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8432), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n8433) );
  NAND2_X1 U10909 ( .A1(n8433), .A2(n8449), .ZN(n10763) );
  OR2_X1 U10910 ( .A1(n6425), .A2(n10770), .ZN(n8434) );
  INV_X1 U10911 ( .A(n11403), .ZN(n11676) );
  NAND2_X1 U10912 ( .A1(n12144), .A2(n11676), .ZN(n12605) );
  OR2_X1 U10913 ( .A1(n8436), .A2(n12605), .ZN(n8438) );
  OR2_X1 U10914 ( .A1(n11398), .A2(n15137), .ZN(n8437) );
  AND2_X1 U10915 ( .A1(n8438), .A2(n8437), .ZN(n11310) );
  NAND2_X1 U10916 ( .A1(n8269), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8446) );
  INV_X1 U10917 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n8439) );
  OR2_X1 U10918 ( .A1(n8710), .A2(n8439), .ZN(n8445) );
  NAND2_X1 U10919 ( .A1(n8440), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8441) );
  AND2_X1 U10920 ( .A1(n8462), .A2(n8441), .ZN(n11317) );
  OR2_X1 U10921 ( .A1(n6430), .A2(n11317), .ZN(n8444) );
  INV_X1 U10922 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n8442) );
  OR2_X1 U10923 ( .A1(n11655), .A2(n8442), .ZN(n8443) );
  XNOR2_X1 U10924 ( .A(n8448), .B(n8447), .ZN(n9259) );
  NAND2_X1 U10925 ( .A1(n11663), .A2(n9259), .ZN(n8454) );
  OR2_X1 U10926 ( .A1(n8310), .A2(SI_11_), .ZN(n8453) );
  OAI21_X1 U10927 ( .B1(n8449), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8451) );
  INV_X1 U10928 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n8450) );
  XNOR2_X1 U10929 ( .A(n8451), .B(n8450), .ZN(n14982) );
  OR2_X1 U10930 ( .A1(n6425), .A2(n12333), .ZN(n8452) );
  INV_X1 U10931 ( .A(n11316), .ZN(n8734) );
  OR2_X1 U10932 ( .A1(n12611), .A2(n8734), .ZN(n8455) );
  AND2_X1 U10933 ( .A1(n11310), .A2(n8455), .ZN(n8457) );
  AND2_X1 U10934 ( .A1(n11307), .A2(n8457), .ZN(n8456) );
  INV_X1 U10935 ( .A(n8457), .ZN(n8458) );
  XNOR2_X1 U10936 ( .A(n12144), .B(n11403), .ZN(n12603) );
  AND2_X1 U10937 ( .A1(n12603), .A2(n12607), .ZN(n11309) );
  OR2_X1 U10938 ( .A1(n8458), .A2(n11309), .ZN(n8459) );
  NAND2_X1 U10939 ( .A1(n12611), .A2(n8734), .ZN(n8460) );
  NAND2_X1 U10940 ( .A1(n11653), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8468) );
  INV_X1 U10941 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n8461) );
  OR2_X1 U10942 ( .A1(n8710), .A2(n8461), .ZN(n8467) );
  AND2_X1 U10943 ( .A1(n8462), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8463) );
  NOR2_X1 U10944 ( .A1(n8492), .A2(n8463), .ZN(n11389) );
  OR2_X1 U10945 ( .A1(n6430), .A2(n11389), .ZN(n8466) );
  INV_X1 U10946 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n8464) );
  OR2_X1 U10947 ( .A1(n11655), .A2(n8464), .ZN(n8465) );
  NAND4_X1 U10948 ( .A1(n8468), .A2(n8467), .A3(n8466), .A4(n8465), .ZN(n12141) );
  XNOR2_X1 U10949 ( .A(n8469), .B(n6609), .ZN(n9242) );
  NAND2_X1 U10950 ( .A1(n9242), .A2(n8430), .ZN(n8480) );
  INV_X1 U10951 ( .A(n8470), .ZN(n8471) );
  NOR2_X1 U10952 ( .A1(n8472), .A2(n8471), .ZN(n8476) );
  INV_X1 U10953 ( .A(n8476), .ZN(n8473) );
  NAND2_X1 U10954 ( .A1(n8473), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8474) );
  MUX2_X1 U10955 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8474), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n8477) );
  INV_X1 U10956 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10957 ( .A1(n8476), .A2(n8475), .ZN(n8484) );
  NAND2_X1 U10958 ( .A1(n8477), .A2(n8484), .ZN(n15001) );
  OR2_X1 U10959 ( .A1(n6425), .A2(n15001), .ZN(n8479) );
  OR2_X1 U10960 ( .A1(n8310), .A2(n9244), .ZN(n8478) );
  INV_X1 U10961 ( .A(n14477), .ZN(n8481) );
  NAND2_X1 U10962 ( .A1(n12596), .A2(n8481), .ZN(n11736) );
  NAND2_X1 U10963 ( .A1(n12141), .A2(n14477), .ZN(n11735) );
  OR2_X2 U10964 ( .A1(n11382), .A2(n11827), .ZN(n11383) );
  NAND2_X1 U10965 ( .A1(n12141), .A2(n8481), .ZN(n8482) );
  XNOR2_X1 U10966 ( .A(n8483), .B(n12205), .ZN(n9331) );
  NAND2_X1 U10967 ( .A1(n9331), .A2(n8430), .ZN(n8488) );
  NAND2_X1 U10968 ( .A1(n8484), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8485) );
  XNOR2_X1 U10969 ( .A(n8485), .B(P3_IR_REG_13__SCAN_IN), .ZN(n15024) );
  INV_X1 U10970 ( .A(n15024), .ZN(n12339) );
  OAI22_X1 U10971 ( .A1(n8310), .A2(n9333), .B1(n6425), .B2(n12339), .ZN(n8486) );
  INV_X1 U10972 ( .A(n8486), .ZN(n8487) );
  NAND2_X1 U10973 ( .A1(n11653), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8498) );
  INV_X1 U10974 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n8489) );
  OR2_X1 U10975 ( .A1(n8490), .A2(n8489), .ZN(n8497) );
  OR2_X1 U10976 ( .A1(n8492), .A2(n8491), .ZN(n8493) );
  AND2_X1 U10977 ( .A1(n8493), .A2(n8507), .ZN(n12598) );
  OR2_X1 U10978 ( .A1(n6430), .A2(n12598), .ZN(n8496) );
  INV_X1 U10979 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n8494) );
  OR2_X1 U10980 ( .A1(n11655), .A2(n8494), .ZN(n8495) );
  NAND2_X1 U10981 ( .A1(n14475), .A2(n12140), .ZN(n8499) );
  INV_X1 U10982 ( .A(n8500), .ZN(n8501) );
  XNOR2_X1 U10983 ( .A(n8502), .B(n8501), .ZN(n9368) );
  NAND2_X1 U10984 ( .A1(n9368), .A2(n8430), .ZN(n8506) );
  INV_X1 U10985 ( .A(SI_14_), .ZN(n12263) );
  XNOR2_X1 U10986 ( .A(n8503), .B(n7199), .ZN(n15033) );
  OAI22_X1 U10987 ( .A1(n8310), .A2(n12263), .B1(n6425), .B2(n15033), .ZN(
        n8504) );
  INV_X1 U10988 ( .A(n8504), .ZN(n8505) );
  NAND2_X1 U10989 ( .A1(n8506), .A2(n8505), .ZN(n12005) );
  NAND2_X1 U10990 ( .A1(n11653), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8512) );
  INV_X1 U10991 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n12680) );
  OR2_X1 U10992 ( .A1(n8710), .A2(n12680), .ZN(n8511) );
  NAND2_X1 U10993 ( .A1(n8507), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8508) );
  AND2_X1 U10994 ( .A1(n8534), .A2(n8508), .ZN(n12009) );
  OR2_X1 U10995 ( .A1(n6430), .A2(n12009), .ZN(n8510) );
  INV_X1 U10996 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n12722) );
  OR2_X1 U10997 ( .A1(n11655), .A2(n12722), .ZN(n8509) );
  OR2_X1 U10998 ( .A1(n12005), .A2(n12597), .ZN(n11746) );
  NAND2_X1 U10999 ( .A1(n12005), .A2(n12597), .ZN(n11745) );
  INV_X1 U11000 ( .A(n8513), .ZN(n8514) );
  XNOR2_X1 U11001 ( .A(n8515), .B(n8514), .ZN(n9576) );
  OR2_X1 U11002 ( .A1(n8516), .A2(n8765), .ZN(n8517) );
  XNOR2_X1 U11003 ( .A(n8517), .B(P3_IR_REG_16__SCAN_IN), .ZN(n14428) );
  INV_X1 U11004 ( .A(n14428), .ZN(n12322) );
  OAI22_X1 U11005 ( .A1(n8310), .A2(n12244), .B1(n6425), .B2(n12322), .ZN(
        n8518) );
  AOI21_X1 U11006 ( .B1(n9576), .B2(n11663), .A(n8518), .ZN(n12563) );
  NAND2_X1 U11007 ( .A1(n11653), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8524) );
  INV_X1 U11008 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12347) );
  OR2_X1 U11009 ( .A1(n8490), .A2(n12347), .ZN(n8523) );
  NOR2_X1 U11010 ( .A1(n8536), .A2(n8519), .ZN(n8520) );
  OR2_X1 U11011 ( .A1(n8558), .A2(n8520), .ZN(n12561) );
  INV_X1 U11012 ( .A(n12561), .ZN(n12062) );
  OR2_X1 U11013 ( .A1(n6430), .A2(n12062), .ZN(n8522) );
  INV_X1 U11014 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12177) );
  OR2_X1 U11015 ( .A1(n11655), .A2(n12177), .ZN(n8521) );
  NAND4_X1 U11016 ( .A1(n8524), .A2(n8523), .A3(n8522), .A4(n8521), .ZN(n12572) );
  AND2_X1 U11017 ( .A1(n12563), .A2(n12572), .ZN(n11756) );
  INV_X1 U11018 ( .A(n11756), .ZN(n8525) );
  INV_X1 U11019 ( .A(n12563), .ZN(n12670) );
  INV_X1 U11020 ( .A(n12559), .ZN(n8543) );
  INV_X1 U11021 ( .A(n8526), .ZN(n8527) );
  XNOR2_X1 U11022 ( .A(n8528), .B(n8527), .ZN(n9530) );
  NAND2_X1 U11023 ( .A1(n9530), .A2(n8430), .ZN(n8532) );
  NAND2_X1 U11024 ( .A1(n6599), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8529) );
  XNOR2_X1 U11025 ( .A(n8529), .B(P3_IR_REG_15__SCAN_IN), .ZN(n14413) );
  INV_X1 U11026 ( .A(n14413), .ZN(n12344) );
  OAI22_X1 U11027 ( .A1(n8310), .A2(n9532), .B1(n6425), .B2(n12344), .ZN(n8530) );
  INV_X1 U11028 ( .A(n8530), .ZN(n8531) );
  NAND2_X1 U11029 ( .A1(n8532), .A2(n8531), .ZN(n12674) );
  NAND2_X1 U11030 ( .A1(n11653), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8541) );
  INV_X1 U11031 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n8533) );
  OR2_X1 U11032 ( .A1(n8710), .A2(n8533), .ZN(n8540) );
  AND2_X1 U11033 ( .A1(n8534), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8535) );
  NOR2_X1 U11034 ( .A1(n8536), .A2(n8535), .ZN(n12574) );
  OR2_X1 U11035 ( .A1(n6430), .A2(n12574), .ZN(n8539) );
  INV_X1 U11036 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n8537) );
  OR2_X1 U11037 ( .A1(n11655), .A2(n8537), .ZN(n8538) );
  NAND2_X1 U11038 ( .A1(n12674), .A2(n12556), .ZN(n8545) );
  INV_X1 U11039 ( .A(n8545), .ZN(n8542) );
  OR2_X1 U11040 ( .A1(n12674), .A2(n12582), .ZN(n11751) );
  NAND2_X1 U11041 ( .A1(n12674), .A2(n12582), .ZN(n11750) );
  INV_X1 U11042 ( .A(n12576), .ZN(n11829) );
  OR2_X1 U11043 ( .A1(n8542), .A2(n11829), .ZN(n12553) );
  AND2_X1 U11044 ( .A1(n8543), .A2(n12553), .ZN(n8544) );
  INV_X1 U11045 ( .A(n8544), .ZN(n8546) );
  NAND2_X1 U11046 ( .A1(n12005), .A2(n12570), .ZN(n12566) );
  AND2_X1 U11047 ( .A1(n12566), .A2(n8545), .ZN(n12552) );
  OR2_X1 U11048 ( .A1(n8546), .A2(n12552), .ZN(n8547) );
  OR2_X1 U11049 ( .A1(n12563), .A2(n12070), .ZN(n8549) );
  XOR2_X1 U11050 ( .A(n8552), .B(n8551), .Z(n9655) );
  NAND2_X1 U11051 ( .A1(n8570), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8554) );
  INV_X1 U11052 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n8553) );
  XNOR2_X1 U11053 ( .A(n8554), .B(n8553), .ZN(n12349) );
  OAI22_X1 U11054 ( .A1(n8310), .A2(n9653), .B1(n6425), .B2(n12349), .ZN(n8555) );
  AOI21_X1 U11055 ( .B1(n9655), .B2(n11663), .A(n8555), .ZN(n12546) );
  NAND2_X1 U11056 ( .A1(n11653), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8564) );
  INV_X1 U11057 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n8556) );
  OR2_X1 U11058 ( .A1(n8490), .A2(n8556), .ZN(n8563) );
  NOR2_X1 U11059 ( .A1(n8558), .A2(n8557), .ZN(n8559) );
  NOR2_X1 U11060 ( .A1(n8576), .A2(n8559), .ZN(n12547) );
  OR2_X1 U11061 ( .A1(n6430), .A2(n12547), .ZN(n8562) );
  INV_X1 U11062 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n8560) );
  OR2_X1 U11063 ( .A1(n11655), .A2(n8560), .ZN(n8561) );
  NAND4_X1 U11064 ( .A1(n8564), .A2(n8563), .A3(n8562), .A4(n8561), .ZN(n12557) );
  AND2_X1 U11065 ( .A1(n12546), .A2(n12557), .ZN(n11762) );
  INV_X1 U11066 ( .A(n11762), .ZN(n8565) );
  INV_X1 U11067 ( .A(n12546), .ZN(n12666) );
  INV_X1 U11068 ( .A(n12557), .ZN(n12527) );
  NAND2_X1 U11069 ( .A1(n12666), .A2(n12527), .ZN(n12532) );
  NAND2_X1 U11070 ( .A1(n8565), .A2(n12532), .ZN(n11830) );
  NAND2_X1 U11071 ( .A1(n12666), .A2(n12557), .ZN(n8566) );
  INV_X1 U11072 ( .A(n8567), .ZN(n8568) );
  XNOR2_X1 U11073 ( .A(n8569), .B(n8568), .ZN(n14377) );
  NAND2_X1 U11074 ( .A1(n14377), .A2(n11663), .ZN(n8575) );
  OAI21_X1 U11075 ( .B1(n8570), .B2(P3_IR_REG_17__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8572) );
  INV_X1 U11076 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n8571) );
  XNOR2_X1 U11077 ( .A(n8572), .B(n8571), .ZN(n14379) );
  OAI22_X1 U11078 ( .A1(n8310), .A2(n12267), .B1(n6425), .B2(n14379), .ZN(
        n8573) );
  INV_X1 U11079 ( .A(n8573), .ZN(n8574) );
  NAND2_X1 U11080 ( .A1(n11653), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8581) );
  INV_X1 U11081 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12715) );
  OR2_X1 U11082 ( .A1(n11655), .A2(n12715), .ZN(n8580) );
  OR2_X1 U11083 ( .A1(n8576), .A2(n12106), .ZN(n8577) );
  AND2_X1 U11084 ( .A1(n8577), .A2(n8591), .ZN(n12529) );
  OR2_X1 U11085 ( .A1(n12529), .A2(n6430), .ZN(n8579) );
  INV_X1 U11086 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12664) );
  OR2_X1 U11087 ( .A1(n8710), .A2(n12664), .ZN(n8578) );
  NAND2_X1 U11088 ( .A1(n12539), .A2(n12511), .ZN(n11765) );
  INV_X1 U11089 ( .A(n12525), .ZN(n12534) );
  XNOR2_X1 U11090 ( .A(n8583), .B(n8582), .ZN(n9810) );
  NAND2_X1 U11091 ( .A1(n9810), .A2(n11663), .ZN(n8590) );
  INV_X1 U11092 ( .A(n8584), .ZN(n8585) );
  NAND2_X1 U11093 ( .A1(n8585), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8586) );
  MUX2_X1 U11094 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8586), .S(
        P3_IR_REG_19__SCAN_IN), .Z(n8587) );
  OAI22_X1 U11095 ( .A1(n8310), .A2(SI_19_), .B1(n12375), .B2(n6425), .ZN(
        n8588) );
  INV_X1 U11096 ( .A(n8588), .ZN(n8589) );
  NAND2_X1 U11097 ( .A1(n11653), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8596) );
  INV_X1 U11098 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n12711) );
  OR2_X1 U11099 ( .A1(n11655), .A2(n12711), .ZN(n8595) );
  AND2_X1 U11100 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(n8591), .ZN(n8592) );
  NOR2_X1 U11101 ( .A1(n8600), .A2(n8592), .ZN(n12515) );
  OR2_X1 U11102 ( .A1(n6430), .A2(n12515), .ZN(n8594) );
  INV_X1 U11103 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n12658) );
  OR2_X1 U11104 ( .A1(n8490), .A2(n12658), .ZN(n8593) );
  NAND4_X1 U11105 ( .A1(n8596), .A2(n8595), .A3(n8594), .A4(n8593), .ZN(n12498) );
  INV_X1 U11106 ( .A(n12498), .ZN(n12528) );
  OR2_X1 U11107 ( .A1(n12713), .A2(n12528), .ZN(n12493) );
  NAND2_X1 U11108 ( .A1(n12534), .A2(n12493), .ZN(n8611) );
  XNOR2_X1 U11109 ( .A(n8597), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n10365) );
  NAND2_X1 U11110 ( .A1(n10365), .A2(n8430), .ZN(n8599) );
  INV_X1 U11111 ( .A(SI_20_), .ZN(n10366) );
  NAND2_X1 U11112 ( .A1(n11653), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n8607) );
  OR2_X1 U11113 ( .A1(n8600), .A2(n12091), .ZN(n8601) );
  AND2_X1 U11114 ( .A1(n8601), .A2(n8616), .ZN(n12502) );
  OR2_X1 U11115 ( .A1(n6430), .A2(n12502), .ZN(n8606) );
  INV_X1 U11116 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n8602) );
  OR2_X1 U11117 ( .A1(n11655), .A2(n8602), .ZN(n8605) );
  INV_X1 U11118 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n8603) );
  OR2_X1 U11119 ( .A1(n8490), .A2(n8603), .ZN(n8604) );
  XNOR2_X1 U11120 ( .A(n12505), .B(n12510), .ZN(n12494) );
  AND2_X1 U11121 ( .A1(n12713), .A2(n12498), .ZN(n11770) );
  INV_X1 U11122 ( .A(n11770), .ZN(n8608) );
  NAND2_X1 U11123 ( .A1(n8608), .A2(n11769), .ZN(n12519) );
  OR2_X1 U11124 ( .A1(n12539), .A2(n12543), .ZN(n12492) );
  NAND2_X1 U11125 ( .A1(n12519), .A2(n12492), .ZN(n8609) );
  NAND2_X1 U11126 ( .A1(n8609), .A2(n12493), .ZN(n8610) );
  XOR2_X1 U11127 ( .A(n8613), .B(n8612), .Z(n10615) );
  NAND2_X1 U11128 ( .A1(n10615), .A2(n11663), .ZN(n8615) );
  INV_X1 U11129 ( .A(SI_21_), .ZN(n10617) );
  OR2_X1 U11130 ( .A1(n8310), .A2(n10617), .ZN(n8614) );
  NAND2_X1 U11131 ( .A1(n11653), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n8621) );
  INV_X1 U11132 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12649) );
  OR2_X1 U11133 ( .A1(n8357), .A2(n12649), .ZN(n8620) );
  NAND2_X1 U11134 ( .A1(n8616), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8617) );
  AND2_X1 U11135 ( .A1(n8630), .A2(n8617), .ZN(n12044) );
  OR2_X1 U11136 ( .A1(n6430), .A2(n12044), .ZN(n8619) );
  INV_X1 U11137 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12706) );
  OR2_X1 U11138 ( .A1(n11655), .A2(n12706), .ZN(n8618) );
  NAND2_X1 U11139 ( .A1(n12708), .A2(n12470), .ZN(n8622) );
  NAND2_X1 U11140 ( .A1(n12480), .A2(n8622), .ZN(n8624) );
  NAND2_X1 U11141 ( .A1(n11776), .A2(n12499), .ZN(n8623) );
  XNOR2_X1 U11142 ( .A(n8626), .B(n8625), .ZN(n10656) );
  NAND2_X1 U11143 ( .A1(n10656), .A2(n11663), .ZN(n8629) );
  INV_X1 U11144 ( .A(SI_22_), .ZN(n8627) );
  OR2_X1 U11145 ( .A1(n8310), .A2(n8627), .ZN(n8628) );
  NAND2_X1 U11146 ( .A1(n11653), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n8635) );
  INV_X1 U11147 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12702) );
  OR2_X1 U11148 ( .A1(n11655), .A2(n12702), .ZN(n8634) );
  AND2_X1 U11149 ( .A1(n8630), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8631) );
  NOR2_X1 U11150 ( .A1(n8642), .A2(n8631), .ZN(n12097) );
  OR2_X1 U11151 ( .A1(n6430), .A2(n12097), .ZN(n8633) );
  INV_X1 U11152 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12645) );
  OR2_X1 U11153 ( .A1(n8357), .A2(n12645), .ZN(n8632) );
  INV_X1 U11154 ( .A(n12482), .ZN(n12138) );
  OR2_X1 U11155 ( .A1(n12472), .A2(n12138), .ZN(n8636) );
  NAND2_X1 U11156 ( .A1(n12472), .A2(n12138), .ZN(n8637) );
  XNOR2_X1 U11157 ( .A(n8639), .B(n8638), .ZN(n10797) );
  NAND2_X1 U11158 ( .A1(n10797), .A2(n8430), .ZN(n8641) );
  INV_X1 U11159 ( .A(SI_23_), .ZN(n10799) );
  OR2_X1 U11160 ( .A1(n8310), .A2(n10799), .ZN(n8640) );
  NAND2_X1 U11161 ( .A1(n11653), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n8647) );
  INV_X1 U11162 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12698) );
  OR2_X1 U11163 ( .A1(n11655), .A2(n12698), .ZN(n8646) );
  NOR2_X1 U11164 ( .A1(n8642), .A2(n12014), .ZN(n8643) );
  OR2_X1 U11165 ( .A1(n8655), .A2(n8643), .ZN(n12461) );
  INV_X1 U11166 ( .A(n12461), .ZN(n12017) );
  OR2_X1 U11167 ( .A1(n6430), .A2(n12017), .ZN(n8645) );
  INV_X1 U11168 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12641) );
  OR2_X1 U11169 ( .A1(n8357), .A2(n12641), .ZN(n8644) );
  NAND4_X1 U11170 ( .A1(n8647), .A2(n8646), .A3(n8645), .A4(n8644), .ZN(n12441) );
  NAND2_X1 U11171 ( .A1(n12700), .A2(n12441), .ZN(n12445) );
  NAND2_X1 U11172 ( .A1(n12019), .A2(n12471), .ZN(n8648) );
  NAND2_X1 U11173 ( .A1(n12445), .A2(n8648), .ZN(n12459) );
  NAND2_X1 U11174 ( .A1(n12019), .A2(n12441), .ZN(n8649) );
  XNOR2_X1 U11175 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n8651), .ZN(n11205) );
  NAND2_X1 U11176 ( .A1(n11205), .A2(n8430), .ZN(n8653) );
  INV_X1 U11177 ( .A(SI_24_), .ZN(n11207) );
  OR2_X1 U11178 ( .A1(n8310), .A2(n11207), .ZN(n8652) );
  NAND2_X1 U11179 ( .A1(n11653), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n8661) );
  INV_X1 U11180 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n8654) );
  OR2_X1 U11181 ( .A1(n8710), .A2(n8654), .ZN(n8660) );
  OR2_X1 U11182 ( .A1(n8655), .A2(n12081), .ZN(n8656) );
  AND2_X1 U11183 ( .A1(n8669), .A2(n8656), .ZN(n12449) );
  OR2_X1 U11184 ( .A1(n6430), .A2(n12449), .ZN(n8659) );
  INV_X1 U11185 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n8657) );
  OR2_X1 U11186 ( .A1(n11655), .A2(n8657), .ZN(n8658) );
  NAND4_X1 U11187 ( .A1(n8661), .A2(n8660), .A3(n8659), .A4(n8658), .ZN(n12137) );
  NOR2_X1 U11188 ( .A1(n12638), .A2(n12456), .ZN(n8662) );
  NAND2_X1 U11189 ( .A1(n12638), .A2(n12456), .ZN(n8663) );
  AOI22_X1 U11190 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(
        P1_DATAO_REG_25__SCAN_IN), .B1(n13302), .B2(n14251), .ZN(n8665) );
  XNOR2_X1 U11191 ( .A(n8666), .B(n8665), .ZN(n11291) );
  NAND2_X1 U11192 ( .A1(n11291), .A2(n8430), .ZN(n8668) );
  OR2_X1 U11193 ( .A1(n8310), .A2(n11292), .ZN(n8667) );
  NAND2_X1 U11194 ( .A1(n11653), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n8675) );
  INV_X1 U11195 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12187) );
  OR2_X1 U11196 ( .A1(n8357), .A2(n12187), .ZN(n8674) );
  NAND2_X1 U11197 ( .A1(n8669), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8670) );
  AND2_X1 U11198 ( .A1(n8681), .A2(n8670), .ZN(n12429) );
  OR2_X1 U11199 ( .A1(n6430), .A2(n12429), .ZN(n8673) );
  INV_X1 U11200 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n8671) );
  OR2_X1 U11201 ( .A1(n11655), .A2(n8671), .ZN(n8672) );
  OR2_X1 U11202 ( .A1(n12631), .A2(n12421), .ZN(n11791) );
  NAND2_X1 U11203 ( .A1(n12631), .A2(n12421), .ZN(n11792) );
  NAND2_X1 U11204 ( .A1(n12631), .A2(n12442), .ZN(n8676) );
  XNOR2_X1 U11205 ( .A(n8678), .B(n8677), .ZN(n12743) );
  NAND2_X1 U11206 ( .A1(n12743), .A2(n8430), .ZN(n8680) );
  OR2_X1 U11207 ( .A1(n8310), .A2(n12745), .ZN(n8679) );
  NAND2_X1 U11208 ( .A1(n11653), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n8687) );
  INV_X1 U11209 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12692) );
  OR2_X1 U11210 ( .A1(n11655), .A2(n12692), .ZN(n8686) );
  NAND2_X1 U11211 ( .A1(n8681), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8682) );
  NAND2_X1 U11212 ( .A1(n8694), .A2(n8682), .ZN(n12423) );
  INV_X1 U11213 ( .A(n12423), .ZN(n8683) );
  OR2_X1 U11214 ( .A1(n6430), .A2(n8683), .ZN(n8685) );
  INV_X1 U11215 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12629) );
  OR2_X1 U11216 ( .A1(n8357), .A2(n12629), .ZN(n8684) );
  OR2_X1 U11217 ( .A1(n12422), .A2(n12404), .ZN(n8688) );
  NAND2_X1 U11218 ( .A1(n12422), .A2(n12404), .ZN(n8689) );
  AOI22_X1 U11219 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n13294), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n7070), .ZN(n8691) );
  INV_X1 U11220 ( .A(SI_27_), .ZN(n12741) );
  OR2_X1 U11221 ( .A1(n8310), .A2(n12741), .ZN(n8693) );
  NAND2_X1 U11222 ( .A1(n11653), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n8700) );
  INV_X1 U11223 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12688) );
  OR2_X1 U11224 ( .A1(n11655), .A2(n12688), .ZN(n8699) );
  AND2_X1 U11225 ( .A1(n8694), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8695) );
  NOR2_X1 U11226 ( .A1(n8696), .A2(n8695), .ZN(n12409) );
  OR2_X1 U11227 ( .A1(n6430), .A2(n12409), .ZN(n8698) );
  INV_X1 U11228 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n12625) );
  OR2_X1 U11229 ( .A1(n8710), .A2(n12625), .ZN(n8697) );
  NAND4_X1 U11230 ( .A1(n8700), .A2(n8699), .A3(n8698), .A4(n8697), .ZN(n12388) );
  NAND2_X1 U11231 ( .A1(n12690), .A2(n12388), .ZN(n8701) );
  NAND2_X1 U11232 ( .A1(n12412), .A2(n12420), .ZN(n12383) );
  NAND2_X1 U11233 ( .A1(n8701), .A2(n12383), .ZN(n11800) );
  NAND2_X1 U11234 ( .A1(n12690), .A2(n12420), .ZN(n8702) );
  XNOR2_X2 U11235 ( .A(n8703), .B(n12000), .ZN(n12386) );
  OAI21_X1 U11236 ( .B1(n12686), .B2(n12000), .A(n12385), .ZN(n8714) );
  NAND2_X1 U11237 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n13292), .ZN(n8705) );
  AOI22_X1 U11238 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n14242), .B1(n8705), 
        .B2(n8704), .ZN(n11650) );
  INV_X1 U11239 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n13463) );
  OAI22_X1 U11240 ( .A1(n13463), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n13285), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11649) );
  INV_X1 U11241 ( .A(n11649), .ZN(n8706) );
  XNOR2_X1 U11242 ( .A(n11650), .B(n8706), .ZN(n12733) );
  NAND2_X1 U11243 ( .A1(n12733), .A2(n8293), .ZN(n8708) );
  INV_X1 U11244 ( .A(SI_29_), .ZN(n12734) );
  OR2_X1 U11245 ( .A1(n8310), .A2(n12734), .ZN(n8707) );
  NAND2_X1 U11246 ( .A1(n8708), .A2(n8707), .ZN(n8796) );
  INV_X1 U11247 ( .A(n14459), .ZN(n8709) );
  NAND2_X1 U11248 ( .A1(n11653), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8713) );
  INV_X1 U11249 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8811) );
  OR2_X1 U11250 ( .A1(n11655), .A2(n8811), .ZN(n8712) );
  OR2_X1 U11251 ( .A1(n8710), .A2(n8795), .ZN(n8711) );
  NAND4_X1 U11252 ( .A1(n11659), .A2(n8713), .A3(n8712), .A4(n8711), .ZN(
        n12389) );
  INV_X1 U11253 ( .A(n12389), .ZN(n8908) );
  OR2_X1 U11254 ( .A1(n8796), .A2(n8908), .ZN(n11810) );
  NAND2_X1 U11255 ( .A1(n8796), .A2(n8908), .ZN(n11807) );
  NAND2_X1 U11256 ( .A1(n11810), .A2(n11807), .ZN(n11836) );
  NAND2_X1 U11257 ( .A1(n11848), .A2(n12375), .ZN(n8801) );
  NAND2_X1 U11258 ( .A1(n8715), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8716) );
  MUX2_X1 U11259 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8716), .S(
        P3_IR_REG_20__SCAN_IN), .Z(n8718) );
  NAND2_X1 U11260 ( .A1(n11682), .A2(n8800), .ZN(n11675) );
  NAND2_X1 U11261 ( .A1(n9989), .A2(n6425), .ZN(n8719) );
  INV_X1 U11262 ( .A(P3_B_REG_SCAN_IN), .ZN(n8720) );
  OR2_X1 U11263 ( .A1(n8211), .A2(n8720), .ZN(n8721) );
  NAND2_X1 U11264 ( .A1(n12571), .A2(n8721), .ZN(n14456) );
  NAND2_X1 U11265 ( .A1(n11653), .A2(P3_REG2_REG_30__SCAN_IN), .ZN(n8725) );
  INV_X1 U11266 ( .A(P3_REG1_REG_30__SCAN_IN), .ZN(n14471) );
  OR2_X1 U11267 ( .A1(n8357), .A2(n14471), .ZN(n8724) );
  INV_X1 U11268 ( .A(P3_REG0_REG_30__SCAN_IN), .ZN(n8722) );
  OR2_X1 U11269 ( .A1(n11655), .A2(n8722), .ZN(n8723) );
  NAND4_X1 U11270 ( .A1(n11659), .A2(n8725), .A3(n8724), .A4(n8723), .ZN(
        n12136) );
  INV_X1 U11271 ( .A(n12136), .ZN(n11665) );
  NAND2_X1 U11272 ( .A1(n8817), .A2(n11686), .ZN(n15086) );
  NAND2_X1 U11273 ( .A1(n15086), .A2(n15085), .ZN(n15084) );
  NAND2_X1 U11274 ( .A1(n15084), .A2(n11689), .ZN(n10682) );
  NAND2_X1 U11275 ( .A1(n10681), .A2(n8727), .ZN(n10727) );
  INV_X1 U11276 ( .A(n11696), .ZN(n11817) );
  NAND2_X1 U11277 ( .A1(n10727), .A2(n11817), .ZN(n10726) );
  NAND2_X1 U11278 ( .A1(n10977), .A2(n11707), .ZN(n11053) );
  NAND2_X1 U11279 ( .A1(n11052), .A2(n8728), .ZN(n11172) );
  INV_X1 U11280 ( .A(n11711), .ZN(n11821) );
  NAND2_X1 U11281 ( .A1(n11399), .A2(n12035), .ZN(n11722) );
  NAND2_X1 U11282 ( .A1(n12145), .A2(n8833), .ZN(n11721) );
  NAND2_X1 U11283 ( .A1(n11722), .A2(n11721), .ZN(n11718) );
  INV_X1 U11284 ( .A(n11718), .ZN(n11820) );
  NAND2_X1 U11285 ( .A1(n12144), .A2(n11403), .ZN(n8729) );
  AND2_X1 U11286 ( .A1(n11820), .A2(n8729), .ZN(n8731) );
  INV_X1 U11287 ( .A(n8729), .ZN(n8730) );
  INV_X1 U11288 ( .A(n12144), .ZN(n12610) );
  NAND2_X1 U11289 ( .A1(n12610), .A2(n11676), .ZN(n8732) );
  NAND2_X1 U11290 ( .A1(n12611), .A2(n11316), .ZN(n11730) );
  NAND2_X1 U11291 ( .A1(n12142), .A2(n8734), .ZN(n11728) );
  NAND2_X1 U11292 ( .A1(n11730), .A2(n11728), .ZN(n11732) );
  NAND2_X1 U11293 ( .A1(n8735), .A2(n11730), .ZN(n11388) );
  NAND2_X1 U11294 ( .A1(n14475), .A2(n12581), .ZN(n11740) );
  INV_X1 U11295 ( .A(n11740), .ZN(n8736) );
  OR2_X1 U11296 ( .A1(n14475), .A2(n12581), .ZN(n11741) );
  AND2_X1 U11297 ( .A1(n6970), .A2(n11760), .ZN(n8742) );
  INV_X1 U11298 ( .A(n11760), .ZN(n8741) );
  AND2_X1 U11299 ( .A1(n12525), .A2(n12532), .ZN(n12531) );
  AOI21_X2 U11300 ( .B1(n12545), .B2(n8742), .A(n7451), .ZN(n12520) );
  NAND2_X1 U11301 ( .A1(n12651), .A2(n12139), .ZN(n8743) );
  NAND2_X1 U11302 ( .A1(n12708), .A2(n12499), .ZN(n8744) );
  NAND2_X1 U11303 ( .A1(n12472), .A2(n12482), .ZN(n11780) );
  NAND2_X1 U11304 ( .A1(n12466), .A2(n11780), .ZN(n8745) );
  INV_X1 U11305 ( .A(n12459), .ZN(n8746) );
  NAND2_X1 U11306 ( .A1(n12638), .A2(n12137), .ZN(n11786) );
  INV_X1 U11307 ( .A(n12638), .ZN(n12085) );
  NAND2_X1 U11308 ( .A1(n12085), .A2(n12456), .ZN(n11785) );
  AND2_X1 U11309 ( .A1(n12447), .A2(n12445), .ZN(n8747) );
  NAND2_X1 U11310 ( .A1(n12444), .A2(n8747), .ZN(n12446) );
  NAND2_X1 U11311 ( .A1(n12446), .A2(n11785), .ZN(n12428) );
  NAND2_X1 U11312 ( .A1(n12428), .A2(n12431), .ZN(n8748) );
  NAND2_X1 U11313 ( .A1(n12422), .A2(n12433), .ZN(n11796) );
  INV_X1 U11314 ( .A(n12383), .ZN(n8749) );
  AOI21_X1 U11315 ( .B1(n8703), .B2(n12000), .A(n8749), .ZN(n11803) );
  NOR2_X1 U11316 ( .A1(n8703), .A2(n12000), .ZN(n11802) );
  NAND2_X1 U11317 ( .A1(n11848), .A2(n10368), .ZN(n8750) );
  NAND2_X1 U11318 ( .A1(n8750), .A2(n12375), .ZN(n8751) );
  NAND2_X1 U11319 ( .A1(n8751), .A2(n10616), .ZN(n8753) );
  INV_X1 U11320 ( .A(n11848), .ZN(n11679) );
  OAI21_X1 U11321 ( .B1(n8800), .B2(n11682), .A(n11679), .ZN(n8752) );
  NAND2_X1 U11322 ( .A1(n8753), .A2(n8752), .ZN(n8896) );
  NAND2_X1 U11323 ( .A1(n10368), .A2(n12363), .ZN(n11843) );
  INV_X1 U11324 ( .A(n11843), .ZN(n8754) );
  NAND3_X1 U11325 ( .A1(n8896), .A2(n8754), .A3(n15138), .ZN(n8755) );
  NAND3_X1 U11326 ( .A1(n11848), .A2(n8800), .A3(n12363), .ZN(n8789) );
  XNOR2_X1 U11327 ( .A(n8759), .B(P3_B_REG_SCAN_IN), .ZN(n8762) );
  NOR2_X1 U11328 ( .A1(n8757), .A2(n8765), .ZN(n8760) );
  NOR2_X1 U11329 ( .A1(n8763), .A2(n8765), .ZN(n8764) );
  OAI22_X2 U11330 ( .A1(n9330), .A2(P3_D_REG_0__SCAN_IN), .B1(n6649), .B2(
        n8759), .ZN(n9282) );
  INV_X1 U11331 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n8769) );
  NAND2_X1 U11332 ( .A1(n8780), .A2(n8769), .ZN(n8771) );
  INV_X1 U11333 ( .A(n8783), .ZN(n11294) );
  NAND2_X1 U11334 ( .A1(n12749), .A2(n11294), .ZN(n8770) );
  NAND2_X1 U11335 ( .A1(n9282), .A2(n10183), .ZN(n8804) );
  NOR2_X1 U11336 ( .A1(P3_D_REG_30__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .ZN(
        n8775) );
  NOR4_X1 U11337 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_28__SCAN_IN), .A4(P3_D_REG_22__SCAN_IN), .ZN(n8774) );
  NOR4_X1 U11338 ( .A1(P3_D_REG_18__SCAN_IN), .A2(P3_D_REG_27__SCAN_IN), .A3(
        P3_D_REG_24__SCAN_IN), .A4(P3_D_REG_29__SCAN_IN), .ZN(n8773) );
  NOR4_X1 U11339 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_25__SCAN_IN), .A3(
        P3_D_REG_20__SCAN_IN), .A4(P3_D_REG_19__SCAN_IN), .ZN(n8772) );
  NAND4_X1 U11340 ( .A1(n8775), .A2(n8774), .A3(n8773), .A4(n8772), .ZN(n8782)
         );
  NOR4_X1 U11341 ( .A1(P3_D_REG_12__SCAN_IN), .A2(P3_D_REG_11__SCAN_IN), .A3(
        P3_D_REG_26__SCAN_IN), .A4(P3_D_REG_9__SCAN_IN), .ZN(n8779) );
  NOR4_X1 U11342 ( .A1(P3_D_REG_14__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_21__SCAN_IN), .ZN(n8778) );
  NOR4_X1 U11343 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8777) );
  NOR4_X1 U11344 ( .A1(P3_D_REG_15__SCAN_IN), .A2(P3_D_REG_13__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8776) );
  NAND4_X1 U11345 ( .A1(n8779), .A2(n8778), .A3(n8777), .A4(n8776), .ZN(n8781)
         );
  NAND2_X1 U11346 ( .A1(n8783), .A2(n8759), .ZN(n8784) );
  INV_X1 U11347 ( .A(n8785), .ZN(n8786) );
  NAND2_X1 U11348 ( .A1(n8786), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8787) );
  AND2_X1 U11349 ( .A1(n8802), .A2(n8918), .ZN(n8788) );
  NAND2_X1 U11350 ( .A1(n11808), .A2(n8789), .ZN(n10182) );
  NAND2_X1 U11351 ( .A1(n11804), .A2(n11843), .ZN(n10185) );
  AND2_X1 U11352 ( .A1(n10182), .A2(n10185), .ZN(n8793) );
  NAND2_X1 U11353 ( .A1(n11848), .A2(n12363), .ZN(n8790) );
  OAI21_X1 U11354 ( .B1(n15138), .B2(n8800), .A(n8790), .ZN(n8791) );
  AOI21_X1 U11355 ( .B1(n8791), .B2(n11843), .A(n11804), .ZN(n8792) );
  MUX2_X1 U11356 ( .A(n8793), .B(n8792), .S(n10183), .Z(n8794) );
  INV_X1 U11357 ( .A(n8796), .ZN(n12379) );
  INV_X1 U11358 ( .A(n12682), .ZN(n8797) );
  NAND2_X1 U11359 ( .A1(n8799), .A2(n8802), .ZN(n8916) );
  NAND2_X1 U11360 ( .A1(n10616), .A2(n8800), .ZN(n11841) );
  OR2_X1 U11361 ( .A1(n11841), .A2(n8801), .ZN(n8897) );
  INV_X1 U11362 ( .A(n8802), .ZN(n8803) );
  INV_X1 U11363 ( .A(n8896), .ZN(n8805) );
  OAI22_X1 U11364 ( .A1(n8916), .A2(n8897), .B1(n8910), .B2(n8805), .ZN(n8806)
         );
  NAND2_X1 U11365 ( .A1(n8806), .A2(n8918), .ZN(n8809) );
  INV_X1 U11366 ( .A(n8916), .ZN(n8807) );
  NOR2_X1 U11367 ( .A1(n9971), .A2(n11843), .ZN(n8909) );
  AND2_X1 U11368 ( .A1(n8909), .A2(n11804), .ZN(n8904) );
  NAND2_X1 U11369 ( .A1(n8807), .A2(n8904), .ZN(n8808) );
  INV_X1 U11370 ( .A(n12724), .ZN(n8812) );
  NAND2_X1 U11371 ( .A1(n8796), .A2(n8812), .ZN(n8813) );
  NAND2_X1 U11372 ( .A1(n8814), .A2(n8813), .ZN(P3_U3456) );
  OAI21_X1 U11373 ( .B1(n11682), .B2(n12363), .A(n10368), .ZN(n8815) );
  XNOR2_X1 U11374 ( .A(n12638), .B(n10202), .ZN(n12078) );
  XNOR2_X1 U11375 ( .A(n12700), .B(n8852), .ZN(n8884) );
  INV_X1 U11376 ( .A(n15103), .ZN(n8816) );
  XNOR2_X1 U11377 ( .A(n10087), .B(n15100), .ZN(n8818) );
  XNOR2_X1 U11378 ( .A(n8852), .B(n15100), .ZN(n8820) );
  NAND2_X1 U11379 ( .A1(n8820), .A2(n15088), .ZN(n8821) );
  NAND2_X1 U11380 ( .A1(n10204), .A2(n8821), .ZN(n10430) );
  XNOR2_X1 U11381 ( .A(n8822), .B(n6670), .ZN(n10431) );
  XNOR2_X1 U11382 ( .A(n6427), .B(n10892), .ZN(n8825) );
  INV_X1 U11383 ( .A(n12149), .ZN(n15087) );
  XNOR2_X1 U11384 ( .A(n8825), .B(n15087), .ZN(n10529) );
  INV_X1 U11385 ( .A(n8822), .ZN(n8823) );
  NAND2_X1 U11386 ( .A1(n8823), .A2(n6670), .ZN(n10526) );
  AND2_X1 U11387 ( .A1(n10529), .A2(n10526), .ZN(n8824) );
  NAND2_X1 U11388 ( .A1(n8825), .A2(n12149), .ZN(n8826) );
  XNOR2_X1 U11389 ( .A(n8852), .B(n8827), .ZN(n8828) );
  NAND2_X1 U11390 ( .A1(n11704), .A2(n8828), .ZN(n8830) );
  INV_X1 U11391 ( .A(n8828), .ZN(n8829) );
  NAND2_X1 U11392 ( .A1(n8829), .A2(n10685), .ZN(n8832) );
  NAND2_X1 U11393 ( .A1(n8830), .A2(n8832), .ZN(n10745) );
  XNOR2_X1 U11394 ( .A(n8852), .B(n15072), .ZN(n8834) );
  XNOR2_X1 U11395 ( .A(n8834), .B(n10747), .ZN(n10801) );
  XNOR2_X1 U11396 ( .A(n11711), .B(n8852), .ZN(n8839) );
  XNOR2_X1 U11397 ( .A(n8833), .B(n10202), .ZN(n8840) );
  XNOR2_X1 U11398 ( .A(n8840), .B(n11399), .ZN(n8837) );
  INV_X1 U11399 ( .A(n8834), .ZN(n8835) );
  NAND2_X1 U11400 ( .A1(n8835), .A2(n10747), .ZN(n10955) );
  XNOR2_X1 U11401 ( .A(n8852), .B(n11062), .ZN(n10957) );
  INV_X1 U11402 ( .A(n12147), .ZN(n10803) );
  NAND2_X1 U11403 ( .A1(n10957), .A2(n10803), .ZN(n8836) );
  INV_X1 U11404 ( .A(n10957), .ZN(n8838) );
  NAND2_X1 U11405 ( .A1(n8838), .A2(n12147), .ZN(n11105) );
  OAI21_X1 U11406 ( .B1(n12031), .B2(n11105), .A(n8839), .ZN(n8842) );
  OAI21_X1 U11407 ( .B1(n11210), .B2(n12031), .A(n12029), .ZN(n8841) );
  XNOR2_X1 U11408 ( .A(n10202), .B(n11403), .ZN(n8845) );
  XNOR2_X1 U11409 ( .A(n8845), .B(n12144), .ZN(n11069) );
  INV_X1 U11410 ( .A(n11069), .ZN(n8844) );
  XNOR2_X1 U11411 ( .A(n8852), .B(n12615), .ZN(n8848) );
  XNOR2_X1 U11412 ( .A(n8848), .B(n11398), .ZN(n11023) );
  INV_X1 U11413 ( .A(n8845), .ZN(n8846) );
  NAND2_X1 U11414 ( .A1(n8846), .A2(n12610), .ZN(n11024) );
  AND2_X1 U11415 ( .A1(n11023), .A2(n11024), .ZN(n8847) );
  NAND2_X1 U11416 ( .A1(n12143), .A2(n8848), .ZN(n8849) );
  XNOR2_X1 U11417 ( .A(n10202), .B(n11316), .ZN(n11162) );
  NAND2_X1 U11418 ( .A1(n11162), .A2(n12611), .ZN(n8851) );
  NOR2_X1 U11419 ( .A1(n11162), .A2(n12611), .ZN(n8850) );
  XNOR2_X1 U11420 ( .A(n8852), .B(n14477), .ZN(n8853) );
  NAND2_X1 U11421 ( .A1(n8853), .A2(n12596), .ZN(n8856) );
  INV_X1 U11422 ( .A(n8853), .ZN(n8854) );
  NAND2_X1 U11423 ( .A1(n8854), .A2(n12141), .ZN(n8855) );
  AND2_X1 U11424 ( .A1(n8856), .A2(n8855), .ZN(n11256) );
  NAND2_X1 U11425 ( .A1(n11255), .A2(n11256), .ZN(n11254) );
  XNOR2_X1 U11426 ( .A(n14475), .B(n10202), .ZN(n8857) );
  INV_X1 U11427 ( .A(n8857), .ZN(n8858) );
  NAND2_X1 U11428 ( .A1(n8858), .A2(n12140), .ZN(n11299) );
  XNOR2_X1 U11429 ( .A(n12005), .B(n10202), .ZN(n8859) );
  XNOR2_X1 U11430 ( .A(n8859), .B(n12570), .ZN(n12007) );
  NAND2_X1 U11431 ( .A1(n12008), .A2(n12007), .ZN(n12006) );
  INV_X1 U11432 ( .A(n8859), .ZN(n8860) );
  NAND2_X1 U11433 ( .A1(n8860), .A2(n12570), .ZN(n8861) );
  XNOR2_X1 U11434 ( .A(n12674), .B(n10202), .ZN(n12123) );
  NAND2_X1 U11435 ( .A1(n12123), .A2(n12582), .ZN(n8862) );
  INV_X1 U11436 ( .A(n12123), .ZN(n8863) );
  NAND2_X1 U11437 ( .A1(n8863), .A2(n12556), .ZN(n8864) );
  XNOR2_X1 U11438 ( .A(n12563), .B(n10202), .ZN(n12057) );
  AND2_X1 U11439 ( .A1(n12057), .A2(n12572), .ZN(n8865) );
  INV_X1 U11440 ( .A(n12057), .ZN(n8866) );
  NAND2_X1 U11441 ( .A1(n8866), .A2(n12070), .ZN(n8867) );
  XNOR2_X1 U11442 ( .A(n12546), .B(n10202), .ZN(n8868) );
  XNOR2_X1 U11443 ( .A(n8868), .B(n12557), .ZN(n12066) );
  NAND2_X1 U11444 ( .A1(n8868), .A2(n12557), .ZN(n8869) );
  NAND2_X1 U11445 ( .A1(n12068), .A2(n8869), .ZN(n12105) );
  XNOR2_X1 U11446 ( .A(n12539), .B(n10202), .ZN(n8870) );
  XNOR2_X1 U11447 ( .A(n8870), .B(n12543), .ZN(n12104) );
  NAND2_X1 U11448 ( .A1(n12105), .A2(n12104), .ZN(n12103) );
  INV_X1 U11449 ( .A(n8870), .ZN(n8871) );
  NAND2_X1 U11450 ( .A1(n8871), .A2(n12543), .ZN(n8872) );
  NAND2_X1 U11451 ( .A1(n12103), .A2(n8872), .ZN(n12024) );
  XNOR2_X1 U11452 ( .A(n12713), .B(n10202), .ZN(n8873) );
  XNOR2_X1 U11453 ( .A(n8873), .B(n12528), .ZN(n12023) );
  NAND2_X1 U11454 ( .A1(n12024), .A2(n12023), .ZN(n12022) );
  NAND2_X1 U11455 ( .A1(n8873), .A2(n12498), .ZN(n8874) );
  NAND2_X1 U11456 ( .A1(n12022), .A2(n8874), .ZN(n12090) );
  XNOR2_X1 U11457 ( .A(n12505), .B(n10202), .ZN(n8875) );
  XNOR2_X1 U11458 ( .A(n8875), .B(n12139), .ZN(n12089) );
  INV_X1 U11459 ( .A(n8875), .ZN(n8876) );
  NAND2_X1 U11460 ( .A1(n8876), .A2(n12139), .ZN(n8877) );
  XNOR2_X1 U11461 ( .A(n11776), .B(n10202), .ZN(n8878) );
  XNOR2_X1 U11462 ( .A(n8878), .B(n12499), .ZN(n12042) );
  INV_X1 U11463 ( .A(n8878), .ZN(n8879) );
  NAND2_X1 U11464 ( .A1(n8879), .A2(n12499), .ZN(n8880) );
  XNOR2_X1 U11465 ( .A(n12472), .B(n6427), .ZN(n8881) );
  INV_X1 U11466 ( .A(n8881), .ZN(n8882) );
  INV_X1 U11467 ( .A(n12078), .ZN(n8886) );
  OAI21_X1 U11468 ( .B1(n12075), .B2(n12441), .A(n12137), .ZN(n8885) );
  NAND2_X1 U11469 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  XNOR2_X1 U11470 ( .A(n12631), .B(n10202), .ZN(n8889) );
  XNOR2_X1 U11471 ( .A(n8889), .B(n12421), .ZN(n12051) );
  INV_X1 U11472 ( .A(n12051), .ZN(n8888) );
  XNOR2_X1 U11473 ( .A(n12422), .B(n10202), .ZN(n8892) );
  XNOR2_X1 U11474 ( .A(n12690), .B(n10202), .ZN(n8893) );
  XNOR2_X1 U11475 ( .A(n8893), .B(n12388), .ZN(n11999) );
  XNOR2_X1 U11476 ( .A(n12386), .B(n10202), .ZN(n8894) );
  NAND2_X1 U11477 ( .A1(n8896), .A2(n15138), .ZN(n10085) );
  OAI22_X1 U11478 ( .A1(n8916), .A2(n10085), .B1(n8910), .B2(n8897), .ZN(n8895) );
  NAND2_X1 U11479 ( .A1(n8916), .A2(n8896), .ZN(n8900) );
  INV_X1 U11480 ( .A(n8897), .ZN(n8898) );
  NAND2_X1 U11481 ( .A1(n8910), .A2(n8898), .ZN(n8899) );
  NAND4_X1 U11482 ( .A1(n8900), .A2(n9203), .A3(n10185), .A4(n8899), .ZN(n8901) );
  NAND2_X1 U11483 ( .A1(n8901), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8906) );
  INV_X1 U11484 ( .A(n9968), .ZN(n8902) );
  NAND2_X1 U11485 ( .A1(n8902), .A2(P3_STATE_REG_SCAN_IN), .ZN(n11851) );
  INV_X1 U11486 ( .A(n11851), .ZN(n8903) );
  AOI21_X1 U11487 ( .B1(n8910), .B2(n8904), .A(n8903), .ZN(n8905) );
  NAND2_X1 U11488 ( .A1(n8909), .A2(n12571), .ZN(n8907) );
  NOR2_X1 U11489 ( .A1(n8908), .A2(n12109), .ZN(n8913) );
  NAND2_X1 U11490 ( .A1(n8909), .A2(n12569), .ZN(n11847) );
  OAI22_X1 U11491 ( .A1(n12420), .A2(n12126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8911), .ZN(n8912) );
  AOI211_X1 U11492 ( .C1(n12392), .C2(n12117), .A(n8913), .B(n8912), .ZN(n8914) );
  INV_X1 U11493 ( .A(n8914), .ZN(n8920) );
  NAND2_X1 U11494 ( .A1(n8918), .A2(n14476), .ZN(n8915) );
  OR2_X1 U11495 ( .A1(n8916), .A2(n8915), .ZN(n8919) );
  NOR2_X1 U11496 ( .A1(n15138), .A2(n15113), .ZN(n8917) );
  INV_X1 U11497 ( .A(n13230), .ZN(n8922) );
  INV_X1 U11498 ( .A(n12969), .ZN(n12935) );
  OAI22_X1 U11499 ( .A1(n8922), .A2(n9080), .B1(n12935), .B2(n9043), .ZN(n9030) );
  AND2_X1 U11500 ( .A1(n8924), .A2(n8923), .ZN(n8933) );
  INV_X1 U11501 ( .A(n9136), .ZN(n8927) );
  OAI21_X1 U11502 ( .B1(n9129), .B2(n13001), .A(n6485), .ZN(n8925) );
  OAI21_X1 U11503 ( .B1(n12872), .B2(n9091), .A(n8925), .ZN(n8926) );
  NOR2_X1 U11504 ( .A1(n8927), .A2(n8926), .ZN(n8930) );
  NAND2_X1 U11505 ( .A1(n14831), .A2(n9128), .ZN(n8928) );
  OAI21_X1 U11506 ( .B1(n9136), .B2(n9091), .A(n8928), .ZN(n8929) );
  INV_X1 U11507 ( .A(n8931), .ZN(n8932) );
  NAND2_X1 U11508 ( .A1(n8934), .A2(n8933), .ZN(n8935) );
  NAND2_X1 U11509 ( .A1(n8936), .A2(n8935), .ZN(n8942) );
  NAND2_X1 U11510 ( .A1(n6433), .A2(n8937), .ZN(n8939) );
  NAND2_X1 U11511 ( .A1(n8942), .A2(n8943), .ZN(n8941) );
  BUF_X1 U11512 ( .A(n6433), .Z(n9092) );
  INV_X4 U11513 ( .A(n6433), .ZN(n9043) );
  OAI22_X1 U11514 ( .A1(n10545), .A2(n9092), .B1(n11625), .B2(n9043), .ZN(
        n8940) );
  INV_X1 U11515 ( .A(n8942), .ZN(n8945) );
  INV_X1 U11516 ( .A(n8943), .ZN(n8944) );
  INV_X1 U11517 ( .A(n12868), .ZN(n9931) );
  OAI22_X1 U11518 ( .A1(n14879), .A2(n9043), .B1(n9931), .B2(n9092), .ZN(n8946) );
  INV_X1 U11519 ( .A(n10177), .ZN(n14887) );
  INV_X1 U11520 ( .A(n12867), .ZN(n9934) );
  OAI22_X1 U11521 ( .A1(n14887), .A2(n9092), .B1(n9934), .B2(n9043), .ZN(n8948) );
  NAND2_X1 U11522 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  OAI22_X1 U11523 ( .A1(n14895), .A2(n9043), .B1(n10155), .B2(n9080), .ZN(
        n8953) );
  OAI22_X1 U11524 ( .A1(n10247), .A2(n9043), .B1(n10242), .B2(n9080), .ZN(
        n8957) );
  OAI22_X1 U11525 ( .A1(n10247), .A2(n9092), .B1(n10242), .B2(n9043), .ZN(
        n8955) );
  AOI21_X1 U11526 ( .B1(n8958), .B2(n8957), .A(n8956), .ZN(n8959) );
  AOI22_X1 U11527 ( .A1(n10443), .A2(n9091), .B1(n12864), .B2(n9080), .ZN(
        n8963) );
  AOI22_X1 U11528 ( .A1(n10443), .A2(n9080), .B1(n9091), .B2(n12864), .ZN(
        n8961) );
  NAND2_X1 U11529 ( .A1(n8964), .A2(n8963), .ZN(n8965) );
  NAND2_X1 U11530 ( .A1(n8966), .A2(n8965), .ZN(n8969) );
  OAI22_X1 U11531 ( .A1(n10470), .A2(n9043), .B1(n10475), .B2(n9080), .ZN(
        n8968) );
  AOI22_X1 U11532 ( .A1(n14916), .A2(n9091), .B1(n12863), .B2(n9080), .ZN(
        n8967) );
  OAI22_X1 U11533 ( .A1(n14923), .A2(n9092), .B1(n10582), .B2(n9043), .ZN(
        n8972) );
  NAND2_X1 U11534 ( .A1(n10875), .A2(n10736), .ZN(n8970) );
  INV_X1 U11535 ( .A(n14923), .ZN(n10653) );
  AOI22_X1 U11536 ( .A1(n10653), .A2(n9080), .B1(n9091), .B2(n12862), .ZN(
        n8971) );
  INV_X1 U11537 ( .A(n10875), .ZN(n14934) );
  AOI21_X1 U11538 ( .B1(n10736), .B2(n9091), .A(n14934), .ZN(n8974) );
  AOI21_X1 U11539 ( .B1(n12861), .B2(n9080), .A(n10875), .ZN(n8973) );
  AOI22_X1 U11540 ( .A1(n14942), .A2(n9080), .B1(n9091), .B2(n12860), .ZN(
        n8976) );
  INV_X1 U11541 ( .A(n12860), .ZN(n11112) );
  OAI22_X1 U11542 ( .A1(n6956), .A2(n9092), .B1(n11112), .B2(n9043), .ZN(n8975) );
  NAND2_X1 U11543 ( .A1(n8977), .A2(n8976), .ZN(n8978) );
  NAND2_X1 U11544 ( .A1(n8979), .A2(n8978), .ZN(n8980) );
  OAI22_X1 U11545 ( .A1(n14527), .A2(n9092), .B1(n11122), .B2(n9043), .ZN(
        n8981) );
  NAND2_X1 U11546 ( .A1(n8980), .A2(n8981), .ZN(n8985) );
  OAI22_X1 U11547 ( .A1(n14527), .A2(n9043), .B1(n11122), .B2(n9080), .ZN(
        n8984) );
  INV_X1 U11548 ( .A(n8980), .ZN(n8983) );
  INV_X1 U11549 ( .A(n8981), .ZN(n8982) );
  AOI22_X1 U11550 ( .A1(n11152), .A2(n9080), .B1(n9091), .B2(n12858), .ZN(
        n8988) );
  INV_X1 U11551 ( .A(n8988), .ZN(n8987) );
  AOI22_X1 U11552 ( .A1(n11152), .A2(n9091), .B1(n12858), .B2(n9080), .ZN(
        n8986) );
  INV_X1 U11553 ( .A(n12857), .ZN(n11273) );
  OAI22_X1 U11554 ( .A1(n14520), .A2(n9092), .B1(n11273), .B2(n9043), .ZN(
        n8994) );
  OAI22_X1 U11555 ( .A1(n14520), .A2(n9043), .B1(n11273), .B2(n9080), .ZN(
        n8991) );
  NAND2_X1 U11556 ( .A1(n8992), .A2(n8991), .ZN(n8998) );
  INV_X1 U11557 ( .A(n8993), .ZN(n8996) );
  INV_X1 U11558 ( .A(n8994), .ZN(n8995) );
  NAND2_X1 U11559 ( .A1(n8996), .A2(n8995), .ZN(n8997) );
  NAND2_X1 U11560 ( .A1(n8998), .A2(n8997), .ZN(n9002) );
  OAI22_X1 U11561 ( .A1(n11375), .A2(n9043), .B1(n11364), .B2(n9080), .ZN(
        n9001) );
  OAI22_X1 U11562 ( .A1(n11375), .A2(n9092), .B1(n11364), .B2(n9043), .ZN(
        n8999) );
  INV_X1 U11563 ( .A(n8999), .ZN(n9000) );
  AOI21_X1 U11564 ( .B1(n9002), .B2(n9001), .A(n9000), .ZN(n9003) );
  AOI22_X1 U11565 ( .A1(n13258), .A2(n9091), .B1(n12956), .B2(n9080), .ZN(
        n9006) );
  INV_X1 U11566 ( .A(n9006), .ZN(n9005) );
  AOI22_X1 U11567 ( .A1(n13258), .A2(n9080), .B1(n9091), .B2(n12956), .ZN(
        n9004) );
  OAI22_X1 U11568 ( .A1(n13174), .A2(n9043), .B1(n12958), .B2(n9080), .ZN(
        n9010) );
  NAND2_X1 U11569 ( .A1(n9009), .A2(n9010), .ZN(n9008) );
  OAI22_X1 U11570 ( .A1(n13174), .A2(n9080), .B1(n12958), .B2(n9043), .ZN(
        n9007) );
  NAND2_X1 U11571 ( .A1(n9008), .A2(n9007), .ZN(n9014) );
  INV_X1 U11572 ( .A(n9009), .ZN(n9012) );
  INV_X1 U11573 ( .A(n9010), .ZN(n9011) );
  NAND2_X1 U11574 ( .A1(n9012), .A2(n9011), .ZN(n9013) );
  OAI22_X1 U11575 ( .A1(n13155), .A2(n9092), .B1(n12961), .B2(n9043), .ZN(
        n9016) );
  OAI22_X1 U11576 ( .A1(n13155), .A2(n9043), .B1(n12961), .B2(n9080), .ZN(
        n9018) );
  INV_X1 U11577 ( .A(n9016), .ZN(n9017) );
  OAI22_X1 U11578 ( .A1(n13244), .A2(n9043), .B1(n12964), .B2(n9080), .ZN(
        n9020) );
  INV_X1 U11579 ( .A(n9020), .ZN(n9019) );
  OAI22_X1 U11580 ( .A1(n13244), .A2(n9080), .B1(n12964), .B2(n9043), .ZN(
        n9021) );
  OAI22_X1 U11581 ( .A1(n13122), .A2(n9080), .B1(n12967), .B2(n9043), .ZN(
        n9024) );
  INV_X1 U11582 ( .A(n9024), .ZN(n9023) );
  OAI22_X1 U11583 ( .A1(n13122), .A2(n9043), .B1(n12967), .B2(n6433), .ZN(
        n9022) );
  NAND2_X1 U11584 ( .A1(n9025), .A2(n9023), .ZN(n9026) );
  NAND2_X1 U11585 ( .A1(n9027), .A2(n9026), .ZN(n9028) );
  AOI22_X1 U11586 ( .A1(n13230), .A2(n9080), .B1(n9091), .B2(n12969), .ZN(
        n9029) );
  AOI22_X1 U11587 ( .A1(n13226), .A2(n9091), .B1(n12972), .B2(n9080), .ZN(
        n9032) );
  INV_X1 U11588 ( .A(n13226), .ZN(n12826) );
  INV_X1 U11589 ( .A(n12972), .ZN(n12921) );
  OAI22_X1 U11590 ( .A1(n12826), .A2(n9043), .B1(n12921), .B2(n9080), .ZN(
        n9031) );
  OAI22_X1 U11591 ( .A1(n13220), .A2(n9043), .B1(n12974), .B2(n6433), .ZN(
        n9034) );
  INV_X1 U11592 ( .A(n12974), .ZN(n12854) );
  AOI22_X1 U11593 ( .A1(n13081), .A2(n9091), .B1(n12854), .B2(n9080), .ZN(
        n9033) );
  OAI22_X1 U11594 ( .A1(n13054), .A2(n9092), .B1(n12977), .B2(n9043), .ZN(
        n9038) );
  OAI22_X1 U11595 ( .A1(n13054), .A2(n9043), .B1(n12977), .B2(n9092), .ZN(
        n9037) );
  INV_X1 U11596 ( .A(n9038), .ZN(n9039) );
  OAI22_X1 U11597 ( .A1(n13039), .A2(n9043), .B1(n12980), .B2(n6433), .ZN(
        n9041) );
  AOI22_X1 U11598 ( .A1(n13208), .A2(n9091), .B1(n12853), .B2(n9080), .ZN(
        n9040) );
  NOR2_X1 U11599 ( .A1(n9042), .A2(n9041), .ZN(n9048) );
  AOI22_X1 U11600 ( .A1(n13202), .A2(n9091), .B1(n12941), .B2(n9080), .ZN(
        n9097) );
  OAI22_X1 U11601 ( .A1(n13028), .A2(n9043), .B1(n12983), .B2(n6433), .ZN(
        n9096) );
  AND2_X1 U11602 ( .A1(n12985), .A2(n9091), .ZN(n9044) );
  AOI21_X1 U11603 ( .B1(n13196), .B2(n9080), .A(n9044), .ZN(n9094) );
  NAND2_X1 U11604 ( .A1(n13196), .A2(n9091), .ZN(n9046) );
  NAND2_X1 U11605 ( .A1(n12985), .A2(n9080), .ZN(n9045) );
  NAND2_X1 U11606 ( .A1(n9046), .A2(n9045), .ZN(n9093) );
  NOR2_X1 U11607 ( .A1(n9094), .A2(n9093), .ZN(n9095) );
  AOI21_X1 U11608 ( .B1(n9097), .B2(n9096), .A(n9095), .ZN(n9047) );
  OAI21_X1 U11609 ( .B1(n9049), .B2(n9048), .A(n9047), .ZN(n9106) );
  INV_X1 U11610 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9053) );
  NAND2_X1 U11611 ( .A1(n7550), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9052) );
  NAND2_X1 U11612 ( .A1(n9050), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9051) );
  OAI211_X1 U11613 ( .C1(n9078), .C2(n9053), .A(n9052), .B(n9051), .ZN(n12914)
         );
  INV_X1 U11614 ( .A(n9056), .ZN(n9057) );
  MUX2_X1 U11615 ( .A(n13463), .B(n13285), .S(n11553), .Z(n9058) );
  XNOR2_X1 U11616 ( .A(n9058), .B(SI_29_), .ZN(n9083) );
  NAND2_X1 U11617 ( .A1(n9084), .A2(n9083), .ZN(n9060) );
  NAND2_X1 U11618 ( .A1(n9058), .A2(n12734), .ZN(n9059) );
  MUX2_X1 U11619 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11553), .Z(n9061) );
  XNOR2_X1 U11620 ( .A(n9061), .B(SI_30_), .ZN(n9069) );
  NAND2_X1 U11621 ( .A1(n9061), .A2(SI_30_), .ZN(n9062) );
  MUX2_X1 U11622 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11553), .Z(n9063) );
  INV_X1 U11623 ( .A(SI_31_), .ZN(n12727) );
  XNOR2_X1 U11624 ( .A(n9063), .B(n12727), .ZN(n9064) );
  INV_X1 U11625 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n9065) );
  AOI22_X1 U11626 ( .A1(n9107), .A2(n9080), .B1(n9091), .B2(n12914), .ZN(n9067) );
  OAI21_X1 U11627 ( .B1(n12914), .B2(n9107), .A(n9067), .ZN(n9090) );
  INV_X1 U11628 ( .A(n9069), .ZN(n9070) );
  NAND2_X1 U11629 ( .A1(n13445), .A2(n9085), .ZN(n9072) );
  INV_X1 U11630 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11648) );
  OR2_X1 U11631 ( .A1(n7943), .A2(n11648), .ZN(n9071) );
  INV_X1 U11632 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n9077) );
  NAND2_X1 U11633 ( .A1(n9073), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9076) );
  NAND2_X1 U11634 ( .A1(n9074), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9075) );
  OAI211_X1 U11635 ( .C1(n9078), .C2(n9077), .A(n9076), .B(n9075), .ZN(n12948)
         );
  NAND2_X1 U11636 ( .A1(n9080), .A2(n12914), .ZN(n9122) );
  NAND2_X1 U11637 ( .A1(n9129), .A2(n12903), .ZN(n9938) );
  OR2_X1 U11638 ( .A1(n9938), .A2(n9160), .ZN(n9161) );
  NAND4_X1 U11639 ( .A1(n9122), .A2(n6464), .A3(n9171), .A4(n9161), .ZN(n9079)
         );
  AOI22_X1 U11640 ( .A1(n9151), .A2(n9091), .B1(n12948), .B2(n9079), .ZN(n9116) );
  NAND2_X1 U11641 ( .A1(n9151), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U11642 ( .A1(n9091), .A2(n12948), .ZN(n9081) );
  NAND2_X1 U11643 ( .A1(n9082), .A2(n9081), .ZN(n9117) );
  NAND2_X1 U11644 ( .A1(n13462), .A2(n9085), .ZN(n9087) );
  OR2_X1 U11645 ( .A1(n7943), .A2(n13285), .ZN(n9086) );
  INV_X1 U11646 ( .A(n9088), .ZN(n12852) );
  AOI22_X1 U11647 ( .A1(n13185), .A2(n9091), .B1(n12852), .B2(n9080), .ZN(
        n9108) );
  OAI22_X1 U11648 ( .A1(n12955), .A2(n9043), .B1(n9088), .B2(n9092), .ZN(n9109) );
  OAI22_X1 U11649 ( .A1(n9116), .A2(n9117), .B1(n9108), .B2(n9109), .ZN(n9089)
         );
  NAND2_X1 U11650 ( .A1(n9090), .A2(n9089), .ZN(n9114) );
  AOI22_X1 U11651 ( .A1(n13190), .A2(n9080), .B1(n9091), .B2(n12946), .ZN(
        n9111) );
  OAI22_X1 U11652 ( .A1(n12909), .A2(n9092), .B1(n12943), .B2(n9043), .ZN(
        n9110) );
  INV_X1 U11653 ( .A(n9093), .ZN(n9103) );
  INV_X1 U11654 ( .A(n9094), .ZN(n9102) );
  INV_X1 U11655 ( .A(n9095), .ZN(n9100) );
  INV_X1 U11656 ( .A(n9096), .ZN(n9099) );
  INV_X1 U11657 ( .A(n9097), .ZN(n9098) );
  NAND3_X1 U11658 ( .A1(n9100), .A2(n9099), .A3(n9098), .ZN(n9101) );
  OAI21_X1 U11659 ( .B1(n9103), .B2(n9102), .A(n9101), .ZN(n9104) );
  AOI21_X1 U11660 ( .B1(n9111), .B2(n9110), .A(n9104), .ZN(n9105) );
  NAND2_X1 U11661 ( .A1(n9106), .A2(n7449), .ZN(n9121) );
  XNOR2_X1 U11662 ( .A(n13180), .B(n12914), .ZN(n9130) );
  INV_X1 U11663 ( .A(n9108), .ZN(n9113) );
  INV_X1 U11664 ( .A(n9109), .ZN(n9112) );
  OAI22_X1 U11665 ( .A1(n9113), .A2(n9112), .B1(n9111), .B2(n9110), .ZN(n9115)
         );
  OAI21_X1 U11666 ( .B1(n9130), .B2(n9115), .A(n9114), .ZN(n9119) );
  NAND2_X1 U11667 ( .A1(n9121), .A2(n9120), .ZN(n9126) );
  NAND2_X1 U11668 ( .A1(n9122), .A2(n6433), .ZN(n9124) );
  NAND2_X1 U11669 ( .A1(n9043), .A2(n12914), .ZN(n9123) );
  MUX2_X1 U11670 ( .A(n9124), .B(n9123), .S(n13180), .Z(n9125) );
  INV_X1 U11671 ( .A(n9162), .ZN(n9157) );
  NAND2_X1 U11672 ( .A1(n6464), .A2(n13001), .ZN(n9127) );
  OAI211_X1 U11673 ( .C1(n9129), .C2(n9128), .A(n9171), .B(n9127), .ZN(n9156)
         );
  INV_X1 U11674 ( .A(n9130), .ZN(n9148) );
  INV_X1 U11675 ( .A(n12985), .ZN(n12942) );
  XNOR2_X1 U11676 ( .A(n13196), .B(n12942), .ZN(n13016) );
  NAND2_X1 U11677 ( .A1(n13190), .A2(n12946), .ZN(n12987) );
  XNOR2_X1 U11678 ( .A(n13214), .B(n12977), .ZN(n13053) );
  XNOR2_X1 U11679 ( .A(n13226), .B(n12921), .ZN(n13092) );
  NAND2_X1 U11680 ( .A1(n13081), .A2(n12974), .ZN(n12938) );
  OR2_X1 U11681 ( .A1(n13081), .A2(n12974), .ZN(n9132) );
  NAND2_X1 U11682 ( .A1(n12938), .A2(n9132), .ZN(n13066) );
  NAND2_X1 U11683 ( .A1(n13237), .A2(n12967), .ZN(n12933) );
  OR2_X1 U11684 ( .A1(n13237), .A2(n12967), .ZN(n9133) );
  XNOR2_X1 U11685 ( .A(n13248), .B(n12961), .ZN(n13157) );
  INV_X1 U11686 ( .A(n12956), .ZN(n12924) );
  XNOR2_X1 U11687 ( .A(n13258), .B(n12924), .ZN(n11362) );
  NAND2_X1 U11688 ( .A1(n13255), .A2(n12958), .ZN(n12927) );
  OR2_X1 U11689 ( .A1(n13255), .A2(n12958), .ZN(n9134) );
  NAND2_X1 U11690 ( .A1(n12927), .A2(n9134), .ZN(n13165) );
  XNOR2_X1 U11691 ( .A(n11287), .B(n12856), .ZN(n11358) );
  INV_X1 U11692 ( .A(n12864), .ZN(n9773) );
  OR2_X1 U11693 ( .A1(n10443), .A2(n9773), .ZN(n10249) );
  NAND2_X1 U11694 ( .A1(n10443), .A2(n9773), .ZN(n9135) );
  NAND2_X1 U11695 ( .A1(n10249), .A2(n9135), .ZN(n10448) );
  XNOR2_X1 U11696 ( .A(n14916), .B(n10475), .ZN(n10246) );
  XNOR2_X1 U11697 ( .A(n14901), .B(n10242), .ZN(n10240) );
  NAND2_X1 U11698 ( .A1(n9927), .A2(n9136), .ZN(n14858) );
  NOR4_X1 U11699 ( .A1(n9918), .A2(n7504), .A3(n10539), .A4(n14858), .ZN(n9137) );
  XNOR2_X1 U11700 ( .A(n10177), .B(n12867), .ZN(n10170) );
  XNOR2_X1 U11701 ( .A(n9932), .B(n12868), .ZN(n14810) );
  NAND4_X1 U11702 ( .A1(n10152), .A2(n9137), .A3(n10170), .A4(n14810), .ZN(
        n9138) );
  NOR4_X1 U11703 ( .A1(n10448), .A2(n10246), .A3(n10240), .A4(n9138), .ZN(
        n9139) );
  XNOR2_X1 U11704 ( .A(n14942), .B(n12860), .ZN(n10878) );
  XNOR2_X1 U11705 ( .A(n10653), .B(n12862), .ZN(n10465) );
  NAND4_X1 U11706 ( .A1(n10578), .A2(n9139), .A3(n10878), .A4(n10465), .ZN(
        n9141) );
  INV_X1 U11707 ( .A(n12858), .ZN(n11116) );
  OR2_X1 U11708 ( .A1(n11152), .A2(n11116), .ZN(n11115) );
  NAND2_X1 U11709 ( .A1(n11152), .A2(n11116), .ZN(n9140) );
  NAND2_X1 U11710 ( .A1(n11115), .A2(n9140), .ZN(n11138) );
  NOR2_X1 U11711 ( .A1(n9141), .A2(n11138), .ZN(n9142) );
  XNOR2_X1 U11712 ( .A(n14498), .B(n12857), .ZN(n11125) );
  INV_X1 U11713 ( .A(n14527), .ZN(n11019) );
  XNOR2_X1 U11714 ( .A(n11019), .B(n12859), .ZN(n14508) );
  NAND4_X1 U11715 ( .A1(n11358), .A2(n9142), .A3(n11125), .A4(n14508), .ZN(
        n9143) );
  NOR4_X1 U11716 ( .A1(n13157), .A2(n11362), .A3(n13165), .A4(n9143), .ZN(
        n9144) );
  XNOR2_X1 U11717 ( .A(n13230), .B(n12969), .ZN(n13109) );
  XNOR2_X1 U11718 ( .A(n6949), .B(n12930), .ZN(n13135) );
  NAND4_X1 U11719 ( .A1(n13125), .A2(n9144), .A3(n13109), .A4(n13135), .ZN(
        n9145) );
  NOR4_X1 U11720 ( .A1(n13053), .A2(n13092), .A3(n13066), .A4(n9145), .ZN(
        n9146) );
  XNOR2_X1 U11721 ( .A(n13202), .B(n12941), .ZN(n13030) );
  NAND4_X1 U11722 ( .A1(n12986), .A2(n9146), .A3(n13030), .A4(n13037), .ZN(
        n9147) );
  XNOR2_X1 U11723 ( .A(n13185), .B(n12852), .ZN(n12988) );
  INV_X1 U11724 ( .A(n12948), .ZN(n9152) );
  NAND3_X1 U11725 ( .A1(n9151), .A2(n9152), .A3(n13001), .ZN(n9150) );
  NOR2_X1 U11726 ( .A1(n13001), .A2(n9160), .ZN(n11150) );
  INV_X1 U11727 ( .A(n11150), .ZN(n9149) );
  NAND3_X1 U11728 ( .A1(n9150), .A2(n11050), .A3(n9149), .ZN(n9154) );
  INV_X1 U11729 ( .A(n9158), .ZN(n9159) );
  NOR3_X1 U11730 ( .A1(n9159), .A2(n6464), .A3(n13001), .ZN(n9164) );
  NAND2_X1 U11731 ( .A1(n6464), .A2(n9160), .ZN(n9937) );
  OAI21_X1 U11732 ( .B1(n13001), .B2(n9937), .A(n9161), .ZN(n9163) );
  OAI21_X1 U11733 ( .B1(n9164), .B2(n9163), .A(n9162), .ZN(n9165) );
  NAND2_X1 U11734 ( .A1(n9166), .A2(n9165), .ZN(n9168) );
  OR2_X1 U11735 ( .A1(n9377), .A2(P2_U3088), .ZN(n11295) );
  NAND2_X1 U11736 ( .A1(n9168), .A2(n9167), .ZN(n9175) );
  NAND2_X1 U11737 ( .A1(n9170), .A2(n9169), .ZN(n13295) );
  NOR4_X1 U11738 ( .A1(n14851), .A2(n12843), .A3(n9171), .A4(n13295), .ZN(
        n9172) );
  AOI211_X1 U11739 ( .C1(n9167), .C2(n6700), .A(n12911), .B(n9172), .ZN(n9173)
         );
  INV_X1 U11740 ( .A(n9173), .ZN(n9174) );
  NAND2_X1 U11741 ( .A1(n9175), .A2(n9174), .ZN(P2_U3328) );
  INV_X1 U11742 ( .A(n9176), .ZN(n9177) );
  NAND2_X1 U11743 ( .A1(n9177), .A2(n9377), .ZN(n9382) );
  NOR2_X1 U11744 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), 
        .ZN(n9180) );
  NAND4_X1 U11745 ( .A1(n9183), .A2(n9182), .A3(n9181), .A4(n9223), .ZN(n9273)
         );
  NAND2_X1 U11746 ( .A1(n9276), .A2(n9185), .ZN(n9186) );
  OAI21_X1 U11747 ( .B1(n9200), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9189) );
  MUX2_X1 U11748 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9189), .S(
        P1_IR_REG_24__SCAN_IN), .Z(n9196) );
  NAND3_X1 U11749 ( .A1(n12257), .A2(n9191), .A3(n9190), .ZN(n9192) );
  OAI21_X1 U11750 ( .B1(n9294), .B2(P1_IR_REG_25__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U11751 ( .A1(n9294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9198) );
  NAND2_X1 U11752 ( .A1(n9200), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9201) );
  NAND2_X2 U11753 ( .A1(n11553), .A2(P2_U3088), .ZN(n13301) );
  OAI222_X1 U11754 ( .A1(n13303), .A2(n9204), .B1(n13301), .B2(n9618), .C1(
        n9372), .C2(P2_U3088), .ZN(P2_U3326) );
  AND2_X1 U11755 ( .A1(n11553), .A2(P1_U3086), .ZN(n10039) );
  INV_X2 U11756 ( .A(n10039), .ZN(n14252) );
  INV_X1 U11757 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n9209) );
  NOR2_X1 U11758 ( .A1(n11553), .A2(P1_STATE_REG_SCAN_IN), .ZN(n14238) );
  NOR2_X1 U11759 ( .A1(n9205), .A2(n10377), .ZN(n9206) );
  MUX2_X1 U11760 ( .A(n10377), .B(n9206), .S(P1_IR_REG_2__SCAN_IN), .Z(n9208)
         );
  INV_X1 U11761 ( .A(n9274), .ZN(n9207) );
  INV_X1 U11762 ( .A(n13767), .ZN(n9301) );
  OAI222_X1 U11763 ( .A1(n14252), .A2(n9209), .B1(n10724), .B2(n9674), .C1(
        n9301), .C2(P1_U3086), .ZN(P1_U3353) );
  NAND2_X1 U11764 ( .A1(n9274), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9210) );
  XNOR2_X1 U11765 ( .A(n9210), .B(P1_IR_REG_3__SCAN_IN), .ZN(n9833) );
  INV_X1 U11766 ( .A(n9833), .ZN(n13778) );
  INV_X1 U11767 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n9211) );
  OAI222_X1 U11768 ( .A1(P1_U3086), .A2(n13778), .B1(n10724), .B2(n9832), .C1(
        n9211), .C2(n14252), .ZN(P1_U3352) );
  NAND2_X1 U11769 ( .A1(n11553), .A2(P3_U3151), .ZN(n12744) );
  INV_X2 U11770 ( .A(n14376), .ZN(n12747) );
  INV_X1 U11771 ( .A(n9213), .ZN(n9214) );
  OAI222_X1 U11772 ( .A1(P3_U3151), .A2(n10666), .B1(n12744), .B2(n9215), .C1(
        n12747), .C2(n9214), .ZN(P3_U3287) );
  INV_X1 U11773 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n9217) );
  NAND2_X1 U11774 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n9216) );
  XNOR2_X1 U11775 ( .A(n9217), .B(n9216), .ZN(n13754) );
  OAI222_X1 U11776 ( .A1(P1_U3086), .A2(n13754), .B1(n10724), .B2(n9618), .C1(
        n6935), .C2(n14252), .ZN(P1_U3354) );
  OAI222_X1 U11777 ( .A1(n13303), .A2(n12233), .B1(n13301), .B2(n9832), .C1(
        n9388), .C2(P2_U3088), .ZN(P2_U3324) );
  OAI222_X1 U11778 ( .A1(n13303), .A2(n9218), .B1(n13301), .B2(n9674), .C1(
        n7546), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U11779 ( .A(n12744), .ZN(n14375) );
  AOI22_X1 U11780 ( .A1(n10108), .A2(P3_STATE_REG_SCAN_IN), .B1(SI_4_), .B2(
        n14375), .ZN(n9219) );
  OAI21_X1 U11781 ( .B1(n9220), .B2(n12747), .A(n9219), .ZN(P3_U3291) );
  OR2_X1 U11782 ( .A1(n9274), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n9222) );
  NAND2_X1 U11783 ( .A1(n9222), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9221) );
  MUX2_X1 U11784 ( .A(n9221), .B(P1_IR_REG_31__SCAN_IN), .S(n9223), .Z(n9225)
         );
  INV_X1 U11785 ( .A(n9222), .ZN(n9224) );
  NAND2_X1 U11786 ( .A1(n9224), .A2(n9223), .ZN(n9232) );
  NAND2_X1 U11787 ( .A1(n9225), .A2(n9232), .ZN(n9312) );
  INV_X1 U11788 ( .A(n9836), .ZN(n9226) );
  OAI222_X1 U11789 ( .A1(P1_U3086), .A2(n9312), .B1(n10724), .B2(n9226), .C1(
        n6693), .C2(n14252), .ZN(P1_U3351) );
  INV_X1 U11790 ( .A(n9390), .ZN(n9430) );
  OAI222_X1 U11791 ( .A1(n13303), .A2(n9227), .B1(n13301), .B2(n9226), .C1(
        n9430), .C2(P2_U3088), .ZN(P2_U3323) );
  NAND2_X1 U11792 ( .A1(n9245), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9228) );
  XNOR2_X1 U11793 ( .A(n9228), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10263) );
  INV_X1 U11794 ( .A(n10263), .ZN(n9470) );
  OAI222_X1 U11795 ( .A1(P1_U3086), .A2(n9470), .B1(n10724), .B2(n10262), .C1(
        n9229), .C2(n14252), .ZN(P1_U3349) );
  INV_X1 U11796 ( .A(n9561), .ZN(n9402) );
  OAI222_X1 U11797 ( .A1(n13303), .A2(n9230), .B1(n13301), .B2(n10262), .C1(
        n9402), .C2(P2_U3088), .ZN(P2_U3321) );
  INV_X1 U11798 ( .A(n9391), .ZN(n9445) );
  OAI222_X1 U11799 ( .A1(n13303), .A2(n9231), .B1(n13301), .B2(n10213), .C1(
        n9445), .C2(P2_U3088), .ZN(P2_U3322) );
  NAND2_X1 U11800 ( .A1(n9232), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9233) );
  MUX2_X1 U11801 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9233), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n9234) );
  INV_X1 U11802 ( .A(n10214), .ZN(n9342) );
  OAI222_X1 U11803 ( .A1(n14252), .A2(n6710), .B1(n10724), .B2(n10213), .C1(
        n9342), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U11804 ( .A(n13715), .ZN(n9542) );
  INV_X1 U11805 ( .A(P1_B_REG_SCAN_IN), .ZN(n13864) );
  NAND2_X1 U11806 ( .A1(n11448), .A2(n13864), .ZN(n9236) );
  AND2_X2 U11807 ( .A1(n9542), .A2(n9499), .ZN(n14704) );
  OR2_X1 U11808 ( .A1(n14244), .A2(P1_U3086), .ZN(n9238) );
  OR2_X1 U11809 ( .A1(n9238), .A2(n9288), .ZN(n9240) );
  OAI22_X1 U11810 ( .A1(n14704), .A2(P1_D_REG_0__SCAN_IN), .B1(n11448), .B2(
        n9240), .ZN(n9239) );
  INV_X1 U11811 ( .A(n9239), .ZN(P1_U3445) );
  OAI22_X1 U11812 ( .A1(n14704), .A2(P1_D_REG_1__SCAN_IN), .B1(n14248), .B2(
        n9240), .ZN(n9241) );
  INV_X1 U11813 ( .A(n9241), .ZN(P1_U3446) );
  INV_X1 U11814 ( .A(n9242), .ZN(n9243) );
  OAI222_X1 U11815 ( .A1(n12744), .A2(n9244), .B1(n12747), .B2(n9243), .C1(
        n15001), .C2(P3_U3151), .ZN(P3_U3283) );
  OAI21_X1 U11816 ( .B1(n9245), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9246) );
  XNOR2_X1 U11817 ( .A(n9246), .B(P1_IR_REG_7__SCAN_IN), .ZN(n10268) );
  INV_X1 U11818 ( .A(n10268), .ZN(n9457) );
  OAI222_X1 U11819 ( .A1(n14252), .A2(n9247), .B1(n10724), .B2(n10267), .C1(
        n9457), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U11820 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n9249) );
  INV_X1 U11821 ( .A(n14785), .ZN(n9248) );
  OAI222_X1 U11822 ( .A1(n13303), .A2(n9249), .B1(n13301), .B2(n10267), .C1(
        n9248), .C2(P2_U3088), .ZN(P2_U3320) );
  INV_X1 U11823 ( .A(SI_9_), .ZN(n9251) );
  OAI222_X1 U11824 ( .A1(P3_U3151), .A2(n10763), .B1(n12726), .B2(n9251), .C1(
        n12747), .C2(n9250), .ZN(P3_U3286) );
  INV_X1 U11825 ( .A(n9252), .ZN(n9254) );
  OAI222_X1 U11826 ( .A1(n12747), .A2(n9254), .B1(n12726), .B2(n9253), .C1(
        P3_U3151), .C2(n9974), .ZN(P3_U3294) );
  INV_X1 U11827 ( .A(SI_7_), .ZN(n9256) );
  OAI222_X1 U11828 ( .A1(P3_U3151), .A2(n10388), .B1(n12726), .B2(n9256), .C1(
        n12747), .C2(n9255), .ZN(P3_U3288) );
  INV_X1 U11829 ( .A(SI_10_), .ZN(n9258) );
  OAI222_X1 U11830 ( .A1(P3_U3151), .A2(n12314), .B1(n12726), .B2(n9258), .C1(
        n12747), .C2(n9257), .ZN(P3_U3285) );
  OAI222_X1 U11831 ( .A1(P3_U3151), .A2(n14982), .B1(n12726), .B2(n9260), .C1(
        n12747), .C2(n9259), .ZN(P3_U3284) );
  INV_X1 U11832 ( .A(n9261), .ZN(n9263) );
  OAI222_X1 U11833 ( .A1(P3_U3151), .A2(n10354), .B1(n12747), .B2(n9263), .C1(
        n9262), .C2(n12726), .ZN(P3_U3289) );
  INV_X1 U11834 ( .A(n9264), .ZN(n9265) );
  OAI222_X1 U11835 ( .A1(P3_U3151), .A2(n9994), .B1(n12747), .B2(n9265), .C1(
        n9515), .C2(n12726), .ZN(P3_U3295) );
  INV_X1 U11836 ( .A(SI_5_), .ZN(n9266) );
  OAI222_X1 U11837 ( .A1(n10003), .A2(P3_U3151), .B1(n12747), .B2(n9267), .C1(
        n9266), .C2(n12726), .ZN(P3_U3290) );
  INV_X1 U11838 ( .A(SI_3_), .ZN(n9268) );
  OAI222_X1 U11839 ( .A1(n9999), .A2(P3_U3151), .B1(n12747), .B2(n9269), .C1(
        n9268), .C2(n12726), .ZN(P3_U3292) );
  INV_X1 U11840 ( .A(n6431), .ZN(n9976) );
  INV_X1 U11841 ( .A(SI_2_), .ZN(n9270) );
  OAI222_X1 U11842 ( .A1(n9976), .A2(P3_U3151), .B1(n12747), .B2(n9271), .C1(
        n9270), .C2(n12726), .ZN(P3_U3293) );
  INV_X1 U11843 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n9272) );
  INV_X1 U11844 ( .A(n9590), .ZN(n9568) );
  OAI222_X1 U11845 ( .A1(n13303), .A2(n9272), .B1(n13301), .B2(n10487), .C1(
        n9568), .C2(P2_U3088), .ZN(P2_U3319) );
  NOR2_X1 U11846 ( .A1(n9274), .A2(n9273), .ZN(n9277) );
  NOR2_X1 U11847 ( .A1(n9277), .A2(n10377), .ZN(n9275) );
  MUX2_X1 U11848 ( .A(n10377), .B(n9275), .S(P1_IR_REG_8__SCAN_IN), .Z(n9279)
         );
  NAND2_X1 U11849 ( .A1(n9277), .A2(n9276), .ZN(n10035) );
  INV_X1 U11850 ( .A(n10035), .ZN(n9278) );
  OAI222_X1 U11851 ( .A1(n14252), .A2(n9280), .B1(n10724), .B2(n10487), .C1(
        n9406), .C2(P1_U3086), .ZN(P1_U3347) );
  NAND2_X1 U11852 ( .A1(n9325), .A2(P3_D_REG_0__SCAN_IN), .ZN(n9281) );
  OAI21_X1 U11853 ( .B1(n9282), .B2(n9325), .A(n9281), .ZN(P3_U3376) );
  AND2_X1 U11854 ( .A1(n9288), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13726) );
  INV_X1 U11855 ( .A(n13726), .ZN(n13717) );
  AND2_X1 U11856 ( .A1(n13715), .A2(n13717), .ZN(n9318) );
  XNOR2_X1 U11857 ( .A(n9283), .B(n9284), .ZN(n9500) );
  INV_X1 U11858 ( .A(n9500), .ZN(n9508) );
  OR2_X1 U11859 ( .A1(n13457), .A2(n9288), .ZN(n9298) );
  NAND2_X1 U11860 ( .A1(n9357), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9290) );
  AND3_X1 U11861 ( .A1(n9292), .A2(n9291), .A3(P1_IR_REG_27__SCAN_IN), .ZN(
        n9297) );
  XNOR2_X1 U11862 ( .A(n9293), .B(P1_IR_REG_31__SCAN_IN), .ZN(n9296) );
  NAND3_X1 U11863 ( .A1(n9294), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n9295) );
  OR2_X1 U11864 ( .A1(n9318), .A2(n9320), .ZN(n14630) );
  NOR2_X1 U11865 ( .A1(n14630), .A2(n9525), .ZN(n14637) );
  INV_X1 U11866 ( .A(n14619), .ZN(n9300) );
  NOR2_X2 U11867 ( .A1(n14630), .A2(n9300), .ZN(n14640) );
  INV_X1 U11868 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9302) );
  INV_X1 U11869 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9633) );
  MUX2_X1 U11870 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9633), .S(n13767), .Z(
        n13773) );
  INV_X1 U11871 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9520) );
  XNOR2_X1 U11872 ( .A(n13754), .B(P1_REG1_REG_1__SCAN_IN), .ZN(n13761) );
  NAND3_X1 U11873 ( .A1(n13761), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n13759) );
  OAI21_X1 U11874 ( .B1(n13754), .B2(n9520), .A(n13759), .ZN(n13772) );
  NAND2_X1 U11875 ( .A1(n13773), .A2(n13772), .ZN(n13771) );
  OAI21_X1 U11876 ( .B1(n9301), .B2(n9633), .A(n13771), .ZN(n13782) );
  XOR2_X1 U11877 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9833), .Z(n13783) );
  NAND2_X1 U11878 ( .A1(n13782), .A2(n13783), .ZN(n13781) );
  OAI21_X1 U11879 ( .B1(n9302), .B2(n13778), .A(n13781), .ZN(n9661) );
  XNOR2_X1 U11880 ( .A(n9312), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9662) );
  INV_X1 U11881 ( .A(n9312), .ZN(n9837) );
  INV_X1 U11882 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9857) );
  MUX2_X1 U11883 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n9857), .S(n10214), .Z(n9303) );
  NAND2_X1 U11884 ( .A1(n9304), .A2(n9303), .ZN(n9336) );
  OAI21_X1 U11885 ( .B1(n9304), .B2(n9303), .A(n9336), .ZN(n9317) );
  INV_X1 U11886 ( .A(n14630), .ZN(n9306) );
  NOR2_X1 U11887 ( .A1(n6468), .A2(n14619), .ZN(n9305) );
  NAND2_X1 U11888 ( .A1(n9306), .A2(n9305), .ZN(n13851) );
  INV_X1 U11889 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9307) );
  MUX2_X1 U11890 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n9307), .S(n13754), .Z(n9309) );
  INV_X1 U11891 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n9308) );
  INV_X1 U11892 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n14621) );
  NOR3_X1 U11893 ( .A1(n9309), .A2(n9308), .A3(n14621), .ZN(n13755) );
  AOI21_X1 U11894 ( .B1(n7362), .B2(P1_REG2_REG_1__SCAN_IN), .A(n13755), .ZN(
        n13769) );
  INV_X1 U11895 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n9310) );
  MUX2_X1 U11896 ( .A(n9310), .B(P1_REG2_REG_2__SCAN_IN), .S(n13767), .Z(
        n13768) );
  OR2_X1 U11897 ( .A1(n13769), .A2(n13768), .ZN(n13787) );
  NAND2_X1 U11898 ( .A1(n13767), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13786) );
  INV_X1 U11899 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9311) );
  MUX2_X1 U11900 ( .A(n9311), .B(P1_REG2_REG_3__SCAN_IN), .S(n9833), .Z(n13785) );
  AOI21_X1 U11901 ( .B1(n13787), .B2(n13786), .A(n13785), .ZN(n13784) );
  NOR2_X1 U11902 ( .A1(n13778), .A2(n9311), .ZN(n9668) );
  INV_X1 U11903 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9840) );
  MUX2_X1 U11904 ( .A(n9840), .B(P1_REG2_REG_4__SCAN_IN), .S(n9312), .Z(n9667)
         );
  OAI21_X1 U11905 ( .B1(n13784), .B2(n9668), .A(n9667), .ZN(n9666) );
  NAND2_X1 U11906 ( .A1(n9837), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n9314) );
  INV_X1 U11907 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n9341) );
  MUX2_X1 U11908 ( .A(n9341), .B(P1_REG2_REG_5__SCAN_IN), .S(n10214), .Z(n9313) );
  AOI21_X1 U11909 ( .B1(n9666), .B2(n9314), .A(n9313), .ZN(n9466) );
  AND3_X1 U11910 ( .A1(n9666), .A2(n9314), .A3(n9313), .ZN(n9315) );
  NOR3_X1 U11911 ( .A1(n13851), .A2(n9466), .A3(n9315), .ZN(n9316) );
  AOI21_X1 U11912 ( .B1(n14640), .B2(n9317), .A(n9316), .ZN(n9323) );
  INV_X1 U11913 ( .A(n9318), .ZN(n9319) );
  AND2_X1 U11914 ( .A1(n9320), .A2(n9319), .ZN(n14627) );
  NAND2_X1 U11915 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10337) );
  INV_X1 U11916 ( .A(n10337), .ZN(n9321) );
  AOI21_X1 U11917 ( .B1(n14627), .B2(P1_ADDR_REG_5__SCAN_IN), .A(n9321), .ZN(
        n9322) );
  OAI211_X1 U11918 ( .C1(n9342), .C2(n13807), .A(n9323), .B(n9322), .ZN(
        P1_U3248) );
  NAND2_X1 U11919 ( .A1(n9325), .A2(P3_D_REG_1__SCAN_IN), .ZN(n9324) );
  OAI21_X1 U11920 ( .B1(n10183), .B2(n9325), .A(n9324), .ZN(P3_U3377) );
  NAND2_X1 U11921 ( .A1(n10035), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9326) );
  MUX2_X1 U11922 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9326), .S(
        P1_IR_REG_9__SCAN_IN), .Z(n9327) );
  INV_X1 U11923 ( .A(n10493), .ZN(n9605) );
  OAI222_X1 U11924 ( .A1(n14252), .A2(n12253), .B1(n10724), .B2(n10492), .C1(
        n9605), .C2(P1_U3086), .ZN(P1_U3346) );
  INV_X1 U11925 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n9328) );
  OAI222_X1 U11926 ( .A1(n13303), .A2(n9328), .B1(n13301), .B2(n10492), .C1(
        n9591), .C2(P2_U3088), .ZN(P2_U3318) );
  AND2_X1 U11927 ( .A1(n9334), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U11928 ( .A1(n9334), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U11929 ( .A1(n9334), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U11930 ( .A1(n9334), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U11931 ( .A1(n9334), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U11932 ( .A1(n9334), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U11933 ( .A1(n9334), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U11934 ( .A1(n9334), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U11935 ( .A1(n9334), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U11936 ( .A1(n9334), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U11937 ( .A1(n9334), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U11938 ( .A1(n9334), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U11939 ( .A1(n9334), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U11940 ( .A1(n9334), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U11941 ( .A1(n9334), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U11942 ( .A1(n9334), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U11943 ( .A1(n9334), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U11944 ( .A1(n9334), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U11945 ( .A1(n9334), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U11946 ( .A1(n9334), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U11947 ( .A1(n9334), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U11948 ( .A1(n9334), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U11949 ( .A1(n9334), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U11950 ( .A1(n9334), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  AND2_X1 U11951 ( .A1(n9334), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U11952 ( .A1(n9334), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  INV_X1 U11953 ( .A(P1_U4016), .ZN(n13751) );
  INV_X1 U11954 ( .A(n13751), .ZN(n13750) );
  NOR2_X1 U11955 ( .A1(n14627), .A2(n13750), .ZN(P1_U3085) );
  INV_X1 U11956 ( .A(n9331), .ZN(n9332) );
  OAI222_X1 U11957 ( .A1(n12744), .A2(n9333), .B1(n12747), .B2(n9332), .C1(
        P3_U3151), .C2(n12339), .ZN(P3_U3282) );
  INV_X1 U11958 ( .A(n9334), .ZN(n9335) );
  INV_X1 U11959 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n12209) );
  NOR2_X1 U11960 ( .A1(n9335), .A2(n12209), .ZN(P3_U3235) );
  INV_X1 U11961 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n12227) );
  NOR2_X1 U11962 ( .A1(n9335), .A2(n12227), .ZN(P3_U3249) );
  INV_X1 U11963 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n12269) );
  NOR2_X1 U11964 ( .A1(n9335), .A2(n12269), .ZN(P3_U3243) );
  INV_X1 U11965 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n12239) );
  NOR2_X1 U11966 ( .A1(n9335), .A2(n12239), .ZN(P3_U3237) );
  OAI21_X1 U11967 ( .B1(n10214), .B2(P1_REG1_REG_5__SCAN_IN), .A(n9336), .ZN(
        n9461) );
  INV_X1 U11968 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10226) );
  MUX2_X1 U11969 ( .A(n10226), .B(P1_REG1_REG_6__SCAN_IN), .S(n10263), .Z(
        n9462) );
  NOR2_X1 U11970 ( .A1(n9461), .A2(n9462), .ZN(n9460) );
  INV_X1 U11971 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n10273) );
  MUX2_X1 U11972 ( .A(n10273), .B(P1_REG1_REG_7__SCAN_IN), .S(n10268), .Z(
        n9448) );
  NOR2_X1 U11973 ( .A1(n9449), .A2(n9448), .ZN(n9447) );
  AOI21_X1 U11974 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(n10268), .A(n9447), .ZN(
        n9338) );
  INV_X1 U11975 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10289) );
  MUX2_X1 U11976 ( .A(n10289), .B(P1_REG1_REG_8__SCAN_IN), .S(n9406), .Z(n9337) );
  NAND2_X1 U11977 ( .A1(n9338), .A2(n9337), .ZN(n9411) );
  OAI21_X1 U11978 ( .B1(n9338), .B2(n9337), .A(n9411), .ZN(n9350) );
  AND2_X1 U11979 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9339) );
  AOI21_X1 U11980 ( .B1(n14627), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n9339), .ZN(
        n9340) );
  OAI21_X1 U11981 ( .B1(n13807), .B2(n9406), .A(n9340), .ZN(n9349) );
  NOR2_X1 U11982 ( .A1(n9342), .A2(n9341), .ZN(n9465) );
  INV_X1 U11983 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10222) );
  MUX2_X1 U11984 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10222), .S(n10263), .Z(
        n9464) );
  OAI21_X1 U11985 ( .B1(n9466), .B2(n9465), .A(n9464), .ZN(n9463) );
  NAND2_X1 U11986 ( .A1(n10263), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n9452) );
  INV_X1 U11987 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n9343) );
  MUX2_X1 U11988 ( .A(n9343), .B(P1_REG2_REG_7__SCAN_IN), .S(n10268), .Z(n9451) );
  AOI21_X1 U11989 ( .B1(n9463), .B2(n9452), .A(n9451), .ZN(n9450) );
  NOR2_X1 U11990 ( .A1(n9457), .A2(n9343), .ZN(n9345) );
  INV_X1 U11991 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10285) );
  MUX2_X1 U11992 ( .A(n10285), .B(P1_REG2_REG_8__SCAN_IN), .S(n9406), .Z(n9344) );
  OAI21_X1 U11993 ( .B1(n9450), .B2(n9345), .A(n9344), .ZN(n9409) );
  INV_X1 U11994 ( .A(n9409), .ZN(n9347) );
  NOR3_X1 U11995 ( .A1(n9450), .A2(n9345), .A3(n9344), .ZN(n9346) );
  NOR3_X1 U11996 ( .A1(n9347), .A2(n9346), .A3(n13851), .ZN(n9348) );
  AOI211_X1 U11997 ( .C1(n14640), .C2(n9350), .A(n9349), .B(n9348), .ZN(n9351)
         );
  INV_X1 U11998 ( .A(n9351), .ZN(P1_U3251) );
  INV_X1 U11999 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n9352) );
  INV_X1 U12000 ( .A(n10137), .ZN(n9805) );
  OAI222_X1 U12001 ( .A1(n13303), .A2(n9352), .B1(n13301), .B2(n10821), .C1(
        n9805), .C2(P2_U3088), .ZN(P2_U3317) );
  NAND2_X1 U12002 ( .A1(n9354), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9353) );
  MUX2_X1 U12003 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9353), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n9355) );
  NAND2_X1 U12004 ( .A1(n9355), .A2(n9876), .ZN(n9727) );
  OAI222_X1 U12005 ( .A1(n14252), .A2(n9356), .B1(n10724), .B2(n10821), .C1(
        n9727), .C2(P1_U3086), .ZN(P1_U3345) );
  NAND2_X1 U12006 ( .A1(n9360), .A2(n9358), .ZN(n14236) );
  XNOR2_X2 U12007 ( .A(n9359), .B(n14233), .ZN(n9363) );
  XNOR2_X2 U12008 ( .A(n9361), .B(P1_IR_REG_29__SCAN_IN), .ZN(n9474) );
  NAND2_X2 U12009 ( .A1(n9363), .A2(n9474), .ZN(n11608) );
  INV_X1 U12010 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14094) );
  OR2_X1 U12011 ( .A1(n6426), .A2(n14094), .ZN(n9366) );
  INV_X1 U12012 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n9362) );
  OR2_X1 U12013 ( .A1(n6467), .A2(n9362), .ZN(n9365) );
  INV_X1 U12014 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14201) );
  OR2_X1 U12015 ( .A1(n13453), .A2(n14201), .ZN(n9364) );
  AND3_X1 U12016 ( .A1(n9366), .A2(n9365), .A3(n9364), .ZN(n13503) );
  NAND2_X1 U12017 ( .A1(n13866), .A2(n13750), .ZN(n9367) );
  OAI21_X1 U12018 ( .B1(n9065), .B2(n13750), .A(n9367), .ZN(P1_U3591) );
  INV_X1 U12019 ( .A(n9368), .ZN(n9369) );
  OAI222_X1 U12020 ( .A1(P3_U3151), .A2(n15033), .B1(n12744), .B2(n12263), 
        .C1(n12747), .C2(n9369), .ZN(P3_U3281) );
  INV_X1 U12021 ( .A(n9388), .ZN(n14770) );
  INV_X1 U12022 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n9370) );
  XNOR2_X1 U12023 ( .A(n14755), .B(n9370), .ZN(n14753) );
  XNOR2_X1 U12024 ( .A(n9372), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n14741) );
  NAND2_X1 U12025 ( .A1(n14739), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n14740) );
  INV_X1 U12026 ( .A(n14740), .ZN(n9371) );
  NAND2_X1 U12027 ( .A1(n14741), .A2(n9371), .ZN(n9374) );
  NAND2_X1 U12028 ( .A1(n14742), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n9373) );
  NAND2_X1 U12029 ( .A1(n9374), .A2(n9373), .ZN(n14752) );
  NAND2_X1 U12030 ( .A1(n14755), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9375) );
  XNOR2_X1 U12031 ( .A(n9388), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n14767) );
  XNOR2_X1 U12032 ( .A(n9390), .B(P2_REG1_REG_4__SCAN_IN), .ZN(n9421) );
  NOR2_X1 U12033 ( .A1(n9422), .A2(n9421), .ZN(n9420) );
  XNOR2_X1 U12034 ( .A(n9391), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n9432) );
  INV_X1 U12035 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9376) );
  MUX2_X1 U12036 ( .A(n9376), .B(P2_REG1_REG_6__SCAN_IN), .S(n9561), .Z(n9385)
         );
  NAND2_X1 U12037 ( .A1(n9378), .A2(n9377), .ZN(n9380) );
  NAND2_X1 U12038 ( .A1(n9380), .A2(n9379), .ZN(n9381) );
  NAND2_X1 U12039 ( .A1(n9382), .A2(n9381), .ZN(n9399) );
  NAND2_X1 U12040 ( .A1(n9397), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13290) );
  INV_X1 U12041 ( .A(n13290), .ZN(n9383) );
  NAND2_X1 U12042 ( .A1(n9399), .A2(n9383), .ZN(n9393) );
  INV_X1 U12043 ( .A(n9393), .ZN(n9384) );
  AOI211_X1 U12044 ( .C1(n9386), .C2(n9385), .A(n14795), .B(n9555), .ZN(n9405)
         );
  NAND2_X1 U12045 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14739), .ZN(n14745) );
  NOR2_X1 U12046 ( .A1(n14746), .A2(n14745), .ZN(n14744) );
  AOI21_X1 U12047 ( .B1(n14742), .B2(P2_REG2_REG_1__SCAN_IN), .A(n14744), .ZN(
        n14757) );
  XNOR2_X1 U12048 ( .A(n14755), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n14758) );
  INV_X1 U12049 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9387) );
  INV_X1 U12050 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n9389) );
  MUX2_X1 U12051 ( .A(n9389), .B(P2_REG2_REG_3__SCAN_IN), .S(n9388), .Z(n14774) );
  NAND2_X1 U12052 ( .A1(n14775), .A2(n14774), .ZN(n14773) );
  NAND2_X1 U12053 ( .A1(n14770), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9424) );
  INV_X1 U12054 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n12175) );
  MUX2_X1 U12055 ( .A(n12175), .B(P2_REG2_REG_4__SCAN_IN), .S(n9390), .Z(n9423) );
  NOR2_X1 U12056 ( .A1(n9430), .A2(n12175), .ZN(n9436) );
  INV_X1 U12057 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9941) );
  MUX2_X1 U12058 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n9941), .S(n9391), .Z(n9435)
         );
  OAI21_X1 U12059 ( .B1(n9437), .B2(n9436), .A(n9435), .ZN(n9434) );
  NAND2_X1 U12060 ( .A1(n9391), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9395) );
  INV_X1 U12061 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n9392) );
  MUX2_X1 U12062 ( .A(n9392), .B(P2_REG2_REG_6__SCAN_IN), .S(n9561), .Z(n9394)
         );
  AOI21_X1 U12063 ( .B1(n9434), .B2(n9395), .A(n9394), .ZN(n9560) );
  AND3_X1 U12064 ( .A1(n9434), .A2(n9395), .A3(n9394), .ZN(n9396) );
  NOR3_X1 U12065 ( .A1(n9560), .A2(n14786), .A3(n9396), .ZN(n9404) );
  NOR2_X1 U12066 ( .A1(n9397), .A2(P2_U3088), .ZN(n9398) );
  AND2_X1 U12067 ( .A1(n9399), .A2(n9398), .ZN(n14805) );
  OR2_X1 U12068 ( .A1(n9399), .A2(P2_U3088), .ZN(n14793) );
  INV_X1 U12069 ( .A(n14793), .ZN(n14799) );
  NAND2_X1 U12070 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3088), .ZN(n9774) );
  INV_X1 U12071 ( .A(n9774), .ZN(n9400) );
  AOI21_X1 U12072 ( .B1(n14799), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n9400), .ZN(
        n9401) );
  OAI21_X1 U12073 ( .B1(n9402), .B2(n12878), .A(n9401), .ZN(n9403) );
  OR3_X1 U12074 ( .A1(n9405), .A2(n9404), .A3(n9403), .ZN(P2_U3220) );
  INV_X1 U12075 ( .A(n9406), .ZN(n10488) );
  NAND2_X1 U12076 ( .A1(n10488), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n9408) );
  INV_X1 U12077 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9604) );
  MUX2_X1 U12078 ( .A(n9604), .B(P1_REG2_REG_9__SCAN_IN), .S(n10493), .Z(n9407) );
  AOI21_X1 U12079 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n9611) );
  NAND3_X1 U12080 ( .A1(n9409), .A2(n9408), .A3(n9407), .ZN(n9410) );
  INV_X1 U12081 ( .A(n13851), .ZN(n14641) );
  NAND2_X1 U12082 ( .A1(n9410), .A2(n14641), .ZN(n9419) );
  INV_X1 U12083 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10498) );
  MUX2_X1 U12084 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10498), .S(n10493), .Z(
        n9413) );
  OAI21_X1 U12085 ( .B1(n9413), .B2(n9412), .A(n9601), .ZN(n9414) );
  NAND2_X1 U12086 ( .A1(n9414), .A2(n14640), .ZN(n9418) );
  NOR2_X1 U12087 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11044), .ZN(n9416) );
  NOR2_X1 U12088 ( .A1(n13807), .A2(n9605), .ZN(n9415) );
  AOI211_X1 U12089 ( .C1(n14627), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n9416), .B(
        n9415), .ZN(n9417) );
  OAI211_X1 U12090 ( .C1(n9611), .C2(n9419), .A(n9418), .B(n9417), .ZN(
        P1_U3252) );
  AOI211_X1 U12091 ( .C1(n9422), .C2(n9421), .A(n9420), .B(n14795), .ZN(n9427)
         );
  AND3_X1 U12092 ( .A1(n14773), .A2(n9424), .A3(n9423), .ZN(n9425) );
  NOR3_X1 U12093 ( .A1(n14786), .A2(n9437), .A3(n9425), .ZN(n9426) );
  NOR2_X1 U12094 ( .A1(n9427), .A2(n9426), .ZN(n9429) );
  AND2_X1 U12095 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n9691) );
  AOI21_X1 U12096 ( .B1(n14799), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n9691), .ZN(
        n9428) );
  OAI211_X1 U12097 ( .C1(n9430), .C2(n12878), .A(n9429), .B(n9428), .ZN(
        P2_U3218) );
  AOI211_X1 U12098 ( .C1(n9433), .C2(n9432), .A(n9431), .B(n14795), .ZN(n9441)
         );
  INV_X1 U12099 ( .A(n9434), .ZN(n9439) );
  NOR3_X1 U12100 ( .A1(n9437), .A2(n9436), .A3(n9435), .ZN(n9438) );
  NOR3_X1 U12101 ( .A1(n14786), .A2(n9439), .A3(n9438), .ZN(n9440) );
  NOR2_X1 U12102 ( .A1(n9441), .A2(n9440), .ZN(n9444) );
  NAND2_X1 U12103 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n9758) );
  INV_X1 U12104 ( .A(n9758), .ZN(n9442) );
  AOI21_X1 U12105 ( .B1(n14799), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n9442), .ZN(
        n9443) );
  OAI211_X1 U12106 ( .C1(n9445), .C2(n12878), .A(n9444), .B(n9443), .ZN(
        P2_U3219) );
  INV_X1 U12107 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n14234) );
  NAND2_X1 U12108 ( .A1(n12914), .A2(n12871), .ZN(n9446) );
  OAI21_X1 U12109 ( .B1(n14234), .B2(n12871), .A(n9446), .ZN(P2_U3562) );
  INV_X1 U12110 ( .A(n14640), .ZN(n13819) );
  AOI211_X1 U12111 ( .C1(n9449), .C2(n9448), .A(n13819), .B(n9447), .ZN(n9459)
         );
  INV_X1 U12112 ( .A(n9450), .ZN(n9454) );
  NAND3_X1 U12113 ( .A1(n9463), .A2(n9452), .A3(n9451), .ZN(n9453) );
  NAND3_X1 U12114 ( .A1(n9454), .A2(n14641), .A3(n9453), .ZN(n9456) );
  AND2_X1 U12115 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10719) );
  AOI21_X1 U12116 ( .B1(n14627), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10719), .ZN(
        n9455) );
  OAI211_X1 U12117 ( .C1(n13807), .C2(n9457), .A(n9456), .B(n9455), .ZN(n9458)
         );
  OR2_X1 U12118 ( .A1(n9459), .A2(n9458), .ZN(P1_U3250) );
  AOI211_X1 U12119 ( .C1(n9462), .C2(n9461), .A(n9460), .B(n13819), .ZN(n9473)
         );
  INV_X1 U12120 ( .A(n9463), .ZN(n9468) );
  NOR3_X1 U12121 ( .A1(n9466), .A2(n9465), .A3(n9464), .ZN(n9467) );
  NOR3_X1 U12122 ( .A1(n9468), .A2(n9467), .A3(n13851), .ZN(n9472) );
  NOR2_X1 U12123 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10223), .ZN(n10629) );
  AOI21_X1 U12124 ( .B1(n14627), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n10629), .ZN(
        n9469) );
  OAI21_X1 U12125 ( .B1(n13807), .B2(n9470), .A(n9469), .ZN(n9471) );
  OR3_X1 U12126 ( .A1(n9473), .A2(n9472), .A3(n9471), .ZN(P1_U3249) );
  NAND2_X1 U12127 ( .A1(n13450), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n9480) );
  OR2_X1 U12128 ( .A1(n6465), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9479) );
  INV_X1 U12129 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9476) );
  OR2_X1 U12130 ( .A1(n6428), .A2(n9476), .ZN(n9478) );
  OR2_X1 U12131 ( .A1(n6467), .A2(n9311), .ZN(n9477) );
  AND4_X2 U12132 ( .A1(n9480), .A2(n9479), .A3(n9478), .A4(n9477), .ZN(n9883)
         );
  MUX2_X1 U12133 ( .A(n12233), .B(n9883), .S(n13750), .Z(n9481) );
  INV_X1 U12134 ( .A(n9481), .ZN(P1_U3563) );
  INV_X1 U12135 ( .A(n9499), .ZN(n9505) );
  NOR2_X1 U12136 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .ZN(
        n9485) );
  NOR4_X1 U12137 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_29__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n9484) );
  NOR4_X1 U12138 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9483) );
  NOR4_X1 U12139 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9482) );
  AND4_X1 U12140 ( .A1(n9485), .A2(n9484), .A3(n9483), .A4(n9482), .ZN(n9491)
         );
  NOR4_X1 U12141 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n9489) );
  NOR4_X1 U12142 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n9488) );
  NOR4_X1 U12143 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n9487) );
  NOR4_X1 U12144 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n9486) );
  AND4_X1 U12145 ( .A1(n9489), .A2(n9488), .A3(n9487), .A4(n9486), .ZN(n9490)
         );
  NAND2_X1 U12146 ( .A1(n9491), .A2(n9490), .ZN(n9492) );
  NAND2_X1 U12147 ( .A1(n9505), .A2(n9492), .ZN(n9539) );
  NAND2_X1 U12148 ( .A1(n9539), .A2(n9542), .ZN(n9538) );
  INV_X1 U12149 ( .A(n13457), .ZN(n9498) );
  NAND2_X1 U12150 ( .A1(n10460), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9494) );
  MUX2_X1 U12151 ( .A(P1_IR_REG_31__SCAN_IN), .B(n9494), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n9496) );
  NAND2_X1 U12152 ( .A1(n10954), .A2(n13920), .ZN(n9497) );
  AND2_X1 U12153 ( .A1(n9498), .A2(n9497), .ZN(n13716) );
  OAI22_X1 U12154 ( .A1(n9499), .A2(P1_D_REG_1__SCAN_IN), .B1(n14244), .B2(
        n14248), .ZN(n9781) );
  NAND2_X1 U12155 ( .A1(n10954), .A2(n9526), .ZN(n13456) );
  INV_X1 U12156 ( .A(n13456), .ZN(n9501) );
  NAND2_X1 U12157 ( .A1(n9781), .A2(n9785), .ZN(n9502) );
  INV_X1 U12158 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n9504) );
  NOR2_X1 U12159 ( .A1(n11448), .A2(n14244), .ZN(n9503) );
  INV_X1 U12160 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n14618) );
  AND2_X1 U12161 ( .A1(n13457), .A2(n13920), .ZN(n9507) );
  NAND2_X1 U12162 ( .A1(n14254), .A2(n13920), .ZN(n9506) );
  OR2_X1 U12163 ( .A1(n13456), .A2(n13920), .ZN(n14716) );
  NAND2_X1 U12164 ( .A1(n9508), .A2(n13442), .ZN(n13441) );
  INV_X1 U12165 ( .A(n13920), .ZN(n11513) );
  NAND2_X1 U12166 ( .A1(n11513), .A2(n14254), .ZN(n9509) );
  NOR2_X1 U12167 ( .A1(n14725), .A2(n14183), .ZN(n9528) );
  NAND2_X1 U12168 ( .A1(n9632), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9514) );
  INV_X1 U12169 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10635) );
  OR2_X1 U12170 ( .A1(n6465), .A2(n10635), .ZN(n9513) );
  INV_X1 U12171 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9510) );
  OR2_X1 U12172 ( .A1(n6428), .A2(n9510), .ZN(n9511) );
  NOR2_X1 U12173 ( .A1(n11553), .A2(n9515), .ZN(n9516) );
  XNOR2_X1 U12174 ( .A(n9516), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14255) );
  NAND2_X1 U12175 ( .A1(n9745), .A2(n6434), .ZN(n9711) );
  INV_X1 U12176 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n9518) );
  INV_X1 U12177 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9519) );
  OR2_X1 U12178 ( .A1(n11606), .A2(n9519), .ZN(n9523) );
  NAND2_X1 U12179 ( .A1(n9710), .A2(n14083), .ZN(n10636) );
  NAND3_X1 U12180 ( .A1(n6434), .A2(n13440), .A3(n9526), .ZN(n9527) );
  OAI211_X1 U12181 ( .C1(n9528), .C2(n13524), .A(n10636), .B(n9527), .ZN(n9574) );
  NAND2_X1 U12182 ( .A1(n9574), .A2(n14734), .ZN(n9529) );
  OAI21_X1 U12183 ( .B1(n14734), .B2(n14618), .A(n9529), .ZN(P1_U3528) );
  INV_X1 U12184 ( .A(n9530), .ZN(n9531) );
  OAI222_X1 U12185 ( .A1(n12744), .A2(n9532), .B1(n12747), .B2(n9531), .C1(
        n12344), .C2(P3_U3151), .ZN(P3_U3280) );
  OAI222_X1 U12186 ( .A1(n9544), .A2(n14618), .B1(n11979), .B2(n6666), .C1(
        n9744), .C2(n10324), .ZN(n9627) );
  INV_X2 U12187 ( .A(n9623), .ZN(n11930) );
  AOI222_X1 U12188 ( .A1(n13752), .A2(n11930), .B1(n6434), .B2(n11932), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(n9534), .ZN(n9626) );
  XOR2_X1 U12189 ( .A(n9627), .B(n9626), .Z(n9657) );
  INV_X1 U12190 ( .A(n9781), .ZN(n9535) );
  NAND2_X1 U12191 ( .A1(n9782), .A2(n9535), .ZN(n9548) );
  NAND2_X1 U12192 ( .A1(n13505), .A2(n9526), .ZN(n9786) );
  NAND3_X1 U12193 ( .A1(n13440), .A2(n11513), .A3(n9526), .ZN(n9536) );
  NAND2_X1 U12194 ( .A1(n14587), .A2(n13457), .ZN(n9537) );
  INV_X1 U12195 ( .A(n9539), .ZN(n9540) );
  OR2_X1 U12196 ( .A1(n9548), .A2(n9540), .ZN(n9541) );
  NAND2_X1 U12197 ( .A1(n9541), .A2(n9785), .ZN(n9547) );
  AND2_X1 U12198 ( .A1(n9547), .A2(n9542), .ZN(n13422) );
  NAND2_X1 U12199 ( .A1(n9544), .A2(n9543), .ZN(n9545) );
  NOR2_X1 U12200 ( .A1(n13716), .A2(n9545), .ZN(n9546) );
  NAND2_X1 U12201 ( .A1(n9547), .A2(n9546), .ZN(n9891) );
  NOR2_X1 U12202 ( .A1(n9891), .A2(P1_U3086), .ZN(n9685) );
  INV_X1 U12203 ( .A(n9710), .ZN(n9716) );
  OAI22_X1 U12204 ( .A1(n9685), .A2(n10635), .B1(n14565), .B2(n9716), .ZN(
        n9549) );
  AOI21_X1 U12205 ( .B1(n6434), .B2(n14576), .A(n9549), .ZN(n9550) );
  OAI21_X1 U12206 ( .B1(n9657), .B2(n14570), .A(n9550), .ZN(P1_U3232) );
  INV_X1 U12207 ( .A(n10912), .ZN(n9553) );
  NAND2_X1 U12208 ( .A1(n9876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9551) );
  XNOR2_X1 U12209 ( .A(n9551), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10913) );
  INV_X1 U12210 ( .A(n10913), .ZN(n9817) );
  OAI222_X1 U12211 ( .A1(n14252), .A2(n9552), .B1(n10724), .B2(n9553), .C1(
        P1_U3086), .C2(n9817), .ZN(P1_U3344) );
  INV_X1 U12212 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n9554) );
  INV_X1 U12213 ( .A(n10308), .ZN(n10135) );
  OAI222_X1 U12214 ( .A1(n13303), .A2(n9554), .B1(n13301), .B2(n9553), .C1(
        P2_U3088), .C2(n10135), .ZN(P2_U3316) );
  AOI21_X1 U12215 ( .B1(P2_REG1_REG_6__SCAN_IN), .B2(n9561), .A(n9555), .ZN(
        n14782) );
  INV_X1 U12216 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9556) );
  MUX2_X1 U12217 ( .A(n9556), .B(P2_REG1_REG_7__SCAN_IN), .S(n14785), .Z(
        n14781) );
  NOR2_X1 U12218 ( .A1(n14782), .A2(n14781), .ZN(n14780) );
  AOI21_X1 U12219 ( .B1(P2_REG1_REG_7__SCAN_IN), .B2(n14785), .A(n14780), .ZN(
        n9559) );
  INV_X1 U12220 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n9557) );
  MUX2_X1 U12221 ( .A(n9557), .B(P2_REG1_REG_8__SCAN_IN), .S(n9590), .Z(n9558)
         );
  AOI211_X1 U12222 ( .C1(n9559), .C2(n9558), .A(n14795), .B(n9584), .ZN(n9571)
         );
  AOI21_X1 U12223 ( .B1(P2_REG2_REG_6__SCAN_IN), .B2(n9561), .A(n9560), .ZN(
        n14788) );
  INV_X1 U12224 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n9562) );
  MUX2_X1 U12225 ( .A(n9562), .B(P2_REG2_REG_7__SCAN_IN), .S(n14785), .Z(
        n14787) );
  OR2_X1 U12226 ( .A1(n14788), .A2(n14787), .ZN(n14789) );
  NAND2_X1 U12227 ( .A1(n14785), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9565) );
  INV_X1 U12228 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9563) );
  MUX2_X1 U12229 ( .A(n9563), .B(P2_REG2_REG_8__SCAN_IN), .S(n9590), .Z(n9564)
         );
  AND3_X1 U12230 ( .A1(n14789), .A2(n9565), .A3(n9564), .ZN(n9566) );
  NOR3_X1 U12231 ( .A1(n9589), .A2(n9566), .A3(n14786), .ZN(n9570) );
  NAND2_X1 U12232 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n10147) );
  NAND2_X1 U12233 ( .A1(n14799), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9567) );
  OAI211_X1 U12234 ( .C1(n12878), .C2(n9568), .A(n10147), .B(n9567), .ZN(n9569) );
  OR3_X1 U12235 ( .A1(n9571), .A2(n9570), .A3(n9569), .ZN(P2_U3222) );
  INV_X1 U12236 ( .A(n9782), .ZN(n9572) );
  NAND2_X1 U12237 ( .A1(n9574), .A2(n14729), .ZN(n9575) );
  OAI21_X1 U12238 ( .B1(n14729), .B2(n9510), .A(n9575), .ZN(P1_U3459) );
  INV_X1 U12239 ( .A(n9576), .ZN(n9577) );
  OAI222_X1 U12240 ( .A1(n12744), .A2(n12244), .B1(n12747), .B2(n9577), .C1(
        n12322), .C2(P3_U3151), .ZN(P3_U3279) );
  INV_X1 U12241 ( .A(n14499), .ZN(n12846) );
  INV_X1 U12242 ( .A(n12783), .ZN(n14496) );
  OAI22_X1 U12243 ( .A1(n9931), .A2(n12913), .B1(n12843), .B2(n11471), .ZN(
        n10537) );
  OR2_X1 U12244 ( .A1(n9578), .A2(P2_U3088), .ZN(n11626) );
  AOI22_X1 U12245 ( .A1(n14496), .A2(n10537), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n11626), .ZN(n9583) );
  OAI21_X1 U12246 ( .B1(n9580), .B2(n9579), .A(n9647), .ZN(n9581) );
  NAND2_X1 U12247 ( .A1(n9581), .A2(n14494), .ZN(n9582) );
  OAI211_X1 U12248 ( .C1(n10545), .C2(n12846), .A(n9583), .B(n9582), .ZN(
        P2_U3209) );
  INV_X1 U12249 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9585) );
  MUX2_X1 U12250 ( .A(n9585), .B(P2_REG1_REG_9__SCAN_IN), .S(n9591), .Z(n9586)
         );
  OAI21_X1 U12251 ( .B1(n9587), .B2(n9586), .A(n9795), .ZN(n9588) );
  NAND2_X1 U12252 ( .A1(n9588), .A2(n14765), .ZN(n9600) );
  AOI21_X1 U12253 ( .B1(n9590), .B2(P2_REG2_REG_8__SCAN_IN), .A(n9589), .ZN(
        n9594) );
  INV_X1 U12254 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U12255 ( .A(n9592), .B(P2_REG2_REG_9__SCAN_IN), .S(n9591), .Z(n9593)
         );
  NAND2_X1 U12256 ( .A1(n9594), .A2(n9593), .ZN(n9798) );
  OAI21_X1 U12257 ( .B1(n9594), .B2(n9593), .A(n9798), .ZN(n9598) );
  INV_X1 U12258 ( .A(n14786), .ZN(n14800) );
  INV_X1 U12259 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U12260 ( .A1(n14805), .A2(n9799), .ZN(n9595) );
  NAND2_X1 U12261 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10642) );
  OAI211_X1 U12262 ( .C1(n14793), .C2(n9596), .A(n9595), .B(n10642), .ZN(n9597) );
  AOI21_X1 U12263 ( .B1(n9598), .B2(n14800), .A(n9597), .ZN(n9599) );
  NAND2_X1 U12264 ( .A1(n9600), .A2(n9599), .ZN(P2_U3223) );
  INV_X1 U12265 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n10514) );
  MUX2_X1 U12266 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n10514), .S(n9727), .Z(
        n9603) );
  OAI21_X1 U12267 ( .B1(n10493), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9601), .ZN(
        n9602) );
  NOR2_X1 U12268 ( .A1(n9602), .A2(n9603), .ZN(n9728) );
  AOI211_X1 U12269 ( .C1(n9603), .C2(n9602), .A(n13819), .B(n9728), .ZN(n9616)
         );
  INV_X1 U12270 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9726) );
  MUX2_X1 U12271 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9726), .S(n9727), .Z(n9607) );
  NOR2_X1 U12272 ( .A1(n9605), .A2(n9604), .ZN(n9609) );
  INV_X1 U12273 ( .A(n9609), .ZN(n9606) );
  NAND2_X1 U12274 ( .A1(n9607), .A2(n9606), .ZN(n9610) );
  MUX2_X1 U12275 ( .A(n9726), .B(P1_REG2_REG_10__SCAN_IN), .S(n9727), .Z(n9608) );
  OAI21_X1 U12276 ( .B1(n9611), .B2(n9609), .A(n9608), .ZN(n9725) );
  OAI211_X1 U12277 ( .C1(n9611), .C2(n9610), .A(n9725), .B(n14641), .ZN(n9614)
         );
  INV_X1 U12278 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n14550) );
  NOR2_X1 U12279 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14550), .ZN(n9612) );
  AOI21_X1 U12280 ( .B1(n14627), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9612), .ZN(
        n9613) );
  OAI211_X1 U12281 ( .C1(n13807), .C2(n9727), .A(n9614), .B(n9613), .ZN(n9615)
         );
  OR2_X1 U12282 ( .A1(n9616), .A2(n9615), .ZN(P1_U3253) );
  OR2_X1 U12283 ( .A1(n13464), .A2(n6935), .ZN(n9620) );
  AND3_X2 U12284 ( .A1(n9621), .A2(n9620), .A3(n9619), .ZN(n13523) );
  INV_X1 U12285 ( .A(n13523), .ZN(n9737) );
  XOR2_X1 U12286 ( .A(n11853), .B(n9622), .Z(n9625) );
  OAI22_X1 U12287 ( .A1(n9716), .A2(n11978), .B1(n13523), .B2(n11979), .ZN(
        n9624) );
  OAI21_X1 U12288 ( .B1(n6487), .B2(n9630), .A(n9679), .ZN(n9631) );
  NAND2_X1 U12289 ( .A1(n9631), .A2(n14553), .ZN(n9642) );
  INV_X1 U12290 ( .A(n9685), .ZN(n9640) );
  INV_X1 U12291 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9684) );
  OR2_X1 U12292 ( .A1(n11606), .A2(n9684), .ZN(n9637) );
  INV_X1 U12293 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9634) );
  OR2_X1 U12294 ( .A1(n13453), .A2(n9634), .ZN(n9635) );
  NAND2_X1 U12295 ( .A1(n13332), .A2(n14085), .ZN(n14562) );
  OAI22_X1 U12296 ( .A1(n14565), .A2(n7348), .B1(n6666), .B2(n14562), .ZN(
        n9639) );
  AOI21_X1 U12297 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n9640), .A(n9639), .ZN(
        n9641) );
  OAI211_X1 U12298 ( .C1(n13523), .C2(n13434), .A(n9642), .B(n9641), .ZN(
        P1_U3222) );
  INV_X1 U12299 ( .A(n10929), .ZN(n9644) );
  OAI21_X1 U12300 ( .B1(n9876), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9702) );
  XNOR2_X1 U12301 ( .A(n9702), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10930) );
  INV_X1 U12302 ( .A(n10930), .ZN(n9820) );
  OAI222_X1 U12303 ( .A1(n14252), .A2(n9643), .B1(n10724), .B2(n9644), .C1(
        n9820), .C2(P1_U3086), .ZN(P1_U3343) );
  INV_X1 U12304 ( .A(n10696), .ZN(n10304) );
  OAI222_X1 U12305 ( .A1(n13303), .A2(n9645), .B1(n13301), .B2(n9644), .C1(
        n10304), .C2(P2_U3088), .ZN(P2_U3315) );
  AND2_X1 U12306 ( .A1(n9647), .A2(n9646), .ZN(n9694) );
  XNOR2_X1 U12307 ( .A(n9693), .B(n9694), .ZN(n9652) );
  INV_X1 U12308 ( .A(n12913), .ZN(n12781) );
  AOI22_X1 U12309 ( .A1(n12781), .A2(n12867), .B1(n12947), .B2(n12869), .ZN(
        n14812) );
  NAND2_X1 U12310 ( .A1(n14499), .A2(n9932), .ZN(n9648) );
  NAND2_X1 U12311 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n14768) );
  OAI211_X1 U12312 ( .C1(n14812), .C2(n12783), .A(n9648), .B(n14768), .ZN(
        n9649) );
  AOI21_X1 U12313 ( .B1(n12842), .B2(n9650), .A(n9649), .ZN(n9651) );
  OAI21_X1 U12314 ( .B1(n9652), .B2(n12816), .A(n9651), .ZN(P2_U3190) );
  OAI22_X1 U12315 ( .A1(n12349), .A2(P3_U3151), .B1(n9653), .B2(n12726), .ZN(
        n9654) );
  AOI21_X1 U12316 ( .B1(n9655), .B2(n14376), .A(n9654), .ZN(n9656) );
  INV_X1 U12317 ( .A(n9656), .ZN(P3_U3278) );
  NAND2_X1 U12318 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n13753) );
  INV_X1 U12319 ( .A(n9657), .ZN(n9658) );
  MUX2_X1 U12320 ( .A(n13753), .B(n9658), .S(n14619), .Z(n9660) );
  NOR2_X1 U12321 ( .A1(n14619), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9659) );
  OR2_X1 U12322 ( .A1(n6468), .A2(n9659), .ZN(n14617) );
  NAND2_X1 U12323 ( .A1(n14617), .A2(n14621), .ZN(n14624) );
  OAI211_X1 U12324 ( .C1(n9660), .C2(n6468), .A(n13750), .B(n14624), .ZN(
        n13777) );
  INV_X1 U12325 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9665) );
  XOR2_X1 U12326 ( .A(n9662), .B(n9661), .Z(n9663) );
  NAND2_X1 U12327 ( .A1(n14640), .A2(n9663), .ZN(n9664) );
  NAND2_X1 U12328 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10410) );
  OAI211_X1 U12329 ( .C1(n9665), .C2(n14645), .A(n9664), .B(n10410), .ZN(n9672) );
  INV_X1 U12330 ( .A(n9666), .ZN(n9670) );
  NOR3_X1 U12331 ( .A1(n13784), .A2(n9668), .A3(n9667), .ZN(n9669) );
  NOR3_X1 U12332 ( .A1(n13851), .A2(n9670), .A3(n9669), .ZN(n9671) );
  AOI211_X1 U12333 ( .C1(n14637), .C2(n9837), .A(n9672), .B(n9671), .ZN(n9673)
         );
  NAND2_X1 U12334 ( .A1(n13777), .A2(n9673), .ZN(P1_U3247) );
  AOI22_X1 U12335 ( .A1(n7349), .A2(n11966), .B1(n13749), .B2(n11932), .ZN(
        n9677) );
  XNOR2_X1 U12336 ( .A(n9677), .B(n11853), .ZN(n9884) );
  NAND2_X1 U12337 ( .A1(n11930), .A2(n13749), .ZN(n9678) );
  OAI21_X1 U12338 ( .B1(n10597), .B2(n11979), .A(n9678), .ZN(n9885) );
  XNOR2_X1 U12339 ( .A(n9884), .B(n9885), .ZN(n9681) );
  NAND2_X1 U12340 ( .A1(n9680), .A2(n9681), .ZN(n9888) );
  OAI21_X1 U12341 ( .B1(n9681), .B2(n9680), .A(n9888), .ZN(n9687) );
  INV_X1 U12342 ( .A(n14562), .ZN(n13409) );
  AOI22_X1 U12343 ( .A1(n13409), .A2(n9710), .B1(n13418), .B2(n9835), .ZN(
        n9683) );
  NAND2_X1 U12344 ( .A1(n14576), .A2(n7349), .ZN(n9682) );
  OAI211_X1 U12345 ( .C1(n9685), .C2(n9684), .A(n9683), .B(n9682), .ZN(n9686)
         );
  AOI21_X1 U12346 ( .B1(n9687), .B2(n14553), .A(n9686), .ZN(n9688) );
  INV_X1 U12347 ( .A(n9688), .ZN(P1_U3237) );
  INV_X1 U12348 ( .A(n9689), .ZN(n10175) );
  OAI22_X1 U12349 ( .A1(n10155), .A2(n12913), .B1(n12843), .B2(n9931), .ZN(
        n10172) );
  NOR2_X1 U12350 ( .A1(n12846), .A2(n14887), .ZN(n9690) );
  AOI211_X1 U12351 ( .C1(n14496), .C2(n10172), .A(n9691), .B(n9690), .ZN(n9701) );
  AOI21_X1 U12352 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9698) );
  INV_X1 U12353 ( .A(n9695), .ZN(n9697) );
  OAI21_X1 U12354 ( .B1(n9698), .B2(n9697), .A(n9696), .ZN(n9699) );
  NAND2_X1 U12355 ( .A1(n9699), .A2(n14494), .ZN(n9700) );
  OAI211_X1 U12356 ( .C1(n14502), .C2(n10175), .A(n9701), .B(n9700), .ZN(
        P2_U3202) );
  INV_X1 U12357 ( .A(n11091), .ZN(n9706) );
  INV_X1 U12358 ( .A(n10868), .ZN(n10703) );
  OAI222_X1 U12359 ( .A1(n13303), .A2(n12205), .B1(n13301), .B2(n9706), .C1(
        n10703), .C2(P2_U3088), .ZN(P2_U3314) );
  INV_X1 U12360 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9873) );
  NAND2_X1 U12361 ( .A1(n9702), .A2(n9873), .ZN(n9703) );
  NAND2_X1 U12362 ( .A1(n9703), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9704) );
  INV_X1 U12363 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n9872) );
  NAND2_X1 U12364 ( .A1(n9704), .A2(n9872), .ZN(n9763) );
  OR2_X1 U12365 ( .A1(n9704), .A2(n9872), .ZN(n9705) );
  INV_X1 U12366 ( .A(n13802), .ZN(n10421) );
  OAI222_X1 U12367 ( .A1(n14252), .A2(n9707), .B1(n10724), .B2(n9706), .C1(
        n10421), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12368 ( .A(P3_DATAO_REG_1__SCAN_IN), .ZN(n9709) );
  NAND2_X1 U12369 ( .A1(n10087), .A2(n12284), .ZN(n9708) );
  OAI21_X1 U12370 ( .B1(P3_U3897), .B2(n9709), .A(n9708), .ZN(P3_U3492) );
  NAND2_X1 U12371 ( .A1(n9710), .A2(n13523), .ZN(n13530) );
  INV_X1 U12372 ( .A(n9711), .ZN(n9714) );
  INV_X1 U12373 ( .A(n9739), .ZN(n9713) );
  AOI21_X1 U12374 ( .B1(n13469), .B2(n9714), .A(n9713), .ZN(n9790) );
  AOI21_X1 U12375 ( .B1(n13469), .B2(n13752), .A(n14166), .ZN(n9715) );
  NOR2_X1 U12376 ( .A1(n9715), .A2(n14085), .ZN(n9719) );
  AOI21_X1 U12377 ( .B1(n6434), .B2(n9737), .A(n9742), .ZN(n9720) );
  XNOR2_X1 U12378 ( .A(n9720), .B(n9716), .ZN(n9717) );
  AOI21_X1 U12379 ( .B1(n9717), .B2(n14183), .A(n13752), .ZN(n9718) );
  OAI222_X1 U12380 ( .A1(n14060), .A2(n7348), .B1(n13957), .B2(n9790), .C1(
        n9719), .C2(n9718), .ZN(n9787) );
  INV_X1 U12381 ( .A(n9787), .ZN(n9723) );
  INV_X1 U12382 ( .A(n9720), .ZN(n9721) );
  NOR2_X1 U12383 ( .A1(n9721), .A2(n14075), .ZN(n9788) );
  AOI21_X1 U12384 ( .B1(n9737), .B2(n14712), .A(n9788), .ZN(n9722) );
  OAI211_X1 U12385 ( .C1(n9790), .C2(n14716), .A(n9723), .B(n9722), .ZN(n14199) );
  NAND2_X1 U12386 ( .A1(n14199), .A2(n14729), .ZN(n9724) );
  OAI21_X1 U12387 ( .B1(n14729), .B2(n9518), .A(n9724), .ZN(P1_U3462) );
  INV_X1 U12388 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9816) );
  MUX2_X1 U12389 ( .A(n9816), .B(P1_REG2_REG_11__SCAN_IN), .S(n10913), .Z(
        n9812) );
  OAI21_X1 U12390 ( .B1(n9726), .B2(n9727), .A(n9725), .ZN(n9814) );
  XOR2_X1 U12391 ( .A(n9812), .B(n9814), .Z(n9736) );
  INV_X1 U12392 ( .A(n9727), .ZN(n10822) );
  INV_X1 U12393 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10830) );
  MUX2_X1 U12394 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10830), .S(n10913), .Z(
        n9729) );
  NAND2_X1 U12395 ( .A1(n9730), .A2(n9729), .ZN(n9821) );
  OAI21_X1 U12396 ( .B1(n9730), .B2(n9729), .A(n9821), .ZN(n9731) );
  NAND2_X1 U12397 ( .A1(n9731), .A2(n14640), .ZN(n9735) );
  NAND2_X1 U12398 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n14577)
         );
  INV_X1 U12399 ( .A(n14577), .ZN(n9733) );
  NOR2_X1 U12400 ( .A1(n13807), .A2(n9817), .ZN(n9732) );
  AOI211_X1 U12401 ( .C1(n14627), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n9733), .B(
        n9732), .ZN(n9734) );
  OAI211_X1 U12402 ( .C1(n13851), .C2(n9736), .A(n9735), .B(n9734), .ZN(
        P1_U3254) );
  OR2_X1 U12403 ( .A1(n9737), .A2(n9710), .ZN(n9738) );
  NAND2_X1 U12404 ( .A1(n13749), .A2(n10597), .ZN(n13535) );
  OAI21_X1 U12405 ( .B1(n9741), .B2(n9740), .A(n9831), .ZN(n10601) );
  INV_X1 U12406 ( .A(n9742), .ZN(n9743) );
  AND2_X1 U12407 ( .A1(n9742), .A2(n10597), .ZN(n10119) );
  AOI211_X1 U12408 ( .C1(n7349), .C2(n9743), .A(n14075), .B(n10119), .ZN(
        n10595) );
  OAI21_X1 U12409 ( .B1(n13533), .B2(n9747), .A(n9852), .ZN(n9748) );
  AOI222_X1 U12410 ( .A1(n14183), .A2(n9748), .B1(n9710), .B2(n14085), .C1(
        n9835), .C2(n14083), .ZN(n9749) );
  INV_X1 U12411 ( .A(n9749), .ZN(n10598) );
  AOI211_X1 U12412 ( .C1(n14725), .C2(n10601), .A(n10595), .B(n10598), .ZN(
        n9753) );
  NAND2_X1 U12413 ( .A1(n14729), .A2(n14712), .ZN(n14227) );
  OAI22_X1 U12414 ( .A1(n14227), .A2(n10597), .B1(n14729), .B2(n9634), .ZN(
        n9750) );
  INV_X1 U12415 ( .A(n9750), .ZN(n9751) );
  OAI21_X1 U12416 ( .B1(n9753), .B2(n14727), .A(n9751), .ZN(P1_U3465) );
  NAND2_X1 U12417 ( .A1(n14734), .A2(n14712), .ZN(n14172) );
  INV_X1 U12418 ( .A(n14172), .ZN(n10857) );
  AOI22_X1 U12419 ( .A1(n10857), .A2(n7349), .B1(n14732), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n9752) );
  OAI21_X1 U12420 ( .B1(n9753), .B2(n14732), .A(n9752), .ZN(P1_U3530) );
  OAI21_X1 U12421 ( .B1(n9756), .B2(n9755), .A(n9754), .ZN(n9757) );
  NAND2_X1 U12422 ( .A1(n9757), .A2(n14494), .ZN(n9762) );
  OAI22_X1 U12423 ( .A1(n10242), .A2(n12913), .B1(n12843), .B2(n9934), .ZN(
        n9939) );
  INV_X1 U12424 ( .A(n9939), .ZN(n9759) );
  OAI21_X1 U12425 ( .B1(n12783), .B2(n9759), .A(n9758), .ZN(n9760) );
  AOI21_X1 U12426 ( .B1(n9942), .B2(n14499), .A(n9760), .ZN(n9761) );
  OAI211_X1 U12427 ( .C1(n14502), .C2(n9944), .A(n9762), .B(n9761), .ZN(
        P2_U3199) );
  INV_X1 U12428 ( .A(n11185), .ZN(n11188) );
  INV_X1 U12429 ( .A(n11220), .ZN(n9765) );
  OAI222_X1 U12430 ( .A1(P2_U3088), .A2(n11188), .B1(n13301), .B2(n9765), .C1(
        n12226), .C2(n13303), .ZN(P2_U3313) );
  NAND2_X1 U12431 ( .A1(n9763), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9764) );
  XNOR2_X1 U12432 ( .A(n9764), .B(P1_IR_REG_14__SCAN_IN), .ZN(n11221) );
  INV_X1 U12433 ( .A(n11221), .ZN(n10998) );
  OAI222_X1 U12434 ( .A1(n14252), .A2(n9766), .B1(n10724), .B2(n9765), .C1(
        n10998), .C2(P1_U3086), .ZN(P1_U3341) );
  INV_X1 U12435 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n9768) );
  NAND2_X1 U12436 ( .A1(n11704), .A2(P3_U3897), .ZN(n9767) );
  OAI21_X1 U12437 ( .B1(P3_U3897), .B2(n9768), .A(n9767), .ZN(P3_U3495) );
  XNOR2_X1 U12438 ( .A(n9770), .B(n9769), .ZN(n9779) );
  INV_X1 U12439 ( .A(n9771), .ZN(n10165) );
  NOR2_X1 U12440 ( .A1(n14502), .A2(n10165), .ZN(n9777) );
  OR2_X1 U12441 ( .A1(n10155), .A2(n12843), .ZN(n9772) );
  OAI21_X1 U12442 ( .B1(n12913), .B2(n9773), .A(n9772), .ZN(n10161) );
  INV_X1 U12443 ( .A(n10161), .ZN(n9775) );
  OAI21_X1 U12444 ( .B1(n12783), .B2(n9775), .A(n9774), .ZN(n9776) );
  AOI211_X1 U12445 ( .C1(n14901), .C2(n14499), .A(n9777), .B(n9776), .ZN(n9778) );
  OAI21_X1 U12446 ( .B1(n9779), .B2(n12816), .A(n9778), .ZN(P2_U3211) );
  INV_X1 U12447 ( .A(n9780), .ZN(n9784) );
  NOR2_X1 U12448 ( .A1(n9782), .A2(n9781), .ZN(n9783) );
  NAND2_X1 U12449 ( .A1(n9784), .A2(n9783), .ZN(n13887) );
  AOI21_X1 U12450 ( .B1(n9788), .B2(n13920), .A(n9787), .ZN(n9789) );
  MUX2_X1 U12451 ( .A(n9307), .B(n9789), .S(n14047), .Z(n9793) );
  OR2_X1 U12452 ( .A1(n9533), .A2(n13920), .ZN(n13459) );
  NOR2_X1 U12453 ( .A1(n14650), .A2(n13459), .ZN(n14669) );
  INV_X1 U12454 ( .A(n9790), .ZN(n9791) );
  INV_X1 U12455 ( .A(n14044), .ZN(n14662) );
  AOI22_X1 U12456 ( .A1(n14669), .A2(n9791), .B1(P1_REG3_REG_1__SCAN_IN), .B2(
        n14662), .ZN(n9792) );
  OAI211_X1 U12457 ( .C1(n13523), .C2(n14666), .A(n9793), .B(n9792), .ZN(
        P1_U3292) );
  INV_X1 U12458 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9794) );
  MUX2_X1 U12459 ( .A(n9794), .B(P2_REG1_REG_10__SCAN_IN), .S(n10137), .Z(
        n9797) );
  NOR2_X1 U12460 ( .A1(n9796), .A2(n9797), .ZN(n10136) );
  AOI211_X1 U12461 ( .C1(n9797), .C2(n9796), .A(n14795), .B(n10136), .ZN(n9808) );
  OAI21_X1 U12462 ( .B1(n9799), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9798), .ZN(
        n9802) );
  INV_X1 U12463 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n9800) );
  MUX2_X1 U12464 ( .A(n9800), .B(P2_REG2_REG_10__SCAN_IN), .S(n10137), .Z(
        n9801) );
  AOI211_X1 U12465 ( .C1(n9802), .C2(n9801), .A(n14786), .B(n10128), .ZN(n9807) );
  NAND2_X1 U12466 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n10787)
         );
  INV_X1 U12467 ( .A(n10787), .ZN(n9803) );
  AOI21_X1 U12468 ( .B1(n14799), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n9803), .ZN(
        n9804) );
  OAI21_X1 U12469 ( .B1(n9805), .B2(n12878), .A(n9804), .ZN(n9806) );
  OR3_X1 U12470 ( .A1(n9808), .A2(n9807), .A3(n9806), .ZN(P2_U3224) );
  OAI222_X1 U12471 ( .A1(n12747), .A2(n9810), .B1(n12744), .B2(n9809), .C1(
        P3_U3151), .C2(n12363), .ZN(P3_U3276) );
  INV_X1 U12472 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9811) );
  AOI22_X1 U12473 ( .A1(n10930), .A2(n9811), .B1(P1_REG2_REG_12__SCAN_IN), 
        .B2(n9820), .ZN(n9819) );
  INV_X1 U12474 ( .A(n9812), .ZN(n9813) );
  NAND2_X1 U12475 ( .A1(n9814), .A2(n9813), .ZN(n9815) );
  OAI21_X1 U12476 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9818) );
  NOR2_X1 U12477 ( .A1(n9819), .A2(n9818), .ZN(n10419) );
  AOI21_X1 U12478 ( .B1(n9819), .B2(n9818), .A(n10419), .ZN(n9829) );
  INV_X1 U12479 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14390) );
  AOI22_X1 U12480 ( .A1(n10930), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n14390), 
        .B2(n9820), .ZN(n9823) );
  OAI21_X1 U12481 ( .B1(n9823), .B2(n9822), .A(n10415), .ZN(n9824) );
  NAND2_X1 U12482 ( .A1(n9824), .A2(n14640), .ZN(n9828) );
  NAND2_X1 U12483 ( .A1(n14627), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n9825) );
  NAND2_X1 U12484 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n13342)
         );
  NAND2_X1 U12485 ( .A1(n9825), .A2(n13342), .ZN(n9826) );
  AOI21_X1 U12486 ( .B1(n14637), .B2(n10930), .A(n9826), .ZN(n9827) );
  OAI211_X1 U12487 ( .C1(n9829), .C2(n13851), .A(n9828), .B(n9827), .ZN(
        P1_U3255) );
  OR2_X1 U12488 ( .A1(n7349), .A2(n13749), .ZN(n9830) );
  OR2_X1 U12489 ( .A1(n9832), .A2(n13436), .ZN(n9834) );
  NAND2_X1 U12490 ( .A1(n9883), .A2(n14706), .ZN(n13543) );
  INV_X1 U12491 ( .A(n14706), .ZN(n10124) );
  NAND2_X1 U12492 ( .A1(n10124), .A2(n9835), .ZN(n13544) );
  NAND2_X1 U12493 ( .A1(n9836), .A2(n13461), .ZN(n9839) );
  AOI22_X1 U12494 ( .A1(n11515), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n11514), 
        .B2(n9837), .ZN(n9838) );
  NAND2_X1 U12495 ( .A1(n9839), .A2(n9838), .ZN(n13548) );
  NAND2_X1 U12496 ( .A1(n11600), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9849) );
  OR2_X1 U12497 ( .A1(n6467), .A2(n9840), .ZN(n9848) );
  INV_X1 U12498 ( .A(n9856), .ZN(n9844) );
  INV_X1 U12499 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9842) );
  INV_X1 U12500 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9841) );
  NAND2_X1 U12501 ( .A1(n9842), .A2(n9841), .ZN(n9843) );
  NAND2_X1 U12502 ( .A1(n9844), .A2(n9843), .ZN(n10606) );
  OR2_X1 U12503 ( .A1(n6465), .A2(n10606), .ZN(n9847) );
  INV_X1 U12504 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9845) );
  OR2_X1 U12505 ( .A1(n6426), .A2(n9845), .ZN(n9846) );
  NAND4_X1 U12506 ( .A1(n9849), .A2(n9848), .A3(n9847), .A4(n9846), .ZN(n13748) );
  NAND2_X1 U12507 ( .A1(n10604), .A2(n13748), .ZN(n9850) );
  NAND2_X1 U12508 ( .A1(n13548), .A2(n10338), .ZN(n10220) );
  NAND2_X1 U12509 ( .A1(n9850), .A2(n10220), .ZN(n13471) );
  OAI21_X1 U12510 ( .B1(n9851), .B2(n13471), .A(n10212), .ZN(n10613) );
  INV_X1 U12511 ( .A(n13471), .ZN(n9854) );
  AND2_X1 U12512 ( .A1(n9855), .A2(n14183), .ZN(n10609) );
  NAND2_X1 U12513 ( .A1(n10119), .A2(n10124), .ZN(n10120) );
  AOI211_X1 U12514 ( .C1(n13548), .C2(n10120), .A(n14075), .B(n10234), .ZN(
        n10603) );
  OR2_X1 U12515 ( .A1(n9883), .A2(n14020), .ZN(n9863) );
  NAND2_X1 U12516 ( .A1(n11600), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9861) );
  OR2_X1 U12517 ( .A1(n6467), .A2(n9341), .ZN(n9860) );
  NAND2_X1 U12518 ( .A1(n9856), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10224) );
  OAI21_X1 U12519 ( .B1(n9856), .B2(P1_REG3_REG_5__SCAN_IN), .A(n10224), .ZN(
        n10341) );
  OR2_X1 U12520 ( .A1(n6465), .A2(n10341), .ZN(n9859) );
  OR2_X1 U12521 ( .A1(n6426), .A2(n9857), .ZN(n9858) );
  NAND4_X1 U12522 ( .A1(n9861), .A2(n9860), .A3(n9859), .A4(n9858), .ZN(n13747) );
  NAND2_X1 U12523 ( .A1(n13747), .A2(n14083), .ZN(n9862) );
  NAND2_X1 U12524 ( .A1(n9863), .A2(n9862), .ZN(n10607) );
  OR3_X1 U12525 ( .A1(n10609), .A2(n10603), .A3(n10607), .ZN(n9864) );
  AOI21_X1 U12526 ( .B1(n14725), .B2(n10613), .A(n9864), .ZN(n9870) );
  INV_X1 U12527 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n9865) );
  OAI22_X1 U12528 ( .A1(n14227), .A2(n10604), .B1(n14729), .B2(n9865), .ZN(
        n9866) );
  INV_X1 U12529 ( .A(n9866), .ZN(n9867) );
  OAI21_X1 U12530 ( .B1(n9870), .B2(n14727), .A(n9867), .ZN(P1_U3471) );
  OAI22_X1 U12531 ( .A1(n14172), .A2(n10604), .B1(n14734), .B2(n9845), .ZN(
        n9868) );
  INV_X1 U12532 ( .A(n9868), .ZN(n9869) );
  OAI21_X1 U12533 ( .B1(n9870), .B2(n14732), .A(n9869), .ZN(P1_U3532) );
  INV_X1 U12534 ( .A(n11225), .ZN(n9879) );
  INV_X1 U12535 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n9871) );
  NAND4_X1 U12536 ( .A1(n9874), .A2(n9873), .A3(n9872), .A4(n9871), .ZN(n9875)
         );
  OAI21_X1 U12537 ( .B1(n9876), .B2(n9875), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n9877) );
  XNOR2_X1 U12538 ( .A(n9877), .B(P1_IR_REG_15__SCAN_IN), .ZN(n14638) );
  INV_X1 U12539 ( .A(n14638), .ZN(n11000) );
  OAI222_X1 U12540 ( .A1(n14252), .A2(n9878), .B1(n10724), .B2(n9879), .C1(
        P1_U3086), .C2(n11000), .ZN(P1_U3340) );
  INV_X1 U12541 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9880) );
  INV_X1 U12542 ( .A(n11342), .ZN(n11335) );
  OAI222_X1 U12543 ( .A1(n13303), .A2(n9880), .B1(n13301), .B2(n9879), .C1(
        P2_U3088), .C2(n11335), .ZN(P2_U3312) );
  NAND2_X1 U12544 ( .A1(n14706), .A2(n11966), .ZN(n9881) );
  OAI21_X1 U12545 ( .B1(n9883), .B2(n11979), .A(n9881), .ZN(n9882) );
  XNOR2_X1 U12546 ( .A(n9882), .B(n11853), .ZN(n10322) );
  OAI22_X1 U12547 ( .A1(n10124), .A2(n11979), .B1(n9883), .B2(n11978), .ZN(
        n10323) );
  XNOR2_X1 U12548 ( .A(n10322), .B(n10323), .ZN(n9890) );
  NAND2_X1 U12549 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  NOR2_X1 U12550 ( .A1(n9889), .A2(n9890), .ZN(n10321) );
  AOI211_X1 U12551 ( .C1(n9890), .C2(n9889), .A(n14570), .B(n10321), .ZN(n9895) );
  AOI22_X1 U12552 ( .A1(n13409), .A2(n13749), .B1(n13418), .B2(n13748), .ZN(
        n9893) );
  MUX2_X1 U12553 ( .A(n14580), .B(P1_STATE_REG_SCAN_IN), .S(
        P1_REG3_REG_3__SCAN_IN), .Z(n9892) );
  OAI211_X1 U12554 ( .C1(n13434), .C2(n10124), .A(n9893), .B(n9892), .ZN(n9894) );
  OR2_X1 U12555 ( .A1(n9895), .A2(n9894), .ZN(P1_U3218) );
  XNOR2_X1 U12556 ( .A(n9897), .B(n9896), .ZN(n9903) );
  OR2_X1 U12557 ( .A1(n10242), .A2(n12843), .ZN(n9898) );
  OAI21_X1 U12558 ( .B1(n12913), .B2(n10475), .A(n9898), .ZN(n9899) );
  INV_X1 U12559 ( .A(n9899), .ZN(n10452) );
  INV_X1 U12560 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n14779) );
  OAI22_X1 U12561 ( .A1(n12783), .A2(n10452), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n14779), .ZN(n9901) );
  INV_X1 U12562 ( .A(n10443), .ZN(n14909) );
  NOR2_X1 U12563 ( .A1(n12846), .A2(n14909), .ZN(n9900) );
  AOI211_X1 U12564 ( .C1(n12842), .C2(n10442), .A(n9901), .B(n9900), .ZN(n9902) );
  OAI21_X1 U12565 ( .B1(n9903), .B2(n12816), .A(n9902), .ZN(P2_U3185) );
  NOR2_X1 U12566 ( .A1(n12117), .A2(P3_U3151), .ZN(n10438) );
  NAND2_X1 U12567 ( .A1(n12285), .A2(n10785), .ZN(n11678) );
  AND2_X1 U12568 ( .A1(n11681), .A2(n11678), .ZN(n11819) );
  INV_X1 U12569 ( .A(n11819), .ZN(n9905) );
  INV_X1 U12570 ( .A(n12132), .ZN(n12114) );
  OAI22_X1 U12571 ( .A1(n12114), .A2(n10785), .B1(n15088), .B2(n12109), .ZN(
        n9904) );
  AOI21_X1 U12572 ( .B1(n6997), .B2(n9905), .A(n9904), .ZN(n9906) );
  OAI21_X1 U12573 ( .B1(n10438), .B2(n9907), .A(n9906), .ZN(P3_U3172) );
  NAND2_X1 U12574 ( .A1(n9909), .A2(n9908), .ZN(n11148) );
  INV_X1 U12575 ( .A(n11148), .ZN(n9912) );
  INV_X1 U12576 ( .A(n14853), .ZN(n9910) );
  AND3_X1 U12577 ( .A1(n9910), .A2(n14854), .A3(n14850), .ZN(n9911) );
  NAND2_X1 U12578 ( .A1(n9912), .A2(n9911), .ZN(n9915) );
  INV_X1 U12579 ( .A(n9913), .ZN(n9914) );
  OR2_X1 U12580 ( .A1(n14844), .A2(n9914), .ZN(n14840) );
  NAND2_X1 U12581 ( .A1(n14507), .A2(n9916), .ZN(n9917) );
  NAND2_X1 U12582 ( .A1(n14855), .A2(n12872), .ZN(n11633) );
  NAND2_X1 U12583 ( .A1(n9918), .A2(n11633), .ZN(n9920) );
  NAND2_X1 U12584 ( .A1(n14865), .A2(n11471), .ZN(n9919) );
  NAND2_X1 U12585 ( .A1(n10540), .A2(n10539), .ZN(n9922) );
  NAND2_X1 U12586 ( .A1(n10545), .A2(n11625), .ZN(n9921) );
  NAND2_X1 U12587 ( .A1(n9922), .A2(n9921), .ZN(n14827) );
  INV_X1 U12588 ( .A(n14810), .ZN(n14826) );
  NAND2_X1 U12589 ( .A1(n14827), .A2(n14826), .ZN(n9924) );
  NAND2_X1 U12590 ( .A1(n14879), .A2(n9931), .ZN(n9923) );
  INV_X1 U12591 ( .A(n10170), .ZN(n9925) );
  NAND2_X1 U12592 ( .A1(n14887), .A2(n9934), .ZN(n9926) );
  XNOR2_X1 U12593 ( .A(n10154), .B(n10152), .ZN(n14896) );
  INV_X1 U12594 ( .A(n9927), .ZN(n11638) );
  NAND2_X1 U12595 ( .A1(n11644), .A2(n11471), .ZN(n9928) );
  INV_X1 U12596 ( .A(n10539), .ZN(n10535) );
  NAND2_X1 U12597 ( .A1(n10536), .A2(n10535), .ZN(n9930) );
  NAND2_X1 U12598 ( .A1(n8937), .A2(n11625), .ZN(n9929) );
  NAND2_X1 U12599 ( .A1(n9932), .A2(n9931), .ZN(n9933) );
  NAND2_X1 U12600 ( .A1(n10177), .A2(n9934), .ZN(n9935) );
  NAND2_X1 U12601 ( .A1(n9936), .A2(n9935), .ZN(n10158) );
  XNOR2_X1 U12602 ( .A(n10158), .B(n10152), .ZN(n9940) );
  AOI21_X1 U12603 ( .B1(n9940), .B2(n14814), .A(n9939), .ZN(n14894) );
  MUX2_X1 U12604 ( .A(n9941), .B(n14894), .S(n14515), .Z(n9947) );
  NAND2_X1 U12605 ( .A1(n14865), .A2(n14831), .ZN(n11634) );
  NOR2_X1 U12606 ( .A1(n11634), .A2(n8937), .ZN(n14818) );
  NAND2_X1 U12607 ( .A1(n14818), .A2(n14879), .ZN(n14817) );
  AOI211_X1 U12608 ( .C1(n9942), .C2(n10174), .A(n13169), .B(n10163), .ZN(
        n14892) );
  INV_X1 U12609 ( .A(n9943), .ZN(n14832) );
  OAI22_X1 U12610 ( .A1(n14824), .A2(n14895), .B1(n14819), .B2(n9944), .ZN(
        n9945) );
  AOI21_X1 U12611 ( .B1(n14892), .B2(n14507), .A(n9945), .ZN(n9946) );
  OAI211_X1 U12612 ( .C1(n13178), .C2(n14896), .A(n9947), .B(n9946), .ZN(
        P2_U3260) );
  MUX2_X1 U12613 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12304), .Z(n10347) );
  INV_X1 U12614 ( .A(n10354), .ZN(n10348) );
  XNOR2_X1 U12615 ( .A(n10347), .B(n10348), .ZN(n10345) );
  MUX2_X1 U12616 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n8210), .Z(n9948) );
  INV_X1 U12617 ( .A(n9974), .ZN(n10051) );
  XNOR2_X1 U12618 ( .A(n9948), .B(n10051), .ZN(n10041) );
  INV_X1 U12619 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n10188) );
  MUX2_X1 U12620 ( .A(n10188), .B(n10782), .S(n12304), .Z(n10191) );
  AND2_X1 U12621 ( .A1(n10191), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10200) );
  NAND2_X1 U12622 ( .A1(n10041), .A2(n10200), .ZN(n9951) );
  INV_X1 U12623 ( .A(n9948), .ZN(n9949) );
  NAND2_X1 U12624 ( .A1(n9949), .A2(n10051), .ZN(n9950) );
  NAND2_X1 U12625 ( .A1(n9951), .A2(n9950), .ZN(n10054) );
  MUX2_X1 U12626 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12304), .Z(n9952) );
  XNOR2_X1 U12627 ( .A(n9952), .B(n6431), .ZN(n10055) );
  NAND2_X1 U12628 ( .A1(n10054), .A2(n10055), .ZN(n9955) );
  INV_X1 U12629 ( .A(n9952), .ZN(n9953) );
  NAND2_X1 U12630 ( .A1(n9953), .A2(n6431), .ZN(n9954) );
  NAND2_X1 U12631 ( .A1(n9955), .A2(n9954), .ZN(n10070) );
  MUX2_X1 U12632 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12304), .Z(n9956) );
  XNOR2_X1 U12633 ( .A(n9956), .B(n10082), .ZN(n10071) );
  NAND2_X1 U12634 ( .A1(n10070), .A2(n10071), .ZN(n9959) );
  INV_X1 U12635 ( .A(n9956), .ZN(n9957) );
  NAND2_X1 U12636 ( .A1(n9957), .A2(n10082), .ZN(n9958) );
  NAND2_X1 U12637 ( .A1(n9959), .A2(n9958), .ZN(n10092) );
  MUX2_X1 U12638 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12304), .Z(n9960) );
  XNOR2_X1 U12639 ( .A(n9960), .B(n10108), .ZN(n10093) );
  NAND2_X1 U12640 ( .A1(n10092), .A2(n10093), .ZN(n9963) );
  INV_X1 U12641 ( .A(n9960), .ZN(n9961) );
  NAND2_X1 U12642 ( .A1(n9961), .A2(n10108), .ZN(n9962) );
  MUX2_X1 U12643 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12304), .Z(n9964) );
  XNOR2_X1 U12644 ( .A(n9964), .B(n6695), .ZN(n10021) );
  NAND2_X1 U12645 ( .A1(n10020), .A2(n10021), .ZN(n9967) );
  INV_X1 U12646 ( .A(n9964), .ZN(n9965) );
  NAND2_X1 U12647 ( .A1(n9965), .A2(n6695), .ZN(n9966) );
  NAND2_X1 U12648 ( .A1(n9967), .A2(n9966), .ZN(n10346) );
  XOR2_X1 U12649 ( .A(n10346), .B(n10345), .Z(n10019) );
  NAND2_X1 U12650 ( .A1(n11804), .A2(n9968), .ZN(n9969) );
  AND2_X1 U12651 ( .A1(n6425), .A2(n9969), .ZN(n10010) );
  NAND2_X1 U12652 ( .A1(n9971), .A2(n11851), .ZN(n10011) );
  AND2_X1 U12653 ( .A1(n10010), .A2(n10011), .ZN(n9991) );
  INV_X1 U12654 ( .A(n8211), .ZN(n9972) );
  MUX2_X1 U12655 ( .A(n9991), .B(P3_U3897), .S(n9972), .Z(n15035) );
  INV_X1 U12656 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n12189) );
  NOR2_X1 U12657 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n10188), .ZN(n10193) );
  NAND2_X1 U12658 ( .A1(n9975), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n9973) );
  OAI21_X1 U12659 ( .B1(n9974), .B2(n10193), .A(n9973), .ZN(n10043) );
  INV_X1 U12660 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n15119) );
  NOR2_X1 U12661 ( .A1(n9977), .A2(n10082), .ZN(n9979) );
  INV_X1 U12662 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n9980) );
  OR2_X1 U12663 ( .A1(n10108), .A2(n9980), .ZN(n9983) );
  NAND2_X1 U12664 ( .A1(n10108), .A2(n9980), .ZN(n9981) );
  NAND2_X1 U12665 ( .A1(n9983), .A2(n9981), .ZN(n10097) );
  INV_X1 U12666 ( .A(n10097), .ZN(n9982) );
  INV_X1 U12667 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n10023) );
  NAND2_X1 U12668 ( .A1(n10354), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n10352) );
  OR2_X1 U12669 ( .A1(n10354), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n9985) );
  NAND2_X1 U12670 ( .A1(n10352), .A2(n9985), .ZN(n9987) );
  INV_X1 U12671 ( .A(n10353), .ZN(n9986) );
  AOI21_X1 U12672 ( .B1(n9988), .B2(n9987), .A(n9986), .ZN(n10016) );
  INV_X1 U12673 ( .A(n9989), .ZN(n9990) );
  NAND2_X1 U12674 ( .A1(n9991), .A2(n6717), .ZN(n12367) );
  INV_X1 U12675 ( .A(n10108), .ZN(n9992) );
  NAND2_X1 U12676 ( .A1(n9992), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n10002) );
  MUX2_X1 U12677 ( .A(n9993), .B(P3_REG1_REG_4__SCAN_IN), .S(n10108), .Z(
        n10100) );
  NAND2_X1 U12678 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n9994), .ZN(n10196) );
  INV_X1 U12679 ( .A(n10196), .ZN(n9996) );
  NOR2_X1 U12680 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10196), .ZN(n9995) );
  AOI21_X1 U12681 ( .B1(n9997), .B2(n9996), .A(n10046), .ZN(n10061) );
  MUX2_X1 U12682 ( .A(P3_REG1_REG_2__SCAN_IN), .B(n9998), .S(n6431), .Z(n10062) );
  NAND2_X1 U12683 ( .A1(n9999), .A2(n10000), .ZN(n10001) );
  XNOR2_X1 U12684 ( .A(n10000), .B(n10082), .ZN(n10075) );
  NAND2_X1 U12685 ( .A1(P3_REG1_REG_3__SCAN_IN), .A2(n10075), .ZN(n10074) );
  NAND2_X1 U12686 ( .A1(n10003), .A2(n10004), .ZN(n10005) );
  NAND2_X1 U12687 ( .A1(P3_REG1_REG_5__SCAN_IN), .A2(n10026), .ZN(n10025) );
  NAND2_X1 U12688 ( .A1(n10005), .A2(n10025), .ZN(n10008) );
  MUX2_X1 U12689 ( .A(P3_REG1_REG_6__SCAN_IN), .B(n10006), .S(n10354), .Z(
        n10007) );
  OAI21_X1 U12690 ( .B1(n10008), .B2(n10007), .A(n10355), .ZN(n10009) );
  NAND2_X1 U12691 ( .A1(n15048), .A2(n10009), .ZN(n10015) );
  INV_X1 U12692 ( .A(n10010), .ZN(n10012) );
  INV_X1 U12693 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n10013) );
  NOR2_X1 U12694 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10013), .ZN(n10961) );
  AOI21_X1 U12695 ( .B1(n14998), .B2(P3_ADDR_REG_6__SCAN_IN), .A(n10961), .ZN(
        n10014) );
  OAI211_X1 U12696 ( .C1(n10016), .C2(n15050), .A(n10015), .B(n10014), .ZN(
        n10017) );
  AOI21_X1 U12697 ( .B1(n10348), .B2(n15035), .A(n10017), .ZN(n10018) );
  OAI21_X1 U12698 ( .B1(n10019), .B2(n15042), .A(n10018), .ZN(P3_U3188) );
  XOR2_X1 U12699 ( .A(n10021), .B(n10020), .Z(n10033) );
  INV_X1 U12700 ( .A(n15050), .ZN(n12328) );
  XNOR2_X1 U12701 ( .A(n10023), .B(n10022), .ZN(n10024) );
  NAND2_X1 U12702 ( .A1(n12328), .A2(n10024), .ZN(n10030) );
  OAI21_X1 U12703 ( .B1(P3_REG1_REG_5__SCAN_IN), .B2(n10026), .A(n10025), .ZN(
        n10027) );
  NAND2_X1 U12704 ( .A1(n15048), .A2(n10027), .ZN(n10029) );
  AND2_X1 U12705 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10805) );
  AOI21_X1 U12706 ( .B1(n14998), .B2(P3_ADDR_REG_5__SCAN_IN), .A(n10805), .ZN(
        n10028) );
  NAND3_X1 U12707 ( .A1(n10030), .A2(n10029), .A3(n10028), .ZN(n10031) );
  AOI21_X1 U12708 ( .B1(n6695), .B2(n15035), .A(n10031), .ZN(n10032) );
  OAI21_X1 U12709 ( .B1(n10033), .B2(n15042), .A(n10032), .ZN(P3_U3187) );
  INV_X1 U12710 ( .A(n11418), .ZN(n10181) );
  OAI21_X1 U12711 ( .B1(n10035), .B2(n10034), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n10036) );
  MUX2_X1 U12712 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10036), .S(
        P1_IR_REG_16__SCAN_IN), .Z(n10038) );
  AOI22_X1 U12713 ( .A1(n13818), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10039), .ZN(n10040) );
  OAI21_X1 U12714 ( .B1(n10181), .B2(n10724), .A(n10040), .ZN(P1_U3339) );
  XOR2_X1 U12715 ( .A(n10200), .B(n10041), .Z(n10053) );
  AOI21_X1 U12716 ( .B1(n15119), .B2(n10043), .A(n10042), .ZN(n10049) );
  NOR2_X1 U12717 ( .A1(n10044), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10045) );
  OAI21_X1 U12718 ( .B1(n10046), .B2(n10045), .A(n15048), .ZN(n10048) );
  AOI22_X1 U12719 ( .A1(n14998), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10047) );
  OAI211_X1 U12720 ( .C1(n10049), .C2(n15050), .A(n10048), .B(n10047), .ZN(
        n10050) );
  AOI21_X1 U12721 ( .B1(n10051), .B2(n15035), .A(n10050), .ZN(n10052) );
  OAI21_X1 U12722 ( .B1(n15042), .B2(n10053), .A(n10052), .ZN(P3_U3183) );
  XOR2_X1 U12723 ( .A(n10055), .B(n10054), .Z(n10069) );
  AOI21_X1 U12724 ( .B1(n10058), .B2(n10057), .A(n10056), .ZN(n10059) );
  NOR2_X1 U12725 ( .A1(n15050), .A2(n10059), .ZN(n10066) );
  AOI21_X1 U12726 ( .B1(n10062), .B2(n10061), .A(n10060), .ZN(n10064) );
  AOI22_X1 U12727 ( .A1(n14998), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10063) );
  OAI21_X1 U12728 ( .B1(n10064), .B2(n12367), .A(n10063), .ZN(n10065) );
  AOI211_X1 U12729 ( .C1(n15035), .C2(n6431), .A(n10066), .B(n10065), .ZN(
        n10068) );
  OAI21_X1 U12730 ( .B1(n10069), .B2(n15042), .A(n10068), .ZN(P3_U3184) );
  XOR2_X1 U12731 ( .A(n10071), .B(n10070), .Z(n10084) );
  AOI21_X1 U12732 ( .B1(n10073), .B2(n12189), .A(n10072), .ZN(n10080) );
  OAI21_X1 U12733 ( .B1(P3_REG1_REG_3__SCAN_IN), .B2(n10075), .A(n10074), .ZN(
        n10076) );
  NAND2_X1 U12734 ( .A1(n15048), .A2(n10076), .ZN(n10079) );
  INV_X1 U12735 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n10077) );
  NOR2_X1 U12736 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10077), .ZN(n10532) );
  AOI21_X1 U12737 ( .B1(n14998), .B2(P3_ADDR_REG_3__SCAN_IN), .A(n10532), .ZN(
        n10078) );
  OAI211_X1 U12738 ( .C1(n10080), .C2(n15050), .A(n10079), .B(n10078), .ZN(
        n10081) );
  AOI21_X1 U12739 ( .B1(n10082), .B2(n15035), .A(n10081), .ZN(n10083) );
  OAI21_X1 U12740 ( .B1(n10084), .B2(n15042), .A(n10083), .ZN(P3_U3185) );
  AND2_X1 U12741 ( .A1(n10085), .A2(n15093), .ZN(n10086) );
  OR2_X1 U12742 ( .A1(n11819), .A2(n10086), .ZN(n10089) );
  NAND2_X1 U12743 ( .A1(n10087), .A2(n12571), .ZN(n10088) );
  NAND2_X1 U12744 ( .A1(n10089), .A2(n10088), .ZN(n10781) );
  OAI22_X1 U12745 ( .A1(n10785), .A2(n12724), .B1(n15143), .B2(n8274), .ZN(
        n10090) );
  AOI21_X1 U12746 ( .B1(n15143), .B2(n10781), .A(n10090), .ZN(n10091) );
  INV_X1 U12747 ( .A(n10091), .ZN(P3_U3390) );
  XOR2_X1 U12748 ( .A(n10093), .B(n10092), .Z(n10110) );
  INV_X1 U12749 ( .A(n10094), .ZN(n10098) );
  INV_X1 U12750 ( .A(n10095), .ZN(n10096) );
  AOI21_X1 U12751 ( .B1(n10098), .B2(n10097), .A(n10096), .ZN(n10106) );
  OAI21_X1 U12752 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10102) );
  NAND2_X1 U12753 ( .A1(n15048), .A2(n10102), .ZN(n10105) );
  INV_X1 U12754 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n10103) );
  NOR2_X1 U12755 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10103), .ZN(n10749) );
  AOI21_X1 U12756 ( .B1(n14998), .B2(P3_ADDR_REG_4__SCAN_IN), .A(n10749), .ZN(
        n10104) );
  OAI211_X1 U12757 ( .C1(n10106), .C2(n15050), .A(n10105), .B(n10104), .ZN(
        n10107) );
  AOI21_X1 U12758 ( .B1(n10108), .B2(n15035), .A(n10107), .ZN(n10109) );
  OAI21_X1 U12759 ( .B1(n10110), .B2(n15042), .A(n10109), .ZN(P3_U3186) );
  OAI21_X1 U12760 ( .B1(n10112), .B2(n13539), .A(n10111), .ZN(n10113) );
  INV_X1 U12761 ( .A(n10113), .ZN(n14709) );
  INV_X1 U12762 ( .A(n14669), .ZN(n14072) );
  OAI21_X1 U12763 ( .B1(n13470), .B2(n10115), .A(n10114), .ZN(n10118) );
  OAI22_X1 U12764 ( .A1(n7348), .A2(n14020), .B1(n10338), .B2(n14060), .ZN(
        n10117) );
  NOR2_X1 U12765 ( .A1(n14709), .A2(n13957), .ZN(n10116) );
  AOI211_X1 U12766 ( .C1(n14183), .C2(n10118), .A(n10117), .B(n10116), .ZN(
        n14708) );
  MUX2_X1 U12767 ( .A(n9311), .B(n14708), .S(n14047), .Z(n10127) );
  INV_X1 U12768 ( .A(n10119), .ZN(n10122) );
  INV_X1 U12769 ( .A(n10120), .ZN(n10121) );
  AOI211_X1 U12770 ( .C1(n14706), .C2(n10122), .A(n14075), .B(n10121), .ZN(
        n14705) );
  INV_X1 U12771 ( .A(n13887), .ZN(n10123) );
  OAI22_X1 U12772 ( .A1(n14666), .A2(n10124), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14044), .ZN(n10125) );
  AOI21_X1 U12773 ( .B1(n14705), .B2(n14659), .A(n10125), .ZN(n10126) );
  OAI211_X1 U12774 ( .C1(n14709), .C2(n14072), .A(n10127), .B(n10126), .ZN(
        P1_U3290) );
  AOI21_X1 U12775 ( .B1(n10137), .B2(P2_REG2_REG_10__SCAN_IN), .A(n10128), 
        .ZN(n10132) );
  INV_X1 U12776 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10129) );
  MUX2_X1 U12777 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10129), .S(n10308), .Z(
        n10131) );
  INV_X1 U12778 ( .A(n10314), .ZN(n10130) );
  OAI21_X1 U12779 ( .B1(n10132), .B2(n10131), .A(n10130), .ZN(n10143) );
  INV_X1 U12780 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10740) );
  NOR2_X1 U12781 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10740), .ZN(n10133) );
  AOI21_X1 U12782 ( .B1(n14799), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n10133), 
        .ZN(n10134) );
  OAI21_X1 U12783 ( .B1(n10135), .B2(n12878), .A(n10134), .ZN(n10142) );
  INV_X1 U12784 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10138) );
  MUX2_X1 U12785 ( .A(n10138), .B(P2_REG1_REG_11__SCAN_IN), .S(n10308), .Z(
        n10139) );
  AOI211_X1 U12786 ( .C1(n10140), .C2(n10139), .A(n14795), .B(n10305), .ZN(
        n10141) );
  AOI211_X1 U12787 ( .C1(n14800), .C2(n10143), .A(n10142), .B(n10141), .ZN(
        n10144) );
  INV_X1 U12788 ( .A(n10144), .ZN(P2_U3225) );
  XOR2_X1 U12789 ( .A(n10145), .B(n10646), .Z(n10146) );
  XNOR2_X1 U12790 ( .A(n10647), .B(n10146), .ZN(n10151) );
  AOI22_X1 U12791 ( .A1(n12781), .A2(n12862), .B1(n12947), .B2(n12864), .ZN(
        n10250) );
  NAND2_X1 U12792 ( .A1(n12842), .A2(n10253), .ZN(n10148) );
  OAI211_X1 U12793 ( .C1(n10250), .C2(n12783), .A(n10148), .B(n10147), .ZN(
        n10149) );
  AOI21_X1 U12794 ( .B1(n14916), .B2(n14499), .A(n10149), .ZN(n10150) );
  OAI21_X1 U12795 ( .B1(n10151), .B2(n12816), .A(n10150), .ZN(P2_U3193) );
  INV_X1 U12796 ( .A(n10152), .ZN(n10153) );
  NAND2_X1 U12797 ( .A1(n14895), .A2(n10155), .ZN(n10156) );
  XOR2_X1 U12798 ( .A(n10240), .B(n10241), .Z(n14904) );
  NOR2_X1 U12799 ( .A1(n14895), .A2(n12866), .ZN(n10157) );
  NAND2_X1 U12800 ( .A1(n14895), .A2(n12866), .ZN(n10159) );
  INV_X1 U12801 ( .A(n10240), .ZN(n10160) );
  OAI21_X1 U12802 ( .B1(n6612), .B2(n10160), .A(n10447), .ZN(n10162) );
  AOI21_X1 U12803 ( .B1(n10162), .B2(n14814), .A(n10161), .ZN(n14902) );
  MUX2_X1 U12804 ( .A(n9392), .B(n14902), .S(n14515), .Z(n10168) );
  INV_X1 U12805 ( .A(n10163), .ZN(n10164) );
  AOI211_X1 U12806 ( .C1(n14901), .C2(n10164), .A(n13169), .B(n10441), .ZN(
        n14900) );
  OAI22_X1 U12807 ( .A1(n14824), .A2(n10247), .B1(n14819), .B2(n10165), .ZN(
        n10166) );
  AOI21_X1 U12808 ( .B1(n14900), .B2(n14507), .A(n10166), .ZN(n10167) );
  OAI211_X1 U12809 ( .C1(n13178), .C2(n14904), .A(n10168), .B(n10167), .ZN(
        P2_U3259) );
  XNOR2_X1 U12810 ( .A(n10169), .B(n10170), .ZN(n14888) );
  XNOR2_X1 U12811 ( .A(n10171), .B(n10170), .ZN(n10173) );
  AOI21_X1 U12812 ( .B1(n10173), .B2(n14814), .A(n10172), .ZN(n14886) );
  MUX2_X1 U12813 ( .A(n12175), .B(n14886), .S(n14515), .Z(n10179) );
  OAI211_X1 U12814 ( .C1(n6944), .C2(n14887), .A(n14816), .B(n10174), .ZN(
        n14885) );
  OAI22_X1 U12815 ( .A1(n14885), .A2(n14820), .B1(n10175), .B2(n14819), .ZN(
        n10176) );
  AOI21_X1 U12816 ( .B1(n13141), .B2(n10177), .A(n10176), .ZN(n10178) );
  OAI211_X1 U12817 ( .C1(n13178), .C2(n14888), .A(n10179), .B(n10178), .ZN(
        P2_U3261) );
  OAI222_X1 U12818 ( .A1(P2_U3088), .A2(n12874), .B1(n13301), .B2(n10181), 
        .C1(n10180), .C2(n13303), .ZN(P2_U3311) );
  XNOR2_X1 U12819 ( .A(n10183), .B(n10182), .ZN(n10184) );
  NAND3_X1 U12820 ( .A1(n10186), .A2(n10185), .A3(n10184), .ZN(n10187) );
  INV_X1 U12821 ( .A(n15113), .ZN(n10896) );
  OR2_X1 U12822 ( .A1(n10187), .A2(n10896), .ZN(n11406) );
  AOI21_X1 U12823 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(n15098), .A(n10781), .ZN(
        n10189) );
  MUX2_X1 U12824 ( .A(n10189), .B(n10188), .S(n14462), .Z(n10190) );
  OAI21_X1 U12825 ( .B1(n10785), .B2(n12587), .A(n10190), .ZN(P3_U3233) );
  NAND3_X1 U12826 ( .A1(n15050), .A2(n12367), .A3(n15042), .ZN(n10199) );
  NOR2_X1 U12827 ( .A1(n15042), .A2(n10191), .ZN(n10192) );
  MUX2_X1 U12828 ( .A(n10192), .B(n15035), .S(P3_IR_REG_0__SCAN_IN), .Z(n10198) );
  AOI22_X1 U12829 ( .A1(n14998), .A2(P3_ADDR_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(P3_U3151), .ZN(n10195) );
  NAND2_X1 U12830 ( .A1(n12328), .A2(n10193), .ZN(n10194) );
  OAI211_X1 U12831 ( .C1(n10196), .C2(n12367), .A(n10195), .B(n10194), .ZN(
        n10197) );
  AOI211_X1 U12832 ( .C1(n10200), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10201) );
  INV_X1 U12833 ( .A(n10201), .ZN(P3_U3182) );
  NAND3_X1 U12834 ( .A1(n15102), .A2(n11681), .A3(n10202), .ZN(n10203) );
  OAI211_X1 U12835 ( .C1(n10205), .C2(n15103), .A(n10204), .B(n10203), .ZN(
        n10206) );
  NAND2_X1 U12836 ( .A1(n10206), .A2(n6997), .ZN(n10210) );
  OAI22_X1 U12837 ( .A1(n15107), .A2(n12126), .B1(n6670), .B2(n12109), .ZN(
        n10207) );
  AOI21_X1 U12838 ( .B1(n10208), .B2(n12132), .A(n10207), .ZN(n10209) );
  OAI211_X1 U12839 ( .C1(n10438), .C2(n15115), .A(n10210), .B(n10209), .ZN(
        P3_U3162) );
  NAND2_X1 U12840 ( .A1(n10604), .A2(n10338), .ZN(n10211) );
  OR2_X1 U12841 ( .A1(n10213), .A2(n13436), .ZN(n10216) );
  AOI22_X1 U12842 ( .A1(n11515), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11514), 
        .B2(n10214), .ZN(n10215) );
  NAND2_X1 U12843 ( .A1(n10216), .A2(n10215), .ZN(n14713) );
  XNOR2_X1 U12844 ( .A(n14713), .B(n13747), .ZN(n13473) );
  INV_X1 U12845 ( .A(n13473), .ZN(n10217) );
  OAI21_X1 U12846 ( .B1(n10218), .B2(n10217), .A(n10261), .ZN(n10219) );
  INV_X1 U12847 ( .A(n10219), .ZN(n14717) );
  OAI21_X1 U12848 ( .B1(n10221), .B2(n13473), .A(n10281), .ZN(n10233) );
  NAND2_X1 U12849 ( .A1(n11600), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n10230) );
  OR2_X1 U12850 ( .A1(n6467), .A2(n10222), .ZN(n10229) );
  AND2_X1 U12851 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  NOR2_X1 U12852 ( .A1(n10224), .A2(n10223), .ZN(n10271) );
  OR2_X1 U12853 ( .A1(n10225), .A2(n10271), .ZN(n14661) );
  OR2_X1 U12854 ( .A1(n6465), .A2(n14661), .ZN(n10228) );
  OR2_X1 U12855 ( .A1(n6426), .A2(n10226), .ZN(n10227) );
  NAND4_X1 U12856 ( .A1(n10230), .A2(n10229), .A3(n10228), .A4(n10227), .ZN(
        n13746) );
  INV_X1 U12857 ( .A(n13746), .ZN(n10624) );
  OAI22_X1 U12858 ( .A1(n10624), .A2(n14060), .B1(n10338), .B2(n14020), .ZN(
        n10232) );
  NOR2_X1 U12859 ( .A1(n14717), .A2(n13957), .ZN(n10231) );
  AOI211_X1 U12860 ( .C1(n14183), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n14715) );
  MUX2_X1 U12861 ( .A(n9341), .B(n14715), .S(n14047), .Z(n10239) );
  INV_X1 U12862 ( .A(n10234), .ZN(n10236) );
  INV_X1 U12863 ( .A(n14713), .ZN(n10259) );
  NAND2_X1 U12864 ( .A1(n10259), .A2(n10234), .ZN(n10551) );
  INV_X1 U12865 ( .A(n10551), .ZN(n10235) );
  AOI211_X1 U12866 ( .C1(n14713), .C2(n10236), .A(n14075), .B(n10235), .ZN(
        n14711) );
  OAI22_X1 U12867 ( .A1(n14666), .A2(n10259), .B1(n14044), .B2(n10341), .ZN(
        n10237) );
  AOI21_X1 U12868 ( .B1(n14711), .B2(n14659), .A(n10237), .ZN(n10238) );
  OAI211_X1 U12869 ( .C1(n14717), .C2(n14072), .A(n10239), .B(n10238), .ZN(
        P1_U3288) );
  NAND2_X1 U12870 ( .A1(n10241), .A2(n10240), .ZN(n10244) );
  NAND2_X1 U12871 ( .A1(n10247), .A2(n10242), .ZN(n10243) );
  INV_X1 U12872 ( .A(n10246), .ZN(n10468) );
  OAI21_X1 U12873 ( .B1(n6610), .B2(n10246), .A(n10464), .ZN(n14918) );
  NOR2_X1 U12874 ( .A1(n10247), .A2(n12865), .ZN(n10445) );
  NOR2_X1 U12875 ( .A1(n10448), .A2(n10445), .ZN(n10248) );
  NAND2_X1 U12876 ( .A1(n10450), .A2(n10249), .ZN(n10469) );
  XNOR2_X1 U12877 ( .A(n10469), .B(n10468), .ZN(n10251) );
  OAI21_X1 U12878 ( .B1(n10251), .B2(n14834), .A(n10250), .ZN(n14920) );
  NAND2_X1 U12879 ( .A1(n14920), .A2(n14515), .ZN(n10257) );
  INV_X1 U12880 ( .A(n10252), .ZN(n10440) );
  AOI211_X1 U12881 ( .C1(n14916), .C2(n10440), .A(n13169), .B(n10479), .ZN(
        n14915) );
  AOI22_X1 U12882 ( .A1(n14844), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n10253), 
        .B2(n14839), .ZN(n10254) );
  OAI21_X1 U12883 ( .B1(n10470), .B2(n14824), .A(n10254), .ZN(n10255) );
  AOI21_X1 U12884 ( .B1(n14915), .B2(n14507), .A(n10255), .ZN(n10256) );
  OAI211_X1 U12885 ( .C1(n13178), .C2(n14918), .A(n10257), .B(n10256), .ZN(
        P2_U3257) );
  AND2_X1 U12886 ( .A1(n13957), .A2(n13459), .ZN(n10258) );
  INV_X1 U12887 ( .A(n13747), .ZN(n10279) );
  NAND2_X1 U12888 ( .A1(n10259), .A2(n10279), .ZN(n10260) );
  AOI22_X1 U12889 ( .A1(n11515), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11514), 
        .B2(n10263), .ZN(n10264) );
  XNOR2_X1 U12890 ( .A(n13556), .B(n13746), .ZN(n13474) );
  OR2_X1 U12891 ( .A1(n13556), .A2(n13746), .ZN(n10266) );
  OR2_X1 U12892 ( .A1(n10267), .A2(n13436), .ZN(n10270) );
  AOI22_X1 U12893 ( .A1(n11515), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11514), 
        .B2(n10268), .ZN(n10269) );
  NAND2_X1 U12894 ( .A1(n10270), .A2(n10269), .ZN(n13563) );
  NAND2_X1 U12895 ( .A1(n11600), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n10277) );
  OR2_X1 U12896 ( .A1(n6467), .A2(n9343), .ZN(n10276) );
  NAND2_X1 U12897 ( .A1(n10271), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10287) );
  OR2_X1 U12898 ( .A1(n10271), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U12899 ( .A1(n10287), .A2(n10272), .ZN(n10717) );
  OR2_X1 U12900 ( .A1(n6465), .A2(n10717), .ZN(n10275) );
  OR2_X1 U12901 ( .A1(n6426), .A2(n10273), .ZN(n10274) );
  NAND4_X1 U12902 ( .A1(n10277), .A2(n10276), .A3(n10275), .A4(n10274), .ZN(
        n13745) );
  XNOR2_X1 U12903 ( .A(n13563), .B(n13745), .ZN(n13476) );
  INV_X1 U12904 ( .A(n13476), .ZN(n10284) );
  OAI21_X1 U12905 ( .B1(n10278), .B2(n10284), .A(n10486), .ZN(n10371) );
  INV_X1 U12906 ( .A(n10371), .ZN(n10302) );
  NAND2_X1 U12907 ( .A1(n14713), .A2(n10279), .ZN(n10280) );
  INV_X1 U12908 ( .A(n13556), .ZN(n14667) );
  NAND2_X1 U12909 ( .A1(n14667), .A2(n13746), .ZN(n10282) );
  NAND2_X1 U12910 ( .A1(n13556), .A2(n10624), .ZN(n10283) );
  XNOR2_X1 U12911 ( .A(n10507), .B(n10284), .ZN(n10295) );
  NAND2_X1 U12912 ( .A1(n11600), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10293) );
  OR2_X1 U12913 ( .A1(n6467), .A2(n10285), .ZN(n10292) );
  NAND2_X1 U12914 ( .A1(n10287), .A2(n10286), .ZN(n10288) );
  NAND2_X1 U12915 ( .A1(n10496), .A2(n10288), .ZN(n14648) );
  OR2_X1 U12916 ( .A1(n6465), .A2(n14648), .ZN(n10291) );
  OR2_X1 U12917 ( .A1(n6426), .A2(n10289), .ZN(n10290) );
  NAND4_X1 U12918 ( .A1(n10293), .A2(n10292), .A3(n10291), .A4(n10290), .ZN(
        n13744) );
  INV_X1 U12919 ( .A(n13744), .ZN(n10508) );
  OAI22_X1 U12920 ( .A1(n10508), .A2(n14060), .B1(n10624), .B2(n14020), .ZN(
        n10720) );
  INV_X1 U12921 ( .A(n10720), .ZN(n10294) );
  OAI21_X1 U12922 ( .B1(n10295), .B2(n14166), .A(n10294), .ZN(n10369) );
  INV_X1 U12923 ( .A(n10369), .ZN(n10296) );
  MUX2_X1 U12924 ( .A(n9343), .B(n10296), .S(n14047), .Z(n10301) );
  INV_X1 U12925 ( .A(n13563), .ZN(n10723) );
  INV_X1 U12926 ( .A(n10567), .ZN(n10297) );
  AOI211_X1 U12927 ( .C1(n13563), .C2(n10298), .A(n14075), .B(n10297), .ZN(
        n10370) );
  OAI22_X1 U12928 ( .A1(n10723), .A2(n14666), .B1(n14044), .B2(n10717), .ZN(
        n10299) );
  AOI21_X1 U12929 ( .B1(n10370), .B2(n14659), .A(n10299), .ZN(n10300) );
  OAI211_X1 U12930 ( .C1(n14091), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        P1_U3286) );
  INV_X1 U12931 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14531) );
  NOR2_X1 U12932 ( .A1(n10304), .A2(n14531), .ZN(n10303) );
  AOI21_X1 U12933 ( .B1(n14531), .B2(n10304), .A(n10303), .ZN(n10307) );
  OAI21_X1 U12934 ( .B1(n10307), .B2(n10306), .A(n10692), .ZN(n10319) );
  NOR2_X1 U12935 ( .A1(n10308), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n10313) );
  INV_X1 U12936 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10309) );
  OR2_X1 U12937 ( .A1(n10696), .A2(n10309), .ZN(n10311) );
  NAND2_X1 U12938 ( .A1(n10696), .A2(n10309), .ZN(n10310) );
  NAND2_X1 U12939 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  OR3_X1 U12940 ( .A1(n10314), .A2(n10313), .A3(n10312), .ZN(n10315) );
  AOI21_X1 U12941 ( .B1(n10695), .B2(n10315), .A(n14786), .ZN(n10318) );
  INV_X1 U12942 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n14601) );
  NAND2_X1 U12943 ( .A1(n14805), .A2(n10696), .ZN(n10316) );
  NAND2_X1 U12944 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11009)
         );
  OAI211_X1 U12945 ( .C1(n14601), .C2(n14793), .A(n10316), .B(n11009), .ZN(
        n10317) );
  AOI211_X1 U12946 ( .C1(n10319), .C2(n14765), .A(n10318), .B(n10317), .ZN(
        n10320) );
  INV_X1 U12947 ( .A(n10320), .ZN(P2_U3226) );
  AOI22_X1 U12948 ( .A1(n13548), .A2(n11967), .B1(n11930), .B2(n13748), .ZN(
        n10326) );
  OAI22_X1 U12949 ( .A1(n10604), .A2(n10324), .B1(n10338), .B2(n11979), .ZN(
        n10325) );
  XOR2_X1 U12950 ( .A(n11853), .B(n10325), .Z(n10408) );
  NAND2_X1 U12951 ( .A1(n14713), .A2(n11966), .ZN(n10329) );
  NAND2_X1 U12952 ( .A1(n13747), .A2(n11967), .ZN(n10328) );
  NAND2_X1 U12953 ( .A1(n10329), .A2(n10328), .ZN(n10330) );
  XNOR2_X1 U12954 ( .A(n10330), .B(n11853), .ZN(n10334) );
  NAND2_X1 U12955 ( .A1(n14713), .A2(n11967), .ZN(n10332) );
  NAND2_X1 U12956 ( .A1(n11930), .A2(n13747), .ZN(n10331) );
  NAND2_X1 U12957 ( .A1(n10332), .A2(n10331), .ZN(n10333) );
  NOR2_X1 U12958 ( .A1(n10334), .A2(n10333), .ZN(n10619) );
  NAND2_X1 U12959 ( .A1(n10334), .A2(n10333), .ZN(n10622) );
  INV_X1 U12960 ( .A(n10622), .ZN(n10335) );
  NOR2_X1 U12961 ( .A1(n10619), .A2(n10335), .ZN(n10336) );
  XNOR2_X1 U12962 ( .A(n10621), .B(n10336), .ZN(n10344) );
  OAI21_X1 U12963 ( .B1(n14562), .B2(n10338), .A(n10337), .ZN(n10339) );
  AOI21_X1 U12964 ( .B1(n13418), .B2(n13746), .A(n10339), .ZN(n10340) );
  OAI21_X1 U12965 ( .B1(n10341), .B2(n14580), .A(n10340), .ZN(n10342) );
  AOI21_X1 U12966 ( .B1(n14576), .B2(n14713), .A(n10342), .ZN(n10343) );
  OAI21_X1 U12967 ( .B1(n10344), .B2(n14570), .A(n10343), .ZN(P1_U3227) );
  MUX2_X1 U12968 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12304), .Z(n10383) );
  XNOR2_X1 U12969 ( .A(n10383), .B(n10396), .ZN(n10381) );
  NAND2_X1 U12970 ( .A1(n10346), .A2(n10345), .ZN(n10351) );
  INV_X1 U12971 ( .A(n10347), .ZN(n10349) );
  NAND2_X1 U12972 ( .A1(n10349), .A2(n10348), .ZN(n10350) );
  NAND2_X1 U12973 ( .A1(n10351), .A2(n10350), .ZN(n10382) );
  XOR2_X1 U12974 ( .A(n10381), .B(n10382), .Z(n10364) );
  INV_X1 U12975 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15060) );
  XNOR2_X1 U12976 ( .A(n15060), .B(n10397), .ZN(n10362) );
  INV_X1 U12977 ( .A(n15035), .ZN(n15002) );
  NAND2_X1 U12978 ( .A1(n10354), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n10356) );
  XNOR2_X1 U12979 ( .A(n10387), .B(n10396), .ZN(n10357) );
  NAND2_X1 U12980 ( .A1(P3_REG1_REG_7__SCAN_IN), .A2(n10357), .ZN(n10389) );
  OAI21_X1 U12981 ( .B1(P3_REG1_REG_7__SCAN_IN), .B2(n10357), .A(n10389), .ZN(
        n10358) );
  NAND2_X1 U12982 ( .A1(n10358), .A2(n15048), .ZN(n10360) );
  AND2_X1 U12983 ( .A1(P3_U3151), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n11109) );
  AOI21_X1 U12984 ( .B1(n14998), .B2(P3_ADDR_REG_7__SCAN_IN), .A(n11109), .ZN(
        n10359) );
  OAI211_X1 U12985 ( .C1(n15002), .C2(n10388), .A(n10360), .B(n10359), .ZN(
        n10361) );
  AOI21_X1 U12986 ( .B1(n10362), .B2(n12328), .A(n10361), .ZN(n10363) );
  OAI21_X1 U12987 ( .B1(n10364), .B2(n15042), .A(n10363), .ZN(P3_U3189) );
  INV_X1 U12988 ( .A(n10365), .ZN(n10367) );
  OAI222_X1 U12989 ( .A1(P3_U3151), .A2(n10368), .B1(n12747), .B2(n10367), 
        .C1(n10366), .C2(n12726), .ZN(P3_U3275) );
  AOI211_X1 U12990 ( .C1(n14725), .C2(n10371), .A(n10370), .B(n10369), .ZN(
        n10376) );
  AOI22_X1 U12991 ( .A1(n13563), .A2(n10857), .B1(n14732), .B2(
        P1_REG1_REG_7__SCAN_IN), .ZN(n10372) );
  OAI21_X1 U12992 ( .B1(n10376), .B2(n14732), .A(n10372), .ZN(P1_U3535) );
  INV_X1 U12993 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10373) );
  OAI22_X1 U12994 ( .A1(n10723), .A2(n14227), .B1(n14729), .B2(n10373), .ZN(
        n10374) );
  INV_X1 U12995 ( .A(n10374), .ZN(n10375) );
  OAI21_X1 U12996 ( .B1(n10376), .B2(n14727), .A(n10375), .ZN(P1_U3480) );
  INV_X1 U12997 ( .A(n11424), .ZN(n10379) );
  XNOR2_X1 U12998 ( .A(n10378), .B(P1_IR_REG_17__SCAN_IN), .ZN(n13833) );
  INV_X1 U12999 ( .A(n13833), .ZN(n13830) );
  OAI222_X1 U13000 ( .A1(n14252), .A2(n7040), .B1(n10724), .B2(n10379), .C1(
        n13830), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U13001 ( .A(n14804), .ZN(n12876) );
  OAI222_X1 U13002 ( .A1(n13303), .A2(n10380), .B1(n13301), .B2(n10379), .C1(
        n12876), .C2(P2_U3088), .ZN(P2_U3310) );
  MUX2_X1 U13003 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12304), .Z(n10661) );
  INV_X1 U13004 ( .A(n10666), .ZN(n10662) );
  XNOR2_X1 U13005 ( .A(n10661), .B(n10662), .ZN(n10659) );
  NAND2_X1 U13006 ( .A1(n10382), .A2(n10381), .ZN(n10386) );
  INV_X1 U13007 ( .A(n10383), .ZN(n10384) );
  NAND2_X1 U13008 ( .A1(n10384), .A2(n10396), .ZN(n10385) );
  NAND2_X1 U13009 ( .A1(n10386), .A2(n10385), .ZN(n10660) );
  XOR2_X1 U13010 ( .A(n10659), .B(n10660), .Z(n10406) );
  NAND2_X1 U13011 ( .A1(n10388), .A2(n10387), .ZN(n10390) );
  MUX2_X1 U13012 ( .A(P3_REG1_REG_8__SCAN_IN), .B(n10391), .S(n10666), .Z(
        n10392) );
  OAI21_X1 U13013 ( .B1(n10393), .B2(n10392), .A(n10667), .ZN(n10404) );
  NOR2_X1 U13014 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12217), .ZN(n12034) );
  AOI21_X1 U13015 ( .B1(n14998), .B2(P3_ADDR_REG_8__SCAN_IN), .A(n12034), .ZN(
        n10394) );
  OAI21_X1 U13016 ( .B1(n15002), .B2(n10666), .A(n10394), .ZN(n10403) );
  NAND2_X1 U13017 ( .A1(n10666), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10671) );
  OR2_X1 U13018 ( .A1(n10666), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U13019 ( .A1(n10671), .A2(n10398), .ZN(n10399) );
  NAND2_X1 U13020 ( .A1(n10400), .A2(n10399), .ZN(n10401) );
  AOI21_X1 U13021 ( .B1(n10672), .B2(n10401), .A(n15050), .ZN(n10402) );
  AOI211_X1 U13022 ( .C1(n15048), .C2(n10404), .A(n10403), .B(n10402), .ZN(
        n10405) );
  OAI21_X1 U13023 ( .B1(n10406), .B2(n15042), .A(n10405), .ZN(P3_U3190) );
  XOR2_X1 U13024 ( .A(n10408), .B(n10407), .Z(n10409) );
  NAND2_X1 U13025 ( .A1(n10409), .A2(n14553), .ZN(n10414) );
  NAND2_X1 U13026 ( .A1(n13332), .A2(n10607), .ZN(n10411) );
  NAND2_X1 U13027 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  AOI21_X1 U13028 ( .B1(n14576), .B2(n13548), .A(n10412), .ZN(n10413) );
  OAI211_X1 U13029 ( .C1(n14580), .C2(n10606), .A(n10414), .B(n10413), .ZN(
        P1_U3230) );
  INV_X1 U13030 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n11081) );
  XNOR2_X1 U13031 ( .A(n11221), .B(n11081), .ZN(n10417) );
  OAI21_X1 U13032 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10930), .A(n10415), 
        .ZN(n13795) );
  INV_X1 U13033 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10940) );
  MUX2_X1 U13034 ( .A(n10940), .B(P1_REG1_REG_13__SCAN_IN), .S(n13802), .Z(
        n13794) );
  NOR2_X1 U13035 ( .A1(n13795), .A2(n13794), .ZN(n13793) );
  NAND2_X1 U13036 ( .A1(n10417), .A2(n10416), .ZN(n10990) );
  OAI21_X1 U13037 ( .B1(n10417), .B2(n10416), .A(n10990), .ZN(n10428) );
  XNOR2_X1 U13038 ( .A(n10998), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n10423) );
  INV_X1 U13039 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n10420) );
  MUX2_X1 U13040 ( .A(P1_REG2_REG_13__SCAN_IN), .B(n10420), .S(n13802), .Z(
        n13800) );
  NOR2_X1 U13041 ( .A1(n10930), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n10418) );
  NOR2_X1 U13042 ( .A1(n10419), .A2(n10418), .ZN(n13801) );
  NAND2_X1 U13043 ( .A1(n13800), .A2(n13801), .ZN(n13799) );
  OAI21_X1 U13044 ( .B1(n10421), .B2(n10420), .A(n13799), .ZN(n10422) );
  NAND2_X1 U13045 ( .A1(n10423), .A2(n10422), .ZN(n10997) );
  OAI211_X1 U13046 ( .C1(n10423), .C2(n10422), .A(n14641), .B(n10997), .ZN(
        n10426) );
  NAND2_X1 U13047 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n14547)
         );
  INV_X1 U13048 ( .A(n14547), .ZN(n10424) );
  AOI21_X1 U13049 ( .B1(n14627), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n10424), 
        .ZN(n10425) );
  OAI211_X1 U13050 ( .C1(n13807), .C2(n10998), .A(n10426), .B(n10425), .ZN(
        n10427) );
  AOI21_X1 U13051 ( .B1(n14640), .B2(n10428), .A(n10427), .ZN(n10429) );
  INV_X1 U13052 ( .A(n10429), .ZN(P1_U3257) );
  OAI21_X1 U13053 ( .B1(n10431), .B2(n10430), .A(n10527), .ZN(n10432) );
  NAND2_X1 U13054 ( .A1(n10432), .A2(n6997), .ZN(n10436) );
  OAI22_X1 U13055 ( .A1(n15088), .A2(n12126), .B1(n15087), .B2(n12109), .ZN(
        n10433) );
  AOI21_X1 U13056 ( .B1(n10434), .B2(n12132), .A(n10433), .ZN(n10435) );
  OAI211_X1 U13057 ( .C1(n10438), .C2(n10437), .A(n10436), .B(n10435), .ZN(
        P3_U3177) );
  XNOR2_X1 U13058 ( .A(n10439), .B(n10448), .ZN(n14912) );
  OAI211_X1 U13059 ( .C1(n14909), .C2(n10441), .A(n10440), .B(n14816), .ZN(
        n14908) );
  AOI22_X1 U13060 ( .A1(n13141), .A2(n10443), .B1(n14839), .B2(n10442), .ZN(
        n10444) );
  OAI21_X1 U13061 ( .B1(n14908), .B2(n14820), .A(n10444), .ZN(n10455) );
  INV_X1 U13062 ( .A(n10445), .ZN(n10446) );
  NAND2_X1 U13063 ( .A1(n10447), .A2(n10446), .ZN(n10449) );
  NAND2_X1 U13064 ( .A1(n10449), .A2(n10448), .ZN(n10451) );
  NAND3_X1 U13065 ( .A1(n10451), .A2(n14814), .A3(n10450), .ZN(n10453) );
  NAND2_X1 U13066 ( .A1(n10453), .A2(n10452), .ZN(n14910) );
  MUX2_X1 U13067 ( .A(n14910), .B(P2_REG2_REG_7__SCAN_IN), .S(n14844), .Z(
        n10454) );
  AOI211_X1 U13068 ( .C1(n14828), .C2(n14912), .A(n10455), .B(n10454), .ZN(
        n10456) );
  INV_X1 U13069 ( .A(n10456), .ZN(P2_U3258) );
  INV_X1 U13070 ( .A(n11507), .ZN(n10462) );
  INV_X1 U13071 ( .A(n12891), .ZN(n12895) );
  OAI222_X1 U13072 ( .A1(n13303), .A2(n10457), .B1(n13301), .B2(n10462), .C1(
        P2_U3088), .C2(n12895), .ZN(P2_U3309) );
  NAND2_X1 U13073 ( .A1(n10458), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10459) );
  MUX2_X1 U13074 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10459), .S(
        P1_IR_REG_18__SCAN_IN), .Z(n10461) );
  AND2_X1 U13075 ( .A1(n10461), .A2(n10460), .ZN(n13847) );
  INV_X1 U13076 ( .A(n13847), .ZN(n13841) );
  OAI222_X1 U13077 ( .A1(n14252), .A2(n7037), .B1(n10724), .B2(n10462), .C1(
        P1_U3086), .C2(n13841), .ZN(P1_U3337) );
  OR2_X1 U13078 ( .A1(n10470), .A2(n10475), .ZN(n10463) );
  NAND2_X1 U13079 ( .A1(n10464), .A2(n10463), .ZN(n10466) );
  INV_X1 U13080 ( .A(n10465), .ZN(n10473) );
  NAND2_X1 U13081 ( .A1(n10466), .A2(n10473), .ZN(n10584) );
  OR2_X1 U13082 ( .A1(n10466), .A2(n10473), .ZN(n10467) );
  NAND2_X1 U13083 ( .A1(n10584), .A2(n10467), .ZN(n14926) );
  NAND2_X1 U13084 ( .A1(n10469), .A2(n10468), .ZN(n10472) );
  NAND2_X1 U13085 ( .A1(n10470), .A2(n12863), .ZN(n10471) );
  XNOR2_X1 U13086 ( .A(n10577), .B(n10473), .ZN(n10474) );
  NAND2_X1 U13087 ( .A1(n10474), .A2(n14814), .ZN(n10478) );
  OR2_X1 U13088 ( .A1(n10475), .A2(n12843), .ZN(n10476) );
  OAI21_X1 U13089 ( .B1(n12913), .B2(n10736), .A(n10476), .ZN(n10477) );
  INV_X1 U13090 ( .A(n10477), .ZN(n10644) );
  NAND2_X1 U13091 ( .A1(n10478), .A2(n10644), .ZN(n14928) );
  NAND2_X1 U13092 ( .A1(n14928), .A2(n14515), .ZN(n10484) );
  OAI211_X1 U13093 ( .C1(n10479), .C2(n14923), .A(n14816), .B(n10587), .ZN(
        n14925) );
  INV_X1 U13094 ( .A(n14925), .ZN(n10482) );
  AOI22_X1 U13095 ( .A1(n14844), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n10641), 
        .B2(n14839), .ZN(n10480) );
  OAI21_X1 U13096 ( .B1(n14923), .B2(n14824), .A(n10480), .ZN(n10481) );
  AOI21_X1 U13097 ( .B1(n10482), .B2(n14507), .A(n10481), .ZN(n10483) );
  OAI211_X1 U13098 ( .C1(n13178), .C2(n14926), .A(n10484), .B(n10483), .ZN(
        P2_U3256) );
  OR2_X1 U13099 ( .A1(n13563), .A2(n13745), .ZN(n10485) );
  NAND2_X1 U13100 ( .A1(n10486), .A2(n10485), .ZN(n10565) );
  OR2_X1 U13101 ( .A1(n10487), .A2(n13436), .ZN(n10490) );
  AOI22_X1 U13102 ( .A1(n11515), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11514), 
        .B2(n10488), .ZN(n10489) );
  XNOR2_X1 U13103 ( .A(n13572), .B(n10508), .ZN(n13478) );
  OR2_X1 U13104 ( .A1(n13572), .A2(n13744), .ZN(n10491) );
  OR2_X1 U13105 ( .A1(n10492), .A2(n13436), .ZN(n10495) );
  AOI22_X1 U13106 ( .A1(n11515), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11514), 
        .B2(n10493), .ZN(n10494) );
  NAND2_X1 U13107 ( .A1(n11600), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10502) );
  OR2_X1 U13108 ( .A1(n6467), .A2(n9604), .ZN(n10501) );
  AND2_X1 U13109 ( .A1(n10496), .A2(n11044), .ZN(n10497) );
  OR2_X1 U13110 ( .A1(n10497), .A2(n10828), .ZN(n11043) );
  OR2_X1 U13111 ( .A1(n6465), .A2(n11043), .ZN(n10500) );
  OR2_X1 U13112 ( .A1(n6426), .A2(n10498), .ZN(n10499) );
  NAND4_X1 U13113 ( .A1(n10502), .A2(n10501), .A3(n10500), .A4(n10499), .ZN(
        n13743) );
  XNOR2_X1 U13114 ( .A(n13576), .B(n13743), .ZN(n13479) );
  OAI21_X1 U13115 ( .B1(n10503), .B2(n10511), .A(n10845), .ZN(n14726) );
  INV_X1 U13116 ( .A(n14726), .ZN(n10525) );
  OAI22_X1 U13117 ( .A1(n14047), .A2(n9604), .B1(n11043), .B2(n14044), .ZN(
        n10506) );
  INV_X1 U13118 ( .A(n13576), .ZN(n10504) );
  NAND2_X1 U13119 ( .A1(n10504), .A2(n10566), .ZN(n10825) );
  OAI211_X1 U13120 ( .C1(n10504), .C2(n10566), .A(n14163), .B(n10825), .ZN(
        n14722) );
  INV_X1 U13121 ( .A(n14659), .ZN(n13975) );
  NOR2_X1 U13122 ( .A1(n14722), .A2(n13975), .ZN(n10505) );
  AOI211_X1 U13123 ( .C1(n13994), .C2(n13576), .A(n10506), .B(n10505), .ZN(
        n10524) );
  INV_X1 U13124 ( .A(n13745), .ZN(n10712) );
  OR2_X1 U13125 ( .A1(n13572), .A2(n10508), .ZN(n10509) );
  NAND2_X1 U13126 ( .A1(n10512), .A2(n10511), .ZN(n10513) );
  AOI21_X1 U13127 ( .B1(n10840), .B2(n10513), .A(n14166), .ZN(n14723) );
  NAND2_X1 U13128 ( .A1(n6688), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10519) );
  XNOR2_X1 U13129 ( .A(n10828), .B(P1_REG3_REG_10__SCAN_IN), .ZN(n14561) );
  OR2_X1 U13130 ( .A1(n6465), .A2(n14561), .ZN(n10518) );
  OR2_X1 U13131 ( .A1(n6426), .A2(n10514), .ZN(n10517) );
  INV_X1 U13132 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10515) );
  OR2_X1 U13133 ( .A1(n6428), .A2(n10515), .ZN(n10516) );
  NAND4_X1 U13134 ( .A1(n10519), .A2(n10518), .A3(n10517), .A4(n10516), .ZN(
        n13742) );
  NAND2_X1 U13135 ( .A1(n13742), .A2(n14083), .ZN(n10521) );
  NAND2_X1 U13136 ( .A1(n13744), .A2(n14085), .ZN(n10520) );
  AND2_X1 U13137 ( .A1(n10521), .A2(n10520), .ZN(n14721) );
  INV_X1 U13138 ( .A(n14721), .ZN(n10522) );
  OAI21_X1 U13139 ( .B1(n14723), .B2(n10522), .A(n14047), .ZN(n10523) );
  OAI211_X1 U13140 ( .C1(n10525), .C2(n14091), .A(n10524), .B(n10523), .ZN(
        P1_U3284) );
  AND2_X1 U13141 ( .A1(n10527), .A2(n10526), .ZN(n10530) );
  OAI211_X1 U13142 ( .C1(n10530), .C2(n10529), .A(n6997), .B(n10528), .ZN(
        n10534) );
  OAI22_X1 U13143 ( .A1(n12114), .A2(n10892), .B1(n10685), .B2(n12109), .ZN(
        n10531) );
  AOI211_X1 U13144 ( .C1(n12107), .C2(n12283), .A(n10532), .B(n10531), .ZN(
        n10533) );
  OAI211_X1 U13145 ( .C1(P3_REG3_REG_3__SCAN_IN), .C2(n12130), .A(n10534), .B(
        n10533), .ZN(P3_U3158) );
  XNOR2_X1 U13146 ( .A(n10536), .B(n10535), .ZN(n10538) );
  AOI21_X1 U13147 ( .B1(n10538), .B2(n14814), .A(n10537), .ZN(n14873) );
  XNOR2_X1 U13148 ( .A(n10540), .B(n10539), .ZN(n14876) );
  NAND2_X1 U13149 ( .A1(n11634), .A2(n8937), .ZN(n10541) );
  NAND2_X1 U13150 ( .A1(n10541), .A2(n14816), .ZN(n10542) );
  NOR2_X1 U13151 ( .A1(n14818), .A2(n10542), .ZN(n14870) );
  AOI22_X1 U13152 ( .A1(n14507), .A2(n14870), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n14839), .ZN(n10544) );
  NAND2_X1 U13153 ( .A1(n14844), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n10543) );
  OAI211_X1 U13154 ( .C1(n10545), .C2(n14824), .A(n10544), .B(n10543), .ZN(
        n10546) );
  AOI21_X1 U13155 ( .B1(n14876), .B2(n14828), .A(n10546), .ZN(n10547) );
  OAI21_X1 U13156 ( .B1(n14844), .B2(n14873), .A(n10547), .ZN(P2_U3263) );
  INV_X1 U13157 ( .A(n14716), .ZN(n14385) );
  OAI21_X1 U13158 ( .B1(n10549), .B2(n10554), .A(n10548), .ZN(n14670) );
  AOI211_X1 U13159 ( .C1(n13556), .C2(n10551), .A(n14075), .B(n10550), .ZN(
        n14660) );
  NAND2_X1 U13160 ( .A1(n13745), .A2(n14083), .ZN(n10553) );
  NAND2_X1 U13161 ( .A1(n13747), .A2(n14085), .ZN(n10552) );
  NAND2_X1 U13162 ( .A1(n10553), .A2(n10552), .ZN(n10630) );
  XNOR2_X1 U13163 ( .A(n10555), .B(n10554), .ZN(n10556) );
  NOR2_X1 U13164 ( .A1(n10556), .A2(n14166), .ZN(n10557) );
  AOI211_X1 U13165 ( .C1(n6436), .C2(n14670), .A(n10630), .B(n10557), .ZN(
        n14672) );
  INV_X1 U13166 ( .A(n14672), .ZN(n10558) );
  AOI211_X1 U13167 ( .C1(n14385), .C2(n14670), .A(n14660), .B(n10558), .ZN(
        n10563) );
  AOI22_X1 U13168 ( .A1(n10857), .A2(n13556), .B1(n14732), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n10559) );
  OAI21_X1 U13169 ( .B1(n10563), .B2(n14732), .A(n10559), .ZN(P1_U3534) );
  INV_X1 U13170 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10560) );
  OAI22_X1 U13171 ( .A1(n14667), .A2(n14227), .B1(n14729), .B2(n10560), .ZN(
        n10561) );
  INV_X1 U13172 ( .A(n10561), .ZN(n10562) );
  OAI21_X1 U13173 ( .B1(n10563), .B2(n14727), .A(n10562), .ZN(P1_U3477) );
  OAI21_X1 U13174 ( .B1(n10565), .B2(n13478), .A(n10564), .ZN(n14656) );
  AOI211_X1 U13175 ( .C1(n13572), .C2(n10567), .A(n14075), .B(n10566), .ZN(
        n14647) );
  XOR2_X1 U13176 ( .A(n13478), .B(n10568), .Z(n10569) );
  INV_X1 U13177 ( .A(n13743), .ZN(n10838) );
  OAI22_X1 U13178 ( .A1(n10838), .A2(n14060), .B1(n10712), .B2(n14020), .ZN(
        n10816) );
  AOI21_X1 U13179 ( .B1(n10569), .B2(n14183), .A(n10816), .ZN(n14658) );
  INV_X1 U13180 ( .A(n14658), .ZN(n10570) );
  AOI211_X1 U13181 ( .C1(n14725), .C2(n14656), .A(n14647), .B(n10570), .ZN(
        n10575) );
  AOI22_X1 U13182 ( .A1(n13572), .A2(n10857), .B1(n14732), .B2(
        P1_REG1_REG_8__SCAN_IN), .ZN(n10571) );
  OAI21_X1 U13183 ( .B1(n10575), .B2(n14732), .A(n10571), .ZN(P1_U3536) );
  INV_X1 U13184 ( .A(n13572), .ZN(n14653) );
  INV_X1 U13185 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10572) );
  OAI22_X1 U13186 ( .A1(n14653), .A2(n14227), .B1(n14729), .B2(n10572), .ZN(
        n10573) );
  INV_X1 U13187 ( .A(n10573), .ZN(n10574) );
  OAI21_X1 U13188 ( .B1(n10575), .B2(n14727), .A(n10574), .ZN(P1_U3483) );
  AND2_X1 U13189 ( .A1(n14923), .A2(n12862), .ZN(n10576) );
  OAI22_X1 U13190 ( .A1(n10577), .A2(n10576), .B1(n14923), .B2(n12862), .ZN(
        n10579) );
  AOI21_X1 U13191 ( .B1(n10579), .B2(n10585), .A(n14834), .ZN(n10581) );
  OR2_X1 U13192 ( .A1(n10582), .A2(n12843), .ZN(n10580) );
  OAI21_X1 U13193 ( .B1(n12913), .B2(n11112), .A(n10580), .ZN(n10786) );
  AOI21_X1 U13194 ( .B1(n10581), .B2(n10880), .A(n10786), .ZN(n14932) );
  OR2_X1 U13195 ( .A1(n14923), .A2(n10582), .ZN(n10583) );
  NAND2_X1 U13196 ( .A1(n10584), .A2(n10583), .ZN(n10586) );
  NAND2_X1 U13197 ( .A1(n10586), .A2(n10585), .ZN(n10877) );
  OAI21_X1 U13198 ( .B1(n10586), .B2(n10585), .A(n10877), .ZN(n14935) );
  INV_X1 U13199 ( .A(n14935), .ZN(n10593) );
  INV_X1 U13200 ( .A(n10587), .ZN(n10588) );
  OAI211_X1 U13201 ( .C1(n10588), .C2(n14934), .A(n14816), .B(n10885), .ZN(
        n14931) );
  AOI22_X1 U13202 ( .A1(n14844), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n10589), 
        .B2(n14839), .ZN(n10591) );
  NAND2_X1 U13203 ( .A1(n10875), .A2(n13141), .ZN(n10590) );
  OAI211_X1 U13204 ( .C1(n14931), .C2(n14820), .A(n10591), .B(n10590), .ZN(
        n10592) );
  AOI21_X1 U13205 ( .B1(n10593), .B2(n14828), .A(n10592), .ZN(n10594) );
  OAI21_X1 U13206 ( .B1(n14932), .B2(n14844), .A(n10594), .ZN(P2_U3255) );
  AOI22_X1 U13207 ( .A1(n10595), .A2(n14659), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n14662), .ZN(n10596) );
  OAI21_X1 U13208 ( .B1(n10597), .B2(n14666), .A(n10596), .ZN(n10600) );
  MUX2_X1 U13209 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10598), .S(n14047), .Z(
        n10599) );
  AOI211_X1 U13210 ( .C1(n14655), .C2(n10601), .A(n10600), .B(n10599), .ZN(
        n10602) );
  INV_X1 U13211 ( .A(n10602), .ZN(P1_U3291) );
  INV_X1 U13212 ( .A(n10603), .ZN(n10605) );
  OAI22_X1 U13213 ( .A1(n10605), .A2(n13975), .B1(n10604), .B2(n14666), .ZN(
        n10612) );
  NOR2_X1 U13214 ( .A1(n14044), .A2(n10606), .ZN(n10608) );
  OR3_X1 U13215 ( .A1(n10609), .A2(n10608), .A3(n10607), .ZN(n10610) );
  MUX2_X1 U13216 ( .A(n10610), .B(P1_REG2_REG_4__SCAN_IN), .S(n14673), .Z(
        n10611) );
  AOI211_X1 U13217 ( .C1(n14655), .C2(n10613), .A(n10612), .B(n10611), .ZN(
        n10614) );
  INV_X1 U13218 ( .A(n10614), .ZN(P1_U3289) );
  INV_X1 U13219 ( .A(n10615), .ZN(n10618) );
  OAI222_X1 U13220 ( .A1(n12747), .A2(n10618), .B1(n12744), .B2(n10617), .C1(
        P3_U3151), .C2(n10616), .ZN(P3_U3274) );
  INV_X1 U13221 ( .A(n10619), .ZN(n10620) );
  OAI22_X1 U13222 ( .A1(n14667), .A2(n10324), .B1(n10624), .B2(n11979), .ZN(
        n10625) );
  XNOR2_X1 U13223 ( .A(n10625), .B(n11853), .ZN(n10707) );
  AND2_X1 U13224 ( .A1(n11930), .A2(n13746), .ZN(n10626) );
  AOI21_X1 U13225 ( .B1(n13556), .B2(n11932), .A(n10626), .ZN(n10708) );
  XNOR2_X1 U13226 ( .A(n10707), .B(n10708), .ZN(n10627) );
  OAI211_X1 U13227 ( .C1(n10628), .C2(n10627), .A(n10711), .B(n14553), .ZN(
        n10634) );
  AOI21_X1 U13228 ( .B1(n13332), .B2(n10630), .A(n10629), .ZN(n10631) );
  OAI21_X1 U13229 ( .B1(n14580), .B2(n14661), .A(n10631), .ZN(n10632) );
  INV_X1 U13230 ( .A(n10632), .ZN(n10633) );
  OAI211_X1 U13231 ( .C1(n14667), .C2(n13434), .A(n10634), .B(n10633), .ZN(
        P1_U3239) );
  NOR2_X1 U13232 ( .A1(n14650), .A2(n14166), .ZN(n13896) );
  NOR2_X1 U13233 ( .A1(n13896), .A2(n14655), .ZN(n10640) );
  NOR2_X1 U13234 ( .A1(n13975), .A2(n14075), .ZN(n14051) );
  OAI21_X1 U13235 ( .B1(n14051), .B2(n13994), .A(n6434), .ZN(n10639) );
  OAI22_X1 U13236 ( .A1(n14650), .A2(n10636), .B1(n10635), .B2(n14044), .ZN(
        n10637) );
  AOI21_X1 U13237 ( .B1(P1_REG2_REG_0__SCAN_IN), .B2(n14650), .A(n10637), .ZN(
        n10638) );
  OAI211_X1 U13238 ( .C1(n10640), .C2(n13524), .A(n10639), .B(n10638), .ZN(
        P1_U3293) );
  NAND2_X1 U13239 ( .A1(n12842), .A2(n10641), .ZN(n10643) );
  OAI211_X1 U13240 ( .C1(n10644), .C2(n12783), .A(n10643), .B(n10642), .ZN(
        n10652) );
  NAND2_X1 U13241 ( .A1(n14494), .A2(n14833), .ZN(n12837) );
  INV_X1 U13242 ( .A(n12837), .ZN(n12822) );
  NAND3_X1 U13243 ( .A1(n10645), .A2(n12822), .A3(n12863), .ZN(n10650) );
  NAND3_X1 U13244 ( .A1(n10647), .A2(n14494), .A3(n10646), .ZN(n10649) );
  AOI21_X1 U13245 ( .B1(n10650), .B2(n10649), .A(n10648), .ZN(n10651) );
  AOI211_X1 U13246 ( .C1(n10653), .C2(n14499), .A(n10652), .B(n10651), .ZN(
        n10654) );
  OAI21_X1 U13247 ( .B1(n10655), .B2(n12816), .A(n10654), .ZN(P2_U3203) );
  INV_X1 U13248 ( .A(n10656), .ZN(n10658) );
  OAI22_X1 U13249 ( .A1(n11848), .A2(P3_U3151), .B1(SI_22_), .B2(n12726), .ZN(
        n10657) );
  AOI21_X1 U13250 ( .B1(n10658), .B2(n14376), .A(n10657), .ZN(P3_U3273) );
  MUX2_X1 U13251 ( .A(P3_REG2_REG_9__SCAN_IN), .B(P3_REG1_REG_9__SCAN_IN), .S(
        n12304), .Z(n10758) );
  XNOR2_X1 U13252 ( .A(n10758), .B(n10770), .ZN(n10756) );
  NAND2_X1 U13253 ( .A1(n10660), .A2(n10659), .ZN(n10665) );
  INV_X1 U13254 ( .A(n10661), .ZN(n10663) );
  NAND2_X1 U13255 ( .A1(n10663), .A2(n10662), .ZN(n10664) );
  NAND2_X1 U13256 ( .A1(n10665), .A2(n10664), .ZN(n10757) );
  XOR2_X1 U13257 ( .A(n10756), .B(n10757), .Z(n10680) );
  NAND2_X1 U13258 ( .A1(n10666), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U13259 ( .A1(P3_REG1_REG_9__SCAN_IN), .A2(n10669), .ZN(n10764) );
  OAI21_X1 U13260 ( .B1(P3_REG1_REG_9__SCAN_IN), .B2(n10669), .A(n10764), .ZN(
        n10678) );
  AND2_X1 U13261 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11071) );
  AOI21_X1 U13262 ( .B1(n14998), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n11071), .ZN(
        n10670) );
  OAI21_X1 U13263 ( .B1(n15002), .B2(n10763), .A(n10670), .ZN(n10677) );
  INV_X1 U13264 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10673) );
  NOR2_X1 U13265 ( .A1(n10673), .A2(n10674), .ZN(n10771) );
  AOI21_X1 U13266 ( .B1(n10674), .B2(n10673), .A(n10771), .ZN(n10675) );
  NOR2_X1 U13267 ( .A1(n10675), .A2(n15050), .ZN(n10676) );
  AOI211_X1 U13268 ( .C1(n15048), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10679) );
  OAI21_X1 U13269 ( .B1(n10680), .B2(n15042), .A(n10679), .ZN(P3_U3191) );
  OAI21_X1 U13270 ( .B1(n10682), .B2(n11815), .A(n10681), .ZN(n10683) );
  INV_X1 U13271 ( .A(n10683), .ZN(n15077) );
  AOI21_X1 U13272 ( .B1(n10684), .B2(n11815), .A(n15093), .ZN(n10688) );
  OAI22_X1 U13273 ( .A1(n6670), .A2(n15106), .B1(n10685), .B2(n15104), .ZN(
        n10686) );
  AOI21_X1 U13274 ( .B1(n10688), .B2(n10687), .A(n10686), .ZN(n15075) );
  OAI21_X1 U13275 ( .B1(n15077), .B2(n15139), .A(n15075), .ZN(n10894) );
  OAI22_X1 U13276 ( .A1(n10892), .A2(n12724), .B1(n15143), .B2(n8304), .ZN(
        n10689) );
  AOI21_X1 U13277 ( .B1(n10894), .B2(n15143), .A(n10689), .ZN(n10690) );
  INV_X1 U13278 ( .A(n10690), .ZN(P3_U3399) );
  INV_X1 U13279 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n11157) );
  NOR2_X1 U13280 ( .A1(n10868), .A2(n11157), .ZN(n10691) );
  AOI21_X1 U13281 ( .B1(n11157), .B2(n10868), .A(n10691), .ZN(n10694) );
  OAI21_X1 U13282 ( .B1(n10696), .B2(P2_REG1_REG_12__SCAN_IN), .A(n10692), 
        .ZN(n10693) );
  NOR2_X1 U13283 ( .A1(n10693), .A2(n10694), .ZN(n10867) );
  AOI211_X1 U13284 ( .C1(n10694), .C2(n10693), .A(n14795), .B(n10867), .ZN(
        n10706) );
  INV_X1 U13285 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10698) );
  MUX2_X1 U13286 ( .A(n10698), .B(P2_REG2_REG_13__SCAN_IN), .S(n10868), .Z(
        n10700) );
  OAI21_X1 U13287 ( .B1(n10696), .B2(P2_REG2_REG_12__SCAN_IN), .A(n10695), 
        .ZN(n10699) );
  AND2_X1 U13288 ( .A1(n10868), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10697) );
  AOI211_X1 U13289 ( .C1(n10700), .C2(n10699), .A(n14786), .B(n10863), .ZN(
        n10705) );
  NOR2_X1 U13290 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10970), .ZN(n10701) );
  AOI21_X1 U13291 ( .B1(n14799), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n10701), 
        .ZN(n10702) );
  OAI21_X1 U13292 ( .B1(n10703), .B2(n12878), .A(n10702), .ZN(n10704) );
  OR3_X1 U13293 ( .A1(n10706), .A2(n10705), .A3(n10704), .ZN(P2_U3227) );
  INV_X1 U13294 ( .A(n10708), .ZN(n10709) );
  OAI22_X1 U13295 ( .A1(n10723), .A2(n10324), .B1(n10712), .B2(n11979), .ZN(
        n10713) );
  XNOR2_X1 U13296 ( .A(n10713), .B(n11853), .ZN(n10809) );
  AND2_X1 U13297 ( .A1(n11930), .A2(n13745), .ZN(n10714) );
  AOI21_X1 U13298 ( .B1(n13563), .B2(n11932), .A(n10714), .ZN(n10810) );
  XNOR2_X1 U13299 ( .A(n10809), .B(n10810), .ZN(n10715) );
  OAI211_X1 U13300 ( .C1(n10716), .C2(n10715), .A(n10813), .B(n14553), .ZN(
        n10722) );
  NOR2_X1 U13301 ( .A1(n14580), .A2(n10717), .ZN(n10718) );
  AOI211_X1 U13302 ( .C1(n13332), .C2(n10720), .A(n10719), .B(n10718), .ZN(
        n10721) );
  OAI211_X1 U13303 ( .C1(n10723), .C2(n13434), .A(n10722), .B(n10721), .ZN(
        P1_U3213) );
  INV_X1 U13304 ( .A(n11512), .ZN(n10754) );
  OAI222_X1 U13305 ( .A1(n14252), .A2(n10725), .B1(n10724), .B2(n10754), .C1(
        n13920), .C2(P1_U3086), .ZN(P1_U3336) );
  OAI21_X1 U13306 ( .B1(n10727), .B2(n11817), .A(n10726), .ZN(n10902) );
  OAI211_X1 U13307 ( .C1(n10729), .C2(n11696), .A(n10728), .B(n15109), .ZN(
        n10731) );
  AOI22_X1 U13308 ( .A1(n12148), .A2(n12571), .B1(n12569), .B2(n12149), .ZN(
        n10730) );
  NAND2_X1 U13309 ( .A1(n10731), .A2(n10730), .ZN(n10899) );
  AOI21_X1 U13310 ( .B1(n14482), .B2(n10902), .A(n10899), .ZN(n10862) );
  OAI22_X1 U13311 ( .A1(n11703), .A2(n12724), .B1(n15143), .B2(n8322), .ZN(
        n10732) );
  INV_X1 U13312 ( .A(n10732), .ZN(n10733) );
  OAI21_X1 U13313 ( .B1(n10862), .B2(n15144), .A(n10733), .ZN(P3_U3402) );
  INV_X1 U13314 ( .A(n10734), .ZN(n10735) );
  AOI21_X1 U13315 ( .B1(n10735), .B2(n10790), .A(n12816), .ZN(n10739) );
  NOR3_X1 U13316 ( .A1(n10737), .A2(n10736), .A3(n12837), .ZN(n10738) );
  OAI21_X1 U13317 ( .B1(n10739), .B2(n10738), .A(n11011), .ZN(n10743) );
  AOI22_X1 U13318 ( .A1(n12781), .A2(n12859), .B1(n12947), .B2(n12861), .ZN(
        n10883) );
  OAI22_X1 U13319 ( .A1(n12783), .A2(n10883), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10740), .ZN(n10741) );
  AOI21_X1 U13320 ( .B1(n7446), .B2(n12842), .A(n10741), .ZN(n10742) );
  OAI211_X1 U13321 ( .C1(n6956), .C2(n12846), .A(n10743), .B(n10742), .ZN(
        P2_U3208) );
  AOI21_X1 U13322 ( .B1(n10746), .B2(n10745), .A(n6455), .ZN(n10753) );
  OAI22_X1 U13323 ( .A1(n12114), .A2(n11703), .B1(n10747), .B2(n12109), .ZN(
        n10748) );
  AOI211_X1 U13324 ( .C1(n12107), .C2(n12149), .A(n10749), .B(n10748), .ZN(
        n10752) );
  INV_X1 U13325 ( .A(n10898), .ZN(n10750) );
  NAND2_X1 U13326 ( .A1(n12117), .A2(n10750), .ZN(n10751) );
  OAI211_X1 U13327 ( .C1(n10753), .C2(n12134), .A(n10752), .B(n10751), .ZN(
        P3_U3170) );
  OAI222_X1 U13328 ( .A1(n13303), .A2(n10755), .B1(P2_U3088), .B2(n13001), 
        .C1(n13301), .C2(n10754), .ZN(P2_U3308) );
  MUX2_X1 U13329 ( .A(P3_REG2_REG_10__SCAN_IN), .B(P3_REG1_REG_10__SCAN_IN), 
        .S(n12304), .Z(n12288) );
  XNOR2_X1 U13330 ( .A(n12288), .B(n12332), .ZN(n12286) );
  NAND2_X1 U13331 ( .A1(n10757), .A2(n10756), .ZN(n10761) );
  INV_X1 U13332 ( .A(n10758), .ZN(n10759) );
  NAND2_X1 U13333 ( .A1(n10759), .A2(n10770), .ZN(n10760) );
  XOR2_X1 U13334 ( .A(n12286), .B(n12287), .Z(n10780) );
  AOI22_X1 U13335 ( .A1(n12332), .A2(n8404), .B1(P3_REG1_REG_10__SCAN_IN), 
        .B2(n12314), .ZN(n10767) );
  NAND2_X1 U13336 ( .A1(n10763), .A2(n10762), .ZN(n10765) );
  NAND2_X1 U13337 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  OAI21_X1 U13338 ( .B1(n10767), .B2(n10766), .A(n12331), .ZN(n10778) );
  AND2_X1 U13339 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n11025) );
  AOI21_X1 U13340 ( .B1(n14998), .B2(P3_ADDR_REG_10__SCAN_IN), .A(n11025), 
        .ZN(n10768) );
  OAI21_X1 U13341 ( .B1(n15002), .B2(n12314), .A(n10768), .ZN(n10777) );
  NOR2_X1 U13342 ( .A1(n10770), .A2(n10769), .ZN(n10772) );
  INV_X1 U13343 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n12613) );
  AOI22_X1 U13344 ( .A1(n12332), .A2(P3_REG2_REG_10__SCAN_IN), .B1(n12613), 
        .B2(n12314), .ZN(n10773) );
  AOI21_X1 U13345 ( .B1(n10774), .B2(n10773), .A(n12313), .ZN(n10775) );
  NOR2_X1 U13346 ( .A1(n10775), .A2(n15050), .ZN(n10776) );
  AOI211_X1 U13347 ( .C1(n15048), .C2(n10778), .A(n10777), .B(n10776), .ZN(
        n10779) );
  OAI21_X1 U13348 ( .B1(n10780), .B2(n15042), .A(n10779), .ZN(P3_U3192) );
  INV_X1 U13349 ( .A(n10781), .ZN(n10783) );
  MUX2_X1 U13350 ( .A(n10783), .B(n10782), .S(n15150), .Z(n10784) );
  OAI21_X1 U13351 ( .B1(n10785), .B2(n12682), .A(n10784), .ZN(P3_U3459) );
  NAND2_X1 U13352 ( .A1(n14496), .A2(n10786), .ZN(n10788) );
  OAI211_X1 U13353 ( .C1(n14502), .C2(n10789), .A(n10788), .B(n10787), .ZN(
        n10795) );
  INV_X1 U13354 ( .A(n10790), .ZN(n10791) );
  AOI211_X1 U13355 ( .C1(n10793), .C2(n10792), .A(n12816), .B(n10791), .ZN(
        n10794) );
  AOI211_X1 U13356 ( .C1(n10875), .C2(n14499), .A(n10795), .B(n10794), .ZN(
        n10796) );
  INV_X1 U13357 ( .A(n10796), .ZN(P2_U3189) );
  NAND2_X1 U13358 ( .A1(n10797), .A2(n14376), .ZN(n10798) );
  OAI211_X1 U13359 ( .C1(n10799), .C2(n12726), .A(n10798), .B(n11851), .ZN(
        P3_U3272) );
  OAI21_X1 U13360 ( .B1(n10801), .B2(n10800), .A(n10956), .ZN(n10802) );
  NAND2_X1 U13361 ( .A1(n10802), .A2(n6997), .ZN(n10807) );
  OAI22_X1 U13362 ( .A1(n12114), .A2(n10984), .B1(n10803), .B2(n12109), .ZN(
        n10804) );
  AOI211_X1 U13363 ( .C1(n12107), .C2(n11704), .A(n10805), .B(n10804), .ZN(
        n10806) );
  OAI211_X1 U13364 ( .C1(n15074), .C2(n12130), .A(n10807), .B(n10806), .ZN(
        P3_U3167) );
  AOI22_X1 U13365 ( .A1(n13572), .A2(n11966), .B1(n11932), .B2(n13744), .ZN(
        n10808) );
  XNOR2_X1 U13366 ( .A(n10808), .B(n11853), .ZN(n11034) );
  AOI22_X1 U13367 ( .A1(n13572), .A2(n11932), .B1(n11930), .B2(n13744), .ZN(
        n11033) );
  XNOR2_X1 U13368 ( .A(n11034), .B(n11033), .ZN(n10815) );
  NAND2_X1 U13369 ( .A1(n10809), .A2(n10811), .ZN(n10812) );
  AOI21_X1 U13370 ( .B1(n10815), .B2(n10814), .A(n11036), .ZN(n10820) );
  AOI22_X1 U13371 ( .A1(n10816), .A2(n13332), .B1(P1_REG3_REG_8__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10817) );
  OAI21_X1 U13372 ( .B1(n14580), .B2(n14648), .A(n10817), .ZN(n10818) );
  AOI21_X1 U13373 ( .B1(n13572), .B2(n14576), .A(n10818), .ZN(n10819) );
  OAI21_X1 U13374 ( .B1(n10820), .B2(n14570), .A(n10819), .ZN(P1_U3221) );
  OR2_X1 U13375 ( .A1(n10821), .A2(n13436), .ZN(n10824) );
  AOI22_X1 U13376 ( .A1(n11515), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11514), 
        .B2(n10822), .ZN(n10823) );
  NAND2_X1 U13377 ( .A1(n10825), .A2(n14559), .ZN(n10826) );
  NAND3_X1 U13378 ( .A1(n10920), .A2(n14163), .A3(n10826), .ZN(n10837) );
  NAND2_X1 U13379 ( .A1(n11600), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n10834) );
  OR2_X1 U13380 ( .A1(n6467), .A2(n9816), .ZN(n10833) );
  AND2_X1 U13381 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_10__SCAN_IN), 
        .ZN(n10827) );
  AOI21_X1 U13382 ( .B1(n10828), .B2(P1_REG3_REG_10__SCAN_IN), .A(
        P1_REG3_REG_11__SCAN_IN), .ZN(n10829) );
  OR2_X1 U13383 ( .A1(n10904), .A2(n10829), .ZN(n14579) );
  OR2_X1 U13384 ( .A1(n6465), .A2(n14579), .ZN(n10832) );
  OR2_X1 U13385 ( .A1(n6426), .A2(n10830), .ZN(n10831) );
  NAND4_X1 U13386 ( .A1(n10834), .A2(n10833), .A3(n10832), .A4(n10831), .ZN(
        n13741) );
  NAND2_X1 U13387 ( .A1(n13741), .A2(n14083), .ZN(n10836) );
  NAND2_X1 U13388 ( .A1(n13743), .A2(n14085), .ZN(n10835) );
  AND2_X1 U13389 ( .A1(n10836), .A2(n10835), .ZN(n14551) );
  NAND2_X1 U13390 ( .A1(n10837), .A2(n14551), .ZN(n10852) );
  NOR2_X1 U13391 ( .A1(n14044), .A2(n14561), .ZN(n10843) );
  XNOR2_X1 U13392 ( .A(n14559), .B(n13742), .ZN(n13480) );
  NAND2_X1 U13393 ( .A1(n13576), .A2(n10838), .ZN(n10839) );
  INV_X1 U13394 ( .A(n10911), .ZN(n10841) );
  AOI211_X1 U13395 ( .C1(n10846), .C2(n10842), .A(n14166), .B(n10841), .ZN(
        n10851) );
  AOI211_X1 U13396 ( .C1(n13920), .C2(n10852), .A(n10843), .B(n10851), .ZN(
        n10850) );
  AOI22_X1 U13397 ( .A1(n14559), .A2(n13994), .B1(P1_REG2_REG_10__SCAN_IN), 
        .B2(n14650), .ZN(n10849) );
  OR2_X1 U13398 ( .A1(n13576), .A2(n13743), .ZN(n10844) );
  OAI21_X1 U13399 ( .B1(n10847), .B2(n10846), .A(n10918), .ZN(n10853) );
  NAND2_X1 U13400 ( .A1(n10853), .A2(n14655), .ZN(n10848) );
  OAI211_X1 U13401 ( .C1(n10850), .C2(n14673), .A(n10849), .B(n10848), .ZN(
        P1_U3283) );
  AOI211_X1 U13402 ( .C1(n14725), .C2(n10853), .A(n10852), .B(n10851), .ZN(
        n10859) );
  INV_X1 U13403 ( .A(n14559), .ZN(n10854) );
  OAI22_X1 U13404 ( .A1(n10854), .A2(n14227), .B1(n14729), .B2(n10515), .ZN(
        n10855) );
  INV_X1 U13405 ( .A(n10855), .ZN(n10856) );
  OAI21_X1 U13406 ( .B1(n10859), .B2(n14727), .A(n10856), .ZN(P1_U3489) );
  AOI22_X1 U13407 ( .A1(n14559), .A2(n10857), .B1(n14732), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n10858) );
  OAI21_X1 U13408 ( .B1(n10859), .B2(n14732), .A(n10858), .ZN(P1_U3538) );
  OAI22_X1 U13409 ( .A1(n12682), .A2(n11703), .B1(n15149), .B2(n9993), .ZN(
        n10860) );
  INV_X1 U13410 ( .A(n10860), .ZN(n10861) );
  OAI21_X1 U13411 ( .B1(n10862), .B2(n15150), .A(n10861), .ZN(P3_U3463) );
  AOI21_X1 U13412 ( .B1(P2_REG2_REG_13__SCAN_IN), .B2(n10868), .A(n10863), 
        .ZN(n11189) );
  XNOR2_X1 U13413 ( .A(n11189), .B(n11188), .ZN(n11190) );
  XNOR2_X1 U13414 ( .A(n11190), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n10873) );
  NAND2_X1 U13415 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14500)
         );
  INV_X1 U13416 ( .A(n14500), .ZN(n10864) );
  AOI21_X1 U13417 ( .B1(n14799), .B2(P2_ADDR_REG_14__SCAN_IN), .A(n10864), 
        .ZN(n10865) );
  OAI21_X1 U13418 ( .B1(n11188), .B2(n12878), .A(n10865), .ZN(n10872) );
  INV_X1 U13419 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n14525) );
  NOR2_X1 U13420 ( .A1(n11185), .A2(n14525), .ZN(n10866) );
  AOI21_X1 U13421 ( .B1(n11185), .B2(n14525), .A(n10866), .ZN(n10870) );
  AOI211_X1 U13422 ( .C1(n10870), .C2(n10869), .A(n14795), .B(n11184), .ZN(
        n10871) );
  AOI211_X1 U13423 ( .C1(n14800), .C2(n10873), .A(n10872), .B(n10871), .ZN(
        n10874) );
  INV_X1 U13424 ( .A(n10874), .ZN(P2_U3228) );
  NAND2_X1 U13425 ( .A1(n10875), .A2(n12861), .ZN(n10876) );
  NAND2_X1 U13426 ( .A1(n10877), .A2(n10876), .ZN(n11119) );
  XNOR2_X1 U13427 ( .A(n11119), .B(n10882), .ZN(n14946) );
  AOI21_X1 U13428 ( .B1(n10882), .B2(n10881), .A(n6597), .ZN(n10884) );
  OAI21_X1 U13429 ( .B1(n10884), .B2(n14834), .A(n10883), .ZN(n14940) );
  NAND2_X1 U13430 ( .A1(n14942), .A2(n10885), .ZN(n10886) );
  NAND2_X1 U13431 ( .A1(n10886), .A2(n14816), .ZN(n10887) );
  NOR2_X1 U13432 ( .A1(n6606), .A2(n10887), .ZN(n14941) );
  NAND2_X1 U13433 ( .A1(n14941), .A2(n14507), .ZN(n10889) );
  AOI22_X1 U13434 ( .A1(n14844), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7446), 
        .B2(n14839), .ZN(n10888) );
  OAI211_X1 U13435 ( .C1(n6956), .C2(n14824), .A(n10889), .B(n10888), .ZN(
        n10890) );
  AOI21_X1 U13436 ( .B1(n14940), .B2(n14515), .A(n10890), .ZN(n10891) );
  OAI21_X1 U13437 ( .B1(n13178), .B2(n14946), .A(n10891), .ZN(P2_U3254) );
  OAI22_X1 U13438 ( .A1(n12682), .A2(n10892), .B1(n15149), .B2(n8305), .ZN(
        n10893) );
  AOI21_X1 U13439 ( .B1(n10894), .B2(n15149), .A(n10893), .ZN(n10895) );
  INV_X1 U13440 ( .A(n10895), .ZN(P3_U3462) );
  AND2_X1 U13441 ( .A1(n10896), .A2(n11682), .ZN(n15095) );
  NAND2_X1 U13442 ( .A1(n15120), .A2(n15090), .ZN(n10897) );
  OAI22_X1 U13443 ( .A1(n12587), .A2(n11703), .B1(n10898), .B2(n15114), .ZN(
        n10901) );
  MUX2_X1 U13444 ( .A(n10899), .B(P3_REG2_REG_4__SCAN_IN), .S(n14462), .Z(
        n10900) );
  AOI211_X1 U13445 ( .C1(n12589), .C2(n10902), .A(n10901), .B(n10900), .ZN(
        n10903) );
  INV_X1 U13446 ( .A(n10903), .ZN(P3_U3229) );
  INV_X1 U13447 ( .A(n13742), .ZN(n14563) );
  NAND2_X1 U13448 ( .A1(n11600), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10909) );
  OR2_X1 U13449 ( .A1(n6467), .A2(n9811), .ZN(n10908) );
  OR2_X1 U13450 ( .A1(n10904), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n10905) );
  NAND2_X1 U13451 ( .A1(n10938), .A2(n10905), .ZN(n13344) );
  OR2_X1 U13452 ( .A1(n6465), .A2(n13344), .ZN(n10907) );
  OR2_X1 U13453 ( .A1(n6426), .A2(n14390), .ZN(n10906) );
  NAND4_X1 U13454 ( .A1(n10909), .A2(n10908), .A3(n10907), .A4(n10906), .ZN(
        n13740) );
  OR2_X1 U13455 ( .A1(n14559), .A2(n14563), .ZN(n10910) );
  NAND2_X1 U13456 ( .A1(n10912), .A2(n13461), .ZN(n10915) );
  AOI22_X1 U13457 ( .A1(n11515), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11514), 
        .B2(n10913), .ZN(n10914) );
  XNOR2_X1 U13458 ( .A(n14575), .B(n13741), .ZN(n13482) );
  XNOR2_X1 U13459 ( .A(n10934), .B(n13482), .ZN(n10916) );
  OAI222_X1 U13460 ( .A1(n14020), .A2(n14563), .B1(n14060), .B2(n14564), .C1(
        n10916), .C2(n14166), .ZN(n14589) );
  INV_X1 U13461 ( .A(n14589), .ZN(n10927) );
  OR2_X1 U13462 ( .A1(n14559), .A2(n13742), .ZN(n10917) );
  XOR2_X1 U13463 ( .A(n10928), .B(n13482), .Z(n14591) );
  INV_X1 U13464 ( .A(n14575), .ZN(n14588) );
  NAND2_X1 U13465 ( .A1(n14588), .A2(n10919), .ZN(n10948) );
  AOI21_X1 U13466 ( .B1(n14575), .B2(n10920), .A(n14075), .ZN(n10921) );
  NAND2_X1 U13467 ( .A1(n10948), .A2(n10921), .ZN(n14586) );
  NAND2_X1 U13468 ( .A1(n14673), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10922) );
  OAI21_X1 U13469 ( .B1(n14044), .B2(n14579), .A(n10922), .ZN(n10923) );
  AOI21_X1 U13470 ( .B1(n14575), .B2(n13994), .A(n10923), .ZN(n10924) );
  OAI21_X1 U13471 ( .B1(n14586), .B2(n13975), .A(n10924), .ZN(n10925) );
  AOI21_X1 U13472 ( .B1(n14591), .B2(n14655), .A(n10925), .ZN(n10926) );
  OAI21_X1 U13473 ( .B1(n14650), .B2(n10927), .A(n10926), .ZN(P1_U3282) );
  INV_X1 U13474 ( .A(n13741), .ZN(n13343) );
  NAND2_X1 U13475 ( .A1(n10929), .A2(n13461), .ZN(n10932) );
  AOI22_X1 U13476 ( .A1(n11515), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10930), 
        .B2(n11514), .ZN(n10931) );
  XNOR2_X1 U13477 ( .A(n13601), .B(n14564), .ZN(n13485) );
  XNOR2_X1 U13478 ( .A(n11095), .B(n13485), .ZN(n14386) );
  NAND2_X1 U13479 ( .A1(n14575), .A2(n13343), .ZN(n10933) );
  NAND2_X1 U13480 ( .A1(n10934), .A2(n10933), .ZN(n10936) );
  OR2_X1 U13481 ( .A1(n14575), .A2(n13343), .ZN(n10935) );
  INV_X1 U13482 ( .A(n13485), .ZN(n11087) );
  XNOR2_X1 U13483 ( .A(n11088), .B(n11087), .ZN(n10946) );
  NAND2_X1 U13484 ( .A1(n11600), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10944) );
  OR2_X1 U13485 ( .A1(n6467), .A2(n10420), .ZN(n10943) );
  NAND2_X1 U13486 ( .A1(n10938), .A2(n10937), .ZN(n10939) );
  NAND2_X1 U13487 ( .A1(n11077), .A2(n10939), .ZN(n13393) );
  OR2_X1 U13488 ( .A1(n6465), .A2(n13393), .ZN(n10942) );
  OR2_X1 U13489 ( .A1(n6426), .A2(n10940), .ZN(n10941) );
  NAND4_X1 U13490 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n13739) );
  AOI22_X1 U13491 ( .A1(n14085), .A2(n13741), .B1(n13739), .B2(n14083), .ZN(
        n10945) );
  OAI21_X1 U13492 ( .B1(n10946), .B2(n14166), .A(n10945), .ZN(n10947) );
  AOI21_X1 U13493 ( .B1(n14386), .B2(n6436), .A(n10947), .ZN(n14388) );
  NAND2_X1 U13494 ( .A1(n10948), .A2(n13601), .ZN(n10949) );
  NAND3_X1 U13495 ( .A1(n11097), .A2(n14163), .A3(n10949), .ZN(n14382) );
  OAI22_X1 U13496 ( .A1(n14047), .A2(n9811), .B1(n13344), .B2(n14044), .ZN(
        n10950) );
  AOI21_X1 U13497 ( .B1(n13601), .B2(n13994), .A(n10950), .ZN(n10951) );
  OAI21_X1 U13498 ( .B1(n14382), .B2(n13975), .A(n10951), .ZN(n10952) );
  AOI21_X1 U13499 ( .B1(n14386), .B2(n14669), .A(n10952), .ZN(n10953) );
  OAI21_X1 U13500 ( .B1(n14388), .B2(n14673), .A(n10953), .ZN(P1_U3281) );
  INV_X1 U13501 ( .A(n11526), .ZN(n10975) );
  OAI222_X1 U13502 ( .A1(n14252), .A2(n11527), .B1(n10724), .B2(n10975), .C1(
        n10954), .C2(P1_U3086), .ZN(P1_U3335) );
  AND2_X1 U13503 ( .A1(n10956), .A2(n10955), .ZN(n10959) );
  XNOR2_X1 U13504 ( .A(n10957), .B(n12147), .ZN(n10958) );
  NAND2_X1 U13505 ( .A1(n10959), .A2(n10958), .ZN(n11106) );
  OAI211_X1 U13506 ( .C1(n10959), .C2(n10958), .A(n11106), .B(n6997), .ZN(
        n10963) );
  OAI22_X1 U13507 ( .A1(n12114), .A2(n11062), .B1(n11210), .B2(n12109), .ZN(
        n10960) );
  AOI211_X1 U13508 ( .C1(n12107), .C2(n12148), .A(n10961), .B(n10960), .ZN(
        n10962) );
  OAI211_X1 U13509 ( .C1(n15067), .C2(n12130), .A(n10963), .B(n10962), .ZN(
        P3_U3179) );
  INV_X1 U13510 ( .A(n11152), .ZN(n11141) );
  AOI21_X1 U13511 ( .B1(n10965), .B2(n10964), .A(n12816), .ZN(n10967) );
  NAND2_X1 U13512 ( .A1(n10967), .A2(n10966), .ZN(n10974) );
  NAND2_X1 U13513 ( .A1(n12781), .A2(n12857), .ZN(n10969) );
  OR2_X1 U13514 ( .A1(n11122), .A2(n12843), .ZN(n10968) );
  NAND2_X1 U13515 ( .A1(n10969), .A2(n10968), .ZN(n11134) );
  INV_X1 U13516 ( .A(n11134), .ZN(n10971) );
  OAI22_X1 U13517 ( .A1(n12783), .A2(n10971), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10970), .ZN(n10972) );
  AOI21_X1 U13518 ( .B1(n11139), .B2(n12842), .A(n10972), .ZN(n10973) );
  OAI211_X1 U13519 ( .C1(n11141), .C2(n12846), .A(n10974), .B(n10973), .ZN(
        P2_U3206) );
  OAI222_X1 U13520 ( .A1(n13303), .A2(n10976), .B1(P2_U3088), .B2(n7504), .C1(
        n13301), .C2(n10975), .ZN(P2_U3307) );
  OAI21_X1 U13521 ( .B1(n10978), .B2(n11822), .A(n10977), .ZN(n10979) );
  INV_X1 U13522 ( .A(n10979), .ZN(n15069) );
  OAI21_X1 U13523 ( .B1(n6611), .B2(n11698), .A(n10980), .ZN(n10981) );
  AOI222_X1 U13524 ( .A1(n15109), .A2(n10981), .B1(n12147), .B2(n12571), .C1(
        n11704), .C2(n12569), .ZN(n15068) );
  OAI21_X1 U13525 ( .B1(n15139), .B2(n15069), .A(n15068), .ZN(n10986) );
  OAI22_X1 U13526 ( .A1(n10984), .A2(n12724), .B1(n15143), .B2(n8342), .ZN(
        n10982) );
  AOI21_X1 U13527 ( .B1(n10986), .B2(n15143), .A(n10982), .ZN(n10983) );
  INV_X1 U13528 ( .A(n10983), .ZN(P3_U3405) );
  OAI22_X1 U13529 ( .A1(n12682), .A2(n10984), .B1(n15149), .B2(n8344), .ZN(
        n10985) );
  AOI21_X1 U13530 ( .B1(n10986), .B2(n15149), .A(n10985), .ZN(n10987) );
  INV_X1 U13531 ( .A(n10987), .ZN(P3_U3464) );
  AND2_X1 U13532 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n10988) );
  AOI21_X1 U13533 ( .B1(n14627), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10988), 
        .ZN(n10989) );
  INV_X1 U13534 ( .A(n10989), .ZN(n10996) );
  OAI21_X1 U13535 ( .B1(n11221), .B2(P1_REG1_REG_14__SCAN_IN), .A(n10990), 
        .ZN(n10991) );
  NAND2_X1 U13536 ( .A1(n11000), .A2(n10991), .ZN(n10992) );
  XNOR2_X1 U13537 ( .A(n10991), .B(n14638), .ZN(n14636) );
  INV_X1 U13538 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U13539 ( .A1(n14636), .A2(n14635), .ZN(n14634) );
  NAND2_X1 U13540 ( .A1(n10992), .A2(n14634), .ZN(n10994) );
  XNOR2_X1 U13541 ( .A(n13818), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n10993) );
  NOR2_X1 U13542 ( .A1(n10993), .A2(n10994), .ZN(n13817) );
  AOI211_X1 U13543 ( .C1(n10994), .C2(n10993), .A(n13817), .B(n13819), .ZN(
        n10995) );
  AOI211_X1 U13544 ( .C1(n14637), .C2(n13818), .A(n10996), .B(n10995), .ZN(
        n11006) );
  INV_X1 U13545 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n11080) );
  OAI21_X1 U13546 ( .B1(n11080), .B2(n10998), .A(n10997), .ZN(n10999) );
  NOR2_X1 U13547 ( .A1(n14638), .A2(n10999), .ZN(n11001) );
  XOR2_X1 U13548 ( .A(n11000), .B(n10999), .Z(n14632) );
  NOR2_X1 U13549 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n14632), .ZN(n14631) );
  NOR2_X1 U13550 ( .A1(n11001), .A2(n14631), .ZN(n11004) );
  NOR2_X1 U13551 ( .A1(n13818), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n11002) );
  AOI21_X1 U13552 ( .B1(n13818), .B2(P1_REG2_REG_16__SCAN_IN), .A(n11002), 
        .ZN(n11003) );
  NAND2_X1 U13553 ( .A1(n11003), .A2(n11004), .ZN(n13812) );
  OAI211_X1 U13554 ( .C1(n11004), .C2(n11003), .A(n14641), .B(n13812), .ZN(
        n11005) );
  NAND2_X1 U13555 ( .A1(n11006), .A2(n11005), .ZN(P1_U3259) );
  NAND2_X1 U13556 ( .A1(n12781), .A2(n12858), .ZN(n11008) );
  NAND2_X1 U13557 ( .A1(n12947), .A2(n12860), .ZN(n11007) );
  AND2_X1 U13558 ( .A1(n11008), .A2(n11007), .ZN(n14510) );
  NAND2_X1 U13559 ( .A1(n12842), .A2(n14512), .ZN(n11010) );
  OAI211_X1 U13560 ( .C1(n14510), .C2(n12783), .A(n11010), .B(n11009), .ZN(
        n11018) );
  INV_X1 U13561 ( .A(n11011), .ZN(n11014) );
  NOR3_X1 U13562 ( .A1(n11012), .A2(n11112), .A3(n12837), .ZN(n11013) );
  AOI21_X1 U13563 ( .B1(n11014), .B2(n14494), .A(n11013), .ZN(n11016) );
  NOR2_X1 U13564 ( .A1(n11016), .A2(n11015), .ZN(n11017) );
  AOI211_X1 U13565 ( .C1(n11019), .C2(n14499), .A(n11018), .B(n11017), .ZN(
        n11020) );
  OAI21_X1 U13566 ( .B1(n11021), .B2(n12816), .A(n11020), .ZN(P2_U3196) );
  NAND2_X1 U13567 ( .A1(n11022), .A2(n6997), .ZN(n11032) );
  AOI21_X1 U13568 ( .B1(n11066), .B2(n11024), .A(n11023), .ZN(n11031) );
  NAND2_X1 U13569 ( .A1(n12107), .A2(n12144), .ZN(n11027) );
  INV_X1 U13570 ( .A(n11025), .ZN(n11026) );
  OAI211_X1 U13571 ( .C1(n12611), .C2(n12109), .A(n11027), .B(n11026), .ZN(
        n11029) );
  NOR2_X1 U13572 ( .A1(n12130), .A2(n12612), .ZN(n11028) );
  AOI211_X1 U13573 ( .C1(n12615), .C2(n12132), .A(n11029), .B(n11028), .ZN(
        n11030) );
  OAI21_X1 U13574 ( .B1(n11032), .B2(n11031), .A(n11030), .ZN(P3_U3157) );
  INV_X1 U13575 ( .A(n13422), .ZN(n11049) );
  NAND2_X1 U13576 ( .A1(n13576), .A2(n14712), .ZN(n14720) );
  AND2_X1 U13577 ( .A1(n11034), .A2(n11033), .ZN(n11035) );
  NAND2_X1 U13578 ( .A1(n13576), .A2(n11966), .ZN(n11038) );
  NAND2_X1 U13579 ( .A1(n13743), .A2(n11967), .ZN(n11037) );
  NAND2_X1 U13580 ( .A1(n11038), .A2(n11037), .ZN(n11039) );
  XNOR2_X1 U13581 ( .A(n11039), .B(n11853), .ZN(n11855) );
  AND2_X1 U13582 ( .A1(n11930), .A2(n13743), .ZN(n11040) );
  AOI21_X1 U13583 ( .B1(n13576), .B2(n11932), .A(n11040), .ZN(n11856) );
  XNOR2_X1 U13584 ( .A(n11855), .B(n11856), .ZN(n11041) );
  OAI211_X1 U13585 ( .C1(n11042), .C2(n11041), .A(n11859), .B(n14553), .ZN(
        n11048) );
  INV_X1 U13586 ( .A(n11043), .ZN(n11046) );
  INV_X1 U13587 ( .A(n14580), .ZN(n13430) );
  INV_X1 U13588 ( .A(n13332), .ZN(n14552) );
  OAI22_X1 U13589 ( .A1(n14552), .A2(n14721), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n11044), .ZN(n11045) );
  AOI21_X1 U13590 ( .B1(n11046), .B2(n13430), .A(n11045), .ZN(n11047) );
  OAI211_X1 U13591 ( .C1(n11049), .C2(n14720), .A(n11048), .B(n11047), .ZN(
        P1_U3231) );
  INV_X1 U13592 ( .A(n11539), .ZN(n11995) );
  OAI222_X1 U13593 ( .A1(n13303), .A2(n11051), .B1(n13301), .B2(n11995), .C1(
        n11050), .C2(P2_U3088), .ZN(P2_U3306) );
  OAI21_X1 U13594 ( .B1(n11053), .B2(n11814), .A(n11052), .ZN(n11054) );
  INV_X1 U13595 ( .A(n11054), .ZN(n15062) );
  OAI211_X1 U13596 ( .C1(n11057), .C2(n11056), .A(n11055), .B(n15109), .ZN(
        n11059) );
  AOI22_X1 U13597 ( .A1(n12569), .A2(n12148), .B1(n12146), .B2(n12571), .ZN(
        n11058) );
  AND2_X1 U13598 ( .A1(n11059), .A2(n11058), .ZN(n15061) );
  OAI21_X1 U13599 ( .B1(n15139), .B2(n15062), .A(n15061), .ZN(n11064) );
  OAI22_X1 U13600 ( .A1(n11062), .A2(n12724), .B1(n15143), .B2(n8360), .ZN(
        n11060) );
  AOI21_X1 U13601 ( .B1(n11064), .B2(n15143), .A(n11060), .ZN(n11061) );
  INV_X1 U13602 ( .A(n11061), .ZN(P3_U3408) );
  OAI22_X1 U13603 ( .A1(n12682), .A2(n11062), .B1(n15149), .B2(n10006), .ZN(
        n11063) );
  AOI21_X1 U13604 ( .B1(n11064), .B2(n15149), .A(n11063), .ZN(n11065) );
  INV_X1 U13605 ( .A(n11065), .ZN(P3_U3465) );
  INV_X1 U13606 ( .A(n11066), .ZN(n11067) );
  AOI21_X1 U13607 ( .B1(n11069), .B2(n11068), .A(n11067), .ZN(n11075) );
  OAI22_X1 U13608 ( .A1(n12114), .A2(n11403), .B1(n11398), .B2(n12109), .ZN(
        n11070) );
  AOI211_X1 U13609 ( .C1(n12107), .C2(n12145), .A(n11071), .B(n11070), .ZN(
        n11074) );
  INV_X1 U13610 ( .A(n11404), .ZN(n11072) );
  NAND2_X1 U13611 ( .A1(n12117), .A2(n11072), .ZN(n11073) );
  OAI211_X1 U13612 ( .C1(n11075), .C2(n12134), .A(n11074), .B(n11073), .ZN(
        P3_U3171) );
  INV_X1 U13613 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n11076) );
  NAND2_X1 U13614 ( .A1(n11077), .A2(n11076), .ZN(n11078) );
  NAND2_X1 U13615 ( .A1(n11229), .A2(n11078), .ZN(n14549) );
  INV_X1 U13616 ( .A(n14549), .ZN(n11079) );
  NAND2_X1 U13617 ( .A1(n11545), .A2(n11079), .ZN(n11086) );
  OR2_X1 U13618 ( .A1(n6467), .A2(n11080), .ZN(n11085) );
  OR2_X1 U13619 ( .A1(n6426), .A2(n11081), .ZN(n11084) );
  INV_X1 U13620 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n11082) );
  OR2_X1 U13621 ( .A1(n6428), .A2(n11082), .ZN(n11083) );
  OR2_X1 U13622 ( .A1(n13601), .A2(n14564), .ZN(n11089) );
  NAND2_X1 U13623 ( .A1(n11091), .A2(n13461), .ZN(n11093) );
  AOI22_X1 U13624 ( .A1(n13802), .A2(n11514), .B1(n11515), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n11092) );
  INV_X1 U13625 ( .A(n13739), .ZN(n14536) );
  XNOR2_X1 U13626 ( .A(n13607), .B(n14536), .ZN(n13484) );
  XNOR2_X1 U13627 ( .A(n11219), .B(n6435), .ZN(n11094) );
  OAI222_X1 U13628 ( .A1(n14020), .A2(n14564), .B1(n14060), .B2(n11885), .C1(
        n11094), .C2(n14166), .ZN(n14583) );
  INV_X1 U13629 ( .A(n14583), .ZN(n11104) );
  XNOR2_X1 U13630 ( .A(n11242), .B(n13484), .ZN(n14585) );
  AOI21_X1 U13631 ( .B1(n13607), .B2(n11097), .A(n14075), .ZN(n11098) );
  NAND2_X1 U13632 ( .A1(n11324), .A2(n11098), .ZN(n14581) );
  NAND2_X1 U13633 ( .A1(n14673), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n11099) );
  OAI21_X1 U13634 ( .B1(n14044), .B2(n13393), .A(n11099), .ZN(n11100) );
  AOI21_X1 U13635 ( .B1(n13607), .B2(n13994), .A(n11100), .ZN(n11101) );
  OAI21_X1 U13636 ( .B1(n14581), .B2(n13975), .A(n11101), .ZN(n11102) );
  AOI21_X1 U13637 ( .B1(n14585), .B2(n14655), .A(n11102), .ZN(n11103) );
  OAI21_X1 U13638 ( .B1(n11104), .B2(n14673), .A(n11103), .ZN(P1_U3280) );
  NAND2_X1 U13639 ( .A1(n11106), .A2(n11105), .ZN(n12030) );
  XNOR2_X1 U13640 ( .A(n12030), .B(n12029), .ZN(n11107) );
  NAND2_X1 U13641 ( .A1(n11107), .A2(n6997), .ZN(n11111) );
  OAI22_X1 U13642 ( .A1(n12114), .A2(n11180), .B1(n11399), .B2(n12109), .ZN(
        n11108) );
  AOI211_X1 U13643 ( .C1(n12107), .C2(n12147), .A(n11109), .B(n11108), .ZN(
        n11110) );
  OAI211_X1 U13644 ( .C1(n15054), .C2(n12130), .A(n11111), .B(n11110), .ZN(
        P3_U3153) );
  NAND2_X1 U13645 ( .A1(n14509), .A2(n14508), .ZN(n11114) );
  OR2_X1 U13646 ( .A1(n14527), .A2(n12859), .ZN(n11113) );
  INV_X1 U13647 ( .A(n11125), .ZN(n11271) );
  XNOR2_X1 U13648 ( .A(n11265), .B(n11271), .ZN(n11117) );
  OAI22_X1 U13649 ( .A1(n11364), .A2(n12913), .B1(n11116), .B2(n12843), .ZN(
        n14497) );
  AOI21_X1 U13650 ( .B1(n11117), .B2(n14814), .A(n14497), .ZN(n14521) );
  OR2_X1 U13651 ( .A1(n14942), .A2(n12860), .ZN(n11118) );
  NAND2_X1 U13652 ( .A1(n14942), .A2(n12860), .ZN(n11120) );
  NAND2_X1 U13653 ( .A1(n14527), .A2(n11122), .ZN(n11123) );
  NOR2_X1 U13654 ( .A1(n11152), .A2(n12858), .ZN(n11124) );
  XNOR2_X1 U13655 ( .A(n11272), .B(n11125), .ZN(n14524) );
  OR2_X1 U13656 ( .A1(n11152), .A2(n14505), .ZN(n11126) );
  INV_X1 U13657 ( .A(n11126), .ZN(n11132) );
  AOI211_X1 U13658 ( .C1(n14498), .C2(n11126), .A(n13169), .B(n11276), .ZN(
        n14518) );
  NAND2_X1 U13659 ( .A1(n14518), .A2(n14507), .ZN(n11129) );
  INV_X1 U13660 ( .A(n14503), .ZN(n11127) );
  AOI22_X1 U13661 ( .A1(n14844), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n11127), 
        .B2(n14839), .ZN(n11128) );
  OAI211_X1 U13662 ( .C1(n14520), .C2(n14824), .A(n11129), .B(n11128), .ZN(
        n11130) );
  AOI21_X1 U13663 ( .B1(n14828), .B2(n14524), .A(n11130), .ZN(n11131) );
  OAI21_X1 U13664 ( .B1(n14844), .B2(n14521), .A(n11131), .ZN(P2_U3251) );
  AOI211_X1 U13665 ( .C1(n11152), .C2(n14505), .A(n13169), .B(n11132), .ZN(
        n11151) );
  XOR2_X1 U13666 ( .A(n11138), .B(n11133), .Z(n11135) );
  AOI21_X1 U13667 ( .B1(n11135), .B2(n14814), .A(n11134), .ZN(n11154) );
  INV_X1 U13668 ( .A(n11154), .ZN(n11136) );
  AOI21_X1 U13669 ( .B1(n11151), .B2(n13001), .A(n11136), .ZN(n11145) );
  XOR2_X1 U13670 ( .A(n11138), .B(n11137), .Z(n11155) );
  INV_X1 U13671 ( .A(n11155), .ZN(n11143) );
  AOI22_X1 U13672 ( .A1(n14844), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11139), 
        .B2(n14839), .ZN(n11140) );
  OAI21_X1 U13673 ( .B1(n11141), .B2(n14824), .A(n11140), .ZN(n11142) );
  AOI21_X1 U13674 ( .B1(n11143), .B2(n14828), .A(n11142), .ZN(n11144) );
  OAI21_X1 U13675 ( .B1(n11145), .B2(n14844), .A(n11144), .ZN(P2_U3252) );
  NAND3_X1 U13676 ( .A1(n14854), .A2(n14853), .A3(n11146), .ZN(n11147) );
  INV_X1 U13677 ( .A(n14850), .ZN(n11149) );
  AND2_X1 U13678 ( .A1(n11150), .A2(n6700), .ZN(n14857) );
  INV_X1 U13679 ( .A(n14857), .ZN(n14945) );
  AOI21_X1 U13680 ( .B1(n14943), .B2(n11152), .A(n11151), .ZN(n11153) );
  OAI211_X1 U13681 ( .C1(n13261), .C2(n11155), .A(n11154), .B(n11153), .ZN(
        n11159) );
  NAND2_X1 U13682 ( .A1(n11159), .A2(n14970), .ZN(n11156) );
  OAI21_X1 U13683 ( .B1(n14970), .B2(n11157), .A(n11156), .ZN(P2_U3512) );
  INV_X1 U13684 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U13685 ( .A1(n11159), .A2(n14952), .ZN(n11160) );
  OAI21_X1 U13686 ( .B1(n14952), .B2(n11161), .A(n11160), .ZN(P2_U3469) );
  XNOR2_X1 U13687 ( .A(n12142), .B(n11162), .ZN(n11163) );
  XNOR2_X1 U13688 ( .A(n11164), .B(n11163), .ZN(n11170) );
  INV_X1 U13689 ( .A(n11317), .ZN(n11165) );
  NAND2_X1 U13690 ( .A1(n12117), .A2(n11165), .ZN(n11167) );
  AND2_X1 U13691 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n14979) );
  AOI21_X1 U13692 ( .B1(n12143), .B2(n12107), .A(n14979), .ZN(n11166) );
  OAI211_X1 U13693 ( .C1(n12596), .C2(n12109), .A(n11167), .B(n11166), .ZN(
        n11168) );
  AOI21_X1 U13694 ( .B1(n11316), .B2(n12132), .A(n11168), .ZN(n11169) );
  OAI21_X1 U13695 ( .B1(n11170), .B2(n12134), .A(n11169), .ZN(P3_U3176) );
  OAI21_X1 U13696 ( .B1(n11172), .B2(n11821), .A(n11171), .ZN(n15056) );
  INV_X1 U13697 ( .A(n15056), .ZN(n11177) );
  OAI211_X1 U13698 ( .C1(n11174), .C2(n11711), .A(n11173), .B(n15109), .ZN(
        n11176) );
  AOI22_X1 U13699 ( .A1(n12145), .A2(n12571), .B1(n12569), .B2(n12147), .ZN(
        n11175) );
  AND2_X1 U13700 ( .A1(n11176), .A2(n11175), .ZN(n15053) );
  OAI21_X1 U13701 ( .B1(n15139), .B2(n11177), .A(n15053), .ZN(n11182) );
  OAI22_X1 U13702 ( .A1(n11180), .A2(n12724), .B1(n15143), .B2(n8376), .ZN(
        n11178) );
  AOI21_X1 U13703 ( .B1(n11182), .B2(n15143), .A(n11178), .ZN(n11179) );
  INV_X1 U13704 ( .A(n11179), .ZN(P3_U3411) );
  OAI22_X1 U13705 ( .A1(n12682), .A2(n11180), .B1(n15149), .B2(n8373), .ZN(
        n11181) );
  AOI21_X1 U13706 ( .B1(n11182), .B2(n15149), .A(n11181), .ZN(n11183) );
  INV_X1 U13707 ( .A(n11183), .ZN(P3_U3466) );
  INV_X1 U13708 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n11186) );
  NOR2_X1 U13709 ( .A1(n11186), .A2(n11187), .ZN(n11337) );
  AOI211_X1 U13710 ( .C1(n11187), .C2(n11186), .A(n11337), .B(n14795), .ZN(
        n11200) );
  OR2_X1 U13711 ( .A1(n11189), .A2(n11188), .ZN(n11193) );
  INV_X1 U13712 ( .A(n11190), .ZN(n11191) );
  NAND2_X1 U13713 ( .A1(n11193), .A2(n11192), .ZN(n11341) );
  XNOR2_X1 U13714 ( .A(n11335), .B(n11341), .ZN(n11194) );
  NAND2_X1 U13715 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11194), .ZN(n11343) );
  OAI211_X1 U13716 ( .C1(P2_REG2_REG_15__SCAN_IN), .C2(n11194), .A(n14800), 
        .B(n11343), .ZN(n11198) );
  NOR2_X1 U13717 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n11195), .ZN(n11196) );
  AOI21_X1 U13718 ( .B1(n14799), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n11196), 
        .ZN(n11197) );
  OAI211_X1 U13719 ( .C1(n12878), .C2(n11335), .A(n11198), .B(n11197), .ZN(
        n11199) );
  OR2_X1 U13720 ( .A1(n11200), .A2(n11199), .ZN(P2_U3229) );
  INV_X1 U13721 ( .A(n11201), .ZN(n11203) );
  OAI222_X1 U13722 ( .A1(n13303), .A2(n11204), .B1(n13301), .B2(n11203), .C1(
        n6700), .C2(P2_U3088), .ZN(P2_U3305) );
  INV_X1 U13723 ( .A(n8759), .ZN(n11208) );
  INV_X1 U13724 ( .A(n11205), .ZN(n11206) );
  OAI222_X1 U13725 ( .A1(P3_U3151), .A2(n11208), .B1(n12744), .B2(n11207), 
        .C1(n12747), .C2(n11206), .ZN(P3_U3271) );
  XNOR2_X1 U13726 ( .A(n11395), .B(n11718), .ZN(n15129) );
  INV_X1 U13727 ( .A(n15090), .ZN(n15112) );
  XNOR2_X1 U13728 ( .A(n11209), .B(n11820), .ZN(n11212) );
  OAI22_X1 U13729 ( .A1(n12610), .A2(n15104), .B1(n11210), .B2(n15106), .ZN(
        n11211) );
  AOI21_X1 U13730 ( .B1(n11212), .B2(n15109), .A(n11211), .ZN(n11213) );
  OAI21_X1 U13731 ( .B1(n15112), .B2(n15129), .A(n11213), .ZN(n15130) );
  NAND2_X1 U13732 ( .A1(n15130), .A2(n15120), .ZN(n11218) );
  AND2_X1 U13733 ( .A1(n12035), .A2(n14476), .ZN(n15131) );
  INV_X1 U13734 ( .A(n15131), .ZN(n11215) );
  OAI22_X1 U13735 ( .A1(n11406), .A2(n11215), .B1(n11214), .B2(n15114), .ZN(
        n11216) );
  AOI21_X1 U13736 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n14462), .A(n11216), .ZN(
        n11217) );
  OAI211_X1 U13737 ( .C1(n15129), .C2(n15116), .A(n11218), .B(n11217), .ZN(
        P3_U3225) );
  NAND2_X1 U13738 ( .A1(n11220), .A2(n13461), .ZN(n11223) );
  AOI22_X1 U13739 ( .A1(n11221), .A2(n11514), .B1(n11515), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n11222) );
  OR2_X1 U13740 ( .A1(n14546), .A2(n11885), .ZN(n13604) );
  NAND2_X1 U13741 ( .A1(n14546), .A2(n11885), .ZN(n13610) );
  NAND2_X1 U13742 ( .A1(n11225), .A2(n13461), .ZN(n11227) );
  AOI22_X1 U13743 ( .A1(n11515), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11514), 
        .B2(n14638), .ZN(n11226) );
  AND2_X1 U13744 ( .A1(n11229), .A2(n11228), .ZN(n11230) );
  OR2_X1 U13745 ( .A1(n11230), .A2(n11237), .ZN(n11248) );
  INV_X1 U13746 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11415) );
  OR2_X1 U13747 ( .A1(n6428), .A2(n11415), .ZN(n11233) );
  INV_X1 U13748 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11231) );
  OR2_X1 U13749 ( .A1(n6467), .A2(n11231), .ZN(n11232) );
  AND2_X1 U13750 ( .A1(n11233), .A2(n11232), .ZN(n11235) );
  OR2_X1 U13751 ( .A1(n6426), .A2(n14635), .ZN(n11234) );
  OAI211_X1 U13752 ( .C1(n11248), .C2(n6465), .A(n11235), .B(n11234), .ZN(
        n14086) );
  INV_X1 U13753 ( .A(n14086), .ZN(n14537) );
  NAND2_X1 U13754 ( .A1(n13612), .A2(n14537), .ZN(n13623) );
  NAND2_X1 U13755 ( .A1(n13616), .A2(n13623), .ZN(n13487) );
  OAI211_X1 U13756 ( .C1(n6603), .C2(n11236), .A(n11433), .B(n14183), .ZN(
        n11241) );
  OR2_X1 U13757 ( .A1(n11237), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n11238) );
  NAND2_X1 U13758 ( .A1(n11437), .A2(n11238), .ZN(n14077) );
  AOI22_X1 U13759 ( .A1(n11600), .A2(P1_REG0_REG_16__SCAN_IN), .B1(n6688), 
        .B2(P1_REG2_REG_16__SCAN_IN), .ZN(n11240) );
  NAND2_X1 U13760 ( .A1(n13450), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n11239) );
  OAI211_X1 U13761 ( .C1(n14077), .C2(n6465), .A(n11240), .B(n11239), .ZN(
        n13737) );
  INV_X1 U13762 ( .A(n11885), .ZN(n13738) );
  AOI22_X1 U13763 ( .A1(n14083), .A2(n13737), .B1(n13738), .B2(n14085), .ZN(
        n13428) );
  NAND2_X1 U13764 ( .A1(n11241), .A2(n13428), .ZN(n11410) );
  INV_X1 U13765 ( .A(n11410), .ZN(n11253) );
  OR2_X1 U13766 ( .A1(n13607), .A2(n13739), .ZN(n11243) );
  NAND2_X1 U13767 ( .A1(n14546), .A2(n13738), .ZN(n11246) );
  OAI21_X1 U13768 ( .B1(n6596), .B2(n13487), .A(n11417), .ZN(n11412) );
  OR2_X1 U13769 ( .A1(n13435), .A2(n6607), .ZN(n11247) );
  AND3_X1 U13770 ( .A1(n14076), .A2(n11247), .A3(n14163), .ZN(n11411) );
  NAND2_X1 U13771 ( .A1(n11411), .A2(n14659), .ZN(n11250) );
  INV_X1 U13772 ( .A(n11248), .ZN(n13431) );
  AOI22_X1 U13773 ( .A1(n14673), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n13431), 
        .B2(n14662), .ZN(n11249) );
  OAI211_X1 U13774 ( .C1(n13435), .C2(n14666), .A(n11250), .B(n11249), .ZN(
        n11251) );
  AOI21_X1 U13775 ( .B1(n11412), .B2(n14655), .A(n11251), .ZN(n11252) );
  OAI21_X1 U13776 ( .B1(n14673), .B2(n11253), .A(n11252), .ZN(P1_U3278) );
  OAI21_X1 U13777 ( .B1(n11256), .B2(n11255), .A(n11254), .ZN(n11257) );
  NAND2_X1 U13778 ( .A1(n11257), .A2(n6997), .ZN(n11263) );
  INV_X1 U13779 ( .A(n11389), .ZN(n11261) );
  INV_X1 U13780 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n11258) );
  NOR2_X1 U13781 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n11258), .ZN(n14997) );
  AOI21_X1 U13782 ( .B1(n12142), .B2(n12107), .A(n14997), .ZN(n11259) );
  OAI21_X1 U13783 ( .B1(n12581), .B2(n12109), .A(n11259), .ZN(n11260) );
  AOI21_X1 U13784 ( .B1(n11261), .B2(n12117), .A(n11260), .ZN(n11262) );
  OAI211_X1 U13785 ( .C1(n14477), .C2(n12114), .A(n11263), .B(n11262), .ZN(
        P3_U3164) );
  INV_X1 U13786 ( .A(n11285), .ZN(n11270) );
  OR2_X1 U13787 ( .A1(n14520), .A2(n12857), .ZN(n11264) );
  NAND2_X1 U13788 ( .A1(n14520), .A2(n12857), .ZN(n11266) );
  NAND2_X1 U13789 ( .A1(n11267), .A2(n11266), .ZN(n11359) );
  XNOR2_X1 U13790 ( .A(n11359), .B(n11358), .ZN(n11269) );
  OAI22_X1 U13791 ( .A1(n12924), .A2(n12913), .B1(n11273), .B2(n12843), .ZN(
        n11283) );
  INV_X1 U13792 ( .A(n11283), .ZN(n11268) );
  OAI21_X1 U13793 ( .B1(n11269), .B2(n14834), .A(n11268), .ZN(n11376) );
  AOI21_X1 U13794 ( .B1(n11270), .B2(n14839), .A(n11376), .ZN(n11280) );
  OR2_X1 U13795 ( .A1(n14520), .A2(n11273), .ZN(n11274) );
  NAND2_X1 U13796 ( .A1(n11275), .A2(n11274), .ZN(n11354) );
  XNOR2_X1 U13797 ( .A(n11354), .B(n11358), .ZN(n11378) );
  NAND2_X1 U13798 ( .A1(n11375), .A2(n11276), .ZN(n11368) );
  OAI211_X1 U13799 ( .C1(n11375), .C2(n11276), .A(n14816), .B(n11368), .ZN(
        n11374) );
  AOI22_X1 U13800 ( .A1(n11287), .A2(n13141), .B1(n14844), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n11277) );
  OAI21_X1 U13801 ( .B1(n11374), .B2(n14820), .A(n11277), .ZN(n11278) );
  AOI21_X1 U13802 ( .B1(n11378), .B2(n14828), .A(n11278), .ZN(n11279) );
  OAI21_X1 U13803 ( .B1(n11280), .B2(n14844), .A(n11279), .ZN(P2_U3250) );
  AOI22_X1 U13804 ( .A1(n11281), .A2(n14494), .B1(n12822), .B2(n12856), .ZN(
        n11290) );
  INV_X1 U13805 ( .A(n11282), .ZN(n11289) );
  AOI22_X1 U13806 ( .A1(n14496), .A2(n11283), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11284) );
  OAI21_X1 U13807 ( .B1(n11285), .B2(n14502), .A(n11284), .ZN(n11286) );
  AOI21_X1 U13808 ( .B1(n11287), .B2(n14499), .A(n11286), .ZN(n11288) );
  OAI21_X1 U13809 ( .B1(n11290), .B2(n11289), .A(n11288), .ZN(P2_U3213) );
  INV_X1 U13810 ( .A(n11291), .ZN(n11293) );
  OAI222_X1 U13811 ( .A1(n11294), .A2(P3_U3151), .B1(n12747), .B2(n11293), 
        .C1(n11292), .C2(n12726), .ZN(P3_U3270) );
  NAND2_X1 U13812 ( .A1(n11566), .A2(n13289), .ZN(n11296) );
  OAI211_X1 U13813 ( .C1(n11297), .C2(n13303), .A(n11296), .B(n11295), .ZN(
        P2_U3304) );
  NAND2_X1 U13814 ( .A1(n11566), .A2(n14238), .ZN(n11298) );
  OAI211_X1 U13815 ( .C1(n11567), .C2(n14252), .A(n11298), .B(n13717), .ZN(
        P1_U3332) );
  NAND2_X1 U13816 ( .A1(n7450), .A2(n11299), .ZN(n11300) );
  XNOR2_X1 U13817 ( .A(n11301), .B(n11300), .ZN(n11306) );
  AND2_X1 U13818 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n15014) );
  NOR2_X1 U13819 ( .A1(n12597), .A2(n12109), .ZN(n11302) );
  AOI211_X1 U13820 ( .C1(n12107), .C2(n12141), .A(n15014), .B(n11302), .ZN(
        n11303) );
  OAI21_X1 U13821 ( .B1(n12598), .B2(n12130), .A(n11303), .ZN(n11304) );
  AOI21_X1 U13822 ( .B1(n14475), .B2(n12132), .A(n11304), .ZN(n11305) );
  OAI21_X1 U13823 ( .B1(n11306), .B2(n12134), .A(n11305), .ZN(P3_U3174) );
  NAND2_X1 U13824 ( .A1(n11308), .A2(n11307), .ZN(n12604) );
  NAND2_X1 U13825 ( .A1(n12604), .A2(n11309), .ZN(n11311) );
  NAND2_X1 U13826 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  XNOR2_X1 U13827 ( .A(n11312), .B(n11320), .ZN(n11315) );
  NAND2_X1 U13828 ( .A1(n12141), .A2(n12571), .ZN(n11313) );
  OAI21_X1 U13829 ( .B1(n11398), .B2(n15106), .A(n11313), .ZN(n11314) );
  AOI21_X1 U13830 ( .B1(n11315), .B2(n15109), .A(n11314), .ZN(n14485) );
  AND2_X1 U13831 ( .A1(n11316), .A2(n14476), .ZN(n14481) );
  INV_X1 U13832 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14973) );
  OAI22_X1 U13833 ( .A1(n15120), .A2(n14973), .B1(n11317), .B2(n15114), .ZN(
        n11318) );
  AOI21_X1 U13834 ( .B1(n11319), .B2(n14481), .A(n11318), .ZN(n11323) );
  XNOR2_X1 U13835 ( .A(n11321), .B(n11320), .ZN(n14483) );
  NAND2_X1 U13836 ( .A1(n14483), .A2(n12589), .ZN(n11322) );
  OAI211_X1 U13837 ( .C1(n14485), .C2(n14462), .A(n11323), .B(n11322), .ZN(
        P3_U3222) );
  NAND2_X1 U13838 ( .A1(n11324), .A2(n14546), .ZN(n11325) );
  NAND2_X1 U13839 ( .A1(n11325), .A2(n14163), .ZN(n11326) );
  NOR2_X1 U13840 ( .A1(n6607), .A2(n11326), .ZN(n14193) );
  NOR2_X1 U13841 ( .A1(n14044), .A2(n14549), .ZN(n11330) );
  XNOR2_X1 U13842 ( .A(n11327), .B(n11244), .ZN(n11328) );
  AOI222_X1 U13843 ( .A1(n14183), .A2(n11328), .B1(n14086), .B2(n14083), .C1(
        n13739), .C2(n14085), .ZN(n14198) );
  INV_X1 U13844 ( .A(n14198), .ZN(n11329) );
  AOI211_X1 U13845 ( .C1(n14193), .C2(n13920), .A(n11330), .B(n11329), .ZN(
        n11334) );
  AOI22_X1 U13846 ( .A1(n14546), .A2(n13994), .B1(n14673), .B2(
        P1_REG2_REG_14__SCAN_IN), .ZN(n11333) );
  NAND2_X1 U13847 ( .A1(n11331), .A2(n13617), .ZN(n14194) );
  NAND3_X1 U13848 ( .A1(n14195), .A2(n14194), .A3(n14655), .ZN(n11332) );
  OAI211_X1 U13849 ( .C1(n11334), .C2(n14650), .A(n11333), .B(n11332), .ZN(
        P1_U3279) );
  NOR2_X1 U13850 ( .A1(n11336), .A2(n11335), .ZN(n11338) );
  NOR2_X1 U13851 ( .A1(n11338), .A2(n11337), .ZN(n11340) );
  XNOR2_X1 U13852 ( .A(n12882), .B(P2_REG1_REG_16__SCAN_IN), .ZN(n11339) );
  NOR2_X1 U13853 ( .A1(n11340), .A2(n11339), .ZN(n12881) );
  AOI211_X1 U13854 ( .C1(n11340), .C2(n11339), .A(n14795), .B(n12881), .ZN(
        n11353) );
  NAND2_X1 U13855 ( .A1(n11342), .A2(n11341), .ZN(n11344) );
  NAND2_X1 U13856 ( .A1(n11344), .A2(n11343), .ZN(n11348) );
  NAND2_X1 U13857 ( .A1(n12882), .A2(n11367), .ZN(n11345) );
  OAI21_X1 U13858 ( .B1(n12882), .B2(n11367), .A(n11345), .ZN(n11347) );
  NAND2_X1 U13859 ( .A1(n12874), .A2(n11367), .ZN(n11346) );
  OAI211_X1 U13860 ( .C1(n12874), .C2(n11367), .A(n11348), .B(n11346), .ZN(
        n12873) );
  OAI211_X1 U13861 ( .C1(n11348), .C2(n11347), .A(n12873), .B(n14800), .ZN(
        n11351) );
  NAND2_X1 U13862 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3088), .ZN(n11464)
         );
  INV_X1 U13863 ( .A(n11464), .ZN(n11349) );
  AOI21_X1 U13864 ( .B1(n14799), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n11349), 
        .ZN(n11350) );
  OAI211_X1 U13865 ( .C1(n12878), .C2(n12874), .A(n11351), .B(n11350), .ZN(
        n11352) );
  OR2_X1 U13866 ( .A1(n11353), .A2(n11352), .ZN(P2_U3230) );
  NAND2_X1 U13867 ( .A1(n11375), .A2(n11364), .ZN(n11355) );
  INV_X1 U13868 ( .A(n11362), .ZN(n12922) );
  NAND2_X1 U13869 ( .A1(n11356), .A2(n12922), .ZN(n11357) );
  NAND2_X1 U13870 ( .A1(n12957), .A2(n11357), .ZN(n13262) );
  NAND2_X1 U13871 ( .A1(n11359), .A2(n11358), .ZN(n11361) );
  NAND2_X1 U13872 ( .A1(n11375), .A2(n12856), .ZN(n11360) );
  NAND2_X1 U13873 ( .A1(n11361), .A2(n11360), .ZN(n12923) );
  XNOR2_X1 U13874 ( .A(n12923), .B(n11362), .ZN(n11363) );
  NAND2_X1 U13875 ( .A1(n11363), .A2(n14814), .ZN(n11366) );
  INV_X1 U13876 ( .A(n12958), .ZN(n12959) );
  NOR2_X1 U13877 ( .A1(n11364), .A2(n12843), .ZN(n11365) );
  AOI21_X1 U13878 ( .B1(n12959), .B2(n12781), .A(n11365), .ZN(n11465) );
  NAND2_X1 U13879 ( .A1(n11366), .A2(n11465), .ZN(n13264) );
  NAND2_X1 U13880 ( .A1(n13264), .A2(n14515), .ZN(n11373) );
  OAI22_X1 U13881 ( .A1(n14515), .A2(n11367), .B1(n11463), .B2(n14819), .ZN(
        n11371) );
  AND2_X1 U13882 ( .A1(n13258), .A2(n11368), .ZN(n11369) );
  OR3_X1 U13883 ( .A1(n13168), .A2(n11369), .A3(n13169), .ZN(n13260) );
  NOR2_X1 U13884 ( .A1(n13260), .A2(n14820), .ZN(n11370) );
  AOI211_X1 U13885 ( .C1(n13141), .C2(n13258), .A(n11371), .B(n11370), .ZN(
        n11372) );
  OAI211_X1 U13886 ( .C1(n13178), .C2(n13262), .A(n11373), .B(n11372), .ZN(
        P2_U3249) );
  OAI21_X1 U13887 ( .B1(n11375), .B2(n14933), .A(n11374), .ZN(n11377) );
  AOI211_X1 U13888 ( .C1(n14913), .C2(n11378), .A(n11377), .B(n11376), .ZN(
        n11381) );
  NAND2_X1 U13889 ( .A1(n14950), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n11379) );
  OAI21_X1 U13890 ( .B1(n11381), .B2(n14950), .A(n11379), .ZN(P2_U3475) );
  NAND2_X1 U13891 ( .A1(n14968), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n11380) );
  OAI21_X1 U13892 ( .B1(n11381), .B2(n14968), .A(n11380), .ZN(P2_U3514) );
  INV_X1 U13893 ( .A(n11382), .ZN(n11384) );
  OAI211_X1 U13894 ( .C1(n11384), .C2(n7189), .A(n15109), .B(n11383), .ZN(
        n11386) );
  AOI22_X1 U13895 ( .A1(n12569), .A2(n12142), .B1(n12140), .B2(n12571), .ZN(
        n11385) );
  NAND2_X1 U13896 ( .A1(n11386), .A2(n11385), .ZN(n14478) );
  INV_X1 U13897 ( .A(n14478), .ZN(n11394) );
  OAI21_X1 U13898 ( .B1(n11388), .B2(n11827), .A(n11387), .ZN(n14480) );
  NOR2_X1 U13899 ( .A1(n12587), .A2(n14477), .ZN(n11392) );
  INV_X1 U13900 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n11390) );
  OAI22_X1 U13901 ( .A1(n15120), .A2(n11390), .B1(n11389), .B2(n15114), .ZN(
        n11391) );
  AOI211_X1 U13902 ( .C1(n14480), .C2(n12589), .A(n11392), .B(n11391), .ZN(
        n11393) );
  OAI21_X1 U13903 ( .B1(n11394), .B2(n14462), .A(n11393), .ZN(P3_U3221) );
  NAND2_X1 U13904 ( .A1(n11395), .A2(n11820), .ZN(n11396) );
  NAND2_X1 U13905 ( .A1(n11396), .A2(n11722), .ZN(n11397) );
  XNOR2_X1 U13906 ( .A(n11397), .B(n12603), .ZN(n15133) );
  XOR2_X1 U13907 ( .A(n12603), .B(n12604), .Z(n11401) );
  OAI22_X1 U13908 ( .A1(n11399), .A2(n15106), .B1(n11398), .B2(n15104), .ZN(
        n11400) );
  AOI21_X1 U13909 ( .B1(n11401), .B2(n15109), .A(n11400), .ZN(n11402) );
  OAI21_X1 U13910 ( .B1(n15112), .B2(n15133), .A(n11402), .ZN(n15134) );
  NAND2_X1 U13911 ( .A1(n15134), .A2(n15120), .ZN(n11409) );
  NOR2_X1 U13912 ( .A1(n11403), .A2(n15138), .ZN(n15135) );
  INV_X1 U13913 ( .A(n15135), .ZN(n11405) );
  OAI22_X1 U13914 ( .A1(n11406), .A2(n11405), .B1(n11404), .B2(n15114), .ZN(
        n11407) );
  AOI21_X1 U13915 ( .B1(n14462), .B2(P3_REG2_REG_9__SCAN_IN), .A(n11407), .ZN(
        n11408) );
  OAI211_X1 U13916 ( .C1(n15133), .C2(n15116), .A(n11409), .B(n11408), .ZN(
        P3_U3224) );
  AOI211_X1 U13917 ( .C1(n11412), .C2(n14725), .A(n11411), .B(n11410), .ZN(
        n11414) );
  MUX2_X1 U13918 ( .A(n14635), .B(n11414), .S(n14734), .Z(n11413) );
  OAI21_X1 U13919 ( .B1(n13435), .B2(n14172), .A(n11413), .ZN(P1_U3543) );
  MUX2_X1 U13920 ( .A(n11415), .B(n11414), .S(n14729), .Z(n11416) );
  OAI21_X1 U13921 ( .B1(n13435), .B2(n14227), .A(n11416), .ZN(P1_U3504) );
  NAND2_X1 U13922 ( .A1(n11418), .A2(n13461), .ZN(n11420) );
  AOI22_X1 U13923 ( .A1(n11515), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11514), 
        .B2(n13818), .ZN(n11419) );
  XNOR2_X1 U13924 ( .A(n14188), .B(n13737), .ZN(n14081) );
  INV_X1 U13925 ( .A(n14081), .ZN(n11421) );
  NAND2_X1 U13926 ( .A1(n14073), .A2(n11421), .ZN(n11423) );
  OR2_X1 U13927 ( .A1(n14188), .A2(n13737), .ZN(n11422) );
  NAND2_X1 U13928 ( .A1(n11424), .A2(n13461), .ZN(n11426) );
  AOI22_X1 U13929 ( .A1(n11515), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11514), 
        .B2(n13833), .ZN(n11425) );
  XNOR2_X1 U13930 ( .A(n11437), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n13374) );
  NAND2_X1 U13931 ( .A1(n13374), .A2(n11545), .ZN(n11432) );
  INV_X1 U13932 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n13810) );
  NAND2_X1 U13933 ( .A1(n11600), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11429) );
  INV_X1 U13934 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11427) );
  OR2_X1 U13935 ( .A1(n6426), .A2(n11427), .ZN(n11428) );
  OAI211_X1 U13936 ( .C1(n6467), .C2(n13810), .A(n11429), .B(n11428), .ZN(
        n11430) );
  INV_X1 U13937 ( .A(n11430), .ZN(n11431) );
  NAND2_X1 U13938 ( .A1(n13638), .A2(n14084), .ZN(n11506) );
  NAND2_X1 U13939 ( .A1(n11503), .A2(n11506), .ZN(n13489) );
  XNOR2_X1 U13940 ( .A(n11505), .B(n13489), .ZN(n14186) );
  INV_X1 U13941 ( .A(n13737), .ZN(n11434) );
  NAND2_X1 U13942 ( .A1(n14188), .A2(n11434), .ZN(n11435) );
  NAND2_X1 U13943 ( .A1(n14080), .A2(n11435), .ZN(n11592) );
  XNOR2_X1 U13944 ( .A(n11592), .B(n13489), .ZN(n14184) );
  NAND2_X1 U13945 ( .A1(n14181), .A2(n14074), .ZN(n14065) );
  OAI211_X1 U13946 ( .C1(n14181), .C2(n14074), .A(n14163), .B(n14065), .ZN(
        n14180) );
  NOR2_X1 U13947 ( .A1(n14047), .A2(n13810), .ZN(n11443) );
  INV_X1 U13948 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n13835) );
  INV_X1 U13949 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n13370) );
  OAI21_X1 U13950 ( .B1(n11437), .B2(n13370), .A(n12188), .ZN(n11438) );
  NAND2_X1 U13951 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n11436) );
  AND2_X1 U13952 ( .A1(n11438), .A2(n11518), .ZN(n14066) );
  NAND2_X1 U13953 ( .A1(n14066), .A2(n11545), .ZN(n11440) );
  AOI22_X1 U13954 ( .A1(n11600), .A2(P1_REG0_REG_18__SCAN_IN), .B1(n6688), 
        .B2(P1_REG2_REG_18__SCAN_IN), .ZN(n11439) );
  OAI211_X1 U13955 ( .C1(n6426), .C2(n13835), .A(n11440), .B(n11439), .ZN(
        n13736) );
  AOI22_X1 U13956 ( .A1(n13736), .A2(n14083), .B1(n14085), .B2(n13737), .ZN(
        n14179) );
  INV_X1 U13957 ( .A(n13374), .ZN(n11441) );
  OAI22_X1 U13958 ( .A1(n14179), .A2(n14650), .B1(n11441), .B2(n14044), .ZN(
        n11442) );
  AOI211_X1 U13959 ( .C1(n13638), .C2(n13994), .A(n11443), .B(n11442), .ZN(
        n11444) );
  OAI21_X1 U13960 ( .B1(n14180), .B2(n13975), .A(n11444), .ZN(n11445) );
  AOI21_X1 U13961 ( .B1(n14184), .B2(n13896), .A(n11445), .ZN(n11446) );
  OAI21_X1 U13962 ( .B1(n14186), .B2(n14091), .A(n11446), .ZN(P1_U3276) );
  INV_X1 U13963 ( .A(n11499), .ZN(n11450) );
  OAI222_X1 U13964 ( .A1(n13303), .A2(n7046), .B1(n13301), .B2(n11450), .C1(
        P2_U3088), .C2(n11447), .ZN(P2_U3303) );
  INV_X1 U13965 ( .A(n11448), .ZN(n11449) );
  OAI222_X1 U13966 ( .A1(n14252), .A2(n11500), .B1(n10724), .B2(n11450), .C1(
        n11449), .C2(P1_U3086), .ZN(P1_U3331) );
  INV_X1 U13967 ( .A(n12961), .ZN(n12928) );
  AOI22_X1 U13968 ( .A1(n12928), .A2(n12781), .B1(n12947), .B2(n12956), .ZN(
        n13166) );
  NAND2_X1 U13969 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n14808)
         );
  NAND2_X1 U13970 ( .A1(n12842), .A2(n13172), .ZN(n11451) );
  OAI211_X1 U13971 ( .C1(n13166), .C2(n12783), .A(n14808), .B(n11451), .ZN(
        n11452) );
  AOI21_X1 U13972 ( .B1(n13255), .B2(n14499), .A(n11452), .ZN(n11457) );
  OAI22_X1 U13973 ( .A1(n11454), .A2(n12816), .B1(n12924), .B2(n12837), .ZN(
        n11455) );
  NAND3_X1 U13974 ( .A1(n11459), .A2(n7152), .A3(n11455), .ZN(n11456) );
  OAI211_X1 U13975 ( .C1(n11458), .C2(n12816), .A(n11457), .B(n11456), .ZN(
        P2_U3200) );
  INV_X1 U13976 ( .A(n11459), .ZN(n11460) );
  AOI21_X1 U13977 ( .B1(n11462), .B2(n11461), .A(n11460), .ZN(n11469) );
  NOR2_X1 U13978 ( .A1(n14502), .A2(n11463), .ZN(n11467) );
  OAI21_X1 U13979 ( .B1(n12783), .B2(n11465), .A(n11464), .ZN(n11466) );
  AOI211_X1 U13980 ( .C1(n13258), .C2(n14499), .A(n11467), .B(n11466), .ZN(
        n11468) );
  OAI21_X1 U13981 ( .B1(n11469), .B2(n12816), .A(n11468), .ZN(P2_U3198) );
  INV_X1 U13982 ( .A(n13445), .ZN(n11646) );
  OAI222_X1 U13983 ( .A1(n13301), .A2(n11646), .B1(P2_U3088), .B2(n11470), 
        .C1(n11648), .C2(n13303), .ZN(P2_U3297) );
  NOR2_X1 U13984 ( .A1(n12913), .A2(n11471), .ZN(n14835) );
  AOI22_X1 U13985 ( .A1(n14496), .A2(n14835), .B1(n14494), .B2(n11472), .ZN(
        n11474) );
  AOI22_X1 U13986 ( .A1(n14499), .A2(n14855), .B1(P2_REG3_REG_0__SCAN_IN), 
        .B2(n11626), .ZN(n11473) );
  OAI211_X1 U13987 ( .C1(n9136), .C2(n12837), .A(n11474), .B(n11473), .ZN(
        P2_U3204) );
  NAND2_X1 U13988 ( .A1(n13296), .A2(n13461), .ZN(n11476) );
  OR2_X1 U13989 ( .A1(n13464), .A2(n14245), .ZN(n11475) );
  NAND2_X1 U13990 ( .A1(n11600), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n11482) );
  INV_X1 U13991 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13922) );
  OR2_X1 U13992 ( .A1(n6467), .A2(n13922), .ZN(n11481) );
  NAND2_X1 U13993 ( .A1(n11494), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U13994 ( .A1(n11485), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11484) );
  NAND2_X1 U13995 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n11477), .ZN(n11582) );
  OAI21_X1 U13996 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n11477), .A(n11582), 
        .ZN(n13921) );
  OR2_X1 U13997 ( .A1(n6465), .A2(n13921), .ZN(n11480) );
  INV_X1 U13998 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n11478) );
  OR2_X1 U13999 ( .A1(n6426), .A2(n11478), .ZN(n11479) );
  NAND4_X1 U14000 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n13934) );
  NAND2_X1 U14001 ( .A1(n11600), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n11490) );
  INV_X1 U14002 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n11483) );
  OR2_X1 U14003 ( .A1(n6467), .A2(n11483), .ZN(n11489) );
  OAI21_X1 U14004 ( .B1(P1_REG3_REG_25__SCAN_IN), .B2(n11485), .A(n11484), 
        .ZN(n13941) );
  OR2_X1 U14005 ( .A1(n6465), .A2(n13941), .ZN(n11488) );
  INV_X1 U14006 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11486) );
  OR2_X1 U14007 ( .A1(n6426), .A2(n11486), .ZN(n11487) );
  NAND4_X1 U14008 ( .A1(n11490), .A2(n11489), .A3(n11488), .A4(n11487), .ZN(
        n13731) );
  INV_X1 U14009 ( .A(n13731), .ZN(n13953) );
  NAND2_X1 U14010 ( .A1(n13299), .A2(n13461), .ZN(n11492) );
  OR2_X1 U14011 ( .A1(n13464), .A2(n14251), .ZN(n11491) );
  NAND2_X1 U14012 ( .A1(n11600), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n11498) );
  INV_X1 U14013 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13963) );
  OR2_X1 U14014 ( .A1(n6467), .A2(n13963), .ZN(n11497) );
  OAI21_X1 U14015 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11494), .A(n11493), 
        .ZN(n13962) );
  OR2_X1 U14016 ( .A1(n6465), .A2(n13962), .ZN(n11496) );
  INV_X1 U14017 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n14138) );
  OR2_X1 U14018 ( .A1(n6426), .A2(n14138), .ZN(n11495) );
  NAND4_X1 U14019 ( .A1(n11498), .A2(n11497), .A3(n11496), .A4(n11495), .ZN(
        n13983) );
  NAND2_X1 U14020 ( .A1(n11499), .A2(n13461), .ZN(n11502) );
  OR2_X1 U14021 ( .A1(n13464), .A2(n11500), .ZN(n11501) );
  INV_X1 U14022 ( .A(n11503), .ZN(n11504) );
  NAND2_X1 U14023 ( .A1(n11507), .A2(n13461), .ZN(n11509) );
  AOI22_X1 U14024 ( .A1(n11515), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11514), 
        .B2(n13847), .ZN(n11508) );
  AND2_X1 U14025 ( .A1(n14175), .A2(n13736), .ZN(n11511) );
  OR2_X1 U14026 ( .A1(n14175), .A2(n13736), .ZN(n11510) );
  NAND2_X1 U14027 ( .A1(n11512), .A2(n13461), .ZN(n11517) );
  AOI22_X1 U14028 ( .A1(n11515), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11514), 
        .B2(n11513), .ZN(n11516) );
  AND2_X1 U14029 ( .A1(n11518), .A2(n13325), .ZN(n11519) );
  OR2_X1 U14030 ( .A1(n11519), .A2(n11530), .ZN(n14045) );
  INV_X1 U14031 ( .A(n14045), .ZN(n11523) );
  INV_X1 U14032 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n14046) );
  NAND2_X1 U14033 ( .A1(n11600), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11521) );
  NAND2_X1 U14034 ( .A1(n13450), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n11520) );
  OAI211_X1 U14035 ( .C1(n6467), .C2(n14046), .A(n11521), .B(n11520), .ZN(
        n11522) );
  AOI21_X1 U14036 ( .B1(n11523), .B2(n11545), .A(n11522), .ZN(n14061) );
  OR2_X1 U14037 ( .A1(n14043), .A2(n14061), .ZN(n13655) );
  AND2_X1 U14038 ( .A1(n14043), .A2(n14061), .ZN(n13642) );
  NAND2_X1 U14039 ( .A1(n13655), .A2(n13659), .ZN(n14040) );
  INV_X1 U14040 ( .A(n14061), .ZN(n13735) );
  OR2_X1 U14041 ( .A1(n14043), .A2(n13735), .ZN(n11524) );
  NAND2_X1 U14042 ( .A1(n11526), .A2(n13461), .ZN(n11529) );
  OR2_X1 U14043 ( .A1(n13464), .A2(n11527), .ZN(n11528) );
  NOR2_X1 U14044 ( .A1(n11530), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n11531) );
  NOR2_X1 U14045 ( .A1(n11542), .A2(n11531), .ZN(n14026) );
  NAND2_X1 U14046 ( .A1(n14026), .A2(n11545), .ZN(n11536) );
  INV_X1 U14047 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n12203) );
  NAND2_X1 U14048 ( .A1(n13450), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U14049 ( .A1(n6688), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11532) );
  OAI211_X1 U14050 ( .C1(n6428), .C2(n12203), .A(n11533), .B(n11532), .ZN(
        n11534) );
  INV_X1 U14051 ( .A(n11534), .ZN(n11535) );
  XNOR2_X1 U14052 ( .A(n14157), .B(n13734), .ZN(n14033) );
  OR2_X1 U14053 ( .A1(n14028), .A2(n13522), .ZN(n11538) );
  NAND2_X1 U14054 ( .A1(n11539), .A2(n13461), .ZN(n11541) );
  OR2_X1 U14055 ( .A1(n13464), .A2(n6752), .ZN(n11540) );
  OR2_X1 U14056 ( .A1(n11542), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n11544) );
  AND2_X1 U14057 ( .A1(n11544), .A2(n11543), .ZN(n14013) );
  NAND2_X1 U14058 ( .A1(n14013), .A2(n11545), .ZN(n11550) );
  INV_X1 U14059 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U14060 ( .A1(n13450), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n11547) );
  NAND2_X1 U14061 ( .A1(n6688), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11546) );
  OAI211_X1 U14062 ( .C1(n6428), .C2(n14220), .A(n11547), .B(n11546), .ZN(
        n11548) );
  INV_X1 U14063 ( .A(n11548), .ZN(n11549) );
  NAND2_X1 U14064 ( .A1(n11550), .A2(n11549), .ZN(n13733) );
  OR2_X1 U14065 ( .A1(n14010), .A2(n13733), .ZN(n11552) );
  NAND2_X1 U14066 ( .A1(n14010), .A2(n13733), .ZN(n11551) );
  NAND2_X1 U14067 ( .A1(n11552), .A2(n11551), .ZN(n14008) );
  OR2_X1 U14068 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  XNOR2_X1 U14069 ( .A(n11555), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14253) );
  NAND2_X1 U14070 ( .A1(n11600), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11563) );
  INV_X1 U14071 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n11556) );
  OR2_X1 U14072 ( .A1(n6467), .A2(n11556), .ZN(n11562) );
  OAI21_X1 U14073 ( .B1(P1_REG3_REG_22__SCAN_IN), .B2(n11559), .A(n11558), 
        .ZN(n13992) );
  OR2_X1 U14074 ( .A1(n6465), .A2(n13992), .ZN(n11561) );
  INV_X1 U14075 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14149) );
  OR2_X1 U14076 ( .A1(n6426), .A2(n14149), .ZN(n11560) );
  NAND4_X1 U14077 ( .A1(n11563), .A2(n11562), .A3(n11561), .A4(n11560), .ZN(
        n13982) );
  XNOR2_X1 U14078 ( .A(n7363), .B(n13982), .ZN(n13996) );
  OR2_X1 U14079 ( .A1(n13997), .A2(n13982), .ZN(n11564) );
  NAND2_X1 U14080 ( .A1(n11566), .A2(n13461), .ZN(n11569) );
  OR2_X1 U14081 ( .A1(n13464), .A2(n11567), .ZN(n11568) );
  NAND2_X1 U14082 ( .A1(n6688), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11576) );
  INV_X1 U14083 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n12215) );
  OR2_X1 U14084 ( .A1(n6428), .A2(n12215), .ZN(n11575) );
  OAI21_X1 U14085 ( .B1(P1_REG3_REG_23__SCAN_IN), .B2(n11571), .A(n11570), 
        .ZN(n13971) );
  OR2_X1 U14086 ( .A1(n6465), .A2(n13971), .ZN(n11574) );
  INV_X1 U14087 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11572) );
  OR2_X1 U14088 ( .A1(n6426), .A2(n11572), .ZN(n11573) );
  NAND4_X1 U14089 ( .A1(n11576), .A2(n11575), .A3(n11574), .A4(n11573), .ZN(
        n13732) );
  XNOR2_X1 U14090 ( .A(n13978), .B(n13990), .ZN(n13493) );
  XNOR2_X1 U14091 ( .A(n13961), .B(n13352), .ZN(n13952) );
  INV_X1 U14092 ( .A(n13952), .ZN(n13949) );
  XNOR2_X1 U14093 ( .A(n13943), .B(n13731), .ZN(n13932) );
  INV_X1 U14094 ( .A(n13932), .ZN(n13938) );
  NAND2_X1 U14095 ( .A1(n13928), .A2(n13310), .ZN(n11598) );
  OR2_X1 U14096 ( .A1(n13928), .A2(n13310), .ZN(n11577) );
  NAND2_X1 U14097 ( .A1(n11598), .A2(n11577), .ZN(n13924) );
  NAND2_X1 U14098 ( .A1(n13293), .A2(n13461), .ZN(n11579) );
  OR2_X1 U14099 ( .A1(n13464), .A2(n7070), .ZN(n11578) );
  NAND2_X1 U14100 ( .A1(n11600), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n11588) );
  INV_X1 U14101 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n11618) );
  OR2_X1 U14102 ( .A1(n6467), .A2(n11618), .ZN(n11587) );
  INV_X1 U14103 ( .A(n11582), .ZN(n11580) );
  NAND2_X1 U14104 ( .A1(n11580), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11604) );
  INV_X1 U14105 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14106 ( .A1(n11582), .A2(n11581), .ZN(n11583) );
  NAND2_X1 U14107 ( .A1(n11604), .A2(n11583), .ZN(n13308) );
  OR2_X1 U14108 ( .A1(n6465), .A2(n13308), .ZN(n11586) );
  INV_X1 U14109 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n11584) );
  OR2_X1 U14110 ( .A1(n6426), .A2(n11584), .ZN(n11585) );
  NAND4_X1 U14111 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n13903) );
  NOR2_X1 U14112 ( .A1(n14181), .A2(n14084), .ZN(n11591) );
  NAND2_X1 U14113 ( .A1(n14181), .A2(n14084), .ZN(n11590) );
  XNOR2_X1 U14114 ( .A(n14175), .B(n13736), .ZN(n14056) );
  INV_X1 U14115 ( .A(n13736), .ZN(n13372) );
  NOR2_X1 U14116 ( .A1(n14175), .A2(n13372), .ZN(n11593) );
  INV_X1 U14117 ( .A(n14040), .ZN(n14037) );
  NAND2_X1 U14118 ( .A1(n14028), .A2(n13734), .ZN(n11594) );
  NAND2_X1 U14119 ( .A1(n14004), .A2(n14008), .ZN(n11596) );
  INV_X1 U14120 ( .A(n13733), .ZN(n14021) );
  OR2_X1 U14121 ( .A1(n14010), .A2(n14021), .ZN(n11595) );
  INV_X1 U14122 ( .A(n13982), .ZN(n13331) );
  NAND2_X1 U14123 ( .A1(n13997), .A2(n13331), .ZN(n11597) );
  INV_X1 U14124 ( .A(n13924), .ZN(n13917) );
  OAI21_X1 U14125 ( .B1(n11599), .B2(n13495), .A(n13876), .ZN(n11614) );
  NAND2_X1 U14126 ( .A1(n11600), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n11612) );
  INV_X1 U14127 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11601) );
  OR2_X1 U14128 ( .A1(n6467), .A2(n11601), .ZN(n11611) );
  INV_X1 U14129 ( .A(n11604), .ZN(n11602) );
  NAND2_X1 U14130 ( .A1(n11602), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n13886) );
  INV_X1 U14131 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14132 ( .A1(n11604), .A2(n11603), .ZN(n11605) );
  NAND2_X1 U14133 ( .A1(n13886), .A2(n11605), .ZN(n13906) );
  OR2_X1 U14134 ( .A1(n6465), .A2(n13906), .ZN(n11610) );
  INV_X1 U14135 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n11607) );
  OR2_X1 U14136 ( .A1(n6426), .A2(n11607), .ZN(n11609) );
  NAND4_X1 U14137 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n13888) );
  INV_X1 U14138 ( .A(n13888), .ZN(n13878) );
  OAI22_X1 U14139 ( .A1(n13878), .A2(n14060), .B1(n13310), .B2(n14020), .ZN(
        n11613) );
  AOI21_X1 U14140 ( .B1(n14115), .B2(n11617), .A(n13861), .ZN(n14116) );
  NOR2_X1 U14141 ( .A1(n13877), .A2(n14666), .ZN(n11620) );
  OAI22_X1 U14142 ( .A1(n14047), .A2(n11618), .B1(n13308), .B2(n14044), .ZN(
        n11619) );
  AOI211_X1 U14143 ( .C1(n14116), .C2(n14051), .A(n11620), .B(n11619), .ZN(
        n11623) );
  INV_X1 U14144 ( .A(n14118), .ZN(n11621) );
  NAND2_X1 U14145 ( .A1(n11621), .A2(n14669), .ZN(n11622) );
  OAI211_X1 U14146 ( .C1(n14121), .C2(n14650), .A(n11623), .B(n11622), .ZN(
        P1_U3266) );
  OAI22_X1 U14147 ( .A1(n11625), .A2(n12913), .B1(n12843), .B2(n11624), .ZN(
        n11639) );
  AOI22_X1 U14148 ( .A1(n14496), .A2(n11639), .B1(P2_REG3_REG_1__SCAN_IN), 
        .B2(n11626), .ZN(n11632) );
  OAI21_X1 U14149 ( .B1(n11629), .B2(n11628), .A(n11627), .ZN(n11630) );
  NAND2_X1 U14150 ( .A1(n14494), .A2(n11630), .ZN(n11631) );
  OAI211_X1 U14151 ( .C1(n14865), .C2(n12846), .A(n11632), .B(n11631), .ZN(
        P2_U3194) );
  XNOR2_X1 U14152 ( .A(n11637), .B(n11633), .ZN(n14862) );
  OAI211_X1 U14153 ( .C1(n14865), .C2(n14831), .A(n14816), .B(n11634), .ZN(
        n14863) );
  INV_X1 U14154 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11635) );
  OAI22_X1 U14155 ( .A1(n14820), .A2(n14863), .B1(n11635), .B2(n14819), .ZN(
        n11643) );
  OAI21_X1 U14156 ( .B1(n11638), .B2(n11637), .A(n11636), .ZN(n11640) );
  AOI21_X1 U14157 ( .B1(n11640), .B2(n14814), .A(n11639), .ZN(n14864) );
  NAND2_X1 U14158 ( .A1(n14844), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n11641) );
  OAI21_X1 U14159 ( .B1(n14864), .B2(n14844), .A(n11641), .ZN(n11642) );
  AOI211_X1 U14160 ( .C1(n13141), .C2(n6424), .A(n11643), .B(n11642), .ZN(
        n11645) );
  OAI21_X1 U14161 ( .B1(n13178), .B2(n14862), .A(n11645), .ZN(P2_U3264) );
  INV_X1 U14162 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U14163 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n11648), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n13446), .ZN(n11661) );
  OAI22_X1 U14164 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n13285), .B1(n11650), 
        .B2(n11649), .ZN(n11660) );
  AOI22_X1 U14165 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n9065), .B2(n14234), .ZN(n11651) );
  NAND2_X1 U14166 ( .A1(n11653), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n11658) );
  INV_X1 U14167 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14468) );
  OR2_X1 U14168 ( .A1(n8357), .A2(n14468), .ZN(n11657) );
  INV_X1 U14169 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n11654) );
  OR2_X1 U14170 ( .A1(n11655), .A2(n11654), .ZN(n11656) );
  NAND4_X1 U14171 ( .A1(n11659), .A2(n11658), .A3(n11657), .A4(n11656), .ZN(
        n14458) );
  NAND2_X1 U14172 ( .A1(n14465), .A2(n14458), .ZN(n11667) );
  XNOR2_X1 U14173 ( .A(n11661), .B(n11660), .ZN(n11997) );
  INV_X1 U14174 ( .A(n11997), .ZN(n11664) );
  INV_X1 U14175 ( .A(SI_30_), .ZN(n11996) );
  NOR2_X1 U14176 ( .A1(n8310), .A2(n11996), .ZN(n11662) );
  AOI21_X1 U14177 ( .B1(n11664), .B2(n11663), .A(n11662), .ZN(n11669) );
  INV_X1 U14178 ( .A(n11669), .ZN(n14470) );
  NAND2_X1 U14179 ( .A1(n14470), .A2(n11665), .ZN(n11666) );
  OAI21_X1 U14180 ( .B1(n11669), .B2(n14458), .A(n11807), .ZN(n11668) );
  OR2_X1 U14181 ( .A1(n14465), .A2(n14458), .ZN(n11839) );
  NAND2_X1 U14182 ( .A1(n11669), .A2(n12136), .ZN(n11809) );
  INV_X1 U14183 ( .A(n11809), .ZN(n11837) );
  INV_X1 U14184 ( .A(n14465), .ZN(n14460) );
  INV_X1 U14185 ( .A(n11675), .ZN(n11845) );
  MUX2_X1 U14186 ( .A(n11676), .B(n12144), .S(n11808), .Z(n11727) );
  OR2_X1 U14187 ( .A1(n11732), .A2(n12607), .ZN(n11813) );
  AOI211_X1 U14188 ( .C1(n11682), .C2(n11678), .A(n11804), .B(n11677), .ZN(
        n11684) );
  INV_X1 U14189 ( .A(n11678), .ZN(n11680) );
  NOR3_X1 U14190 ( .A1(n15102), .A2(n11680), .A3(n11679), .ZN(n11683) );
  OAI22_X1 U14191 ( .A1(n11684), .A2(n11683), .B1(n11682), .B2(n11681), .ZN(
        n11688) );
  MUX2_X1 U14192 ( .A(n11686), .B(n11685), .S(n11808), .Z(n11687) );
  NAND3_X1 U14193 ( .A1(n11688), .A2(n15085), .A3(n11687), .ZN(n11692) );
  INV_X1 U14194 ( .A(n11689), .ZN(n11690) );
  OAI21_X1 U14195 ( .B1(n11697), .B2(n11690), .A(n11808), .ZN(n11691) );
  AOI21_X1 U14196 ( .B1(n11695), .B2(n11693), .A(n11808), .ZN(n11694) );
  AOI21_X1 U14197 ( .B1(n11702), .B2(n11699), .A(n11804), .ZN(n11710) );
  AOI21_X1 U14198 ( .B1(n11706), .B2(n11700), .A(n11710), .ZN(n11701) );
  NAND3_X1 U14199 ( .A1(n11704), .A2(n11804), .A3(n11703), .ZN(n11705) );
  NAND2_X1 U14200 ( .A1(n11706), .A2(n11705), .ZN(n11713) );
  INV_X1 U14201 ( .A(n11707), .ZN(n11708) );
  NOR3_X1 U14202 ( .A1(n11710), .A2(n11709), .A3(n11708), .ZN(n11712) );
  AOI21_X1 U14203 ( .B1(n11713), .B2(n11712), .A(n11711), .ZN(n11720) );
  INV_X1 U14204 ( .A(n11714), .ZN(n11717) );
  INV_X1 U14205 ( .A(n11715), .ZN(n11716) );
  MUX2_X1 U14206 ( .A(n11717), .B(n11716), .S(n11808), .Z(n11719) );
  INV_X1 U14207 ( .A(n11721), .ZN(n11724) );
  INV_X1 U14208 ( .A(n11722), .ZN(n11723) );
  MUX2_X1 U14209 ( .A(n11724), .B(n11723), .S(n11808), .Z(n11725) );
  AOI211_X1 U14210 ( .C1(n12605), .C2(n11727), .A(n11813), .B(n11726), .ZN(
        n11739) );
  OAI211_X1 U14211 ( .C1(n11732), .C2(n11729), .A(n11728), .B(n11735), .ZN(
        n11734) );
  OAI211_X1 U14212 ( .C1(n11732), .C2(n11731), .A(n11736), .B(n11730), .ZN(
        n11733) );
  MUX2_X1 U14213 ( .A(n11734), .B(n11733), .S(n11808), .Z(n11738) );
  AND2_X1 U14214 ( .A1(n11741), .A2(n11740), .ZN(n12594) );
  MUX2_X1 U14215 ( .A(n11736), .B(n11735), .S(n11808), .Z(n11737) );
  OAI211_X1 U14216 ( .C1(n11739), .C2(n11738), .A(n12594), .B(n11737), .ZN(
        n11744) );
  MUX2_X1 U14217 ( .A(n11741), .B(n11740), .S(n11808), .Z(n11742) );
  AND3_X1 U14218 ( .A1(n11744), .A2(n11743), .A3(n11742), .ZN(n11749) );
  INV_X1 U14219 ( .A(n11746), .ZN(n11747) );
  MUX2_X1 U14220 ( .A(n7180), .B(n11747), .S(n11808), .Z(n11748) );
  OAI21_X1 U14221 ( .B1(n11749), .B2(n11748), .A(n12576), .ZN(n11759) );
  NOR2_X1 U14222 ( .A1(n11755), .A2(n7179), .ZN(n11754) );
  INV_X1 U14223 ( .A(n11751), .ZN(n11752) );
  NOR2_X1 U14224 ( .A1(n11756), .A2(n11752), .ZN(n11753) );
  MUX2_X1 U14225 ( .A(n11754), .B(n11753), .S(n11808), .Z(n11758) );
  MUX2_X1 U14226 ( .A(n11756), .B(n11755), .S(n11808), .Z(n11757) );
  AOI21_X1 U14227 ( .B1(n11759), .B2(n11758), .A(n11757), .ZN(n11763) );
  NAND2_X1 U14228 ( .A1(n11760), .A2(n11804), .ZN(n11761) );
  AOI211_X1 U14229 ( .C1(n11762), .C2(n11765), .A(n11761), .B(n11770), .ZN(
        n11764) );
  OAI22_X1 U14230 ( .A1(n11763), .A2(n11830), .B1(n11764), .B2(n12532), .ZN(
        n11768) );
  INV_X1 U14231 ( .A(n11764), .ZN(n11767) );
  NAND3_X1 U14232 ( .A1(n11769), .A2(n11765), .A3(n11808), .ZN(n11766) );
  INV_X1 U14233 ( .A(n11769), .ZN(n11771) );
  MUX2_X1 U14234 ( .A(n11771), .B(n11770), .S(n11808), .Z(n11772) );
  XNOR2_X1 U14235 ( .A(n11776), .B(n12470), .ZN(n12479) );
  NOR2_X1 U14236 ( .A1(n12505), .A2(n11808), .ZN(n11774) );
  NOR2_X1 U14237 ( .A1(n12651), .A2(n11804), .ZN(n11773) );
  MUX2_X1 U14238 ( .A(n11774), .B(n11773), .S(n12510), .Z(n11775) );
  NOR3_X1 U14239 ( .A1(n12708), .A2(n12499), .A3(n11808), .ZN(n11778) );
  NOR3_X1 U14240 ( .A1(n11776), .A2(n12470), .A3(n11804), .ZN(n11777) );
  NAND2_X1 U14241 ( .A1(n11779), .A2(n11780), .ZN(n12467) );
  INV_X1 U14242 ( .A(n11779), .ZN(n11782) );
  INV_X1 U14243 ( .A(n11780), .ZN(n11781) );
  MUX2_X1 U14244 ( .A(n11782), .B(n11781), .S(n11808), .Z(n11783) );
  OAI33_X1 U14245 ( .A1(n12441), .A2(n12700), .A3(n11808), .B1(n12459), .B2(
        n11784), .B3(n11783), .ZN(n11790) );
  INV_X1 U14246 ( .A(n11785), .ZN(n11788) );
  AOI21_X1 U14247 ( .B1(n12445), .B2(n11786), .A(n11788), .ZN(n11787) );
  MUX2_X1 U14248 ( .A(n11788), .B(n11787), .S(n11808), .Z(n11789) );
  INV_X1 U14249 ( .A(n11791), .ZN(n11794) );
  INV_X1 U14250 ( .A(n11792), .ZN(n11793) );
  MUX2_X1 U14251 ( .A(n11794), .B(n11793), .S(n11808), .Z(n11795) );
  NAND2_X1 U14252 ( .A1(n11797), .A2(n11796), .ZN(n12417) );
  INV_X1 U14253 ( .A(n11796), .ZN(n11799) );
  INV_X1 U14254 ( .A(n11797), .ZN(n11798) );
  MUX2_X1 U14255 ( .A(n11799), .B(n11798), .S(n11808), .Z(n11801) );
  INV_X1 U14256 ( .A(n11835), .ZN(n11805) );
  OAI22_X1 U14257 ( .A1(n11805), .A2(n11804), .B1(n11803), .B2(n11802), .ZN(
        n11806) );
  AND3_X1 U14258 ( .A1(n11811), .A2(n11810), .A3(n11809), .ZN(n11812) );
  OAI21_X1 U14259 ( .B1(n11812), .B2(n11838), .A(n11839), .ZN(n11844) );
  INV_X1 U14260 ( .A(n11844), .ZN(n11842) );
  INV_X1 U14261 ( .A(n11813), .ZN(n11826) );
  AND2_X1 U14262 ( .A1(n11815), .A2(n11814), .ZN(n11818) );
  INV_X1 U14263 ( .A(n15102), .ZN(n11816) );
  NAND4_X1 U14264 ( .A1(n11818), .A2(n15085), .A3(n11817), .A4(n11816), .ZN(
        n11824) );
  NAND4_X1 U14265 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11823) );
  NOR3_X1 U14266 ( .A1(n11824), .A2(n11823), .A3(n12603), .ZN(n11825) );
  NAND4_X1 U14267 ( .A1(n12594), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11828) );
  NOR4_X1 U14268 ( .A1(n11830), .A2(n11829), .A3(n12583), .A4(n11828), .ZN(
        n11831) );
  NAND3_X1 U14269 ( .A1(n12525), .A2(n12559), .A3(n11831), .ZN(n11832) );
  OR4_X1 U14270 ( .A1(n12467), .A2(n12479), .A3(n12519), .A4(n11832), .ZN(
        n11833) );
  NOR3_X1 U14271 ( .A1(n12494), .A2(n12459), .A3(n11833), .ZN(n11834) );
  INV_X1 U14272 ( .A(n11838), .ZN(n11840) );
  NOR2_X1 U14273 ( .A1(n11847), .A2(n11846), .ZN(n11850) );
  OAI21_X1 U14274 ( .B1(n11848), .B2(n11851), .A(P3_B_REG_SCAN_IN), .ZN(n11849) );
  INV_X1 U14275 ( .A(n13462), .ZN(n13288) );
  OAI222_X1 U14276 ( .A1(n14252), .A2(n13463), .B1(P1_U3086), .B2(n11852), 
        .C1(n10724), .C2(n13288), .ZN(P1_U3326) );
  AOI22_X1 U14277 ( .A1(n14188), .A2(n11967), .B1(n11930), .B2(n13737), .ZN(
        n11901) );
  INV_X1 U14278 ( .A(n11901), .ZN(n11904) );
  AOI22_X1 U14279 ( .A1(n14188), .A2(n11966), .B1(n11967), .B2(n13737), .ZN(
        n11854) );
  XNOR2_X1 U14280 ( .A(n11854), .B(n11853), .ZN(n11902) );
  INV_X1 U14281 ( .A(n11902), .ZN(n11903) );
  AND2_X1 U14282 ( .A1(n11930), .A2(n13742), .ZN(n11860) );
  AOI21_X1 U14283 ( .B1(n14559), .B2(n11932), .A(n11860), .ZN(n11867) );
  AOI22_X1 U14284 ( .A1(n14559), .A2(n11966), .B1(n11932), .B2(n13742), .ZN(
        n11861) );
  XNOR2_X1 U14285 ( .A(n11861), .B(n11853), .ZN(n11866) );
  XOR2_X1 U14286 ( .A(n11867), .B(n11866), .Z(n14554) );
  NAND2_X1 U14287 ( .A1(n14575), .A2(n11966), .ZN(n11863) );
  NAND2_X1 U14288 ( .A1(n13741), .A2(n11932), .ZN(n11862) );
  NAND2_X1 U14289 ( .A1(n11863), .A2(n11862), .ZN(n11864) );
  XNOR2_X1 U14290 ( .A(n11864), .B(n11853), .ZN(n11873) );
  AND2_X1 U14291 ( .A1(n11930), .A2(n13741), .ZN(n11865) );
  AOI21_X1 U14292 ( .B1(n14575), .B2(n11932), .A(n11865), .ZN(n11871) );
  XNOR2_X1 U14293 ( .A(n11873), .B(n11871), .ZN(n14566) );
  INV_X1 U14294 ( .A(n11866), .ZN(n11869) );
  INV_X1 U14295 ( .A(n11867), .ZN(n11868) );
  NAND2_X1 U14296 ( .A1(n11869), .A2(n11868), .ZN(n14567) );
  INV_X1 U14297 ( .A(n11871), .ZN(n11872) );
  AOI22_X1 U14298 ( .A1(n13601), .A2(n11966), .B1(n11932), .B2(n13740), .ZN(
        n11874) );
  XNOR2_X1 U14299 ( .A(n11874), .B(n11853), .ZN(n11875) );
  AOI22_X1 U14300 ( .A1(n13601), .A2(n11967), .B1(n11930), .B2(n13740), .ZN(
        n11876) );
  XNOR2_X1 U14301 ( .A(n11875), .B(n11876), .ZN(n13338) );
  INV_X1 U14302 ( .A(n11875), .ZN(n11878) );
  INV_X1 U14303 ( .A(n11876), .ZN(n11877) );
  OAI22_X1 U14304 ( .A1(n14582), .A2(n10324), .B1(n14536), .B2(n11979), .ZN(
        n11880) );
  XNOR2_X1 U14305 ( .A(n11880), .B(n11853), .ZN(n11889) );
  AND2_X1 U14306 ( .A1(n11930), .A2(n13739), .ZN(n11881) );
  AOI21_X1 U14307 ( .B1(n13607), .B2(n11932), .A(n11881), .ZN(n11887) );
  XNOR2_X1 U14308 ( .A(n11889), .B(n11887), .ZN(n13391) );
  NAND2_X1 U14309 ( .A1(n14546), .A2(n11966), .ZN(n11883) );
  OR2_X1 U14310 ( .A1(n11885), .A2(n11979), .ZN(n11882) );
  NAND2_X1 U14311 ( .A1(n11883), .A2(n11882), .ZN(n11884) );
  XNOR2_X1 U14312 ( .A(n11884), .B(n11853), .ZN(n11890) );
  NOR2_X1 U14313 ( .A1(n11885), .A2(n11978), .ZN(n11886) );
  AOI21_X1 U14314 ( .B1(n14546), .B2(n11932), .A(n11886), .ZN(n11891) );
  XNOR2_X1 U14315 ( .A(n11890), .B(n11891), .ZN(n14538) );
  INV_X1 U14316 ( .A(n11887), .ZN(n11888) );
  NAND2_X1 U14317 ( .A1(n11889), .A2(n11888), .ZN(n14539) );
  INV_X1 U14318 ( .A(n11890), .ZN(n11892) );
  NAND2_X1 U14319 ( .A1(n11892), .A2(n11891), .ZN(n11893) );
  NAND2_X1 U14320 ( .A1(n13612), .A2(n11966), .ZN(n11895) );
  NAND2_X1 U14321 ( .A1(n14086), .A2(n11932), .ZN(n11894) );
  NAND2_X1 U14322 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  XNOR2_X1 U14323 ( .A(n11896), .B(n11853), .ZN(n11897) );
  OAI22_X1 U14324 ( .A1(n13435), .A2(n11979), .B1(n14537), .B2(n11978), .ZN(
        n13426) );
  INV_X1 U14325 ( .A(n11897), .ZN(n11898) );
  OR2_X1 U14326 ( .A1(n11899), .A2(n11898), .ZN(n11900) );
  XNOR2_X1 U14327 ( .A(n11902), .B(n11901), .ZN(n13360) );
  OAI22_X1 U14328 ( .A1(n14181), .A2(n11979), .B1(n13628), .B2(n11978), .ZN(
        n11906) );
  OAI22_X1 U14329 ( .A1(n14181), .A2(n10324), .B1(n13628), .B2(n11979), .ZN(
        n11905) );
  XNOR2_X1 U14330 ( .A(n11905), .B(n11853), .ZN(n11907) );
  XOR2_X1 U14331 ( .A(n11906), .B(n11907), .Z(n13368) );
  INV_X1 U14332 ( .A(n14175), .ZN(n14068) );
  OAI22_X1 U14333 ( .A1(n14068), .A2(n11979), .B1(n13372), .B2(n11978), .ZN(
        n11913) );
  NAND2_X1 U14334 ( .A1(n14175), .A2(n11966), .ZN(n11910) );
  NAND2_X1 U14335 ( .A1(n13736), .A2(n11967), .ZN(n11909) );
  NAND2_X1 U14336 ( .A1(n11910), .A2(n11909), .ZN(n11911) );
  XNOR2_X1 U14337 ( .A(n11911), .B(n11853), .ZN(n11912) );
  XOR2_X1 U14338 ( .A(n11913), .B(n11912), .Z(n13407) );
  INV_X1 U14339 ( .A(n11912), .ZN(n11915) );
  INV_X1 U14340 ( .A(n11913), .ZN(n11914) );
  AOI22_X1 U14341 ( .A1(n14043), .A2(n11967), .B1(n11930), .B2(n13735), .ZN(
        n11918) );
  AOI22_X1 U14342 ( .A1(n14043), .A2(n11966), .B1(n11932), .B2(n13735), .ZN(
        n11916) );
  XNOR2_X1 U14343 ( .A(n11916), .B(n11853), .ZN(n11917) );
  XOR2_X1 U14344 ( .A(n11918), .B(n11917), .Z(n13323) );
  INV_X1 U14345 ( .A(n11917), .ZN(n11920) );
  INV_X1 U14346 ( .A(n11918), .ZN(n11919) );
  NAND2_X1 U14347 ( .A1(n11920), .A2(n11919), .ZN(n11921) );
  OAI22_X1 U14348 ( .A1(n14028), .A2(n11979), .B1(n13522), .B2(n11978), .ZN(
        n11923) );
  OAI22_X1 U14349 ( .A1(n14028), .A2(n10324), .B1(n13522), .B2(n11979), .ZN(
        n11922) );
  XNOR2_X1 U14350 ( .A(n11922), .B(n11853), .ZN(n11924) );
  XOR2_X1 U14351 ( .A(n11923), .B(n11924), .Z(n13385) );
  NAND2_X1 U14352 ( .A1(n11924), .A2(n11923), .ZN(n11925) );
  AOI22_X1 U14353 ( .A1(n14010), .A2(n11966), .B1(n11932), .B2(n13733), .ZN(
        n11926) );
  XNOR2_X1 U14354 ( .A(n11926), .B(n11853), .ZN(n11928) );
  AOI22_X1 U14355 ( .A1(n14010), .A2(n11967), .B1(n11930), .B2(n13733), .ZN(
        n11927) );
  XNOR2_X1 U14356 ( .A(n11928), .B(n11927), .ZN(n13330) );
  OAI22_X1 U14357 ( .A1(n7363), .A2(n10324), .B1(n13331), .B2(n11979), .ZN(
        n11929) );
  XNOR2_X1 U14358 ( .A(n11929), .B(n11853), .ZN(n11933) );
  AND2_X1 U14359 ( .A1(n11930), .A2(n13982), .ZN(n11931) );
  AOI21_X1 U14360 ( .B1(n13997), .B2(n11932), .A(n11931), .ZN(n11934) );
  XNOR2_X1 U14361 ( .A(n11933), .B(n11934), .ZN(n13400) );
  INV_X1 U14362 ( .A(n11933), .ZN(n11935) );
  NAND2_X1 U14363 ( .A1(n11935), .A2(n11934), .ZN(n11936) );
  NAND2_X1 U14364 ( .A1(n13398), .A2(n11936), .ZN(n13315) );
  OAI22_X1 U14365 ( .A1(n14142), .A2(n11979), .B1(n13990), .B2(n11978), .ZN(
        n11941) );
  NAND2_X1 U14366 ( .A1(n13978), .A2(n11966), .ZN(n11938) );
  NAND2_X1 U14367 ( .A1(n13732), .A2(n11932), .ZN(n11937) );
  NAND2_X1 U14368 ( .A1(n11938), .A2(n11937), .ZN(n11939) );
  XNOR2_X1 U14369 ( .A(n11939), .B(n11853), .ZN(n11940) );
  XOR2_X1 U14370 ( .A(n11941), .B(n11940), .Z(n13316) );
  INV_X1 U14371 ( .A(n11940), .ZN(n11943) );
  INV_X1 U14372 ( .A(n11941), .ZN(n11942) );
  NAND2_X1 U14373 ( .A1(n11943), .A2(n11942), .ZN(n11944) );
  OAI22_X1 U14374 ( .A1(n11616), .A2(n11979), .B1(n13352), .B2(n11978), .ZN(
        n11948) );
  NAND2_X1 U14375 ( .A1(n13961), .A2(n11966), .ZN(n11946) );
  NAND2_X1 U14376 ( .A1(n13983), .A2(n11967), .ZN(n11945) );
  NAND2_X1 U14377 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  XNOR2_X1 U14378 ( .A(n11947), .B(n11853), .ZN(n11949) );
  XOR2_X1 U14379 ( .A(n11948), .B(n11949), .Z(n13378) );
  NAND2_X1 U14380 ( .A1(n13943), .A2(n11966), .ZN(n11951) );
  NAND2_X1 U14381 ( .A1(n13731), .A2(n11932), .ZN(n11950) );
  NAND2_X1 U14382 ( .A1(n11951), .A2(n11950), .ZN(n11952) );
  XNOR2_X1 U14383 ( .A(n11952), .B(n11853), .ZN(n11954) );
  OAI22_X1 U14384 ( .A1(n11953), .A2(n11979), .B1(n13953), .B2(n11978), .ZN(
        n11955) );
  XNOR2_X1 U14385 ( .A(n11954), .B(n11955), .ZN(n13350) );
  INV_X1 U14386 ( .A(n11954), .ZN(n11957) );
  INV_X1 U14387 ( .A(n11955), .ZN(n11956) );
  NAND2_X1 U14388 ( .A1(n11957), .A2(n11956), .ZN(n11958) );
  OAI22_X1 U14389 ( .A1(n13417), .A2(n11979), .B1(n13310), .B2(n11978), .ZN(
        n11963) );
  NAND2_X1 U14390 ( .A1(n13928), .A2(n11966), .ZN(n11960) );
  NAND2_X1 U14391 ( .A1(n13934), .A2(n11967), .ZN(n11959) );
  NAND2_X1 U14392 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  XNOR2_X1 U14393 ( .A(n11961), .B(n11853), .ZN(n11962) );
  XOR2_X1 U14394 ( .A(n11963), .B(n11962), .Z(n13416) );
  INV_X1 U14395 ( .A(n11962), .ZN(n11965) );
  INV_X1 U14396 ( .A(n11963), .ZN(n11964) );
  INV_X1 U14397 ( .A(n13903), .ZN(n13913) );
  OAI22_X1 U14398 ( .A1(n13877), .A2(n11979), .B1(n13913), .B2(n11978), .ZN(
        n11972) );
  NAND2_X1 U14399 ( .A1(n14115), .A2(n11966), .ZN(n11969) );
  NAND2_X1 U14400 ( .A1(n13903), .A2(n11967), .ZN(n11968) );
  NAND2_X1 U14401 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  XNOR2_X1 U14402 ( .A(n11970), .B(n11853), .ZN(n11971) );
  XOR2_X1 U14403 ( .A(n11972), .B(n11971), .Z(n13307) );
  INV_X1 U14404 ( .A(n11971), .ZN(n11974) );
  INV_X1 U14405 ( .A(n11972), .ZN(n11973) );
  NAND2_X1 U14406 ( .A1(n11975), .A2(n13461), .ZN(n11977) );
  OR2_X1 U14407 ( .A1(n13464), .A2(n14242), .ZN(n11976) );
  OAI22_X1 U14408 ( .A1(n13860), .A2(n10324), .B1(n13878), .B2(n11979), .ZN(
        n11982) );
  OAI22_X1 U14409 ( .A1(n13860), .A2(n11979), .B1(n13878), .B2(n11978), .ZN(
        n11980) );
  XNOR2_X1 U14410 ( .A(n11980), .B(n11853), .ZN(n11981) );
  XOR2_X1 U14411 ( .A(n11982), .B(n11981), .Z(n11983) );
  XNOR2_X1 U14412 ( .A(n11984), .B(n11983), .ZN(n11994) );
  NOR2_X1 U14413 ( .A1(n14580), .A2(n13906), .ZN(n11992) );
  NAND2_X1 U14414 ( .A1(n6688), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n11989) );
  NAND2_X1 U14415 ( .A1(n13450), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11988) );
  OR2_X1 U14416 ( .A1(n6465), .A2(n13886), .ZN(n11987) );
  INV_X1 U14417 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n11985) );
  OR2_X1 U14418 ( .A1(n13453), .A2(n11985), .ZN(n11986) );
  NAND4_X1 U14419 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n13902) );
  AOI22_X1 U14420 ( .A1(n13418), .A2(n13902), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11990) );
  OAI21_X1 U14421 ( .B1(n13913), .B2(n14562), .A(n11990), .ZN(n11991) );
  AOI211_X1 U14422 ( .C1(n14111), .C2(n14576), .A(n11992), .B(n11991), .ZN(
        n11993) );
  OAI21_X1 U14423 ( .B1(n11994), .B2(n14570), .A(n11993), .ZN(P1_U3220) );
  OAI222_X1 U14424 ( .A1(n14252), .A2(n6752), .B1(n10724), .B2(n11995), .C1(
        P1_U3086), .C2(n13440), .ZN(P1_U3334) );
  OAI222_X1 U14425 ( .A1(P3_U3151), .A2(n11998), .B1(n12747), .B2(n11997), 
        .C1(n11996), .C2(n12744), .ZN(P3_U3265) );
  NOR2_X1 U14426 ( .A1(n12130), .A2(n12409), .ZN(n12003) );
  INV_X1 U14427 ( .A(n12000), .ZN(n12405) );
  AOI22_X1 U14428 ( .A1(n12405), .A2(n12128), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12001) );
  OAI21_X1 U14429 ( .B1(n12433), .B2(n12126), .A(n12001), .ZN(n12002) );
  AOI211_X1 U14430 ( .C1(n12412), .C2(n12132), .A(n12003), .B(n12002), .ZN(
        n12004) );
  INV_X1 U14431 ( .A(n12005), .ZN(n12725) );
  OAI211_X1 U14432 ( .C1(n12008), .C2(n12007), .A(n12006), .B(n6997), .ZN(
        n12013) );
  INV_X1 U14433 ( .A(n12009), .ZN(n12585) );
  NAND2_X1 U14434 ( .A1(n12140), .A2(n12107), .ZN(n12010) );
  NAND2_X1 U14435 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n15036)
         );
  OAI211_X1 U14436 ( .C1(n12582), .C2(n12109), .A(n12010), .B(n15036), .ZN(
        n12011) );
  AOI21_X1 U14437 ( .B1(n12585), .B2(n12117), .A(n12011), .ZN(n12012) );
  OAI211_X1 U14438 ( .C1(n12725), .C2(n12114), .A(n12013), .B(n12012), .ZN(
        P3_U3155) );
  XNOR2_X1 U14439 ( .A(n12076), .B(n12075), .ZN(n12077) );
  XNOR2_X1 U14440 ( .A(n12077), .B(n12471), .ZN(n12021) );
  OAI22_X1 U14441 ( .A1(n12482), .A2(n12126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12014), .ZN(n12015) );
  AOI21_X1 U14442 ( .B1(n12128), .B2(n12137), .A(n12015), .ZN(n12016) );
  OAI21_X1 U14443 ( .B1(n12130), .B2(n12017), .A(n12016), .ZN(n12018) );
  AOI21_X1 U14444 ( .B1(n12019), .B2(n12132), .A(n12018), .ZN(n12020) );
  OAI21_X1 U14445 ( .B1(n12021), .B2(n12134), .A(n12020), .ZN(P3_U3156) );
  OAI211_X1 U14446 ( .C1(n12024), .C2(n12023), .A(n12022), .B(n6997), .ZN(
        n12028) );
  NAND2_X1 U14447 ( .A1(P3_U3151), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n12365)
         );
  OAI21_X1 U14448 ( .B1(n12511), .B2(n12126), .A(n12365), .ZN(n12026) );
  NOR2_X1 U14449 ( .A1(n12130), .A2(n12515), .ZN(n12025) );
  AOI211_X1 U14450 ( .C1(n12128), .C2(n12139), .A(n12026), .B(n12025), .ZN(
        n12027) );
  OAI211_X1 U14451 ( .C1(n12114), .C2(n12713), .A(n12028), .B(n12027), .ZN(
        P3_U3159) );
  MUX2_X1 U14452 ( .A(n12030), .B(n12146), .S(n12029), .Z(n12032) );
  XNOR2_X1 U14453 ( .A(n12032), .B(n12031), .ZN(n12033) );
  NAND2_X1 U14454 ( .A1(n12033), .A2(n6997), .ZN(n12040) );
  AOI21_X1 U14455 ( .B1(n12146), .B2(n12107), .A(n12034), .ZN(n12039) );
  AOI22_X1 U14456 ( .A1(n12132), .A2(n12035), .B1(n12128), .B2(n12144), .ZN(
        n12038) );
  NAND2_X1 U14457 ( .A1(n12117), .A2(n12036), .ZN(n12037) );
  NAND4_X1 U14458 ( .A1(n12040), .A2(n12039), .A3(n12038), .A4(n12037), .ZN(
        P3_U3161) );
  OAI211_X1 U14459 ( .C1(n12043), .C2(n12042), .A(n12041), .B(n6997), .ZN(
        n12048) );
  INV_X1 U14460 ( .A(n12044), .ZN(n12483) );
  AOI22_X1 U14461 ( .A1(n12139), .A2(n12107), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12045) );
  OAI21_X1 U14462 ( .B1(n12482), .B2(n12109), .A(n12045), .ZN(n12046) );
  AOI21_X1 U14463 ( .B1(n12483), .B2(n12117), .A(n12046), .ZN(n12047) );
  OAI211_X1 U14464 ( .C1(n12708), .C2(n12114), .A(n12048), .B(n12047), .ZN(
        P3_U3163) );
  XOR2_X1 U14465 ( .A(n12051), .B(n12050), .Z(n12056) );
  AOI22_X1 U14466 ( .A1(n12107), .A2(n12137), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12053) );
  NAND2_X1 U14467 ( .A1(n12404), .A2(n12128), .ZN(n12052) );
  OAI211_X1 U14468 ( .C1(n12130), .C2(n12429), .A(n12053), .B(n12052), .ZN(
        n12054) );
  AOI21_X1 U14469 ( .B1(n12631), .B2(n12132), .A(n12054), .ZN(n12055) );
  OAI21_X1 U14470 ( .B1(n12056), .B2(n12134), .A(n12055), .ZN(P3_U3165) );
  XNOR2_X1 U14471 ( .A(n12057), .B(n12070), .ZN(n12058) );
  XNOR2_X1 U14472 ( .A(n6454), .B(n12058), .ZN(n12065) );
  NAND2_X1 U14473 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n14429)
         );
  OAI21_X1 U14474 ( .B1(n12582), .B2(n12126), .A(n14429), .ZN(n12060) );
  AOI21_X1 U14475 ( .B1(n12128), .B2(n12557), .A(n12060), .ZN(n12061) );
  OAI21_X1 U14476 ( .B1(n12130), .B2(n12062), .A(n12061), .ZN(n12063) );
  AOI21_X1 U14477 ( .B1(n12670), .B2(n12132), .A(n12063), .ZN(n12064) );
  OAI21_X1 U14478 ( .B1(n12065), .B2(n12134), .A(n12064), .ZN(P3_U3166) );
  AOI21_X1 U14479 ( .B1(n12067), .B2(n12066), .A(n12134), .ZN(n12069) );
  NAND2_X1 U14480 ( .A1(n12069), .A2(n12068), .ZN(n12074) );
  NAND2_X1 U14481 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n14447)
         );
  OAI21_X1 U14482 ( .B1(n12070), .B2(n12126), .A(n14447), .ZN(n12072) );
  NOR2_X1 U14483 ( .A1(n12130), .A2(n12547), .ZN(n12071) );
  AOI211_X1 U14484 ( .C1(n12128), .C2(n12543), .A(n12072), .B(n12071), .ZN(
        n12073) );
  OAI211_X1 U14485 ( .C1(n12546), .C2(n12114), .A(n12074), .B(n12073), .ZN(
        P3_U3168) );
  OAI22_X1 U14486 ( .A1(n12077), .A2(n12441), .B1(n12076), .B2(n12075), .ZN(
        n12080) );
  XNOR2_X1 U14487 ( .A(n12078), .B(n12137), .ZN(n12079) );
  XNOR2_X1 U14488 ( .A(n12080), .B(n12079), .ZN(n12087) );
  OAI22_X1 U14489 ( .A1(n12471), .A2(n12126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12081), .ZN(n12082) );
  AOI21_X1 U14490 ( .B1(n12128), .B2(n12442), .A(n12082), .ZN(n12083) );
  OAI21_X1 U14491 ( .B1(n12130), .B2(n12449), .A(n12083), .ZN(n12084) );
  AOI21_X1 U14492 ( .B1(n12085), .B2(n12132), .A(n12084), .ZN(n12086) );
  OAI21_X1 U14493 ( .B1(n12087), .B2(n12134), .A(n12086), .ZN(P3_U3169) );
  OAI211_X1 U14494 ( .C1(n12090), .C2(n12089), .A(n12088), .B(n6997), .ZN(
        n12095) );
  OAI22_X1 U14495 ( .A1(n12528), .A2(n12126), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12091), .ZN(n12093) );
  NOR2_X1 U14496 ( .A1(n12130), .A2(n12502), .ZN(n12092) );
  AOI211_X1 U14497 ( .C1(n12128), .C2(n12499), .A(n12093), .B(n12092), .ZN(
        n12094) );
  OAI211_X1 U14498 ( .C1(n12651), .C2(n12114), .A(n12095), .B(n12094), .ZN(
        P3_U3173) );
  XNOR2_X1 U14499 ( .A(n6459), .B(n12138), .ZN(n12102) );
  INV_X1 U14500 ( .A(n12097), .ZN(n12473) );
  NAND2_X1 U14501 ( .A1(n12117), .A2(n12473), .ZN(n12099) );
  AOI22_X1 U14502 ( .A1(n12499), .A2(n12107), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12098) );
  OAI211_X1 U14503 ( .C1(n12471), .C2(n12109), .A(n12099), .B(n12098), .ZN(
        n12100) );
  AOI21_X1 U14504 ( .B1(n12472), .B2(n12132), .A(n12100), .ZN(n12101) );
  OAI21_X1 U14505 ( .B1(n12102), .B2(n12134), .A(n12101), .ZN(P3_U3175) );
  INV_X1 U14506 ( .A(n12539), .ZN(n12717) );
  OAI211_X1 U14507 ( .C1(n12105), .C2(n12104), .A(n12103), .B(n6997), .ZN(
        n12113) );
  INV_X1 U14508 ( .A(n12529), .ZN(n12111) );
  NOR2_X1 U14509 ( .A1(n12106), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12350) );
  AOI21_X1 U14510 ( .B1(n12107), .B2(n12557), .A(n12350), .ZN(n12108) );
  OAI21_X1 U14511 ( .B1(n12528), .B2(n12109), .A(n12108), .ZN(n12110) );
  AOI21_X1 U14512 ( .B1(n12111), .B2(n12117), .A(n12110), .ZN(n12112) );
  OAI211_X1 U14513 ( .C1(n12717), .C2(n12114), .A(n12113), .B(n12112), .ZN(
        P3_U3178) );
  NAND2_X1 U14514 ( .A1(n12117), .A2(n12423), .ZN(n12119) );
  AOI22_X1 U14515 ( .A1(n12128), .A2(n12388), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12118) );
  OAI211_X1 U14516 ( .C1(n12421), .C2(n12126), .A(n12119), .B(n12118), .ZN(
        n12120) );
  AOI21_X1 U14517 ( .B1(n12422), .B2(n12132), .A(n12120), .ZN(n12121) );
  OAI21_X1 U14518 ( .B1(n12122), .B2(n12134), .A(n12121), .ZN(P3_U3180) );
  XNOR2_X1 U14519 ( .A(n12123), .B(n12556), .ZN(n12124) );
  XNOR2_X1 U14520 ( .A(n12125), .B(n12124), .ZN(n12135) );
  NAND2_X1 U14521 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14414)
         );
  OAI21_X1 U14522 ( .B1(n12597), .B2(n12126), .A(n14414), .ZN(n12127) );
  AOI21_X1 U14523 ( .B1(n12128), .B2(n12572), .A(n12127), .ZN(n12129) );
  OAI21_X1 U14524 ( .B1(n12130), .B2(n12574), .A(n12129), .ZN(n12131) );
  AOI21_X1 U14525 ( .B1(n12674), .B2(n12132), .A(n12131), .ZN(n12133) );
  OAI21_X1 U14526 ( .B1(n12135), .B2(n12134), .A(n12133), .ZN(P3_U3181) );
  MUX2_X1 U14527 ( .A(P3_DATAO_REG_31__SCAN_IN), .B(n14458), .S(P3_U3897), .Z(
        P3_U3522) );
  MUX2_X1 U14528 ( .A(P3_DATAO_REG_30__SCAN_IN), .B(n12136), .S(P3_U3897), .Z(
        P3_U3521) );
  MUX2_X1 U14529 ( .A(P3_DATAO_REG_29__SCAN_IN), .B(n12389), .S(P3_U3897), .Z(
        P3_U3520) );
  MUX2_X1 U14530 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12405), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14531 ( .A(P3_DATAO_REG_27__SCAN_IN), .B(n12388), .S(P3_U3897), .Z(
        P3_U3518) );
  MUX2_X1 U14532 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12404), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14533 ( .A(P3_DATAO_REG_25__SCAN_IN), .B(n12442), .S(P3_U3897), .Z(
        P3_U3516) );
  MUX2_X1 U14534 ( .A(P3_DATAO_REG_24__SCAN_IN), .B(n12137), .S(P3_U3897), .Z(
        P3_U3515) );
  MUX2_X1 U14535 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12441), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14536 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12138), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14537 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12499), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14538 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12139), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14539 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12498), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14540 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12543), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14541 ( .A(P3_DATAO_REG_17__SCAN_IN), .B(n12557), .S(P3_U3897), .Z(
        P3_U3508) );
  MUX2_X1 U14542 ( .A(P3_DATAO_REG_16__SCAN_IN), .B(n12572), .S(P3_U3897), .Z(
        P3_U3507) );
  MUX2_X1 U14543 ( .A(P3_DATAO_REG_15__SCAN_IN), .B(n12556), .S(P3_U3897), .Z(
        P3_U3506) );
  MUX2_X1 U14544 ( .A(P3_DATAO_REG_14__SCAN_IN), .B(n12570), .S(P3_U3897), .Z(
        P3_U3505) );
  MUX2_X1 U14545 ( .A(P3_DATAO_REG_13__SCAN_IN), .B(n12140), .S(P3_U3897), .Z(
        P3_U3504) );
  MUX2_X1 U14546 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n12141), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U14547 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12142), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14548 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12143), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14549 ( .A(P3_DATAO_REG_9__SCAN_IN), .B(n12144), .S(n12284), .Z(
        P3_U3500) );
  MUX2_X1 U14550 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12145), .S(n12284), .Z(
        P3_U3499) );
  MUX2_X1 U14551 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12146), .S(n12284), .Z(
        P3_U3498) );
  MUX2_X1 U14552 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n12147), .S(n12284), .Z(
        P3_U3497) );
  MUX2_X1 U14553 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12148), .S(n12284), .Z(
        P3_U3496) );
  MUX2_X1 U14554 ( .A(P3_DATAO_REG_3__SCAN_IN), .B(n12149), .S(n12284), .Z(
        n12282) );
  NOR4_X1 U14555 ( .A1(keyinput13), .A2(keyinput9), .A3(keyinput5), .A4(
        keyinput1), .ZN(n12153) );
  NOR4_X1 U14556 ( .A1(keyinput21), .A2(keyinput24), .A3(keyinput40), .A4(
        keyinput60), .ZN(n12152) );
  NOR4_X1 U14557 ( .A1(keyinput52), .A2(keyinput32), .A3(keyinput38), .A4(
        keyinput59), .ZN(n12151) );
  NOR4_X1 U14558 ( .A1(keyinput51), .A2(keyinput26), .A3(keyinput30), .A4(
        keyinput18), .ZN(n12150) );
  NAND4_X1 U14559 ( .A1(n12153), .A2(n12152), .A3(n12151), .A4(n12150), .ZN(
        n12201) );
  NOR2_X1 U14560 ( .A1(keyinput62), .A2(keyinput22), .ZN(n12154) );
  NAND3_X1 U14561 ( .A1(keyinput42), .A2(keyinput36), .A3(n12154), .ZN(n12159)
         );
  NAND3_X1 U14562 ( .A1(keyinput48), .A2(keyinput14), .A3(keyinput25), .ZN(
        n12158) );
  NOR3_X1 U14563 ( .A1(keyinput20), .A2(keyinput10), .A3(keyinput39), .ZN(
        n12156) );
  NOR3_X1 U14564 ( .A1(keyinput31), .A2(keyinput44), .A3(keyinput4), .ZN(
        n12155) );
  NAND4_X1 U14565 ( .A1(keyinput16), .A2(n12156), .A3(keyinput41), .A4(n12155), 
        .ZN(n12157) );
  NOR4_X1 U14566 ( .A1(keyinput7), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12173) );
  NAND2_X1 U14567 ( .A1(keyinput47), .A2(keyinput17), .ZN(n12160) );
  NOR3_X1 U14568 ( .A1(keyinput12), .A2(keyinput0), .A3(n12160), .ZN(n12172)
         );
  NAND2_X1 U14569 ( .A1(keyinput34), .A2(keyinput54), .ZN(n12165) );
  NOR3_X1 U14570 ( .A1(keyinput53), .A2(keyinput27), .A3(keyinput57), .ZN(
        n12163) );
  INV_X1 U14571 ( .A(keyinput29), .ZN(n12161) );
  NOR3_X1 U14572 ( .A1(keyinput8), .A2(keyinput50), .A3(n12161), .ZN(n12162)
         );
  NAND4_X1 U14573 ( .A1(keyinput43), .A2(n12163), .A3(keyinput2), .A4(n12162), 
        .ZN(n12164) );
  NOR4_X1 U14574 ( .A1(keyinput49), .A2(keyinput6), .A3(n12165), .A4(n12164), 
        .ZN(n12171) );
  NAND4_X1 U14575 ( .A1(keyinput37), .A2(keyinput45), .A3(keyinput33), .A4(
        keyinput61), .ZN(n12169) );
  NAND4_X1 U14576 ( .A1(keyinput28), .A2(keyinput56), .A3(keyinput35), .A4(
        keyinput46), .ZN(n12168) );
  NAND4_X1 U14577 ( .A1(keyinput58), .A2(keyinput55), .A3(keyinput63), .A4(
        keyinput11), .ZN(n12167) );
  NAND4_X1 U14578 ( .A1(keyinput15), .A2(keyinput3), .A3(keyinput23), .A4(
        keyinput19), .ZN(n12166) );
  NOR4_X1 U14579 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12170) );
  NAND4_X1 U14580 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12200) );
  AOI22_X1 U14581 ( .A1(n15017), .A2(keyinput51), .B1(n12175), .B2(keyinput33), 
        .ZN(n12174) );
  OAI221_X1 U14582 ( .B1(n15017), .B2(keyinput51), .C1(n12175), .C2(keyinput33), .A(n12174), .ZN(n12184) );
  AOI22_X1 U14583 ( .A1(n12177), .A2(keyinput45), .B1(keyinput46), .B2(n8418), 
        .ZN(n12176) );
  OAI221_X1 U14584 ( .B1(n12177), .B2(keyinput45), .C1(n8418), .C2(keyinput46), 
        .A(n12176), .ZN(n12183) );
  AOI22_X1 U14585 ( .A1(n12613), .A2(keyinput52), .B1(keyinput19), .B2(n12645), 
        .ZN(n12178) );
  OAI221_X1 U14586 ( .B1(n12613), .B2(keyinput52), .C1(n12645), .C2(keyinput19), .A(n12178), .ZN(n12182) );
  XOR2_X1 U14587 ( .A(n9362), .B(keyinput1), .Z(n12180) );
  XNOR2_X1 U14588 ( .A(P3_IR_REG_23__SCAN_IN), .B(keyinput28), .ZN(n12179) );
  NAND2_X1 U14589 ( .A1(n12180), .A2(n12179), .ZN(n12181) );
  NOR4_X1 U14590 ( .A1(n12184), .A2(n12183), .A3(n12182), .A4(n12181), .ZN(
        n12199) );
  INV_X1 U14591 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U14592 ( .A1(n12187), .A2(keyinput60), .B1(keyinput37), .B2(n12186), 
        .ZN(n12185) );
  OAI221_X1 U14593 ( .B1(n12187), .B2(keyinput60), .C1(n12186), .C2(keyinput37), .A(n12185), .ZN(n12197) );
  INV_X1 U14594 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n12188) );
  XNOR2_X1 U14595 ( .A(keyinput32), .B(n12188), .ZN(n12196) );
  XNOR2_X1 U14596 ( .A(keyinput3), .B(n12189), .ZN(n12195) );
  XNOR2_X1 U14597 ( .A(P2_IR_REG_12__SCAN_IN), .B(keyinput23), .ZN(n12193) );
  XNOR2_X1 U14598 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput18), .ZN(n12192)
         );
  XNOR2_X1 U14599 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput55), .ZN(n12191)
         );
  XNOR2_X1 U14600 ( .A(P3_IR_REG_10__SCAN_IN), .B(keyinput30), .ZN(n12190) );
  NAND4_X1 U14601 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12194) );
  NOR4_X1 U14602 ( .A1(n12197), .A2(n12196), .A3(n12195), .A4(n12194), .ZN(
        n12198) );
  OAI211_X1 U14603 ( .C1(n12201), .C2(n12200), .A(n12199), .B(n12198), .ZN(
        n12280) );
  INV_X1 U14604 ( .A(P1_D_REG_10__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U14605 ( .A1(n12203), .A2(keyinput20), .B1(n14695), .B2(keyinput16), 
        .ZN(n12202) );
  OAI221_X1 U14606 ( .B1(n12203), .B2(keyinput20), .C1(n14695), .C2(keyinput16), .A(n12202), .ZN(n12213) );
  AOI22_X1 U14607 ( .A1(n14601), .A2(keyinput10), .B1(n12205), .B2(keyinput39), 
        .ZN(n12204) );
  OAI221_X1 U14608 ( .B1(n14601), .B2(keyinput10), .C1(n12205), .C2(keyinput39), .A(n12204), .ZN(n12212) );
  INV_X1 U14609 ( .A(keyinput31), .ZN(n12207) );
  AOI22_X1 U14610 ( .A1(n8627), .A2(keyinput44), .B1(P3_DATAO_REG_1__SCAN_IN), 
        .B2(n12207), .ZN(n12206) );
  OAI221_X1 U14611 ( .B1(n8627), .B2(keyinput44), .C1(n12207), .C2(
        P3_DATAO_REG_1__SCAN_IN), .A(n12206), .ZN(n12211) );
  INV_X1 U14612 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n14847) );
  AOI22_X1 U14613 ( .A1(n12209), .A2(keyinput4), .B1(keyinput41), .B2(n14847), 
        .ZN(n12208) );
  OAI221_X1 U14614 ( .B1(n12209), .B2(keyinput4), .C1(n14847), .C2(keyinput41), 
        .A(n12208), .ZN(n12210) );
  NOR4_X1 U14615 ( .A1(n12213), .A2(n12212), .A3(n12211), .A4(n12210), .ZN(
        n12252) );
  AOI22_X1 U14616 ( .A1(n8305), .A2(keyinput36), .B1(keyinput22), .B2(n12215), 
        .ZN(n12214) );
  OAI221_X1 U14617 ( .B1(n8305), .B2(keyinput36), .C1(n12215), .C2(keyinput22), 
        .A(n12214), .ZN(n12224) );
  AOI22_X1 U14618 ( .A1(n12217), .A2(keyinput14), .B1(keyinput25), .B2(n13325), 
        .ZN(n12216) );
  OAI221_X1 U14619 ( .B1(n12217), .B2(keyinput14), .C1(n13325), .C2(keyinput25), .A(n12216), .ZN(n12223) );
  XNOR2_X1 U14620 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput62), .ZN(n12221) );
  XNOR2_X1 U14621 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(keyinput42), .ZN(n12220)
         );
  XNOR2_X1 U14622 ( .A(P3_IR_REG_15__SCAN_IN), .B(keyinput7), .ZN(n12219) );
  XNOR2_X1 U14623 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput48), .ZN(n12218) );
  NAND4_X1 U14624 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n12222) );
  NOR3_X1 U14625 ( .A1(n12224), .A2(n12223), .A3(n12222), .ZN(n12251) );
  AOI22_X1 U14626 ( .A1(n12227), .A2(keyinput27), .B1(keyinput57), .B2(n12226), 
        .ZN(n12225) );
  OAI221_X1 U14627 ( .B1(n12227), .B2(keyinput27), .C1(n12226), .C2(keyinput57), .A(n12225), .ZN(n12237) );
  XNOR2_X1 U14628 ( .A(n12228), .B(keyinput43), .ZN(n12236) );
  XNOR2_X1 U14629 ( .A(P3_REG1_REG_0__SCAN_IN), .B(keyinput17), .ZN(n12232) );
  XNOR2_X1 U14630 ( .A(P2_IR_REG_8__SCAN_IN), .B(keyinput47), .ZN(n12231) );
  XNOR2_X1 U14631 ( .A(P2_REG0_REG_28__SCAN_IN), .B(keyinput12), .ZN(n12230)
         );
  XNOR2_X1 U14632 ( .A(P2_IR_REG_3__SCAN_IN), .B(keyinput0), .ZN(n12229) );
  NAND4_X1 U14633 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12235) );
  XNOR2_X1 U14634 ( .A(n12233), .B(keyinput53), .ZN(n12234) );
  NOR4_X1 U14635 ( .A1(n12237), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n12250) );
  AOI22_X1 U14636 ( .A1(n12240), .A2(keyinput34), .B1(n12239), .B2(keyinput49), 
        .ZN(n12238) );
  OAI221_X1 U14637 ( .B1(n12240), .B2(keyinput34), .C1(n12239), .C2(keyinput49), .A(n12238), .ZN(n12248) );
  AOI22_X1 U14638 ( .A1(n7037), .A2(keyinput6), .B1(keyinput54), .B2(n9794), 
        .ZN(n12241) );
  OAI221_X1 U14639 ( .B1(n7037), .B2(keyinput6), .C1(n9794), .C2(keyinput54), 
        .A(n12241), .ZN(n12247) );
  INV_X1 U14640 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n14443) );
  AOI22_X1 U14641 ( .A1(n14443), .A2(keyinput8), .B1(keyinput2), .B2(n7818), 
        .ZN(n12242) );
  OAI221_X1 U14642 ( .B1(n14443), .B2(keyinput8), .C1(n7818), .C2(keyinput2), 
        .A(n12242), .ZN(n12246) );
  AOI22_X1 U14643 ( .A1(n12244), .A2(keyinput29), .B1(n8450), .B2(keyinput50), 
        .ZN(n12243) );
  OAI221_X1 U14644 ( .B1(n12244), .B2(keyinput29), .C1(n8450), .C2(keyinput50), 
        .A(n12243), .ZN(n12245) );
  NOR4_X1 U14645 ( .A1(n12248), .A2(n12247), .A3(n12246), .A4(n12245), .ZN(
        n12249) );
  NAND4_X1 U14646 ( .A1(n12252), .A2(n12251), .A3(n12250), .A4(n12249), .ZN(
        n12279) );
  INV_X1 U14647 ( .A(P1_D_REG_25__SCAN_IN), .ZN(n14680) );
  XNOR2_X1 U14648 ( .A(n14680), .B(keyinput58), .ZN(n12261) );
  XNOR2_X1 U14649 ( .A(n12253), .B(keyinput21), .ZN(n12260) );
  XNOR2_X1 U14650 ( .A(P1_STATE_REG_SCAN_IN), .B(keyinput15), .ZN(n12256) );
  XNOR2_X1 U14651 ( .A(SI_1_), .B(keyinput56), .ZN(n12255) );
  XNOR2_X1 U14652 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput9), .ZN(n12254) );
  NAND3_X1 U14653 ( .A1(n12256), .A2(n12255), .A3(n12254), .ZN(n12259) );
  XNOR2_X1 U14654 ( .A(n12257), .B(keyinput63), .ZN(n12258) );
  NOR4_X1 U14655 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12265) );
  OAI22_X1 U14656 ( .A1(n14251), .A2(keyinput24), .B1(n12263), .B2(keyinput11), 
        .ZN(n12262) );
  AOI221_X1 U14657 ( .B1(n14251), .B2(keyinput24), .C1(keyinput11), .C2(n12263), .A(n12262), .ZN(n12264) );
  NAND2_X1 U14658 ( .A1(n12265), .A2(n12264), .ZN(n12278) );
  INV_X1 U14659 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14287) );
  OAI22_X1 U14660 ( .A1(n12267), .A2(keyinput38), .B1(n14287), .B2(keyinput61), 
        .ZN(n12266) );
  AOI221_X1 U14661 ( .B1(n12267), .B2(keyinput38), .C1(keyinput61), .C2(n14287), .A(n12266), .ZN(n12276) );
  OAI22_X1 U14662 ( .A1(n12269), .A2(keyinput26), .B1(n10289), .B2(keyinput35), 
        .ZN(n12268) );
  AOI221_X1 U14663 ( .B1(n12269), .B2(keyinput26), .C1(keyinput35), .C2(n10289), .A(n12268), .ZN(n12275) );
  INV_X1 U14664 ( .A(P1_D_REG_24__SCAN_IN), .ZN(n14681) );
  OAI22_X1 U14665 ( .A1(n15119), .A2(keyinput13), .B1(n14681), .B2(keyinput40), 
        .ZN(n12270) );
  AOI221_X1 U14666 ( .B1(n15119), .B2(keyinput13), .C1(keyinput40), .C2(n14681), .A(n12270), .ZN(n12274) );
  INV_X1 U14667 ( .A(P1_D_REG_31__SCAN_IN), .ZN(n14674) );
  INV_X1 U14668 ( .A(keyinput5), .ZN(n12272) );
  OAI22_X1 U14669 ( .A1(n14674), .A2(keyinput59), .B1(n12272), .B2(
        P3_DATAO_REG_4__SCAN_IN), .ZN(n12271) );
  AOI221_X1 U14670 ( .B1(n14674), .B2(keyinput59), .C1(P3_DATAO_REG_4__SCAN_IN), .C2(n12272), .A(n12271), .ZN(n12273) );
  NAND4_X1 U14671 ( .A1(n12276), .A2(n12275), .A3(n12274), .A4(n12273), .ZN(
        n12277) );
  NOR4_X1 U14672 ( .A1(n12280), .A2(n12279), .A3(n12278), .A4(n12277), .ZN(
        n12281) );
  XOR2_X1 U14673 ( .A(n12282), .B(n12281), .Z(P3_U3494) );
  MUX2_X1 U14674 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12283), .S(n12284), .Z(
        P3_U3493) );
  MUX2_X1 U14675 ( .A(P3_DATAO_REG_0__SCAN_IN), .B(n12285), .S(n12284), .Z(
        P3_U3491) );
  MUX2_X1 U14676 ( .A(P3_REG2_REG_18__SCAN_IN), .B(P3_REG1_REG_18__SCAN_IN), 
        .S(n6717), .Z(n12312) );
  MUX2_X1 U14677 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n6717), .Z(n12310) );
  MUX2_X1 U14678 ( .A(P3_REG2_REG_16__SCAN_IN), .B(P3_REG1_REG_16__SCAN_IN), 
        .S(n6717), .Z(n12309) );
  NAND2_X1 U14679 ( .A1(n12287), .A2(n12286), .ZN(n12291) );
  INV_X1 U14680 ( .A(n12288), .ZN(n12289) );
  NAND2_X1 U14681 ( .A1(n12289), .A2(n12332), .ZN(n12290) );
  NAND2_X1 U14682 ( .A1(n12291), .A2(n12290), .ZN(n14975) );
  MUX2_X1 U14683 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n6717), .Z(n12292) );
  XNOR2_X1 U14684 ( .A(n12292), .B(n12333), .ZN(n14974) );
  NAND2_X1 U14685 ( .A1(n14975), .A2(n14974), .ZN(n12295) );
  INV_X1 U14686 ( .A(n12292), .ZN(n12293) );
  NAND2_X1 U14687 ( .A1(n12293), .A2(n12333), .ZN(n12294) );
  NAND2_X1 U14688 ( .A1(n12295), .A2(n12294), .ZN(n14991) );
  MUX2_X1 U14689 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n6717), .Z(n12296) );
  XNOR2_X1 U14690 ( .A(n12296), .B(n15001), .ZN(n14992) );
  OR2_X1 U14691 ( .A1(n14991), .A2(n14992), .ZN(n12298) );
  NAND2_X1 U14692 ( .A1(n12296), .A2(n15001), .ZN(n12297) );
  NAND2_X1 U14693 ( .A1(n12298), .A2(n12297), .ZN(n15019) );
  MUX2_X1 U14694 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n6717), .Z(n12299) );
  XNOR2_X1 U14695 ( .A(n12299), .B(n12339), .ZN(n15018) );
  INV_X1 U14696 ( .A(n12299), .ZN(n12300) );
  NAND2_X1 U14697 ( .A1(n12300), .A2(n15024), .ZN(n12301) );
  AND2_X1 U14698 ( .A1(n15033), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12319) );
  NOR2_X1 U14699 ( .A1(n15033), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n12302) );
  OR2_X1 U14700 ( .A1(n12319), .A2(n12302), .ZN(n15028) );
  AND2_X1 U14701 ( .A1(n15033), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12343) );
  NOR2_X1 U14702 ( .A1(n15033), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n12303) );
  OR2_X1 U14703 ( .A1(n12343), .A2(n12303), .ZN(n12330) );
  MUX2_X1 U14704 ( .A(n15028), .B(n12330), .S(n6717), .Z(n15044) );
  INV_X1 U14705 ( .A(n12319), .ZN(n12306) );
  INV_X1 U14706 ( .A(n12343), .ZN(n12305) );
  MUX2_X1 U14707 ( .A(n12306), .B(n12305), .S(n12304), .Z(n12307) );
  NAND2_X1 U14708 ( .A1(n15040), .A2(n12307), .ZN(n12308) );
  XNOR2_X1 U14709 ( .A(n12308), .B(n14413), .ZN(n14410) );
  MUX2_X1 U14710 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n6717), .Z(n14409) );
  XNOR2_X1 U14711 ( .A(n12309), .B(n14428), .ZN(n14432) );
  NAND2_X1 U14712 ( .A1(n14433), .A2(n14432), .ZN(n14435) );
  OAI21_X1 U14713 ( .B1(n12309), .B2(n12322), .A(n14435), .ZN(n14450) );
  XNOR2_X1 U14714 ( .A(n12310), .B(n12349), .ZN(n14451) );
  NOR2_X1 U14715 ( .A1(n14450), .A2(n14451), .ZN(n14449) );
  AOI21_X1 U14716 ( .B1(n12310), .B2(n12349), .A(n14449), .ZN(n12372) );
  XOR2_X1 U14717 ( .A(n14379), .B(n12372), .Z(n12311) );
  NOR2_X1 U14718 ( .A1(n12311), .A2(n12312), .ZN(n12370) );
  AOI21_X1 U14719 ( .B1(n12312), .B2(n12311), .A(n12370), .ZN(n12356) );
  INV_X1 U14720 ( .A(n14379), .ZN(n12371) );
  INV_X1 U14721 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n12530) );
  AND2_X1 U14722 ( .A1(n14379), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n12357) );
  AOI21_X1 U14723 ( .B1(n12371), .B2(n12530), .A(n12357), .ZN(n12327) );
  NOR2_X1 U14724 ( .A1(n12333), .A2(n12315), .ZN(n12316) );
  NOR2_X1 U14725 ( .A1(n14973), .A2(n14972), .ZN(n14971) );
  NAND2_X1 U14726 ( .A1(n15001), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n12317) );
  OAI21_X1 U14727 ( .B1(n15001), .B2(P3_REG2_REG_12__SCAN_IN), .A(n12317), 
        .ZN(n14989) );
  INV_X1 U14728 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n15010) );
  INV_X1 U14729 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n14406) );
  INV_X1 U14730 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n12321) );
  AOI22_X1 U14731 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n14428), .B1(n12322), 
        .B2(n12321), .ZN(n14423) );
  NOR2_X1 U14732 ( .A1(n14428), .A2(n12321), .ZN(n12323) );
  OAI21_X1 U14733 ( .B1(n6698), .B2(n12325), .A(n12324), .ZN(n12326) );
  NAND2_X1 U14734 ( .A1(n12326), .A2(n12327), .ZN(n12359) );
  OAI21_X1 U14735 ( .B1(n12327), .B2(n12326), .A(n12359), .ZN(n12329) );
  NAND2_X1 U14736 ( .A1(n12329), .A2(n12328), .ZN(n12355) );
  XNOR2_X1 U14737 ( .A(n14379), .B(P3_REG1_REG_18__SCAN_IN), .ZN(n12361) );
  XNOR2_X1 U14738 ( .A(n14428), .B(P3_REG1_REG_16__SCAN_IN), .ZN(n14426) );
  INV_X1 U14739 ( .A(n12330), .ZN(n15031) );
  NAND2_X1 U14740 ( .A1(n15001), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U14741 ( .A1(n14982), .A2(n12334), .ZN(n12335) );
  NAND2_X1 U14742 ( .A1(P3_REG1_REG_11__SCAN_IN), .A2(n14977), .ZN(n14976) );
  NAND2_X1 U14743 ( .A1(n12335), .A2(n14976), .ZN(n14994) );
  INV_X1 U14744 ( .A(n15001), .ZN(n12337) );
  INV_X1 U14745 ( .A(n12338), .ZN(n12336) );
  AOI21_X1 U14746 ( .B1(n12337), .B2(n8461), .A(n12336), .ZN(n14995) );
  NAND2_X1 U14747 ( .A1(n14994), .A2(n14995), .ZN(n14993) );
  NAND2_X1 U14748 ( .A1(n12338), .A2(n14993), .ZN(n12340) );
  NAND2_X1 U14749 ( .A1(n12339), .A2(n12340), .ZN(n12341) );
  NAND2_X1 U14750 ( .A1(n12341), .A2(n15011), .ZN(n15032) );
  NAND2_X1 U14751 ( .A1(n15031), .A2(n15032), .ZN(n15030) );
  INV_X1 U14752 ( .A(n15030), .ZN(n12342) );
  OR2_X1 U14753 ( .A1(n14413), .A2(n12345), .ZN(n12346) );
  XNOR2_X1 U14754 ( .A(n12345), .B(n12344), .ZN(n14408) );
  NAND2_X1 U14755 ( .A1(n14426), .A2(n14427), .ZN(n14425) );
  XOR2_X1 U14756 ( .A(n12361), .B(n12362), .Z(n12352) );
  AOI21_X1 U14757 ( .B1(n14998), .B2(P3_ADDR_REG_18__SCAN_IN), .A(n12350), 
        .ZN(n12351) );
  OAI21_X1 U14758 ( .B1(n12352), .B2(n12367), .A(n12351), .ZN(n12353) );
  AOI21_X1 U14759 ( .B1(n12371), .B2(n15035), .A(n12353), .ZN(n12354) );
  OAI211_X1 U14760 ( .C1(n12356), .C2(n15042), .A(n12355), .B(n12354), .ZN(
        P3_U3200) );
  INV_X1 U14761 ( .A(n12357), .ZN(n12358) );
  NAND2_X1 U14762 ( .A1(n12359), .A2(n12358), .ZN(n12360) );
  XNOR2_X1 U14763 ( .A(n12363), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n12369) );
  XNOR2_X1 U14764 ( .A(n12360), .B(n12369), .ZN(n12377) );
  XNOR2_X1 U14765 ( .A(n12363), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n12368) );
  XNOR2_X1 U14766 ( .A(n12364), .B(n12368), .ZN(n12366) );
  MUX2_X1 U14767 ( .A(n12369), .B(n12368), .S(n6717), .Z(n12373) );
  OAI21_X1 U14768 ( .B1(n12377), .B2(n15050), .A(n12376), .ZN(P3_U3201) );
  AOI22_X1 U14769 ( .A1(n14462), .A2(P3_REG2_REG_29__SCAN_IN), .B1(n14459), 
        .B2(n15098), .ZN(n12378) );
  OAI21_X1 U14770 ( .B1(n12379), .B2(n12587), .A(n12378), .ZN(n12380) );
  AOI21_X1 U14771 ( .B1(n12381), .B2(n12589), .A(n12380), .ZN(n12382) );
  OAI21_X1 U14772 ( .B1(n6525), .B2(n14462), .A(n12382), .ZN(P3_U3204) );
  NAND2_X1 U14773 ( .A1(n12399), .A2(n12383), .ZN(n12384) );
  XNOR2_X1 U14774 ( .A(n12384), .B(n12386), .ZN(n12619) );
  OAI211_X1 U14775 ( .C1(n12387), .C2(n12386), .A(n12385), .B(n15109), .ZN(
        n12391) );
  AOI22_X1 U14776 ( .A1(n12571), .A2(n12389), .B1(n12388), .B2(n12569), .ZN(
        n12390) );
  AND2_X1 U14777 ( .A1(n12391), .A2(n12390), .ZN(n12620) );
  INV_X1 U14778 ( .A(n12620), .ZN(n12395) );
  AOI22_X1 U14779 ( .A1(n14462), .A2(P3_REG2_REG_28__SCAN_IN), .B1(n15098), 
        .B2(n12392), .ZN(n12393) );
  OAI21_X1 U14780 ( .B1(n12686), .B2(n12587), .A(n12393), .ZN(n12394) );
  AOI21_X1 U14781 ( .B1(n12395), .B2(n15120), .A(n12394), .ZN(n12396) );
  OAI21_X1 U14782 ( .B1(n12619), .B2(n12618), .A(n12396), .ZN(P3_U3205) );
  NAND2_X1 U14783 ( .A1(n12399), .A2(n12398), .ZN(n12624) );
  INV_X1 U14784 ( .A(n12624), .ZN(n12415) );
  INV_X1 U14785 ( .A(n12400), .ZN(n12401) );
  AOI21_X1 U14786 ( .B1(n12403), .B2(n12402), .A(n12401), .ZN(n12408) );
  AOI22_X1 U14787 ( .A1(n12571), .A2(n12405), .B1(n12404), .B2(n12569), .ZN(
        n12407) );
  NAND2_X1 U14788 ( .A1(n12624), .A2(n15090), .ZN(n12406) );
  NAND2_X1 U14789 ( .A1(n12623), .A2(n15120), .ZN(n12414) );
  INV_X1 U14790 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n12410) );
  OAI22_X1 U14791 ( .A1(n15120), .A2(n12410), .B1(n12409), .B2(n15114), .ZN(
        n12411) );
  AOI21_X1 U14792 ( .B1(n12412), .B2(n15081), .A(n12411), .ZN(n12413) );
  OAI211_X1 U14793 ( .C1(n12415), .C2(n15116), .A(n12414), .B(n12413), .ZN(
        P3_U3206) );
  XOR2_X1 U14794 ( .A(n12416), .B(n12417), .Z(n12628) );
  INV_X1 U14795 ( .A(n12628), .ZN(n12427) );
  XNOR2_X1 U14796 ( .A(n12418), .B(n12417), .ZN(n12419) );
  OAI222_X1 U14797 ( .A1(n15106), .A2(n12421), .B1(n15104), .B2(n12420), .C1(
        n12419), .C2(n15093), .ZN(n12627) );
  INV_X1 U14798 ( .A(n12422), .ZN(n12694) );
  AOI22_X1 U14799 ( .A1(n14462), .A2(P3_REG2_REG_26__SCAN_IN), .B1(n15098), 
        .B2(n12423), .ZN(n12424) );
  OAI21_X1 U14800 ( .B1(n12694), .B2(n12587), .A(n12424), .ZN(n12425) );
  AOI21_X1 U14801 ( .B1(n12627), .B2(n15120), .A(n12425), .ZN(n12426) );
  OAI21_X1 U14802 ( .B1(n12618), .B2(n12427), .A(n12426), .ZN(P3_U3207) );
  XOR2_X1 U14803 ( .A(n12428), .B(n12431), .Z(n12634) );
  INV_X1 U14804 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n12430) );
  OAI22_X1 U14805 ( .A1(n15120), .A2(n12430), .B1(n12429), .B2(n15114), .ZN(
        n12438) );
  AOI21_X1 U14806 ( .B1(n12432), .B2(n12431), .A(n15093), .ZN(n12436) );
  OAI22_X1 U14807 ( .A1(n12456), .A2(n15106), .B1(n12433), .B2(n15104), .ZN(
        n12434) );
  AOI21_X1 U14808 ( .B1(n12436), .B2(n12435), .A(n12434), .ZN(n12633) );
  NOR2_X1 U14809 ( .A1(n12633), .A2(n14462), .ZN(n12437) );
  AOI211_X1 U14810 ( .C1(n15081), .C2(n12631), .A(n12438), .B(n12437), .ZN(
        n12439) );
  OAI21_X1 U14811 ( .B1(n12618), .B2(n12634), .A(n12439), .ZN(P3_U3208) );
  XNOR2_X1 U14812 ( .A(n12440), .B(n12447), .ZN(n12443) );
  AOI222_X1 U14813 ( .A1(n15109), .A2(n12443), .B1(n12442), .B2(n12571), .C1(
        n12441), .C2(n12569), .ZN(n12637) );
  AND2_X1 U14814 ( .A1(n12444), .A2(n12445), .ZN(n12448) );
  OAI21_X1 U14815 ( .B1(n12448), .B2(n12447), .A(n12446), .ZN(n12635) );
  INV_X1 U14816 ( .A(n12449), .ZN(n12450) );
  AOI22_X1 U14817 ( .A1(n14462), .A2(P3_REG2_REG_24__SCAN_IN), .B1(n15098), 
        .B2(n12450), .ZN(n12451) );
  OAI21_X1 U14818 ( .B1(n12638), .B2(n12587), .A(n12451), .ZN(n12452) );
  AOI21_X1 U14819 ( .B1(n12635), .B2(n12589), .A(n12452), .ZN(n12453) );
  OAI21_X1 U14820 ( .B1(n12637), .B2(n14462), .A(n12453), .ZN(P3_U3209) );
  XNOR2_X1 U14821 ( .A(n12454), .B(n12459), .ZN(n12455) );
  OAI222_X1 U14822 ( .A1(n15104), .A2(n12456), .B1(n15106), .B2(n12482), .C1(
        n12455), .C2(n15093), .ZN(n12639) );
  INV_X1 U14823 ( .A(n12639), .ZN(n12465) );
  INV_X1 U14824 ( .A(n12457), .ZN(n12460) );
  INV_X1 U14825 ( .A(n12444), .ZN(n12458) );
  AOI21_X1 U14826 ( .B1(n12460), .B2(n12459), .A(n12458), .ZN(n12640) );
  AOI22_X1 U14827 ( .A1(n14462), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n15098), 
        .B2(n12461), .ZN(n12462) );
  OAI21_X1 U14828 ( .B1(n12700), .B2(n12587), .A(n12462), .ZN(n12463) );
  AOI21_X1 U14829 ( .B1(n12640), .B2(n12589), .A(n12463), .ZN(n12464) );
  OAI21_X1 U14830 ( .B1(n14462), .B2(n12465), .A(n12464), .ZN(P3_U3210) );
  XNOR2_X1 U14831 ( .A(n12466), .B(n12467), .ZN(n12644) );
  INV_X1 U14832 ( .A(n12644), .ZN(n12477) );
  XNOR2_X1 U14833 ( .A(n12468), .B(n12467), .ZN(n12469) );
  OAI222_X1 U14834 ( .A1(n15104), .A2(n12471), .B1(n15106), .B2(n12470), .C1(
        n12469), .C2(n15093), .ZN(n12643) );
  INV_X1 U14835 ( .A(n12472), .ZN(n12704) );
  AOI22_X1 U14836 ( .A1(n14462), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n15098), 
        .B2(n12473), .ZN(n12474) );
  OAI21_X1 U14837 ( .B1(n12704), .B2(n12587), .A(n12474), .ZN(n12475) );
  AOI21_X1 U14838 ( .B1(n12643), .B2(n15120), .A(n12475), .ZN(n12476) );
  OAI21_X1 U14839 ( .B1(n12618), .B2(n12477), .A(n12476), .ZN(P3_U3211) );
  XNOR2_X1 U14840 ( .A(n12478), .B(n12479), .ZN(n12648) );
  INV_X1 U14841 ( .A(n12648), .ZN(n12487) );
  XNOR2_X1 U14842 ( .A(n12480), .B(n12479), .ZN(n12481) );
  OAI222_X1 U14843 ( .A1(n15104), .A2(n12482), .B1(n15106), .B2(n12510), .C1(
        n15093), .C2(n12481), .ZN(n12647) );
  AOI22_X1 U14844 ( .A1(n14462), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n15098), 
        .B2(n12483), .ZN(n12484) );
  OAI21_X1 U14845 ( .B1(n12708), .B2(n12587), .A(n12484), .ZN(n12485) );
  AOI21_X1 U14846 ( .B1(n12647), .B2(n15120), .A(n12485), .ZN(n12486) );
  OAI21_X1 U14847 ( .B1(n12618), .B2(n12487), .A(n12486), .ZN(P3_U3212) );
  NAND2_X1 U14848 ( .A1(n12488), .A2(n12494), .ZN(n12489) );
  NAND2_X1 U14849 ( .A1(n12490), .A2(n12489), .ZN(n12652) );
  NAND2_X1 U14850 ( .A1(n12523), .A2(n12492), .ZN(n12509) );
  INV_X1 U14851 ( .A(n12519), .ZN(n12508) );
  NAND2_X1 U14852 ( .A1(n12513), .A2(n12493), .ZN(n12496) );
  INV_X1 U14853 ( .A(n12494), .ZN(n12495) );
  XNOR2_X1 U14854 ( .A(n12496), .B(n12495), .ZN(n12497) );
  NAND2_X1 U14855 ( .A1(n12497), .A2(n15109), .ZN(n12501) );
  AOI22_X1 U14856 ( .A1(n12499), .A2(n12571), .B1(n12569), .B2(n12498), .ZN(
        n12500) );
  NAND2_X1 U14857 ( .A1(n12501), .A2(n12500), .ZN(n12654) );
  NAND2_X1 U14858 ( .A1(n12654), .A2(n15120), .ZN(n12507) );
  INV_X1 U14859 ( .A(P3_REG2_REG_20__SCAN_IN), .ZN(n12503) );
  OAI22_X1 U14860 ( .A1(n15120), .A2(n12503), .B1(n12502), .B2(n15114), .ZN(
        n12504) );
  AOI21_X1 U14861 ( .B1(n12505), .B2(n15081), .A(n12504), .ZN(n12506) );
  OAI211_X1 U14862 ( .C1(n12618), .C2(n12652), .A(n12507), .B(n12506), .ZN(
        P3_U3213) );
  AOI21_X1 U14863 ( .B1(n12509), .B2(n12508), .A(n15093), .ZN(n12514) );
  OAI22_X1 U14864 ( .A1(n12511), .A2(n15106), .B1(n12510), .B2(n15104), .ZN(
        n12512) );
  AOI21_X1 U14865 ( .B1(n12514), .B2(n12513), .A(n12512), .ZN(n12657) );
  INV_X1 U14866 ( .A(n12713), .ZN(n12518) );
  INV_X1 U14867 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n12516) );
  OAI22_X1 U14868 ( .A1(n15120), .A2(n12516), .B1(n12515), .B2(n15114), .ZN(
        n12517) );
  AOI21_X1 U14869 ( .B1(n12518), .B2(n15081), .A(n12517), .ZN(n12522) );
  XNOR2_X1 U14870 ( .A(n12520), .B(n12519), .ZN(n12655) );
  NAND2_X1 U14871 ( .A1(n12655), .A2(n12589), .ZN(n12521) );
  OAI211_X1 U14872 ( .C1(n12657), .C2(n14462), .A(n12522), .B(n12521), .ZN(
        P3_U3214) );
  INV_X1 U14873 ( .A(n12523), .ZN(n12524) );
  AOI21_X1 U14874 ( .B1(n12525), .B2(n12491), .A(n12524), .ZN(n12526) );
  OAI222_X1 U14875 ( .A1(n15104), .A2(n12528), .B1(n15106), .B2(n12527), .C1(
        n15093), .C2(n12526), .ZN(n12661) );
  INV_X1 U14876 ( .A(n12661), .ZN(n12541) );
  OAI22_X1 U14877 ( .A1(n15120), .A2(n12530), .B1(n12529), .B2(n15114), .ZN(
        n12538) );
  NAND2_X1 U14878 ( .A1(n12545), .A2(n6970), .ZN(n12533) );
  NAND2_X1 U14879 ( .A1(n12533), .A2(n12531), .ZN(n12662) );
  INV_X1 U14880 ( .A(n12662), .ZN(n12536) );
  NAND2_X1 U14881 ( .A1(n12533), .A2(n12532), .ZN(n12535) );
  NOR3_X1 U14882 ( .A1(n12536), .A2(n12660), .A3(n12618), .ZN(n12537) );
  AOI211_X1 U14883 ( .C1(n15081), .C2(n12539), .A(n12538), .B(n12537), .ZN(
        n12540) );
  OAI21_X1 U14884 ( .B1(n12541), .B2(n14462), .A(n12540), .ZN(P3_U3215) );
  XNOR2_X1 U14885 ( .A(n12542), .B(n6970), .ZN(n12544) );
  AOI222_X1 U14886 ( .A1(n15109), .A2(n12544), .B1(n12543), .B2(n12571), .C1(
        n12572), .C2(n12569), .ZN(n12669) );
  XNOR2_X1 U14887 ( .A(n12545), .B(n6970), .ZN(n12667) );
  NOR2_X1 U14888 ( .A1(n12546), .A2(n12587), .ZN(n12549) );
  OAI22_X1 U14889 ( .A1(n15120), .A2(n14443), .B1(n12547), .B2(n15114), .ZN(
        n12548) );
  AOI211_X1 U14890 ( .C1(n12667), .C2(n12589), .A(n12549), .B(n12548), .ZN(
        n12550) );
  OAI21_X1 U14891 ( .B1(n12669), .B2(n14462), .A(n12550), .ZN(P3_U3216) );
  NAND2_X1 U14892 ( .A1(n12551), .A2(n12583), .ZN(n12567) );
  NAND2_X1 U14893 ( .A1(n12567), .A2(n12552), .ZN(n12554) );
  AND2_X1 U14894 ( .A1(n12554), .A2(n12553), .ZN(n12555) );
  XNOR2_X1 U14895 ( .A(n12555), .B(n12559), .ZN(n12558) );
  AOI222_X1 U14896 ( .A1(n15109), .A2(n12558), .B1(n12557), .B2(n12571), .C1(
        n12556), .C2(n12569), .ZN(n12673) );
  XNOR2_X1 U14897 ( .A(n12560), .B(n12559), .ZN(n12671) );
  AOI22_X1 U14898 ( .A1(n14462), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n15098), 
        .B2(n12561), .ZN(n12562) );
  OAI21_X1 U14899 ( .B1(n12563), .B2(n12587), .A(n12562), .ZN(n12564) );
  AOI21_X1 U14900 ( .B1(n12671), .B2(n12589), .A(n12564), .ZN(n12565) );
  OAI21_X1 U14901 ( .B1(n12673), .B2(n14462), .A(n12565), .ZN(P3_U3217) );
  NAND2_X1 U14902 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  XNOR2_X1 U14903 ( .A(n12568), .B(n12576), .ZN(n12573) );
  AOI222_X1 U14904 ( .A1(n15109), .A2(n12573), .B1(n12572), .B2(n12571), .C1(
        n12570), .C2(n12569), .ZN(n12677) );
  OAI22_X1 U14905 ( .A1(n15120), .A2(n14406), .B1(n12574), .B2(n15114), .ZN(
        n12575) );
  AOI21_X1 U14906 ( .B1(n12674), .B2(n15081), .A(n12575), .ZN(n12579) );
  XNOR2_X1 U14907 ( .A(n12577), .B(n12576), .ZN(n12675) );
  NAND2_X1 U14908 ( .A1(n12675), .A2(n12589), .ZN(n12578) );
  OAI211_X1 U14909 ( .C1(n12677), .C2(n14462), .A(n12579), .B(n12578), .ZN(
        P3_U3218) );
  XNOR2_X1 U14910 ( .A(n12551), .B(n12583), .ZN(n12580) );
  OAI222_X1 U14911 ( .A1(n15104), .A2(n12582), .B1(n15106), .B2(n12581), .C1(
        n12580), .C2(n15093), .ZN(n12678) );
  INV_X1 U14912 ( .A(n12678), .ZN(n12591) );
  XNOR2_X1 U14913 ( .A(n12584), .B(n12583), .ZN(n12679) );
  AOI22_X1 U14914 ( .A1(n14462), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n15098), 
        .B2(n12585), .ZN(n12586) );
  OAI21_X1 U14915 ( .B1(n12725), .B2(n12587), .A(n12586), .ZN(n12588) );
  AOI21_X1 U14916 ( .B1(n12679), .B2(n12589), .A(n12588), .ZN(n12590) );
  OAI21_X1 U14917 ( .B1(n12591), .B2(n14462), .A(n12590), .ZN(P3_U3219) );
  XOR2_X1 U14918 ( .A(n12594), .B(n12592), .Z(n14472) );
  XOR2_X1 U14919 ( .A(n12594), .B(n12593), .Z(n12595) );
  OAI222_X1 U14920 ( .A1(n15104), .A2(n12597), .B1(n15106), .B2(n12596), .C1(
        n12595), .C2(n15093), .ZN(n14473) );
  NAND2_X1 U14921 ( .A1(n14473), .A2(n15120), .ZN(n12601) );
  OAI22_X1 U14922 ( .A1(n15120), .A2(n15010), .B1(n12598), .B2(n15114), .ZN(
        n12599) );
  AOI21_X1 U14923 ( .B1(n14475), .B2(n15081), .A(n12599), .ZN(n12600) );
  OAI211_X1 U14924 ( .C1(n12618), .C2(n14472), .A(n12601), .B(n12600), .ZN(
        P3_U3220) );
  XNOR2_X1 U14925 ( .A(n12602), .B(n12607), .ZN(n15140) );
  NAND2_X1 U14926 ( .A1(n12604), .A2(n12603), .ZN(n12606) );
  NAND2_X1 U14927 ( .A1(n12606), .A2(n12605), .ZN(n12608) );
  XNOR2_X1 U14928 ( .A(n12608), .B(n12607), .ZN(n12609) );
  OAI222_X1 U14929 ( .A1(n15104), .A2(n12611), .B1(n15106), .B2(n12610), .C1(
        n12609), .C2(n15093), .ZN(n15142) );
  NAND2_X1 U14930 ( .A1(n15142), .A2(n15120), .ZN(n12617) );
  OAI22_X1 U14931 ( .A1(n15120), .A2(n12613), .B1(n12612), .B2(n15114), .ZN(
        n12614) );
  AOI21_X1 U14932 ( .B1(n15081), .B2(n12615), .A(n12614), .ZN(n12616) );
  OAI211_X1 U14933 ( .C1(n12618), .C2(n15140), .A(n12617), .B(n12616), .ZN(
        P3_U3223) );
  MUX2_X1 U14934 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n12683), .S(n15149), .Z(
        n12621) );
  INV_X1 U14935 ( .A(n12621), .ZN(n12622) );
  OAI21_X1 U14936 ( .B1(n12686), .B2(n12682), .A(n12622), .ZN(P3_U3487) );
  MUX2_X1 U14937 ( .A(n12625), .B(n12687), .S(n15149), .Z(n12626) );
  OAI21_X1 U14938 ( .B1(n12690), .B2(n12682), .A(n12626), .ZN(P3_U3486) );
  AOI21_X1 U14939 ( .B1(n12628), .B2(n14482), .A(n12627), .ZN(n12691) );
  MUX2_X1 U14940 ( .A(n12629), .B(n12691), .S(n15149), .Z(n12630) );
  OAI21_X1 U14941 ( .B1(n12694), .B2(n12682), .A(n12630), .ZN(P3_U3485) );
  NAND2_X1 U14942 ( .A1(n12631), .A2(n14476), .ZN(n12632) );
  OAI211_X1 U14943 ( .C1(n12634), .C2(n15139), .A(n12633), .B(n12632), .ZN(
        n12695) );
  MUX2_X1 U14944 ( .A(P3_REG1_REG_25__SCAN_IN), .B(n12695), .S(n15149), .Z(
        P3_U3484) );
  NAND2_X1 U14945 ( .A1(n12635), .A2(n14482), .ZN(n12636) );
  OAI211_X1 U14946 ( .C1(n12638), .C2(n15138), .A(n12637), .B(n12636), .ZN(
        n12696) );
  MUX2_X1 U14947 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12696), .S(n15149), .Z(
        P3_U3483) );
  AOI21_X1 U14948 ( .B1(n12640), .B2(n14482), .A(n12639), .ZN(n12697) );
  MUX2_X1 U14949 ( .A(n12641), .B(n12697), .S(n15149), .Z(n12642) );
  OAI21_X1 U14950 ( .B1(n12700), .B2(n12682), .A(n12642), .ZN(P3_U3482) );
  AOI21_X1 U14951 ( .B1(n14482), .B2(n12644), .A(n12643), .ZN(n12701) );
  MUX2_X1 U14952 ( .A(n12645), .B(n12701), .S(n15149), .Z(n12646) );
  OAI21_X1 U14953 ( .B1(n12704), .B2(n12682), .A(n12646), .ZN(P3_U3481) );
  AOI21_X1 U14954 ( .B1(n12648), .B2(n14482), .A(n12647), .ZN(n12705) );
  MUX2_X1 U14955 ( .A(n12649), .B(n12705), .S(n15149), .Z(n12650) );
  OAI21_X1 U14956 ( .B1(n12708), .B2(n12682), .A(n12650), .ZN(P3_U3480) );
  OAI22_X1 U14957 ( .A1(n12652), .A2(n15139), .B1(n12651), .B2(n15138), .ZN(
        n12653) );
  MUX2_X1 U14958 ( .A(P3_REG1_REG_20__SCAN_IN), .B(n12709), .S(n15149), .Z(
        P3_U3479) );
  NAND2_X1 U14959 ( .A1(n12655), .A2(n14482), .ZN(n12656) );
  AND2_X1 U14960 ( .A1(n12657), .A2(n12656), .ZN(n12710) );
  MUX2_X1 U14961 ( .A(n12658), .B(n12710), .S(n15149), .Z(n12659) );
  OAI21_X1 U14962 ( .B1(n12682), .B2(n12713), .A(n12659), .ZN(P3_U3478) );
  NOR2_X1 U14963 ( .A1(n12660), .A2(n15139), .ZN(n12663) );
  AOI21_X1 U14964 ( .B1(n12663), .B2(n12662), .A(n12661), .ZN(n12714) );
  MUX2_X1 U14965 ( .A(n12664), .B(n12714), .S(n15149), .Z(n12665) );
  OAI21_X1 U14966 ( .B1(n12717), .B2(n12682), .A(n12665), .ZN(P3_U3477) );
  AOI22_X1 U14967 ( .A1(n12667), .A2(n14482), .B1(n14476), .B2(n12666), .ZN(
        n12668) );
  NAND2_X1 U14968 ( .A1(n12669), .A2(n12668), .ZN(n12718) );
  MUX2_X1 U14969 ( .A(P3_REG1_REG_17__SCAN_IN), .B(n12718), .S(n15149), .Z(
        P3_U3476) );
  AOI22_X1 U14970 ( .A1(n12671), .A2(n14482), .B1(n14476), .B2(n12670), .ZN(
        n12672) );
  NAND2_X1 U14971 ( .A1(n12673), .A2(n12672), .ZN(n12719) );
  MUX2_X1 U14972 ( .A(P3_REG1_REG_16__SCAN_IN), .B(n12719), .S(n15149), .Z(
        P3_U3475) );
  AOI22_X1 U14973 ( .A1(n12675), .A2(n14482), .B1(n14476), .B2(n12674), .ZN(
        n12676) );
  NAND2_X1 U14974 ( .A1(n12677), .A2(n12676), .ZN(n12720) );
  MUX2_X1 U14975 ( .A(P3_REG1_REG_15__SCAN_IN), .B(n12720), .S(n15149), .Z(
        P3_U3474) );
  AOI21_X1 U14976 ( .B1(n14482), .B2(n12679), .A(n12678), .ZN(n12721) );
  MUX2_X1 U14977 ( .A(n12680), .B(n12721), .S(n15149), .Z(n12681) );
  OAI21_X1 U14978 ( .B1(n12725), .B2(n12682), .A(n12681), .ZN(P3_U3473) );
  INV_X1 U14979 ( .A(n12683), .ZN(n12685) );
  MUX2_X1 U14980 ( .A(n12688), .B(n12687), .S(n15143), .Z(n12689) );
  OAI21_X1 U14981 ( .B1(n12690), .B2(n12724), .A(n12689), .ZN(P3_U3454) );
  MUX2_X1 U14982 ( .A(n12692), .B(n12691), .S(n15143), .Z(n12693) );
  OAI21_X1 U14983 ( .B1(n12694), .B2(n12724), .A(n12693), .ZN(P3_U3453) );
  MUX2_X1 U14984 ( .A(P3_REG0_REG_25__SCAN_IN), .B(n12695), .S(n15143), .Z(
        P3_U3452) );
  MUX2_X1 U14985 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12696), .S(n15143), .Z(
        P3_U3451) );
  MUX2_X1 U14986 ( .A(n12698), .B(n12697), .S(n15143), .Z(n12699) );
  OAI21_X1 U14987 ( .B1(n12700), .B2(n12724), .A(n12699), .ZN(P3_U3450) );
  MUX2_X1 U14988 ( .A(n12702), .B(n12701), .S(n15143), .Z(n12703) );
  OAI21_X1 U14989 ( .B1(n12704), .B2(n12724), .A(n12703), .ZN(P3_U3449) );
  MUX2_X1 U14990 ( .A(n12706), .B(n12705), .S(n15143), .Z(n12707) );
  OAI21_X1 U14991 ( .B1(n12708), .B2(n12724), .A(n12707), .ZN(P3_U3448) );
  MUX2_X1 U14992 ( .A(n12709), .B(P3_REG0_REG_20__SCAN_IN), .S(n15144), .Z(
        P3_U3447) );
  MUX2_X1 U14993 ( .A(n12711), .B(n12710), .S(n15143), .Z(n12712) );
  OAI21_X1 U14994 ( .B1(n12724), .B2(n12713), .A(n12712), .ZN(P3_U3446) );
  MUX2_X1 U14995 ( .A(n12715), .B(n12714), .S(n15143), .Z(n12716) );
  OAI21_X1 U14996 ( .B1(n12717), .B2(n12724), .A(n12716), .ZN(P3_U3444) );
  MUX2_X1 U14997 ( .A(P3_REG0_REG_17__SCAN_IN), .B(n12718), .S(n15143), .Z(
        P3_U3441) );
  MUX2_X1 U14998 ( .A(P3_REG0_REG_16__SCAN_IN), .B(n12719), .S(n15143), .Z(
        P3_U3438) );
  MUX2_X1 U14999 ( .A(P3_REG0_REG_15__SCAN_IN), .B(n12720), .S(n15143), .Z(
        P3_U3435) );
  MUX2_X1 U15000 ( .A(n12722), .B(n12721), .S(n15143), .Z(n12723) );
  OAI21_X1 U15001 ( .B1(n12725), .B2(n12724), .A(n12723), .ZN(P3_U3432) );
  NAND3_X1 U15002 ( .A1(n6624), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n12728) );
  OAI22_X1 U15003 ( .A1(n12729), .A2(n12728), .B1(n12727), .B2(n12726), .ZN(
        n12730) );
  AOI21_X1 U15004 ( .B1(n12731), .B2(n14376), .A(n12730), .ZN(n12732) );
  INV_X1 U15005 ( .A(n12732), .ZN(P3_U3264) );
  INV_X1 U15006 ( .A(n12733), .ZN(n12735) );
  OAI222_X1 U15007 ( .A1(P3_U3151), .A2(n12736), .B1(n12747), .B2(n12735), 
        .C1(n12734), .C2(n12744), .ZN(P3_U3266) );
  INV_X1 U15008 ( .A(n12737), .ZN(n12738) );
  INV_X1 U15009 ( .A(n12740), .ZN(n12742) );
  OAI222_X1 U15010 ( .A1(P3_U3151), .A2(n6717), .B1(n12747), .B2(n12742), .C1(
        n12741), .C2(n12744), .ZN(P3_U3268) );
  INV_X1 U15011 ( .A(n12743), .ZN(n12746) );
  OAI222_X1 U15012 ( .A1(n12749), .A2(P3_U3151), .B1(n12747), .B2(n12746), 
        .C1(n12745), .C2(n12744), .ZN(P3_U3269) );
  NAND2_X1 U15013 ( .A1(n12751), .A2(n12750), .ZN(n12752) );
  NAND3_X1 U15014 ( .A1(n12753), .A2(n14494), .A3(n12752), .ZN(n12758) );
  OAI22_X1 U15015 ( .A1(n12943), .A2(n12913), .B1(n12983), .B2(n12843), .ZN(
        n13008) );
  INV_X1 U15016 ( .A(n13012), .ZN(n12755) );
  OAI22_X1 U15017 ( .A1(n12755), .A2(n14502), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12754), .ZN(n12756) );
  AOI21_X1 U15018 ( .B1(n13008), .B2(n14496), .A(n12756), .ZN(n12757) );
  OAI211_X1 U15019 ( .C1(n6953), .C2(n12846), .A(n12758), .B(n12757), .ZN(
        P2_U3186) );
  AOI22_X1 U15020 ( .A1(n12759), .A2(n14494), .B1(n12822), .B2(n12854), .ZN(
        n12768) );
  INV_X1 U15021 ( .A(n12760), .ZN(n12767) );
  OR2_X1 U15022 ( .A1(n12977), .A2(n12913), .ZN(n12762) );
  NAND2_X1 U15023 ( .A1(n12972), .A2(n12947), .ZN(n12761) );
  AND2_X1 U15024 ( .A1(n12762), .A2(n12761), .ZN(n13070) );
  INV_X1 U15025 ( .A(n13078), .ZN(n12763) );
  AOI22_X1 U15026 ( .A1(n12763), .A2(n12842), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12764) );
  OAI21_X1 U15027 ( .B1(n13070), .B2(n12783), .A(n12764), .ZN(n12765) );
  AOI21_X1 U15028 ( .B1(n13081), .B2(n14499), .A(n12765), .ZN(n12766) );
  OAI21_X1 U15029 ( .B1(n12768), .B2(n12767), .A(n12766), .ZN(P2_U3188) );
  INV_X1 U15030 ( .A(n12769), .ZN(n12772) );
  NOR3_X1 U15031 ( .A1(n12770), .A2(n12961), .A3(n12837), .ZN(n12771) );
  AOI21_X1 U15032 ( .B1(n12772), .B2(n14494), .A(n12771), .ZN(n12780) );
  INV_X1 U15033 ( .A(n12773), .ZN(n12812) );
  INV_X1 U15034 ( .A(n12967), .ZN(n12855) );
  NOR2_X1 U15035 ( .A1(n12961), .A2(n12843), .ZN(n12774) );
  AOI21_X1 U15036 ( .B1(n12855), .B2(n12781), .A(n12774), .ZN(n13133) );
  NAND2_X1 U15037 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n12906)
         );
  OAI21_X1 U15038 ( .B1(n13133), .B2(n12783), .A(n12906), .ZN(n12775) );
  AOI21_X1 U15039 ( .B1(n13140), .B2(n12842), .A(n12775), .ZN(n12776) );
  OAI21_X1 U15040 ( .B1(n13244), .B2(n12846), .A(n12776), .ZN(n12777) );
  AOI21_X1 U15041 ( .B1(n12812), .B2(n14494), .A(n12777), .ZN(n12778) );
  OAI21_X1 U15042 ( .B1(n12780), .B2(n12779), .A(n12778), .ZN(P2_U3191) );
  AOI22_X1 U15043 ( .A1(n12972), .A2(n12781), .B1(n12947), .B2(n12855), .ZN(
        n13112) );
  AOI22_X1 U15044 ( .A1(n12842), .A2(n13102), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12782) );
  OAI21_X1 U15045 ( .B1(n13112), .B2(n12783), .A(n12782), .ZN(n12789) );
  INV_X1 U15046 ( .A(n12784), .ZN(n12785) );
  AOI211_X1 U15047 ( .C1(n12787), .C2(n12786), .A(n12816), .B(n12785), .ZN(
        n12788) );
  AOI211_X1 U15048 ( .C1(n13230), .C2(n14499), .A(n12789), .B(n12788), .ZN(
        n12790) );
  INV_X1 U15049 ( .A(n12790), .ZN(P2_U3195) );
  INV_X1 U15050 ( .A(n12791), .ZN(n12792) );
  AOI21_X1 U15051 ( .B1(n12801), .B2(n12792), .A(n12816), .ZN(n12796) );
  NOR3_X1 U15052 ( .A1(n12793), .A2(n12977), .A3(n12837), .ZN(n12795) );
  OAI21_X1 U15053 ( .B1(n12796), .B2(n12795), .A(n12794), .ZN(n12800) );
  OAI22_X1 U15054 ( .A1(n12983), .A2(n12913), .B1(n12977), .B2(n12843), .ZN(
        n13035) );
  OAI22_X1 U15055 ( .A1(n13043), .A2(n14502), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12797), .ZN(n12798) );
  AOI21_X1 U15056 ( .B1(n13035), .B2(n14496), .A(n12798), .ZN(n12799) );
  OAI211_X1 U15057 ( .C1(n13039), .C2(n12846), .A(n12800), .B(n12799), .ZN(
        P2_U3197) );
  OAI211_X1 U15058 ( .C1(n12803), .C2(n12802), .A(n12801), .B(n14494), .ZN(
        n12807) );
  OAI22_X1 U15059 ( .A1(n12980), .A2(n12913), .B1(n12974), .B2(n12843), .ZN(
        n13050) );
  OAI22_X1 U15060 ( .A1(n13058), .A2(n14502), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12804), .ZN(n12805) );
  AOI21_X1 U15061 ( .B1(n13050), .B2(n14496), .A(n12805), .ZN(n12806) );
  OAI211_X1 U15062 ( .C1(n13054), .C2(n12846), .A(n12807), .B(n12806), .ZN(
        P2_U3201) );
  OAI22_X1 U15063 ( .A1(n12935), .A2(n12913), .B1(n12964), .B2(n12843), .ZN(
        n13126) );
  AOI22_X1 U15064 ( .A1(n13126), .A2(n14496), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12808) );
  OAI21_X1 U15065 ( .B1(n13119), .B2(n14502), .A(n12808), .ZN(n12814) );
  AOI22_X1 U15066 ( .A1(n12809), .A2(n14494), .B1(n12822), .B2(n12930), .ZN(
        n12811) );
  NOR3_X1 U15067 ( .A1(n12812), .A2(n12811), .A3(n12810), .ZN(n12813) );
  AOI211_X1 U15068 ( .C1(n13237), .C2(n14499), .A(n12814), .B(n12813), .ZN(
        n12815) );
  OAI21_X1 U15069 ( .B1(n12817), .B2(n12816), .A(n12815), .ZN(P2_U3205) );
  XNOR2_X1 U15070 ( .A(n12819), .B(n12818), .ZN(n12821) );
  NAND3_X1 U15071 ( .A1(n12821), .A2(n14494), .A3(n12820), .ZN(n12831) );
  INV_X1 U15072 ( .A(n12821), .ZN(n12823) );
  NAND3_X1 U15073 ( .A1(n12823), .A2(n12822), .A3(n12972), .ZN(n12830) );
  OAI22_X1 U15074 ( .A1(n12974), .A2(n12913), .B1(n12935), .B2(n12843), .ZN(
        n13087) );
  INV_X1 U15075 ( .A(n13095), .ZN(n12825) );
  OAI22_X1 U15076 ( .A1(n12825), .A2(n14502), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12824), .ZN(n12828) );
  NOR2_X1 U15077 ( .A1(n12826), .A2(n12846), .ZN(n12827) );
  AOI211_X1 U15078 ( .C1(n14496), .C2(n13087), .A(n12828), .B(n12827), .ZN(
        n12829) );
  NAND3_X1 U15079 ( .A1(n12831), .A2(n12830), .A3(n12829), .ZN(P2_U3207) );
  OAI211_X1 U15080 ( .C1(n12833), .C2(n12832), .A(n12769), .B(n14494), .ZN(
        n12836) );
  OAI22_X1 U15081 ( .A1(n12964), .A2(n12913), .B1(n12958), .B2(n12843), .ZN(
        n13148) );
  AND2_X1 U15082 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n12880) );
  NOR2_X1 U15083 ( .A1(n14502), .A2(n13152), .ZN(n12834) );
  AOI211_X1 U15084 ( .C1(n14496), .C2(n13148), .A(n12880), .B(n12834), .ZN(
        n12835) );
  OAI211_X1 U15085 ( .C1(n13155), .C2(n12846), .A(n12836), .B(n12835), .ZN(
        P2_U3210) );
  INV_X1 U15086 ( .A(n12794), .ZN(n12840) );
  NOR3_X1 U15087 ( .A1(n12838), .A2(n12980), .A3(n12837), .ZN(n12839) );
  AOI21_X1 U15088 ( .B1(n12840), .B2(n14494), .A(n12839), .ZN(n12851) );
  INV_X1 U15089 ( .A(n12841), .ZN(n12848) );
  AOI22_X1 U15090 ( .A1(n13026), .A2(n12842), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12845) );
  OAI22_X1 U15091 ( .A1(n12942), .A2(n12913), .B1(n12980), .B2(n12843), .ZN(
        n13021) );
  NAND2_X1 U15092 ( .A1(n13021), .A2(n14496), .ZN(n12844) );
  OAI211_X1 U15093 ( .C1(n13028), .C2(n12846), .A(n12845), .B(n12844), .ZN(
        n12847) );
  AOI21_X1 U15094 ( .B1(n12848), .B2(n14494), .A(n12847), .ZN(n12849) );
  OAI21_X1 U15095 ( .B1(n12851), .B2(n12850), .A(n12849), .ZN(P2_U3212) );
  MUX2_X1 U15096 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n12948), .S(n12871), .Z(
        P2_U3561) );
  MUX2_X1 U15097 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n12852), .S(n12871), .Z(
        P2_U3560) );
  MUX2_X1 U15098 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n12946), .S(P2_U3947), .Z(
        P2_U3559) );
  MUX2_X1 U15099 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n12985), .S(P2_U3947), .Z(
        P2_U3558) );
  MUX2_X1 U15100 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n12941), .S(P2_U3947), .Z(
        P2_U3557) );
  MUX2_X1 U15101 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n12853), .S(P2_U3947), .Z(
        P2_U3556) );
  INV_X1 U15102 ( .A(n12977), .ZN(n12940) );
  MUX2_X1 U15103 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n12940), .S(P2_U3947), .Z(
        P2_U3555) );
  MUX2_X1 U15104 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n12854), .S(n12871), .Z(
        P2_U3554) );
  MUX2_X1 U15105 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n12972), .S(n12871), .Z(
        P2_U3553) );
  MUX2_X1 U15106 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n12969), .S(n12871), .Z(
        P2_U3552) );
  MUX2_X1 U15107 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n12855), .S(n12871), .Z(
        P2_U3551) );
  MUX2_X1 U15108 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n12930), .S(n12871), .Z(
        P2_U3550) );
  MUX2_X1 U15109 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n12928), .S(n12871), .Z(
        P2_U3549) );
  MUX2_X1 U15110 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n12959), .S(n12871), .Z(
        P2_U3548) );
  MUX2_X1 U15111 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n12956), .S(n12871), .Z(
        P2_U3547) );
  MUX2_X1 U15112 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n12856), .S(n12871), .Z(
        P2_U3546) );
  MUX2_X1 U15113 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n12857), .S(n12871), .Z(
        P2_U3545) );
  MUX2_X1 U15114 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n12858), .S(n12871), .Z(
        P2_U3544) );
  MUX2_X1 U15115 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n12859), .S(n12871), .Z(
        P2_U3543) );
  MUX2_X1 U15116 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n12860), .S(n12871), .Z(
        P2_U3542) );
  MUX2_X1 U15117 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n12861), .S(n12871), .Z(
        P2_U3541) );
  MUX2_X1 U15118 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n12862), .S(n12871), .Z(
        P2_U3540) );
  MUX2_X1 U15119 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n12863), .S(n12871), .Z(
        P2_U3539) );
  MUX2_X1 U15120 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n12864), .S(n12871), .Z(
        P2_U3538) );
  MUX2_X1 U15121 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n12865), .S(n12871), .Z(
        P2_U3537) );
  MUX2_X1 U15122 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n12866), .S(n12871), .Z(
        P2_U3536) );
  MUX2_X1 U15123 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n12867), .S(n12871), .Z(
        P2_U3535) );
  MUX2_X1 U15124 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n12868), .S(n12871), .Z(
        P2_U3534) );
  MUX2_X1 U15125 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n12869), .S(n12871), .Z(
        P2_U3533) );
  MUX2_X1 U15126 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n12870), .S(n12871), .Z(
        P2_U3532) );
  MUX2_X1 U15127 ( .A(P2_DATAO_REG_0__SCAN_IN), .B(n12872), .S(n12871), .Z(
        P2_U3531) );
  OAI21_X1 U15128 ( .B1(n11367), .B2(n12874), .A(n12873), .ZN(n14803) );
  MUX2_X1 U15129 ( .A(P2_REG2_REG_17__SCAN_IN), .B(n12875), .S(n14804), .Z(
        n14802) );
  NAND2_X1 U15130 ( .A1(n14803), .A2(n14802), .ZN(n14801) );
  XNOR2_X1 U15131 ( .A(n12890), .B(n12891), .ZN(n12877) );
  NOR2_X1 U15132 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12877), .ZN(n12893) );
  AOI21_X1 U15133 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12877), .A(n12893), 
        .ZN(n12889) );
  NOR2_X1 U15134 ( .A1(n12878), .A2(n12895), .ZN(n12879) );
  AOI211_X1 U15135 ( .C1(n14799), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n12880), 
        .B(n12879), .ZN(n12888) );
  AOI21_X1 U15136 ( .B1(n12882), .B2(P2_REG1_REG_16__SCAN_IN), .A(n12881), 
        .ZN(n14797) );
  XNOR2_X1 U15137 ( .A(n14804), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n14796) );
  NOR2_X1 U15138 ( .A1(n14797), .A2(n14796), .ZN(n14794) );
  INV_X1 U15139 ( .A(n12883), .ZN(n12886) );
  INV_X1 U15140 ( .A(n12898), .ZN(n12885) );
  OAI211_X1 U15141 ( .C1(P2_REG1_REG_18__SCAN_IN), .C2(n12886), .A(n14765), 
        .B(n12885), .ZN(n12887) );
  OAI211_X1 U15142 ( .C1(n12889), .C2(n14786), .A(n12888), .B(n12887), .ZN(
        P2_U3232) );
  NOR2_X1 U15143 ( .A1(n12891), .A2(n12890), .ZN(n12892) );
  XOR2_X1 U15144 ( .A(n12894), .B(P2_REG2_REG_19__SCAN_IN), .Z(n12901) );
  NOR2_X1 U15145 ( .A1(n12896), .A2(n12895), .ZN(n12897) );
  XNOR2_X1 U15146 ( .A(n12899), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U15147 ( .A1(n12901), .A2(n14800), .B1(n14765), .B2(n12900), .ZN(
        n12905) );
  INV_X1 U15148 ( .A(n12900), .ZN(n12902) );
  MUX2_X1 U15149 ( .A(n12905), .B(n12904), .S(n12903), .Z(n12907) );
  OAI211_X1 U15150 ( .C1(n12908), .C2(n14793), .A(n12907), .B(n12906), .ZN(
        P2_U3233) );
  NAND2_X1 U15151 ( .A1(n13122), .A2(n13139), .ZN(n13118) );
  OR2_X1 U15152 ( .A1(n13230), .A2(n13118), .ZN(n13106) );
  NOR2_X1 U15153 ( .A1(n13226), .A2(n13106), .ZN(n13094) );
  NOR2_X1 U15154 ( .A1(n13185), .A2(n12998), .ZN(n12952) );
  NAND2_X1 U15155 ( .A1(n12952), .A2(n13183), .ZN(n12917) );
  XNOR2_X1 U15156 ( .A(n13180), .B(n12917), .ZN(n12910) );
  NAND2_X1 U15157 ( .A1(n12910), .A2(n14816), .ZN(n13179) );
  NOR2_X1 U15158 ( .A1(n13295), .A2(n12911), .ZN(n12912) );
  NOR2_X1 U15159 ( .A1(n12913), .A2(n12912), .ZN(n12949) );
  NAND2_X1 U15160 ( .A1(n12949), .A2(n12914), .ZN(n13181) );
  NOR2_X1 U15161 ( .A1(n14844), .A2(n13181), .ZN(n12919) );
  NOR2_X1 U15162 ( .A1(n13180), .A2(n14824), .ZN(n12915) );
  AOI211_X1 U15163 ( .C1(n14844), .C2(P2_REG2_REG_31__SCAN_IN), .A(n12919), 
        .B(n12915), .ZN(n12916) );
  OAI21_X1 U15164 ( .B1(n13179), .B2(n14820), .A(n12916), .ZN(P2_U3234) );
  OAI211_X1 U15165 ( .C1(n12952), .C2(n13183), .A(n14816), .B(n12917), .ZN(
        n13182) );
  NOR2_X1 U15166 ( .A1(n13183), .A2(n14824), .ZN(n12918) );
  AOI211_X1 U15167 ( .C1(n14844), .C2(P2_REG2_REG_30__SCAN_IN), .A(n12919), 
        .B(n12918), .ZN(n12920) );
  OAI21_X1 U15168 ( .B1(n14820), .B2(n13182), .A(n12920), .ZN(P2_U3235) );
  NOR2_X1 U15169 ( .A1(n13226), .A2(n12921), .ZN(n13064) );
  NOR2_X1 U15170 ( .A1(n13066), .A2(n13064), .ZN(n12937) );
  NAND2_X1 U15171 ( .A1(n12923), .A2(n12922), .ZN(n12926) );
  OR2_X1 U15172 ( .A1(n13258), .A2(n12924), .ZN(n12925) );
  NAND2_X1 U15173 ( .A1(n12926), .A2(n12925), .ZN(n13164) );
  NOR2_X1 U15174 ( .A1(n13244), .A2(n12930), .ZN(n12929) );
  NAND2_X1 U15175 ( .A1(n13244), .A2(n12930), .ZN(n12931) );
  NAND2_X1 U15176 ( .A1(n13124), .A2(n13125), .ZN(n13123) );
  NAND2_X1 U15177 ( .A1(n13123), .A2(n12933), .ZN(n13110) );
  OR2_X1 U15178 ( .A1(n13230), .A2(n12935), .ZN(n12934) );
  NAND2_X1 U15179 ( .A1(n13230), .A2(n12935), .ZN(n12936) );
  INV_X1 U15180 ( .A(n12938), .ZN(n12939) );
  INV_X1 U15181 ( .A(n13016), .ZN(n13006) );
  NAND2_X1 U15182 ( .A1(n12949), .A2(n12948), .ZN(n12950) );
  AOI211_X1 U15183 ( .C1(n13185), .C2(n12998), .A(n13169), .B(n12952), .ZN(
        n13184) );
  AOI22_X1 U15184 ( .A1(n12953), .A2(n14839), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n14844), .ZN(n12954) );
  OAI21_X1 U15185 ( .B1(n12955), .B2(n14824), .A(n12954), .ZN(n12989) );
  INV_X1 U15186 ( .A(n13066), .ZN(n13073) );
  INV_X1 U15187 ( .A(n13109), .ZN(n12971) );
  NOR2_X1 U15188 ( .A1(n13174), .A2(n12958), .ZN(n12960) );
  NAND2_X1 U15189 ( .A1(n13155), .A2(n12961), .ZN(n12962) );
  AND2_X1 U15190 ( .A1(n13244), .A2(n12964), .ZN(n12965) );
  NOR2_X1 U15191 ( .A1(n13122), .A2(n12967), .ZN(n12966) );
  NAND2_X1 U15192 ( .A1(n13122), .A2(n12967), .ZN(n12968) );
  NOR2_X1 U15193 ( .A1(n13230), .A2(n12969), .ZN(n12970) );
  NAND2_X1 U15194 ( .A1(n13091), .A2(n13092), .ZN(n13090) );
  NAND2_X1 U15195 ( .A1(n13226), .A2(n12972), .ZN(n12973) );
  NAND2_X1 U15196 ( .A1(n13090), .A2(n12973), .ZN(n13072) );
  NAND2_X1 U15197 ( .A1(n13220), .A2(n12974), .ZN(n12975) );
  OR2_X1 U15198 ( .A1(n13054), .A2(n12977), .ZN(n12978) );
  NAND2_X1 U15199 ( .A1(n13039), .A2(n12980), .ZN(n12979) );
  OR2_X1 U15200 ( .A1(n13039), .A2(n12980), .ZN(n12981) );
  NOR2_X1 U15201 ( .A1(n13028), .A2(n12983), .ZN(n12982) );
  NAND2_X1 U15202 ( .A1(n13028), .A2(n12983), .ZN(n12984) );
  NAND2_X1 U15203 ( .A1(n12992), .A2(n12994), .ZN(n12991) );
  OAI21_X1 U15204 ( .B1(n13187), .B2(n14844), .A(n12990), .ZN(P2_U3236) );
  OAI21_X1 U15205 ( .B1(n12992), .B2(n12994), .A(n12991), .ZN(n13193) );
  AOI21_X1 U15206 ( .B1(n6696), .B2(n12994), .A(n14834), .ZN(n12997) );
  AOI21_X1 U15207 ( .B1(n12997), .B2(n12996), .A(n12995), .ZN(n13192) );
  INV_X1 U15208 ( .A(n12998), .ZN(n12999) );
  AOI211_X1 U15209 ( .C1(n13190), .C2(n6955), .A(n13169), .B(n12999), .ZN(
        n13189) );
  AOI22_X1 U15210 ( .A1(n13189), .A2(n13001), .B1(n14839), .B2(n13000), .ZN(
        n13002) );
  AOI21_X1 U15211 ( .B1(n13192), .B2(n13002), .A(n14844), .ZN(n13003) );
  INV_X1 U15212 ( .A(n13003), .ZN(n13005) );
  AOI22_X1 U15213 ( .A1(n13190), .A2(n13141), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n14844), .ZN(n13004) );
  OAI211_X1 U15214 ( .C1(n13178), .C2(n13193), .A(n13005), .B(n13004), .ZN(
        P2_U3237) );
  XNOR2_X1 U15215 ( .A(n13007), .B(n13006), .ZN(n13009) );
  AOI21_X1 U15216 ( .B1(n13009), .B2(n14814), .A(n13008), .ZN(n13200) );
  AND2_X1 U15217 ( .A1(n13196), .A2(n13023), .ZN(n13010) );
  OR3_X1 U15218 ( .A1(n13011), .A2(n13010), .A3(n13169), .ZN(n13199) );
  AOI22_X1 U15219 ( .A1(n13012), .A2(n14839), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n14844), .ZN(n13014) );
  NAND2_X1 U15220 ( .A1(n13196), .A2(n13141), .ZN(n13013) );
  OAI211_X1 U15221 ( .C1(n13199), .C2(n14820), .A(n13014), .B(n13013), .ZN(
        n13015) );
  INV_X1 U15222 ( .A(n13015), .ZN(n13019) );
  OR2_X1 U15223 ( .A1(n13017), .A2(n13016), .ZN(n13195) );
  NAND3_X1 U15224 ( .A1(n13195), .A2(n13194), .A3(n14828), .ZN(n13018) );
  OAI211_X1 U15225 ( .C1(n13200), .C2(n14844), .A(n13019), .B(n13018), .ZN(
        P2_U3238) );
  XOR2_X1 U15226 ( .A(n13030), .B(n13020), .Z(n13022) );
  AOI21_X1 U15227 ( .B1(n13022), .B2(n14814), .A(n13021), .ZN(n13204) );
  INV_X1 U15228 ( .A(n13040), .ZN(n13025) );
  INV_X1 U15229 ( .A(n13023), .ZN(n13024) );
  AOI211_X1 U15230 ( .C1(n13202), .C2(n13025), .A(n13169), .B(n13024), .ZN(
        n13201) );
  AOI22_X1 U15231 ( .A1(n13026), .A2(n14839), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n14844), .ZN(n13027) );
  OAI21_X1 U15232 ( .B1(n13028), .B2(n14824), .A(n13027), .ZN(n13032) );
  XOR2_X1 U15233 ( .A(n13030), .B(n13029), .Z(n13205) );
  NOR2_X1 U15234 ( .A1(n13205), .A2(n13178), .ZN(n13031) );
  AOI211_X1 U15235 ( .C1(n13201), .C2(n14507), .A(n13032), .B(n13031), .ZN(
        n13033) );
  OAI21_X1 U15236 ( .B1(n14844), .B2(n13204), .A(n13033), .ZN(P2_U3239) );
  XNOR2_X1 U15237 ( .A(n13034), .B(n13037), .ZN(n13036) );
  AOI21_X1 U15238 ( .B1(n13036), .B2(n14814), .A(n13035), .ZN(n13210) );
  XOR2_X1 U15239 ( .A(n13037), .B(n13038), .Z(n13211) );
  INV_X1 U15240 ( .A(n13211), .ZN(n13047) );
  NOR2_X1 U15241 ( .A1(n13039), .A2(n13055), .ZN(n13041) );
  INV_X1 U15242 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13042) );
  OAI22_X1 U15243 ( .A1(n13043), .A2(n14819), .B1(n13042), .B2(n14515), .ZN(
        n13044) );
  AOI21_X1 U15244 ( .B1(n13208), .B2(n13141), .A(n13044), .ZN(n13045) );
  OAI21_X1 U15245 ( .B1(n13206), .B2(n14820), .A(n13045), .ZN(n13046) );
  AOI21_X1 U15246 ( .B1(n13047), .B2(n14828), .A(n13046), .ZN(n13048) );
  OAI21_X1 U15247 ( .B1(n13210), .B2(n14844), .A(n13048), .ZN(P2_U3240) );
  XNOR2_X1 U15248 ( .A(n13049), .B(n12976), .ZN(n13051) );
  AOI21_X1 U15249 ( .B1(n13051), .B2(n14814), .A(n13050), .ZN(n13216) );
  OAI21_X1 U15250 ( .B1(n6488), .B2(n13053), .A(n13052), .ZN(n13217) );
  INV_X1 U15251 ( .A(n13217), .ZN(n13062) );
  NOR2_X1 U15252 ( .A1(n13054), .A2(n13077), .ZN(n13056) );
  OAI22_X1 U15253 ( .A1(n13058), .A2(n14819), .B1(n14515), .B2(n13057), .ZN(
        n13059) );
  AOI21_X1 U15254 ( .B1(n13214), .B2(n13141), .A(n13059), .ZN(n13060) );
  OAI21_X1 U15255 ( .B1(n13212), .B2(n14820), .A(n13060), .ZN(n13061) );
  AOI21_X1 U15256 ( .B1(n13062), .B2(n14828), .A(n13061), .ZN(n13063) );
  OAI21_X1 U15257 ( .B1(n13216), .B2(n14844), .A(n13063), .ZN(P2_U3241) );
  INV_X1 U15258 ( .A(n13064), .ZN(n13065) );
  NAND2_X1 U15259 ( .A1(n13089), .A2(n13065), .ZN(n13067) );
  AND2_X1 U15260 ( .A1(n13067), .A2(n13066), .ZN(n13068) );
  OAI21_X1 U15261 ( .B1(n13069), .B2(n13068), .A(n14814), .ZN(n13071) );
  NAND2_X1 U15262 ( .A1(n13071), .A2(n13070), .ZN(n13223) );
  INV_X1 U15263 ( .A(n13223), .ZN(n13085) );
  NAND2_X1 U15264 ( .A1(n13073), .A2(n13072), .ZN(n13074) );
  NAND2_X1 U15265 ( .A1(n13075), .A2(n13074), .ZN(n13218) );
  NOR2_X1 U15266 ( .A1(n13220), .A2(n13094), .ZN(n13076) );
  OAI22_X1 U15267 ( .A1(n14515), .A2(n13079), .B1(n13078), .B2(n14819), .ZN(
        n13080) );
  AOI21_X1 U15268 ( .B1(n13081), .B2(n13141), .A(n13080), .ZN(n13082) );
  OAI21_X1 U15269 ( .B1(n13219), .B2(n14820), .A(n13082), .ZN(n13083) );
  AOI21_X1 U15270 ( .B1(n14828), .B2(n13218), .A(n13083), .ZN(n13084) );
  OAI21_X1 U15271 ( .B1(n13085), .B2(n14844), .A(n13084), .ZN(P2_U3242) );
  AOI21_X1 U15272 ( .B1(n13086), .B2(n13092), .A(n14834), .ZN(n13088) );
  AOI21_X1 U15273 ( .B1(n13089), .B2(n13088), .A(n13087), .ZN(n13228) );
  OAI21_X1 U15274 ( .B1(n13092), .B2(n13091), .A(n13090), .ZN(n13229) );
  INV_X1 U15275 ( .A(n13229), .ZN(n13099) );
  AND2_X1 U15276 ( .A1(n13226), .A2(n13106), .ZN(n13093) );
  OR3_X1 U15277 ( .A1(n13094), .A2(n13093), .A3(n13169), .ZN(n13224) );
  AOI22_X1 U15278 ( .A1(n13095), .A2(n14839), .B1(n14844), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n13097) );
  NAND2_X1 U15279 ( .A1(n13226), .A2(n13141), .ZN(n13096) );
  OAI211_X1 U15280 ( .C1(n13224), .C2(n14820), .A(n13097), .B(n13096), .ZN(
        n13098) );
  AOI21_X1 U15281 ( .B1(n13099), .B2(n14828), .A(n13098), .ZN(n13100) );
  OAI21_X1 U15282 ( .B1(n13228), .B2(n14844), .A(n13100), .ZN(P2_U3243) );
  XNOR2_X1 U15283 ( .A(n13109), .B(n13101), .ZN(n13233) );
  INV_X1 U15284 ( .A(n13102), .ZN(n13103) );
  OAI22_X1 U15285 ( .A1(n14515), .A2(n13104), .B1(n13103), .B2(n14819), .ZN(
        n13108) );
  NAND2_X1 U15286 ( .A1(n13230), .A2(n13118), .ZN(n13105) );
  NAND3_X1 U15287 ( .A1(n13106), .A2(n14816), .A3(n13105), .ZN(n13232) );
  NOR2_X1 U15288 ( .A1(n13232), .A2(n14820), .ZN(n13107) );
  AOI211_X1 U15289 ( .C1(n13141), .C2(n13230), .A(n13108), .B(n13107), .ZN(
        n13115) );
  XNOR2_X1 U15290 ( .A(n13110), .B(n13109), .ZN(n13111) );
  NAND2_X1 U15291 ( .A1(n13111), .A2(n14814), .ZN(n13113) );
  NAND2_X1 U15292 ( .A1(n13113), .A2(n13112), .ZN(n13235) );
  NAND2_X1 U15293 ( .A1(n13235), .A2(n14515), .ZN(n13114) );
  OAI211_X1 U15294 ( .C1(n13178), .C2(n13233), .A(n13115), .B(n13114), .ZN(
        P2_U3244) );
  XOR2_X1 U15295 ( .A(n13116), .B(n13125), .Z(n13240) );
  OR2_X1 U15296 ( .A1(n13122), .A2(n13139), .ZN(n13117) );
  AND3_X1 U15297 ( .A1(n13118), .A2(n13117), .A3(n14816), .ZN(n13236) );
  NOR2_X1 U15298 ( .A1(n13119), .A2(n14819), .ZN(n13120) );
  AOI21_X1 U15299 ( .B1(n14844), .B2(P2_REG2_REG_20__SCAN_IN), .A(n13120), 
        .ZN(n13121) );
  OAI21_X1 U15300 ( .B1(n13122), .B2(n14824), .A(n13121), .ZN(n13129) );
  OAI21_X1 U15301 ( .B1(n13125), .B2(n13124), .A(n13123), .ZN(n13127) );
  AOI21_X1 U15302 ( .B1(n13127), .B2(n14814), .A(n13126), .ZN(n13239) );
  NOR2_X1 U15303 ( .A1(n13239), .A2(n14844), .ZN(n13128) );
  AOI211_X1 U15304 ( .C1(n13236), .C2(n14507), .A(n13129), .B(n13128), .ZN(
        n13130) );
  OAI21_X1 U15305 ( .B1(n13178), .B2(n13240), .A(n13130), .ZN(P2_U3245) );
  XNOR2_X1 U15306 ( .A(n13131), .B(n13135), .ZN(n13132) );
  NAND2_X1 U15307 ( .A1(n13132), .A2(n14814), .ZN(n13134) );
  NAND2_X1 U15308 ( .A1(n13134), .A2(n13133), .ZN(n13246) );
  INV_X1 U15309 ( .A(n13246), .ZN(n13146) );
  INV_X1 U15310 ( .A(n13135), .ZN(n13136) );
  XNOR2_X1 U15311 ( .A(n13137), .B(n13136), .ZN(n13241) );
  NOR2_X1 U15312 ( .A1(n13244), .A2(n13150), .ZN(n13138) );
  AOI22_X1 U15313 ( .A1(n14844), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n13140), 
        .B2(n14839), .ZN(n13143) );
  NAND2_X1 U15314 ( .A1(n6949), .A2(n13141), .ZN(n13142) );
  OAI211_X1 U15315 ( .C1(n13242), .C2(n14820), .A(n13143), .B(n13142), .ZN(
        n13144) );
  AOI21_X1 U15316 ( .B1(n13241), .B2(n14828), .A(n13144), .ZN(n13145) );
  OAI21_X1 U15317 ( .B1(n13146), .B2(n14844), .A(n13145), .ZN(P2_U3246) );
  XOR2_X1 U15318 ( .A(n13147), .B(n13157), .Z(n13149) );
  AOI21_X1 U15319 ( .B1(n13149), .B2(n14814), .A(n13148), .ZN(n13250) );
  INV_X1 U15320 ( .A(n13171), .ZN(n13151) );
  AOI211_X1 U15321 ( .C1(n13248), .C2(n13151), .A(n13169), .B(n13150), .ZN(
        n13247) );
  INV_X1 U15322 ( .A(n13152), .ZN(n13153) );
  AOI22_X1 U15323 ( .A1(n14844), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n13153), 
        .B2(n14839), .ZN(n13154) );
  OAI21_X1 U15324 ( .B1(n13155), .B2(n14824), .A(n13154), .ZN(n13159) );
  XOR2_X1 U15325 ( .A(n13157), .B(n13156), .Z(n13251) );
  NOR2_X1 U15326 ( .A1(n13251), .A2(n13178), .ZN(n13158) );
  AOI211_X1 U15327 ( .C1(n13247), .C2(n14507), .A(n13159), .B(n13158), .ZN(
        n13160) );
  OAI21_X1 U15328 ( .B1(n14844), .B2(n13250), .A(n13160), .ZN(P2_U3247) );
  XNOR2_X1 U15329 ( .A(n13161), .B(n13165), .ZN(n13257) );
  INV_X1 U15330 ( .A(n13162), .ZN(n13163) );
  AOI21_X1 U15331 ( .B1(n13165), .B2(n13164), .A(n13163), .ZN(n13167) );
  OAI21_X1 U15332 ( .B1(n13167), .B2(n14834), .A(n13166), .ZN(n13253) );
  NOR2_X1 U15333 ( .A1(n13174), .A2(n13168), .ZN(n13170) );
  NOR2_X1 U15334 ( .A1(n13252), .A2(n14820), .ZN(n13176) );
  AOI22_X1 U15335 ( .A1(n14844), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13172), 
        .B2(n14839), .ZN(n13173) );
  OAI21_X1 U15336 ( .B1(n13174), .B2(n14824), .A(n13173), .ZN(n13175) );
  AOI211_X1 U15337 ( .C1(n13253), .C2(n14515), .A(n13176), .B(n13175), .ZN(
        n13177) );
  OAI21_X1 U15338 ( .B1(n13178), .B2(n13257), .A(n13177), .ZN(P2_U3248) );
  OAI211_X1 U15339 ( .C1(n13180), .C2(n14933), .A(n13179), .B(n13181), .ZN(
        n13265) );
  MUX2_X1 U15340 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13265), .S(n14970), .Z(
        P2_U3530) );
  OAI211_X1 U15341 ( .C1(n13183), .C2(n14933), .A(n13182), .B(n13181), .ZN(
        n13266) );
  MUX2_X1 U15342 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13266), .S(n14970), .Z(
        P2_U3529) );
  AOI21_X1 U15343 ( .B1(n14943), .B2(n13185), .A(n13184), .ZN(n13186) );
  AOI21_X1 U15344 ( .B1(n14943), .B2(n13190), .A(n13189), .ZN(n13191) );
  OAI211_X1 U15345 ( .C1(n13261), .C2(n13193), .A(n13192), .B(n13191), .ZN(
        n13268) );
  MUX2_X1 U15346 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13268), .S(n14970), .Z(
        P2_U3527) );
  NAND3_X1 U15347 ( .A1(n13195), .A2(n14913), .A3(n13194), .ZN(n13198) );
  NAND2_X1 U15348 ( .A1(n13196), .A2(n14943), .ZN(n13197) );
  NAND4_X1 U15349 ( .A1(n13200), .A2(n13199), .A3(n13198), .A4(n13197), .ZN(
        n13269) );
  MUX2_X1 U15350 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13269), .S(n14970), .Z(
        P2_U3526) );
  AOI21_X1 U15351 ( .B1(n14943), .B2(n13202), .A(n13201), .ZN(n13203) );
  OAI211_X1 U15352 ( .C1(n13261), .C2(n13205), .A(n13204), .B(n13203), .ZN(
        n13270) );
  MUX2_X1 U15353 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13270), .S(n14970), .Z(
        P2_U3525) );
  INV_X1 U15354 ( .A(n13206), .ZN(n13207) );
  AOI21_X1 U15355 ( .B1(n14943), .B2(n13208), .A(n13207), .ZN(n13209) );
  OAI211_X1 U15356 ( .C1(n13261), .C2(n13211), .A(n13210), .B(n13209), .ZN(
        n13271) );
  MUX2_X1 U15357 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13271), .S(n14970), .Z(
        P2_U3524) );
  INV_X1 U15358 ( .A(n13212), .ZN(n13213) );
  AOI21_X1 U15359 ( .B1(n14943), .B2(n13214), .A(n13213), .ZN(n13215) );
  OAI211_X1 U15360 ( .C1(n13261), .C2(n13217), .A(n13216), .B(n13215), .ZN(
        n13272) );
  MUX2_X1 U15361 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13272), .S(n14970), .Z(
        P2_U3523) );
  AND2_X1 U15362 ( .A1(n13218), .A2(n14913), .ZN(n13222) );
  OAI21_X1 U15363 ( .B1(n13220), .B2(n14933), .A(n13219), .ZN(n13221) );
  MUX2_X1 U15364 ( .A(n13273), .B(P2_REG1_REG_23__SCAN_IN), .S(n14968), .Z(
        P2_U3522) );
  INV_X1 U15365 ( .A(n13224), .ZN(n13225) );
  AOI21_X1 U15366 ( .B1(n14943), .B2(n13226), .A(n13225), .ZN(n13227) );
  OAI211_X1 U15367 ( .C1(n13261), .C2(n13229), .A(n13228), .B(n13227), .ZN(
        n13274) );
  MUX2_X1 U15368 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13274), .S(n14970), .Z(
        P2_U3521) );
  NAND2_X1 U15369 ( .A1(n13230), .A2(n14943), .ZN(n13231) );
  OAI211_X1 U15370 ( .C1(n13233), .C2(n13261), .A(n13232), .B(n13231), .ZN(
        n13234) );
  MUX2_X1 U15371 ( .A(n13275), .B(P2_REG1_REG_21__SCAN_IN), .S(n14968), .Z(
        P2_U3520) );
  AOI21_X1 U15372 ( .B1(n14943), .B2(n13237), .A(n13236), .ZN(n13238) );
  OAI211_X1 U15373 ( .C1(n13261), .C2(n13240), .A(n13239), .B(n13238), .ZN(
        n13276) );
  MUX2_X1 U15374 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13276), .S(n14970), .Z(
        P2_U3519) );
  NAND2_X1 U15375 ( .A1(n13241), .A2(n14913), .ZN(n13243) );
  OAI211_X1 U15376 ( .C1(n13244), .C2(n14933), .A(n13243), .B(n13242), .ZN(
        n13245) );
  MUX2_X1 U15377 ( .A(n13277), .B(P2_REG1_REG_19__SCAN_IN), .S(n14968), .Z(
        P2_U3518) );
  AOI21_X1 U15378 ( .B1(n14943), .B2(n13248), .A(n13247), .ZN(n13249) );
  OAI211_X1 U15379 ( .C1(n13261), .C2(n13251), .A(n13250), .B(n13249), .ZN(
        n13278) );
  MUX2_X1 U15380 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13278), .S(n14970), .Z(
        P2_U3517) );
  INV_X1 U15381 ( .A(n13252), .ZN(n13254) );
  AOI211_X1 U15382 ( .C1(n14943), .C2(n13255), .A(n13254), .B(n13253), .ZN(
        n13256) );
  OAI21_X1 U15383 ( .B1(n13261), .B2(n13257), .A(n13256), .ZN(n13279) );
  MUX2_X1 U15384 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13279), .S(n14970), .Z(
        P2_U3516) );
  NAND2_X1 U15385 ( .A1(n13258), .A2(n14943), .ZN(n13259) );
  OAI211_X1 U15386 ( .C1(n13262), .C2(n13261), .A(n13260), .B(n13259), .ZN(
        n13263) );
  OR2_X1 U15387 ( .A1(n13264), .A2(n13263), .ZN(n13280) );
  MUX2_X1 U15388 ( .A(n13280), .B(P2_REG1_REG_16__SCAN_IN), .S(n14968), .Z(
        P2_U3515) );
  MUX2_X1 U15389 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13265), .S(n14952), .Z(
        P2_U3498) );
  MUX2_X1 U15390 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13266), .S(n14952), .Z(
        P2_U3497) );
  MUX2_X1 U15391 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13267), .S(n14952), .Z(
        P2_U3496) );
  MUX2_X1 U15392 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n13268), .S(n14952), .Z(
        P2_U3495) );
  MUX2_X1 U15393 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13269), .S(n14952), .Z(
        P2_U3494) );
  MUX2_X1 U15394 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13270), .S(n14952), .Z(
        P2_U3493) );
  MUX2_X1 U15395 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13271), .S(n14952), .Z(
        P2_U3492) );
  MUX2_X1 U15396 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13272), .S(n14952), .Z(
        P2_U3491) );
  MUX2_X1 U15397 ( .A(n13273), .B(P2_REG0_REG_23__SCAN_IN), .S(n14950), .Z(
        P2_U3490) );
  MUX2_X1 U15398 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13274), .S(n14952), .Z(
        P2_U3489) );
  MUX2_X1 U15399 ( .A(n13275), .B(P2_REG0_REG_21__SCAN_IN), .S(n14950), .Z(
        P2_U3488) );
  MUX2_X1 U15400 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13276), .S(n14952), .Z(
        P2_U3487) );
  MUX2_X1 U15401 ( .A(n13277), .B(P2_REG0_REG_19__SCAN_IN), .S(n14950), .Z(
        P2_U3486) );
  MUX2_X1 U15402 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13278), .S(n14952), .Z(
        P2_U3484) );
  MUX2_X1 U15403 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13279), .S(n14952), .Z(
        P2_U3481) );
  MUX2_X1 U15404 ( .A(n13280), .B(P2_REG0_REG_16__SCAN_IN), .S(n14950), .Z(
        P2_U3478) );
  INV_X1 U15405 ( .A(n13437), .ZN(n14239) );
  NAND2_X1 U15406 ( .A1(n14239), .A2(n13289), .ZN(n13284) );
  OR4_X1 U15407 ( .A1(n13282), .A2(P2_IR_REG_30__SCAN_IN), .A3(n13281), .A4(
        P2_U3088), .ZN(n13283) );
  OAI211_X1 U15408 ( .C1(n9065), .C2(n13303), .A(n13284), .B(n13283), .ZN(
        P2_U3296) );
  OAI222_X1 U15409 ( .A1(n13301), .A2(n13288), .B1(P2_U3088), .B2(n13286), 
        .C1(n13285), .C2(n13303), .ZN(P2_U3298) );
  NAND2_X1 U15410 ( .A1(n11975), .A2(n13289), .ZN(n13291) );
  OAI211_X1 U15411 ( .C1(n13303), .C2(n13292), .A(n13291), .B(n13290), .ZN(
        P2_U3299) );
  INV_X1 U15412 ( .A(n13293), .ZN(n14243) );
  OAI222_X1 U15413 ( .A1(n13295), .A2(P2_U3088), .B1(n13301), .B2(n14243), 
        .C1(n13294), .C2(n13303), .ZN(P2_U3300) );
  INV_X1 U15414 ( .A(n13296), .ZN(n14246) );
  OAI222_X1 U15415 ( .A1(P2_U3088), .A2(n13298), .B1(n13301), .B2(n14246), 
        .C1(n13297), .C2(n13303), .ZN(P2_U3301) );
  INV_X1 U15416 ( .A(n13299), .ZN(n14250) );
  OAI222_X1 U15417 ( .A1(n13303), .A2(n13302), .B1(n13301), .B2(n14250), .C1(
        P2_U3088), .C2(n13300), .ZN(P2_U3302) );
  INV_X1 U15418 ( .A(n13304), .ZN(n13305) );
  MUX2_X1 U15419 ( .A(n13305), .B(n14739), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3327) );
  XOR2_X1 U15420 ( .A(n13307), .B(n13306), .Z(n13314) );
  NOR2_X1 U15421 ( .A1(n14580), .A2(n13308), .ZN(n13312) );
  AOI22_X1 U15422 ( .A1(n13418), .A2(n13888), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13309) );
  OAI21_X1 U15423 ( .B1(n13310), .B2(n14562), .A(n13309), .ZN(n13311) );
  AOI211_X1 U15424 ( .C1(n14115), .C2(n14576), .A(n13312), .B(n13311), .ZN(
        n13313) );
  OAI21_X1 U15425 ( .B1(n13314), .B2(n14570), .A(n13313), .ZN(P1_U3214) );
  XOR2_X1 U15426 ( .A(n13316), .B(n13315), .Z(n13321) );
  NOR2_X1 U15427 ( .A1(n14580), .A2(n13971), .ZN(n13319) );
  AOI22_X1 U15428 ( .A1(n13418), .A2(n13983), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13317) );
  OAI21_X1 U15429 ( .B1(n13331), .B2(n14562), .A(n13317), .ZN(n13318) );
  AOI211_X1 U15430 ( .C1(n13978), .C2(n14576), .A(n13319), .B(n13318), .ZN(
        n13320) );
  OAI21_X1 U15431 ( .B1(n13321), .B2(n14570), .A(n13320), .ZN(P1_U3216) );
  OAI211_X1 U15432 ( .C1(n13324), .C2(n13323), .A(n13322), .B(n14553), .ZN(
        n13328) );
  OAI22_X1 U15433 ( .A1(n13522), .A2(n14060), .B1(n13372), .B2(n14020), .ZN(
        n14162) );
  NOR2_X1 U15434 ( .A1(n13325), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13857) );
  NOR2_X1 U15435 ( .A1(n14580), .A2(n14045), .ZN(n13326) );
  AOI211_X1 U15436 ( .C1(n14162), .C2(n13332), .A(n13857), .B(n13326), .ZN(
        n13327) );
  OAI211_X1 U15437 ( .C1(n14228), .C2(n13434), .A(n13328), .B(n13327), .ZN(
        P1_U3219) );
  AOI21_X1 U15438 ( .B1(n13330), .B2(n13329), .A(n6530), .ZN(n13337) );
  INV_X1 U15439 ( .A(n14013), .ZN(n13334) );
  OAI22_X1 U15440 ( .A1(n13522), .A2(n14020), .B1(n13331), .B2(n14060), .ZN(
        n14005) );
  AOI22_X1 U15441 ( .A1(n14005), .A2(n13332), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13333) );
  OAI21_X1 U15442 ( .B1(n13334), .B2(n14580), .A(n13333), .ZN(n13335) );
  AOI21_X1 U15443 ( .B1(n14010), .B2(n14576), .A(n13335), .ZN(n13336) );
  OAI21_X1 U15444 ( .B1(n13337), .B2(n14570), .A(n13336), .ZN(P1_U3223) );
  INV_X1 U15445 ( .A(n13601), .ZN(n14383) );
  AOI21_X1 U15446 ( .B1(n13339), .B2(n13338), .A(n14570), .ZN(n13341) );
  NAND2_X1 U15447 ( .A1(n13341), .A2(n13340), .ZN(n13348) );
  OAI21_X1 U15448 ( .B1(n14562), .B2(n13343), .A(n13342), .ZN(n13346) );
  NOR2_X1 U15449 ( .A1(n14580), .A2(n13344), .ZN(n13345) );
  AOI211_X1 U15450 ( .C1(n13418), .C2(n13739), .A(n13346), .B(n13345), .ZN(
        n13347) );
  OAI211_X1 U15451 ( .C1(n14383), .C2(n13434), .A(n13348), .B(n13347), .ZN(
        P1_U3224) );
  XOR2_X1 U15452 ( .A(n13350), .B(n13349), .Z(n13356) );
  AND2_X1 U15453 ( .A1(n13943), .A2(n14712), .ZN(n14127) );
  NOR2_X1 U15454 ( .A1(n14580), .A2(n13941), .ZN(n13354) );
  AOI22_X1 U15455 ( .A1(n13418), .A2(n13934), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13351) );
  OAI21_X1 U15456 ( .B1(n13352), .B2(n14562), .A(n13351), .ZN(n13353) );
  AOI211_X1 U15457 ( .C1(n14127), .C2(n13422), .A(n13354), .B(n13353), .ZN(
        n13355) );
  OAI21_X1 U15458 ( .B1(n13356), .B2(n14570), .A(n13355), .ZN(P1_U3225) );
  INV_X1 U15459 ( .A(n13357), .ZN(n13358) );
  AOI21_X1 U15460 ( .B1(n13360), .B2(n13359), .A(n13358), .ZN(n13365) );
  AOI22_X1 U15461 ( .A1(n13409), .A2(n14086), .B1(P1_REG3_REG_16__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13362) );
  NAND2_X1 U15462 ( .A1(n13418), .A2(n14084), .ZN(n13361) );
  OAI211_X1 U15463 ( .C1(n14580), .C2(n14077), .A(n13362), .B(n13361), .ZN(
        n13363) );
  AOI21_X1 U15464 ( .B1(n14188), .B2(n14576), .A(n13363), .ZN(n13364) );
  OAI21_X1 U15465 ( .B1(n13365), .B2(n14570), .A(n13364), .ZN(P1_U3226) );
  OAI21_X1 U15466 ( .B1(n13368), .B2(n13367), .A(n13366), .ZN(n13369) );
  NAND2_X1 U15467 ( .A1(n13369), .A2(n14553), .ZN(n13376) );
  NOR2_X1 U15468 ( .A1(n13370), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13809) );
  AOI21_X1 U15469 ( .B1(n13409), .B2(n13737), .A(n13809), .ZN(n13371) );
  OAI21_X1 U15470 ( .B1(n13372), .B2(n14565), .A(n13371), .ZN(n13373) );
  AOI21_X1 U15471 ( .B1(n13374), .B2(n13430), .A(n13373), .ZN(n13375) );
  OAI211_X1 U15472 ( .C1(n14181), .C2(n13434), .A(n13376), .B(n13375), .ZN(
        P1_U3228) );
  XOR2_X1 U15473 ( .A(n13378), .B(n13377), .Z(n13383) );
  NOR2_X1 U15474 ( .A1(n14580), .A2(n13962), .ZN(n13381) );
  AOI22_X1 U15475 ( .A1(n13418), .A2(n13731), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13379) );
  OAI21_X1 U15476 ( .B1(n13990), .B2(n14562), .A(n13379), .ZN(n13380) );
  AOI211_X1 U15477 ( .C1(n13961), .C2(n14576), .A(n13381), .B(n13380), .ZN(
        n13382) );
  OAI21_X1 U15478 ( .B1(n13383), .B2(n14570), .A(n13382), .ZN(P1_U3229) );
  OAI211_X1 U15479 ( .C1(n13386), .C2(n13385), .A(n13384), .B(n14553), .ZN(
        n13390) );
  AOI22_X1 U15480 ( .A1(n13735), .A2(n13409), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13387) );
  OAI21_X1 U15481 ( .B1(n14021), .B2(n14565), .A(n13387), .ZN(n13388) );
  AOI21_X1 U15482 ( .B1(n14026), .B2(n13430), .A(n13388), .ZN(n13389) );
  OAI211_X1 U15483 ( .C1(n14028), .C2(n13434), .A(n13390), .B(n13389), .ZN(
        P1_U3233) );
  OAI211_X1 U15484 ( .C1(n13392), .C2(n13391), .A(n14540), .B(n14553), .ZN(
        n13397) );
  NAND2_X1 U15485 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n13797)
         );
  OAI21_X1 U15486 ( .B1(n14562), .B2(n14564), .A(n13797), .ZN(n13395) );
  NOR2_X1 U15487 ( .A1(n14580), .A2(n13393), .ZN(n13394) );
  AOI211_X1 U15488 ( .C1(n13418), .C2(n13738), .A(n13395), .B(n13394), .ZN(
        n13396) );
  OAI211_X1 U15489 ( .C1(n14582), .C2(n13434), .A(n13397), .B(n13396), .ZN(
        P1_U3234) );
  OAI21_X1 U15490 ( .B1(n13400), .B2(n13399), .A(n13398), .ZN(n13401) );
  NAND2_X1 U15491 ( .A1(n13401), .A2(n14553), .ZN(n13406) );
  NOR2_X1 U15492 ( .A1(n14580), .A2(n13992), .ZN(n13404) );
  INV_X1 U15493 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n13402) );
  OAI22_X1 U15494 ( .A1(n14021), .A2(n14562), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13402), .ZN(n13403) );
  AOI211_X1 U15495 ( .C1(n13418), .C2(n13732), .A(n13404), .B(n13403), .ZN(
        n13405) );
  OAI211_X1 U15496 ( .C1(n13434), .C2(n7363), .A(n13406), .B(n13405), .ZN(
        P1_U3235) );
  XOR2_X1 U15497 ( .A(n13408), .B(n13407), .Z(n13414) );
  NAND2_X1 U15498 ( .A1(n13409), .A2(n14084), .ZN(n13410) );
  NAND2_X1 U15499 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13826)
         );
  OAI211_X1 U15500 ( .C1(n14061), .C2(n14565), .A(n13410), .B(n13826), .ZN(
        n13412) );
  NOR2_X1 U15501 ( .A1(n14068), .A2(n13434), .ZN(n13411) );
  AOI211_X1 U15502 ( .C1(n13430), .C2(n14066), .A(n13412), .B(n13411), .ZN(
        n13413) );
  OAI21_X1 U15503 ( .B1(n13414), .B2(n14570), .A(n13413), .ZN(P1_U3238) );
  XOR2_X1 U15504 ( .A(n13416), .B(n13415), .Z(n13424) );
  NOR2_X1 U15505 ( .A1(n13417), .A2(n14587), .ZN(n14122) );
  NOR2_X1 U15506 ( .A1(n14580), .A2(n13921), .ZN(n13421) );
  AOI22_X1 U15507 ( .A1(n13418), .A2(n13903), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13419) );
  OAI21_X1 U15508 ( .B1(n13953), .B2(n14562), .A(n13419), .ZN(n13420) );
  AOI211_X1 U15509 ( .C1(n14122), .C2(n13422), .A(n13421), .B(n13420), .ZN(
        n13423) );
  OAI21_X1 U15510 ( .B1(n13424), .B2(n14570), .A(n13423), .ZN(P1_U3240) );
  OAI211_X1 U15511 ( .C1(n13427), .C2(n13426), .A(n13425), .B(n14553), .ZN(
        n13433) );
  NAND2_X1 U15512 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n14643)
         );
  OAI21_X1 U15513 ( .B1(n13428), .B2(n14552), .A(n14643), .ZN(n13429) );
  AOI21_X1 U15514 ( .B1(n13431), .B2(n13430), .A(n13429), .ZN(n13432) );
  OAI211_X1 U15515 ( .C1(n13435), .C2(n13434), .A(n13433), .B(n13432), .ZN(
        P1_U3241) );
  OR2_X1 U15516 ( .A1(n13464), .A2(n14234), .ZN(n13438) );
  XNOR2_X1 U15517 ( .A(n14254), .B(n13920), .ZN(n13443) );
  NAND2_X1 U15518 ( .A1(n13443), .A2(n13440), .ZN(n13516) );
  NAND2_X1 U15519 ( .A1(n13516), .A2(n13441), .ZN(n13449) );
  NAND2_X1 U15520 ( .A1(n13443), .A2(n13442), .ZN(n13444) );
  NAND2_X1 U15521 ( .A1(n13862), .A2(n6466), .ZN(n13502) );
  NAND2_X1 U15522 ( .A1(n13445), .A2(n13461), .ZN(n13448) );
  OR2_X1 U15523 ( .A1(n13464), .A2(n13446), .ZN(n13447) );
  INV_X1 U15524 ( .A(n13449), .ZN(n13454) );
  INV_X1 U15525 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14204) );
  NAND2_X1 U15526 ( .A1(n6688), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n13452) );
  NAND2_X1 U15527 ( .A1(n13450), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n13451) );
  OAI211_X1 U15528 ( .C1(n6428), .C2(n14204), .A(n13452), .B(n13451), .ZN(
        n13884) );
  OAI21_X1 U15529 ( .B1(n13866), .B2(n13454), .A(n13884), .ZN(n13455) );
  MUX2_X1 U15530 ( .A(n14206), .B(n13455), .S(n6591), .Z(n13710) );
  NOR2_X1 U15531 ( .A1(n13506), .A2(n13710), .ZN(n13460) );
  NAND2_X1 U15532 ( .A1(n13457), .A2(n13456), .ZN(n13458) );
  AND2_X1 U15533 ( .A1(n13459), .A2(n13458), .ZN(n13711) );
  NOR2_X1 U15534 ( .A1(n13711), .A2(n13505), .ZN(n13725) );
  OAI211_X1 U15535 ( .C1(n13866), .C2(n13502), .A(n13460), .B(n13725), .ZN(
        n13721) );
  INV_X1 U15536 ( .A(n13721), .ZN(n13521) );
  XNOR2_X1 U15537 ( .A(n13862), .B(n13866), .ZN(n13724) );
  NAND2_X1 U15538 ( .A1(n13462), .A2(n13461), .ZN(n13466) );
  OR2_X1 U15539 ( .A1(n13464), .A2(n13463), .ZN(n13465) );
  INV_X1 U15540 ( .A(n13902), .ZN(n13467) );
  XNOR2_X1 U15541 ( .A(n13883), .B(n13467), .ZN(n13880) );
  NAND2_X1 U15542 ( .A1(n14111), .A2(n13888), .ZN(n13874) );
  OR2_X1 U15543 ( .A1(n14111), .A2(n13888), .ZN(n13468) );
  NAND2_X1 U15544 ( .A1(n13874), .A2(n13468), .ZN(n13873) );
  NAND4_X1 U15545 ( .A1(n13470), .A2(n13533), .A3(n13469), .A4(n13524), .ZN(
        n13472) );
  NOR2_X1 U15546 ( .A1(n13472), .A2(n13471), .ZN(n13475) );
  NAND4_X1 U15547 ( .A1(n13476), .A2(n13475), .A3(n13474), .A4(n13473), .ZN(
        n13477) );
  NOR2_X1 U15548 ( .A1(n13478), .A2(n13477), .ZN(n13481) );
  NAND4_X1 U15549 ( .A1(n13482), .A2(n13481), .A3(n13480), .A4(n13479), .ZN(
        n13483) );
  OR4_X1 U15550 ( .A1(n11244), .A2(n13485), .A3(n13484), .A4(n13483), .ZN(
        n13486) );
  NOR2_X1 U15551 ( .A1(n13487), .A2(n13486), .ZN(n13488) );
  NAND3_X1 U15552 ( .A1(n13489), .A2(n13488), .A3(n14081), .ZN(n13490) );
  NOR2_X1 U15553 ( .A1(n14040), .A2(n13490), .ZN(n13491) );
  NAND4_X1 U15554 ( .A1(n14008), .A2(n13491), .A3(n14033), .A4(n14056), .ZN(
        n13492) );
  OR4_X1 U15555 ( .A1(n13952), .A2(n13493), .A3(n13996), .A4(n13492), .ZN(
        n13494) );
  NOR2_X1 U15556 ( .A1(n13924), .A2(n13494), .ZN(n13496) );
  NAND4_X1 U15557 ( .A1(n13873), .A2(n13496), .A3(n13495), .A4(n13932), .ZN(
        n13497) );
  NOR2_X1 U15558 ( .A1(n13880), .A2(n13497), .ZN(n13499) );
  INV_X1 U15559 ( .A(n14206), .ZN(n13519) );
  XNOR2_X1 U15560 ( .A(n13519), .B(n13884), .ZN(n13498) );
  NAND3_X1 U15561 ( .A1(n13724), .A2(n13499), .A3(n13498), .ZN(n13500) );
  XNOR2_X1 U15562 ( .A(n13500), .B(n13920), .ZN(n13501) );
  NAND2_X1 U15563 ( .A1(n13501), .A2(n13505), .ZN(n13514) );
  INV_X1 U15564 ( .A(n13711), .ZN(n13507) );
  XNOR2_X1 U15565 ( .A(n13502), .B(n13507), .ZN(n13504) );
  NAND2_X1 U15566 ( .A1(n13504), .A2(n13503), .ZN(n13512) );
  INV_X1 U15567 ( .A(n13505), .ZN(n13511) );
  NAND3_X1 U15568 ( .A1(n13508), .A2(n13866), .A3(n13507), .ZN(n13509) );
  NAND4_X1 U15569 ( .A1(n13512), .A2(n13511), .A3(n13510), .A4(n13509), .ZN(
        n13513) );
  NAND2_X1 U15570 ( .A1(n6466), .A2(n13866), .ZN(n13517) );
  INV_X1 U15571 ( .A(n13884), .ZN(n13515) );
  AOI21_X1 U15572 ( .B1(n13517), .B2(n13516), .A(n13515), .ZN(n13518) );
  AOI21_X1 U15573 ( .B1(n13519), .B2(n7235), .A(n13518), .ZN(n13713) );
  NAND2_X1 U15574 ( .A1(n13713), .A2(n13726), .ZN(n13720) );
  INV_X1 U15575 ( .A(n13720), .ZN(n13520) );
  AOI22_X1 U15576 ( .A1(n13726), .A2(n13521), .B1(n13727), .B2(n13520), .ZN(
        n13730) );
  MUX2_X1 U15577 ( .A(n13982), .B(n13997), .S(n7235), .Z(n13672) );
  MUX2_X1 U15578 ( .A(n13522), .B(n14028), .S(n7235), .Z(n13664) );
  OAI211_X1 U15579 ( .C1(n13527), .C2(n9710), .A(n13703), .B(n13523), .ZN(
        n13526) );
  NAND2_X1 U15580 ( .A1(n13524), .A2(n6779), .ZN(n13525) );
  OAI211_X1 U15581 ( .C1(n6466), .C2(n13527), .A(n13526), .B(n13525), .ZN(
        n13532) );
  NAND3_X1 U15582 ( .A1(n13527), .A2(n13703), .A3(n9710), .ZN(n13528) );
  OAI21_X1 U15583 ( .B1(n6466), .B2(n13529), .A(n13528), .ZN(n13531) );
  OAI22_X1 U15584 ( .A1(n13532), .A2(n13531), .B1(n6466), .B2(n13530), .ZN(
        n13534) );
  NAND2_X1 U15585 ( .A1(n13534), .A2(n13533), .ZN(n13542) );
  INV_X1 U15586 ( .A(n13535), .ZN(n13538) );
  INV_X1 U15587 ( .A(n13536), .ZN(n13537) );
  MUX2_X1 U15588 ( .A(n13538), .B(n13537), .S(n13703), .Z(n13540) );
  NOR2_X1 U15589 ( .A1(n13540), .A2(n13539), .ZN(n13541) );
  NAND2_X1 U15590 ( .A1(n13542), .A2(n13541), .ZN(n13546) );
  MUX2_X1 U15591 ( .A(n13544), .B(n13543), .S(n6591), .Z(n13545) );
  NAND2_X1 U15592 ( .A1(n13546), .A2(n13545), .ZN(n13551) );
  MUX2_X1 U15593 ( .A(n13548), .B(n13748), .S(n6591), .Z(n13547) );
  INV_X1 U15594 ( .A(n13547), .ZN(n13550) );
  MUX2_X1 U15595 ( .A(n13548), .B(n13748), .S(n6466), .Z(n13549) );
  OAI21_X1 U15596 ( .B1(n13551), .B2(n13550), .A(n13549), .ZN(n13553) );
  NAND2_X1 U15597 ( .A1(n13551), .A2(n13550), .ZN(n13552) );
  MUX2_X1 U15598 ( .A(n14713), .B(n13747), .S(n6466), .Z(n13555) );
  MUX2_X1 U15599 ( .A(n14713), .B(n13747), .S(n6591), .Z(n13554) );
  MUX2_X1 U15600 ( .A(n13556), .B(n13746), .S(n6591), .Z(n13559) );
  NAND2_X1 U15601 ( .A1(n13560), .A2(n13559), .ZN(n13558) );
  MUX2_X1 U15602 ( .A(n13556), .B(n13746), .S(n6466), .Z(n13557) );
  NAND2_X1 U15603 ( .A1(n13558), .A2(n13557), .ZN(n13562) );
  NAND2_X1 U15604 ( .A1(n13562), .A2(n13561), .ZN(n13566) );
  MUX2_X1 U15605 ( .A(n13745), .B(n13563), .S(n6591), .Z(n13567) );
  NAND2_X1 U15606 ( .A1(n13566), .A2(n13567), .ZN(n13565) );
  MUX2_X1 U15607 ( .A(n13563), .B(n13745), .S(n7235), .Z(n13564) );
  NAND2_X1 U15608 ( .A1(n13565), .A2(n13564), .ZN(n13571) );
  INV_X1 U15609 ( .A(n13566), .ZN(n13569) );
  INV_X1 U15610 ( .A(n13567), .ZN(n13568) );
  NAND2_X1 U15611 ( .A1(n13569), .A2(n13568), .ZN(n13570) );
  NAND2_X1 U15612 ( .A1(n13571), .A2(n13570), .ZN(n13575) );
  MUX2_X1 U15613 ( .A(n13744), .B(n13572), .S(n6466), .Z(n13574) );
  MUX2_X1 U15614 ( .A(n13744), .B(n13572), .S(n6591), .Z(n13573) );
  MUX2_X1 U15615 ( .A(n13743), .B(n13576), .S(n6591), .Z(n13580) );
  MUX2_X1 U15616 ( .A(n13743), .B(n13576), .S(n6466), .Z(n13577) );
  NAND2_X1 U15617 ( .A1(n13578), .A2(n13577), .ZN(n13584) );
  INV_X1 U15618 ( .A(n13579), .ZN(n13582) );
  INV_X1 U15619 ( .A(n13580), .ZN(n13581) );
  NAND2_X1 U15620 ( .A1(n13582), .A2(n13581), .ZN(n13583) );
  NAND2_X1 U15621 ( .A1(n13584), .A2(n13583), .ZN(n13587) );
  MUX2_X1 U15622 ( .A(n13742), .B(n14559), .S(n6466), .Z(n13588) );
  NAND2_X1 U15623 ( .A1(n13587), .A2(n13588), .ZN(n13586) );
  MUX2_X1 U15624 ( .A(n13742), .B(n14559), .S(n6591), .Z(n13585) );
  NAND2_X1 U15625 ( .A1(n13586), .A2(n13585), .ZN(n13592) );
  INV_X1 U15626 ( .A(n13587), .ZN(n13590) );
  INV_X1 U15627 ( .A(n13588), .ZN(n13589) );
  NAND2_X1 U15628 ( .A1(n13590), .A2(n13589), .ZN(n13591) );
  NAND2_X1 U15629 ( .A1(n13592), .A2(n13591), .ZN(n13595) );
  MUX2_X1 U15630 ( .A(n13741), .B(n14575), .S(n6591), .Z(n13596) );
  NAND2_X1 U15631 ( .A1(n13595), .A2(n13596), .ZN(n13594) );
  MUX2_X1 U15632 ( .A(n13741), .B(n14575), .S(n6466), .Z(n13593) );
  NAND2_X1 U15633 ( .A1(n13594), .A2(n13593), .ZN(n13600) );
  INV_X1 U15634 ( .A(n13595), .ZN(n13598) );
  INV_X1 U15635 ( .A(n13596), .ZN(n13597) );
  NAND2_X1 U15636 ( .A1(n13598), .A2(n13597), .ZN(n13599) );
  MUX2_X1 U15637 ( .A(n13740), .B(n13601), .S(n6466), .Z(n13603) );
  MUX2_X1 U15638 ( .A(n13740), .B(n13601), .S(n7235), .Z(n13602) );
  MUX2_X1 U15639 ( .A(n13739), .B(n13607), .S(n7235), .Z(n13615) );
  AND2_X1 U15640 ( .A1(n13616), .A2(n13604), .ZN(n13605) );
  AND4_X1 U15641 ( .A1(n13616), .A2(n6466), .A3(n13617), .A4(n13607), .ZN(
        n13608) );
  NAND2_X1 U15642 ( .A1(n13609), .A2(n13608), .ZN(n13622) );
  NOR2_X1 U15643 ( .A1(n13610), .A2(n14086), .ZN(n13613) );
  AOI21_X1 U15644 ( .B1(n13610), .B2(n14086), .A(n7235), .ZN(n13611) );
  OAI21_X1 U15645 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n13621) );
  INV_X1 U15646 ( .A(n13614), .ZN(n13619) );
  INV_X1 U15647 ( .A(n13615), .ZN(n13618) );
  NAND4_X1 U15648 ( .A1(n13619), .A2(n13618), .A3(n13617), .A4(n13616), .ZN(
        n13620) );
  NAND3_X1 U15649 ( .A1(n13622), .A2(n13621), .A3(n13620), .ZN(n13624) );
  OAI22_X1 U15650 ( .A1(n13625), .A2(n13624), .B1(n6466), .B2(n13623), .ZN(
        n13634) );
  MUX2_X1 U15651 ( .A(n13737), .B(n14188), .S(n7235), .Z(n13646) );
  AOI21_X1 U15652 ( .B1(n13646), .B2(n14084), .A(n6592), .ZN(n13632) );
  NAND2_X1 U15653 ( .A1(n14084), .A2(n6466), .ZN(n13647) );
  OR2_X1 U15654 ( .A1(n14188), .A2(n13647), .ZN(n13627) );
  NAND2_X1 U15655 ( .A1(n6592), .A2(n13628), .ZN(n13626) );
  AND2_X1 U15656 ( .A1(n13627), .A2(n13626), .ZN(n13636) );
  NAND2_X1 U15657 ( .A1(n13646), .A2(n13628), .ZN(n13629) );
  OR2_X1 U15658 ( .A1(n14188), .A2(n7235), .ZN(n13644) );
  NAND2_X1 U15659 ( .A1(n13629), .A2(n13644), .ZN(n13630) );
  NAND2_X1 U15660 ( .A1(n13630), .A2(n14181), .ZN(n13631) );
  OAI211_X1 U15661 ( .C1(n13632), .C2(n14181), .A(n13636), .B(n13631), .ZN(
        n13633) );
  NAND2_X1 U15662 ( .A1(n13646), .A2(n6592), .ZN(n13635) );
  OAI21_X1 U15663 ( .B1(n6466), .B2(n14084), .A(n13635), .ZN(n13639) );
  INV_X1 U15664 ( .A(n13636), .ZN(n13637) );
  AOI22_X1 U15665 ( .A1(n13639), .A2(n13638), .B1(n13646), .B2(n13637), .ZN(
        n13652) );
  XNOR2_X1 U15666 ( .A(n13736), .B(n7235), .ZN(n13656) );
  NOR2_X1 U15667 ( .A1(n14175), .A2(n6466), .ZN(n13640) );
  AOI21_X1 U15668 ( .B1(n13655), .B2(n13656), .A(n13640), .ZN(n13643) );
  NAND3_X1 U15669 ( .A1(n13655), .A2(n6466), .A3(n14175), .ZN(n13641) );
  OAI21_X1 U15670 ( .B1(n13643), .B2(n13642), .A(n13641), .ZN(n13651) );
  INV_X1 U15671 ( .A(n13644), .ZN(n13645) );
  NAND2_X1 U15672 ( .A1(n13646), .A2(n13645), .ZN(n13648) );
  NAND2_X1 U15673 ( .A1(n13648), .A2(n13647), .ZN(n13649) );
  NAND2_X1 U15674 ( .A1(n13649), .A2(n14181), .ZN(n13650) );
  NAND3_X1 U15675 ( .A1(n14175), .A2(n6466), .A3(n13656), .ZN(n13653) );
  NAND2_X1 U15676 ( .A1(n13655), .A2(n13653), .ZN(n13654) );
  OAI21_X1 U15677 ( .B1(n13655), .B2(n7235), .A(n13654), .ZN(n13658) );
  NAND4_X1 U15678 ( .A1(n13659), .A2(n14068), .A3(n7235), .A4(n13656), .ZN(
        n13657) );
  OAI211_X1 U15679 ( .C1(n13659), .C2(n7235), .A(n13658), .B(n13657), .ZN(
        n13660) );
  INV_X1 U15680 ( .A(n13660), .ZN(n13661) );
  MUX2_X1 U15681 ( .A(n13734), .B(n14157), .S(n6466), .Z(n13663) );
  MUX2_X1 U15682 ( .A(n13733), .B(n14010), .S(n6466), .Z(n13667) );
  MUX2_X1 U15683 ( .A(n13733), .B(n14010), .S(n7235), .Z(n13665) );
  NAND2_X1 U15684 ( .A1(n13666), .A2(n13665), .ZN(n13669) );
  MUX2_X1 U15685 ( .A(n13982), .B(n13997), .S(n6466), .Z(n13670) );
  MUX2_X1 U15686 ( .A(n13732), .B(n13978), .S(n6466), .Z(n13676) );
  MUX2_X1 U15687 ( .A(n13732), .B(n13978), .S(n7235), .Z(n13675) );
  MUX2_X1 U15688 ( .A(n13983), .B(n13961), .S(n7235), .Z(n13679) );
  NAND2_X1 U15689 ( .A1(n13680), .A2(n13679), .ZN(n13678) );
  MUX2_X1 U15690 ( .A(n13983), .B(n13961), .S(n6466), .Z(n13677) );
  NAND2_X1 U15691 ( .A1(n13678), .A2(n13677), .ZN(n13682) );
  NAND2_X1 U15692 ( .A1(n13682), .A2(n13681), .ZN(n13685) );
  MUX2_X1 U15693 ( .A(n13731), .B(n13943), .S(n6466), .Z(n13686) );
  NAND2_X1 U15694 ( .A1(n13685), .A2(n13686), .ZN(n13684) );
  MUX2_X1 U15695 ( .A(n13731), .B(n13943), .S(n7235), .Z(n13683) );
  NAND2_X1 U15696 ( .A1(n13684), .A2(n13683), .ZN(n13690) );
  INV_X1 U15697 ( .A(n13685), .ZN(n13688) );
  INV_X1 U15698 ( .A(n13686), .ZN(n13687) );
  NAND2_X1 U15699 ( .A1(n13688), .A2(n13687), .ZN(n13689) );
  NAND2_X1 U15700 ( .A1(n13690), .A2(n13689), .ZN(n13693) );
  MUX2_X1 U15701 ( .A(n13934), .B(n13928), .S(n7235), .Z(n13692) );
  MUX2_X1 U15702 ( .A(n13934), .B(n13928), .S(n6466), .Z(n13691) );
  MUX2_X1 U15703 ( .A(n13903), .B(n14115), .S(n6466), .Z(n13696) );
  MUX2_X1 U15704 ( .A(n13903), .B(n14115), .S(n7235), .Z(n13694) );
  NAND2_X1 U15705 ( .A1(n13695), .A2(n13694), .ZN(n13699) );
  INV_X1 U15706 ( .A(n13696), .ZN(n13697) );
  MUX2_X1 U15707 ( .A(n13888), .B(n14111), .S(n7235), .Z(n13701) );
  MUX2_X1 U15708 ( .A(n13888), .B(n14111), .S(n6466), .Z(n13700) );
  INV_X1 U15709 ( .A(n13701), .ZN(n13702) );
  MUX2_X1 U15710 ( .A(n13902), .B(n13883), .S(n6466), .Z(n13707) );
  NAND2_X1 U15711 ( .A1(n13706), .A2(n13707), .ZN(n13705) );
  MUX2_X1 U15712 ( .A(n13902), .B(n13883), .S(n6591), .Z(n13704) );
  INV_X1 U15713 ( .A(n13706), .ZN(n13709) );
  INV_X1 U15714 ( .A(n13707), .ZN(n13708) );
  INV_X1 U15715 ( .A(n13710), .ZN(n13712) );
  NAND2_X1 U15716 ( .A1(n13724), .A2(n13711), .ZN(n13714) );
  AOI211_X1 U15717 ( .C1(n13713), .C2(n13712), .A(n13717), .B(n13714), .ZN(
        n13723) );
  NOR4_X1 U15718 ( .A1(n13716), .A2(n14020), .A3(n14619), .A4(n13715), .ZN(
        n13719) );
  OAI21_X1 U15719 ( .B1(n14254), .B2(n13717), .A(P1_B_REG_SCAN_IN), .ZN(n13718) );
  OAI22_X1 U15720 ( .A1(n13721), .A2(n13720), .B1(n13719), .B2(n13718), .ZN(
        n13722) );
  INV_X1 U15721 ( .A(n13724), .ZN(n13729) );
  INV_X1 U15722 ( .A(n13725), .ZN(n13728) );
  MUX2_X1 U15723 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n13884), .S(n13750), .Z(
        P1_U3590) );
  MUX2_X1 U15724 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13902), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15725 ( .A(n13888), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13751), .Z(
        P1_U3588) );
  MUX2_X1 U15726 ( .A(n13903), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13751), .Z(
        P1_U3587) );
  MUX2_X1 U15727 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n13934), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U15728 ( .A(n13731), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13751), .Z(
        P1_U3585) );
  MUX2_X1 U15729 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n13983), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U15730 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n13732), .S(n13750), .Z(
        P1_U3583) );
  MUX2_X1 U15731 ( .A(n13982), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13751), .Z(
        P1_U3582) );
  MUX2_X1 U15732 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n13733), .S(P1_U4016), .Z(
        P1_U3581) );
  MUX2_X1 U15733 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13734), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15734 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13735), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15735 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n13736), .S(P1_U4016), .Z(
        P1_U3578) );
  MUX2_X1 U15736 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14084), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U15737 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n13737), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U15738 ( .A(n14086), .B(P1_DATAO_REG_15__SCAN_IN), .S(n13751), .Z(
        P1_U3575) );
  MUX2_X1 U15739 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n13738), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U15740 ( .A(n13739), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13751), .Z(
        P1_U3573) );
  MUX2_X1 U15741 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n13740), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U15742 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n13741), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U15743 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n13742), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U15744 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n13743), .S(P1_U4016), .Z(
        P1_U3569) );
  MUX2_X1 U15745 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n13744), .S(n13750), .Z(
        P1_U3568) );
  MUX2_X1 U15746 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n13745), .S(n13750), .Z(
        P1_U3567) );
  MUX2_X1 U15747 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n13746), .S(n13750), .Z(
        P1_U3566) );
  MUX2_X1 U15748 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n13747), .S(P1_U4016), .Z(
        P1_U3565) );
  MUX2_X1 U15749 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n13748), .S(n13750), .Z(
        P1_U3564) );
  MUX2_X1 U15750 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n13749), .S(n13750), .Z(
        P1_U3562) );
  MUX2_X1 U15751 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9710), .S(n13750), .Z(
        P1_U3561) );
  MUX2_X1 U15752 ( .A(n13752), .B(P1_DATAO_REG_0__SCAN_IN), .S(n13751), .Z(
        P1_U3560) );
  INV_X1 U15753 ( .A(n13753), .ZN(n13758) );
  MUX2_X1 U15754 ( .A(n9307), .B(P1_REG2_REG_1__SCAN_IN), .S(n13754), .Z(
        n13757) );
  INV_X1 U15755 ( .A(n13755), .ZN(n13756) );
  OAI211_X1 U15756 ( .C1(n13758), .C2(n13757), .A(n14641), .B(n13756), .ZN(
        n13765) );
  AOI22_X1 U15757 ( .A1(n14627), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13764) );
  NAND2_X1 U15758 ( .A1(n14637), .A2(n7362), .ZN(n13763) );
  AND2_X1 U15759 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n13760) );
  OAI211_X1 U15760 ( .C1(n13761), .C2(n13760), .A(n14640), .B(n13759), .ZN(
        n13762) );
  NAND4_X1 U15761 ( .A1(n13765), .A2(n13764), .A3(n13763), .A4(n13762), .ZN(
        P1_U3244) );
  OAI22_X1 U15762 ( .A1(n14645), .A2(n14259), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9684), .ZN(n13766) );
  AOI21_X1 U15763 ( .B1(n13767), .B2(n14637), .A(n13766), .ZN(n13776) );
  NAND2_X1 U15764 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  NAND3_X1 U15765 ( .A1(n14641), .A2(n13787), .A3(n13770), .ZN(n13775) );
  OAI211_X1 U15766 ( .C1(n13773), .C2(n13772), .A(n14640), .B(n13771), .ZN(
        n13774) );
  NAND4_X1 U15767 ( .A1(n13777), .A2(n13776), .A3(n13775), .A4(n13774), .ZN(
        P1_U3245) );
  AND2_X1 U15768 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13780) );
  NOR2_X1 U15769 ( .A1(n13807), .A2(n13778), .ZN(n13779) );
  AOI211_X1 U15770 ( .C1(n14627), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n13780), .B(
        n13779), .ZN(n13792) );
  OAI211_X1 U15771 ( .C1(n13783), .C2(n13782), .A(n14640), .B(n13781), .ZN(
        n13791) );
  INV_X1 U15772 ( .A(n13784), .ZN(n13789) );
  NAND3_X1 U15773 ( .A1(n13787), .A2(n13786), .A3(n13785), .ZN(n13788) );
  NAND3_X1 U15774 ( .A1(n14641), .A2(n13789), .A3(n13788), .ZN(n13790) );
  NAND3_X1 U15775 ( .A1(n13792), .A2(n13791), .A3(n13790), .ZN(P1_U3246) );
  AOI211_X1 U15776 ( .C1(n13795), .C2(n13794), .A(n13793), .B(n13819), .ZN(
        n13796) );
  INV_X1 U15777 ( .A(n13796), .ZN(n13806) );
  INV_X1 U15778 ( .A(n13797), .ZN(n13798) );
  AOI21_X1 U15779 ( .B1(n14627), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n13798), 
        .ZN(n13805) );
  OAI211_X1 U15780 ( .C1(n13801), .C2(n13800), .A(n14641), .B(n13799), .ZN(
        n13804) );
  NAND2_X1 U15781 ( .A1(n14637), .A2(n13802), .ZN(n13803) );
  NAND4_X1 U15782 ( .A1(n13806), .A2(n13805), .A3(n13804), .A4(n13803), .ZN(
        P1_U3256) );
  NOR2_X1 U15783 ( .A1(n13807), .A2(n13830), .ZN(n13808) );
  AOI211_X1 U15784 ( .C1(n14627), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n13809), 
        .B(n13808), .ZN(n13825) );
  NOR2_X1 U15785 ( .A1(n13830), .A2(n13810), .ZN(n13811) );
  AOI21_X1 U15786 ( .B1(n13810), .B2(n13830), .A(n13811), .ZN(n13816) );
  INV_X1 U15787 ( .A(n13818), .ZN(n13814) );
  INV_X1 U15788 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n13813) );
  OAI21_X1 U15789 ( .B1(n13814), .B2(n13813), .A(n13812), .ZN(n13815) );
  NAND2_X1 U15790 ( .A1(n13816), .A2(n13815), .ZN(n13829) );
  OAI211_X1 U15791 ( .C1(n13816), .C2(n13815), .A(n14641), .B(n13829), .ZN(
        n13824) );
  XNOR2_X1 U15792 ( .A(n13833), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n13820) );
  NOR2_X1 U15793 ( .A1(n13821), .A2(n13820), .ZN(n13832) );
  AOI211_X1 U15794 ( .C1(n13821), .C2(n13820), .A(n13832), .B(n13819), .ZN(
        n13822) );
  INV_X1 U15795 ( .A(n13822), .ZN(n13823) );
  NAND3_X1 U15796 ( .A1(n13825), .A2(n13824), .A3(n13823), .ZN(P1_U3260) );
  INV_X1 U15797 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n13827) );
  OAI21_X1 U15798 ( .B1(n14645), .B2(n13827), .A(n13826), .ZN(n13828) );
  AOI21_X1 U15799 ( .B1(n13847), .B2(n14637), .A(n13828), .ZN(n13840) );
  OAI21_X1 U15800 ( .B1(n13810), .B2(n13830), .A(n13829), .ZN(n13846) );
  XNOR2_X1 U15801 ( .A(n13841), .B(n13846), .ZN(n13831) );
  NAND2_X1 U15802 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n13831), .ZN(n13849) );
  OAI211_X1 U15803 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n13831), .A(n14641), 
        .B(n13849), .ZN(n13839) );
  XNOR2_X1 U15804 ( .A(n13841), .B(n13842), .ZN(n13834) );
  INV_X1 U15805 ( .A(n13834), .ZN(n13837) );
  NOR2_X1 U15806 ( .A1(n13835), .A2(n13834), .ZN(n13844) );
  INV_X1 U15807 ( .A(n13844), .ZN(n13836) );
  OAI211_X1 U15808 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n13837), .A(n14640), 
        .B(n13836), .ZN(n13838) );
  NAND3_X1 U15809 ( .A1(n13840), .A2(n13839), .A3(n13838), .ZN(P1_U3261) );
  NOR2_X1 U15810 ( .A1(n13842), .A2(n13841), .ZN(n13843) );
  NOR2_X1 U15811 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  XNOR2_X1 U15812 ( .A(n13845), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n13855) );
  INV_X1 U15813 ( .A(n13855), .ZN(n13853) );
  NAND2_X1 U15814 ( .A1(n13847), .A2(n13846), .ZN(n13848) );
  NAND2_X1 U15815 ( .A1(n13849), .A2(n13848), .ZN(n13850) );
  XOR2_X1 U15816 ( .A(n13850), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13854) );
  NOR2_X1 U15817 ( .A1(n13854), .A2(n13851), .ZN(n13852) );
  AOI22_X1 U15818 ( .A1(n13855), .A2(n14640), .B1(n14641), .B2(n13854), .ZN(
        n13856) );
  INV_X1 U15819 ( .A(n13857), .ZN(n13858) );
  OAI211_X1 U15820 ( .C1(n7474), .C2(n14645), .A(n13859), .B(n13858), .ZN(
        P1_U3262) );
  NAND2_X1 U15821 ( .A1(n14206), .A2(n13882), .ZN(n13869) );
  XNOR2_X1 U15822 ( .A(n13862), .B(n13869), .ZN(n13863) );
  NAND2_X1 U15823 ( .A1(n14093), .A2(n14659), .ZN(n13868) );
  NOR2_X1 U15824 ( .A1(n14619), .A2(n13864), .ZN(n13865) );
  NOR2_X1 U15825 ( .A1(n14060), .A2(n13865), .ZN(n13885) );
  AND2_X1 U15826 ( .A1(n13866), .A2(n13885), .ZN(n14092) );
  INV_X1 U15827 ( .A(n14092), .ZN(n14096) );
  NOR2_X1 U15828 ( .A1(n14650), .A2(n14096), .ZN(n13871) );
  AOI21_X1 U15829 ( .B1(n14673), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13871), 
        .ZN(n13867) );
  OAI211_X1 U15830 ( .C1(n7236), .C2(n14666), .A(n13868), .B(n13867), .ZN(
        P1_U3263) );
  OAI211_X1 U15831 ( .C1(n14206), .C2(n13882), .A(n14163), .B(n13869), .ZN(
        n14097) );
  NOR2_X1 U15832 ( .A1(n14206), .A2(n14666), .ZN(n13870) );
  AOI211_X1 U15833 ( .C1(n14650), .C2(P1_REG2_REG_30__SCAN_IN), .A(n13871), 
        .B(n13870), .ZN(n13872) );
  OAI21_X1 U15834 ( .B1(n13975), .B2(n14097), .A(n13872), .ZN(P1_U3264) );
  NAND2_X1 U15835 ( .A1(n14107), .A2(n13874), .ZN(n13875) );
  NAND2_X1 U15836 ( .A1(n13860), .A2(n13888), .ZN(n13879) );
  INV_X1 U15837 ( .A(n13883), .ZN(n14102) );
  AOI211_X1 U15838 ( .C1(n13883), .C2(n13900), .A(n14075), .B(n13882), .ZN(
        n14104) );
  NAND2_X1 U15839 ( .A1(n14104), .A2(n14659), .ZN(n13892) );
  NAND2_X1 U15840 ( .A1(n13885), .A2(n13884), .ZN(n14100) );
  OAI22_X1 U15841 ( .A1(n13887), .A2(n14100), .B1(n13886), .B2(n14044), .ZN(
        n13890) );
  NAND2_X1 U15842 ( .A1(n13888), .A2(n14085), .ZN(n14101) );
  NOR2_X1 U15843 ( .A1(n14673), .A2(n14101), .ZN(n13889) );
  AOI211_X1 U15844 ( .C1(n14673), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13890), 
        .B(n13889), .ZN(n13891) );
  OAI211_X1 U15845 ( .C1(n14102), .C2(n14666), .A(n13892), .B(n13891), .ZN(
        n13893) );
  AOI21_X1 U15846 ( .B1(n14105), .B2(n13896), .A(n13893), .ZN(n13894) );
  OAI21_X1 U15847 ( .B1(n14106), .B2(n14091), .A(n13894), .ZN(P1_U3356) );
  XNOR2_X1 U15848 ( .A(n13895), .B(n13897), .ZN(n14114) );
  INV_X1 U15849 ( .A(n13896), .ZN(n14054) );
  NAND3_X1 U15850 ( .A1(n14108), .A2(n14107), .A3(n14655), .ZN(n13912) );
  AOI21_X1 U15851 ( .B1(n14111), .B2(n13899), .A(n14075), .ZN(n13901) );
  NAND2_X1 U15852 ( .A1(n13902), .A2(n14083), .ZN(n13905) );
  NAND2_X1 U15853 ( .A1(n13903), .A2(n14085), .ZN(n13904) );
  NAND2_X1 U15854 ( .A1(n13905), .A2(n13904), .ZN(n14110) );
  INV_X1 U15855 ( .A(n14110), .ZN(n13907) );
  OAI22_X1 U15856 ( .A1(n14673), .A2(n13907), .B1(n13906), .B2(n14044), .ZN(
        n13908) );
  AOI21_X1 U15857 ( .B1(P1_REG2_REG_28__SCAN_IN), .B2(n14650), .A(n13908), 
        .ZN(n13909) );
  OAI21_X1 U15858 ( .B1(n13860), .B2(n14666), .A(n13909), .ZN(n13910) );
  AOI21_X1 U15859 ( .B1(n14109), .B2(n14659), .A(n13910), .ZN(n13911) );
  OAI211_X1 U15860 ( .C1(n14114), .C2(n14054), .A(n13912), .B(n13911), .ZN(
        P1_U3265) );
  XNOR2_X1 U15861 ( .A(n13928), .B(n13936), .ZN(n13914) );
  OAI222_X1 U15862 ( .A1(n14075), .A2(n13914), .B1(n14060), .B2(n13913), .C1(
        n14020), .C2(n13953), .ZN(n14123) );
  OAI21_X1 U15863 ( .B1(n13917), .B2(n13916), .A(n13915), .ZN(n13918) );
  NAND2_X1 U15864 ( .A1(n13918), .A2(n14183), .ZN(n14124) );
  INV_X1 U15865 ( .A(n14124), .ZN(n13919) );
  AOI21_X1 U15866 ( .B1(n13920), .B2(n14123), .A(n13919), .ZN(n13930) );
  OAI22_X1 U15867 ( .A1(n14047), .A2(n13922), .B1(n13921), .B2(n14044), .ZN(
        n13927) );
  OAI21_X1 U15868 ( .B1(n13925), .B2(n13924), .A(n13923), .ZN(n14126) );
  NOR2_X1 U15869 ( .A1(n14126), .A2(n14091), .ZN(n13926) );
  AOI211_X1 U15870 ( .C1(n13994), .C2(n13928), .A(n13927), .B(n13926), .ZN(
        n13929) );
  OAI21_X1 U15871 ( .B1(n14673), .B2(n13930), .A(n13929), .ZN(P1_U3267) );
  OAI21_X1 U15872 ( .B1(n13933), .B2(n13932), .A(n13931), .ZN(n13935) );
  AOI222_X1 U15873 ( .A1(n14183), .A2(n13935), .B1(n13983), .B2(n14085), .C1(
        n13934), .C2(n14083), .ZN(n14133) );
  AOI21_X1 U15874 ( .B1(n13943), .B2(n13959), .A(n14075), .ZN(n13937) );
  NAND2_X1 U15875 ( .A1(n13937), .A2(n13936), .ZN(n14130) );
  OR2_X1 U15876 ( .A1(n13939), .A2(n13938), .ZN(n14129) );
  NAND3_X1 U15877 ( .A1(n14129), .A2(n14128), .A3(n14655), .ZN(n13945) );
  NAND2_X1 U15878 ( .A1(n14673), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13940) );
  OAI21_X1 U15879 ( .B1(n14044), .B2(n13941), .A(n13940), .ZN(n13942) );
  AOI21_X1 U15880 ( .B1(n13943), .B2(n13994), .A(n13942), .ZN(n13944) );
  OAI211_X1 U15881 ( .C1(n14130), .C2(n13975), .A(n13945), .B(n13944), .ZN(
        n13946) );
  INV_X1 U15882 ( .A(n13946), .ZN(n13947) );
  OAI21_X1 U15883 ( .B1(n14133), .B2(n14673), .A(n13947), .ZN(P1_U3268) );
  AOI21_X1 U15884 ( .B1(n13949), .B2(n13948), .A(n6423), .ZN(n14134) );
  AOI211_X1 U15885 ( .C1(n13952), .C2(n13951), .A(n14166), .B(n13950), .ZN(
        n13955) );
  OAI22_X1 U15886 ( .A1(n13953), .A2(n14060), .B1(n13990), .B2(n14020), .ZN(
        n13954) );
  NOR2_X1 U15887 ( .A1(n13955), .A2(n13954), .ZN(n13956) );
  OAI21_X1 U15888 ( .B1(n14134), .B2(n13957), .A(n13956), .ZN(n14135) );
  NAND2_X1 U15889 ( .A1(n14135), .A2(n14047), .ZN(n13967) );
  INV_X1 U15890 ( .A(n13959), .ZN(n13960) );
  AOI211_X1 U15891 ( .C1(n13961), .C2(n13974), .A(n14075), .B(n13960), .ZN(
        n14136) );
  NOR2_X1 U15892 ( .A1(n11616), .A2(n14666), .ZN(n13965) );
  OAI22_X1 U15893 ( .A1(n14047), .A2(n13963), .B1(n13962), .B2(n14044), .ZN(
        n13964) );
  AOI211_X1 U15894 ( .C1(n14136), .C2(n14659), .A(n13965), .B(n13964), .ZN(
        n13966) );
  OAI211_X1 U15895 ( .C1(n14134), .C2(n14072), .A(n13967), .B(n13966), .ZN(
        P1_U3269) );
  NAND2_X1 U15896 ( .A1(n13968), .A2(n7434), .ZN(n13969) );
  NAND2_X1 U15897 ( .A1(n13970), .A2(n13969), .ZN(n14140) );
  INV_X1 U15898 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n13972) );
  OAI22_X1 U15899 ( .A1(n14047), .A2(n13972), .B1(n13971), .B2(n14044), .ZN(
        n13977) );
  NAND2_X1 U15900 ( .A1(n13978), .A2(n13998), .ZN(n13973) );
  NAND3_X1 U15901 ( .A1(n13974), .A2(n14163), .A3(n13973), .ZN(n14141) );
  NOR2_X1 U15902 ( .A1(n14141), .A2(n13975), .ZN(n13976) );
  AOI211_X1 U15903 ( .C1(n13994), .C2(n13978), .A(n13977), .B(n13976), .ZN(
        n13987) );
  OAI21_X1 U15904 ( .B1(n13980), .B2(n7434), .A(n13979), .ZN(n13981) );
  NAND2_X1 U15905 ( .A1(n13981), .A2(n14183), .ZN(n13985) );
  AOI22_X1 U15906 ( .A1(n14083), .A2(n13983), .B1(n13982), .B2(n14085), .ZN(
        n13984) );
  NAND2_X1 U15907 ( .A1(n13985), .A2(n13984), .ZN(n14144) );
  NAND2_X1 U15908 ( .A1(n14144), .A2(n14047), .ZN(n13986) );
  OAI211_X1 U15909 ( .C1(n14140), .C2(n14091), .A(n13987), .B(n13986), .ZN(
        P1_U3270) );
  XOR2_X1 U15910 ( .A(n13988), .B(n13996), .Z(n13989) );
  OAI222_X1 U15911 ( .A1(n14020), .A2(n14021), .B1(n14060), .B2(n13990), .C1(
        n14166), .C2(n13989), .ZN(n14146) );
  NAND2_X1 U15912 ( .A1(n14146), .A2(n14047), .ZN(n14003) );
  NAND2_X1 U15913 ( .A1(n14650), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n13991) );
  OAI21_X1 U15914 ( .B1(n14044), .B2(n13992), .A(n13991), .ZN(n13993) );
  AOI21_X1 U15915 ( .B1(n13997), .B2(n13994), .A(n13993), .ZN(n14002) );
  XNOR2_X1 U15916 ( .A(n13995), .B(n13996), .ZN(n14148) );
  NAND2_X1 U15917 ( .A1(n14148), .A2(n14655), .ZN(n14001) );
  AOI21_X1 U15918 ( .B1(n13997), .B2(n14012), .A(n14075), .ZN(n13999) );
  AND2_X1 U15919 ( .A1(n13999), .A2(n13998), .ZN(n14147) );
  NAND2_X1 U15920 ( .A1(n14147), .A2(n14659), .ZN(n14000) );
  NAND4_X1 U15921 ( .A1(n14003), .A2(n14002), .A3(n14001), .A4(n14000), .ZN(
        P1_U3271) );
  XNOR2_X1 U15922 ( .A(n14004), .B(n14008), .ZN(n14007) );
  INV_X1 U15923 ( .A(n14005), .ZN(n14006) );
  OAI21_X1 U15924 ( .B1(n14007), .B2(n14166), .A(n14006), .ZN(n14151) );
  INV_X1 U15925 ( .A(n14151), .ZN(n14018) );
  OAI21_X1 U15926 ( .B1(n6528), .B2(n7423), .A(n14009), .ZN(n14153) );
  INV_X1 U15927 ( .A(n14010), .ZN(n14222) );
  NAND2_X1 U15928 ( .A1(n14010), .A2(n14025), .ZN(n14011) );
  AND3_X1 U15929 ( .A1(n14012), .A2(n14163), .A3(n14011), .ZN(n14152) );
  NAND2_X1 U15930 ( .A1(n14152), .A2(n14659), .ZN(n14015) );
  AOI22_X1 U15931 ( .A1(n14013), .A2(n14662), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n14650), .ZN(n14014) );
  OAI211_X1 U15932 ( .C1(n14222), .C2(n14666), .A(n14015), .B(n14014), .ZN(
        n14016) );
  AOI21_X1 U15933 ( .B1(n14153), .B2(n14655), .A(n14016), .ZN(n14017) );
  OAI21_X1 U15934 ( .B1(n14650), .B2(n14018), .A(n14017), .ZN(P1_U3272) );
  AOI21_X1 U15935 ( .B1(n11537), .B2(n14019), .A(n14166), .ZN(n14024) );
  OAI22_X1 U15936 ( .A1(n14021), .A2(n14060), .B1(n14061), .B2(n14020), .ZN(
        n14022) );
  AOI21_X1 U15937 ( .B1(n14024), .B2(n14023), .A(n14022), .ZN(n14161) );
  OAI211_X1 U15938 ( .C1(n14028), .C2(n14042), .A(n14163), .B(n14025), .ZN(
        n14158) );
  INV_X1 U15939 ( .A(n14158), .ZN(n14030) );
  AOI22_X1 U15940 ( .A1(n14026), .A2(n14662), .B1(n14673), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n14027) );
  OAI21_X1 U15941 ( .B1(n14028), .B2(n14666), .A(n14027), .ZN(n14029) );
  AOI21_X1 U15942 ( .B1(n14030), .B2(n14659), .A(n14029), .ZN(n14035) );
  NAND2_X1 U15943 ( .A1(n14032), .A2(n14033), .ZN(n14156) );
  NAND3_X1 U15944 ( .A1(n14031), .A2(n14156), .A3(n14655), .ZN(n14034) );
  OAI211_X1 U15945 ( .C1(n14161), .C2(n14650), .A(n14035), .B(n14034), .ZN(
        P1_U3273) );
  OAI21_X1 U15946 ( .B1(n14038), .B2(n14037), .A(n14036), .ZN(n14039) );
  INV_X1 U15947 ( .A(n14039), .ZN(n14167) );
  XNOR2_X1 U15948 ( .A(n14041), .B(n14040), .ZN(n14169) );
  NAND2_X1 U15949 ( .A1(n14169), .A2(n14655), .ZN(n14053) );
  AOI21_X1 U15950 ( .B1(n14043), .B2(n14063), .A(n14042), .ZN(n14164) );
  OAI22_X1 U15951 ( .A1(n14047), .A2(n14046), .B1(n14045), .B2(n14044), .ZN(
        n14048) );
  AOI21_X1 U15952 ( .B1(n14162), .B2(n14047), .A(n14048), .ZN(n14049) );
  OAI21_X1 U15953 ( .B1(n14228), .B2(n14666), .A(n14049), .ZN(n14050) );
  AOI21_X1 U15954 ( .B1(n14164), .B2(n14051), .A(n14050), .ZN(n14052) );
  OAI211_X1 U15955 ( .C1(n14167), .C2(n14054), .A(n14053), .B(n14052), .ZN(
        P1_U3274) );
  XNOR2_X1 U15956 ( .A(n14055), .B(n14056), .ZN(n14058) );
  INV_X1 U15957 ( .A(n14058), .ZN(n14178) );
  XOR2_X1 U15958 ( .A(n14057), .B(n14056), .Z(n14059) );
  AOI222_X1 U15959 ( .A1(n14183), .A2(n14059), .B1(n14058), .B2(n6436), .C1(
        n14084), .C2(n14085), .ZN(n14177) );
  INV_X1 U15960 ( .A(n14177), .ZN(n14062) );
  NOR2_X1 U15961 ( .A1(n14061), .A2(n14060), .ZN(n14174) );
  OAI21_X1 U15962 ( .B1(n14062), .B2(n14174), .A(n14047), .ZN(n14071) );
  INV_X1 U15963 ( .A(n14063), .ZN(n14064) );
  AOI211_X1 U15964 ( .C1(n14175), .C2(n14065), .A(n14075), .B(n14064), .ZN(
        n14173) );
  AOI22_X1 U15965 ( .A1(n14650), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n14066), 
        .B2(n14662), .ZN(n14067) );
  OAI21_X1 U15966 ( .B1(n14068), .B2(n14666), .A(n14067), .ZN(n14069) );
  AOI21_X1 U15967 ( .B1(n14173), .B2(n14659), .A(n14069), .ZN(n14070) );
  OAI211_X1 U15968 ( .C1(n14178), .C2(n14072), .A(n14071), .B(n14070), .ZN(
        P1_U3275) );
  XNOR2_X1 U15969 ( .A(n14073), .B(n14081), .ZN(n14191) );
  AOI211_X1 U15970 ( .C1(n14188), .C2(n14076), .A(n14075), .B(n14074), .ZN(
        n14187) );
  INV_X1 U15971 ( .A(n14077), .ZN(n14078) );
  AOI22_X1 U15972 ( .A1(n14673), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n14078), 
        .B2(n14662), .ZN(n14079) );
  OAI21_X1 U15973 ( .B1(n6938), .B2(n14666), .A(n14079), .ZN(n14089) );
  OAI21_X1 U15974 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(n14087) );
  AOI222_X1 U15975 ( .A1(n14183), .A2(n14087), .B1(n14086), .B2(n14085), .C1(
        n14084), .C2(n14083), .ZN(n14190) );
  NOR2_X1 U15976 ( .A1(n14190), .A2(n14650), .ZN(n14088) );
  AOI211_X1 U15977 ( .C1(n14187), .C2(n14659), .A(n14089), .B(n14088), .ZN(
        n14090) );
  OAI21_X1 U15978 ( .B1(n14091), .B2(n14191), .A(n14090), .ZN(P1_U3277) );
  NOR2_X1 U15979 ( .A1(n14093), .A2(n14092), .ZN(n14200) );
  MUX2_X1 U15980 ( .A(n14094), .B(n14200), .S(n14734), .Z(n14095) );
  OAI21_X1 U15981 ( .B1(n7236), .B2(n14172), .A(n14095), .ZN(P1_U3559) );
  INV_X1 U15982 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14098) );
  AND2_X1 U15983 ( .A1(n14097), .A2(n14096), .ZN(n14203) );
  MUX2_X1 U15984 ( .A(n14098), .B(n14203), .S(n14734), .Z(n14099) );
  OAI21_X1 U15985 ( .B1(n14206), .B2(n14172), .A(n14099), .ZN(P1_U3558) );
  OAI211_X1 U15986 ( .C1(n14102), .C2(n14587), .A(n14101), .B(n14100), .ZN(
        n14103) );
  NAND3_X1 U15987 ( .A1(n14108), .A2(n14107), .A3(n14725), .ZN(n14113) );
  AOI211_X1 U15988 ( .C1(n14111), .C2(n14712), .A(n14110), .B(n14109), .ZN(
        n14112) );
  OAI211_X1 U15989 ( .C1(n14166), .C2(n14114), .A(n14113), .B(n14112), .ZN(
        n14208) );
  MUX2_X1 U15990 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14208), .S(n14734), .Z(
        P1_U3556) );
  AOI22_X1 U15991 ( .A1(n14116), .A2(n14163), .B1(n14115), .B2(n14712), .ZN(
        n14117) );
  MUX2_X1 U15992 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14209), .S(n14734), .Z(
        P1_U3555) );
  NOR2_X1 U15993 ( .A1(n14123), .A2(n14122), .ZN(n14125) );
  OAI211_X1 U15994 ( .C1(n14126), .C2(n14192), .A(n14125), .B(n14124), .ZN(
        n14210) );
  MUX2_X1 U15995 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14210), .S(n14734), .Z(
        P1_U3554) );
  INV_X1 U15996 ( .A(n14127), .ZN(n14132) );
  NAND3_X1 U15997 ( .A1(n14129), .A2(n14128), .A3(n14725), .ZN(n14131) );
  NAND4_X1 U15998 ( .A1(n14133), .A2(n14132), .A3(n14131), .A4(n14130), .ZN(
        n14211) );
  MUX2_X1 U15999 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14211), .S(n14734), .Z(
        P1_U3553) );
  INV_X1 U16000 ( .A(n14134), .ZN(n14137) );
  AOI211_X1 U16001 ( .C1(n14385), .C2(n14137), .A(n14136), .B(n14135), .ZN(
        n14212) );
  MUX2_X1 U16002 ( .A(n14138), .B(n14212), .S(n14734), .Z(n14139) );
  OAI21_X1 U16003 ( .B1(n11616), .B2(n14172), .A(n14139), .ZN(P1_U3552) );
  NOR2_X1 U16004 ( .A1(n14140), .A2(n14192), .ZN(n14145) );
  OAI21_X1 U16005 ( .B1(n14142), .B2(n14587), .A(n14141), .ZN(n14143) );
  MUX2_X1 U16006 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14215), .S(n14734), .Z(
        P1_U3551) );
  AOI211_X1 U16007 ( .C1(n14725), .C2(n14148), .A(n14147), .B(n14146), .ZN(
        n14216) );
  MUX2_X1 U16008 ( .A(n14149), .B(n14216), .S(n14734), .Z(n14150) );
  OAI21_X1 U16009 ( .B1(n14172), .B2(n7363), .A(n14150), .ZN(P1_U3550) );
  INV_X1 U16010 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n14154) );
  AOI211_X1 U16011 ( .C1(n14725), .C2(n14153), .A(n14152), .B(n14151), .ZN(
        n14219) );
  MUX2_X1 U16012 ( .A(n14154), .B(n14219), .S(n14734), .Z(n14155) );
  OAI21_X1 U16013 ( .B1(n14222), .B2(n14172), .A(n14155), .ZN(P1_U3549) );
  NAND3_X1 U16014 ( .A1(n14031), .A2(n14156), .A3(n14725), .ZN(n14160) );
  NAND2_X1 U16015 ( .A1(n14157), .A2(n14712), .ZN(n14159) );
  NAND4_X1 U16016 ( .A1(n14161), .A2(n14160), .A3(n14159), .A4(n14158), .ZN(
        n14223) );
  MUX2_X1 U16017 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14223), .S(n14734), .Z(
        P1_U3548) );
  INV_X1 U16018 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14170) );
  AOI21_X1 U16019 ( .B1(n14164), .B2(n14163), .A(n14162), .ZN(n14165) );
  OAI21_X1 U16020 ( .B1(n14167), .B2(n14166), .A(n14165), .ZN(n14168) );
  AOI21_X1 U16021 ( .B1(n14725), .B2(n14169), .A(n14168), .ZN(n14224) );
  MUX2_X1 U16022 ( .A(n14170), .B(n14224), .S(n14734), .Z(n14171) );
  OAI21_X1 U16023 ( .B1(n14228), .B2(n14172), .A(n14171), .ZN(P1_U3547) );
  AOI211_X1 U16024 ( .C1(n14175), .C2(n14712), .A(n14174), .B(n14173), .ZN(
        n14176) );
  OAI211_X1 U16025 ( .C1(n14178), .C2(n14716), .A(n14177), .B(n14176), .ZN(
        n14229) );
  MUX2_X1 U16026 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14229), .S(n14734), .Z(
        P1_U3546) );
  OAI211_X1 U16027 ( .C1(n14181), .C2(n14587), .A(n14180), .B(n14179), .ZN(
        n14182) );
  AOI21_X1 U16028 ( .B1(n14184), .B2(n14183), .A(n14182), .ZN(n14185) );
  OAI21_X1 U16029 ( .B1(n14186), .B2(n14192), .A(n14185), .ZN(n14230) );
  MUX2_X1 U16030 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14230), .S(n14734), .Z(
        P1_U3545) );
  AOI21_X1 U16031 ( .B1(n14188), .B2(n14712), .A(n14187), .ZN(n14189) );
  OAI211_X1 U16032 ( .C1(n14192), .C2(n14191), .A(n14190), .B(n14189), .ZN(
        n14231) );
  MUX2_X1 U16033 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14231), .S(n14734), .Z(
        P1_U3544) );
  AOI21_X1 U16034 ( .B1(n14546), .B2(n14712), .A(n14193), .ZN(n14197) );
  NAND3_X1 U16035 ( .A1(n14195), .A2(n14194), .A3(n14725), .ZN(n14196) );
  NAND3_X1 U16036 ( .A1(n14198), .A2(n14197), .A3(n14196), .ZN(n14232) );
  MUX2_X1 U16037 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n14232), .S(n14734), .Z(
        P1_U3542) );
  MUX2_X1 U16038 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n14199), .S(n14734), .Z(
        P1_U3529) );
  MUX2_X1 U16039 ( .A(n14201), .B(n14200), .S(n14729), .Z(n14202) );
  OAI21_X1 U16040 ( .B1(n7236), .B2(n14227), .A(n14202), .ZN(P1_U3527) );
  MUX2_X1 U16041 ( .A(n14204), .B(n14203), .S(n14729), .Z(n14205) );
  OAI21_X1 U16042 ( .B1(n14206), .B2(n14227), .A(n14205), .ZN(P1_U3526) );
  MUX2_X1 U16043 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14208), .S(n14729), .Z(
        P1_U3524) );
  MUX2_X1 U16044 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14210), .S(n14729), .Z(
        P1_U3522) );
  MUX2_X1 U16045 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14211), .S(n14729), .Z(
        P1_U3521) );
  INV_X1 U16046 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n14213) );
  MUX2_X1 U16047 ( .A(n14213), .B(n14212), .S(n14729), .Z(n14214) );
  OAI21_X1 U16048 ( .B1(n11616), .B2(n14227), .A(n14214), .ZN(P1_U3520) );
  MUX2_X1 U16049 ( .A(n14215), .B(P1_REG0_REG_23__SCAN_IN), .S(n14727), .Z(
        P1_U3519) );
  INV_X1 U16050 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n14217) );
  MUX2_X1 U16051 ( .A(n14217), .B(n14216), .S(n14729), .Z(n14218) );
  OAI21_X1 U16052 ( .B1(n14227), .B2(n7363), .A(n14218), .ZN(P1_U3518) );
  MUX2_X1 U16053 ( .A(n14220), .B(n14219), .S(n14729), .Z(n14221) );
  OAI21_X1 U16054 ( .B1(n14222), .B2(n14227), .A(n14221), .ZN(P1_U3517) );
  MUX2_X1 U16055 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14223), .S(n14729), .Z(
        P1_U3516) );
  INV_X1 U16056 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14225) );
  MUX2_X1 U16057 ( .A(n14225), .B(n14224), .S(n14729), .Z(n14226) );
  OAI21_X1 U16058 ( .B1(n14228), .B2(n14227), .A(n14226), .ZN(P1_U3515) );
  MUX2_X1 U16059 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14229), .S(n14729), .Z(
        P1_U3513) );
  MUX2_X1 U16060 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14230), .S(n14729), .Z(
        P1_U3510) );
  MUX2_X1 U16061 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14231), .S(n14729), .Z(
        P1_U3507) );
  MUX2_X1 U16062 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n14232), .S(n14729), .Z(
        P1_U3501) );
  NAND3_X1 U16063 ( .A1(n14233), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n14235) );
  OAI22_X1 U16064 ( .A1(n14236), .A2(n14235), .B1(n14234), .B2(n14252), .ZN(
        n14237) );
  AOI21_X1 U16065 ( .B1(n14239), .B2(n14238), .A(n14237), .ZN(n14240) );
  INV_X1 U16066 ( .A(n14240), .ZN(P1_U3324) );
  INV_X1 U16067 ( .A(n11975), .ZN(n14241) );
  OAI222_X1 U16068 ( .A1(n14252), .A2(n14242), .B1(n10724), .B2(n14241), .C1(
        P1_U3086), .C2(n6468), .ZN(P1_U3327) );
  OAI222_X1 U16069 ( .A1(n14252), .A2(n7070), .B1(n10724), .B2(n14243), .C1(
        n14619), .C2(P1_U3086), .ZN(P1_U3328) );
  INV_X1 U16070 ( .A(n14244), .ZN(n14247) );
  OAI222_X1 U16071 ( .A1(n14247), .A2(P1_U3086), .B1(n10724), .B2(n14246), 
        .C1(n14245), .C2(n14252), .ZN(P1_U3329) );
  INV_X1 U16072 ( .A(n14248), .ZN(n14249) );
  OAI222_X1 U16073 ( .A1(n14252), .A2(n14251), .B1(n10724), .B2(n14250), .C1(
        n14249), .C2(P1_U3086), .ZN(P1_U3330) );
  MUX2_X1 U16074 ( .A(n14254), .B(n14253), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16075 ( .A(n14255), .ZN(n14256) );
  MUX2_X1 U16076 ( .A(n14256), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  XNOR2_X1 U16077 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(P3_ADDR_REG_15__SCAN_IN), 
        .ZN(n14292) );
  INV_X1 U16078 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n15039) );
  NOR2_X1 U16079 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(n15039), .ZN(n14291) );
  INV_X1 U16080 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14285) );
  INV_X1 U16081 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14281) );
  INV_X1 U16082 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14279) );
  XOR2_X1 U16083 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P3_ADDR_REG_2__SCAN_IN), .Z(
        n14297) );
  NOR2_X1 U16084 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(n14305), .ZN(n14262) );
  NOR2_X1 U16085 ( .A1(n14266), .A2(n14267), .ZN(n14269) );
  AND2_X1 U16086 ( .A1(n14270), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n14271) );
  NOR2_X1 U16087 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14272), .ZN(n14275) );
  XNOR2_X1 U16088 ( .A(P3_ADDR_REG_7__SCAN_IN), .B(n14272), .ZN(n14315) );
  INV_X1 U16089 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14273) );
  XNOR2_X1 U16090 ( .A(n14277), .B(P1_ADDR_REG_8__SCAN_IN), .ZN(n14293) );
  XNOR2_X1 U16091 ( .A(P3_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n14321) );
  NAND2_X1 U16092 ( .A1(n14322), .A2(n14321), .ZN(n14278) );
  NAND2_X1 U16093 ( .A1(n14281), .A2(n14280), .ZN(n14327) );
  NAND2_X1 U16094 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n14328), .ZN(n14282) );
  NAND2_X1 U16095 ( .A1(n14327), .A2(n14282), .ZN(n14332) );
  INV_X1 U16096 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14283) );
  NAND2_X1 U16097 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(n14283), .ZN(n14284) );
  XOR2_X1 U16098 ( .A(P3_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .Z(n14337) );
  INV_X1 U16099 ( .A(n14340), .ZN(n14289) );
  AND2_X1 U16100 ( .A1(n15017), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14288) );
  INV_X1 U16101 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14290) );
  OAI22_X1 U16102 ( .A1(n14291), .A2(n14345), .B1(P3_ADDR_REG_14__SCAN_IN), 
        .B2(n14290), .ZN(n14350) );
  XOR2_X1 U16103 ( .A(n14292), .B(n14350), .Z(n14347) );
  INV_X1 U16104 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14609) );
  XOR2_X1 U16105 ( .A(n14294), .B(n14293), .Z(n14320) );
  NAND2_X1 U16106 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14296), .ZN(n14307) );
  INV_X1 U16107 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14370) );
  XNOR2_X1 U16108 ( .A(n14298), .B(n14297), .ZN(n14368) );
  NAND2_X1 U16109 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14301), .ZN(n14303) );
  AOI21_X1 U16110 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14300), .A(n7137), .ZN(
        n15156) );
  INV_X1 U16111 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15155) );
  NOR2_X1 U16112 ( .A1(n15156), .A2(n15155), .ZN(n15164) );
  XOR2_X1 U16113 ( .A(n14301), .B(P2_ADDR_REG_1__SCAN_IN), .Z(n15163) );
  NAND2_X1 U16114 ( .A1(n15164), .A2(n15163), .ZN(n14302) );
  NAND2_X1 U16115 ( .A1(n14368), .A2(n14369), .ZN(n14304) );
  NOR2_X1 U16116 ( .A1(n14368), .A2(n14369), .ZN(n14367) );
  XNOR2_X1 U16117 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14305), .ZN(n15161) );
  NOR2_X1 U16118 ( .A1(n15160), .A2(n15161), .ZN(n14306) );
  INV_X1 U16119 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n14778) );
  NAND2_X1 U16120 ( .A1(n15160), .A2(n15161), .ZN(n15159) );
  XNOR2_X1 U16121 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14308), .ZN(n14309) );
  XNOR2_X1 U16122 ( .A(n14310), .B(n14309), .ZN(n15154) );
  NAND2_X1 U16123 ( .A1(n14311), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14314) );
  XNOR2_X1 U16124 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(P3_ADDR_REG_6__SCAN_IN), 
        .ZN(n14313) );
  XOR2_X1 U16125 ( .A(n14313), .B(n14312), .Z(n14372) );
  XNOR2_X1 U16126 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14315), .ZN(n15158) );
  NAND2_X1 U16127 ( .A1(n15157), .A2(n15158), .ZN(n14318) );
  NAND2_X1 U16128 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14316), .ZN(n14317) );
  XNOR2_X1 U16129 ( .A(n14322), .B(n14321), .ZN(n14324) );
  NAND2_X1 U16130 ( .A1(n14323), .A2(n14324), .ZN(n14326) );
  NAND2_X1 U16131 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n14380), .ZN(n14325) );
  NAND2_X1 U16132 ( .A1(n14328), .A2(n14327), .ZN(n14329) );
  XOR2_X1 U16133 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n14329), .Z(n14330) );
  XNOR2_X1 U16134 ( .A(P3_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n14333) );
  XOR2_X1 U16135 ( .A(n14333), .B(n14332), .Z(n14334) );
  XNOR2_X1 U16136 ( .A(n14338), .B(n14337), .ZN(n14599) );
  NAND2_X1 U16137 ( .A1(n14600), .A2(n14599), .ZN(n14339) );
  XNOR2_X1 U16138 ( .A(P3_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n14341) );
  XNOR2_X1 U16139 ( .A(n14341), .B(n14340), .ZN(n14342) );
  XNOR2_X1 U16140 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n14346) );
  XNOR2_X1 U16141 ( .A(n14346), .B(n14345), .ZN(n14608) );
  XNOR2_X1 U16142 ( .A(P1_ADDR_REG_16__SCAN_IN), .B(P3_ADDR_REG_16__SCAN_IN), 
        .ZN(n14352) );
  INV_X1 U16143 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n14646) );
  NOR2_X1 U16144 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n14646), .ZN(n14351) );
  INV_X1 U16145 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14416) );
  OAI22_X1 U16146 ( .A1(n14351), .A2(n14350), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14416), .ZN(n14355) );
  XOR2_X1 U16147 ( .A(n14352), .B(n14355), .Z(n14353) );
  INV_X1 U16148 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n14357) );
  INV_X1 U16149 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14431) );
  NOR2_X1 U16150 ( .A1(P1_ADDR_REG_16__SCAN_IN), .A2(n14431), .ZN(n14356) );
  OAI22_X1 U16151 ( .A1(P3_ADDR_REG_16__SCAN_IN), .A2(n14357), .B1(n14356), 
        .B2(n14355), .ZN(n14361) );
  XNOR2_X1 U16152 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n14361), .ZN(n14362) );
  XOR2_X1 U16153 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14362), .Z(n14359) );
  NOR2_X1 U16154 ( .A1(n14358), .A2(n14359), .ZN(n14393) );
  NOR2_X1 U16155 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n14361), .ZN(n14364) );
  INV_X1 U16156 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n14448) );
  NOR2_X1 U16157 ( .A1(n14448), .A2(n14362), .ZN(n14363) );
  NOR2_X1 U16158 ( .A1(n14364), .A2(n14363), .ZN(n14398) );
  XOR2_X1 U16159 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), 
        .Z(n14397) );
  XNOR2_X1 U16160 ( .A(n14398), .B(n14397), .ZN(n14396) );
  XNOR2_X1 U16161 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14395), .ZN(SUB_1596_U62)
         );
  AOI21_X1 U16162 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14365) );
  OAI21_X1 U16163 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14365), 
        .ZN(U28) );
  AOI21_X1 U16164 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(
        P3_RD_REG_SCAN_IN), .ZN(n14366) );
  OAI21_X1 U16165 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .A(n14366), 
        .ZN(U29) );
  AOI21_X1 U16166 ( .B1(n14369), .B2(n14368), .A(n14367), .ZN(n14371) );
  XNOR2_X1 U16167 ( .A(n14371), .B(n14370), .ZN(SUB_1596_U61) );
  XOR2_X1 U16168 ( .A(n14373), .B(n14372), .Z(SUB_1596_U57) );
  XNOR2_X1 U16169 ( .A(n14374), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  AOI22_X1 U16170 ( .A1(n14377), .A2(n14376), .B1(SI_18_), .B2(n14375), .ZN(
        n14378) );
  OAI21_X1 U16171 ( .B1(P3_U3151), .B2(n14379), .A(n14378), .ZN(P3_U3277) );
  XOR2_X1 U16172 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n14380), .Z(SUB_1596_U54) );
  XNOR2_X1 U16173 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14381), .ZN(SUB_1596_U70)
         );
  OAI21_X1 U16174 ( .B1(n14383), .B2(n14587), .A(n14382), .ZN(n14384) );
  AOI21_X1 U16175 ( .B1(n14386), .B2(n14385), .A(n14384), .ZN(n14387) );
  AND2_X1 U16176 ( .A1(n14388), .A2(n14387), .ZN(n14391) );
  INV_X1 U16177 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14389) );
  AOI22_X1 U16178 ( .A1(n14729), .A2(n14391), .B1(n14389), .B2(n14727), .ZN(
        P1_U3495) );
  AOI22_X1 U16179 ( .A1(n14734), .A2(n14391), .B1(n14390), .B2(n14732), .ZN(
        P1_U3540) );
  NOR2_X1 U16180 ( .A1(n14393), .A2(n14392), .ZN(n14394) );
  XOR2_X1 U16181 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14394), .Z(SUB_1596_U63)
         );
  NOR2_X1 U16182 ( .A1(n14398), .A2(n14397), .ZN(n14399) );
  AOI21_X1 U16183 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n13827), .A(n14399), 
        .ZN(n14403) );
  XNOR2_X1 U16184 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n14400) );
  XNOR2_X1 U16185 ( .A(n14401), .B(n14400), .ZN(n14402) );
  AOI21_X1 U16186 ( .B1(n14406), .B2(n14405), .A(n14404), .ZN(n14421) );
  OAI21_X1 U16187 ( .B1(n14408), .B2(P3_REG1_REG_15__SCAN_IN), .A(n14407), 
        .ZN(n14419) );
  INV_X1 U16188 ( .A(n15042), .ZN(n15005) );
  OAI21_X1 U16189 ( .B1(n14410), .B2(n14409), .A(n15005), .ZN(n14412) );
  NOR2_X1 U16190 ( .A1(n14412), .A2(n14411), .ZN(n14418) );
  INV_X1 U16191 ( .A(n14998), .ZN(n15038) );
  NAND2_X1 U16192 ( .A1(n15035), .A2(n14413), .ZN(n14415) );
  OAI211_X1 U16193 ( .C1(n14416), .C2(n15038), .A(n14415), .B(n14414), .ZN(
        n14417) );
  AOI211_X1 U16194 ( .C1(n14419), .C2(n15048), .A(n14418), .B(n14417), .ZN(
        n14420) );
  OAI21_X1 U16195 ( .B1(n14421), .B2(n15050), .A(n14420), .ZN(P3_U3197) );
  AOI21_X1 U16196 ( .B1(n14424), .B2(n14423), .A(n14422), .ZN(n14440) );
  OAI21_X1 U16197 ( .B1(n14427), .B2(n14426), .A(n14425), .ZN(n14438) );
  NAND2_X1 U16198 ( .A1(n15035), .A2(n14428), .ZN(n14430) );
  OAI211_X1 U16199 ( .C1(n14431), .C2(n15038), .A(n14430), .B(n14429), .ZN(
        n14437) );
  OR2_X1 U16200 ( .A1(n14433), .A2(n14432), .ZN(n14434) );
  AOI21_X1 U16201 ( .B1(n14435), .B2(n14434), .A(n15042), .ZN(n14436) );
  AOI211_X1 U16202 ( .C1(n15048), .C2(n14438), .A(n14437), .B(n14436), .ZN(
        n14439) );
  OAI21_X1 U16203 ( .B1(n14440), .B2(n15050), .A(n14439), .ZN(P3_U3198) );
  AOI21_X1 U16204 ( .B1(n14443), .B2(n14442), .A(n14441), .ZN(n14455) );
  XNOR2_X1 U16205 ( .A(n14444), .B(P3_REG1_REG_17__SCAN_IN), .ZN(n14445) );
  NAND2_X1 U16206 ( .A1(n15048), .A2(n14445), .ZN(n14446) );
  OAI211_X1 U16207 ( .C1(n15038), .C2(n14448), .A(n14447), .B(n14446), .ZN(
        n14453) );
  AOI211_X1 U16208 ( .C1(n14451), .C2(n14450), .A(n15042), .B(n14449), .ZN(
        n14452) );
  AOI211_X1 U16209 ( .C1(n15035), .C2(n6698), .A(n14453), .B(n14452), .ZN(
        n14454) );
  OAI21_X1 U16210 ( .B1(n14455), .B2(n15050), .A(n14454), .ZN(P3_U3199) );
  INV_X1 U16211 ( .A(n14456), .ZN(n14457) );
  AOI22_X1 U16212 ( .A1(n14459), .A2(n15098), .B1(n14469), .B2(n15120), .ZN(
        n14464) );
  AOI22_X1 U16213 ( .A1(n14460), .A2(n15081), .B1(n14462), .B2(
        P3_REG2_REG_31__SCAN_IN), .ZN(n14461) );
  NAND2_X1 U16214 ( .A1(n14464), .A2(n14461), .ZN(P3_U3202) );
  AOI22_X1 U16215 ( .A1(n14470), .A2(n15081), .B1(P3_REG2_REG_30__SCAN_IN), 
        .B2(n14462), .ZN(n14463) );
  NAND2_X1 U16216 ( .A1(n14464), .A2(n14463), .ZN(P3_U3203) );
  OR2_X1 U16217 ( .A1(n14465), .A2(n15138), .ZN(n14467) );
  INV_X1 U16218 ( .A(n14469), .ZN(n14466) );
  AOI22_X1 U16219 ( .A1(n15149), .A2(n14486), .B1(n14468), .B2(n15150), .ZN(
        P3_U3490) );
  AOI21_X1 U16220 ( .B1(n14470), .B2(n14476), .A(n14469), .ZN(n14487) );
  AOI22_X1 U16221 ( .A1(n15149), .A2(n14487), .B1(n14471), .B2(n15150), .ZN(
        P3_U3489) );
  NOR2_X1 U16222 ( .A1(n14472), .A2(n15139), .ZN(n14474) );
  AOI211_X1 U16223 ( .C1(n14476), .C2(n14475), .A(n14474), .B(n14473), .ZN(
        n14488) );
  AOI22_X1 U16224 ( .A1(n15149), .A2(n14488), .B1(n8489), .B2(n15150), .ZN(
        P3_U3472) );
  NOR2_X1 U16225 ( .A1(n14477), .A2(n15138), .ZN(n14479) );
  AOI211_X1 U16226 ( .C1(n14482), .C2(n14480), .A(n14479), .B(n14478), .ZN(
        n14489) );
  AOI22_X1 U16227 ( .A1(n15149), .A2(n14489), .B1(n8461), .B2(n15150), .ZN(
        P3_U3471) );
  AOI21_X1 U16228 ( .B1(n14483), .B2(n14482), .A(n14481), .ZN(n14484) );
  AND2_X1 U16229 ( .A1(n14485), .A2(n14484), .ZN(n14490) );
  AOI22_X1 U16230 ( .A1(n15149), .A2(n14490), .B1(n8439), .B2(n15150), .ZN(
        P3_U3470) );
  AOI22_X1 U16231 ( .A1(n15144), .A2(n11654), .B1(n14486), .B2(n15143), .ZN(
        P3_U3458) );
  AOI22_X1 U16232 ( .A1(n15144), .A2(n8722), .B1(n14487), .B2(n15143), .ZN(
        P3_U3457) );
  AOI22_X1 U16233 ( .A1(n15144), .A2(n8494), .B1(n14488), .B2(n15143), .ZN(
        P3_U3429) );
  AOI22_X1 U16234 ( .A1(n15144), .A2(n8464), .B1(n14489), .B2(n15143), .ZN(
        P3_U3426) );
  AOI22_X1 U16235 ( .A1(n15144), .A2(n8442), .B1(n14490), .B2(n15143), .ZN(
        P3_U3423) );
  OAI21_X1 U16236 ( .B1(n14493), .B2(n14492), .A(n14491), .ZN(n14495) );
  AOI222_X1 U16237 ( .A1(n14499), .A2(n14498), .B1(n14497), .B2(n14496), .C1(
        n14495), .C2(n14494), .ZN(n14501) );
  OAI211_X1 U16238 ( .C1(n14503), .C2(n14502), .A(n14501), .B(n14500), .ZN(
        P2_U3187) );
  XNOR2_X1 U16239 ( .A(n14504), .B(n14508), .ZN(n14530) );
  OAI211_X1 U16240 ( .C1(n14527), .C2(n6606), .A(n14816), .B(n14505), .ZN(
        n14526) );
  INV_X1 U16241 ( .A(n14526), .ZN(n14506) );
  AOI22_X1 U16242 ( .A1(n14530), .A2(n14828), .B1(n14507), .B2(n14506), .ZN(
        n14517) );
  XOR2_X1 U16243 ( .A(n14509), .B(n14508), .Z(n14511) );
  OAI21_X1 U16244 ( .B1(n14511), .B2(n14834), .A(n14510), .ZN(n14528) );
  AOI22_X1 U16245 ( .A1(n14844), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n14512), 
        .B2(n14839), .ZN(n14513) );
  OAI21_X1 U16246 ( .B1(n14527), .B2(n14824), .A(n14513), .ZN(n14514) );
  AOI21_X1 U16247 ( .B1(n14528), .B2(n14515), .A(n14514), .ZN(n14516) );
  NAND2_X1 U16248 ( .A1(n14517), .A2(n14516), .ZN(P2_U3253) );
  INV_X1 U16249 ( .A(n14518), .ZN(n14519) );
  OAI21_X1 U16250 ( .B1(n14520), .B2(n14933), .A(n14519), .ZN(n14523) );
  INV_X1 U16251 ( .A(n14521), .ZN(n14522) );
  AOI211_X1 U16252 ( .C1(n14913), .C2(n14524), .A(n14523), .B(n14522), .ZN(
        n14533) );
  AOI22_X1 U16253 ( .A1(n14970), .A2(n14533), .B1(n14525), .B2(n14968), .ZN(
        P2_U3513) );
  OAI21_X1 U16254 ( .B1(n14527), .B2(n14933), .A(n14526), .ZN(n14529) );
  AOI211_X1 U16255 ( .C1(n14913), .C2(n14530), .A(n14529), .B(n14528), .ZN(
        n14535) );
  AOI22_X1 U16256 ( .A1(n14970), .A2(n14535), .B1(n14531), .B2(n14968), .ZN(
        P2_U3511) );
  INV_X1 U16257 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14532) );
  AOI22_X1 U16258 ( .A1(n14952), .A2(n14533), .B1(n14532), .B2(n14950), .ZN(
        P2_U3472) );
  INV_X1 U16259 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14534) );
  AOI22_X1 U16260 ( .A1(n14952), .A2(n14535), .B1(n14534), .B2(n14950), .ZN(
        P2_U3466) );
  OAI22_X1 U16261 ( .A1(n14565), .A2(n14537), .B1(n14536), .B2(n14562), .ZN(
        n14545) );
  AOI21_X1 U16262 ( .B1(n14540), .B2(n14539), .A(n14538), .ZN(n14541) );
  INV_X1 U16263 ( .A(n14541), .ZN(n14543) );
  AOI21_X1 U16264 ( .B1(n14543), .B2(n14542), .A(n14570), .ZN(n14544) );
  AOI211_X1 U16265 ( .C1(n14576), .C2(n14546), .A(n14545), .B(n14544), .ZN(
        n14548) );
  OAI211_X1 U16266 ( .C1(n14580), .C2(n14549), .A(n14548), .B(n14547), .ZN(
        P1_U3215) );
  OAI22_X1 U16267 ( .A1(n14552), .A2(n14551), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14550), .ZN(n14558) );
  OAI211_X1 U16268 ( .C1(n14555), .C2(n14554), .A(n14568), .B(n14553), .ZN(
        n14556) );
  INV_X1 U16269 ( .A(n14556), .ZN(n14557) );
  AOI211_X1 U16270 ( .C1(n14576), .C2(n14559), .A(n14558), .B(n14557), .ZN(
        n14560) );
  OAI21_X1 U16271 ( .B1(n14561), .B2(n14580), .A(n14560), .ZN(P1_U3217) );
  OAI22_X1 U16272 ( .A1(n14565), .A2(n14564), .B1(n14563), .B2(n14562), .ZN(
        n14574) );
  AOI21_X1 U16273 ( .B1(n14568), .B2(n14567), .A(n14566), .ZN(n14569) );
  INV_X1 U16274 ( .A(n14569), .ZN(n14572) );
  AOI21_X1 U16275 ( .B1(n14572), .B2(n14571), .A(n14570), .ZN(n14573) );
  AOI211_X1 U16276 ( .C1(n14576), .C2(n14575), .A(n14574), .B(n14573), .ZN(
        n14578) );
  OAI211_X1 U16277 ( .C1(n14580), .C2(n14579), .A(n14578), .B(n14577), .ZN(
        P1_U3236) );
  OAI21_X1 U16278 ( .B1(n14582), .B2(n14587), .A(n14581), .ZN(n14584) );
  AOI211_X1 U16279 ( .C1(n14585), .C2(n14725), .A(n14584), .B(n14583), .ZN(
        n14593) );
  AOI22_X1 U16280 ( .A1(n14734), .A2(n14593), .B1(n10940), .B2(n14732), .ZN(
        P1_U3541) );
  OAI21_X1 U16281 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(n14590) );
  AOI211_X1 U16282 ( .C1(n14591), .C2(n14725), .A(n14590), .B(n14589), .ZN(
        n14595) );
  AOI22_X1 U16283 ( .A1(n14734), .A2(n14595), .B1(n10830), .B2(n14732), .ZN(
        P1_U3539) );
  INV_X1 U16284 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14592) );
  AOI22_X1 U16285 ( .A1(n14729), .A2(n14593), .B1(n14592), .B2(n14727), .ZN(
        P1_U3498) );
  INV_X1 U16286 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n14594) );
  AOI22_X1 U16287 ( .A1(n14729), .A2(n14595), .B1(n14594), .B2(n14727), .ZN(
        P1_U3492) );
  XOR2_X1 U16288 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(n14597), .Z(SUB_1596_U69)
         );
  AOI21_X1 U16289 ( .B1(n14600), .B2(n14599), .A(n14598), .ZN(n14602) );
  XNOR2_X1 U16290 ( .A(n14602), .B(n14601), .ZN(SUB_1596_U68) );
  NOR2_X1 U16291 ( .A1(n14604), .A2(n14603), .ZN(n14605) );
  XOR2_X1 U16292 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(n14605), .Z(SUB_1596_U67)
         );
  AOI21_X1 U16293 ( .B1(n14608), .B2(n14607), .A(n14606), .ZN(n14610) );
  XNOR2_X1 U16294 ( .A(n14610), .B(n14609), .ZN(SUB_1596_U66) );
  NOR2_X1 U16295 ( .A1(n14612), .A2(n14611), .ZN(n14613) );
  XOR2_X1 U16296 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n14613), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16297 ( .A1(n14615), .A2(n14614), .ZN(n14616) );
  XOR2_X1 U16298 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(n14616), .Z(SUB_1596_U64)
         );
  INV_X1 U16299 ( .A(n14617), .ZN(n14620) );
  NAND2_X1 U16300 ( .A1(n14619), .A2(n14618), .ZN(n14622) );
  NAND2_X1 U16301 ( .A1(n14620), .A2(n14622), .ZN(n14623) );
  MUX2_X1 U16302 ( .A(n14623), .B(n14622), .S(n14621), .Z(n14625) );
  NAND2_X1 U16303 ( .A1(n14625), .A2(n14624), .ZN(n14629) );
  AOI22_X1 U16304 ( .A1(n14627), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n14628) );
  OAI21_X1 U16305 ( .B1(n14630), .B2(n14629), .A(n14628), .ZN(P1_U3243) );
  AOI21_X1 U16306 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n14632), .A(n14631), 
        .ZN(n14633) );
  INV_X1 U16307 ( .A(n14633), .ZN(n14642) );
  OAI21_X1 U16308 ( .B1(n14636), .B2(n14635), .A(n14634), .ZN(n14639) );
  AOI222_X1 U16309 ( .A1(n14642), .A2(n14641), .B1(n14640), .B2(n14639), .C1(
        n14638), .C2(n14637), .ZN(n14644) );
  OAI211_X1 U16310 ( .C1(n14646), .C2(n14645), .A(n14644), .B(n14643), .ZN(
        P1_U3258) );
  NAND2_X1 U16311 ( .A1(n14647), .A2(n14659), .ZN(n14652) );
  INV_X1 U16312 ( .A(n14648), .ZN(n14649) );
  AOI22_X1 U16313 ( .A1(n14650), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n14649), 
        .B2(n14662), .ZN(n14651) );
  OAI211_X1 U16314 ( .C1(n14653), .C2(n14666), .A(n14652), .B(n14651), .ZN(
        n14654) );
  AOI21_X1 U16315 ( .B1(n14656), .B2(n14655), .A(n14654), .ZN(n14657) );
  OAI21_X1 U16316 ( .B1(n14673), .B2(n14658), .A(n14657), .ZN(P1_U3285) );
  NAND2_X1 U16317 ( .A1(n14660), .A2(n14659), .ZN(n14665) );
  INV_X1 U16318 ( .A(n14661), .ZN(n14663) );
  AOI22_X1 U16319 ( .A1(n14673), .A2(P1_REG2_REG_6__SCAN_IN), .B1(n14663), 
        .B2(n14662), .ZN(n14664) );
  OAI211_X1 U16320 ( .C1(n14667), .C2(n14666), .A(n14665), .B(n14664), .ZN(
        n14668) );
  AOI21_X1 U16321 ( .B1(n14670), .B2(n14669), .A(n14668), .ZN(n14671) );
  OAI21_X1 U16322 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(P1_U3287) );
  NOR2_X1 U16323 ( .A1(n14704), .A2(n14674), .ZN(P1_U3294) );
  INV_X1 U16324 ( .A(P1_D_REG_30__SCAN_IN), .ZN(n14675) );
  NOR2_X1 U16325 ( .A1(n14704), .A2(n14675), .ZN(P1_U3295) );
  INV_X1 U16326 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n14676) );
  NOR2_X1 U16327 ( .A1(n14704), .A2(n14676), .ZN(P1_U3296) );
  INV_X1 U16328 ( .A(P1_D_REG_28__SCAN_IN), .ZN(n14677) );
  NOR2_X1 U16329 ( .A1(n14704), .A2(n14677), .ZN(P1_U3297) );
  INV_X1 U16330 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n14678) );
  NOR2_X1 U16331 ( .A1(n14704), .A2(n14678), .ZN(P1_U3298) );
  INV_X1 U16332 ( .A(P1_D_REG_26__SCAN_IN), .ZN(n14679) );
  NOR2_X1 U16333 ( .A1(n14704), .A2(n14679), .ZN(P1_U3299) );
  NOR2_X1 U16334 ( .A1(n14704), .A2(n14680), .ZN(P1_U3300) );
  NOR2_X1 U16335 ( .A1(n14704), .A2(n14681), .ZN(P1_U3301) );
  INV_X1 U16336 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n14682) );
  NOR2_X1 U16337 ( .A1(n14704), .A2(n14682), .ZN(P1_U3302) );
  INV_X1 U16338 ( .A(P1_D_REG_22__SCAN_IN), .ZN(n14683) );
  NOR2_X1 U16339 ( .A1(n14704), .A2(n14683), .ZN(P1_U3303) );
  INV_X1 U16340 ( .A(P1_D_REG_21__SCAN_IN), .ZN(n14684) );
  NOR2_X1 U16341 ( .A1(n14704), .A2(n14684), .ZN(P1_U3304) );
  INV_X1 U16342 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n14685) );
  NOR2_X1 U16343 ( .A1(n14704), .A2(n14685), .ZN(P1_U3305) );
  INV_X1 U16344 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n14686) );
  NOR2_X1 U16345 ( .A1(n14704), .A2(n14686), .ZN(P1_U3306) );
  INV_X1 U16346 ( .A(P1_D_REG_18__SCAN_IN), .ZN(n14687) );
  NOR2_X1 U16347 ( .A1(n14704), .A2(n14687), .ZN(P1_U3307) );
  INV_X1 U16348 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n14688) );
  NOR2_X1 U16349 ( .A1(n14704), .A2(n14688), .ZN(P1_U3308) );
  INV_X1 U16350 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n14689) );
  NOR2_X1 U16351 ( .A1(n14704), .A2(n14689), .ZN(P1_U3309) );
  INV_X1 U16352 ( .A(P1_D_REG_15__SCAN_IN), .ZN(n14690) );
  NOR2_X1 U16353 ( .A1(n14704), .A2(n14690), .ZN(P1_U3310) );
  INV_X1 U16354 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n14691) );
  NOR2_X1 U16355 ( .A1(n14704), .A2(n14691), .ZN(P1_U3311) );
  INV_X1 U16356 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n14692) );
  NOR2_X1 U16357 ( .A1(n14704), .A2(n14692), .ZN(P1_U3312) );
  INV_X1 U16358 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n14693) );
  NOR2_X1 U16359 ( .A1(n14704), .A2(n14693), .ZN(P1_U3313) );
  INV_X1 U16360 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n14694) );
  NOR2_X1 U16361 ( .A1(n14704), .A2(n14694), .ZN(P1_U3314) );
  NOR2_X1 U16362 ( .A1(n14704), .A2(n14695), .ZN(P1_U3315) );
  INV_X1 U16363 ( .A(P1_D_REG_9__SCAN_IN), .ZN(n14696) );
  NOR2_X1 U16364 ( .A1(n14704), .A2(n14696), .ZN(P1_U3316) );
  INV_X1 U16365 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n14697) );
  NOR2_X1 U16366 ( .A1(n14704), .A2(n14697), .ZN(P1_U3317) );
  INV_X1 U16367 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n14698) );
  NOR2_X1 U16368 ( .A1(n14704), .A2(n14698), .ZN(P1_U3318) );
  INV_X1 U16369 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n14699) );
  NOR2_X1 U16370 ( .A1(n14704), .A2(n14699), .ZN(P1_U3319) );
  INV_X1 U16371 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n14700) );
  NOR2_X1 U16372 ( .A1(n14704), .A2(n14700), .ZN(P1_U3320) );
  INV_X1 U16373 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n14701) );
  NOR2_X1 U16374 ( .A1(n14704), .A2(n14701), .ZN(P1_U3321) );
  INV_X1 U16375 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n14702) );
  NOR2_X1 U16376 ( .A1(n14704), .A2(n14702), .ZN(P1_U3322) );
  INV_X1 U16377 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n14703) );
  NOR2_X1 U16378 ( .A1(n14704), .A2(n14703), .ZN(P1_U3323) );
  AOI21_X1 U16379 ( .B1(n14706), .B2(n14712), .A(n14705), .ZN(n14707) );
  OAI211_X1 U16380 ( .C1(n14709), .C2(n14716), .A(n14708), .B(n14707), .ZN(
        n14710) );
  INV_X1 U16381 ( .A(n14710), .ZN(n14730) );
  AOI22_X1 U16382 ( .A1(n14729), .A2(n14730), .B1(n9476), .B2(n14727), .ZN(
        P1_U3468) );
  AOI21_X1 U16383 ( .B1(n14713), .B2(n14712), .A(n14711), .ZN(n14714) );
  OAI211_X1 U16384 ( .C1(n14717), .C2(n14716), .A(n14715), .B(n14714), .ZN(
        n14718) );
  INV_X1 U16385 ( .A(n14718), .ZN(n14731) );
  INV_X1 U16386 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14719) );
  AOI22_X1 U16387 ( .A1(n14729), .A2(n14731), .B1(n14719), .B2(n14727), .ZN(
        P1_U3474) );
  NAND3_X1 U16388 ( .A1(n14722), .A2(n14721), .A3(n14720), .ZN(n14724) );
  AOI211_X1 U16389 ( .C1(n14726), .C2(n14725), .A(n14724), .B(n14723), .ZN(
        n14733) );
  INV_X1 U16390 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14728) );
  AOI22_X1 U16391 ( .A1(n14729), .A2(n14733), .B1(n14728), .B2(n14727), .ZN(
        P1_U3486) );
  AOI22_X1 U16392 ( .A1(n14734), .A2(n14730), .B1(n9302), .B2(n14732), .ZN(
        P1_U3531) );
  AOI22_X1 U16393 ( .A1(n14734), .A2(n14731), .B1(n9857), .B2(n14732), .ZN(
        P1_U3533) );
  AOI22_X1 U16394 ( .A1(n14734), .A2(n14733), .B1(n10498), .B2(n14732), .ZN(
        P1_U3537) );
  NOR2_X1 U16395 ( .A1(n14799), .A2(P2_U3947), .ZN(P2_U3087) );
  AOI22_X1 U16396 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n14800), .B1(n14765), 
        .B2(P2_REG1_REG_0__SCAN_IN), .ZN(n14738) );
  AOI22_X1 U16397 ( .A1(n14799), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3088), .ZN(n14737) );
  OAI22_X1 U16398 ( .A1(n14795), .A2(P2_REG1_REG_0__SCAN_IN), .B1(
        P2_REG2_REG_0__SCAN_IN), .B2(n14786), .ZN(n14735) );
  OAI21_X1 U16399 ( .B1(n14805), .B2(n14735), .A(n14739), .ZN(n14736) );
  OAI211_X1 U16400 ( .C1(n14739), .C2(n14738), .A(n14737), .B(n14736), .ZN(
        P2_U3214) );
  AOI22_X1 U16401 ( .A1(n14799), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3088), .ZN(n14750) );
  XNOR2_X1 U16402 ( .A(n14741), .B(n14740), .ZN(n14743) );
  AOI22_X1 U16403 ( .A1(n14765), .A2(n14743), .B1(n14742), .B2(n14805), .ZN(
        n14749) );
  AOI211_X1 U16404 ( .C1(n14746), .C2(n14745), .A(n14744), .B(n14786), .ZN(
        n14747) );
  INV_X1 U16405 ( .A(n14747), .ZN(n14748) );
  NAND3_X1 U16406 ( .A1(n14750), .A2(n14749), .A3(n14748), .ZN(P2_U3215) );
  AOI22_X1 U16407 ( .A1(n14799), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3088), .ZN(n14762) );
  OAI21_X1 U16408 ( .B1(n14753), .B2(n14752), .A(n14751), .ZN(n14754) );
  INV_X1 U16409 ( .A(n14754), .ZN(n14756) );
  AOI22_X1 U16410 ( .A1(n14765), .A2(n14756), .B1(n14755), .B2(n14805), .ZN(
        n14761) );
  XOR2_X1 U16411 ( .A(n14758), .B(n14757), .Z(n14759) );
  NAND2_X1 U16412 ( .A1(n14800), .A2(n14759), .ZN(n14760) );
  NAND3_X1 U16413 ( .A1(n14762), .A2(n14761), .A3(n14760), .ZN(P2_U3216) );
  INV_X1 U16414 ( .A(n14763), .ZN(n14764) );
  OAI211_X1 U16415 ( .C1(n14767), .C2(n14766), .A(n14765), .B(n14764), .ZN(
        n14772) );
  INV_X1 U16416 ( .A(n14768), .ZN(n14769) );
  AOI21_X1 U16417 ( .B1(n14805), .B2(n14770), .A(n14769), .ZN(n14771) );
  AND2_X1 U16418 ( .A1(n14772), .A2(n14771), .ZN(n14777) );
  OAI211_X1 U16419 ( .C1(n14775), .C2(n14774), .A(n14800), .B(n14773), .ZN(
        n14776) );
  OAI211_X1 U16420 ( .C1(n14793), .C2(n14778), .A(n14777), .B(n14776), .ZN(
        P2_U3217) );
  NOR2_X1 U16421 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n14779), .ZN(n14784) );
  AOI211_X1 U16422 ( .C1(n14782), .C2(n14781), .A(n14795), .B(n14780), .ZN(
        n14783) );
  AOI211_X1 U16423 ( .C1(n14805), .C2(n14785), .A(n14784), .B(n14783), .ZN(
        n14792) );
  AOI21_X1 U16424 ( .B1(n14788), .B2(n14787), .A(n14786), .ZN(n14790) );
  NAND2_X1 U16425 ( .A1(n14790), .A2(n14789), .ZN(n14791) );
  OAI211_X1 U16426 ( .C1(n14793), .C2(n7140), .A(n14792), .B(n14791), .ZN(
        P2_U3221) );
  AOI211_X1 U16427 ( .C1(n14797), .C2(n14796), .A(n14795), .B(n14794), .ZN(
        n14798) );
  AOI21_X1 U16428 ( .B1(n14799), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n14798), 
        .ZN(n14809) );
  OAI211_X1 U16429 ( .C1(n14803), .C2(n14802), .A(n14801), .B(n14800), .ZN(
        n14807) );
  NAND2_X1 U16430 ( .A1(n14805), .A2(n14804), .ZN(n14806) );
  NAND4_X1 U16431 ( .A1(n14809), .A2(n14808), .A3(n14807), .A4(n14806), .ZN(
        P2_U3231) );
  XNOR2_X1 U16432 ( .A(n14811), .B(n14810), .ZN(n14815) );
  INV_X1 U16433 ( .A(n14812), .ZN(n14813) );
  AOI21_X1 U16434 ( .B1(n14815), .B2(n14814), .A(n14813), .ZN(n14880) );
  OAI211_X1 U16435 ( .C1(n14818), .C2(n14879), .A(n14817), .B(n14816), .ZN(
        n14878) );
  OAI22_X1 U16436 ( .A1(n14820), .A2(n14878), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14819), .ZN(n14821) );
  INV_X1 U16437 ( .A(n14821), .ZN(n14823) );
  NAND2_X1 U16438 ( .A1(n14844), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n14822) );
  OAI211_X1 U16439 ( .C1(n14824), .C2(n14879), .A(n14823), .B(n14822), .ZN(
        n14825) );
  INV_X1 U16440 ( .A(n14825), .ZN(n14830) );
  XNOR2_X1 U16441 ( .A(n14827), .B(n14826), .ZN(n14883) );
  NAND2_X1 U16442 ( .A1(n14828), .A2(n14883), .ZN(n14829) );
  OAI211_X1 U16443 ( .C1(n14844), .C2(n14880), .A(n14830), .B(n14829), .ZN(
        P2_U3262) );
  AOI21_X1 U16444 ( .B1(n14833), .B2(n14832), .A(n14831), .ZN(n14838) );
  NAND2_X1 U16445 ( .A1(n6660), .A2(n14834), .ZN(n14836) );
  AOI21_X1 U16446 ( .B1(n14858), .B2(n14836), .A(n14835), .ZN(n14860) );
  INV_X1 U16447 ( .A(n14860), .ZN(n14837) );
  AOI211_X1 U16448 ( .C1(n14839), .C2(P2_REG3_REG_0__SCAN_IN), .A(n14838), .B(
        n14837), .ZN(n14843) );
  INV_X1 U16449 ( .A(n14840), .ZN(n14841) );
  AOI22_X1 U16450 ( .A1(n14841), .A2(n14858), .B1(P2_REG2_REG_0__SCAN_IN), 
        .B2(n14844), .ZN(n14842) );
  OAI21_X1 U16451 ( .B1(n14844), .B2(n14843), .A(n14842), .ZN(P2_U3265) );
  NOR2_X1 U16452 ( .A1(n14851), .A2(n14845), .ZN(n14848) );
  AND2_X1 U16453 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14846), .ZN(P2_U3266) );
  AND2_X1 U16454 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14846), .ZN(P2_U3267) );
  AND2_X1 U16455 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14846), .ZN(P2_U3268) );
  AND2_X1 U16456 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14846), .ZN(P2_U3269) );
  AND2_X1 U16457 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14846), .ZN(P2_U3270) );
  AND2_X1 U16458 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14846), .ZN(P2_U3271) );
  AND2_X1 U16459 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14846), .ZN(P2_U3272) );
  AND2_X1 U16460 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14846), .ZN(P2_U3273) );
  AND2_X1 U16461 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14846), .ZN(P2_U3274) );
  AND2_X1 U16462 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14846), .ZN(P2_U3275) );
  AND2_X1 U16463 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14846), .ZN(P2_U3276) );
  AND2_X1 U16464 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14846), .ZN(P2_U3277) );
  AND2_X1 U16465 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14846), .ZN(P2_U3278) );
  AND2_X1 U16466 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14846), .ZN(P2_U3279) );
  AND2_X1 U16467 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14846), .ZN(P2_U3280) );
  AND2_X1 U16468 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14846), .ZN(P2_U3281) );
  AND2_X1 U16469 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14846), .ZN(P2_U3282) );
  AND2_X1 U16470 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14846), .ZN(P2_U3283) );
  AND2_X1 U16471 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14846), .ZN(P2_U3284) );
  AND2_X1 U16472 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14846), .ZN(P2_U3285) );
  AND2_X1 U16473 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14846), .ZN(P2_U3286) );
  AND2_X1 U16474 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14846), .ZN(P2_U3287) );
  AND2_X1 U16475 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14846), .ZN(P2_U3288) );
  AND2_X1 U16476 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14846), .ZN(P2_U3289) );
  AND2_X1 U16477 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14846), .ZN(P2_U3290) );
  AND2_X1 U16478 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14846), .ZN(P2_U3291) );
  AND2_X1 U16479 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14846), .ZN(P2_U3292) );
  AND2_X1 U16480 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14846), .ZN(P2_U3293) );
  AND2_X1 U16481 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14846), .ZN(P2_U3294) );
  NOR2_X1 U16482 ( .A1(n14848), .A2(n14847), .ZN(P2_U3295) );
  AOI22_X1 U16483 ( .A1(n14854), .A2(n14850), .B1(n14849), .B2(n14851), .ZN(
        P2_U3416) );
  AOI22_X1 U16484 ( .A1(n14854), .A2(n14853), .B1(n14852), .B2(n14851), .ZN(
        P2_U3417) );
  AOI22_X1 U16485 ( .A1(n14858), .A2(n14857), .B1(n14856), .B2(n14855), .ZN(
        n14859) );
  AND2_X1 U16486 ( .A1(n14860), .A2(n14859), .ZN(n14954) );
  INV_X1 U16487 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14861) );
  AOI22_X1 U16488 ( .A1(n14952), .A2(n14954), .B1(n14861), .B2(n14950), .ZN(
        P2_U3430) );
  INV_X1 U16489 ( .A(n14862), .ZN(n14868) );
  INV_X1 U16490 ( .A(n6660), .ZN(n14949) );
  NOR2_X1 U16491 ( .A1(n14862), .A2(n14945), .ZN(n14867) );
  OAI211_X1 U16492 ( .C1(n14865), .C2(n14933), .A(n14864), .B(n14863), .ZN(
        n14866) );
  AOI211_X1 U16493 ( .C1(n14868), .C2(n14949), .A(n14867), .B(n14866), .ZN(
        n14956) );
  INV_X1 U16494 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14869) );
  AOI22_X1 U16495 ( .A1(n14952), .A2(n14956), .B1(n14869), .B2(n14950), .ZN(
        P2_U3433) );
  INV_X1 U16496 ( .A(n14876), .ZN(n14872) );
  AOI21_X1 U16497 ( .B1(n14943), .B2(n8937), .A(n14870), .ZN(n14871) );
  OAI21_X1 U16498 ( .B1(n14872), .B2(n14945), .A(n14871), .ZN(n14875) );
  INV_X1 U16499 ( .A(n14873), .ZN(n14874) );
  AOI211_X1 U16500 ( .C1(n14949), .C2(n14876), .A(n14875), .B(n14874), .ZN(
        n14957) );
  INV_X1 U16501 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14877) );
  AOI22_X1 U16502 ( .A1(n14952), .A2(n14957), .B1(n14877), .B2(n14950), .ZN(
        P2_U3436) );
  OAI21_X1 U16503 ( .B1(n14879), .B2(n14933), .A(n14878), .ZN(n14882) );
  INV_X1 U16504 ( .A(n14880), .ZN(n14881) );
  AOI211_X1 U16505 ( .C1(n14883), .C2(n14913), .A(n14882), .B(n14881), .ZN(
        n14958) );
  INV_X1 U16506 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U16507 ( .A1(n14952), .A2(n14958), .B1(n14884), .B2(n14950), .ZN(
        P2_U3439) );
  OAI211_X1 U16508 ( .C1(n14887), .C2(n14933), .A(n14886), .B(n14885), .ZN(
        n14890) );
  AOI21_X1 U16509 ( .B1(n6660), .B2(n14945), .A(n14888), .ZN(n14889) );
  NOR2_X1 U16510 ( .A1(n14890), .A2(n14889), .ZN(n14960) );
  INV_X1 U16511 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14891) );
  AOI22_X1 U16512 ( .A1(n14952), .A2(n14960), .B1(n14891), .B2(n14950), .ZN(
        P2_U3442) );
  INV_X1 U16513 ( .A(n14892), .ZN(n14893) );
  OAI211_X1 U16514 ( .C1(n14895), .C2(n14933), .A(n14894), .B(n14893), .ZN(
        n14898) );
  AOI21_X1 U16515 ( .B1(n6660), .B2(n14945), .A(n14896), .ZN(n14897) );
  NOR2_X1 U16516 ( .A1(n14898), .A2(n14897), .ZN(n14962) );
  INV_X1 U16517 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U16518 ( .A1(n14952), .A2(n14962), .B1(n14899), .B2(n14950), .ZN(
        P2_U3445) );
  INV_X1 U16519 ( .A(n14904), .ZN(n14906) );
  AOI21_X1 U16520 ( .B1(n14943), .B2(n14901), .A(n14900), .ZN(n14903) );
  OAI211_X1 U16521 ( .C1(n14945), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        n14905) );
  AOI21_X1 U16522 ( .B1(n14949), .B2(n14906), .A(n14905), .ZN(n14963) );
  INV_X1 U16523 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n14907) );
  AOI22_X1 U16524 ( .A1(n14952), .A2(n14963), .B1(n14907), .B2(n14950), .ZN(
        P2_U3448) );
  OAI21_X1 U16525 ( .B1(n14909), .B2(n14933), .A(n14908), .ZN(n14911) );
  AOI211_X1 U16526 ( .C1(n14913), .C2(n14912), .A(n14911), .B(n14910), .ZN(
        n14964) );
  INV_X1 U16527 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n14914) );
  AOI22_X1 U16528 ( .A1(n14952), .A2(n14964), .B1(n14914), .B2(n14950), .ZN(
        P2_U3451) );
  INV_X1 U16529 ( .A(n14918), .ZN(n14921) );
  AOI21_X1 U16530 ( .B1(n14943), .B2(n14916), .A(n14915), .ZN(n14917) );
  OAI21_X1 U16531 ( .B1(n14945), .B2(n14918), .A(n14917), .ZN(n14919) );
  AOI211_X1 U16532 ( .C1(n14949), .C2(n14921), .A(n14920), .B(n14919), .ZN(
        n14965) );
  INV_X1 U16533 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14922) );
  AOI22_X1 U16534 ( .A1(n14952), .A2(n14965), .B1(n14922), .B2(n14950), .ZN(
        P2_U3454) );
  OR2_X1 U16535 ( .A1(n14923), .A2(n14933), .ZN(n14924) );
  OAI211_X1 U16536 ( .C1(n14926), .C2(n14945), .A(n14925), .B(n14924), .ZN(
        n14929) );
  NOR2_X1 U16537 ( .A1(n14926), .A2(n6660), .ZN(n14927) );
  NOR3_X1 U16538 ( .A1(n14929), .A2(n14928), .A3(n14927), .ZN(n14966) );
  INV_X1 U16539 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n14930) );
  AOI22_X1 U16540 ( .A1(n14952), .A2(n14966), .B1(n14930), .B2(n14950), .ZN(
        P2_U3457) );
  OAI211_X1 U16541 ( .C1(n14934), .C2(n14933), .A(n14932), .B(n14931), .ZN(
        n14938) );
  AOI21_X1 U16542 ( .B1(n6660), .B2(n14945), .A(n14935), .ZN(n14937) );
  NOR2_X1 U16543 ( .A1(n14938), .A2(n14937), .ZN(n14967) );
  INV_X1 U16544 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14939) );
  AOI22_X1 U16545 ( .A1(n14952), .A2(n14967), .B1(n14939), .B2(n14950), .ZN(
        P2_U3460) );
  INV_X1 U16546 ( .A(n14946), .ZN(n14948) );
  AOI211_X1 U16547 ( .C1(n14943), .C2(n14942), .A(n14941), .B(n14940), .ZN(
        n14944) );
  OAI21_X1 U16548 ( .B1(n14946), .B2(n14945), .A(n14944), .ZN(n14947) );
  AOI21_X1 U16549 ( .B1(n14949), .B2(n14948), .A(n14947), .ZN(n14969) );
  INV_X1 U16550 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n14951) );
  AOI22_X1 U16551 ( .A1(n14952), .A2(n14969), .B1(n14951), .B2(n14950), .ZN(
        P2_U3463) );
  INV_X1 U16552 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14953) );
  AOI22_X1 U16553 ( .A1(n14970), .A2(n14954), .B1(n14953), .B2(n14968), .ZN(
        P2_U3499) );
  INV_X1 U16554 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n14955) );
  AOI22_X1 U16555 ( .A1(n14970), .A2(n14956), .B1(n14955), .B2(n14968), .ZN(
        P2_U3500) );
  AOI22_X1 U16556 ( .A1(n14970), .A2(n14957), .B1(n9370), .B2(n14968), .ZN(
        P2_U3501) );
  AOI22_X1 U16557 ( .A1(n14970), .A2(n14958), .B1(n6840), .B2(n14968), .ZN(
        P2_U3502) );
  INV_X1 U16558 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U16559 ( .A1(n14970), .A2(n14960), .B1(n14959), .B2(n14968), .ZN(
        P2_U3503) );
  INV_X1 U16560 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U16561 ( .A1(n14970), .A2(n14962), .B1(n14961), .B2(n14968), .ZN(
        P2_U3504) );
  AOI22_X1 U16562 ( .A1(n14970), .A2(n14963), .B1(n9376), .B2(n14968), .ZN(
        P2_U3505) );
  AOI22_X1 U16563 ( .A1(n14970), .A2(n14964), .B1(n9556), .B2(n14968), .ZN(
        P2_U3506) );
  AOI22_X1 U16564 ( .A1(n14970), .A2(n14965), .B1(n9557), .B2(n14968), .ZN(
        P2_U3507) );
  AOI22_X1 U16565 ( .A1(n14970), .A2(n14966), .B1(n9585), .B2(n14968), .ZN(
        P2_U3508) );
  AOI22_X1 U16566 ( .A1(n14970), .A2(n14967), .B1(n9794), .B2(n14968), .ZN(
        P2_U3509) );
  AOI22_X1 U16567 ( .A1(n14970), .A2(n14969), .B1(n10138), .B2(n14968), .ZN(
        P2_U3510) );
  NOR2_X1 U16568 ( .A1(P3_U3897), .A2(n14998), .ZN(P3_U3150) );
  AOI21_X1 U16569 ( .B1(n14973), .B2(n14972), .A(n14971), .ZN(n14986) );
  XNOR2_X1 U16570 ( .A(n14975), .B(n14974), .ZN(n14984) );
  OAI21_X1 U16571 ( .B1(n14977), .B2(P3_REG1_REG_11__SCAN_IN), .A(n14976), 
        .ZN(n14978) );
  NAND2_X1 U16572 ( .A1(n14978), .A2(n15048), .ZN(n14981) );
  AOI21_X1 U16573 ( .B1(n14998), .B2(P3_ADDR_REG_11__SCAN_IN), .A(n14979), 
        .ZN(n14980) );
  OAI211_X1 U16574 ( .C1(n15002), .C2(n14982), .A(n14981), .B(n14980), .ZN(
        n14983) );
  AOI21_X1 U16575 ( .B1(n15005), .B2(n14984), .A(n14983), .ZN(n14985) );
  OAI21_X1 U16576 ( .B1(n14986), .B2(n15050), .A(n14985), .ZN(P3_U3193) );
  INV_X1 U16577 ( .A(n14987), .ZN(n14988) );
  AOI21_X1 U16578 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n15007) );
  XOR2_X1 U16579 ( .A(n14992), .B(n14991), .Z(n15004) );
  OAI21_X1 U16580 ( .B1(n14995), .B2(n14994), .A(n14993), .ZN(n14996) );
  NAND2_X1 U16581 ( .A1(n14996), .A2(n15048), .ZN(n15000) );
  AOI21_X1 U16582 ( .B1(n14998), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n14997), 
        .ZN(n14999) );
  OAI211_X1 U16583 ( .C1(n15002), .C2(n15001), .A(n15000), .B(n14999), .ZN(
        n15003) );
  AOI21_X1 U16584 ( .B1(n15005), .B2(n15004), .A(n15003), .ZN(n15006) );
  OAI21_X1 U16585 ( .B1(n15007), .B2(n15050), .A(n15006), .ZN(P3_U3194) );
  AOI21_X1 U16586 ( .B1(n15010), .B2(n15009), .A(n15008), .ZN(n15026) );
  OAI21_X1 U16587 ( .B1(n15012), .B2(P3_REG1_REG_13__SCAN_IN), .A(n15011), 
        .ZN(n15013) );
  NAND2_X1 U16588 ( .A1(n15048), .A2(n15013), .ZN(n15016) );
  INV_X1 U16589 ( .A(n15014), .ZN(n15015) );
  OAI211_X1 U16590 ( .C1(n15038), .C2(n15017), .A(n15016), .B(n15015), .ZN(
        n15023) );
  NAND2_X1 U16591 ( .A1(n15019), .A2(n15018), .ZN(n15020) );
  AOI21_X1 U16592 ( .B1(n15021), .B2(n15020), .A(n15042), .ZN(n15022) );
  AOI211_X1 U16593 ( .C1(n15035), .C2(n15024), .A(n15023), .B(n15022), .ZN(
        n15025) );
  OAI21_X1 U16594 ( .B1(n15026), .B2(n15050), .A(n15025), .ZN(P3_U3195) );
  AOI21_X1 U16595 ( .B1(n15029), .B2(n15028), .A(n15027), .ZN(n15051) );
  OAI21_X1 U16596 ( .B1(n15032), .B2(n15031), .A(n15030), .ZN(n15047) );
  INV_X1 U16597 ( .A(n15033), .ZN(n15034) );
  NAND2_X1 U16598 ( .A1(n15035), .A2(n15034), .ZN(n15037) );
  OAI211_X1 U16599 ( .C1(n15039), .C2(n15038), .A(n15037), .B(n15036), .ZN(
        n15046) );
  INV_X1 U16600 ( .A(n15040), .ZN(n15041) );
  AOI211_X1 U16601 ( .C1(n15044), .C2(n15043), .A(n15042), .B(n15041), .ZN(
        n15045) );
  AOI211_X1 U16602 ( .C1(n15048), .C2(n15047), .A(n15046), .B(n15045), .ZN(
        n15049) );
  OAI21_X1 U16603 ( .B1(n15051), .B2(n15050), .A(n15049), .ZN(P3_U3196) );
  NAND2_X1 U16604 ( .A1(n15056), .A2(n15090), .ZN(n15052) );
  OAI211_X1 U16605 ( .C1(n15054), .C2(n15114), .A(n15053), .B(n15052), .ZN(
        n15058) );
  INV_X1 U16606 ( .A(n15116), .ZN(n15055) );
  AOI222_X1 U16607 ( .A1(n15058), .A2(n15120), .B1(n15081), .B2(n15057), .C1(
        n15056), .C2(n15055), .ZN(n15059) );
  OAI21_X1 U16608 ( .B1(n15120), .B2(n15060), .A(n15059), .ZN(P3_U3226) );
  NOR2_X1 U16609 ( .A1(n15090), .A2(n15095), .ZN(n15076) );
  OAI21_X1 U16610 ( .B1(n15062), .B2(n15076), .A(n15061), .ZN(n15063) );
  MUX2_X1 U16611 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n15063), .S(n15120), .Z(
        n15064) );
  AOI21_X1 U16612 ( .B1(n15081), .B2(n15065), .A(n15064), .ZN(n15066) );
  OAI21_X1 U16613 ( .B1(n15067), .B2(n15114), .A(n15066), .ZN(P3_U3227) );
  OAI21_X1 U16614 ( .B1(n15076), .B2(n15069), .A(n15068), .ZN(n15070) );
  MUX2_X1 U16615 ( .A(P3_REG2_REG_5__SCAN_IN), .B(n15070), .S(n15120), .Z(
        n15071) );
  AOI21_X1 U16616 ( .B1(n15081), .B2(n15072), .A(n15071), .ZN(n15073) );
  OAI21_X1 U16617 ( .B1(n15074), .B2(n15114), .A(n15073), .ZN(P3_U3228) );
  OAI21_X1 U16618 ( .B1(n15077), .B2(n15076), .A(n15075), .ZN(n15078) );
  MUX2_X1 U16619 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n15078), .S(n15120), .Z(
        n15079) );
  AOI21_X1 U16620 ( .B1(n15081), .B2(n15080), .A(n15079), .ZN(n15082) );
  OAI21_X1 U16621 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15114), .A(n15082), .ZN(
        P3_U3230) );
  XNOR2_X1 U16622 ( .A(n15083), .B(n15085), .ZN(n15092) );
  OAI21_X1 U16623 ( .B1(n15086), .B2(n15085), .A(n15084), .ZN(n15128) );
  OAI22_X1 U16624 ( .A1(n15088), .A2(n15106), .B1(n15087), .B2(n15104), .ZN(
        n15089) );
  AOI21_X1 U16625 ( .B1(n15128), .B2(n15090), .A(n15089), .ZN(n15091) );
  OAI21_X1 U16626 ( .B1(n15093), .B2(n15092), .A(n15091), .ZN(n15126) );
  NOR2_X1 U16627 ( .A1(n15094), .A2(n15138), .ZN(n15127) );
  AOI22_X1 U16628 ( .A1(n15128), .A2(n15095), .B1(n15127), .B2(n15113), .ZN(
        n15096) );
  INV_X1 U16629 ( .A(n15096), .ZN(n15097) );
  AOI211_X1 U16630 ( .C1(P3_REG3_REG_2__SCAN_IN), .C2(n15098), .A(n15126), .B(
        n15097), .ZN(n15099) );
  AOI22_X1 U16631 ( .A1(n14462), .A2(n7017), .B1(n15099), .B2(n15120), .ZN(
        P3_U3231) );
  NOR2_X1 U16632 ( .A1(n15100), .A2(n15138), .ZN(n15124) );
  XNOR2_X1 U16633 ( .A(n15102), .B(n15101), .ZN(n15122) );
  XNOR2_X1 U16634 ( .A(n15103), .B(n15102), .ZN(n15110) );
  OAI22_X1 U16635 ( .A1(n15107), .A2(n15106), .B1(n6670), .B2(n15104), .ZN(
        n15108) );
  AOI21_X1 U16636 ( .B1(n15110), .B2(n15109), .A(n15108), .ZN(n15111) );
  OAI21_X1 U16637 ( .B1(n15122), .B2(n15112), .A(n15111), .ZN(n15123) );
  AOI21_X1 U16638 ( .B1(n15124), .B2(n15113), .A(n15123), .ZN(n15121) );
  OAI22_X1 U16639 ( .A1(n15122), .A2(n15116), .B1(n15115), .B2(n15114), .ZN(
        n15117) );
  INV_X1 U16640 ( .A(n15117), .ZN(n15118) );
  OAI221_X1 U16641 ( .B1(n14462), .B2(n15121), .C1(n15120), .C2(n15119), .A(
        n15118), .ZN(P3_U3232) );
  INV_X1 U16642 ( .A(n15122), .ZN(n15125) );
  AOI211_X1 U16643 ( .C1(n6605), .C2(n15125), .A(n15124), .B(n15123), .ZN(
        n15145) );
  AOI22_X1 U16644 ( .A1(n15144), .A2(n8268), .B1(n15145), .B2(n15143), .ZN(
        P3_U3393) );
  AOI211_X1 U16645 ( .C1(n6605), .C2(n15128), .A(n15127), .B(n15126), .ZN(
        n15146) );
  AOI22_X1 U16646 ( .A1(n15144), .A2(n8288), .B1(n15146), .B2(n15143), .ZN(
        P3_U3396) );
  INV_X1 U16647 ( .A(n15129), .ZN(n15132) );
  AOI211_X1 U16648 ( .C1(n15132), .C2(n6605), .A(n15131), .B(n15130), .ZN(
        n15147) );
  AOI22_X1 U16649 ( .A1(n15144), .A2(n8390), .B1(n15147), .B2(n15143), .ZN(
        P3_U3414) );
  INV_X1 U16650 ( .A(n15133), .ZN(n15136) );
  AOI211_X1 U16651 ( .C1(n15136), .C2(n6605), .A(n15135), .B(n15134), .ZN(
        n15148) );
  AOI22_X1 U16652 ( .A1(n15144), .A2(n8423), .B1(n15148), .B2(n15143), .ZN(
        P3_U3417) );
  OAI22_X1 U16653 ( .A1(n15140), .A2(n15139), .B1(n15138), .B2(n15137), .ZN(
        n15141) );
  NOR2_X1 U16654 ( .A1(n15142), .A2(n15141), .ZN(n15151) );
  AOI22_X1 U16655 ( .A1(n15144), .A2(n8406), .B1(n15151), .B2(n15143), .ZN(
        P3_U3420) );
  AOI22_X1 U16656 ( .A1(n15149), .A2(n15145), .B1(n8270), .B2(n15150), .ZN(
        P3_U3460) );
  AOI22_X1 U16657 ( .A1(n15149), .A2(n15146), .B1(n9998), .B2(n15150), .ZN(
        P3_U3461) );
  AOI22_X1 U16658 ( .A1(n15149), .A2(n15147), .B1(n10391), .B2(n15150), .ZN(
        P3_U3467) );
  AOI22_X1 U16659 ( .A1(n15149), .A2(n15148), .B1(n8418), .B2(n15150), .ZN(
        P3_U3468) );
  AOI22_X1 U16660 ( .A1(n15149), .A2(n15151), .B1(n8404), .B2(n15150), .ZN(
        P3_U3469) );
  XOR2_X1 U16661 ( .A(n15153), .B(n15152), .Z(SUB_1596_U59) );
  XNOR2_X1 U16662 ( .A(n15154), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16663 ( .B1(n15156), .B2(n15155), .A(n15164), .ZN(SUB_1596_U53) );
  XOR2_X1 U16664 ( .A(n15157), .B(n15158), .Z(SUB_1596_U56) );
  OAI21_X1 U16665 ( .B1(n15161), .B2(n15160), .A(n15159), .ZN(n15162) );
  XNOR2_X1 U16666 ( .A(n15162), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  XOR2_X1 U16667 ( .A(n15164), .B(n15163), .Z(SUB_1596_U5) );
  NAND2_X1 U7199 ( .A1(n12041), .A2(n8880), .ZN(n8883) );
  CLKBUF_X1 U7209 ( .A(n6799), .Z(n6716) );
  CLKBUF_X1 U7282 ( .A(n13053), .Z(n12976) );
  CLKBUF_X1 U7322 ( .A(n12096), .Z(n6459) );
  CLKBUF_X1 U7500 ( .A(n10067), .Z(n6431) );
  CLKBUF_X1 U7514 ( .A(n9299), .Z(n6468) );
endmodule

